module basic_2500_25000_3000_125_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_754,In_2257);
nor U1 (N_1,In_1966,In_820);
or U2 (N_2,In_1248,In_73);
or U3 (N_3,In_551,In_2184);
and U4 (N_4,In_636,In_2409);
nand U5 (N_5,In_2248,In_1171);
or U6 (N_6,In_1894,In_331);
or U7 (N_7,In_589,In_1558);
or U8 (N_8,In_350,In_1132);
nor U9 (N_9,In_1193,In_1586);
and U10 (N_10,In_1616,In_498);
or U11 (N_11,In_373,In_144);
or U12 (N_12,In_109,In_1825);
and U13 (N_13,In_2352,In_598);
xor U14 (N_14,In_2094,In_2066);
nor U15 (N_15,In_1094,In_83);
or U16 (N_16,In_943,In_1339);
nor U17 (N_17,In_1938,In_337);
nor U18 (N_18,In_207,In_945);
and U19 (N_19,In_2366,In_789);
and U20 (N_20,In_1968,In_352);
and U21 (N_21,In_524,In_2395);
and U22 (N_22,In_874,In_2107);
nand U23 (N_23,In_986,In_2357);
nand U24 (N_24,In_1170,In_2010);
xnor U25 (N_25,In_2057,In_1503);
nand U26 (N_26,In_1597,In_607);
nor U27 (N_27,In_2283,In_784);
and U28 (N_28,In_2070,In_1533);
and U29 (N_29,In_128,In_1362);
xor U30 (N_30,In_965,In_1693);
nor U31 (N_31,In_984,In_1200);
nor U32 (N_32,In_1054,In_2408);
xor U33 (N_33,In_653,In_948);
xnor U34 (N_34,In_329,In_1677);
nand U35 (N_35,In_2271,In_673);
or U36 (N_36,In_2358,In_1239);
nand U37 (N_37,In_427,In_1466);
nor U38 (N_38,In_2492,In_2085);
nand U39 (N_39,In_2499,In_177);
nor U40 (N_40,In_970,In_343);
nand U41 (N_41,In_918,In_2290);
xnor U42 (N_42,In_2118,In_442);
nor U43 (N_43,In_962,In_1761);
nor U44 (N_44,In_601,In_1845);
nand U45 (N_45,In_1246,In_573);
xnor U46 (N_46,In_2313,In_333);
nor U47 (N_47,In_492,In_1521);
nand U48 (N_48,In_1844,In_1264);
and U49 (N_49,In_595,In_1915);
xnor U50 (N_50,In_2125,In_1724);
or U51 (N_51,In_2008,In_591);
or U52 (N_52,In_2398,In_783);
xnor U53 (N_53,In_707,In_1875);
or U54 (N_54,In_1456,In_1582);
or U55 (N_55,In_2065,In_283);
nor U56 (N_56,In_2350,In_748);
or U57 (N_57,In_96,In_2123);
or U58 (N_58,In_338,In_868);
nand U59 (N_59,In_1139,In_1596);
nor U60 (N_60,In_2335,In_1668);
xnor U61 (N_61,In_2200,In_2153);
nor U62 (N_62,In_712,In_2073);
nand U63 (N_63,In_1283,In_856);
nand U64 (N_64,In_1797,In_1721);
and U65 (N_65,In_2055,In_628);
and U66 (N_66,In_2204,In_664);
nand U67 (N_67,In_2056,In_1899);
nor U68 (N_68,In_1182,In_1853);
and U69 (N_69,In_980,In_2176);
nand U70 (N_70,In_2451,In_930);
nand U71 (N_71,In_98,In_2212);
nor U72 (N_72,In_20,In_830);
and U73 (N_73,In_2020,In_1663);
xor U74 (N_74,In_290,In_2081);
nor U75 (N_75,In_582,In_219);
xor U76 (N_76,In_80,In_94);
nand U77 (N_77,In_2159,In_1902);
nor U78 (N_78,In_1700,In_1891);
nand U79 (N_79,In_471,In_2);
and U80 (N_80,In_1572,In_2321);
nand U81 (N_81,In_2237,In_1169);
or U82 (N_82,In_781,In_1397);
nor U83 (N_83,In_2463,In_1324);
or U84 (N_84,In_1612,In_158);
or U85 (N_85,In_1838,In_1227);
nand U86 (N_86,In_964,In_579);
or U87 (N_87,In_114,In_662);
and U88 (N_88,In_1382,In_1123);
xnor U89 (N_89,In_280,In_1261);
nand U90 (N_90,In_1114,In_835);
nor U91 (N_91,In_1862,In_1633);
nor U92 (N_92,In_1790,In_2496);
and U93 (N_93,In_2019,In_1282);
nor U94 (N_94,In_1457,In_996);
nor U95 (N_95,In_950,In_2268);
nand U96 (N_96,In_496,In_1980);
nand U97 (N_97,In_1958,In_592);
and U98 (N_98,In_1818,In_1629);
nand U99 (N_99,In_2025,In_1743);
xor U100 (N_100,In_143,In_2236);
and U101 (N_101,In_2038,In_1719);
nand U102 (N_102,In_729,In_1691);
nand U103 (N_103,In_1144,In_2262);
xnor U104 (N_104,In_2249,In_49);
xnor U105 (N_105,In_787,In_695);
xor U106 (N_106,In_43,In_2115);
xnor U107 (N_107,In_818,In_1356);
nand U108 (N_108,In_1623,In_328);
or U109 (N_109,In_275,In_927);
nand U110 (N_110,In_1064,In_1660);
xor U111 (N_111,In_1373,In_2468);
or U112 (N_112,In_1219,In_1051);
nand U113 (N_113,In_77,In_661);
or U114 (N_114,In_201,In_1926);
nand U115 (N_115,In_525,In_453);
nor U116 (N_116,In_2027,In_1849);
nand U117 (N_117,In_1177,In_2003);
nand U118 (N_118,In_2060,In_78);
and U119 (N_119,In_249,In_1537);
nand U120 (N_120,In_1292,In_507);
xor U121 (N_121,In_2349,In_1213);
nor U122 (N_122,In_238,In_1727);
nand U123 (N_123,In_2242,In_995);
xnor U124 (N_124,In_1065,In_1712);
or U125 (N_125,In_125,In_1179);
xnor U126 (N_126,In_111,In_1272);
and U127 (N_127,In_91,In_2480);
and U128 (N_128,In_2071,In_155);
nor U129 (N_129,In_2145,In_888);
nand U130 (N_130,In_1458,In_1506);
xnor U131 (N_131,In_1391,In_260);
nand U132 (N_132,In_1780,In_647);
and U133 (N_133,In_923,In_750);
xnor U134 (N_134,In_827,In_1214);
or U135 (N_135,In_1728,In_2078);
nand U136 (N_136,In_1085,In_2269);
or U137 (N_137,In_968,In_1355);
xnor U138 (N_138,In_680,In_1698);
nor U139 (N_139,In_1449,In_195);
nand U140 (N_140,In_1855,In_2014);
nor U141 (N_141,In_604,In_1565);
and U142 (N_142,In_1771,In_771);
nand U143 (N_143,In_705,In_1194);
or U144 (N_144,In_693,In_1235);
nor U145 (N_145,In_51,In_1764);
nor U146 (N_146,In_747,In_1119);
nor U147 (N_147,In_2407,In_2138);
and U148 (N_148,In_1999,In_1071);
nor U149 (N_149,In_222,In_741);
and U150 (N_150,In_132,In_1871);
nor U151 (N_151,In_1931,In_1316);
or U152 (N_152,In_2253,In_30);
nor U153 (N_153,In_718,In_2338);
nand U154 (N_154,In_1075,In_2183);
and U155 (N_155,In_1184,In_1856);
nor U156 (N_156,In_1108,In_2347);
and U157 (N_157,In_226,In_1619);
and U158 (N_158,In_515,In_1545);
or U159 (N_159,In_2105,In_668);
nand U160 (N_160,In_2109,In_1019);
or U161 (N_161,In_278,In_1437);
xnor U162 (N_162,In_404,In_845);
and U163 (N_163,In_1920,In_2354);
or U164 (N_164,In_677,In_1645);
and U165 (N_165,In_1387,In_742);
xor U166 (N_166,In_1304,In_1695);
and U167 (N_167,In_2007,In_183);
and U168 (N_168,In_833,In_149);
nand U169 (N_169,In_616,In_460);
and U170 (N_170,In_1777,In_1905);
nand U171 (N_171,In_1514,In_0);
nand U172 (N_172,In_434,In_457);
and U173 (N_173,In_2053,In_999);
and U174 (N_174,In_184,In_603);
and U175 (N_175,In_436,In_2309);
nand U176 (N_176,In_708,In_920);
nand U177 (N_177,In_1009,In_1671);
nor U178 (N_178,In_1823,In_1626);
xor U179 (N_179,In_1981,In_489);
nor U180 (N_180,In_236,In_1890);
xnor U181 (N_181,In_2048,In_2432);
or U182 (N_182,In_869,In_397);
nor U183 (N_183,In_983,In_90);
nor U184 (N_184,In_2288,In_2491);
nor U185 (N_185,In_549,In_926);
xnor U186 (N_186,In_1518,In_1187);
and U187 (N_187,In_1255,In_1694);
and U188 (N_188,In_288,In_2440);
nor U189 (N_189,In_1794,In_2293);
nor U190 (N_190,In_1296,In_2023);
and U191 (N_191,In_946,In_521);
nand U192 (N_192,In_1000,In_666);
nor U193 (N_193,In_97,In_1010);
nor U194 (N_194,In_1384,In_2052);
nand U195 (N_195,In_656,In_1882);
nand U196 (N_196,In_1953,In_1269);
and U197 (N_197,In_2382,In_1333);
xnor U198 (N_198,In_561,In_368);
and U199 (N_199,In_1829,In_187);
xor U200 (N_200,In_1175,In_1640);
and U201 (N_201,N_128,In_1606);
or U202 (N_202,In_1934,N_124);
xnor U203 (N_203,In_1886,N_46);
and U204 (N_204,In_2301,In_44);
and U205 (N_205,In_1903,In_199);
xnor U206 (N_206,In_2442,In_258);
and U207 (N_207,In_1786,In_1135);
xor U208 (N_208,In_2474,In_1842);
and U209 (N_209,In_1464,In_998);
nand U210 (N_210,In_769,In_1454);
xor U211 (N_211,In_394,In_810);
and U212 (N_212,In_859,N_170);
or U213 (N_213,N_85,In_1013);
and U214 (N_214,In_84,In_430);
or U215 (N_215,In_2475,In_2150);
and U216 (N_216,In_752,N_132);
xnor U217 (N_217,In_475,In_554);
nand U218 (N_218,In_213,In_1375);
xnor U219 (N_219,In_1158,N_5);
nor U220 (N_220,In_295,In_2119);
nor U221 (N_221,In_1232,In_1215);
nand U222 (N_222,In_776,In_755);
nand U223 (N_223,In_2190,In_68);
and U224 (N_224,In_804,In_1634);
nand U225 (N_225,In_847,In_606);
nor U226 (N_226,In_2416,N_15);
nand U227 (N_227,In_354,In_1793);
xnor U228 (N_228,In_889,In_1447);
nand U229 (N_229,In_1628,In_911);
and U230 (N_230,In_1992,In_391);
or U231 (N_231,In_2343,In_1785);
and U232 (N_232,In_216,In_1952);
nand U233 (N_233,In_1080,In_1116);
and U234 (N_234,In_468,In_107);
and U235 (N_235,In_1753,N_99);
or U236 (N_236,In_233,In_2163);
nand U237 (N_237,In_1491,In_1684);
nor U238 (N_238,In_944,In_2302);
nand U239 (N_239,In_958,In_1486);
nor U240 (N_240,In_857,In_2396);
and U241 (N_241,In_2033,In_1432);
nor U242 (N_242,N_149,In_1987);
nand U243 (N_243,In_1035,In_1913);
and U244 (N_244,In_1982,In_1773);
or U245 (N_245,In_2389,In_2273);
or U246 (N_246,In_1138,In_987);
or U247 (N_247,In_1142,In_1251);
nor U248 (N_248,In_1168,In_2486);
nand U249 (N_249,In_2223,In_753);
nor U250 (N_250,In_1395,In_1352);
nor U251 (N_251,In_854,In_376);
xnor U252 (N_252,N_148,In_1320);
and U253 (N_253,In_1118,N_104);
or U254 (N_254,In_1993,In_568);
nor U255 (N_255,In_2326,In_1186);
nor U256 (N_256,In_905,In_1834);
or U257 (N_257,In_1335,In_1520);
nand U258 (N_258,In_1502,In_198);
or U259 (N_259,In_1176,In_72);
xor U260 (N_260,In_370,N_125);
or U261 (N_261,In_735,In_1050);
and U262 (N_262,In_511,In_822);
nand U263 (N_263,In_1476,In_2462);
and U264 (N_264,In_1008,In_1630);
nand U265 (N_265,In_2376,In_1268);
nor U266 (N_266,In_2069,In_1347);
or U267 (N_267,In_168,In_1801);
and U268 (N_268,In_732,In_1331);
xor U269 (N_269,N_198,In_2334);
or U270 (N_270,N_137,In_1429);
nor U271 (N_271,In_982,In_1505);
xor U272 (N_272,In_1133,In_955);
nand U273 (N_273,In_581,In_1519);
and U274 (N_274,In_1542,In_50);
xnor U275 (N_275,In_744,In_396);
or U276 (N_276,In_2022,In_139);
and U277 (N_277,In_1178,N_109);
or U278 (N_278,N_4,In_766);
nand U279 (N_279,In_1569,In_1746);
or U280 (N_280,In_2128,In_466);
nor U281 (N_281,In_2386,In_600);
or U282 (N_282,In_2096,In_2256);
nand U283 (N_283,In_402,In_642);
xnor U284 (N_284,In_702,In_1877);
or U285 (N_285,In_1206,In_472);
or U286 (N_286,In_2045,In_440);
nand U287 (N_287,In_1809,In_54);
xor U288 (N_288,In_1972,In_452);
nand U289 (N_289,In_1602,In_1686);
nor U290 (N_290,In_1702,In_349);
and U291 (N_291,In_4,In_2191);
xnor U292 (N_292,In_1318,In_1897);
nand U293 (N_293,In_1989,In_407);
xnor U294 (N_294,In_2192,In_1441);
and U295 (N_295,N_184,In_1109);
xor U296 (N_296,In_767,In_174);
nand U297 (N_297,N_86,In_2099);
and U298 (N_298,In_1880,In_1427);
nor U299 (N_299,In_38,In_1576);
nand U300 (N_300,In_1067,In_2490);
and U301 (N_301,In_2446,In_649);
xor U302 (N_302,In_1620,In_814);
and U303 (N_303,In_898,In_863);
or U304 (N_304,In_10,In_1507);
and U305 (N_305,In_1613,In_1252);
or U306 (N_306,In_2220,In_2210);
xnor U307 (N_307,In_2077,In_2009);
nand U308 (N_308,In_1016,In_170);
nand U309 (N_309,In_1566,In_1799);
nand U310 (N_310,In_1388,In_850);
or U311 (N_311,In_861,In_978);
xnor U312 (N_312,In_2478,In_1847);
xnor U313 (N_313,In_610,In_1480);
nor U314 (N_314,In_190,In_411);
and U315 (N_315,In_575,In_266);
xor U316 (N_316,N_160,In_2281);
or U317 (N_317,In_795,In_1245);
or U318 (N_318,In_1368,In_1639);
nor U319 (N_319,In_1122,In_2238);
or U320 (N_320,In_1253,In_172);
or U321 (N_321,In_1631,In_8);
or U322 (N_322,In_2298,In_864);
nor U323 (N_323,In_508,In_1775);
nor U324 (N_324,In_1942,In_2084);
nand U325 (N_325,In_2195,In_819);
xor U326 (N_326,In_517,In_660);
xor U327 (N_327,In_2461,In_941);
nor U328 (N_328,In_2227,In_2092);
nor U329 (N_329,In_388,In_2420);
or U330 (N_330,In_178,In_1190);
and U331 (N_331,In_706,In_1153);
or U332 (N_332,In_2481,In_1759);
nor U333 (N_333,In_866,In_2103);
nor U334 (N_334,In_185,In_640);
xnor U335 (N_335,In_104,In_1451);
nor U336 (N_336,N_49,In_2181);
and U337 (N_337,In_1812,In_65);
nor U338 (N_338,In_157,In_896);
or U339 (N_339,In_2277,In_336);
nor U340 (N_340,In_1311,In_1172);
xor U341 (N_341,In_788,N_93);
nand U342 (N_342,In_234,In_126);
nor U343 (N_343,In_1070,N_120);
nand U344 (N_344,In_270,In_2245);
xnor U345 (N_345,In_1300,In_273);
nor U346 (N_346,In_638,In_317);
xnor U347 (N_347,In_782,In_227);
and U348 (N_348,In_1327,In_448);
nand U349 (N_349,In_1813,N_169);
or U350 (N_350,In_1497,In_1196);
or U351 (N_351,In_1511,In_1939);
and U352 (N_352,In_1509,In_1056);
nand U353 (N_353,N_45,In_537);
nand U354 (N_354,In_1974,In_1651);
xor U355 (N_355,In_1740,In_2209);
or U356 (N_356,In_2470,In_1342);
nor U357 (N_357,In_86,In_532);
nand U358 (N_358,In_1162,In_1650);
nor U359 (N_359,In_2344,In_123);
or U360 (N_360,In_1529,In_812);
and U361 (N_361,In_110,In_1157);
nand U362 (N_362,In_1076,In_657);
nand U363 (N_363,In_900,In_775);
xnor U364 (N_364,In_221,N_191);
nor U365 (N_365,In_1031,In_1416);
or U366 (N_366,In_1493,In_467);
or U367 (N_367,In_2439,In_1111);
or U368 (N_368,In_159,In_1510);
nand U369 (N_369,In_2211,In_1156);
xor U370 (N_370,In_75,In_2421);
nand U371 (N_371,In_1413,N_155);
nand U372 (N_372,In_1453,In_2434);
nand U373 (N_373,In_1303,In_1512);
nor U374 (N_374,In_464,In_1199);
nand U375 (N_375,In_1917,N_185);
xnor U376 (N_376,In_973,N_144);
or U377 (N_377,In_1032,N_139);
or U378 (N_378,In_2263,In_2401);
xnor U379 (N_379,In_1816,In_1925);
xnor U380 (N_380,In_659,In_180);
or U381 (N_381,In_230,In_264);
or U382 (N_382,In_1101,In_1066);
nand U383 (N_383,In_1083,N_145);
and U384 (N_384,In_1238,In_1997);
nand U385 (N_385,In_2013,In_2189);
nor U386 (N_386,In_1549,In_1647);
nor U387 (N_387,In_154,In_1749);
or U388 (N_388,In_2050,In_921);
nor U389 (N_389,In_1125,In_762);
nor U390 (N_390,In_257,In_1185);
nor U391 (N_391,In_2095,In_263);
nor U392 (N_392,In_2032,In_293);
nand U393 (N_393,In_2182,In_1443);
nand U394 (N_394,In_671,N_25);
xor U395 (N_395,In_825,N_154);
nand U396 (N_396,In_2341,In_1137);
and U397 (N_397,In_1014,N_30);
and U398 (N_398,In_1805,In_543);
or U399 (N_399,In_479,N_74);
xnor U400 (N_400,In_1778,N_141);
and U401 (N_401,N_10,In_723);
or U402 (N_402,In_2197,In_959);
or U403 (N_403,In_2002,In_428);
xor U404 (N_404,In_624,In_562);
xor U405 (N_405,In_1709,In_135);
xnor U406 (N_406,In_121,In_1405);
or U407 (N_407,N_33,In_294);
xor U408 (N_408,In_643,In_658);
nand U409 (N_409,In_2291,N_13);
nand U410 (N_410,N_188,In_82);
and U411 (N_411,N_321,In_855);
xnor U412 (N_412,In_381,In_1692);
nand U413 (N_413,In_302,In_2222);
or U414 (N_414,In_1419,In_1475);
nand U415 (N_415,In_612,In_1901);
nand U416 (N_416,In_764,In_1940);
xor U417 (N_417,In_217,In_539);
nor U418 (N_418,In_1411,N_366);
or U419 (N_419,N_295,In_433);
and U420 (N_420,In_1275,In_1751);
or U421 (N_421,In_141,In_1112);
nor U422 (N_422,In_491,In_887);
and U423 (N_423,In_153,In_1947);
or U424 (N_424,In_1979,In_737);
nor U425 (N_425,In_2147,In_1653);
xor U426 (N_426,In_2367,In_1627);
nand U427 (N_427,In_282,In_1929);
nor U428 (N_428,In_719,N_225);
xor U429 (N_429,In_307,In_2117);
nand U430 (N_430,In_904,In_1472);
or U431 (N_431,N_95,In_237);
nand U432 (N_432,In_393,In_485);
or U433 (N_433,In_2443,In_1559);
or U434 (N_434,In_69,In_374);
nor U435 (N_435,In_1970,In_2356);
or U436 (N_436,In_1535,In_1241);
nor U437 (N_437,In_2383,In_1745);
nand U438 (N_438,In_313,In_1039);
and U439 (N_439,In_1930,In_347);
nor U440 (N_440,In_1438,In_406);
nor U441 (N_441,N_190,In_239);
xor U442 (N_442,N_81,In_846);
nand U443 (N_443,In_1365,In_681);
nand U444 (N_444,In_500,In_618);
xnor U445 (N_445,N_224,In_596);
and U446 (N_446,In_1879,N_264);
xnor U447 (N_447,In_1723,In_106);
or U448 (N_448,In_1564,In_76);
nor U449 (N_449,In_935,In_774);
nand U450 (N_450,In_392,In_2384);
xnor U451 (N_451,In_1340,In_2264);
nand U452 (N_452,N_277,N_197);
nor U453 (N_453,In_319,In_203);
nand U454 (N_454,In_2046,In_1423);
xor U455 (N_455,In_2012,In_655);
and U456 (N_456,In_981,N_370);
nor U457 (N_457,In_1442,In_704);
xnor U458 (N_458,In_1490,In_765);
nor U459 (N_459,In_813,In_2448);
and U460 (N_460,In_1450,In_309);
nor U461 (N_461,In_1819,In_1763);
nand U462 (N_462,In_891,In_1059);
and U463 (N_463,N_351,In_1500);
nand U464 (N_464,In_1073,In_1207);
or U465 (N_465,In_1836,In_1937);
xnor U466 (N_466,In_389,In_1688);
or U467 (N_467,In_458,In_169);
or U468 (N_468,In_1782,In_2412);
nor U469 (N_469,In_1583,In_976);
xor U470 (N_470,In_1935,N_189);
nand U471 (N_471,N_349,In_131);
nand U472 (N_472,In_2430,In_1995);
and U473 (N_473,In_1662,N_394);
or U474 (N_474,In_422,In_1312);
or U475 (N_475,In_717,In_1202);
or U476 (N_476,N_42,In_2286);
nor U477 (N_477,In_2088,In_1827);
nor U478 (N_478,In_2308,In_916);
or U479 (N_479,In_639,In_2487);
nor U480 (N_480,In_105,In_1983);
or U481 (N_481,In_2300,In_906);
or U482 (N_482,In_2332,In_1603);
or U483 (N_483,In_1027,In_617);
and U484 (N_484,In_1436,In_2148);
or U485 (N_485,N_118,In_2026);
nor U486 (N_486,In_1591,In_1102);
nor U487 (N_487,In_2040,In_2074);
nor U488 (N_488,In_1965,In_1685);
nand U489 (N_489,In_615,N_17);
and U490 (N_490,In_792,N_12);
or U491 (N_491,In_1426,In_2413);
nor U492 (N_492,In_1605,In_11);
xnor U493 (N_493,In_2377,In_320);
nand U494 (N_494,N_88,N_196);
or U495 (N_495,In_597,In_2403);
xnor U496 (N_496,In_116,In_251);
or U497 (N_497,In_2444,In_2425);
nor U498 (N_498,In_484,In_843);
and U499 (N_499,In_2289,In_298);
xnor U500 (N_500,In_504,In_2390);
xnor U501 (N_501,In_1007,In_2436);
and U502 (N_502,In_1948,In_56);
or U503 (N_503,In_731,In_1143);
and U504 (N_504,In_1174,In_1784);
or U505 (N_505,In_1924,In_182);
nor U506 (N_506,In_366,In_1315);
nor U507 (N_507,In_192,In_117);
xnor U508 (N_508,In_929,N_163);
xnor U509 (N_509,In_586,In_1393);
and U510 (N_510,In_2405,In_1943);
xnor U511 (N_511,N_92,In_1259);
xnor U512 (N_512,In_1739,In_409);
nor U513 (N_513,In_786,N_218);
nor U514 (N_514,In_2162,N_202);
nor U515 (N_515,In_1002,In_477);
xor U516 (N_516,In_966,In_2187);
nor U517 (N_517,In_838,N_143);
nor U518 (N_518,In_2039,In_2059);
xnor U519 (N_519,In_1831,In_495);
xor U520 (N_520,N_179,In_323);
xnor U521 (N_521,In_2274,In_176);
xnor U522 (N_522,In_1840,In_663);
xor U523 (N_523,N_28,In_494);
xor U524 (N_524,In_1460,In_1492);
nor U525 (N_525,In_1036,N_18);
xor U526 (N_526,In_1409,In_879);
nand U527 (N_527,In_676,N_24);
nand U528 (N_528,N_50,In_2016);
or U529 (N_529,In_2454,In_99);
and U530 (N_530,In_2371,N_268);
and U531 (N_531,N_39,N_230);
nand U532 (N_532,N_338,In_1029);
xor U533 (N_533,N_373,In_1479);
nor U534 (N_534,In_572,In_1183);
or U535 (N_535,In_2355,In_299);
and U536 (N_536,In_424,In_1433);
nor U537 (N_537,N_286,In_1220);
nand U538 (N_538,In_1098,In_1286);
nand U539 (N_539,In_291,In_103);
and U540 (N_540,N_223,In_148);
xor U541 (N_541,In_330,In_1004);
or U542 (N_542,In_698,N_353);
nor U543 (N_543,In_2206,In_1755);
nand U544 (N_544,In_429,In_2247);
nor U545 (N_545,In_2328,N_234);
nand U546 (N_546,In_1736,In_853);
nor U547 (N_547,In_2415,N_23);
nand U548 (N_548,In_242,In_1431);
nand U549 (N_549,In_53,In_1689);
or U550 (N_550,N_389,In_2167);
or U551 (N_551,In_851,In_1288);
xor U552 (N_552,N_252,In_691);
nor U553 (N_553,In_1536,In_1681);
nor U554 (N_554,In_700,In_728);
and U555 (N_555,N_269,In_2134);
xor U556 (N_556,In_1762,In_1909);
xnor U557 (N_557,In_756,In_670);
and U558 (N_558,In_1859,In_1040);
nand U559 (N_559,In_1705,In_2467);
or U560 (N_560,N_226,In_1636);
nor U561 (N_561,In_733,In_1747);
and U562 (N_562,In_142,In_1130);
or U563 (N_563,In_36,In_2393);
or U564 (N_564,In_459,In_2111);
xor U565 (N_565,In_1563,In_1149);
or U566 (N_566,In_23,In_1515);
or U567 (N_567,In_538,In_339);
and U568 (N_568,In_160,In_1048);
nand U569 (N_569,In_48,In_1330);
or U570 (N_570,In_474,In_2385);
or U571 (N_571,In_1463,In_1444);
nor U572 (N_572,In_565,In_2174);
nor U573 (N_573,In_481,In_1087);
or U574 (N_574,N_367,In_2331);
and U575 (N_575,N_130,In_346);
and U576 (N_576,In_2151,N_147);
xor U577 (N_577,In_1181,In_483);
or U578 (N_578,In_2374,In_809);
and U579 (N_579,In_2426,In_2258);
and U580 (N_580,In_1725,In_1611);
nand U581 (N_581,In_1146,In_1733);
and U582 (N_582,In_1201,In_1615);
nor U583 (N_583,In_883,In_893);
nand U584 (N_584,In_912,In_848);
xnor U585 (N_585,N_121,In_2124);
nand U586 (N_586,In_1377,N_346);
xor U587 (N_587,In_1390,In_17);
xnor U588 (N_588,In_730,In_1044);
or U589 (N_589,In_25,In_1552);
or U590 (N_590,N_116,In_2255);
and U591 (N_591,In_687,In_1026);
and U592 (N_592,In_1820,In_684);
and U593 (N_593,In_2435,In_1654);
or U594 (N_594,In_2307,In_61);
xor U595 (N_595,N_89,In_1240);
or U596 (N_596,In_2419,In_913);
and U597 (N_597,N_270,In_1389);
nand U598 (N_598,N_117,In_1306);
xnor U599 (N_599,In_1299,In_1731);
and U600 (N_600,In_1770,In_1573);
nor U601 (N_601,N_245,In_908);
nor U602 (N_602,In_204,In_2036);
and U603 (N_603,N_108,N_476);
nor U604 (N_604,N_543,In_2323);
or U605 (N_605,N_481,In_1332);
or U606 (N_606,In_583,N_51);
nor U607 (N_607,N_512,N_253);
nor U608 (N_608,In_310,In_550);
nor U609 (N_609,In_2031,In_1006);
xnor U610 (N_610,In_510,In_2080);
nor U611 (N_611,In_990,N_546);
nor U612 (N_612,In_630,N_31);
nand U613 (N_613,In_1971,In_2106);
nand U614 (N_614,N_560,In_188);
xnor U615 (N_615,In_229,N_323);
nor U616 (N_616,N_249,In_1683);
nor U617 (N_617,In_545,N_164);
xnor U618 (N_618,N_380,N_590);
nand U619 (N_619,In_2041,In_2161);
nand U620 (N_620,N_596,In_1404);
nor U621 (N_621,N_227,N_361);
nand U622 (N_622,In_1508,In_2004);
nand U623 (N_623,In_152,In_214);
or U624 (N_624,N_331,In_714);
and U625 (N_625,In_274,N_281);
or U626 (N_626,N_62,In_1421);
nor U627 (N_627,In_1643,N_376);
xnor U628 (N_628,N_483,In_1374);
nand U629 (N_629,In_1867,In_2104);
nor U630 (N_630,In_2280,N_60);
nand U631 (N_631,In_1600,In_1482);
or U632 (N_632,In_2068,N_369);
nor U633 (N_633,In_1328,In_470);
nand U634 (N_634,In_446,N_181);
nor U635 (N_635,In_650,In_2230);
or U636 (N_636,N_595,In_1922);
xor U637 (N_637,In_1349,In_367);
and U638 (N_638,In_514,N_244);
or U639 (N_639,In_405,In_2306);
nor U640 (N_640,In_1944,In_1380);
and U641 (N_641,N_469,In_870);
nand U642 (N_642,In_2067,N_385);
nand U643 (N_643,In_390,In_993);
or U644 (N_644,N_131,In_1495);
or U645 (N_645,N_87,In_1305);
xor U646 (N_646,In_2482,In_261);
or U647 (N_647,In_1750,In_129);
xor U648 (N_648,In_1795,In_972);
or U649 (N_649,In_418,In_1687);
nor U650 (N_650,In_2231,In_100);
xor U651 (N_651,In_1889,In_1099);
or U652 (N_652,In_335,In_2160);
xor U653 (N_653,In_1949,In_332);
xor U654 (N_654,In_2226,N_496);
and U655 (N_655,In_1941,In_2233);
and U656 (N_656,In_884,In_403);
xnor U657 (N_657,N_431,In_341);
and U658 (N_658,In_1912,N_550);
nand U659 (N_659,N_418,N_516);
nor U660 (N_660,In_1516,N_258);
or U661 (N_661,In_629,N_460);
nor U662 (N_662,In_522,In_1372);
and U663 (N_663,N_97,N_337);
xor U664 (N_664,In_1092,N_311);
or U665 (N_665,In_1163,N_19);
or U666 (N_666,N_211,In_1895);
nand U667 (N_667,N_112,In_2422);
nand U668 (N_668,In_1141,In_880);
nor U669 (N_669,In_1699,In_196);
xnor U670 (N_670,In_1581,In_1560);
or U671 (N_671,In_1211,In_186);
and U672 (N_672,In_832,In_1023);
or U673 (N_673,In_1872,In_1873);
and U674 (N_674,N_263,In_2186);
and U675 (N_675,N_217,In_1927);
nor U676 (N_676,In_553,N_135);
and U677 (N_677,In_365,In_1796);
xor U678 (N_678,In_1410,In_1291);
nand U679 (N_679,N_150,N_363);
and U680 (N_680,In_531,In_529);
xnor U681 (N_681,N_47,In_1900);
nor U682 (N_682,In_778,In_942);
or U683 (N_683,In_2399,N_38);
and U684 (N_684,N_557,N_152);
or U685 (N_685,In_2450,N_241);
nor U686 (N_686,N_326,In_535);
nor U687 (N_687,N_582,N_548);
or U688 (N_688,In_599,In_9);
and U689 (N_689,In_1557,In_1243);
nor U690 (N_690,In_977,N_44);
or U691 (N_691,In_42,In_967);
or U692 (N_692,In_862,In_503);
xor U693 (N_693,N_475,In_285);
or U694 (N_694,In_1624,N_348);
nor U695 (N_695,N_257,In_1674);
nand U696 (N_696,In_1403,In_645);
nor U697 (N_697,In_2311,In_1473);
xor U698 (N_698,N_427,In_145);
nor U699 (N_699,N_166,In_994);
nor U700 (N_700,In_2441,In_1093);
nand U701 (N_701,N_246,In_1789);
xor U702 (N_702,In_798,In_1985);
nand U703 (N_703,N_440,In_2172);
or U704 (N_704,In_1406,In_1539);
nor U705 (N_705,In_101,In_1317);
nor U706 (N_706,In_736,In_871);
and U707 (N_707,In_2157,In_1635);
xnor U708 (N_708,In_1682,In_2232);
xor U709 (N_709,In_1351,N_486);
xnor U710 (N_710,In_1077,N_506);
and U711 (N_711,In_1001,In_1567);
nand U712 (N_712,In_1030,In_975);
nand U713 (N_713,In_1590,N_78);
xnor U714 (N_714,In_1273,In_1089);
xnor U715 (N_715,In_2297,In_1336);
nor U716 (N_716,N_423,In_1621);
and U717 (N_717,In_1256,N_451);
nor U718 (N_718,In_241,In_253);
nor U719 (N_719,In_1072,N_442);
xor U720 (N_720,In_1822,In_6);
nand U721 (N_721,In_1734,In_1237);
and U722 (N_722,In_1329,In_2090);
nand U723 (N_723,N_288,In_523);
and U724 (N_724,In_1212,In_2397);
nor U725 (N_725,In_578,N_443);
or U726 (N_726,In_2287,In_2305);
or U727 (N_727,In_1851,In_1079);
xor U728 (N_728,N_41,N_479);
or U729 (N_729,N_156,In_1341);
xor U730 (N_730,In_1658,N_419);
nor U731 (N_731,In_1817,N_289);
or U732 (N_732,In_594,In_1551);
nor U733 (N_733,N_558,In_444);
nor U734 (N_734,In_308,In_1249);
or U735 (N_735,In_271,In_547);
xnor U736 (N_736,In_2458,In_1810);
and U737 (N_737,In_872,N_523);
or U738 (N_738,N_322,In_2285);
nor U739 (N_739,N_238,In_1936);
or U740 (N_740,In_743,In_2142);
and U741 (N_741,In_1669,N_22);
or U742 (N_742,In_828,In_1348);
and U743 (N_743,N_29,In_1575);
and U744 (N_744,N_549,In_1752);
nor U745 (N_745,In_455,In_1896);
or U746 (N_746,N_371,In_19);
and U747 (N_747,N_57,In_585);
nand U748 (N_748,In_2202,In_15);
nor U749 (N_749,In_1768,In_1078);
or U750 (N_750,In_342,In_1366);
and U751 (N_751,In_609,N_77);
nand U752 (N_752,In_1284,In_1053);
nor U753 (N_753,In_760,In_482);
nand U754 (N_754,N_532,In_1832);
and U755 (N_755,N_448,In_1878);
nor U756 (N_756,In_1226,In_1034);
xnor U757 (N_757,N_36,In_2299);
nor U758 (N_758,N_424,In_548);
nand U759 (N_759,In_1546,In_252);
and U760 (N_760,In_2082,In_1828);
xnor U761 (N_761,In_34,N_140);
xnor U762 (N_762,N_0,In_1910);
xnor U763 (N_763,In_1791,In_1538);
and U764 (N_764,N_195,N_259);
and U765 (N_765,In_2180,In_120);
xnor U766 (N_766,In_2329,In_2208);
nor U767 (N_767,In_165,In_2011);
nor U768 (N_768,N_485,N_445);
or U769 (N_769,N_452,In_39);
nor U770 (N_770,In_699,In_1601);
nand U771 (N_771,In_1541,In_1800);
xor U772 (N_772,In_1846,In_2330);
nor U773 (N_773,In_1888,N_110);
or U774 (N_774,In_210,In_1835);
and U775 (N_775,In_2279,In_89);
nor U776 (N_776,In_1385,N_502);
xor U777 (N_777,N_339,In_1247);
nor U778 (N_778,In_2391,N_79);
xor U779 (N_779,In_1402,In_952);
nor U780 (N_780,In_2152,In_849);
xor U781 (N_781,In_355,N_547);
nand U782 (N_782,N_499,In_2259);
nor U783 (N_783,In_1266,N_474);
or U784 (N_784,In_2051,In_146);
xnor U785 (N_785,In_2089,In_1012);
and U786 (N_786,In_1221,In_369);
nor U787 (N_787,N_530,N_165);
nor U788 (N_788,In_634,In_654);
nand U789 (N_789,In_2216,N_578);
nand U790 (N_790,N_591,In_115);
and U791 (N_791,In_1870,N_75);
nor U792 (N_792,In_1161,N_27);
nand U793 (N_793,N_228,In_1337);
xor U794 (N_794,In_2372,In_2318);
xnor U795 (N_795,In_1151,In_71);
xor U796 (N_796,In_316,N_35);
and U797 (N_797,In_59,N_21);
nand U798 (N_798,In_1969,N_421);
and U799 (N_799,In_2337,In_1531);
nand U800 (N_800,N_235,In_1588);
and U801 (N_801,In_292,In_1865);
nand U802 (N_802,In_534,In_1496);
or U803 (N_803,N_712,In_1732);
xor U804 (N_804,N_618,N_649);
or U805 (N_805,N_538,N_465);
or U806 (N_806,In_858,In_1313);
nand U807 (N_807,In_580,In_1701);
nor U808 (N_808,In_246,In_21);
or U809 (N_809,In_574,In_505);
and U810 (N_810,In_1159,N_216);
nand U811 (N_811,N_393,In_1414);
and U812 (N_812,In_1821,In_1115);
and U813 (N_813,N_727,In_652);
nor U814 (N_814,In_2173,In_1644);
and U815 (N_815,N_702,N_626);
or U816 (N_816,In_1730,In_1302);
and U817 (N_817,In_2100,N_470);
and U818 (N_818,N_436,N_407);
nor U819 (N_819,N_310,In_191);
nand U820 (N_820,N_580,In_1858);
nor U821 (N_821,N_168,N_136);
nor U822 (N_822,In_1735,In_1448);
or U823 (N_823,In_1105,N_344);
xnor U824 (N_824,N_587,N_53);
and U825 (N_825,In_757,N_497);
xor U826 (N_826,In_197,In_1543);
nand U827 (N_827,In_674,N_302);
and U828 (N_828,In_836,In_1587);
or U829 (N_829,In_1197,N_240);
or U830 (N_830,In_626,In_796);
and U831 (N_831,In_465,N_535);
nand U832 (N_832,In_2225,In_2135);
nor U833 (N_833,In_1933,In_2098);
and U834 (N_834,In_35,In_441);
xnor U835 (N_835,N_575,In_1042);
or U836 (N_836,N_774,In_2064);
and U837 (N_837,In_555,In_413);
nor U838 (N_838,N_319,In_899);
nor U839 (N_839,In_915,N_740);
and U840 (N_840,In_2030,In_1043);
nand U841 (N_841,In_2471,In_268);
xnor U842 (N_842,In_2058,In_711);
nand U843 (N_843,N_638,In_408);
or U844 (N_844,N_248,In_1715);
nor U845 (N_845,In_281,N_318);
and U846 (N_846,N_375,In_552);
xnor U847 (N_847,In_57,N_105);
nand U848 (N_848,In_1011,In_1103);
and U849 (N_849,In_1210,N_416);
xnor U850 (N_850,In_749,In_564);
xnor U851 (N_851,In_1883,In_513);
and U852 (N_852,In_665,In_1354);
nor U853 (N_853,In_438,In_1884);
or U854 (N_854,N_350,N_604);
nand U855 (N_855,In_2325,In_588);
nor U856 (N_856,In_802,In_876);
or U857 (N_857,In_2035,In_451);
nor U858 (N_858,In_1097,In_2072);
or U859 (N_859,N_632,N_272);
nand U860 (N_860,N_628,In_1425);
and U861 (N_861,In_1976,In_985);
nand U862 (N_862,In_2063,N_745);
xor U863 (N_863,N_680,In_2265);
nand U864 (N_864,N_518,In_1680);
xor U865 (N_865,In_463,In_2196);
and U866 (N_866,In_1830,In_173);
nor U867 (N_867,In_715,In_1876);
nor U868 (N_868,N_529,N_52);
xor U869 (N_869,In_2373,In_31);
nor U870 (N_870,N_103,In_1488);
nand U871 (N_871,N_400,In_1717);
nand U872 (N_872,In_2402,N_501);
nor U873 (N_873,In_1068,N_644);
nor U874 (N_874,In_2312,In_2378);
xor U875 (N_875,In_1716,In_2234);
or U876 (N_876,N_659,In_1407);
nor U877 (N_877,N_273,In_327);
nor U878 (N_878,In_1468,In_2348);
or U879 (N_879,In_1885,N_384);
nor U880 (N_880,In_2017,In_2155);
nor U881 (N_881,In_1544,In_1994);
and U882 (N_882,In_2361,In_740);
nor U883 (N_883,In_713,In_2087);
or U884 (N_884,In_2282,In_1485);
nand U885 (N_885,In_2459,In_1217);
nor U886 (N_886,In_1487,N_482);
or U887 (N_887,In_1274,In_304);
and U888 (N_888,In_1276,N_343);
xnor U889 (N_889,In_356,In_200);
xnor U890 (N_890,In_1592,N_282);
xor U891 (N_891,In_1499,N_449);
nand U892 (N_892,In_2319,N_720);
xor U893 (N_893,In_171,In_1470);
nand U894 (N_894,N_294,In_487);
and U895 (N_895,In_823,N_83);
nor U896 (N_896,In_7,N_6);
and U897 (N_897,In_829,In_1371);
nor U898 (N_898,N_410,In_1632);
or U899 (N_899,N_603,In_305);
xnor U900 (N_900,In_314,In_1408);
or U901 (N_901,In_1063,N_794);
xor U902 (N_902,In_1738,N_645);
or U903 (N_903,In_576,In_840);
nand U904 (N_904,N_625,In_1265);
nor U905 (N_905,In_751,In_903);
or U906 (N_906,In_2346,In_88);
nand U907 (N_907,N_677,In_26);
nor U908 (N_908,In_1086,In_1703);
nor U909 (N_909,N_608,In_163);
and U910 (N_910,In_2228,In_297);
xnor U911 (N_911,In_2029,N_432);
nor U912 (N_912,In_32,In_841);
or U913 (N_913,In_1594,N_94);
or U914 (N_914,In_2149,N_544);
xnor U915 (N_915,N_707,In_1360);
xor U916 (N_916,In_881,In_2469);
and U917 (N_917,In_1570,N_699);
xor U918 (N_918,N_134,In_1323);
xor U919 (N_919,N_489,N_247);
and U920 (N_920,In_556,N_619);
or U921 (N_921,In_486,N_236);
nand U922 (N_922,N_588,N_98);
nand U923 (N_923,In_1641,N_510);
xor U924 (N_924,N_415,In_939);
xnor U925 (N_925,In_379,In_456);
nand U926 (N_926,N_737,In_364);
nor U927 (N_927,In_2417,N_34);
nand U928 (N_928,In_2404,N_260);
xor U929 (N_929,In_179,N_567);
xor U930 (N_930,N_251,N_171);
xor U931 (N_931,N_161,N_40);
xnor U932 (N_932,In_2219,N_507);
and U933 (N_933,In_1361,In_1129);
or U934 (N_934,In_2037,In_1254);
nand U935 (N_935,N_764,In_520);
and U936 (N_936,In_1236,N_204);
or U937 (N_937,In_821,In_1525);
xor U938 (N_938,In_1547,In_2483);
xor U939 (N_939,N_70,In_1964);
nor U940 (N_940,N_453,In_1205);
and U941 (N_941,N_577,In_1607);
xor U942 (N_942,In_992,N_657);
nand U943 (N_943,In_289,N_133);
or U944 (N_944,In_971,In_1301);
xor U945 (N_945,In_2235,In_1841);
and U946 (N_946,In_1420,In_805);
or U947 (N_947,In_202,N_563);
nand U948 (N_948,N_297,In_1978);
xor U949 (N_949,In_1887,In_235);
nor U950 (N_950,N_377,In_1874);
and U951 (N_951,In_1218,In_873);
and U952 (N_952,N_574,N_682);
xnor U953 (N_953,In_1807,In_60);
xor U954 (N_954,In_2165,In_1524);
nand U955 (N_955,In_1646,N_194);
nand U956 (N_956,N_333,In_1839);
xor U957 (N_957,In_512,N_237);
nand U958 (N_958,In_1287,N_674);
nand U959 (N_959,N_317,In_1088);
or U960 (N_960,In_2075,In_1504);
nand U961 (N_961,In_2363,In_1262);
xnor U962 (N_962,N_82,In_800);
and U963 (N_963,In_1069,In_1697);
and U964 (N_964,In_1338,N_59);
xnor U965 (N_965,N_111,In_807);
xor U966 (N_966,In_228,In_40);
xor U967 (N_967,In_2455,In_2438);
and U968 (N_968,In_2136,In_1769);
nand U969 (N_969,N_606,N_412);
xor U970 (N_970,In_2062,In_399);
and U971 (N_971,In_1445,N_54);
nor U972 (N_972,In_385,N_671);
nand U973 (N_973,In_2175,In_502);
nor U974 (N_974,In_1756,N_327);
or U975 (N_975,N_528,In_1228);
nor U976 (N_976,In_1191,In_2498);
or U977 (N_977,In_739,N_505);
nand U978 (N_978,In_194,In_2112);
or U979 (N_979,In_93,N_636);
xnor U980 (N_980,N_661,In_1779);
nand U981 (N_981,In_208,N_11);
nor U982 (N_982,In_2327,In_380);
xnor U983 (N_983,In_777,In_648);
nor U984 (N_984,In_2171,N_646);
or U985 (N_985,In_449,N_9);
nor U986 (N_986,N_613,In_2083);
nand U987 (N_987,N_692,N_276);
and U988 (N_988,N_313,N_222);
nor U989 (N_989,In_324,In_1672);
nand U990 (N_990,In_2303,In_490);
xor U991 (N_991,N_63,In_345);
and U992 (N_992,In_897,In_675);
nor U993 (N_993,N_688,In_1399);
nor U994 (N_994,In_1638,In_2351);
or U995 (N_995,N_461,N_769);
nand U996 (N_996,N_255,In_1128);
xnor U997 (N_997,N_723,N_472);
nor U998 (N_998,N_434,N_668);
xnor U999 (N_999,In_1675,In_2126);
or U1000 (N_1000,N_200,N_944);
nand U1001 (N_1001,N_684,In_2261);
nand U1002 (N_1002,N_797,In_2394);
xor U1003 (N_1003,N_690,In_1271);
nor U1004 (N_1004,N_663,N_32);
nand U1005 (N_1005,In_81,In_710);
or U1006 (N_1006,In_1860,In_1951);
xnor U1007 (N_1007,In_279,In_2015);
xor U1008 (N_1008,In_357,In_2431);
or U1009 (N_1009,In_2199,In_2054);
xnor U1010 (N_1010,In_963,In_541);
nor U1011 (N_1011,In_1767,N_655);
nor U1012 (N_1012,In_1396,In_2188);
xnor U1013 (N_1013,In_934,In_2392);
nand U1014 (N_1014,In_709,In_1788);
or U1015 (N_1015,In_725,N_988);
or U1016 (N_1016,N_262,In_1041);
or U1017 (N_1017,N_838,N_524);
xor U1018 (N_1018,In_1369,In_1045);
nor U1019 (N_1019,N_275,N_714);
or U1020 (N_1020,In_1160,N_610);
nor U1021 (N_1021,N_926,N_772);
and U1022 (N_1022,N_700,In_2205);
nand U1023 (N_1023,N_979,In_919);
and U1024 (N_1024,In_1074,In_566);
and U1025 (N_1025,In_85,In_801);
and U1026 (N_1026,In_27,In_2169);
or U1027 (N_1027,N_629,N_402);
nand U1028 (N_1028,N_458,N_368);
nand U1029 (N_1029,In_1257,In_250);
nor U1030 (N_1030,N_883,In_488);
nor U1031 (N_1031,In_1188,N_456);
and U1032 (N_1032,In_1711,In_878);
nor U1033 (N_1033,In_1134,N_834);
and U1034 (N_1034,In_1216,In_1);
and U1035 (N_1035,In_1198,In_67);
nand U1036 (N_1036,In_1430,N_328);
nor U1037 (N_1037,In_256,In_1439);
and U1038 (N_1038,In_140,N_492);
and U1039 (N_1039,In_1021,In_2381);
xor U1040 (N_1040,N_809,N_857);
or U1041 (N_1041,In_1474,N_142);
xnor U1042 (N_1042,N_754,In_1803);
or U1043 (N_1043,In_1748,In_2322);
nand U1044 (N_1044,In_2213,In_1148);
or U1045 (N_1045,In_322,In_2427);
and U1046 (N_1046,In_1998,In_940);
and U1047 (N_1047,N_840,N_292);
or U1048 (N_1048,In_1107,In_1852);
nor U1049 (N_1049,N_732,In_842);
and U1050 (N_1050,N_519,In_953);
nand U1051 (N_1051,N_974,In_622);
nand U1052 (N_1052,N_175,N_826);
and U1053 (N_1053,In_2246,In_1359);
nor U1054 (N_1054,In_1154,In_2464);
xnor U1055 (N_1055,In_1033,N_823);
or U1056 (N_1056,In_1147,In_1710);
and U1057 (N_1057,N_330,In_1571);
and U1058 (N_1058,In_773,N_881);
xnor U1059 (N_1059,In_806,In_922);
and U1060 (N_1060,N_783,N_447);
nand U1061 (N_1061,In_1150,In_340);
nand U1062 (N_1062,N_521,N_69);
or U1063 (N_1063,In_1096,N_989);
nor U1064 (N_1064,In_623,N_803);
nor U1065 (N_1065,N_752,N_962);
nor U1066 (N_1066,In_2006,In_1428);
or U1067 (N_1067,N_266,N_387);
nand U1068 (N_1068,In_1868,In_2034);
nor U1069 (N_1069,N_533,In_2370);
or U1070 (N_1070,In_2251,In_1435);
or U1071 (N_1071,In_265,In_363);
nor U1072 (N_1072,N_307,In_682);
and U1073 (N_1073,N_593,In_2447);
xnor U1074 (N_1074,In_1881,N_836);
and U1075 (N_1075,In_785,In_1037);
xnor U1076 (N_1076,In_1517,In_559);
xor U1077 (N_1077,In_1657,N_860);
and U1078 (N_1078,In_2423,N_335);
nand U1079 (N_1079,In_1224,In_2473);
nor U1080 (N_1080,In_118,In_1869);
or U1081 (N_1081,In_722,In_811);
nor U1082 (N_1082,In_1954,N_819);
and U1083 (N_1083,In_2097,N_757);
nand U1084 (N_1084,In_1585,In_1760);
and U1085 (N_1085,N_541,In_1956);
nor U1086 (N_1086,In_635,In_557);
nand U1087 (N_1087,N_561,In_1483);
or U1088 (N_1088,N_791,N_243);
nor U1089 (N_1089,In_1417,In_1540);
nor U1090 (N_1090,N_842,N_945);
nand U1091 (N_1091,In_2304,N_439);
xor U1092 (N_1092,N_695,In_885);
nor U1093 (N_1093,In_1263,N_743);
or U1094 (N_1094,In_419,N_854);
or U1095 (N_1095,N_929,In_1242);
xnor U1096 (N_1096,In_1140,N_818);
nor U1097 (N_1097,N_58,In_2456);
nor U1098 (N_1098,In_1126,In_1229);
nand U1099 (N_1099,N_748,In_794);
and U1100 (N_1100,N_951,N_833);
and U1101 (N_1101,In_1676,In_803);
or U1102 (N_1102,In_2043,In_22);
xor U1103 (N_1103,In_726,In_2091);
nor U1104 (N_1104,N_360,In_686);
or U1105 (N_1105,In_398,In_694);
nand U1106 (N_1106,N_399,In_1110);
nand U1107 (N_1107,N_146,In_961);
xor U1108 (N_1108,In_1267,In_1494);
nand U1109 (N_1109,In_431,In_2494);
nand U1110 (N_1110,N_8,N_500);
nand U1111 (N_1111,N_404,In_834);
and U1112 (N_1112,N_865,N_357);
nor U1113 (N_1113,N_68,N_763);
xor U1114 (N_1114,In_255,N_61);
and U1115 (N_1115,In_14,N_824);
nand U1116 (N_1116,In_223,N_799);
xnor U1117 (N_1117,In_189,In_1164);
and U1118 (N_1118,N_969,N_250);
nand U1119 (N_1119,In_410,In_2493);
nor U1120 (N_1120,N_417,In_1501);
nand U1121 (N_1121,In_2178,N_114);
nor U1122 (N_1122,In_2000,In_425);
nor U1123 (N_1123,In_1637,In_432);
xor U1124 (N_1124,N_662,In_1758);
and U1125 (N_1125,N_893,In_161);
nor U1126 (N_1126,N_630,In_991);
xor U1127 (N_1127,N_701,In_1489);
nand U1128 (N_1128,In_1082,N_765);
nand U1129 (N_1129,In_2270,N_949);
xor U1130 (N_1130,In_1561,N_759);
nor U1131 (N_1131,In_779,N_254);
or U1132 (N_1132,N_579,N_849);
or U1133 (N_1133,N_76,In_2239);
xor U1134 (N_1134,In_1843,In_1018);
xor U1135 (N_1135,N_362,N_271);
nor U1136 (N_1136,N_584,N_274);
and U1137 (N_1137,In_1857,In_720);
or U1138 (N_1138,In_1578,In_1022);
xnor U1139 (N_1139,In_1370,N_219);
xnor U1140 (N_1140,In_1898,In_1314);
nand U1141 (N_1141,N_749,In_1025);
nand U1142 (N_1142,In_1376,N_542);
nor U1143 (N_1143,In_1550,In_937);
nor U1144 (N_1144,N_835,N_571);
or U1145 (N_1145,N_895,In_1364);
nor U1146 (N_1146,In_974,In_1378);
or U1147 (N_1147,In_1381,In_2179);
nor U1148 (N_1148,In_1250,In_679);
or U1149 (N_1149,N_341,N_467);
xor U1150 (N_1150,N_975,N_229);
and U1151 (N_1151,In_1195,In_2127);
or U1152 (N_1152,In_2076,In_1204);
or U1153 (N_1153,In_150,In_892);
or U1154 (N_1154,N_422,In_2144);
or U1155 (N_1155,In_815,N_386);
nor U1156 (N_1156,In_1904,In_1977);
nand U1157 (N_1157,N_444,In_989);
and U1158 (N_1158,In_690,In_1783);
and U1159 (N_1159,In_2449,N_304);
and U1160 (N_1160,N_910,In_1152);
nand U1161 (N_1161,In_1722,In_1707);
nor U1162 (N_1162,In_156,In_1319);
nor U1163 (N_1163,In_2108,N_961);
or U1164 (N_1164,In_18,N_514);
or U1165 (N_1165,In_1837,N_927);
and U1166 (N_1166,In_1911,N_471);
xnor U1167 (N_1167,In_5,In_1363);
nor U1168 (N_1168,N_784,N_811);
nor U1169 (N_1169,In_688,In_1906);
nand U1170 (N_1170,In_584,In_2284);
and U1171 (N_1171,In_956,In_2400);
or U1172 (N_1172,In_506,In_689);
or U1173 (N_1173,In_1833,In_546);
and U1174 (N_1174,N_933,N_186);
and U1175 (N_1175,In_1990,N_581);
nand U1176 (N_1176,N_426,In_1579);
and U1177 (N_1177,N_534,N_435);
or U1178 (N_1178,In_92,N_696);
xnor U1179 (N_1179,In_651,In_768);
or U1180 (N_1180,N_395,N_372);
nor U1181 (N_1181,N_201,In_1599);
nor U1182 (N_1182,In_1120,In_1289);
nand U1183 (N_1183,N_766,In_1052);
xnor U1184 (N_1184,N_209,In_45);
or U1185 (N_1185,N_284,N_685);
or U1186 (N_1186,N_964,In_1704);
and U1187 (N_1187,In_166,N_129);
nand U1188 (N_1188,N_828,N_347);
or U1189 (N_1189,N_793,In_2368);
nor U1190 (N_1190,In_1203,N_859);
and U1191 (N_1191,In_382,N_940);
xnor U1192 (N_1192,In_867,N_607);
nor U1193 (N_1193,N_55,N_739);
xor U1194 (N_1194,N_342,In_1584);
nor U1195 (N_1195,In_1091,N_43);
nor U1196 (N_1196,N_788,N_830);
and U1197 (N_1197,In_1923,In_1060);
nand U1198 (N_1198,In_1418,In_1145);
nor U1199 (N_1199,N_789,In_113);
nand U1200 (N_1200,In_244,N_494);
nand U1201 (N_1201,N_401,In_745);
nor U1202 (N_1202,In_1353,N_672);
and U1203 (N_1203,N_722,In_306);
nand U1204 (N_1204,In_1090,N_1133);
xor U1205 (N_1205,In_1737,N_879);
nand U1206 (N_1206,N_513,N_545);
or U1207 (N_1207,In_2424,N_420);
nor U1208 (N_1208,In_837,In_243);
or U1209 (N_1209,N_1151,N_991);
or U1210 (N_1210,In_439,In_2132);
nor U1211 (N_1211,In_1350,N_733);
or U1212 (N_1212,In_2353,N_352);
or U1213 (N_1213,In_2340,In_954);
nor U1214 (N_1214,N_517,In_1422);
nand U1215 (N_1215,N_1130,N_1070);
nand U1216 (N_1216,N_913,N_1159);
nor U1217 (N_1217,N_686,N_642);
and U1218 (N_1218,In_2275,N_600);
nor U1219 (N_1219,In_1005,In_2437);
xnor U1220 (N_1220,N_637,In_1124);
and U1221 (N_1221,In_2154,In_1580);
nand U1222 (N_1222,In_528,N_598);
or U1223 (N_1223,N_1193,N_1098);
or U1224 (N_1224,N_1061,In_2229);
or U1225 (N_1225,N_71,N_1106);
nor U1226 (N_1226,In_358,In_646);
nand U1227 (N_1227,N_758,N_846);
and U1228 (N_1228,In_577,N_746);
and U1229 (N_1229,N_717,N_1067);
nand U1230 (N_1230,In_614,N_1091);
xor U1231 (N_1231,N_623,N_495);
nand U1232 (N_1232,In_1757,In_1379);
or U1233 (N_1233,N_1163,N_994);
nand U1234 (N_1234,In_62,In_759);
and U1235 (N_1235,In_2116,In_1233);
or U1236 (N_1236,N_667,In_2362);
and U1237 (N_1237,In_2021,In_1893);
nor U1238 (N_1238,N_1166,N_617);
xor U1239 (N_1239,In_1062,N_1108);
or U1240 (N_1240,N_73,N_1114);
and U1241 (N_1241,N_848,N_345);
nand U1242 (N_1242,In_917,N_911);
or U1243 (N_1243,N_820,N_918);
and U1244 (N_1244,In_1618,In_276);
or U1245 (N_1245,In_526,In_1434);
nand U1246 (N_1246,In_95,In_2333);
or U1247 (N_1247,N_1035,In_33);
xor U1248 (N_1248,N_320,In_516);
and U1249 (N_1249,In_527,N_455);
and U1250 (N_1250,In_605,N_1170);
or U1251 (N_1251,In_2429,In_2252);
and U1252 (N_1252,In_692,N_891);
nand U1253 (N_1253,N_1093,In_931);
and U1254 (N_1254,In_519,N_851);
nor U1255 (N_1255,N_1143,N_973);
and U1256 (N_1256,N_735,In_569);
xnor U1257 (N_1257,N_1009,N_1120);
xnor U1258 (N_1258,N_947,In_1720);
xnor U1259 (N_1259,N_889,N_950);
and U1260 (N_1260,N_1122,In_1562);
or U1261 (N_1261,In_1774,N_381);
nand U1262 (N_1262,In_248,N_1010);
and U1263 (N_1263,In_2140,N_503);
xnor U1264 (N_1264,N_627,N_1165);
xnor U1265 (N_1265,In_2418,In_70);
nor U1266 (N_1266,N_935,N_429);
and U1267 (N_1267,In_286,N_462);
xnor U1268 (N_1268,N_670,N_586);
nor U1269 (N_1269,N_437,In_240);
xor U1270 (N_1270,N_976,N_1117);
and U1271 (N_1271,N_1027,N_1110);
nor U1272 (N_1272,N_488,N_728);
nor U1273 (N_1273,In_1962,In_763);
nor U1274 (N_1274,N_1017,In_134);
xor U1275 (N_1275,N_556,N_1191);
nand U1276 (N_1276,In_2244,N_980);
xnor U1277 (N_1277,In_353,N_873);
xnor U1278 (N_1278,N_808,N_938);
or U1279 (N_1279,N_1038,N_614);
and U1280 (N_1280,N_620,N_1043);
xnor U1281 (N_1281,In_1864,N_303);
xor U1282 (N_1282,In_1513,N_314);
xor U1283 (N_1283,In_1963,In_1787);
nor U1284 (N_1284,In_997,In_1279);
or U1285 (N_1285,In_1469,In_215);
nand U1286 (N_1286,N_845,In_770);
xnor U1287 (N_1287,N_526,N_1197);
nand U1288 (N_1288,N_1195,N_1001);
or U1289 (N_1289,N_683,N_869);
or U1290 (N_1290,In_167,In_2101);
xor U1291 (N_1291,N_1155,In_613);
nand U1292 (N_1292,In_1908,In_2102);
nor U1293 (N_1293,In_303,N_1141);
xor U1294 (N_1294,N_954,In_910);
nand U1295 (N_1295,N_1105,In_136);
nor U1296 (N_1296,N_525,N_207);
nor U1297 (N_1297,In_2276,In_1534);
nand U1298 (N_1298,In_138,N_886);
or U1299 (N_1299,In_1655,In_2433);
nor U1300 (N_1300,N_1139,N_1171);
and U1301 (N_1301,N_767,In_1690);
or U1302 (N_1302,N_1138,N_267);
nor U1303 (N_1303,N_934,In_1622);
and U1304 (N_1304,N_66,In_360);
nor U1305 (N_1305,In_1297,N_1062);
nand U1306 (N_1306,In_1670,In_447);
xor U1307 (N_1307,N_634,N_864);
nor U1308 (N_1308,N_858,In_254);
nand U1309 (N_1309,In_1017,N_1044);
nand U1310 (N_1310,N_293,N_878);
and U1311 (N_1311,In_1498,In_401);
xor U1312 (N_1312,N_1148,N_805);
and U1313 (N_1313,N_884,N_192);
xor U1314 (N_1314,In_1661,N_599);
or U1315 (N_1315,N_414,In_509);
nand U1316 (N_1316,In_1325,N_566);
nor U1317 (N_1317,N_1131,N_1127);
nor U1318 (N_1318,In_2170,N_570);
and U1319 (N_1319,N_907,N_1113);
and U1320 (N_1320,In_1679,N_741);
or U1321 (N_1321,In_2137,In_2120);
xnor U1322 (N_1322,N_622,In_2121);
xor U1323 (N_1323,N_127,In_2113);
xor U1324 (N_1324,N_298,In_533);
nand U1325 (N_1325,N_792,In_716);
or U1326 (N_1326,In_205,In_1290);
and U1327 (N_1327,In_1084,N_866);
nor U1328 (N_1328,In_563,N_997);
xor U1329 (N_1329,In_1792,N_871);
nor U1330 (N_1330,In_2359,N_708);
or U1331 (N_1331,N_719,In_2316);
xnor U1332 (N_1332,In_445,N_1095);
nand U1333 (N_1333,N_1198,In_839);
nor U1334 (N_1334,N_1128,N_726);
xor U1335 (N_1335,N_329,N_1005);
xnor U1336 (N_1336,In_824,In_2495);
xnor U1337 (N_1337,N_959,N_536);
and U1338 (N_1338,N_37,N_283);
nor U1339 (N_1339,In_2166,N_762);
nand U1340 (N_1340,N_215,N_1081);
nand U1341 (N_1341,N_1162,In_2479);
and U1342 (N_1342,In_16,N_537);
nand U1343 (N_1343,In_1973,N_968);
and U1344 (N_1344,In_1345,In_1945);
xor U1345 (N_1345,N_430,N_123);
or U1346 (N_1346,In_1918,N_1064);
or U1347 (N_1347,N_770,N_899);
nand U1348 (N_1348,N_554,In_2445);
and U1349 (N_1349,In_2336,N_1154);
nand U1350 (N_1350,In_914,N_721);
nor U1351 (N_1351,N_1182,N_1116);
or U1352 (N_1352,In_2497,N_744);
nor U1353 (N_1353,In_2453,N_378);
or U1354 (N_1354,In_218,In_791);
xnor U1355 (N_1355,In_1424,N_162);
nor U1356 (N_1356,In_2131,In_1477);
nand U1357 (N_1357,In_1165,In_925);
nand U1358 (N_1358,N_1167,N_1181);
nand U1359 (N_1359,N_1109,N_609);
nand U1360 (N_1360,N_564,N_650);
xor U1361 (N_1361,N_1188,N_212);
nand U1362 (N_1362,In_817,N_102);
xor U1363 (N_1363,In_1412,In_1673);
nor U1364 (N_1364,N_90,N_1168);
or U1365 (N_1365,In_1866,N_956);
nand U1366 (N_1366,In_570,In_1781);
xor U1367 (N_1367,In_1815,N_742);
nand U1368 (N_1368,N_1156,In_1824);
and U1369 (N_1369,In_1358,In_450);
or U1370 (N_1370,N_568,N_641);
nor U1371 (N_1371,N_174,In_721);
nor U1372 (N_1372,N_1012,N_1097);
nand U1373 (N_1373,N_80,N_1057);
xnor U1374 (N_1374,In_1459,In_685);
and U1375 (N_1375,N_1190,In_1772);
or U1376 (N_1376,In_164,In_1131);
xor U1377 (N_1377,In_1100,N_936);
or U1378 (N_1378,In_567,N_775);
and U1379 (N_1379,N_559,In_2380);
and U1380 (N_1380,N_912,N_957);
nor U1381 (N_1381,In_2129,In_949);
nand U1382 (N_1382,In_1666,In_1741);
nand U1383 (N_1383,N_1089,In_678);
and U1384 (N_1384,N_231,In_2047);
and U1385 (N_1385,In_696,In_443);
nand U1386 (N_1386,In_797,N_853);
nor U1387 (N_1387,In_633,In_2005);
nand U1388 (N_1388,In_1055,In_703);
nand U1389 (N_1389,In_1467,N_565);
nand U1390 (N_1390,In_1556,N_928);
xor U1391 (N_1391,N_48,In_375);
nor U1392 (N_1392,In_1231,N_522);
or U1393 (N_1393,N_1101,In_58);
nor U1394 (N_1394,N_457,N_909);
and U1395 (N_1395,In_1113,In_259);
nor U1396 (N_1396,In_1180,N_301);
nor U1397 (N_1397,In_437,N_1112);
or U1398 (N_1398,N_562,N_1071);
xor U1399 (N_1399,In_386,In_1742);
nand U1400 (N_1400,N_1073,In_262);
nor U1401 (N_1401,N_1002,In_501);
nor U1402 (N_1402,In_1726,In_232);
nand U1403 (N_1403,In_2114,In_1028);
nor U1404 (N_1404,In_209,In_1610);
or U1405 (N_1405,N_1209,N_1184);
and U1406 (N_1406,N_413,In_2414);
or U1407 (N_1407,N_1176,In_2250);
and U1408 (N_1408,N_605,N_900);
nor U1409 (N_1409,N_868,N_1313);
nand U1410 (N_1410,In_1854,N_498);
or U1411 (N_1411,In_2143,N_583);
nand U1412 (N_1412,N_1219,N_1185);
and U1413 (N_1413,N_1096,N_1327);
and U1414 (N_1414,In_1415,N_982);
nand U1415 (N_1415,In_746,N_585);
xor U1416 (N_1416,N_1199,In_1554);
and U1417 (N_1417,N_316,N_1389);
nor U1418 (N_1418,N_1360,In_1346);
xor U1419 (N_1419,N_678,In_1776);
nor U1420 (N_1420,In_1617,In_1392);
nand U1421 (N_1421,N_1092,N_1066);
xnor U1422 (N_1422,In_151,N_983);
nor U1423 (N_1423,N_1380,N_1223);
nor U1424 (N_1424,N_1008,In_1548);
nor U1425 (N_1425,N_210,N_1213);
xnor U1426 (N_1426,N_572,N_611);
nand U1427 (N_1427,In_2364,N_1282);
xor U1428 (N_1428,In_1598,N_635);
nor U1429 (N_1429,In_2194,N_615);
and U1430 (N_1430,N_151,In_1020);
xnor U1431 (N_1431,In_1826,In_124);
nor U1432 (N_1432,N_1194,In_480);
or U1433 (N_1433,N_356,In_683);
nand U1434 (N_1434,N_1399,In_672);
nand U1435 (N_1435,N_1290,In_558);
nor U1436 (N_1436,In_1106,N_388);
nand U1437 (N_1437,N_1118,In_359);
xor U1438 (N_1438,N_1142,In_1258);
nand U1439 (N_1439,In_641,N_1334);
xor U1440 (N_1440,N_1239,N_665);
xnor U1441 (N_1441,In_1310,N_919);
nor U1442 (N_1442,N_795,N_1058);
and U1443 (N_1443,N_239,N_1186);
and U1444 (N_1444,N_882,In_1166);
nor U1445 (N_1445,In_1244,N_862);
xor U1446 (N_1446,In_1465,N_654);
or U1447 (N_1447,In_530,N_1241);
and U1448 (N_1448,N_300,N_1367);
nor U1449 (N_1449,N_1375,In_2296);
nor U1450 (N_1450,In_1058,N_1090);
or U1451 (N_1451,In_13,In_220);
and U1452 (N_1452,N_1121,In_2477);
xor U1453 (N_1453,N_107,N_290);
and U1454 (N_1454,In_1960,N_1229);
and U1455 (N_1455,N_187,In_137);
and U1456 (N_1456,N_1150,N_1119);
or U1457 (N_1457,N_405,N_955);
nor U1458 (N_1458,In_1121,In_780);
or U1459 (N_1459,N_1179,In_122);
xnor U1460 (N_1460,N_1175,N_1390);
nor U1461 (N_1461,In_2164,N_998);
nand U1462 (N_1462,In_2365,N_924);
and U1463 (N_1463,In_478,N_932);
xnor U1464 (N_1464,In_269,N_221);
nand U1465 (N_1465,N_2,N_480);
xnor U1466 (N_1466,In_2018,N_1272);
or U1467 (N_1467,N_1305,In_1222);
or U1468 (N_1468,In_1230,N_1297);
xnor U1469 (N_1469,In_2215,In_1334);
nand U1470 (N_1470,N_800,In_2272);
and U1471 (N_1471,N_291,N_986);
nand U1472 (N_1472,In_420,N_810);
xnor U1473 (N_1473,In_435,In_321);
nand U1474 (N_1474,N_1326,In_2254);
nand U1475 (N_1475,In_231,N_1080);
or U1476 (N_1476,N_1041,N_1330);
nand U1477 (N_1477,In_1173,In_64);
and U1478 (N_1478,N_1345,N_1161);
nand U1479 (N_1479,In_875,In_1047);
nor U1480 (N_1480,In_1718,N_660);
and U1481 (N_1481,In_620,N_1018);
or U1482 (N_1482,N_334,In_2146);
xnor U1483 (N_1483,In_697,N_1087);
nor U1484 (N_1484,In_372,In_162);
xor U1485 (N_1485,In_1708,N_573);
and U1486 (N_1486,N_428,N_287);
nor U1487 (N_1487,N_778,In_415);
xnor U1488 (N_1488,N_520,N_1054);
or U1489 (N_1489,In_590,N_1357);
and U1490 (N_1490,In_2314,In_1298);
or U1491 (N_1491,N_256,N_681);
nand U1492 (N_1492,In_644,N_1065);
xnor U1493 (N_1493,N_1039,In_2489);
nand U1494 (N_1494,N_875,N_106);
xnor U1495 (N_1495,N_379,N_1385);
and U1496 (N_1496,In_1649,N_1342);
nor U1497 (N_1497,In_1386,In_384);
nor U1498 (N_1498,In_1209,N_939);
xnor U1499 (N_1499,In_87,In_2339);
and U1500 (N_1500,In_499,N_126);
nor U1501 (N_1501,N_1246,N_392);
nand U1502 (N_1502,N_850,N_1205);
xor U1503 (N_1503,In_454,N_473);
nand U1504 (N_1504,In_772,N_1031);
and U1505 (N_1505,In_1471,In_1189);
nor U1506 (N_1506,In_272,In_2410);
xor U1507 (N_1507,N_382,N_1249);
xor U1508 (N_1508,In_1344,In_1861);
and U1509 (N_1509,N_183,N_1078);
or U1510 (N_1510,In_602,In_1167);
nand U1511 (N_1511,N_1354,N_508);
and U1512 (N_1512,In_625,In_1577);
nand U1513 (N_1513,N_1014,N_1020);
xnor U1514 (N_1514,N_1216,In_362);
nor U1515 (N_1515,In_414,In_1604);
and U1516 (N_1516,N_1222,N_324);
nand U1517 (N_1517,N_996,N_639);
nand U1518 (N_1518,N_1203,In_287);
nor U1519 (N_1519,N_96,In_1991);
or U1520 (N_1520,N_1270,In_560);
and U1521 (N_1521,N_902,N_1307);
and U1522 (N_1522,In_928,N_182);
and U1523 (N_1523,In_2406,N_1042);
nand U1524 (N_1524,N_1280,In_758);
nor U1525 (N_1525,N_312,N_1160);
or U1526 (N_1526,N_916,In_2360);
or U1527 (N_1527,N_1136,In_119);
nand U1528 (N_1528,N_852,N_1207);
nor U1529 (N_1529,In_1589,In_2320);
and U1530 (N_1530,In_1568,In_417);
or U1531 (N_1531,In_2168,N_652);
and U1532 (N_1532,N_340,N_901);
nor U1533 (N_1533,N_703,N_1126);
and U1534 (N_1534,N_1111,In_1665);
and U1535 (N_1535,N_694,N_1265);
nand U1536 (N_1536,In_245,N_1377);
or U1537 (N_1537,In_518,N_325);
and U1538 (N_1538,In_2241,In_1555);
nand U1539 (N_1539,N_1317,In_66);
xor U1540 (N_1540,In_877,In_2243);
and U1541 (N_1541,In_1798,N_704);
and U1542 (N_1542,In_793,N_806);
nand U1543 (N_1543,N_1204,N_821);
and U1544 (N_1544,N_1045,N_1228);
nor U1545 (N_1545,In_1714,N_72);
xnor U1546 (N_1546,N_1396,N_1135);
and U1547 (N_1547,In_476,N_1388);
and U1548 (N_1548,N_1394,N_1271);
or U1549 (N_1549,N_1137,N_807);
nand U1550 (N_1550,N_233,In_1278);
nor U1551 (N_1551,In_2310,In_2042);
nor U1552 (N_1552,N_1231,In_1136);
nor U1553 (N_1553,In_1400,N_441);
nand U1554 (N_1554,N_779,N_193);
or U1555 (N_1555,N_406,N_1217);
nand U1556 (N_1556,In_325,N_1333);
or U1557 (N_1557,In_378,N_1304);
xor U1558 (N_1558,N_1259,N_1240);
or U1559 (N_1559,In_1808,N_531);
and U1560 (N_1560,In_1192,In_960);
or U1561 (N_1561,In_2049,N_261);
or U1562 (N_1562,N_1048,N_1315);
nand U1563 (N_1563,In_79,N_1276);
nand U1564 (N_1564,N_1321,N_1079);
xnor U1565 (N_1565,In_2079,In_74);
nor U1566 (N_1566,N_1034,N_1132);
xor U1567 (N_1567,N_214,In_1281);
nor U1568 (N_1568,N_1172,In_2224);
xnor U1569 (N_1569,N_138,N_1256);
and U1570 (N_1570,N_1050,N_1040);
or U1571 (N_1571,N_689,N_761);
nor U1572 (N_1572,N_825,N_1322);
xor U1573 (N_1573,In_2452,In_497);
nor U1574 (N_1574,N_1312,N_942);
nor U1575 (N_1575,N_1147,In_1309);
nor U1576 (N_1576,N_1202,N_113);
nor U1577 (N_1577,N_814,N_1237);
xnor U1578 (N_1578,N_812,In_890);
nor U1579 (N_1579,In_1863,In_1664);
nand U1580 (N_1580,In_2061,N_1033);
xor U1581 (N_1581,In_2133,N_827);
or U1582 (N_1582,In_193,N_906);
nor U1583 (N_1583,In_2472,N_898);
xnor U1584 (N_1584,N_734,N_589);
xor U1585 (N_1585,In_957,In_831);
or U1586 (N_1586,N_552,In_383);
or U1587 (N_1587,N_84,N_278);
and U1588 (N_1588,In_2295,In_387);
and U1589 (N_1589,N_1324,N_172);
or U1590 (N_1590,In_542,N_967);
or U1591 (N_1591,In_1967,In_400);
and U1592 (N_1592,N_676,In_2466);
and U1593 (N_1593,N_1362,N_464);
xnor U1594 (N_1594,N_925,N_602);
nand U1595 (N_1595,N_1075,N_691);
nor U1596 (N_1596,N_511,N_1077);
xor U1597 (N_1597,N_892,N_877);
nor U1598 (N_1598,In_2139,N_1382);
or U1599 (N_1599,N_403,In_361);
or U1600 (N_1600,N_1030,N_1563);
xnor U1601 (N_1601,In_761,N_1374);
or U1602 (N_1602,N_1460,In_2214);
and U1603 (N_1603,N_1541,N_1056);
nand U1604 (N_1604,In_1706,In_1528);
nand U1605 (N_1605,In_108,N_965);
or U1606 (N_1606,N_365,N_1310);
nand U1607 (N_1607,N_914,N_1420);
nand U1608 (N_1608,N_1100,In_1277);
or U1609 (N_1609,N_897,N_798);
nor U1610 (N_1610,In_1522,N_1339);
or U1611 (N_1611,N_711,N_1502);
nor U1612 (N_1612,In_1523,N_1278);
nand U1613 (N_1613,In_1766,N_1466);
nor U1614 (N_1614,N_1047,In_924);
xnor U1615 (N_1615,N_1069,N_832);
xnor U1616 (N_1616,N_777,N_1537);
nand U1617 (N_1617,N_612,In_587);
nor U1618 (N_1618,N_780,N_896);
nand U1619 (N_1619,N_1488,In_727);
xor U1620 (N_1620,In_947,N_1404);
or U1621 (N_1621,N_640,In_1024);
and U1622 (N_1622,N_1084,N_1363);
nor U1623 (N_1623,In_211,N_993);
nor U1624 (N_1624,N_1180,N_1448);
nor U1625 (N_1625,N_653,N_491);
or U1626 (N_1626,N_1115,N_305);
nor U1627 (N_1627,In_667,N_643);
or U1628 (N_1628,N_101,N_729);
nor U1629 (N_1629,N_839,N_1487);
and U1630 (N_1630,N_1449,N_631);
nand U1631 (N_1631,N_1475,N_915);
and U1632 (N_1632,N_1242,N_1371);
nand U1633 (N_1633,N_177,N_890);
nor U1634 (N_1634,N_1419,N_1392);
xnor U1635 (N_1635,In_2379,N_1582);
xor U1636 (N_1636,N_308,N_1293);
nor U1637 (N_1637,In_1950,N_1298);
nand U1638 (N_1638,In_902,N_336);
or U1639 (N_1639,N_3,N_1430);
nand U1640 (N_1640,N_992,N_1003);
xnor U1641 (N_1641,In_1811,In_1892);
and U1642 (N_1642,N_1405,N_894);
xnor U1643 (N_1643,N_1511,N_1243);
nor U1644 (N_1644,N_280,In_2488);
nand U1645 (N_1645,N_1082,N_569);
xnor U1646 (N_1646,N_1004,N_315);
or U1647 (N_1647,N_450,N_1568);
nand U1648 (N_1648,N_715,N_1571);
and U1649 (N_1649,In_28,N_1230);
xor U1650 (N_1650,In_29,N_397);
and U1651 (N_1651,N_1552,N_904);
xor U1652 (N_1652,N_1275,N_937);
and U1653 (N_1653,N_1221,N_265);
or U1654 (N_1654,In_2122,N_725);
nor U1655 (N_1655,N_1158,N_504);
and U1656 (N_1656,N_540,N_1592);
nor U1657 (N_1657,N_1029,In_55);
and U1658 (N_1658,N_1226,N_1547);
or U1659 (N_1659,N_1578,N_425);
nor U1660 (N_1660,N_861,In_826);
and U1661 (N_1661,N_1022,In_1527);
nand U1662 (N_1662,N_1296,N_1489);
xnor U1663 (N_1663,N_199,N_205);
nor U1664 (N_1664,N_1364,N_747);
xor U1665 (N_1665,N_1425,N_1523);
nor U1666 (N_1666,N_180,N_1512);
and U1667 (N_1667,In_1961,N_1470);
nand U1668 (N_1668,N_782,N_1212);
or U1669 (N_1669,N_1257,In_421);
and U1670 (N_1670,In_816,N_1253);
xor U1671 (N_1671,N_887,N_153);
xor U1672 (N_1672,N_1129,N_953);
or U1673 (N_1673,N_1187,N_1444);
nor U1674 (N_1674,N_1427,In_416);
or U1675 (N_1675,N_296,N_411);
and U1676 (N_1676,N_1028,N_981);
nor U1677 (N_1677,In_1484,N_409);
and U1678 (N_1678,In_2387,In_1038);
or U1679 (N_1679,N_16,In_312);
or U1680 (N_1680,N_1588,N_1483);
or U1681 (N_1681,N_1406,N_885);
nor U1682 (N_1682,N_1498,N_706);
nand U1683 (N_1683,N_1196,N_1055);
nand U1684 (N_1684,N_1123,N_1534);
and U1685 (N_1685,In_1916,In_979);
nor U1686 (N_1686,N_1,In_426);
nor U1687 (N_1687,N_1551,N_1232);
xor U1688 (N_1688,In_790,In_24);
nor U1689 (N_1689,N_1140,N_306);
xnor U1690 (N_1690,N_1037,N_1564);
nand U1691 (N_1691,N_1376,In_1455);
nand U1692 (N_1692,In_1656,N_943);
or U1693 (N_1693,N_601,N_1328);
xor U1694 (N_1694,N_1355,N_1189);
nand U1695 (N_1695,N_1235,N_1124);
or U1696 (N_1696,N_675,N_100);
nand U1697 (N_1697,N_159,N_1591);
xor U1698 (N_1698,N_1538,N_509);
or U1699 (N_1699,N_648,In_1530);
or U1700 (N_1700,N_1244,In_2086);
nand U1701 (N_1701,In_52,In_895);
nor U1702 (N_1702,In_2460,N_459);
or U1703 (N_1703,N_1456,N_1350);
nand U1704 (N_1704,N_750,N_1252);
nand U1705 (N_1705,N_309,In_1667);
and U1706 (N_1706,N_870,N_1435);
xnor U1707 (N_1707,N_664,N_1527);
xnor U1708 (N_1708,N_1268,In_1532);
and U1709 (N_1709,N_1440,N_1391);
nor U1710 (N_1710,N_1453,N_1424);
nor U1711 (N_1711,N_1482,N_1545);
and U1712 (N_1712,In_540,N_1583);
nand U1713 (N_1713,N_679,In_412);
xor U1714 (N_1714,N_1289,N_1072);
or U1715 (N_1715,N_1356,N_1201);
nor U1716 (N_1716,N_829,In_2001);
xor U1717 (N_1717,In_936,N_995);
xor U1718 (N_1718,N_1365,N_941);
or U1719 (N_1719,N_1370,N_1254);
xnor U1720 (N_1720,N_1149,In_1642);
nor U1721 (N_1721,In_1481,N_515);
and U1722 (N_1722,N_1273,In_1659);
nand U1723 (N_1723,In_1223,N_438);
nor U1724 (N_1724,In_2457,N_658);
nand U1725 (N_1725,In_808,N_1279);
nor U1726 (N_1726,N_736,N_1245);
xnor U1727 (N_1727,In_1959,N_1255);
or U1728 (N_1728,In_2260,N_1372);
nand U1729 (N_1729,N_1509,N_1585);
xnor U1730 (N_1730,N_1446,N_463);
and U1731 (N_1731,N_1353,In_2267);
or U1732 (N_1732,N_1461,N_1457);
and U1733 (N_1733,N_1284,N_555);
or U1734 (N_1734,N_1491,In_1975);
nand U1735 (N_1735,N_790,N_1418);
or U1736 (N_1736,N_1134,N_972);
or U1737 (N_1737,N_1286,N_1576);
nand U1738 (N_1738,N_801,N_1479);
nand U1739 (N_1739,In_206,N_1384);
xnor U1740 (N_1740,In_619,In_1295);
nand U1741 (N_1741,N_206,N_1525);
xnor U1742 (N_1742,N_831,In_1081);
nor U1743 (N_1743,In_1280,N_1472);
or U1744 (N_1744,N_713,N_1215);
xnor U1745 (N_1745,In_2324,N_1323);
nand U1746 (N_1746,N_822,N_1316);
and U1747 (N_1747,N_1086,N_616);
and U1748 (N_1748,N_1015,N_65);
nand U1749 (N_1749,N_1351,In_2201);
xnor U1750 (N_1750,In_1462,In_1452);
or U1751 (N_1751,In_886,N_946);
and U1752 (N_1752,N_1478,In_284);
nor U1753 (N_1753,N_1346,N_56);
nor U1754 (N_1754,N_1493,N_354);
nand U1755 (N_1755,N_1439,N_157);
or U1756 (N_1756,In_2193,N_1510);
or U1757 (N_1757,In_395,N_279);
or U1758 (N_1758,In_2221,N_119);
or U1759 (N_1759,N_203,N_1540);
or U1760 (N_1760,In_212,N_1349);
or U1761 (N_1761,In_799,N_952);
xnor U1762 (N_1762,N_1451,N_1549);
xor U1763 (N_1763,N_855,In_938);
nor U1764 (N_1764,N_1403,In_348);
and U1765 (N_1765,N_1560,In_315);
xnor U1766 (N_1766,N_1599,N_971);
or U1767 (N_1767,N_1063,N_1565);
and U1768 (N_1768,N_1145,N_1501);
nand U1769 (N_1769,N_1495,N_1238);
and U1770 (N_1770,N_1468,N_1569);
and U1771 (N_1771,In_1765,N_1492);
nand U1772 (N_1772,N_1036,N_710);
or U1773 (N_1773,N_1412,N_1447);
or U1774 (N_1774,N_178,N_1378);
nor U1775 (N_1775,In_738,In_225);
nor U1776 (N_1776,In_1478,N_1400);
and U1777 (N_1777,N_232,N_1021);
xnor U1778 (N_1778,N_1450,N_1575);
xor U1779 (N_1779,N_1299,N_1445);
xor U1780 (N_1780,N_1218,N_1413);
or U1781 (N_1781,N_1026,In_2217);
nor U1782 (N_1782,In_1921,N_1441);
xor U1783 (N_1783,N_1520,N_760);
xnor U1784 (N_1784,N_843,N_1584);
or U1785 (N_1785,N_477,N_1329);
nand U1786 (N_1786,In_1928,In_1996);
xnor U1787 (N_1787,N_923,N_1352);
or U1788 (N_1788,N_1343,N_816);
nor U1789 (N_1789,N_1007,In_631);
or U1790 (N_1790,N_731,N_1422);
nand U1791 (N_1791,In_1003,N_1513);
nor U1792 (N_1792,N_781,N_880);
or U1793 (N_1793,N_1476,In_334);
or U1794 (N_1794,N_785,N_813);
or U1795 (N_1795,N_730,N_1068);
xnor U1796 (N_1796,N_1485,N_1319);
nor U1797 (N_1797,In_544,N_1436);
and U1798 (N_1798,N_1379,N_1521);
nand U1799 (N_1799,N_863,In_701);
or U1800 (N_1800,N_1083,N_716);
nor U1801 (N_1801,In_2185,N_1579);
xor U1802 (N_1802,N_1557,In_852);
or U1803 (N_1803,In_1907,N_1471);
or U1804 (N_1804,In_224,N_786);
and U1805 (N_1805,N_1225,N_1546);
xnor U1806 (N_1806,N_1309,In_894);
or U1807 (N_1807,N_1683,N_1707);
nand U1808 (N_1808,N_1740,N_1177);
nand U1809 (N_1809,N_1013,N_1613);
or U1810 (N_1810,N_1183,N_1503);
and U1811 (N_1811,N_1553,N_1515);
xor U1812 (N_1812,In_296,N_1542);
or U1813 (N_1813,N_1632,N_1369);
nand U1814 (N_1814,N_446,In_1754);
xor U1815 (N_1815,In_1614,N_1768);
nand U1816 (N_1816,In_2485,N_1651);
or U1817 (N_1817,N_1277,In_2266);
nor U1818 (N_1818,N_1780,N_773);
nor U1819 (N_1819,N_987,N_1302);
nor U1820 (N_1820,N_960,N_1301);
or U1821 (N_1821,N_633,N_1516);
nand U1822 (N_1822,In_1307,N_847);
xor U1823 (N_1823,N_1174,In_2158);
nand U1824 (N_1824,In_1957,In_1946);
nand U1825 (N_1825,N_1721,N_383);
xor U1826 (N_1826,N_1500,N_1023);
nand U1827 (N_1827,In_2198,N_359);
xor U1828 (N_1828,N_1397,N_1442);
nor U1829 (N_1829,N_1656,N_1267);
nand U1830 (N_1830,N_115,N_527);
nand U1831 (N_1831,N_771,In_423);
nand U1832 (N_1832,In_2203,N_970);
or U1833 (N_1833,N_1094,N_876);
xnor U1834 (N_1834,N_1672,N_1473);
and U1835 (N_1835,In_669,N_1711);
nand U1836 (N_1836,In_1595,N_1775);
nor U1837 (N_1837,In_1806,N_391);
nor U1838 (N_1838,N_1411,In_1383);
nand U1839 (N_1839,N_1753,N_651);
xor U1840 (N_1840,N_1739,In_2428);
or U1841 (N_1841,N_1517,In_147);
nand U1842 (N_1842,In_301,N_1629);
nor U1843 (N_1843,N_408,In_2130);
or U1844 (N_1844,In_1984,N_1716);
or U1845 (N_1845,N_1556,N_841);
nor U1846 (N_1846,N_1606,N_1587);
nand U1847 (N_1847,In_2218,N_358);
xnor U1848 (N_1848,N_1344,N_1562);
nor U1849 (N_1849,N_1706,N_1595);
nor U1850 (N_1850,In_2024,N_1535);
xor U1851 (N_1851,In_1367,N_1386);
nand U1852 (N_1852,In_1648,N_1477);
xnor U1853 (N_1853,N_26,N_1251);
nand U1854 (N_1854,In_1446,N_1610);
or U1855 (N_1855,N_1720,N_1778);
or U1856 (N_1856,N_1624,In_1814);
or U1857 (N_1857,In_469,N_1717);
or U1858 (N_1858,N_1709,N_990);
xnor U1859 (N_1859,N_1745,N_1496);
and U1860 (N_1860,In_311,N_1596);
nand U1861 (N_1861,N_1335,N_1288);
nor U1862 (N_1862,N_1662,N_1667);
or U1863 (N_1863,N_1438,N_1506);
xor U1864 (N_1864,N_1737,N_1233);
or U1865 (N_1865,N_1715,N_1558);
xnor U1866 (N_1866,N_1608,N_1152);
or U1867 (N_1867,In_2028,N_1710);
xnor U1868 (N_1868,N_755,In_1127);
nand U1869 (N_1869,N_1761,N_1340);
or U1870 (N_1870,N_1734,N_1049);
nand U1871 (N_1871,N_1570,N_1795);
nor U1872 (N_1872,N_1698,N_1642);
nand U1873 (N_1873,N_1671,N_332);
nand U1874 (N_1874,N_1661,N_1532);
nor U1875 (N_1875,N_1722,In_1914);
nand U1876 (N_1876,N_1519,N_1682);
nand U1877 (N_1877,In_1713,N_1742);
or U1878 (N_1878,In_1343,N_1636);
nand U1879 (N_1879,N_1670,N_1758);
nor U1880 (N_1880,N_1793,N_1046);
xor U1881 (N_1881,N_1104,N_1518);
nor U1882 (N_1882,N_1227,N_1623);
nor U1883 (N_1883,N_1408,In_1804);
nand U1884 (N_1884,In_1608,N_1748);
and U1885 (N_1885,In_844,N_355);
or U1886 (N_1886,N_977,N_1689);
nand U1887 (N_1887,N_1153,In_493);
and U1888 (N_1888,N_454,N_1409);
nor U1889 (N_1889,N_1799,N_1645);
and U1890 (N_1890,In_1729,N_490);
nor U1891 (N_1891,In_2484,N_1210);
nand U1892 (N_1892,In_351,N_1770);
or U1893 (N_1893,N_874,N_1401);
xor U1894 (N_1894,N_1702,N_908);
or U1895 (N_1895,N_1431,N_1462);
or U1896 (N_1896,N_1674,N_1416);
and U1897 (N_1897,N_1607,N_1787);
xor U1898 (N_1898,N_1704,N_917);
or U1899 (N_1899,N_1529,N_1773);
or U1900 (N_1900,N_999,N_1474);
xor U1901 (N_1901,N_1393,N_1359);
and U1902 (N_1902,N_1687,N_1025);
nand U1903 (N_1903,N_844,N_1679);
nor U1904 (N_1904,N_1605,N_1732);
nand U1905 (N_1905,N_1347,N_1566);
xnor U1906 (N_1906,N_1263,N_158);
and U1907 (N_1907,N_647,N_1789);
and U1908 (N_1908,N_1628,N_1728);
or U1909 (N_1909,In_1932,N_724);
xnor U1910 (N_1910,N_1220,N_468);
xor U1911 (N_1911,N_1714,N_1703);
or U1912 (N_1912,In_2342,N_1602);
and U1913 (N_1913,N_1784,N_1598);
nor U1914 (N_1914,N_1572,N_1373);
nor U1915 (N_1915,N_478,N_1712);
and U1916 (N_1916,N_1423,N_1590);
nand U1917 (N_1917,N_796,N_1643);
nand U1918 (N_1918,N_1655,In_632);
and U1919 (N_1919,N_1348,N_213);
or U1920 (N_1920,N_718,N_1733);
nand U1921 (N_1921,N_1294,N_1426);
and U1922 (N_1922,In_1357,N_1637);
nand U1923 (N_1923,N_1250,In_2240);
xnor U1924 (N_1924,N_673,In_593);
nand U1925 (N_1925,N_299,N_1266);
and U1926 (N_1926,N_768,In_1294);
nand U1927 (N_1927,N_539,N_1274);
and U1928 (N_1928,N_1586,In_1593);
xnor U1929 (N_1929,In_181,In_1046);
and U1930 (N_1930,N_1368,N_1459);
and U1931 (N_1931,N_1619,N_1783);
nor U1932 (N_1932,N_1724,N_1731);
or U1933 (N_1933,N_1735,N_1781);
or U1934 (N_1934,N_1467,N_1615);
nand U1935 (N_1935,N_1776,N_1291);
nor U1936 (N_1936,N_1200,N_1016);
nor U1937 (N_1937,N_1719,N_493);
nor U1938 (N_1938,N_1308,In_318);
and U1939 (N_1939,N_985,In_1208);
and U1940 (N_1940,N_1214,N_1622);
nor U1941 (N_1941,N_1484,N_1306);
or U1942 (N_1942,N_1785,N_67);
nand U1943 (N_1943,N_1524,In_1988);
xnor U1944 (N_1944,N_1749,N_693);
nand U1945 (N_1945,N_1648,N_592);
or U1946 (N_1946,N_1691,N_1759);
nor U1947 (N_1947,N_122,In_608);
nand U1948 (N_1948,N_1318,N_1051);
nand U1949 (N_1949,In_2093,N_1248);
xor U1950 (N_1950,N_1499,In_37);
xor U1951 (N_1951,In_611,N_669);
and U1952 (N_1952,N_963,N_1762);
xnor U1953 (N_1953,N_398,N_1580);
or U1954 (N_1954,N_1292,N_1641);
nor U1955 (N_1955,N_176,N_922);
or U1956 (N_1956,N_1490,In_1526);
xor U1957 (N_1957,N_1646,N_1164);
xnor U1958 (N_1958,N_285,N_1415);
and U1959 (N_1959,N_1258,N_1633);
xor U1960 (N_1960,N_1531,N_1103);
or U1961 (N_1961,N_1685,In_1104);
nor U1962 (N_1962,N_14,In_1285);
xnor U1963 (N_1963,N_1750,In_882);
nand U1964 (N_1964,N_1574,In_1848);
and U1965 (N_1965,N_1561,N_1688);
xor U1966 (N_1966,N_1443,N_1696);
nand U1967 (N_1967,N_753,N_984);
or U1968 (N_1968,In_1394,N_666);
or U1969 (N_1969,N_1236,N_978);
xor U1970 (N_1970,N_1059,N_374);
xor U1971 (N_1971,In_734,N_1790);
nor U1972 (N_1972,N_1543,In_102);
nand U1973 (N_1973,N_1398,In_1850);
nand U1974 (N_1974,N_1464,N_1539);
or U1975 (N_1975,N_1452,N_1006);
nand U1976 (N_1976,In_1155,In_2317);
and U1977 (N_1977,In_621,N_1777);
nand U1978 (N_1978,N_656,In_1919);
or U1979 (N_1979,N_576,N_1011);
xor U1980 (N_1980,N_1746,N_91);
xor U1981 (N_1981,N_1494,N_1331);
nand U1982 (N_1982,In_1609,N_1211);
nor U1983 (N_1983,In_1293,N_433);
and U1984 (N_1984,N_1508,N_220);
and U1985 (N_1985,N_1727,In_865);
nor U1986 (N_1986,N_1481,N_776);
xnor U1987 (N_1987,N_1465,N_1635);
and U1988 (N_1988,N_1664,In_907);
and U1989 (N_1989,In_1260,In_127);
xor U1990 (N_1990,N_1765,N_921);
xnor U1991 (N_1991,N_1625,In_2141);
xor U1992 (N_1992,N_1763,N_1796);
nand U1993 (N_1993,N_697,N_1402);
and U1994 (N_1994,N_1361,N_1695);
nor U1995 (N_1995,N_1603,N_1612);
and U1996 (N_1996,N_698,N_1264);
nand U1997 (N_1997,N_1486,N_1536);
or U1998 (N_1998,In_1049,N_1208);
xnor U1999 (N_1999,N_687,In_12);
xnor U2000 (N_2000,N_1814,In_2294);
nor U2001 (N_2001,N_1868,N_1387);
and U2002 (N_2002,In_1678,In_1652);
nand U2003 (N_2003,N_1862,N_1887);
xnor U2004 (N_2004,N_1844,N_1332);
nand U2005 (N_2005,N_1910,N_1774);
or U2006 (N_2006,N_1936,N_1756);
nor U2007 (N_2007,N_621,N_1895);
and U2008 (N_2008,N_1897,N_931);
xor U2009 (N_2009,N_1979,N_1974);
nand U2010 (N_2010,N_1019,N_1757);
xor U2011 (N_2011,N_1262,N_1548);
and U2012 (N_2012,N_1769,N_1829);
nor U2013 (N_2013,N_1680,N_1810);
nand U2014 (N_2014,N_1533,N_1822);
nor U2015 (N_2015,N_1530,N_1937);
nand U2016 (N_2016,N_1754,N_1911);
and U2017 (N_2017,In_1061,N_1848);
or U2018 (N_2018,N_705,N_1295);
nor U2019 (N_2019,N_1281,N_1871);
nor U2020 (N_2020,N_1960,N_1863);
nand U2021 (N_2021,N_7,In_462);
xnor U2022 (N_2022,N_1806,N_1882);
nor U2023 (N_2023,N_1866,N_1938);
nor U2024 (N_2024,N_1701,N_1760);
or U2025 (N_2025,N_1300,N_1877);
nor U2026 (N_2026,N_1729,N_1944);
and U2027 (N_2027,N_1983,In_2177);
or U2028 (N_2028,N_1581,N_1808);
xnor U2029 (N_2029,N_1311,N_1157);
nor U2030 (N_2030,N_1060,In_112);
and U2031 (N_2031,N_1692,N_1678);
or U2032 (N_2032,N_1676,N_364);
xnor U2033 (N_2033,N_1992,N_1994);
nand U2034 (N_2034,N_1920,N_1577);
xor U2035 (N_2035,N_1893,N_1803);
or U2036 (N_2036,N_1074,In_2156);
nand U2037 (N_2037,N_1961,N_837);
xnor U2038 (N_2038,N_1809,N_1684);
nand U2039 (N_2039,N_1821,N_1838);
or U2040 (N_2040,N_1982,N_1993);
and U2041 (N_2041,In_1440,In_2110);
nand U2042 (N_2042,N_1800,N_948);
nor U2043 (N_2043,N_1755,N_594);
and U2044 (N_2044,N_1747,N_1169);
xor U2045 (N_2045,N_1969,N_1855);
or U2046 (N_2046,N_1971,In_1234);
nand U2047 (N_2047,N_1366,In_473);
and U2048 (N_2048,N_1978,N_1942);
nand U2049 (N_2049,N_1782,N_1428);
and U2050 (N_2050,N_1660,N_1797);
xnor U2051 (N_2051,N_1432,N_1178);
xnor U2052 (N_2052,N_1338,N_1952);
nand U2053 (N_2053,N_1883,In_951);
nor U2054 (N_2054,N_1935,N_1835);
nor U2055 (N_2055,N_1395,In_175);
and U2056 (N_2056,N_1909,In_1321);
nor U2057 (N_2057,N_1407,N_1843);
nor U2058 (N_2058,N_1550,N_1980);
xor U2059 (N_2059,In_1625,N_751);
nand U2060 (N_2060,N_1997,N_1738);
or U2061 (N_2061,N_466,N_1555);
xnor U2062 (N_2062,N_1954,In_1802);
nand U2063 (N_2063,In_988,N_1975);
xnor U2064 (N_2064,N_1906,N_1878);
nand U2065 (N_2065,N_1833,N_1928);
nor U2066 (N_2066,N_888,In_2476);
or U2067 (N_2067,N_1889,N_1647);
or U2068 (N_2068,N_1959,N_1963);
or U2069 (N_2069,N_1693,N_1973);
nor U2070 (N_2070,N_1052,N_1946);
xor U2071 (N_2071,N_1792,N_1815);
nand U2072 (N_2072,In_2278,N_1681);
or U2073 (N_2073,N_1805,N_787);
and U2074 (N_2074,N_1675,N_1842);
nor U2075 (N_2075,N_1528,N_1864);
xnor U2076 (N_2076,N_1410,N_1247);
and U2077 (N_2077,N_1144,N_1652);
xor U2078 (N_2078,In_371,N_1102);
or U2079 (N_2079,N_1654,N_1955);
xor U2080 (N_2080,In_2369,N_1358);
and U2081 (N_2081,N_1726,N_1522);
or U2082 (N_2082,N_1690,N_1417);
nand U2083 (N_2083,N_1907,N_1986);
and U2084 (N_2084,N_1890,N_1939);
nand U2085 (N_2085,N_1970,N_1836);
or U2086 (N_2086,N_1988,N_738);
and U2087 (N_2087,N_1898,In_1326);
or U2088 (N_2088,N_1665,N_1996);
or U2089 (N_2089,N_1497,N_1966);
xor U2090 (N_2090,N_1597,N_1618);
and U2091 (N_2091,N_1976,N_867);
nor U2092 (N_2092,N_905,N_1837);
or U2093 (N_2093,N_1859,N_1856);
or U2094 (N_2094,N_1891,N_1850);
xnor U2095 (N_2095,In_2207,N_1705);
xnor U2096 (N_2096,N_1314,N_1653);
or U2097 (N_2097,N_1616,N_1206);
nand U2098 (N_2098,N_1626,N_1337);
xnor U2099 (N_2099,In_724,N_1823);
xor U2100 (N_2100,N_1901,N_1224);
or U2101 (N_2101,N_1609,N_1853);
xnor U2102 (N_2102,N_1991,In_969);
and U2103 (N_2103,N_1725,N_1811);
or U2104 (N_2104,In_1117,N_1611);
nand U2105 (N_2105,N_1638,In_2345);
nand U2106 (N_2106,N_1819,N_1865);
nand U2107 (N_2107,N_1567,In_1308);
or U2108 (N_2108,N_1505,N_1896);
nand U2109 (N_2109,N_1791,N_1458);
nand U2110 (N_2110,N_551,N_872);
xor U2111 (N_2111,N_1507,N_856);
xor U2112 (N_2112,N_1285,N_1977);
xor U2113 (N_2113,In_46,N_1916);
or U2114 (N_2114,N_1873,N_390);
nand U2115 (N_2115,N_1779,N_1269);
xnor U2116 (N_2116,N_1950,N_1989);
nor U2117 (N_2117,N_1824,In_2375);
nor U2118 (N_2118,N_487,N_1852);
nor U2119 (N_2119,N_1964,N_1383);
and U2120 (N_2120,N_1744,N_1919);
or U2121 (N_2121,N_1801,N_1669);
nor U2122 (N_2122,N_1925,N_1699);
and U2123 (N_2123,N_958,N_64);
nand U2124 (N_2124,N_1908,N_1767);
or U2125 (N_2125,N_1817,In_1015);
or U2126 (N_2126,N_1930,N_1903);
nor U2127 (N_2127,N_1990,N_1870);
and U2128 (N_2128,N_1650,N_1594);
xnor U2129 (N_2129,N_1984,N_1336);
and U2130 (N_2130,N_1804,In_1696);
and U2131 (N_2131,N_930,N_1621);
xnor U2132 (N_2132,N_1867,N_1934);
nand U2133 (N_2133,In_63,N_1958);
nor U2134 (N_2134,N_1668,N_815);
or U2135 (N_2135,N_1825,N_1924);
xnor U2136 (N_2136,N_1700,N_1469);
nand U2137 (N_2137,N_1968,N_1697);
or U2138 (N_2138,N_1627,In_571);
nor U2139 (N_2139,N_1957,N_1839);
nand U2140 (N_2140,N_1434,N_1433);
nand U2141 (N_2141,In_1270,N_966);
or U2142 (N_2142,N_1663,N_1287);
nor U2143 (N_2143,N_1718,N_1949);
nand U2144 (N_2144,N_1858,N_1751);
and U2145 (N_2145,N_1604,N_1846);
nor U2146 (N_2146,N_1631,N_1283);
nand U2147 (N_2147,N_1559,N_1694);
nor U2148 (N_2148,N_1813,In_932);
nand U2149 (N_2149,N_1723,In_860);
or U2150 (N_2150,N_1857,N_1480);
and U2151 (N_2151,N_173,N_1644);
nor U2152 (N_2152,N_1341,N_1617);
or U2153 (N_2153,N_920,N_1788);
xor U2154 (N_2154,N_1657,N_1686);
and U2155 (N_2155,In_47,N_1912);
xnor U2156 (N_2156,In_536,N_1173);
nand U2157 (N_2157,N_1941,N_1771);
or U2158 (N_2158,N_484,N_167);
and U2159 (N_2159,N_903,In_267);
xnor U2160 (N_2160,N_396,N_1947);
xor U2161 (N_2161,In_130,N_1929);
xor U2162 (N_2162,N_756,N_1713);
or U2163 (N_2163,N_1320,N_1544);
nand U2164 (N_2164,In_2044,N_1831);
nor U2165 (N_2165,N_1965,N_1260);
nand U2166 (N_2166,In_901,N_1830);
xor U2167 (N_2167,N_1807,N_1786);
or U2168 (N_2168,N_1847,N_1640);
or U2169 (N_2169,N_1554,N_1828);
nor U2170 (N_2170,N_1869,In_933);
and U2171 (N_2171,N_1948,N_1927);
xnor U2172 (N_2172,N_1325,In_344);
xnor U2173 (N_2173,N_1854,N_1881);
nor U2174 (N_2174,N_1673,N_1454);
and U2175 (N_2175,N_1381,N_1818);
nand U2176 (N_2176,In_627,N_1940);
and U2177 (N_2177,N_1526,In_377);
xor U2178 (N_2178,In_909,N_1943);
xnor U2179 (N_2179,N_1752,N_1884);
nand U2180 (N_2180,N_1455,N_1614);
nor U2181 (N_2181,N_1845,N_1630);
nand U2182 (N_2182,N_1832,N_1107);
nand U2183 (N_2183,N_1708,N_1851);
or U2184 (N_2184,In_3,In_41);
or U2185 (N_2185,N_1923,N_1914);
or U2186 (N_2186,In_1553,N_1921);
and U2187 (N_2187,N_1860,In_1225);
xor U2188 (N_2188,N_1956,N_208);
nor U2189 (N_2189,N_1834,N_1303);
and U2190 (N_2190,N_1234,N_1894);
and U2191 (N_2191,In_2411,N_1972);
or U2192 (N_2192,N_1634,N_1649);
xnor U2193 (N_2193,N_1926,N_1967);
and U2194 (N_2194,N_1879,In_300);
and U2195 (N_2195,N_1593,N_1874);
nor U2196 (N_2196,N_1917,N_817);
nand U2197 (N_2197,N_1981,N_1812);
nand U2198 (N_2198,N_1933,N_1945);
or U2199 (N_2199,In_247,In_2315);
nor U2200 (N_2200,N_1053,In_2388);
and U2201 (N_2201,N_2114,N_2182);
nor U2202 (N_2202,N_2158,N_2023);
nand U2203 (N_2203,In_277,N_2199);
or U2204 (N_2204,In_1322,N_2197);
and U2205 (N_2205,N_2170,N_2044);
or U2206 (N_2206,N_1902,N_2069);
xnor U2207 (N_2207,In_1095,N_2147);
nor U2208 (N_2208,N_2176,N_2110);
or U2209 (N_2209,In_1744,N_2077);
and U2210 (N_2210,N_2057,In_2292);
and U2211 (N_2211,N_2174,N_2108);
and U2212 (N_2212,N_1899,N_2053);
xnor U2213 (N_2213,N_1743,N_2072);
xor U2214 (N_2214,N_2055,N_2193);
nand U2215 (N_2215,In_1401,N_2092);
xnor U2216 (N_2216,N_1573,N_2076);
and U2217 (N_2217,N_2152,N_2084);
xor U2218 (N_2218,N_1962,N_2156);
nand U2219 (N_2219,N_2121,N_1658);
and U2220 (N_2220,N_1932,N_2062);
and U2221 (N_2221,N_2085,N_2141);
and U2222 (N_2222,N_2154,N_2097);
or U2223 (N_2223,N_2058,N_2167);
xnor U2224 (N_2224,N_1918,N_2031);
or U2225 (N_2225,N_2127,N_2074);
nand U2226 (N_2226,N_2187,N_2148);
xnor U2227 (N_2227,N_242,N_2020);
or U2228 (N_2228,N_1904,N_2136);
or U2229 (N_2229,N_2011,N_1024);
nand U2230 (N_2230,N_2088,N_1985);
and U2231 (N_2231,In_1461,N_2002);
or U2232 (N_2232,N_2063,In_1574);
and U2233 (N_2233,N_1437,N_1730);
nor U2234 (N_2234,N_2161,N_1414);
or U2235 (N_2235,N_2090,N_2185);
xnor U2236 (N_2236,N_2151,N_1999);
and U2237 (N_2237,N_1915,N_2105);
xor U2238 (N_2238,N_2032,N_2071);
or U2239 (N_2239,N_2086,N_2033);
nand U2240 (N_2240,N_2022,N_802);
or U2241 (N_2241,N_2096,N_2171);
and U2242 (N_2242,N_2164,N_2146);
nor U2243 (N_2243,N_1659,N_2054);
and U2244 (N_2244,N_2101,N_2080);
xor U2245 (N_2245,N_2131,N_2112);
nor U2246 (N_2246,N_2021,N_2006);
nand U2247 (N_2247,N_2034,N_2042);
and U2248 (N_2248,N_2153,N_2029);
nor U2249 (N_2249,N_2192,N_2107);
nand U2250 (N_2250,N_2132,N_2070);
nor U2251 (N_2251,N_2130,N_2001);
nor U2252 (N_2252,N_804,N_2091);
nor U2253 (N_2253,N_2026,N_2135);
or U2254 (N_2254,N_2037,N_1892);
and U2255 (N_2255,N_1772,N_2049);
nor U2256 (N_2256,N_2196,N_2036);
xnor U2257 (N_2257,N_1032,N_1620);
nand U2258 (N_2258,N_1000,N_2133);
or U2259 (N_2259,N_1099,N_2004);
nor U2260 (N_2260,N_2051,N_2015);
nor U2261 (N_2261,N_1085,N_1995);
and U2262 (N_2262,N_1088,N_2012);
or U2263 (N_2263,N_2067,N_1639);
nand U2264 (N_2264,N_2082,N_2129);
or U2265 (N_2265,N_1816,N_2188);
xor U2266 (N_2266,N_2104,N_1589);
and U2267 (N_2267,N_2000,N_2008);
and U2268 (N_2268,N_2050,N_2079);
nor U2269 (N_2269,N_1888,N_1876);
or U2270 (N_2270,N_2066,N_2005);
nand U2271 (N_2271,N_2128,N_2116);
xnor U2272 (N_2272,N_1076,N_2035);
and U2273 (N_2273,N_2125,N_2115);
nor U2274 (N_2274,N_2138,N_2043);
xor U2275 (N_2275,N_1886,N_2065);
nor U2276 (N_2276,N_1900,N_1861);
xor U2277 (N_2277,N_2060,N_2059);
nand U2278 (N_2278,N_2142,N_2075);
xnor U2279 (N_2279,N_2089,N_1798);
and U2280 (N_2280,In_637,N_2027);
or U2281 (N_2281,N_1125,N_2064);
nand U2282 (N_2282,N_1802,N_2040);
nor U2283 (N_2283,N_2163,N_2195);
or U2284 (N_2284,N_2109,N_1827);
or U2285 (N_2285,N_709,N_2180);
nand U2286 (N_2286,N_2157,N_1841);
or U2287 (N_2287,N_2019,N_1875);
nor U2288 (N_2288,N_1840,N_2013);
nand U2289 (N_2289,N_2048,N_2081);
xor U2290 (N_2290,N_1953,N_2179);
xor U2291 (N_2291,N_1192,N_2178);
nand U2292 (N_2292,In_461,N_2189);
and U2293 (N_2293,N_2139,N_1504);
or U2294 (N_2294,N_2083,N_1922);
or U2295 (N_2295,N_1987,N_1429);
xnor U2296 (N_2296,N_2168,N_2134);
and U2297 (N_2297,N_2198,N_2118);
and U2298 (N_2298,N_2117,N_2039);
xnor U2299 (N_2299,In_1057,N_2113);
nand U2300 (N_2300,N_1736,N_1820);
nor U2301 (N_2301,N_2093,In_1986);
nand U2302 (N_2302,N_624,N_2194);
xor U2303 (N_2303,N_2123,N_1764);
nor U2304 (N_2304,N_2052,N_553);
and U2305 (N_2305,N_2175,N_2007);
nor U2306 (N_2306,N_2102,N_2106);
or U2307 (N_2307,N_1514,N_2165);
xor U2308 (N_2308,N_2047,N_1677);
and U2309 (N_2309,In_326,N_1601);
and U2310 (N_2310,N_2137,N_1463);
or U2311 (N_2311,N_2038,N_2061);
or U2312 (N_2312,In_1955,N_1826);
xnor U2313 (N_2313,N_2166,N_1666);
or U2314 (N_2314,N_1766,N_2190);
nand U2315 (N_2315,N_2103,N_1931);
xor U2316 (N_2316,N_2172,N_1998);
nor U2317 (N_2317,N_2184,N_2119);
nor U2318 (N_2318,N_1905,N_1600);
nand U2319 (N_2319,N_2145,N_2068);
and U2320 (N_2320,N_2162,N_2159);
nor U2321 (N_2321,N_2149,N_1146);
and U2322 (N_2322,N_2150,N_2025);
and U2323 (N_2323,N_2100,N_2191);
or U2324 (N_2324,N_2173,N_2028);
and U2325 (N_2325,N_2045,N_2016);
nand U2326 (N_2326,N_1951,N_2098);
nand U2327 (N_2327,N_2056,N_2183);
nor U2328 (N_2328,N_2122,N_2126);
and U2329 (N_2329,N_2078,N_1261);
nand U2330 (N_2330,N_2120,N_2073);
and U2331 (N_2331,In_133,N_2181);
or U2332 (N_2332,N_2018,N_2030);
and U2333 (N_2333,N_1880,In_2465);
nor U2334 (N_2334,N_2099,N_597);
nand U2335 (N_2335,N_1741,N_2046);
and U2336 (N_2336,N_2014,N_2177);
and U2337 (N_2337,N_2094,N_1913);
xor U2338 (N_2338,N_2010,N_1872);
xnor U2339 (N_2339,N_2087,In_1398);
or U2340 (N_2340,N_2155,N_1885);
nor U2341 (N_2341,N_2024,N_2111);
xor U2342 (N_2342,N_2003,N_2160);
and U2343 (N_2343,N_2009,N_2144);
or U2344 (N_2344,N_2041,N_1794);
or U2345 (N_2345,N_2143,N_2017);
and U2346 (N_2346,N_1421,N_2124);
and U2347 (N_2347,N_2186,N_20);
nand U2348 (N_2348,N_1849,N_2169);
or U2349 (N_2349,N_2140,N_2095);
xor U2350 (N_2350,N_1743,N_2156);
and U2351 (N_2351,N_2150,N_2010);
nand U2352 (N_2352,N_2069,N_1888);
xor U2353 (N_2353,N_2146,N_2143);
xor U2354 (N_2354,N_2179,N_2126);
xnor U2355 (N_2355,N_2104,N_2084);
and U2356 (N_2356,N_2191,N_2142);
or U2357 (N_2357,In_326,N_2199);
nor U2358 (N_2358,N_2063,N_2153);
or U2359 (N_2359,N_2037,N_2131);
or U2360 (N_2360,N_2063,N_2172);
and U2361 (N_2361,In_637,In_1744);
and U2362 (N_2362,N_1601,N_2150);
nor U2363 (N_2363,N_2163,N_2151);
and U2364 (N_2364,N_2146,N_2142);
or U2365 (N_2365,N_2114,N_2075);
xor U2366 (N_2366,N_804,N_2055);
or U2367 (N_2367,N_2033,N_2101);
or U2368 (N_2368,N_1125,N_2168);
or U2369 (N_2369,N_597,N_709);
or U2370 (N_2370,N_2079,N_1573);
nor U2371 (N_2371,N_1076,N_2178);
xor U2372 (N_2372,N_2047,N_2042);
or U2373 (N_2373,N_2174,N_2076);
or U2374 (N_2374,N_2028,N_2099);
nor U2375 (N_2375,In_1398,N_2165);
or U2376 (N_2376,N_2023,In_1574);
and U2377 (N_2377,N_2084,N_2087);
xnor U2378 (N_2378,N_2072,N_2111);
nand U2379 (N_2379,In_1322,N_1620);
xor U2380 (N_2380,N_2116,N_1995);
or U2381 (N_2381,N_2158,N_2097);
or U2382 (N_2382,N_2056,N_2126);
nor U2383 (N_2383,N_2176,N_1816);
nor U2384 (N_2384,N_2175,N_2140);
or U2385 (N_2385,N_2146,N_1000);
nand U2386 (N_2386,N_2173,N_2146);
xor U2387 (N_2387,N_2122,N_1085);
nand U2388 (N_2388,N_2119,N_1429);
nor U2389 (N_2389,N_2130,N_2133);
or U2390 (N_2390,N_2168,N_1888);
nand U2391 (N_2391,N_2069,N_1841);
and U2392 (N_2392,N_1999,N_2008);
xor U2393 (N_2393,N_2114,N_1880);
xor U2394 (N_2394,N_2158,In_1057);
xor U2395 (N_2395,N_2142,N_2153);
nor U2396 (N_2396,N_2076,N_2083);
nor U2397 (N_2397,N_2158,N_2148);
nand U2398 (N_2398,N_2034,N_2175);
nand U2399 (N_2399,N_2189,N_2075);
nand U2400 (N_2400,N_2219,N_2235);
nand U2401 (N_2401,N_2216,N_2396);
and U2402 (N_2402,N_2316,N_2304);
or U2403 (N_2403,N_2315,N_2390);
or U2404 (N_2404,N_2207,N_2380);
xor U2405 (N_2405,N_2305,N_2352);
or U2406 (N_2406,N_2384,N_2213);
xor U2407 (N_2407,N_2287,N_2246);
and U2408 (N_2408,N_2233,N_2206);
or U2409 (N_2409,N_2342,N_2215);
nor U2410 (N_2410,N_2375,N_2203);
or U2411 (N_2411,N_2221,N_2355);
and U2412 (N_2412,N_2281,N_2383);
nand U2413 (N_2413,N_2373,N_2386);
and U2414 (N_2414,N_2266,N_2237);
and U2415 (N_2415,N_2200,N_2204);
nand U2416 (N_2416,N_2345,N_2256);
nand U2417 (N_2417,N_2269,N_2217);
xor U2418 (N_2418,N_2303,N_2369);
nand U2419 (N_2419,N_2212,N_2344);
nor U2420 (N_2420,N_2299,N_2278);
nor U2421 (N_2421,N_2318,N_2382);
and U2422 (N_2422,N_2357,N_2253);
nand U2423 (N_2423,N_2242,N_2244);
and U2424 (N_2424,N_2343,N_2261);
nand U2425 (N_2425,N_2296,N_2249);
xnor U2426 (N_2426,N_2268,N_2285);
xor U2427 (N_2427,N_2227,N_2209);
xnor U2428 (N_2428,N_2323,N_2310);
nor U2429 (N_2429,N_2363,N_2336);
and U2430 (N_2430,N_2338,N_2326);
or U2431 (N_2431,N_2291,N_2300);
and U2432 (N_2432,N_2379,N_2210);
or U2433 (N_2433,N_2302,N_2348);
or U2434 (N_2434,N_2346,N_2360);
and U2435 (N_2435,N_2341,N_2301);
and U2436 (N_2436,N_2374,N_2262);
xnor U2437 (N_2437,N_2358,N_2329);
nand U2438 (N_2438,N_2214,N_2201);
or U2439 (N_2439,N_2362,N_2255);
nand U2440 (N_2440,N_2208,N_2313);
and U2441 (N_2441,N_2337,N_2236);
xnor U2442 (N_2442,N_2378,N_2397);
xnor U2443 (N_2443,N_2259,N_2319);
xnor U2444 (N_2444,N_2391,N_2228);
nand U2445 (N_2445,N_2312,N_2321);
xor U2446 (N_2446,N_2260,N_2280);
and U2447 (N_2447,N_2317,N_2284);
xnor U2448 (N_2448,N_2271,N_2327);
and U2449 (N_2449,N_2314,N_2325);
or U2450 (N_2450,N_2340,N_2356);
nor U2451 (N_2451,N_2270,N_2250);
nand U2452 (N_2452,N_2311,N_2272);
xnor U2453 (N_2453,N_2361,N_2309);
nor U2454 (N_2454,N_2335,N_2263);
or U2455 (N_2455,N_2243,N_2395);
xor U2456 (N_2456,N_2308,N_2351);
or U2457 (N_2457,N_2251,N_2289);
nand U2458 (N_2458,N_2332,N_2222);
nor U2459 (N_2459,N_2330,N_2365);
and U2460 (N_2460,N_2224,N_2277);
nor U2461 (N_2461,N_2376,N_2241);
and U2462 (N_2462,N_2230,N_2223);
or U2463 (N_2463,N_2324,N_2388);
and U2464 (N_2464,N_2229,N_2275);
nand U2465 (N_2465,N_2385,N_2234);
nor U2466 (N_2466,N_2239,N_2245);
nand U2467 (N_2467,N_2292,N_2240);
nand U2468 (N_2468,N_2381,N_2293);
and U2469 (N_2469,N_2370,N_2307);
nand U2470 (N_2470,N_2364,N_2399);
nand U2471 (N_2471,N_2286,N_2290);
xnor U2472 (N_2472,N_2322,N_2393);
nor U2473 (N_2473,N_2353,N_2247);
or U2474 (N_2474,N_2226,N_2333);
nand U2475 (N_2475,N_2331,N_2218);
and U2476 (N_2476,N_2389,N_2220);
nand U2477 (N_2477,N_2347,N_2320);
nand U2478 (N_2478,N_2354,N_2225);
or U2479 (N_2479,N_2252,N_2306);
nand U2480 (N_2480,N_2265,N_2295);
and U2481 (N_2481,N_2254,N_2294);
or U2482 (N_2482,N_2238,N_2394);
nand U2483 (N_2483,N_2328,N_2273);
xor U2484 (N_2484,N_2339,N_2377);
xnor U2485 (N_2485,N_2367,N_2371);
xnor U2486 (N_2486,N_2298,N_2232);
nor U2487 (N_2487,N_2366,N_2372);
xnor U2488 (N_2488,N_2334,N_2288);
nand U2489 (N_2489,N_2248,N_2267);
or U2490 (N_2490,N_2359,N_2349);
nand U2491 (N_2491,N_2297,N_2257);
nand U2492 (N_2492,N_2276,N_2368);
nor U2493 (N_2493,N_2202,N_2211);
nand U2494 (N_2494,N_2264,N_2398);
nor U2495 (N_2495,N_2205,N_2231);
and U2496 (N_2496,N_2279,N_2274);
nand U2497 (N_2497,N_2387,N_2350);
nand U2498 (N_2498,N_2282,N_2283);
nand U2499 (N_2499,N_2392,N_2258);
nand U2500 (N_2500,N_2273,N_2327);
nand U2501 (N_2501,N_2268,N_2341);
nand U2502 (N_2502,N_2310,N_2347);
xnor U2503 (N_2503,N_2210,N_2250);
or U2504 (N_2504,N_2285,N_2322);
xnor U2505 (N_2505,N_2369,N_2306);
and U2506 (N_2506,N_2393,N_2235);
or U2507 (N_2507,N_2354,N_2295);
nand U2508 (N_2508,N_2211,N_2364);
xnor U2509 (N_2509,N_2275,N_2262);
nor U2510 (N_2510,N_2296,N_2214);
nor U2511 (N_2511,N_2390,N_2223);
xor U2512 (N_2512,N_2257,N_2290);
xnor U2513 (N_2513,N_2287,N_2344);
or U2514 (N_2514,N_2398,N_2323);
xnor U2515 (N_2515,N_2226,N_2343);
or U2516 (N_2516,N_2213,N_2289);
or U2517 (N_2517,N_2384,N_2296);
nor U2518 (N_2518,N_2214,N_2325);
xor U2519 (N_2519,N_2201,N_2321);
or U2520 (N_2520,N_2215,N_2288);
nor U2521 (N_2521,N_2358,N_2328);
nand U2522 (N_2522,N_2349,N_2382);
xnor U2523 (N_2523,N_2326,N_2324);
nand U2524 (N_2524,N_2343,N_2294);
or U2525 (N_2525,N_2366,N_2386);
nand U2526 (N_2526,N_2391,N_2370);
xor U2527 (N_2527,N_2371,N_2273);
and U2528 (N_2528,N_2305,N_2336);
nand U2529 (N_2529,N_2241,N_2399);
nor U2530 (N_2530,N_2287,N_2355);
and U2531 (N_2531,N_2339,N_2313);
and U2532 (N_2532,N_2211,N_2293);
nor U2533 (N_2533,N_2235,N_2285);
nand U2534 (N_2534,N_2310,N_2267);
xor U2535 (N_2535,N_2276,N_2383);
xnor U2536 (N_2536,N_2288,N_2370);
xor U2537 (N_2537,N_2314,N_2234);
nand U2538 (N_2538,N_2333,N_2346);
nand U2539 (N_2539,N_2289,N_2255);
or U2540 (N_2540,N_2249,N_2396);
xor U2541 (N_2541,N_2359,N_2223);
xnor U2542 (N_2542,N_2290,N_2225);
nand U2543 (N_2543,N_2258,N_2264);
nor U2544 (N_2544,N_2313,N_2335);
nor U2545 (N_2545,N_2234,N_2359);
xor U2546 (N_2546,N_2233,N_2316);
nor U2547 (N_2547,N_2203,N_2393);
or U2548 (N_2548,N_2370,N_2329);
nand U2549 (N_2549,N_2299,N_2300);
and U2550 (N_2550,N_2343,N_2366);
xnor U2551 (N_2551,N_2367,N_2239);
xor U2552 (N_2552,N_2214,N_2248);
nor U2553 (N_2553,N_2381,N_2228);
nor U2554 (N_2554,N_2259,N_2341);
or U2555 (N_2555,N_2272,N_2237);
nand U2556 (N_2556,N_2347,N_2366);
nand U2557 (N_2557,N_2307,N_2227);
or U2558 (N_2558,N_2329,N_2217);
nand U2559 (N_2559,N_2221,N_2353);
xor U2560 (N_2560,N_2203,N_2242);
nand U2561 (N_2561,N_2272,N_2264);
nor U2562 (N_2562,N_2276,N_2357);
and U2563 (N_2563,N_2231,N_2312);
and U2564 (N_2564,N_2373,N_2334);
nand U2565 (N_2565,N_2214,N_2259);
and U2566 (N_2566,N_2341,N_2244);
nor U2567 (N_2567,N_2386,N_2240);
xor U2568 (N_2568,N_2371,N_2337);
nand U2569 (N_2569,N_2260,N_2289);
and U2570 (N_2570,N_2222,N_2379);
nor U2571 (N_2571,N_2364,N_2365);
nand U2572 (N_2572,N_2255,N_2383);
nor U2573 (N_2573,N_2293,N_2387);
and U2574 (N_2574,N_2293,N_2252);
or U2575 (N_2575,N_2201,N_2267);
or U2576 (N_2576,N_2201,N_2221);
and U2577 (N_2577,N_2249,N_2394);
nor U2578 (N_2578,N_2385,N_2379);
nor U2579 (N_2579,N_2310,N_2278);
nand U2580 (N_2580,N_2363,N_2217);
nand U2581 (N_2581,N_2205,N_2353);
nand U2582 (N_2582,N_2300,N_2226);
nor U2583 (N_2583,N_2278,N_2338);
xor U2584 (N_2584,N_2227,N_2292);
nor U2585 (N_2585,N_2243,N_2214);
nor U2586 (N_2586,N_2290,N_2359);
nor U2587 (N_2587,N_2382,N_2245);
nand U2588 (N_2588,N_2283,N_2332);
xor U2589 (N_2589,N_2394,N_2339);
and U2590 (N_2590,N_2216,N_2301);
or U2591 (N_2591,N_2349,N_2222);
nand U2592 (N_2592,N_2322,N_2384);
nand U2593 (N_2593,N_2386,N_2258);
nand U2594 (N_2594,N_2379,N_2241);
and U2595 (N_2595,N_2238,N_2340);
nor U2596 (N_2596,N_2327,N_2315);
and U2597 (N_2597,N_2275,N_2225);
nand U2598 (N_2598,N_2355,N_2267);
xnor U2599 (N_2599,N_2269,N_2278);
and U2600 (N_2600,N_2407,N_2422);
nand U2601 (N_2601,N_2485,N_2507);
nand U2602 (N_2602,N_2598,N_2503);
nand U2603 (N_2603,N_2561,N_2466);
xor U2604 (N_2604,N_2567,N_2424);
and U2605 (N_2605,N_2481,N_2555);
xor U2606 (N_2606,N_2583,N_2425);
xnor U2607 (N_2607,N_2509,N_2429);
nand U2608 (N_2608,N_2406,N_2562);
xor U2609 (N_2609,N_2565,N_2504);
nor U2610 (N_2610,N_2537,N_2441);
and U2611 (N_2611,N_2542,N_2401);
xnor U2612 (N_2612,N_2548,N_2426);
or U2613 (N_2613,N_2516,N_2595);
and U2614 (N_2614,N_2433,N_2460);
nand U2615 (N_2615,N_2432,N_2417);
and U2616 (N_2616,N_2591,N_2515);
xor U2617 (N_2617,N_2563,N_2408);
and U2618 (N_2618,N_2511,N_2445);
nand U2619 (N_2619,N_2400,N_2442);
and U2620 (N_2620,N_2524,N_2462);
nor U2621 (N_2621,N_2594,N_2495);
xor U2622 (N_2622,N_2443,N_2519);
and U2623 (N_2623,N_2456,N_2541);
xor U2624 (N_2624,N_2496,N_2517);
nor U2625 (N_2625,N_2420,N_2581);
nor U2626 (N_2626,N_2547,N_2418);
nand U2627 (N_2627,N_2449,N_2568);
nand U2628 (N_2628,N_2437,N_2454);
nand U2629 (N_2629,N_2569,N_2546);
nor U2630 (N_2630,N_2543,N_2451);
xor U2631 (N_2631,N_2578,N_2582);
and U2632 (N_2632,N_2520,N_2414);
nor U2633 (N_2633,N_2573,N_2464);
and U2634 (N_2634,N_2529,N_2486);
and U2635 (N_2635,N_2483,N_2447);
and U2636 (N_2636,N_2539,N_2491);
nor U2637 (N_2637,N_2579,N_2538);
nor U2638 (N_2638,N_2597,N_2455);
and U2639 (N_2639,N_2550,N_2532);
nor U2640 (N_2640,N_2463,N_2501);
nand U2641 (N_2641,N_2593,N_2472);
and U2642 (N_2642,N_2448,N_2430);
nand U2643 (N_2643,N_2514,N_2477);
nor U2644 (N_2644,N_2435,N_2457);
and U2645 (N_2645,N_2572,N_2416);
nor U2646 (N_2646,N_2575,N_2431);
nand U2647 (N_2647,N_2576,N_2508);
or U2648 (N_2648,N_2510,N_2560);
nor U2649 (N_2649,N_2411,N_2484);
and U2650 (N_2650,N_2586,N_2444);
nor U2651 (N_2651,N_2473,N_2469);
or U2652 (N_2652,N_2436,N_2570);
nand U2653 (N_2653,N_2459,N_2453);
or U2654 (N_2654,N_2482,N_2584);
or U2655 (N_2655,N_2489,N_2592);
or U2656 (N_2656,N_2536,N_2412);
and U2657 (N_2657,N_2587,N_2413);
or U2658 (N_2658,N_2558,N_2530);
and U2659 (N_2659,N_2471,N_2450);
and U2660 (N_2660,N_2438,N_2505);
and U2661 (N_2661,N_2404,N_2410);
nand U2662 (N_2662,N_2440,N_2580);
and U2663 (N_2663,N_2552,N_2480);
or U2664 (N_2664,N_2478,N_2461);
nor U2665 (N_2665,N_2476,N_2494);
or U2666 (N_2666,N_2402,N_2564);
or U2667 (N_2667,N_2409,N_2512);
nand U2668 (N_2668,N_2492,N_2589);
nand U2669 (N_2669,N_2533,N_2499);
xor U2670 (N_2670,N_2493,N_2566);
nor U2671 (N_2671,N_2518,N_2528);
or U2672 (N_2672,N_2475,N_2585);
and U2673 (N_2673,N_2534,N_2554);
and U2674 (N_2674,N_2465,N_2551);
nand U2675 (N_2675,N_2452,N_2428);
xnor U2676 (N_2676,N_2458,N_2487);
nor U2677 (N_2677,N_2521,N_2506);
or U2678 (N_2678,N_2527,N_2470);
and U2679 (N_2679,N_2500,N_2526);
nor U2680 (N_2680,N_2502,N_2557);
and U2681 (N_2681,N_2599,N_2556);
nor U2682 (N_2682,N_2479,N_2535);
and U2683 (N_2683,N_2549,N_2525);
or U2684 (N_2684,N_2596,N_2446);
nand U2685 (N_2685,N_2590,N_2403);
nand U2686 (N_2686,N_2571,N_2497);
xnor U2687 (N_2687,N_2467,N_2513);
or U2688 (N_2688,N_2421,N_2523);
xor U2689 (N_2689,N_2544,N_2540);
nor U2690 (N_2690,N_2415,N_2588);
xor U2691 (N_2691,N_2545,N_2434);
nand U2692 (N_2692,N_2577,N_2468);
xor U2693 (N_2693,N_2553,N_2574);
and U2694 (N_2694,N_2490,N_2419);
and U2695 (N_2695,N_2405,N_2498);
nor U2696 (N_2696,N_2559,N_2423);
nand U2697 (N_2697,N_2531,N_2474);
or U2698 (N_2698,N_2439,N_2522);
and U2699 (N_2699,N_2427,N_2488);
or U2700 (N_2700,N_2482,N_2498);
xnor U2701 (N_2701,N_2434,N_2455);
xnor U2702 (N_2702,N_2406,N_2459);
and U2703 (N_2703,N_2491,N_2499);
xor U2704 (N_2704,N_2553,N_2546);
nand U2705 (N_2705,N_2527,N_2539);
or U2706 (N_2706,N_2451,N_2419);
and U2707 (N_2707,N_2423,N_2536);
xor U2708 (N_2708,N_2594,N_2476);
or U2709 (N_2709,N_2572,N_2576);
or U2710 (N_2710,N_2497,N_2405);
and U2711 (N_2711,N_2473,N_2578);
nand U2712 (N_2712,N_2573,N_2459);
and U2713 (N_2713,N_2406,N_2453);
nand U2714 (N_2714,N_2500,N_2426);
nand U2715 (N_2715,N_2525,N_2595);
and U2716 (N_2716,N_2466,N_2462);
and U2717 (N_2717,N_2549,N_2497);
xor U2718 (N_2718,N_2465,N_2587);
nand U2719 (N_2719,N_2578,N_2532);
xnor U2720 (N_2720,N_2529,N_2440);
or U2721 (N_2721,N_2550,N_2425);
nor U2722 (N_2722,N_2410,N_2457);
and U2723 (N_2723,N_2505,N_2433);
or U2724 (N_2724,N_2590,N_2559);
xor U2725 (N_2725,N_2541,N_2460);
xor U2726 (N_2726,N_2443,N_2440);
or U2727 (N_2727,N_2558,N_2529);
nand U2728 (N_2728,N_2477,N_2435);
nand U2729 (N_2729,N_2537,N_2573);
xnor U2730 (N_2730,N_2438,N_2466);
xor U2731 (N_2731,N_2508,N_2564);
or U2732 (N_2732,N_2469,N_2532);
or U2733 (N_2733,N_2438,N_2551);
nor U2734 (N_2734,N_2487,N_2533);
and U2735 (N_2735,N_2478,N_2521);
nand U2736 (N_2736,N_2483,N_2540);
nand U2737 (N_2737,N_2463,N_2432);
or U2738 (N_2738,N_2482,N_2587);
and U2739 (N_2739,N_2431,N_2567);
xnor U2740 (N_2740,N_2562,N_2462);
and U2741 (N_2741,N_2407,N_2484);
nor U2742 (N_2742,N_2547,N_2477);
nor U2743 (N_2743,N_2439,N_2582);
xor U2744 (N_2744,N_2509,N_2535);
and U2745 (N_2745,N_2494,N_2426);
xor U2746 (N_2746,N_2508,N_2596);
nor U2747 (N_2747,N_2451,N_2412);
nand U2748 (N_2748,N_2439,N_2409);
nor U2749 (N_2749,N_2545,N_2414);
nor U2750 (N_2750,N_2425,N_2580);
and U2751 (N_2751,N_2424,N_2572);
and U2752 (N_2752,N_2493,N_2544);
nand U2753 (N_2753,N_2458,N_2457);
or U2754 (N_2754,N_2475,N_2462);
and U2755 (N_2755,N_2462,N_2439);
nand U2756 (N_2756,N_2407,N_2462);
nand U2757 (N_2757,N_2435,N_2432);
nor U2758 (N_2758,N_2516,N_2500);
or U2759 (N_2759,N_2556,N_2521);
or U2760 (N_2760,N_2597,N_2400);
and U2761 (N_2761,N_2585,N_2413);
nor U2762 (N_2762,N_2499,N_2585);
xor U2763 (N_2763,N_2558,N_2512);
nand U2764 (N_2764,N_2442,N_2420);
xnor U2765 (N_2765,N_2525,N_2479);
nor U2766 (N_2766,N_2460,N_2516);
or U2767 (N_2767,N_2417,N_2436);
nand U2768 (N_2768,N_2454,N_2413);
nand U2769 (N_2769,N_2569,N_2459);
or U2770 (N_2770,N_2432,N_2414);
and U2771 (N_2771,N_2514,N_2510);
and U2772 (N_2772,N_2472,N_2550);
or U2773 (N_2773,N_2524,N_2435);
nor U2774 (N_2774,N_2567,N_2530);
xor U2775 (N_2775,N_2545,N_2526);
xor U2776 (N_2776,N_2517,N_2485);
or U2777 (N_2777,N_2505,N_2401);
and U2778 (N_2778,N_2512,N_2450);
nor U2779 (N_2779,N_2597,N_2535);
xnor U2780 (N_2780,N_2402,N_2540);
and U2781 (N_2781,N_2522,N_2510);
nor U2782 (N_2782,N_2519,N_2468);
or U2783 (N_2783,N_2495,N_2499);
or U2784 (N_2784,N_2442,N_2426);
nand U2785 (N_2785,N_2460,N_2542);
nor U2786 (N_2786,N_2531,N_2472);
nand U2787 (N_2787,N_2409,N_2598);
nand U2788 (N_2788,N_2558,N_2436);
nand U2789 (N_2789,N_2597,N_2487);
and U2790 (N_2790,N_2407,N_2589);
xor U2791 (N_2791,N_2508,N_2409);
nor U2792 (N_2792,N_2531,N_2556);
xor U2793 (N_2793,N_2571,N_2414);
xnor U2794 (N_2794,N_2487,N_2428);
and U2795 (N_2795,N_2458,N_2409);
nand U2796 (N_2796,N_2455,N_2541);
xor U2797 (N_2797,N_2430,N_2542);
nand U2798 (N_2798,N_2592,N_2555);
nor U2799 (N_2799,N_2443,N_2487);
and U2800 (N_2800,N_2692,N_2788);
nor U2801 (N_2801,N_2612,N_2627);
and U2802 (N_2802,N_2610,N_2750);
nor U2803 (N_2803,N_2678,N_2677);
or U2804 (N_2804,N_2721,N_2719);
and U2805 (N_2805,N_2734,N_2651);
nand U2806 (N_2806,N_2726,N_2782);
or U2807 (N_2807,N_2689,N_2600);
and U2808 (N_2808,N_2667,N_2776);
and U2809 (N_2809,N_2609,N_2784);
nor U2810 (N_2810,N_2626,N_2696);
or U2811 (N_2811,N_2711,N_2728);
nand U2812 (N_2812,N_2781,N_2765);
nand U2813 (N_2813,N_2698,N_2643);
xor U2814 (N_2814,N_2729,N_2613);
nand U2815 (N_2815,N_2683,N_2771);
nor U2816 (N_2816,N_2702,N_2707);
nor U2817 (N_2817,N_2709,N_2631);
and U2818 (N_2818,N_2701,N_2608);
nand U2819 (N_2819,N_2620,N_2688);
xnor U2820 (N_2820,N_2694,N_2716);
nand U2821 (N_2821,N_2653,N_2796);
xor U2822 (N_2822,N_2706,N_2650);
or U2823 (N_2823,N_2630,N_2679);
and U2824 (N_2824,N_2697,N_2637);
xnor U2825 (N_2825,N_2718,N_2681);
xor U2826 (N_2826,N_2756,N_2703);
nand U2827 (N_2827,N_2684,N_2722);
xor U2828 (N_2828,N_2708,N_2790);
xor U2829 (N_2829,N_2743,N_2783);
or U2830 (N_2830,N_2622,N_2735);
and U2831 (N_2831,N_2648,N_2733);
xnor U2832 (N_2832,N_2699,N_2789);
or U2833 (N_2833,N_2662,N_2685);
nor U2834 (N_2834,N_2601,N_2793);
xor U2835 (N_2835,N_2607,N_2760);
nor U2836 (N_2836,N_2705,N_2621);
xnor U2837 (N_2837,N_2792,N_2611);
or U2838 (N_2838,N_2780,N_2691);
and U2839 (N_2839,N_2604,N_2661);
or U2840 (N_2840,N_2658,N_2766);
nor U2841 (N_2841,N_2740,N_2649);
xnor U2842 (N_2842,N_2695,N_2647);
or U2843 (N_2843,N_2787,N_2723);
xnor U2844 (N_2844,N_2720,N_2639);
and U2845 (N_2845,N_2616,N_2757);
nand U2846 (N_2846,N_2632,N_2670);
or U2847 (N_2847,N_2657,N_2742);
nand U2848 (N_2848,N_2629,N_2725);
nor U2849 (N_2849,N_2798,N_2738);
nand U2850 (N_2850,N_2666,N_2762);
xor U2851 (N_2851,N_2663,N_2713);
and U2852 (N_2852,N_2755,N_2741);
nor U2853 (N_2853,N_2636,N_2777);
nand U2854 (N_2854,N_2791,N_2751);
xor U2855 (N_2855,N_2676,N_2736);
or U2856 (N_2856,N_2619,N_2673);
or U2857 (N_2857,N_2665,N_2749);
or U2858 (N_2858,N_2778,N_2775);
nand U2859 (N_2859,N_2764,N_2772);
xor U2860 (N_2860,N_2794,N_2737);
nor U2861 (N_2861,N_2739,N_2618);
or U2862 (N_2862,N_2686,N_2745);
and U2863 (N_2863,N_2635,N_2652);
and U2864 (N_2864,N_2638,N_2797);
nand U2865 (N_2865,N_2640,N_2642);
nor U2866 (N_2866,N_2704,N_2672);
nor U2867 (N_2867,N_2763,N_2606);
or U2868 (N_2868,N_2680,N_2625);
and U2869 (N_2869,N_2628,N_2759);
or U2870 (N_2870,N_2715,N_2786);
or U2871 (N_2871,N_2654,N_2732);
nand U2872 (N_2872,N_2761,N_2799);
and U2873 (N_2873,N_2671,N_2615);
or U2874 (N_2874,N_2779,N_2717);
and U2875 (N_2875,N_2747,N_2633);
or U2876 (N_2876,N_2795,N_2675);
xor U2877 (N_2877,N_2693,N_2617);
nand U2878 (N_2878,N_2605,N_2769);
nand U2879 (N_2879,N_2646,N_2641);
or U2880 (N_2880,N_2731,N_2614);
nand U2881 (N_2881,N_2767,N_2724);
or U2882 (N_2882,N_2655,N_2754);
and U2883 (N_2883,N_2753,N_2687);
nand U2884 (N_2884,N_2748,N_2682);
or U2885 (N_2885,N_2768,N_2669);
xor U2886 (N_2886,N_2623,N_2602);
nand U2887 (N_2887,N_2712,N_2785);
and U2888 (N_2888,N_2714,N_2656);
and U2889 (N_2889,N_2690,N_2603);
nand U2890 (N_2890,N_2758,N_2730);
or U2891 (N_2891,N_2727,N_2744);
and U2892 (N_2892,N_2659,N_2645);
nand U2893 (N_2893,N_2770,N_2746);
xor U2894 (N_2894,N_2773,N_2752);
and U2895 (N_2895,N_2664,N_2624);
and U2896 (N_2896,N_2660,N_2700);
and U2897 (N_2897,N_2674,N_2644);
nand U2898 (N_2898,N_2710,N_2774);
nor U2899 (N_2899,N_2668,N_2634);
and U2900 (N_2900,N_2794,N_2706);
xor U2901 (N_2901,N_2719,N_2693);
nor U2902 (N_2902,N_2632,N_2745);
or U2903 (N_2903,N_2640,N_2745);
or U2904 (N_2904,N_2730,N_2658);
nor U2905 (N_2905,N_2602,N_2646);
or U2906 (N_2906,N_2628,N_2710);
and U2907 (N_2907,N_2794,N_2789);
nand U2908 (N_2908,N_2795,N_2740);
xor U2909 (N_2909,N_2767,N_2733);
and U2910 (N_2910,N_2696,N_2611);
or U2911 (N_2911,N_2631,N_2638);
or U2912 (N_2912,N_2684,N_2699);
xor U2913 (N_2913,N_2699,N_2666);
or U2914 (N_2914,N_2652,N_2728);
or U2915 (N_2915,N_2744,N_2791);
xor U2916 (N_2916,N_2739,N_2659);
nor U2917 (N_2917,N_2673,N_2734);
or U2918 (N_2918,N_2671,N_2703);
nor U2919 (N_2919,N_2672,N_2767);
or U2920 (N_2920,N_2630,N_2797);
nor U2921 (N_2921,N_2675,N_2747);
xor U2922 (N_2922,N_2718,N_2607);
or U2923 (N_2923,N_2641,N_2713);
nor U2924 (N_2924,N_2706,N_2767);
and U2925 (N_2925,N_2634,N_2670);
and U2926 (N_2926,N_2750,N_2797);
nand U2927 (N_2927,N_2730,N_2789);
or U2928 (N_2928,N_2789,N_2710);
and U2929 (N_2929,N_2684,N_2798);
nand U2930 (N_2930,N_2719,N_2713);
nand U2931 (N_2931,N_2772,N_2699);
nand U2932 (N_2932,N_2744,N_2694);
or U2933 (N_2933,N_2614,N_2777);
nor U2934 (N_2934,N_2761,N_2711);
or U2935 (N_2935,N_2683,N_2648);
and U2936 (N_2936,N_2778,N_2798);
and U2937 (N_2937,N_2680,N_2728);
or U2938 (N_2938,N_2783,N_2647);
nor U2939 (N_2939,N_2783,N_2620);
nor U2940 (N_2940,N_2732,N_2624);
or U2941 (N_2941,N_2641,N_2712);
nand U2942 (N_2942,N_2793,N_2711);
nor U2943 (N_2943,N_2684,N_2690);
nand U2944 (N_2944,N_2652,N_2769);
nand U2945 (N_2945,N_2723,N_2671);
nand U2946 (N_2946,N_2702,N_2689);
and U2947 (N_2947,N_2789,N_2716);
or U2948 (N_2948,N_2686,N_2633);
nand U2949 (N_2949,N_2623,N_2707);
or U2950 (N_2950,N_2627,N_2739);
nor U2951 (N_2951,N_2656,N_2640);
nand U2952 (N_2952,N_2747,N_2716);
xor U2953 (N_2953,N_2747,N_2695);
and U2954 (N_2954,N_2677,N_2704);
or U2955 (N_2955,N_2644,N_2776);
or U2956 (N_2956,N_2654,N_2690);
nor U2957 (N_2957,N_2709,N_2661);
nand U2958 (N_2958,N_2727,N_2650);
nor U2959 (N_2959,N_2735,N_2671);
nand U2960 (N_2960,N_2786,N_2687);
nand U2961 (N_2961,N_2632,N_2744);
xnor U2962 (N_2962,N_2721,N_2783);
nor U2963 (N_2963,N_2682,N_2609);
or U2964 (N_2964,N_2759,N_2611);
or U2965 (N_2965,N_2674,N_2735);
or U2966 (N_2966,N_2765,N_2692);
and U2967 (N_2967,N_2607,N_2743);
nand U2968 (N_2968,N_2637,N_2767);
and U2969 (N_2969,N_2777,N_2618);
xor U2970 (N_2970,N_2723,N_2775);
nor U2971 (N_2971,N_2708,N_2661);
or U2972 (N_2972,N_2790,N_2687);
nor U2973 (N_2973,N_2688,N_2658);
nand U2974 (N_2974,N_2631,N_2629);
nor U2975 (N_2975,N_2741,N_2751);
xor U2976 (N_2976,N_2754,N_2696);
or U2977 (N_2977,N_2738,N_2624);
nor U2978 (N_2978,N_2698,N_2736);
nand U2979 (N_2979,N_2716,N_2604);
and U2980 (N_2980,N_2762,N_2711);
nor U2981 (N_2981,N_2635,N_2677);
nor U2982 (N_2982,N_2601,N_2708);
xor U2983 (N_2983,N_2687,N_2702);
nor U2984 (N_2984,N_2658,N_2732);
and U2985 (N_2985,N_2661,N_2662);
or U2986 (N_2986,N_2687,N_2759);
nor U2987 (N_2987,N_2728,N_2705);
xnor U2988 (N_2988,N_2746,N_2719);
nor U2989 (N_2989,N_2772,N_2703);
nand U2990 (N_2990,N_2673,N_2793);
nor U2991 (N_2991,N_2643,N_2760);
xor U2992 (N_2992,N_2608,N_2660);
and U2993 (N_2993,N_2610,N_2796);
and U2994 (N_2994,N_2733,N_2750);
nor U2995 (N_2995,N_2611,N_2714);
nand U2996 (N_2996,N_2698,N_2700);
or U2997 (N_2997,N_2684,N_2696);
or U2998 (N_2998,N_2607,N_2675);
or U2999 (N_2999,N_2738,N_2665);
xnor U3000 (N_3000,N_2854,N_2988);
nor U3001 (N_3001,N_2915,N_2919);
or U3002 (N_3002,N_2935,N_2874);
xor U3003 (N_3003,N_2906,N_2867);
or U3004 (N_3004,N_2828,N_2989);
and U3005 (N_3005,N_2934,N_2878);
or U3006 (N_3006,N_2925,N_2894);
nor U3007 (N_3007,N_2995,N_2922);
and U3008 (N_3008,N_2967,N_2813);
and U3009 (N_3009,N_2964,N_2857);
nand U3010 (N_3010,N_2852,N_2974);
or U3011 (N_3011,N_2950,N_2877);
nand U3012 (N_3012,N_2817,N_2820);
and U3013 (N_3013,N_2971,N_2947);
nand U3014 (N_3014,N_2962,N_2842);
xnor U3015 (N_3015,N_2969,N_2824);
nor U3016 (N_3016,N_2843,N_2881);
or U3017 (N_3017,N_2865,N_2864);
or U3018 (N_3018,N_2996,N_2999);
or U3019 (N_3019,N_2931,N_2970);
or U3020 (N_3020,N_2923,N_2811);
nor U3021 (N_3021,N_2900,N_2991);
nand U3022 (N_3022,N_2801,N_2916);
xor U3023 (N_3023,N_2993,N_2903);
xor U3024 (N_3024,N_2850,N_2924);
and U3025 (N_3025,N_2836,N_2818);
nand U3026 (N_3026,N_2875,N_2913);
nand U3027 (N_3027,N_2902,N_2805);
or U3028 (N_3028,N_2888,N_2972);
nor U3029 (N_3029,N_2910,N_2914);
xnor U3030 (N_3030,N_2809,N_2961);
and U3031 (N_3031,N_2933,N_2815);
and U3032 (N_3032,N_2833,N_2921);
nand U3033 (N_3033,N_2909,N_2901);
nor U3034 (N_3034,N_2814,N_2855);
and U3035 (N_3035,N_2978,N_2958);
nand U3036 (N_3036,N_2897,N_2955);
nor U3037 (N_3037,N_2835,N_2807);
nor U3038 (N_3038,N_2886,N_2890);
nor U3039 (N_3039,N_2987,N_2968);
and U3040 (N_3040,N_2904,N_2942);
xor U3041 (N_3041,N_2889,N_2837);
nor U3042 (N_3042,N_2912,N_2860);
nor U3043 (N_3043,N_2975,N_2823);
and U3044 (N_3044,N_2868,N_2896);
nor U3045 (N_3045,N_2946,N_2821);
nor U3046 (N_3046,N_2982,N_2840);
xor U3047 (N_3047,N_2976,N_2810);
nor U3048 (N_3048,N_2841,N_2851);
nand U3049 (N_3049,N_2905,N_2939);
xor U3050 (N_3050,N_2907,N_2891);
and U3051 (N_3051,N_2838,N_2803);
or U3052 (N_3052,N_2938,N_2831);
or U3053 (N_3053,N_2927,N_2883);
xor U3054 (N_3054,N_2825,N_2829);
nand U3055 (N_3055,N_2863,N_2990);
nand U3056 (N_3056,N_2918,N_2844);
and U3057 (N_3057,N_2822,N_2959);
nand U3058 (N_3058,N_2917,N_2997);
and U3059 (N_3059,N_2806,N_2856);
nor U3060 (N_3060,N_2928,N_2885);
and U3061 (N_3061,N_2992,N_2966);
or U3062 (N_3062,N_2985,N_2940);
or U3063 (N_3063,N_2952,N_2937);
nor U3064 (N_3064,N_2884,N_2819);
and U3065 (N_3065,N_2949,N_2859);
and U3066 (N_3066,N_2953,N_2930);
nand U3067 (N_3067,N_2957,N_2893);
nor U3068 (N_3068,N_2979,N_2960);
nor U3069 (N_3069,N_2986,N_2846);
nor U3070 (N_3070,N_2853,N_2839);
or U3071 (N_3071,N_2977,N_2869);
and U3072 (N_3072,N_2872,N_2858);
nand U3073 (N_3073,N_2849,N_2984);
nand U3074 (N_3074,N_2936,N_2871);
xnor U3075 (N_3075,N_2954,N_2920);
nor U3076 (N_3076,N_2826,N_2948);
nand U3077 (N_3077,N_2808,N_2847);
nand U3078 (N_3078,N_2861,N_2876);
xor U3079 (N_3079,N_2804,N_2862);
xor U3080 (N_3080,N_2932,N_2834);
or U3081 (N_3081,N_2963,N_2983);
nor U3082 (N_3082,N_2816,N_2908);
and U3083 (N_3083,N_2965,N_2945);
nor U3084 (N_3084,N_2981,N_2926);
nand U3085 (N_3085,N_2895,N_2911);
nand U3086 (N_3086,N_2832,N_2973);
or U3087 (N_3087,N_2998,N_2941);
nor U3088 (N_3088,N_2994,N_2879);
xor U3089 (N_3089,N_2873,N_2800);
nor U3090 (N_3090,N_2892,N_2812);
nand U3091 (N_3091,N_2802,N_2827);
or U3092 (N_3092,N_2956,N_2845);
or U3093 (N_3093,N_2898,N_2944);
and U3094 (N_3094,N_2929,N_2848);
and U3095 (N_3095,N_2951,N_2870);
nor U3096 (N_3096,N_2880,N_2866);
and U3097 (N_3097,N_2887,N_2943);
or U3098 (N_3098,N_2899,N_2830);
nand U3099 (N_3099,N_2882,N_2980);
xnor U3100 (N_3100,N_2944,N_2922);
xor U3101 (N_3101,N_2870,N_2816);
nand U3102 (N_3102,N_2898,N_2838);
nand U3103 (N_3103,N_2847,N_2993);
nor U3104 (N_3104,N_2963,N_2933);
xor U3105 (N_3105,N_2902,N_2951);
nor U3106 (N_3106,N_2834,N_2934);
xnor U3107 (N_3107,N_2936,N_2985);
nor U3108 (N_3108,N_2864,N_2971);
nand U3109 (N_3109,N_2862,N_2919);
or U3110 (N_3110,N_2908,N_2889);
nor U3111 (N_3111,N_2820,N_2855);
and U3112 (N_3112,N_2923,N_2842);
and U3113 (N_3113,N_2907,N_2954);
or U3114 (N_3114,N_2900,N_2845);
nand U3115 (N_3115,N_2860,N_2867);
and U3116 (N_3116,N_2857,N_2954);
and U3117 (N_3117,N_2867,N_2889);
nor U3118 (N_3118,N_2827,N_2839);
and U3119 (N_3119,N_2922,N_2982);
or U3120 (N_3120,N_2887,N_2998);
or U3121 (N_3121,N_2809,N_2902);
and U3122 (N_3122,N_2870,N_2844);
nand U3123 (N_3123,N_2818,N_2986);
nand U3124 (N_3124,N_2950,N_2983);
nor U3125 (N_3125,N_2921,N_2925);
or U3126 (N_3126,N_2909,N_2802);
and U3127 (N_3127,N_2808,N_2917);
and U3128 (N_3128,N_2939,N_2848);
and U3129 (N_3129,N_2985,N_2804);
nor U3130 (N_3130,N_2843,N_2964);
nor U3131 (N_3131,N_2961,N_2866);
xor U3132 (N_3132,N_2878,N_2856);
xnor U3133 (N_3133,N_2836,N_2807);
or U3134 (N_3134,N_2950,N_2888);
nor U3135 (N_3135,N_2941,N_2884);
and U3136 (N_3136,N_2866,N_2983);
nor U3137 (N_3137,N_2813,N_2843);
and U3138 (N_3138,N_2909,N_2938);
and U3139 (N_3139,N_2993,N_2972);
nand U3140 (N_3140,N_2962,N_2826);
and U3141 (N_3141,N_2807,N_2927);
or U3142 (N_3142,N_2861,N_2888);
and U3143 (N_3143,N_2983,N_2973);
and U3144 (N_3144,N_2815,N_2894);
or U3145 (N_3145,N_2852,N_2836);
nor U3146 (N_3146,N_2918,N_2982);
nand U3147 (N_3147,N_2920,N_2948);
and U3148 (N_3148,N_2809,N_2882);
or U3149 (N_3149,N_2921,N_2862);
or U3150 (N_3150,N_2836,N_2837);
nor U3151 (N_3151,N_2880,N_2805);
and U3152 (N_3152,N_2937,N_2851);
xnor U3153 (N_3153,N_2998,N_2942);
nand U3154 (N_3154,N_2927,N_2930);
xnor U3155 (N_3155,N_2862,N_2873);
or U3156 (N_3156,N_2882,N_2964);
nand U3157 (N_3157,N_2887,N_2991);
and U3158 (N_3158,N_2905,N_2858);
and U3159 (N_3159,N_2973,N_2831);
or U3160 (N_3160,N_2968,N_2820);
nand U3161 (N_3161,N_2909,N_2994);
or U3162 (N_3162,N_2922,N_2861);
xor U3163 (N_3163,N_2922,N_2914);
and U3164 (N_3164,N_2839,N_2881);
or U3165 (N_3165,N_2856,N_2986);
xnor U3166 (N_3166,N_2878,N_2846);
or U3167 (N_3167,N_2882,N_2940);
nor U3168 (N_3168,N_2981,N_2950);
and U3169 (N_3169,N_2871,N_2884);
or U3170 (N_3170,N_2920,N_2878);
nor U3171 (N_3171,N_2801,N_2870);
nand U3172 (N_3172,N_2818,N_2882);
nand U3173 (N_3173,N_2955,N_2814);
xnor U3174 (N_3174,N_2930,N_2996);
xnor U3175 (N_3175,N_2842,N_2883);
nor U3176 (N_3176,N_2953,N_2943);
or U3177 (N_3177,N_2891,N_2990);
nand U3178 (N_3178,N_2912,N_2931);
xor U3179 (N_3179,N_2946,N_2902);
nand U3180 (N_3180,N_2816,N_2853);
or U3181 (N_3181,N_2835,N_2899);
xor U3182 (N_3182,N_2887,N_2803);
and U3183 (N_3183,N_2966,N_2872);
nor U3184 (N_3184,N_2941,N_2982);
xnor U3185 (N_3185,N_2973,N_2859);
xnor U3186 (N_3186,N_2974,N_2838);
nor U3187 (N_3187,N_2942,N_2916);
xor U3188 (N_3188,N_2824,N_2838);
and U3189 (N_3189,N_2872,N_2835);
or U3190 (N_3190,N_2823,N_2904);
or U3191 (N_3191,N_2835,N_2841);
or U3192 (N_3192,N_2923,N_2904);
xor U3193 (N_3193,N_2911,N_2929);
xor U3194 (N_3194,N_2917,N_2938);
xnor U3195 (N_3195,N_2961,N_2826);
and U3196 (N_3196,N_2864,N_2956);
nand U3197 (N_3197,N_2900,N_2911);
or U3198 (N_3198,N_2901,N_2890);
and U3199 (N_3199,N_2963,N_2958);
nor U3200 (N_3200,N_3166,N_3132);
nand U3201 (N_3201,N_3056,N_3047);
nor U3202 (N_3202,N_3057,N_3177);
or U3203 (N_3203,N_3176,N_3099);
xnor U3204 (N_3204,N_3042,N_3008);
and U3205 (N_3205,N_3077,N_3088);
nand U3206 (N_3206,N_3139,N_3023);
nor U3207 (N_3207,N_3049,N_3183);
xor U3208 (N_3208,N_3011,N_3193);
nor U3209 (N_3209,N_3004,N_3010);
or U3210 (N_3210,N_3085,N_3178);
or U3211 (N_3211,N_3130,N_3121);
and U3212 (N_3212,N_3180,N_3100);
and U3213 (N_3213,N_3107,N_3189);
nand U3214 (N_3214,N_3138,N_3198);
xor U3215 (N_3215,N_3199,N_3112);
nor U3216 (N_3216,N_3124,N_3046);
or U3217 (N_3217,N_3053,N_3184);
nor U3218 (N_3218,N_3161,N_3172);
nand U3219 (N_3219,N_3186,N_3142);
nor U3220 (N_3220,N_3016,N_3086);
or U3221 (N_3221,N_3167,N_3116);
or U3222 (N_3222,N_3015,N_3170);
nand U3223 (N_3223,N_3129,N_3181);
and U3224 (N_3224,N_3092,N_3187);
xnor U3225 (N_3225,N_3159,N_3014);
or U3226 (N_3226,N_3054,N_3171);
xnor U3227 (N_3227,N_3179,N_3070);
and U3228 (N_3228,N_3148,N_3135);
and U3229 (N_3229,N_3038,N_3102);
nor U3230 (N_3230,N_3191,N_3078);
or U3231 (N_3231,N_3087,N_3064);
or U3232 (N_3232,N_3175,N_3007);
or U3233 (N_3233,N_3145,N_3163);
xnor U3234 (N_3234,N_3105,N_3072);
or U3235 (N_3235,N_3143,N_3034);
xnor U3236 (N_3236,N_3098,N_3106);
and U3237 (N_3237,N_3144,N_3018);
nand U3238 (N_3238,N_3120,N_3156);
nand U3239 (N_3239,N_3160,N_3174);
and U3240 (N_3240,N_3125,N_3022);
nor U3241 (N_3241,N_3122,N_3128);
nor U3242 (N_3242,N_3052,N_3059);
nand U3243 (N_3243,N_3131,N_3157);
and U3244 (N_3244,N_3061,N_3197);
xor U3245 (N_3245,N_3073,N_3089);
nand U3246 (N_3246,N_3152,N_3101);
nor U3247 (N_3247,N_3032,N_3103);
or U3248 (N_3248,N_3019,N_3095);
xnor U3249 (N_3249,N_3025,N_3079);
and U3250 (N_3250,N_3136,N_3063);
nor U3251 (N_3251,N_3123,N_3158);
nor U3252 (N_3252,N_3045,N_3182);
nor U3253 (N_3253,N_3093,N_3060);
and U3254 (N_3254,N_3013,N_3173);
nor U3255 (N_3255,N_3028,N_3006);
xnor U3256 (N_3256,N_3115,N_3062);
or U3257 (N_3257,N_3024,N_3196);
nor U3258 (N_3258,N_3151,N_3058);
or U3259 (N_3259,N_3104,N_3000);
nor U3260 (N_3260,N_3114,N_3068);
xnor U3261 (N_3261,N_3192,N_3033);
and U3262 (N_3262,N_3137,N_3190);
and U3263 (N_3263,N_3067,N_3040);
nor U3264 (N_3264,N_3149,N_3043);
nor U3265 (N_3265,N_3126,N_3076);
nor U3266 (N_3266,N_3127,N_3118);
and U3267 (N_3267,N_3108,N_3066);
nand U3268 (N_3268,N_3017,N_3146);
nand U3269 (N_3269,N_3185,N_3051);
and U3270 (N_3270,N_3050,N_3020);
nor U3271 (N_3271,N_3084,N_3117);
xnor U3272 (N_3272,N_3096,N_3154);
or U3273 (N_3273,N_3164,N_3119);
nor U3274 (N_3274,N_3110,N_3026);
nor U3275 (N_3275,N_3075,N_3001);
or U3276 (N_3276,N_3031,N_3082);
nand U3277 (N_3277,N_3094,N_3035);
xor U3278 (N_3278,N_3133,N_3150);
or U3279 (N_3279,N_3113,N_3162);
or U3280 (N_3280,N_3044,N_3037);
nand U3281 (N_3281,N_3081,N_3188);
nor U3282 (N_3282,N_3169,N_3055);
or U3283 (N_3283,N_3194,N_3090);
xor U3284 (N_3284,N_3069,N_3039);
xnor U3285 (N_3285,N_3155,N_3195);
and U3286 (N_3286,N_3141,N_3134);
xnor U3287 (N_3287,N_3027,N_3030);
nor U3288 (N_3288,N_3140,N_3071);
or U3289 (N_3289,N_3168,N_3029);
nor U3290 (N_3290,N_3111,N_3097);
nand U3291 (N_3291,N_3041,N_3021);
or U3292 (N_3292,N_3005,N_3080);
nand U3293 (N_3293,N_3153,N_3036);
nor U3294 (N_3294,N_3074,N_3009);
and U3295 (N_3295,N_3002,N_3065);
or U3296 (N_3296,N_3048,N_3109);
xnor U3297 (N_3297,N_3147,N_3083);
nand U3298 (N_3298,N_3091,N_3003);
and U3299 (N_3299,N_3165,N_3012);
nand U3300 (N_3300,N_3077,N_3149);
xnor U3301 (N_3301,N_3195,N_3005);
nor U3302 (N_3302,N_3046,N_3099);
xnor U3303 (N_3303,N_3122,N_3067);
xnor U3304 (N_3304,N_3195,N_3154);
and U3305 (N_3305,N_3064,N_3188);
or U3306 (N_3306,N_3095,N_3032);
or U3307 (N_3307,N_3164,N_3014);
nor U3308 (N_3308,N_3105,N_3163);
nand U3309 (N_3309,N_3060,N_3030);
nand U3310 (N_3310,N_3018,N_3048);
nand U3311 (N_3311,N_3057,N_3005);
nand U3312 (N_3312,N_3078,N_3090);
nand U3313 (N_3313,N_3098,N_3184);
and U3314 (N_3314,N_3084,N_3082);
xor U3315 (N_3315,N_3013,N_3106);
nor U3316 (N_3316,N_3025,N_3188);
nand U3317 (N_3317,N_3184,N_3154);
nand U3318 (N_3318,N_3197,N_3187);
or U3319 (N_3319,N_3135,N_3195);
nand U3320 (N_3320,N_3129,N_3145);
xor U3321 (N_3321,N_3144,N_3050);
and U3322 (N_3322,N_3099,N_3094);
nand U3323 (N_3323,N_3093,N_3199);
nor U3324 (N_3324,N_3013,N_3107);
or U3325 (N_3325,N_3080,N_3081);
and U3326 (N_3326,N_3139,N_3059);
nor U3327 (N_3327,N_3095,N_3119);
xnor U3328 (N_3328,N_3167,N_3191);
and U3329 (N_3329,N_3121,N_3191);
xnor U3330 (N_3330,N_3010,N_3071);
or U3331 (N_3331,N_3156,N_3050);
and U3332 (N_3332,N_3155,N_3109);
or U3333 (N_3333,N_3003,N_3183);
nand U3334 (N_3334,N_3008,N_3180);
nor U3335 (N_3335,N_3009,N_3182);
nor U3336 (N_3336,N_3066,N_3181);
and U3337 (N_3337,N_3031,N_3142);
xor U3338 (N_3338,N_3062,N_3008);
nor U3339 (N_3339,N_3199,N_3063);
and U3340 (N_3340,N_3152,N_3049);
xor U3341 (N_3341,N_3051,N_3138);
nand U3342 (N_3342,N_3175,N_3157);
or U3343 (N_3343,N_3045,N_3155);
nor U3344 (N_3344,N_3050,N_3138);
nor U3345 (N_3345,N_3009,N_3100);
nor U3346 (N_3346,N_3150,N_3161);
and U3347 (N_3347,N_3034,N_3182);
and U3348 (N_3348,N_3149,N_3127);
xnor U3349 (N_3349,N_3146,N_3111);
xnor U3350 (N_3350,N_3168,N_3069);
nor U3351 (N_3351,N_3061,N_3049);
nor U3352 (N_3352,N_3162,N_3132);
and U3353 (N_3353,N_3197,N_3167);
or U3354 (N_3354,N_3057,N_3060);
nand U3355 (N_3355,N_3195,N_3181);
and U3356 (N_3356,N_3162,N_3040);
xnor U3357 (N_3357,N_3055,N_3143);
nand U3358 (N_3358,N_3006,N_3142);
xnor U3359 (N_3359,N_3027,N_3168);
nor U3360 (N_3360,N_3044,N_3100);
xnor U3361 (N_3361,N_3135,N_3038);
xnor U3362 (N_3362,N_3036,N_3154);
or U3363 (N_3363,N_3068,N_3059);
or U3364 (N_3364,N_3131,N_3197);
and U3365 (N_3365,N_3198,N_3005);
and U3366 (N_3366,N_3029,N_3174);
nand U3367 (N_3367,N_3049,N_3087);
nor U3368 (N_3368,N_3022,N_3036);
xor U3369 (N_3369,N_3010,N_3169);
or U3370 (N_3370,N_3101,N_3069);
and U3371 (N_3371,N_3029,N_3050);
nand U3372 (N_3372,N_3154,N_3086);
xnor U3373 (N_3373,N_3007,N_3176);
nor U3374 (N_3374,N_3030,N_3089);
xor U3375 (N_3375,N_3034,N_3001);
xor U3376 (N_3376,N_3090,N_3111);
nor U3377 (N_3377,N_3106,N_3117);
or U3378 (N_3378,N_3009,N_3042);
and U3379 (N_3379,N_3046,N_3018);
nand U3380 (N_3380,N_3081,N_3138);
and U3381 (N_3381,N_3117,N_3123);
nor U3382 (N_3382,N_3020,N_3019);
xor U3383 (N_3383,N_3053,N_3146);
nor U3384 (N_3384,N_3102,N_3159);
or U3385 (N_3385,N_3143,N_3099);
nand U3386 (N_3386,N_3047,N_3019);
xor U3387 (N_3387,N_3150,N_3141);
xnor U3388 (N_3388,N_3180,N_3150);
xnor U3389 (N_3389,N_3199,N_3197);
xor U3390 (N_3390,N_3158,N_3112);
and U3391 (N_3391,N_3191,N_3089);
and U3392 (N_3392,N_3129,N_3177);
and U3393 (N_3393,N_3182,N_3007);
xnor U3394 (N_3394,N_3159,N_3189);
nor U3395 (N_3395,N_3025,N_3013);
xnor U3396 (N_3396,N_3019,N_3017);
xor U3397 (N_3397,N_3044,N_3162);
nor U3398 (N_3398,N_3013,N_3112);
nand U3399 (N_3399,N_3040,N_3014);
and U3400 (N_3400,N_3360,N_3240);
nor U3401 (N_3401,N_3338,N_3273);
and U3402 (N_3402,N_3383,N_3297);
xor U3403 (N_3403,N_3361,N_3371);
and U3404 (N_3404,N_3366,N_3239);
or U3405 (N_3405,N_3204,N_3304);
and U3406 (N_3406,N_3315,N_3327);
xor U3407 (N_3407,N_3272,N_3269);
nand U3408 (N_3408,N_3345,N_3339);
xnor U3409 (N_3409,N_3323,N_3291);
nand U3410 (N_3410,N_3265,N_3391);
nand U3411 (N_3411,N_3217,N_3222);
or U3412 (N_3412,N_3318,N_3280);
or U3413 (N_3413,N_3210,N_3375);
nand U3414 (N_3414,N_3238,N_3229);
and U3415 (N_3415,N_3313,N_3295);
nor U3416 (N_3416,N_3247,N_3373);
nand U3417 (N_3417,N_3336,N_3209);
nand U3418 (N_3418,N_3274,N_3332);
xor U3419 (N_3419,N_3224,N_3270);
or U3420 (N_3420,N_3281,N_3250);
or U3421 (N_3421,N_3330,N_3215);
or U3422 (N_3422,N_3368,N_3254);
nor U3423 (N_3423,N_3214,N_3328);
xnor U3424 (N_3424,N_3341,N_3379);
nor U3425 (N_3425,N_3311,N_3301);
xnor U3426 (N_3426,N_3326,N_3230);
and U3427 (N_3427,N_3267,N_3242);
and U3428 (N_3428,N_3226,N_3305);
and U3429 (N_3429,N_3351,N_3282);
nor U3430 (N_3430,N_3329,N_3294);
nor U3431 (N_3431,N_3275,N_3314);
nand U3432 (N_3432,N_3237,N_3356);
and U3433 (N_3433,N_3389,N_3212);
xor U3434 (N_3434,N_3335,N_3298);
or U3435 (N_3435,N_3216,N_3349);
nand U3436 (N_3436,N_3380,N_3261);
xor U3437 (N_3437,N_3398,N_3394);
and U3438 (N_3438,N_3259,N_3288);
and U3439 (N_3439,N_3296,N_3202);
xnor U3440 (N_3440,N_3344,N_3231);
xnor U3441 (N_3441,N_3221,N_3350);
or U3442 (N_3442,N_3365,N_3369);
or U3443 (N_3443,N_3255,N_3355);
nand U3444 (N_3444,N_3225,N_3319);
or U3445 (N_3445,N_3264,N_3310);
or U3446 (N_3446,N_3299,N_3300);
and U3447 (N_3447,N_3354,N_3363);
and U3448 (N_3448,N_3285,N_3279);
nand U3449 (N_3449,N_3289,N_3219);
nand U3450 (N_3450,N_3359,N_3200);
nor U3451 (N_3451,N_3367,N_3251);
xor U3452 (N_3452,N_3347,N_3331);
xor U3453 (N_3453,N_3384,N_3207);
xor U3454 (N_3454,N_3358,N_3244);
or U3455 (N_3455,N_3243,N_3286);
or U3456 (N_3456,N_3324,N_3306);
nand U3457 (N_3457,N_3309,N_3208);
xnor U3458 (N_3458,N_3357,N_3223);
xor U3459 (N_3459,N_3337,N_3290);
or U3460 (N_3460,N_3346,N_3257);
xor U3461 (N_3461,N_3283,N_3340);
or U3462 (N_3462,N_3388,N_3308);
or U3463 (N_3463,N_3271,N_3312);
nand U3464 (N_3464,N_3378,N_3236);
or U3465 (N_3465,N_3235,N_3232);
xnor U3466 (N_3466,N_3348,N_3343);
xor U3467 (N_3467,N_3317,N_3386);
xnor U3468 (N_3468,N_3320,N_3382);
or U3469 (N_3469,N_3253,N_3376);
nand U3470 (N_3470,N_3396,N_3262);
nor U3471 (N_3471,N_3353,N_3241);
xnor U3472 (N_3472,N_3260,N_3390);
xor U3473 (N_3473,N_3256,N_3284);
xor U3474 (N_3474,N_3372,N_3233);
nor U3475 (N_3475,N_3213,N_3364);
nor U3476 (N_3476,N_3205,N_3248);
xor U3477 (N_3477,N_3227,N_3392);
or U3478 (N_3478,N_3316,N_3206);
nand U3479 (N_3479,N_3292,N_3276);
nor U3480 (N_3480,N_3321,N_3377);
or U3481 (N_3481,N_3249,N_3287);
nor U3482 (N_3482,N_3220,N_3374);
nand U3483 (N_3483,N_3395,N_3263);
nor U3484 (N_3484,N_3352,N_3268);
xor U3485 (N_3485,N_3293,N_3381);
and U3486 (N_3486,N_3307,N_3399);
xor U3487 (N_3487,N_3266,N_3278);
xnor U3488 (N_3488,N_3385,N_3218);
and U3489 (N_3489,N_3370,N_3277);
nand U3490 (N_3490,N_3325,N_3203);
and U3491 (N_3491,N_3342,N_3397);
and U3492 (N_3492,N_3211,N_3333);
nor U3493 (N_3493,N_3201,N_3362);
nand U3494 (N_3494,N_3302,N_3334);
and U3495 (N_3495,N_3246,N_3252);
or U3496 (N_3496,N_3322,N_3393);
nor U3497 (N_3497,N_3228,N_3387);
or U3498 (N_3498,N_3303,N_3245);
nand U3499 (N_3499,N_3234,N_3258);
and U3500 (N_3500,N_3252,N_3203);
or U3501 (N_3501,N_3218,N_3397);
and U3502 (N_3502,N_3366,N_3284);
nor U3503 (N_3503,N_3202,N_3320);
xnor U3504 (N_3504,N_3366,N_3357);
xnor U3505 (N_3505,N_3223,N_3206);
or U3506 (N_3506,N_3355,N_3225);
or U3507 (N_3507,N_3264,N_3280);
and U3508 (N_3508,N_3324,N_3332);
nor U3509 (N_3509,N_3308,N_3337);
nor U3510 (N_3510,N_3360,N_3386);
xor U3511 (N_3511,N_3356,N_3302);
nor U3512 (N_3512,N_3224,N_3251);
and U3513 (N_3513,N_3212,N_3286);
nor U3514 (N_3514,N_3255,N_3230);
or U3515 (N_3515,N_3238,N_3213);
or U3516 (N_3516,N_3397,N_3325);
or U3517 (N_3517,N_3254,N_3235);
xor U3518 (N_3518,N_3322,N_3327);
xor U3519 (N_3519,N_3322,N_3399);
or U3520 (N_3520,N_3290,N_3281);
and U3521 (N_3521,N_3350,N_3379);
xnor U3522 (N_3522,N_3343,N_3396);
and U3523 (N_3523,N_3232,N_3397);
nand U3524 (N_3524,N_3323,N_3370);
and U3525 (N_3525,N_3242,N_3364);
nor U3526 (N_3526,N_3205,N_3245);
nand U3527 (N_3527,N_3367,N_3210);
nor U3528 (N_3528,N_3293,N_3296);
xor U3529 (N_3529,N_3379,N_3293);
nor U3530 (N_3530,N_3311,N_3365);
nand U3531 (N_3531,N_3277,N_3281);
xnor U3532 (N_3532,N_3344,N_3356);
and U3533 (N_3533,N_3345,N_3356);
or U3534 (N_3534,N_3373,N_3261);
and U3535 (N_3535,N_3231,N_3220);
and U3536 (N_3536,N_3313,N_3271);
and U3537 (N_3537,N_3275,N_3239);
xnor U3538 (N_3538,N_3257,N_3205);
and U3539 (N_3539,N_3304,N_3280);
xnor U3540 (N_3540,N_3288,N_3308);
or U3541 (N_3541,N_3270,N_3312);
nand U3542 (N_3542,N_3383,N_3253);
nand U3543 (N_3543,N_3261,N_3277);
or U3544 (N_3544,N_3348,N_3217);
nand U3545 (N_3545,N_3229,N_3222);
nor U3546 (N_3546,N_3294,N_3228);
nor U3547 (N_3547,N_3353,N_3243);
and U3548 (N_3548,N_3206,N_3262);
xnor U3549 (N_3549,N_3337,N_3254);
nor U3550 (N_3550,N_3230,N_3398);
and U3551 (N_3551,N_3229,N_3390);
xnor U3552 (N_3552,N_3236,N_3265);
nand U3553 (N_3553,N_3260,N_3265);
nor U3554 (N_3554,N_3272,N_3335);
xor U3555 (N_3555,N_3265,N_3371);
nor U3556 (N_3556,N_3322,N_3364);
xnor U3557 (N_3557,N_3360,N_3328);
or U3558 (N_3558,N_3224,N_3282);
or U3559 (N_3559,N_3218,N_3311);
xnor U3560 (N_3560,N_3259,N_3329);
or U3561 (N_3561,N_3368,N_3237);
nand U3562 (N_3562,N_3282,N_3283);
and U3563 (N_3563,N_3313,N_3209);
nor U3564 (N_3564,N_3276,N_3265);
xnor U3565 (N_3565,N_3381,N_3295);
and U3566 (N_3566,N_3332,N_3364);
nand U3567 (N_3567,N_3271,N_3249);
nand U3568 (N_3568,N_3339,N_3241);
xnor U3569 (N_3569,N_3227,N_3212);
nand U3570 (N_3570,N_3321,N_3250);
xnor U3571 (N_3571,N_3370,N_3394);
xnor U3572 (N_3572,N_3395,N_3335);
or U3573 (N_3573,N_3295,N_3352);
and U3574 (N_3574,N_3225,N_3334);
xnor U3575 (N_3575,N_3242,N_3299);
nor U3576 (N_3576,N_3259,N_3317);
or U3577 (N_3577,N_3340,N_3240);
or U3578 (N_3578,N_3212,N_3325);
nor U3579 (N_3579,N_3205,N_3261);
nor U3580 (N_3580,N_3343,N_3326);
or U3581 (N_3581,N_3295,N_3364);
or U3582 (N_3582,N_3233,N_3263);
nor U3583 (N_3583,N_3269,N_3302);
xor U3584 (N_3584,N_3277,N_3254);
nand U3585 (N_3585,N_3270,N_3358);
or U3586 (N_3586,N_3211,N_3341);
and U3587 (N_3587,N_3210,N_3267);
xnor U3588 (N_3588,N_3381,N_3226);
and U3589 (N_3589,N_3298,N_3267);
nand U3590 (N_3590,N_3343,N_3308);
and U3591 (N_3591,N_3343,N_3223);
nor U3592 (N_3592,N_3231,N_3355);
xnor U3593 (N_3593,N_3294,N_3248);
or U3594 (N_3594,N_3291,N_3283);
xor U3595 (N_3595,N_3396,N_3293);
xnor U3596 (N_3596,N_3356,N_3245);
or U3597 (N_3597,N_3258,N_3319);
nor U3598 (N_3598,N_3299,N_3308);
or U3599 (N_3599,N_3354,N_3373);
nor U3600 (N_3600,N_3527,N_3541);
xnor U3601 (N_3601,N_3469,N_3487);
or U3602 (N_3602,N_3550,N_3587);
or U3603 (N_3603,N_3558,N_3493);
nand U3604 (N_3604,N_3422,N_3444);
nand U3605 (N_3605,N_3472,N_3521);
nand U3606 (N_3606,N_3583,N_3446);
and U3607 (N_3607,N_3442,N_3426);
nor U3608 (N_3608,N_3554,N_3596);
and U3609 (N_3609,N_3559,N_3407);
nand U3610 (N_3610,N_3423,N_3485);
nor U3611 (N_3611,N_3565,N_3402);
or U3612 (N_3612,N_3477,N_3589);
nor U3613 (N_3613,N_3495,N_3547);
xnor U3614 (N_3614,N_3403,N_3525);
xnor U3615 (N_3615,N_3517,N_3597);
xnor U3616 (N_3616,N_3510,N_3545);
or U3617 (N_3617,N_3464,N_3482);
nor U3618 (N_3618,N_3511,N_3453);
and U3619 (N_3619,N_3534,N_3552);
xor U3620 (N_3620,N_3471,N_3501);
nand U3621 (N_3621,N_3484,N_3513);
and U3622 (N_3622,N_3543,N_3439);
xnor U3623 (N_3623,N_3479,N_3451);
xor U3624 (N_3624,N_3560,N_3557);
nand U3625 (N_3625,N_3506,N_3419);
nor U3626 (N_3626,N_3567,N_3467);
nor U3627 (N_3627,N_3412,N_3432);
xor U3628 (N_3628,N_3413,N_3406);
nor U3629 (N_3629,N_3433,N_3519);
nand U3630 (N_3630,N_3490,N_3505);
and U3631 (N_3631,N_3509,N_3568);
xnor U3632 (N_3632,N_3494,N_3458);
or U3633 (N_3633,N_3496,N_3500);
nand U3634 (N_3634,N_3438,N_3538);
xnor U3635 (N_3635,N_3514,N_3572);
and U3636 (N_3636,N_3425,N_3473);
xnor U3637 (N_3637,N_3595,N_3566);
or U3638 (N_3638,N_3470,N_3441);
nand U3639 (N_3639,N_3497,N_3481);
and U3640 (N_3640,N_3588,N_3544);
xnor U3641 (N_3641,N_3591,N_3416);
nor U3642 (N_3642,N_3575,N_3524);
nor U3643 (N_3643,N_3449,N_3551);
nand U3644 (N_3644,N_3576,N_3401);
xor U3645 (N_3645,N_3448,N_3578);
or U3646 (N_3646,N_3593,N_3502);
nand U3647 (N_3647,N_3599,N_3431);
nand U3648 (N_3648,N_3491,N_3592);
nor U3649 (N_3649,N_3580,N_3415);
or U3650 (N_3650,N_3535,N_3480);
and U3651 (N_3651,N_3455,N_3492);
nor U3652 (N_3652,N_3499,N_3507);
nand U3653 (N_3653,N_3555,N_3563);
xor U3654 (N_3654,N_3447,N_3574);
xor U3655 (N_3655,N_3435,N_3585);
and U3656 (N_3656,N_3584,N_3581);
xor U3657 (N_3657,N_3421,N_3504);
nand U3658 (N_3658,N_3465,N_3440);
or U3659 (N_3659,N_3410,N_3540);
and U3660 (N_3660,N_3582,N_3520);
xnor U3661 (N_3661,N_3549,N_3474);
xnor U3662 (N_3662,N_3548,N_3530);
nand U3663 (N_3663,N_3418,N_3586);
xnor U3664 (N_3664,N_3536,N_3539);
nor U3665 (N_3665,N_3443,N_3411);
nand U3666 (N_3666,N_3461,N_3434);
nor U3667 (N_3667,N_3522,N_3508);
or U3668 (N_3668,N_3428,N_3518);
or U3669 (N_3669,N_3409,N_3590);
and U3670 (N_3670,N_3427,N_3537);
and U3671 (N_3671,N_3476,N_3516);
nand U3672 (N_3672,N_3512,N_3526);
or U3673 (N_3673,N_3478,N_3486);
xnor U3674 (N_3674,N_3503,N_3598);
nor U3675 (N_3675,N_3528,N_3562);
xor U3676 (N_3676,N_3457,N_3561);
or U3677 (N_3677,N_3456,N_3436);
or U3678 (N_3678,N_3414,N_3553);
nor U3679 (N_3679,N_3468,N_3533);
nand U3680 (N_3680,N_3573,N_3569);
or U3681 (N_3681,N_3405,N_3579);
nor U3682 (N_3682,N_3445,N_3523);
and U3683 (N_3683,N_3529,N_3594);
xor U3684 (N_3684,N_3450,N_3498);
nand U3685 (N_3685,N_3408,N_3420);
nor U3686 (N_3686,N_3459,N_3542);
xor U3687 (N_3687,N_3556,N_3571);
and U3688 (N_3688,N_3532,N_3400);
nor U3689 (N_3689,N_3429,N_3570);
nor U3690 (N_3690,N_3546,N_3452);
nor U3691 (N_3691,N_3424,N_3577);
or U3692 (N_3692,N_3454,N_3475);
xnor U3693 (N_3693,N_3460,N_3531);
xnor U3694 (N_3694,N_3483,N_3463);
or U3695 (N_3695,N_3417,N_3430);
or U3696 (N_3696,N_3466,N_3404);
or U3697 (N_3697,N_3515,N_3437);
nand U3698 (N_3698,N_3488,N_3462);
xnor U3699 (N_3699,N_3564,N_3489);
nand U3700 (N_3700,N_3587,N_3420);
and U3701 (N_3701,N_3560,N_3570);
nand U3702 (N_3702,N_3470,N_3459);
and U3703 (N_3703,N_3414,N_3555);
or U3704 (N_3704,N_3496,N_3456);
xnor U3705 (N_3705,N_3585,N_3423);
nand U3706 (N_3706,N_3410,N_3554);
nand U3707 (N_3707,N_3594,N_3504);
or U3708 (N_3708,N_3592,N_3546);
and U3709 (N_3709,N_3561,N_3536);
xor U3710 (N_3710,N_3510,N_3579);
nand U3711 (N_3711,N_3545,N_3574);
nand U3712 (N_3712,N_3537,N_3426);
nor U3713 (N_3713,N_3455,N_3511);
nand U3714 (N_3714,N_3412,N_3544);
and U3715 (N_3715,N_3489,N_3453);
and U3716 (N_3716,N_3416,N_3565);
nor U3717 (N_3717,N_3577,N_3471);
nand U3718 (N_3718,N_3527,N_3597);
nor U3719 (N_3719,N_3535,N_3580);
and U3720 (N_3720,N_3527,N_3513);
and U3721 (N_3721,N_3434,N_3531);
nor U3722 (N_3722,N_3543,N_3422);
nand U3723 (N_3723,N_3500,N_3423);
and U3724 (N_3724,N_3542,N_3463);
nand U3725 (N_3725,N_3557,N_3405);
nor U3726 (N_3726,N_3487,N_3413);
xnor U3727 (N_3727,N_3422,N_3498);
nor U3728 (N_3728,N_3411,N_3402);
or U3729 (N_3729,N_3576,N_3463);
or U3730 (N_3730,N_3503,N_3560);
or U3731 (N_3731,N_3407,N_3493);
nand U3732 (N_3732,N_3485,N_3424);
xor U3733 (N_3733,N_3439,N_3502);
and U3734 (N_3734,N_3560,N_3466);
nand U3735 (N_3735,N_3481,N_3454);
or U3736 (N_3736,N_3485,N_3466);
or U3737 (N_3737,N_3507,N_3560);
xnor U3738 (N_3738,N_3465,N_3497);
nor U3739 (N_3739,N_3498,N_3524);
nor U3740 (N_3740,N_3552,N_3509);
or U3741 (N_3741,N_3569,N_3480);
and U3742 (N_3742,N_3501,N_3585);
and U3743 (N_3743,N_3562,N_3432);
nor U3744 (N_3744,N_3559,N_3594);
or U3745 (N_3745,N_3521,N_3594);
nor U3746 (N_3746,N_3525,N_3533);
xor U3747 (N_3747,N_3586,N_3530);
and U3748 (N_3748,N_3432,N_3539);
nand U3749 (N_3749,N_3499,N_3547);
and U3750 (N_3750,N_3513,N_3518);
nor U3751 (N_3751,N_3505,N_3438);
nor U3752 (N_3752,N_3533,N_3540);
nand U3753 (N_3753,N_3540,N_3580);
or U3754 (N_3754,N_3497,N_3526);
xnor U3755 (N_3755,N_3457,N_3554);
or U3756 (N_3756,N_3404,N_3428);
nor U3757 (N_3757,N_3456,N_3421);
xnor U3758 (N_3758,N_3596,N_3451);
or U3759 (N_3759,N_3422,N_3586);
nor U3760 (N_3760,N_3443,N_3475);
and U3761 (N_3761,N_3543,N_3410);
nor U3762 (N_3762,N_3582,N_3405);
xnor U3763 (N_3763,N_3521,N_3548);
nand U3764 (N_3764,N_3468,N_3566);
and U3765 (N_3765,N_3412,N_3503);
or U3766 (N_3766,N_3404,N_3467);
or U3767 (N_3767,N_3417,N_3491);
and U3768 (N_3768,N_3542,N_3569);
nor U3769 (N_3769,N_3480,N_3412);
nand U3770 (N_3770,N_3544,N_3468);
or U3771 (N_3771,N_3480,N_3470);
and U3772 (N_3772,N_3555,N_3536);
or U3773 (N_3773,N_3488,N_3509);
xnor U3774 (N_3774,N_3588,N_3540);
xnor U3775 (N_3775,N_3438,N_3518);
nor U3776 (N_3776,N_3411,N_3533);
or U3777 (N_3777,N_3515,N_3564);
xnor U3778 (N_3778,N_3502,N_3543);
nand U3779 (N_3779,N_3465,N_3424);
and U3780 (N_3780,N_3457,N_3503);
or U3781 (N_3781,N_3500,N_3491);
and U3782 (N_3782,N_3465,N_3593);
xor U3783 (N_3783,N_3460,N_3406);
nand U3784 (N_3784,N_3465,N_3506);
or U3785 (N_3785,N_3579,N_3530);
nor U3786 (N_3786,N_3517,N_3478);
nand U3787 (N_3787,N_3422,N_3431);
or U3788 (N_3788,N_3543,N_3408);
xor U3789 (N_3789,N_3523,N_3521);
and U3790 (N_3790,N_3545,N_3541);
nand U3791 (N_3791,N_3542,N_3588);
xnor U3792 (N_3792,N_3522,N_3416);
xnor U3793 (N_3793,N_3549,N_3550);
nand U3794 (N_3794,N_3430,N_3540);
nor U3795 (N_3795,N_3588,N_3441);
xor U3796 (N_3796,N_3460,N_3501);
nor U3797 (N_3797,N_3506,N_3578);
nand U3798 (N_3798,N_3575,N_3526);
nand U3799 (N_3799,N_3528,N_3571);
nor U3800 (N_3800,N_3646,N_3749);
xnor U3801 (N_3801,N_3756,N_3742);
or U3802 (N_3802,N_3785,N_3625);
xor U3803 (N_3803,N_3763,N_3663);
or U3804 (N_3804,N_3626,N_3620);
nor U3805 (N_3805,N_3787,N_3707);
or U3806 (N_3806,N_3634,N_3619);
nand U3807 (N_3807,N_3669,N_3641);
or U3808 (N_3808,N_3798,N_3685);
and U3809 (N_3809,N_3613,N_3792);
nor U3810 (N_3810,N_3696,N_3778);
nand U3811 (N_3811,N_3672,N_3608);
xor U3812 (N_3812,N_3782,N_3727);
xnor U3813 (N_3813,N_3795,N_3653);
or U3814 (N_3814,N_3766,N_3793);
nand U3815 (N_3815,N_3693,N_3665);
nand U3816 (N_3816,N_3605,N_3691);
xnor U3817 (N_3817,N_3730,N_3639);
or U3818 (N_3818,N_3768,N_3703);
nand U3819 (N_3819,N_3616,N_3751);
nor U3820 (N_3820,N_3681,N_3697);
and U3821 (N_3821,N_3640,N_3732);
nor U3822 (N_3822,N_3773,N_3791);
or U3823 (N_3823,N_3661,N_3740);
nand U3824 (N_3824,N_3704,N_3638);
or U3825 (N_3825,N_3624,N_3769);
xor U3826 (N_3826,N_3666,N_3673);
nor U3827 (N_3827,N_3713,N_3741);
xor U3828 (N_3828,N_3654,N_3761);
or U3829 (N_3829,N_3614,N_3746);
nor U3830 (N_3830,N_3794,N_3676);
nand U3831 (N_3831,N_3757,N_3658);
or U3832 (N_3832,N_3774,N_3758);
nand U3833 (N_3833,N_3765,N_3701);
and U3834 (N_3834,N_3683,N_3747);
nand U3835 (N_3835,N_3627,N_3799);
xnor U3836 (N_3836,N_3790,N_3726);
or U3837 (N_3837,N_3680,N_3717);
and U3838 (N_3838,N_3686,N_3621);
xnor U3839 (N_3839,N_3731,N_3650);
nor U3840 (N_3840,N_3737,N_3622);
and U3841 (N_3841,N_3753,N_3667);
xnor U3842 (N_3842,N_3720,N_3648);
and U3843 (N_3843,N_3702,N_3644);
nor U3844 (N_3844,N_3698,N_3722);
or U3845 (N_3845,N_3700,N_3776);
xnor U3846 (N_3846,N_3652,N_3786);
nor U3847 (N_3847,N_3601,N_3762);
nor U3848 (N_3848,N_3617,N_3796);
xor U3849 (N_3849,N_3708,N_3725);
xor U3850 (N_3850,N_3739,N_3692);
xnor U3851 (N_3851,N_3689,N_3662);
nor U3852 (N_3852,N_3743,N_3682);
or U3853 (N_3853,N_3656,N_3750);
and U3854 (N_3854,N_3715,N_3609);
nor U3855 (N_3855,N_3699,N_3760);
or U3856 (N_3856,N_3735,N_3771);
xor U3857 (N_3857,N_3607,N_3779);
nor U3858 (N_3858,N_3714,N_3695);
xor U3859 (N_3859,N_3612,N_3675);
or U3860 (N_3860,N_3629,N_3755);
or U3861 (N_3861,N_3719,N_3690);
nor U3862 (N_3862,N_3674,N_3645);
or U3863 (N_3863,N_3606,N_3679);
or U3864 (N_3864,N_3780,N_3655);
nand U3865 (N_3865,N_3636,N_3604);
nor U3866 (N_3866,N_3712,N_3660);
xnor U3867 (N_3867,N_3671,N_3723);
or U3868 (N_3868,N_3781,N_3688);
or U3869 (N_3869,N_3721,N_3733);
nor U3870 (N_3870,N_3783,N_3738);
or U3871 (N_3871,N_3632,N_3628);
nor U3872 (N_3872,N_3637,N_3684);
nand U3873 (N_3873,N_3777,N_3694);
or U3874 (N_3874,N_3710,N_3752);
nor U3875 (N_3875,N_3724,N_3797);
nand U3876 (N_3876,N_3748,N_3603);
nor U3877 (N_3877,N_3623,N_3759);
and U3878 (N_3878,N_3767,N_3643);
and U3879 (N_3879,N_3630,N_3600);
xnor U3880 (N_3880,N_3631,N_3687);
nand U3881 (N_3881,N_3716,N_3784);
and U3882 (N_3882,N_3775,N_3764);
and U3883 (N_3883,N_3657,N_3678);
nand U3884 (N_3884,N_3788,N_3610);
nand U3885 (N_3885,N_3772,N_3602);
nand U3886 (N_3886,N_3647,N_3729);
or U3887 (N_3887,N_3642,N_3718);
nand U3888 (N_3888,N_3649,N_3728);
nand U3889 (N_3889,N_3615,N_3734);
nor U3890 (N_3890,N_3668,N_3754);
xnor U3891 (N_3891,N_3770,N_3677);
nand U3892 (N_3892,N_3744,N_3736);
xor U3893 (N_3893,N_3618,N_3789);
or U3894 (N_3894,N_3664,N_3635);
nand U3895 (N_3895,N_3745,N_3711);
xor U3896 (N_3896,N_3651,N_3633);
and U3897 (N_3897,N_3611,N_3670);
nor U3898 (N_3898,N_3706,N_3659);
nor U3899 (N_3899,N_3705,N_3709);
nor U3900 (N_3900,N_3712,N_3750);
nor U3901 (N_3901,N_3733,N_3797);
and U3902 (N_3902,N_3710,N_3705);
nor U3903 (N_3903,N_3787,N_3702);
xor U3904 (N_3904,N_3766,N_3603);
nor U3905 (N_3905,N_3775,N_3698);
nor U3906 (N_3906,N_3731,N_3700);
or U3907 (N_3907,N_3606,N_3751);
nor U3908 (N_3908,N_3683,N_3714);
or U3909 (N_3909,N_3773,N_3691);
nor U3910 (N_3910,N_3737,N_3692);
or U3911 (N_3911,N_3743,N_3770);
and U3912 (N_3912,N_3719,N_3715);
or U3913 (N_3913,N_3618,N_3645);
and U3914 (N_3914,N_3716,N_3747);
nor U3915 (N_3915,N_3781,N_3799);
or U3916 (N_3916,N_3679,N_3759);
or U3917 (N_3917,N_3683,N_3663);
nor U3918 (N_3918,N_3624,N_3699);
nand U3919 (N_3919,N_3764,N_3765);
xnor U3920 (N_3920,N_3685,N_3673);
nand U3921 (N_3921,N_3717,N_3771);
xor U3922 (N_3922,N_3788,N_3631);
nand U3923 (N_3923,N_3728,N_3770);
nor U3924 (N_3924,N_3611,N_3729);
nor U3925 (N_3925,N_3726,N_3799);
xnor U3926 (N_3926,N_3634,N_3668);
nand U3927 (N_3927,N_3742,N_3676);
nand U3928 (N_3928,N_3736,N_3785);
nor U3929 (N_3929,N_3683,N_3765);
and U3930 (N_3930,N_3695,N_3669);
nand U3931 (N_3931,N_3703,N_3620);
xor U3932 (N_3932,N_3683,N_3641);
and U3933 (N_3933,N_3635,N_3605);
nand U3934 (N_3934,N_3700,N_3654);
or U3935 (N_3935,N_3741,N_3659);
and U3936 (N_3936,N_3698,N_3660);
nor U3937 (N_3937,N_3698,N_3656);
or U3938 (N_3938,N_3605,N_3681);
nand U3939 (N_3939,N_3738,N_3605);
nor U3940 (N_3940,N_3611,N_3679);
and U3941 (N_3941,N_3783,N_3709);
nand U3942 (N_3942,N_3747,N_3662);
nand U3943 (N_3943,N_3743,N_3785);
and U3944 (N_3944,N_3613,N_3761);
nand U3945 (N_3945,N_3753,N_3652);
nor U3946 (N_3946,N_3673,N_3655);
or U3947 (N_3947,N_3780,N_3742);
nor U3948 (N_3948,N_3789,N_3749);
and U3949 (N_3949,N_3750,N_3742);
xnor U3950 (N_3950,N_3790,N_3688);
xnor U3951 (N_3951,N_3635,N_3681);
nand U3952 (N_3952,N_3733,N_3737);
nor U3953 (N_3953,N_3682,N_3717);
xor U3954 (N_3954,N_3721,N_3710);
xor U3955 (N_3955,N_3648,N_3608);
nor U3956 (N_3956,N_3608,N_3714);
and U3957 (N_3957,N_3676,N_3633);
xor U3958 (N_3958,N_3708,N_3738);
xor U3959 (N_3959,N_3794,N_3698);
nand U3960 (N_3960,N_3770,N_3644);
xor U3961 (N_3961,N_3712,N_3751);
xor U3962 (N_3962,N_3775,N_3781);
or U3963 (N_3963,N_3658,N_3742);
nand U3964 (N_3964,N_3768,N_3736);
nand U3965 (N_3965,N_3671,N_3748);
nand U3966 (N_3966,N_3645,N_3720);
and U3967 (N_3967,N_3678,N_3600);
and U3968 (N_3968,N_3631,N_3612);
and U3969 (N_3969,N_3727,N_3719);
xnor U3970 (N_3970,N_3672,N_3669);
xor U3971 (N_3971,N_3663,N_3791);
or U3972 (N_3972,N_3669,N_3642);
nor U3973 (N_3973,N_3612,N_3740);
xor U3974 (N_3974,N_3782,N_3627);
nand U3975 (N_3975,N_3690,N_3760);
nor U3976 (N_3976,N_3659,N_3778);
nor U3977 (N_3977,N_3794,N_3715);
or U3978 (N_3978,N_3668,N_3691);
and U3979 (N_3979,N_3658,N_3664);
xnor U3980 (N_3980,N_3790,N_3679);
nand U3981 (N_3981,N_3709,N_3664);
nor U3982 (N_3982,N_3609,N_3763);
or U3983 (N_3983,N_3619,N_3776);
or U3984 (N_3984,N_3775,N_3695);
nor U3985 (N_3985,N_3681,N_3618);
xnor U3986 (N_3986,N_3623,N_3723);
nand U3987 (N_3987,N_3736,N_3748);
nand U3988 (N_3988,N_3657,N_3793);
nand U3989 (N_3989,N_3795,N_3702);
nor U3990 (N_3990,N_3785,N_3616);
and U3991 (N_3991,N_3722,N_3653);
and U3992 (N_3992,N_3618,N_3613);
xor U3993 (N_3993,N_3782,N_3737);
nor U3994 (N_3994,N_3787,N_3616);
nor U3995 (N_3995,N_3798,N_3766);
or U3996 (N_3996,N_3624,N_3780);
nand U3997 (N_3997,N_3712,N_3651);
and U3998 (N_3998,N_3643,N_3605);
nor U3999 (N_3999,N_3761,N_3707);
xnor U4000 (N_4000,N_3868,N_3986);
and U4001 (N_4001,N_3992,N_3853);
xnor U4002 (N_4002,N_3894,N_3842);
nand U4003 (N_4003,N_3957,N_3872);
nand U4004 (N_4004,N_3928,N_3899);
or U4005 (N_4005,N_3873,N_3863);
nand U4006 (N_4006,N_3911,N_3877);
xnor U4007 (N_4007,N_3923,N_3821);
nor U4008 (N_4008,N_3801,N_3944);
nand U4009 (N_4009,N_3898,N_3800);
nand U4010 (N_4010,N_3879,N_3999);
nand U4011 (N_4011,N_3883,N_3964);
and U4012 (N_4012,N_3832,N_3869);
nand U4013 (N_4013,N_3948,N_3865);
or U4014 (N_4014,N_3994,N_3808);
and U4015 (N_4015,N_3910,N_3969);
nand U4016 (N_4016,N_3860,N_3933);
nand U4017 (N_4017,N_3830,N_3946);
or U4018 (N_4018,N_3968,N_3841);
nand U4019 (N_4019,N_3955,N_3813);
nand U4020 (N_4020,N_3838,N_3901);
nor U4021 (N_4021,N_3931,N_3812);
and U4022 (N_4022,N_3980,N_3963);
or U4023 (N_4023,N_3936,N_3858);
xnor U4024 (N_4024,N_3851,N_3849);
xnor U4025 (N_4025,N_3837,N_3970);
nand U4026 (N_4026,N_3884,N_3888);
xor U4027 (N_4027,N_3835,N_3861);
xnor U4028 (N_4028,N_3943,N_3902);
and U4029 (N_4029,N_3859,N_3953);
or U4030 (N_4030,N_3976,N_3991);
and U4031 (N_4031,N_3985,N_3839);
or U4032 (N_4032,N_3989,N_3961);
and U4033 (N_4033,N_3965,N_3891);
nand U4034 (N_4034,N_3874,N_3870);
and U4035 (N_4035,N_3803,N_3952);
xnor U4036 (N_4036,N_3862,N_3940);
and U4037 (N_4037,N_3804,N_3833);
and U4038 (N_4038,N_3922,N_3881);
nor U4039 (N_4039,N_3918,N_3896);
xnor U4040 (N_4040,N_3973,N_3807);
xnor U4041 (N_4041,N_3855,N_3904);
or U4042 (N_4042,N_3826,N_3843);
or U4043 (N_4043,N_3834,N_3981);
xor U4044 (N_4044,N_3810,N_3990);
nor U4045 (N_4045,N_3950,N_3856);
nand U4046 (N_4046,N_3959,N_3958);
nor U4047 (N_4047,N_3988,N_3998);
nor U4048 (N_4048,N_3978,N_3903);
nor U4049 (N_4049,N_3895,N_3814);
xor U4050 (N_4050,N_3993,N_3960);
or U4051 (N_4051,N_3915,N_3947);
or U4052 (N_4052,N_3974,N_3997);
nor U4053 (N_4053,N_3930,N_3967);
nor U4054 (N_4054,N_3817,N_3982);
nand U4055 (N_4055,N_3846,N_3913);
nor U4056 (N_4056,N_3905,N_3828);
xor U4057 (N_4057,N_3937,N_3802);
xnor U4058 (N_4058,N_3889,N_3852);
nor U4059 (N_4059,N_3945,N_3847);
and U4060 (N_4060,N_3920,N_3929);
and U4061 (N_4061,N_3823,N_3880);
nand U4062 (N_4062,N_3939,N_3848);
and U4063 (N_4063,N_3926,N_3857);
xor U4064 (N_4064,N_3977,N_3887);
xor U4065 (N_4065,N_3927,N_3854);
nand U4066 (N_4066,N_3819,N_3951);
nor U4067 (N_4067,N_3956,N_3871);
nand U4068 (N_4068,N_3882,N_3935);
or U4069 (N_4069,N_3890,N_3942);
xnor U4070 (N_4070,N_3987,N_3822);
nand U4071 (N_4071,N_3919,N_3972);
nand U4072 (N_4072,N_3995,N_3941);
nand U4073 (N_4073,N_3949,N_3875);
xnor U4074 (N_4074,N_3892,N_3867);
nor U4075 (N_4075,N_3962,N_3809);
or U4076 (N_4076,N_3820,N_3816);
nand U4077 (N_4077,N_3914,N_3916);
and U4078 (N_4078,N_3827,N_3844);
and U4079 (N_4079,N_3912,N_3831);
nand U4080 (N_4080,N_3954,N_3850);
nand U4081 (N_4081,N_3818,N_3924);
nor U4082 (N_4082,N_3909,N_3829);
nor U4083 (N_4083,N_3979,N_3885);
nand U4084 (N_4084,N_3836,N_3845);
and U4085 (N_4085,N_3906,N_3996);
nor U4086 (N_4086,N_3876,N_3975);
xnor U4087 (N_4087,N_3897,N_3938);
nand U4088 (N_4088,N_3805,N_3815);
nor U4089 (N_4089,N_3864,N_3825);
nor U4090 (N_4090,N_3983,N_3900);
nand U4091 (N_4091,N_3908,N_3878);
and U4092 (N_4092,N_3984,N_3925);
or U4093 (N_4093,N_3966,N_3917);
and U4094 (N_4094,N_3840,N_3806);
and U4095 (N_4095,N_3886,N_3921);
nand U4096 (N_4096,N_3934,N_3893);
nor U4097 (N_4097,N_3907,N_3824);
xnor U4098 (N_4098,N_3811,N_3866);
and U4099 (N_4099,N_3971,N_3932);
or U4100 (N_4100,N_3821,N_3807);
and U4101 (N_4101,N_3898,N_3861);
and U4102 (N_4102,N_3854,N_3824);
nand U4103 (N_4103,N_3807,N_3990);
or U4104 (N_4104,N_3889,N_3999);
or U4105 (N_4105,N_3829,N_3821);
and U4106 (N_4106,N_3891,N_3899);
xor U4107 (N_4107,N_3840,N_3996);
nor U4108 (N_4108,N_3963,N_3920);
nor U4109 (N_4109,N_3817,N_3835);
nand U4110 (N_4110,N_3910,N_3847);
nand U4111 (N_4111,N_3998,N_3936);
xor U4112 (N_4112,N_3915,N_3992);
nand U4113 (N_4113,N_3925,N_3901);
or U4114 (N_4114,N_3869,N_3800);
and U4115 (N_4115,N_3944,N_3985);
or U4116 (N_4116,N_3815,N_3975);
or U4117 (N_4117,N_3840,N_3986);
xor U4118 (N_4118,N_3968,N_3829);
nand U4119 (N_4119,N_3959,N_3932);
xnor U4120 (N_4120,N_3997,N_3964);
nand U4121 (N_4121,N_3866,N_3980);
xor U4122 (N_4122,N_3928,N_3971);
nor U4123 (N_4123,N_3968,N_3881);
nand U4124 (N_4124,N_3957,N_3853);
and U4125 (N_4125,N_3965,N_3958);
nand U4126 (N_4126,N_3914,N_3841);
and U4127 (N_4127,N_3826,N_3931);
nand U4128 (N_4128,N_3953,N_3823);
xnor U4129 (N_4129,N_3951,N_3969);
or U4130 (N_4130,N_3807,N_3998);
xnor U4131 (N_4131,N_3939,N_3842);
xnor U4132 (N_4132,N_3966,N_3816);
nor U4133 (N_4133,N_3988,N_3812);
or U4134 (N_4134,N_3912,N_3925);
xnor U4135 (N_4135,N_3904,N_3818);
nor U4136 (N_4136,N_3932,N_3941);
nand U4137 (N_4137,N_3856,N_3850);
xor U4138 (N_4138,N_3929,N_3909);
xor U4139 (N_4139,N_3927,N_3951);
xor U4140 (N_4140,N_3983,N_3836);
xor U4141 (N_4141,N_3809,N_3937);
or U4142 (N_4142,N_3852,N_3803);
and U4143 (N_4143,N_3858,N_3806);
nand U4144 (N_4144,N_3959,N_3859);
and U4145 (N_4145,N_3901,N_3923);
or U4146 (N_4146,N_3844,N_3869);
or U4147 (N_4147,N_3923,N_3879);
nand U4148 (N_4148,N_3871,N_3965);
xnor U4149 (N_4149,N_3831,N_3926);
nor U4150 (N_4150,N_3903,N_3845);
nor U4151 (N_4151,N_3981,N_3845);
nand U4152 (N_4152,N_3845,N_3939);
or U4153 (N_4153,N_3876,N_3863);
and U4154 (N_4154,N_3968,N_3939);
or U4155 (N_4155,N_3903,N_3874);
nand U4156 (N_4156,N_3969,N_3959);
xor U4157 (N_4157,N_3835,N_3865);
nor U4158 (N_4158,N_3975,N_3940);
or U4159 (N_4159,N_3827,N_3977);
xnor U4160 (N_4160,N_3895,N_3998);
xnor U4161 (N_4161,N_3819,N_3938);
nand U4162 (N_4162,N_3898,N_3869);
nor U4163 (N_4163,N_3929,N_3801);
nand U4164 (N_4164,N_3989,N_3990);
and U4165 (N_4165,N_3961,N_3839);
nor U4166 (N_4166,N_3991,N_3923);
nand U4167 (N_4167,N_3985,N_3914);
xor U4168 (N_4168,N_3893,N_3961);
nand U4169 (N_4169,N_3825,N_3827);
or U4170 (N_4170,N_3806,N_3966);
or U4171 (N_4171,N_3831,N_3965);
nor U4172 (N_4172,N_3902,N_3819);
or U4173 (N_4173,N_3846,N_3866);
nand U4174 (N_4174,N_3915,N_3815);
and U4175 (N_4175,N_3914,N_3829);
nor U4176 (N_4176,N_3965,N_3876);
xor U4177 (N_4177,N_3985,N_3806);
xor U4178 (N_4178,N_3893,N_3811);
xor U4179 (N_4179,N_3914,N_3961);
nor U4180 (N_4180,N_3845,N_3950);
nand U4181 (N_4181,N_3875,N_3858);
or U4182 (N_4182,N_3816,N_3980);
nand U4183 (N_4183,N_3943,N_3990);
xor U4184 (N_4184,N_3909,N_3831);
or U4185 (N_4185,N_3999,N_3906);
nor U4186 (N_4186,N_3936,N_3982);
nor U4187 (N_4187,N_3822,N_3914);
and U4188 (N_4188,N_3829,N_3934);
xnor U4189 (N_4189,N_3821,N_3809);
xor U4190 (N_4190,N_3967,N_3842);
nand U4191 (N_4191,N_3889,N_3877);
nand U4192 (N_4192,N_3807,N_3877);
nand U4193 (N_4193,N_3911,N_3957);
and U4194 (N_4194,N_3937,N_3891);
or U4195 (N_4195,N_3960,N_3895);
and U4196 (N_4196,N_3863,N_3889);
nand U4197 (N_4197,N_3801,N_3928);
xnor U4198 (N_4198,N_3872,N_3905);
and U4199 (N_4199,N_3842,N_3837);
nor U4200 (N_4200,N_4142,N_4018);
xnor U4201 (N_4201,N_4053,N_4138);
nor U4202 (N_4202,N_4177,N_4192);
nand U4203 (N_4203,N_4197,N_4143);
xnor U4204 (N_4204,N_4008,N_4175);
nor U4205 (N_4205,N_4186,N_4141);
or U4206 (N_4206,N_4010,N_4048);
or U4207 (N_4207,N_4068,N_4130);
xor U4208 (N_4208,N_4159,N_4161);
nor U4209 (N_4209,N_4043,N_4120);
xnor U4210 (N_4210,N_4178,N_4070);
xor U4211 (N_4211,N_4193,N_4006);
nand U4212 (N_4212,N_4169,N_4049);
nand U4213 (N_4213,N_4113,N_4093);
and U4214 (N_4214,N_4119,N_4144);
nor U4215 (N_4215,N_4027,N_4055);
and U4216 (N_4216,N_4004,N_4089);
nand U4217 (N_4217,N_4162,N_4009);
xor U4218 (N_4218,N_4154,N_4184);
or U4219 (N_4219,N_4107,N_4050);
nor U4220 (N_4220,N_4045,N_4023);
nor U4221 (N_4221,N_4020,N_4137);
or U4222 (N_4222,N_4153,N_4096);
and U4223 (N_4223,N_4033,N_4047);
xnor U4224 (N_4224,N_4035,N_4031);
or U4225 (N_4225,N_4002,N_4052);
xor U4226 (N_4226,N_4110,N_4126);
xnor U4227 (N_4227,N_4109,N_4037);
or U4228 (N_4228,N_4059,N_4040);
xnor U4229 (N_4229,N_4171,N_4058);
xnor U4230 (N_4230,N_4030,N_4098);
and U4231 (N_4231,N_4199,N_4054);
and U4232 (N_4232,N_4191,N_4145);
nor U4233 (N_4233,N_4014,N_4073);
nor U4234 (N_4234,N_4026,N_4083);
nand U4235 (N_4235,N_4124,N_4038);
nand U4236 (N_4236,N_4081,N_4156);
nor U4237 (N_4237,N_4101,N_4129);
or U4238 (N_4238,N_4097,N_4189);
and U4239 (N_4239,N_4003,N_4167);
nand U4240 (N_4240,N_4180,N_4136);
nand U4241 (N_4241,N_4111,N_4194);
and U4242 (N_4242,N_4057,N_4185);
and U4243 (N_4243,N_4132,N_4176);
and U4244 (N_4244,N_4118,N_4072);
or U4245 (N_4245,N_4117,N_4076);
nor U4246 (N_4246,N_4121,N_4032);
nand U4247 (N_4247,N_4179,N_4105);
nand U4248 (N_4248,N_4108,N_4091);
and U4249 (N_4249,N_4034,N_4085);
nor U4250 (N_4250,N_4077,N_4190);
nor U4251 (N_4251,N_4151,N_4087);
and U4252 (N_4252,N_4021,N_4170);
nor U4253 (N_4253,N_4172,N_4041);
nor U4254 (N_4254,N_4084,N_4078);
nand U4255 (N_4255,N_4125,N_4140);
xnor U4256 (N_4256,N_4067,N_4133);
or U4257 (N_4257,N_4075,N_4123);
or U4258 (N_4258,N_4007,N_4086);
xor U4259 (N_4259,N_4149,N_4039);
or U4260 (N_4260,N_4187,N_4104);
or U4261 (N_4261,N_4061,N_4062);
and U4262 (N_4262,N_4155,N_4188);
xnor U4263 (N_4263,N_4135,N_4195);
and U4264 (N_4264,N_4168,N_4024);
or U4265 (N_4265,N_4128,N_4094);
nor U4266 (N_4266,N_4074,N_4051);
nor U4267 (N_4267,N_4147,N_4100);
xor U4268 (N_4268,N_4127,N_4106);
or U4269 (N_4269,N_4166,N_4163);
xor U4270 (N_4270,N_4099,N_4013);
xor U4271 (N_4271,N_4115,N_4016);
and U4272 (N_4272,N_4012,N_4088);
and U4273 (N_4273,N_4146,N_4095);
xor U4274 (N_4274,N_4066,N_4183);
or U4275 (N_4275,N_4000,N_4102);
or U4276 (N_4276,N_4060,N_4182);
xnor U4277 (N_4277,N_4005,N_4064);
nand U4278 (N_4278,N_4131,N_4001);
and U4279 (N_4279,N_4015,N_4157);
xnor U4280 (N_4280,N_4139,N_4112);
and U4281 (N_4281,N_4134,N_4019);
xor U4282 (N_4282,N_4025,N_4063);
nand U4283 (N_4283,N_4181,N_4160);
nor U4284 (N_4284,N_4036,N_4158);
or U4285 (N_4285,N_4029,N_4152);
or U4286 (N_4286,N_4092,N_4173);
or U4287 (N_4287,N_4079,N_4071);
xor U4288 (N_4288,N_4165,N_4198);
nand U4289 (N_4289,N_4090,N_4017);
xor U4290 (N_4290,N_4082,N_4174);
and U4291 (N_4291,N_4011,N_4044);
or U4292 (N_4292,N_4046,N_4042);
xor U4293 (N_4293,N_4164,N_4116);
nand U4294 (N_4294,N_4122,N_4022);
or U4295 (N_4295,N_4114,N_4056);
or U4296 (N_4296,N_4065,N_4069);
and U4297 (N_4297,N_4080,N_4103);
nand U4298 (N_4298,N_4148,N_4150);
and U4299 (N_4299,N_4196,N_4028);
and U4300 (N_4300,N_4109,N_4108);
xor U4301 (N_4301,N_4023,N_4162);
nor U4302 (N_4302,N_4021,N_4169);
nor U4303 (N_4303,N_4111,N_4058);
nand U4304 (N_4304,N_4089,N_4196);
or U4305 (N_4305,N_4158,N_4067);
nand U4306 (N_4306,N_4138,N_4101);
nand U4307 (N_4307,N_4080,N_4076);
nor U4308 (N_4308,N_4058,N_4080);
and U4309 (N_4309,N_4054,N_4127);
or U4310 (N_4310,N_4176,N_4030);
or U4311 (N_4311,N_4023,N_4176);
and U4312 (N_4312,N_4060,N_4107);
nor U4313 (N_4313,N_4143,N_4064);
xnor U4314 (N_4314,N_4097,N_4134);
or U4315 (N_4315,N_4176,N_4035);
or U4316 (N_4316,N_4016,N_4097);
and U4317 (N_4317,N_4171,N_4045);
nand U4318 (N_4318,N_4049,N_4144);
and U4319 (N_4319,N_4114,N_4127);
nand U4320 (N_4320,N_4098,N_4083);
or U4321 (N_4321,N_4057,N_4149);
xor U4322 (N_4322,N_4182,N_4004);
nand U4323 (N_4323,N_4155,N_4109);
and U4324 (N_4324,N_4063,N_4003);
xor U4325 (N_4325,N_4099,N_4058);
nor U4326 (N_4326,N_4018,N_4182);
or U4327 (N_4327,N_4096,N_4176);
nand U4328 (N_4328,N_4079,N_4024);
xnor U4329 (N_4329,N_4016,N_4010);
nand U4330 (N_4330,N_4083,N_4173);
nand U4331 (N_4331,N_4041,N_4068);
xor U4332 (N_4332,N_4133,N_4058);
xnor U4333 (N_4333,N_4152,N_4125);
nor U4334 (N_4334,N_4199,N_4132);
or U4335 (N_4335,N_4088,N_4063);
or U4336 (N_4336,N_4089,N_4126);
xnor U4337 (N_4337,N_4194,N_4158);
xnor U4338 (N_4338,N_4008,N_4131);
or U4339 (N_4339,N_4115,N_4001);
or U4340 (N_4340,N_4156,N_4160);
nor U4341 (N_4341,N_4157,N_4114);
xor U4342 (N_4342,N_4071,N_4084);
and U4343 (N_4343,N_4100,N_4076);
xnor U4344 (N_4344,N_4067,N_4151);
nor U4345 (N_4345,N_4158,N_4087);
xnor U4346 (N_4346,N_4112,N_4039);
nand U4347 (N_4347,N_4096,N_4157);
and U4348 (N_4348,N_4181,N_4142);
or U4349 (N_4349,N_4036,N_4024);
and U4350 (N_4350,N_4022,N_4064);
xnor U4351 (N_4351,N_4067,N_4026);
or U4352 (N_4352,N_4025,N_4135);
xnor U4353 (N_4353,N_4078,N_4188);
nand U4354 (N_4354,N_4176,N_4121);
xnor U4355 (N_4355,N_4058,N_4117);
nor U4356 (N_4356,N_4089,N_4076);
nand U4357 (N_4357,N_4168,N_4027);
nand U4358 (N_4358,N_4040,N_4090);
nand U4359 (N_4359,N_4066,N_4189);
and U4360 (N_4360,N_4171,N_4040);
xnor U4361 (N_4361,N_4111,N_4170);
nor U4362 (N_4362,N_4025,N_4095);
nor U4363 (N_4363,N_4012,N_4038);
or U4364 (N_4364,N_4001,N_4148);
nor U4365 (N_4365,N_4023,N_4104);
nand U4366 (N_4366,N_4163,N_4137);
xor U4367 (N_4367,N_4079,N_4039);
and U4368 (N_4368,N_4023,N_4095);
nor U4369 (N_4369,N_4052,N_4102);
and U4370 (N_4370,N_4172,N_4095);
nand U4371 (N_4371,N_4078,N_4198);
xor U4372 (N_4372,N_4100,N_4192);
xnor U4373 (N_4373,N_4158,N_4165);
nor U4374 (N_4374,N_4138,N_4103);
or U4375 (N_4375,N_4113,N_4110);
xor U4376 (N_4376,N_4173,N_4196);
and U4377 (N_4377,N_4022,N_4165);
or U4378 (N_4378,N_4169,N_4020);
nand U4379 (N_4379,N_4054,N_4070);
and U4380 (N_4380,N_4077,N_4107);
nand U4381 (N_4381,N_4149,N_4158);
nand U4382 (N_4382,N_4175,N_4067);
and U4383 (N_4383,N_4028,N_4065);
and U4384 (N_4384,N_4080,N_4124);
or U4385 (N_4385,N_4005,N_4037);
nand U4386 (N_4386,N_4001,N_4003);
or U4387 (N_4387,N_4025,N_4088);
xor U4388 (N_4388,N_4011,N_4126);
nand U4389 (N_4389,N_4191,N_4072);
or U4390 (N_4390,N_4084,N_4139);
nor U4391 (N_4391,N_4059,N_4122);
nand U4392 (N_4392,N_4159,N_4037);
xor U4393 (N_4393,N_4056,N_4116);
and U4394 (N_4394,N_4111,N_4108);
nor U4395 (N_4395,N_4139,N_4068);
nor U4396 (N_4396,N_4053,N_4066);
or U4397 (N_4397,N_4192,N_4143);
nand U4398 (N_4398,N_4063,N_4149);
or U4399 (N_4399,N_4188,N_4068);
nand U4400 (N_4400,N_4319,N_4367);
nand U4401 (N_4401,N_4255,N_4365);
nand U4402 (N_4402,N_4304,N_4364);
or U4403 (N_4403,N_4337,N_4240);
or U4404 (N_4404,N_4328,N_4234);
or U4405 (N_4405,N_4315,N_4277);
nand U4406 (N_4406,N_4303,N_4370);
nand U4407 (N_4407,N_4276,N_4244);
nand U4408 (N_4408,N_4326,N_4358);
nand U4409 (N_4409,N_4383,N_4300);
xnor U4410 (N_4410,N_4250,N_4271);
nand U4411 (N_4411,N_4248,N_4292);
nor U4412 (N_4412,N_4274,N_4219);
or U4413 (N_4413,N_4395,N_4203);
xor U4414 (N_4414,N_4212,N_4397);
and U4415 (N_4415,N_4293,N_4317);
and U4416 (N_4416,N_4366,N_4216);
nand U4417 (N_4417,N_4392,N_4230);
or U4418 (N_4418,N_4385,N_4312);
nand U4419 (N_4419,N_4362,N_4207);
xor U4420 (N_4420,N_4252,N_4253);
and U4421 (N_4421,N_4265,N_4291);
nor U4422 (N_4422,N_4272,N_4284);
xor U4423 (N_4423,N_4290,N_4285);
nand U4424 (N_4424,N_4247,N_4261);
nand U4425 (N_4425,N_4345,N_4320);
nand U4426 (N_4426,N_4373,N_4393);
and U4427 (N_4427,N_4281,N_4275);
or U4428 (N_4428,N_4308,N_4324);
or U4429 (N_4429,N_4204,N_4218);
nand U4430 (N_4430,N_4347,N_4269);
and U4431 (N_4431,N_4301,N_4283);
nor U4432 (N_4432,N_4237,N_4214);
xor U4433 (N_4433,N_4297,N_4372);
nor U4434 (N_4434,N_4352,N_4399);
or U4435 (N_4435,N_4295,N_4313);
nor U4436 (N_4436,N_4257,N_4354);
xor U4437 (N_4437,N_4348,N_4310);
nand U4438 (N_4438,N_4227,N_4353);
xor U4439 (N_4439,N_4263,N_4318);
or U4440 (N_4440,N_4391,N_4260);
or U4441 (N_4441,N_4384,N_4349);
and U4442 (N_4442,N_4220,N_4242);
nor U4443 (N_4443,N_4251,N_4369);
xnor U4444 (N_4444,N_4254,N_4338);
and U4445 (N_4445,N_4396,N_4217);
nand U4446 (N_4446,N_4279,N_4343);
nor U4447 (N_4447,N_4389,N_4209);
nand U4448 (N_4448,N_4222,N_4316);
and U4449 (N_4449,N_4371,N_4273);
nand U4450 (N_4450,N_4287,N_4229);
and U4451 (N_4451,N_4355,N_4375);
xnor U4452 (N_4452,N_4238,N_4333);
or U4453 (N_4453,N_4201,N_4330);
and U4454 (N_4454,N_4381,N_4382);
nor U4455 (N_4455,N_4344,N_4243);
xor U4456 (N_4456,N_4377,N_4379);
nor U4457 (N_4457,N_4334,N_4305);
nand U4458 (N_4458,N_4278,N_4233);
xnor U4459 (N_4459,N_4258,N_4256);
and U4460 (N_4460,N_4341,N_4306);
xor U4461 (N_4461,N_4359,N_4378);
or U4462 (N_4462,N_4299,N_4331);
nand U4463 (N_4463,N_4246,N_4245);
and U4464 (N_4464,N_4363,N_4327);
and U4465 (N_4465,N_4374,N_4267);
and U4466 (N_4466,N_4224,N_4208);
and U4467 (N_4467,N_4228,N_4323);
xnor U4468 (N_4468,N_4236,N_4280);
xor U4469 (N_4469,N_4332,N_4206);
nand U4470 (N_4470,N_4262,N_4322);
or U4471 (N_4471,N_4289,N_4351);
or U4472 (N_4472,N_4336,N_4211);
and U4473 (N_4473,N_4270,N_4249);
xor U4474 (N_4474,N_4213,N_4232);
nand U4475 (N_4475,N_4298,N_4210);
nand U4476 (N_4476,N_4239,N_4311);
or U4477 (N_4477,N_4390,N_4225);
xnor U4478 (N_4478,N_4205,N_4226);
xnor U4479 (N_4479,N_4350,N_4266);
nand U4480 (N_4480,N_4259,N_4264);
nand U4481 (N_4481,N_4286,N_4376);
and U4482 (N_4482,N_4380,N_4202);
and U4483 (N_4483,N_4294,N_4329);
or U4484 (N_4484,N_4325,N_4302);
or U4485 (N_4485,N_4241,N_4387);
nor U4486 (N_4486,N_4388,N_4282);
xnor U4487 (N_4487,N_4360,N_4235);
nand U4488 (N_4488,N_4368,N_4335);
and U4489 (N_4489,N_4288,N_4340);
nand U4490 (N_4490,N_4398,N_4339);
nand U4491 (N_4491,N_4314,N_4268);
xor U4492 (N_4492,N_4215,N_4357);
xor U4493 (N_4493,N_4361,N_4307);
nand U4494 (N_4494,N_4394,N_4223);
xor U4495 (N_4495,N_4231,N_4342);
and U4496 (N_4496,N_4309,N_4221);
nor U4497 (N_4497,N_4321,N_4346);
nand U4498 (N_4498,N_4356,N_4386);
or U4499 (N_4499,N_4200,N_4296);
nor U4500 (N_4500,N_4302,N_4385);
or U4501 (N_4501,N_4278,N_4291);
nor U4502 (N_4502,N_4265,N_4249);
and U4503 (N_4503,N_4236,N_4293);
and U4504 (N_4504,N_4282,N_4323);
xnor U4505 (N_4505,N_4376,N_4378);
xnor U4506 (N_4506,N_4286,N_4398);
nand U4507 (N_4507,N_4378,N_4319);
or U4508 (N_4508,N_4381,N_4300);
and U4509 (N_4509,N_4287,N_4392);
nand U4510 (N_4510,N_4200,N_4315);
xor U4511 (N_4511,N_4225,N_4366);
nand U4512 (N_4512,N_4376,N_4353);
nor U4513 (N_4513,N_4319,N_4371);
and U4514 (N_4514,N_4391,N_4247);
nor U4515 (N_4515,N_4241,N_4341);
or U4516 (N_4516,N_4283,N_4221);
or U4517 (N_4517,N_4271,N_4213);
nand U4518 (N_4518,N_4395,N_4391);
or U4519 (N_4519,N_4238,N_4326);
and U4520 (N_4520,N_4295,N_4253);
nand U4521 (N_4521,N_4240,N_4362);
or U4522 (N_4522,N_4350,N_4395);
nor U4523 (N_4523,N_4284,N_4270);
and U4524 (N_4524,N_4269,N_4382);
and U4525 (N_4525,N_4379,N_4365);
xor U4526 (N_4526,N_4280,N_4242);
nand U4527 (N_4527,N_4337,N_4225);
and U4528 (N_4528,N_4353,N_4216);
nand U4529 (N_4529,N_4294,N_4286);
or U4530 (N_4530,N_4277,N_4290);
nor U4531 (N_4531,N_4279,N_4219);
xnor U4532 (N_4532,N_4337,N_4202);
nor U4533 (N_4533,N_4288,N_4259);
xnor U4534 (N_4534,N_4233,N_4287);
or U4535 (N_4535,N_4315,N_4233);
and U4536 (N_4536,N_4383,N_4313);
and U4537 (N_4537,N_4317,N_4267);
xnor U4538 (N_4538,N_4244,N_4334);
and U4539 (N_4539,N_4219,N_4321);
xnor U4540 (N_4540,N_4207,N_4237);
nor U4541 (N_4541,N_4242,N_4264);
nand U4542 (N_4542,N_4314,N_4317);
or U4543 (N_4543,N_4360,N_4309);
xor U4544 (N_4544,N_4273,N_4274);
xor U4545 (N_4545,N_4352,N_4307);
nor U4546 (N_4546,N_4394,N_4235);
nand U4547 (N_4547,N_4238,N_4206);
and U4548 (N_4548,N_4343,N_4231);
nor U4549 (N_4549,N_4336,N_4355);
and U4550 (N_4550,N_4381,N_4263);
nand U4551 (N_4551,N_4389,N_4382);
nand U4552 (N_4552,N_4217,N_4290);
nor U4553 (N_4553,N_4270,N_4253);
xor U4554 (N_4554,N_4338,N_4305);
nor U4555 (N_4555,N_4250,N_4244);
nand U4556 (N_4556,N_4327,N_4226);
and U4557 (N_4557,N_4265,N_4362);
and U4558 (N_4558,N_4263,N_4388);
or U4559 (N_4559,N_4258,N_4210);
nor U4560 (N_4560,N_4228,N_4243);
nand U4561 (N_4561,N_4369,N_4380);
nor U4562 (N_4562,N_4211,N_4251);
and U4563 (N_4563,N_4283,N_4234);
nor U4564 (N_4564,N_4233,N_4220);
or U4565 (N_4565,N_4376,N_4219);
xnor U4566 (N_4566,N_4286,N_4399);
and U4567 (N_4567,N_4252,N_4321);
and U4568 (N_4568,N_4357,N_4205);
or U4569 (N_4569,N_4202,N_4384);
and U4570 (N_4570,N_4308,N_4361);
nand U4571 (N_4571,N_4293,N_4209);
xnor U4572 (N_4572,N_4298,N_4343);
and U4573 (N_4573,N_4243,N_4281);
and U4574 (N_4574,N_4350,N_4325);
nor U4575 (N_4575,N_4261,N_4263);
and U4576 (N_4576,N_4204,N_4327);
and U4577 (N_4577,N_4213,N_4351);
and U4578 (N_4578,N_4308,N_4315);
nor U4579 (N_4579,N_4277,N_4299);
nand U4580 (N_4580,N_4374,N_4216);
xnor U4581 (N_4581,N_4344,N_4382);
or U4582 (N_4582,N_4236,N_4307);
nor U4583 (N_4583,N_4387,N_4265);
nor U4584 (N_4584,N_4308,N_4267);
and U4585 (N_4585,N_4355,N_4224);
nand U4586 (N_4586,N_4220,N_4201);
xnor U4587 (N_4587,N_4314,N_4265);
or U4588 (N_4588,N_4300,N_4295);
and U4589 (N_4589,N_4287,N_4242);
or U4590 (N_4590,N_4364,N_4363);
nand U4591 (N_4591,N_4229,N_4339);
nor U4592 (N_4592,N_4293,N_4224);
or U4593 (N_4593,N_4266,N_4375);
or U4594 (N_4594,N_4389,N_4336);
xor U4595 (N_4595,N_4374,N_4222);
xnor U4596 (N_4596,N_4208,N_4203);
xnor U4597 (N_4597,N_4215,N_4380);
and U4598 (N_4598,N_4268,N_4293);
nor U4599 (N_4599,N_4207,N_4284);
nor U4600 (N_4600,N_4581,N_4448);
nand U4601 (N_4601,N_4546,N_4545);
xnor U4602 (N_4602,N_4404,N_4573);
or U4603 (N_4603,N_4455,N_4419);
nand U4604 (N_4604,N_4489,N_4434);
nor U4605 (N_4605,N_4469,N_4553);
or U4606 (N_4606,N_4454,N_4530);
nor U4607 (N_4607,N_4498,N_4558);
or U4608 (N_4608,N_4430,N_4440);
and U4609 (N_4609,N_4480,N_4538);
or U4610 (N_4610,N_4598,N_4533);
nor U4611 (N_4611,N_4429,N_4442);
nor U4612 (N_4612,N_4518,N_4524);
nand U4613 (N_4613,N_4554,N_4536);
nor U4614 (N_4614,N_4453,N_4523);
or U4615 (N_4615,N_4468,N_4574);
or U4616 (N_4616,N_4499,N_4487);
xor U4617 (N_4617,N_4561,N_4551);
xnor U4618 (N_4618,N_4583,N_4472);
nor U4619 (N_4619,N_4496,N_4566);
and U4620 (N_4620,N_4542,N_4527);
nor U4621 (N_4621,N_4432,N_4426);
nor U4622 (N_4622,N_4579,N_4405);
or U4623 (N_4623,N_4486,N_4417);
and U4624 (N_4624,N_4540,N_4591);
nor U4625 (N_4625,N_4544,N_4473);
or U4626 (N_4626,N_4441,N_4559);
xnor U4627 (N_4627,N_4503,N_4525);
and U4628 (N_4628,N_4413,N_4431);
and U4629 (N_4629,N_4515,N_4436);
nand U4630 (N_4630,N_4437,N_4521);
nor U4631 (N_4631,N_4476,N_4466);
and U4632 (N_4632,N_4443,N_4531);
xor U4633 (N_4633,N_4578,N_4438);
nor U4634 (N_4634,N_4414,N_4411);
nor U4635 (N_4635,N_4457,N_4460);
nor U4636 (N_4636,N_4497,N_4548);
xnor U4637 (N_4637,N_4526,N_4512);
xnor U4638 (N_4638,N_4439,N_4403);
or U4639 (N_4639,N_4471,N_4433);
and U4640 (N_4640,N_4415,N_4479);
nor U4641 (N_4641,N_4425,N_4456);
or U4642 (N_4642,N_4534,N_4450);
and U4643 (N_4643,N_4597,N_4522);
nand U4644 (N_4644,N_4567,N_4416);
and U4645 (N_4645,N_4402,N_4599);
or U4646 (N_4646,N_4595,N_4513);
xnor U4647 (N_4647,N_4409,N_4474);
or U4648 (N_4648,N_4470,N_4594);
xor U4649 (N_4649,N_4504,N_4463);
xor U4650 (N_4650,N_4461,N_4406);
or U4651 (N_4651,N_4452,N_4401);
nor U4652 (N_4652,N_4537,N_4528);
xor U4653 (N_4653,N_4444,N_4477);
and U4654 (N_4654,N_4507,N_4520);
xor U4655 (N_4655,N_4484,N_4576);
xnor U4656 (N_4656,N_4552,N_4421);
nor U4657 (N_4657,N_4575,N_4502);
nor U4658 (N_4658,N_4410,N_4467);
and U4659 (N_4659,N_4400,N_4509);
or U4660 (N_4660,N_4494,N_4451);
and U4661 (N_4661,N_4535,N_4516);
xnor U4662 (N_4662,N_4582,N_4565);
nor U4663 (N_4663,N_4539,N_4590);
nor U4664 (N_4664,N_4493,N_4510);
or U4665 (N_4665,N_4592,N_4412);
nor U4666 (N_4666,N_4459,N_4418);
nand U4667 (N_4667,N_4596,N_4572);
or U4668 (N_4668,N_4481,N_4571);
or U4669 (N_4669,N_4549,N_4483);
nor U4670 (N_4670,N_4501,N_4495);
or U4671 (N_4671,N_4580,N_4541);
nor U4672 (N_4672,N_4407,N_4475);
or U4673 (N_4673,N_4427,N_4585);
xor U4674 (N_4674,N_4556,N_4500);
or U4675 (N_4675,N_4508,N_4555);
xnor U4676 (N_4676,N_4505,N_4420);
xnor U4677 (N_4677,N_4593,N_4446);
xnor U4678 (N_4678,N_4488,N_4532);
nand U4679 (N_4679,N_4449,N_4464);
or U4680 (N_4680,N_4577,N_4422);
or U4681 (N_4681,N_4424,N_4447);
nor U4682 (N_4682,N_4445,N_4519);
or U4683 (N_4683,N_4511,N_4529);
and U4684 (N_4684,N_4482,N_4589);
nor U4685 (N_4685,N_4492,N_4435);
and U4686 (N_4686,N_4408,N_4560);
or U4687 (N_4687,N_4557,N_4563);
or U4688 (N_4688,N_4543,N_4514);
xor U4689 (N_4689,N_4428,N_4462);
xor U4690 (N_4690,N_4478,N_4587);
or U4691 (N_4691,N_4485,N_4586);
or U4692 (N_4692,N_4465,N_4550);
xnor U4693 (N_4693,N_4562,N_4588);
xor U4694 (N_4694,N_4490,N_4491);
nand U4695 (N_4695,N_4569,N_4547);
xnor U4696 (N_4696,N_4506,N_4564);
nor U4697 (N_4697,N_4423,N_4584);
nor U4698 (N_4698,N_4517,N_4458);
nand U4699 (N_4699,N_4568,N_4570);
or U4700 (N_4700,N_4585,N_4547);
xor U4701 (N_4701,N_4437,N_4547);
nand U4702 (N_4702,N_4486,N_4592);
nand U4703 (N_4703,N_4445,N_4571);
nand U4704 (N_4704,N_4487,N_4400);
and U4705 (N_4705,N_4577,N_4435);
nor U4706 (N_4706,N_4440,N_4490);
nand U4707 (N_4707,N_4542,N_4490);
nand U4708 (N_4708,N_4500,N_4490);
nor U4709 (N_4709,N_4402,N_4481);
or U4710 (N_4710,N_4441,N_4446);
or U4711 (N_4711,N_4512,N_4445);
nor U4712 (N_4712,N_4446,N_4507);
nand U4713 (N_4713,N_4471,N_4566);
and U4714 (N_4714,N_4566,N_4440);
nand U4715 (N_4715,N_4536,N_4564);
and U4716 (N_4716,N_4584,N_4469);
nor U4717 (N_4717,N_4585,N_4545);
and U4718 (N_4718,N_4565,N_4581);
or U4719 (N_4719,N_4480,N_4515);
xor U4720 (N_4720,N_4554,N_4599);
and U4721 (N_4721,N_4509,N_4457);
nor U4722 (N_4722,N_4562,N_4536);
and U4723 (N_4723,N_4489,N_4548);
nand U4724 (N_4724,N_4455,N_4450);
nor U4725 (N_4725,N_4550,N_4426);
nor U4726 (N_4726,N_4525,N_4407);
and U4727 (N_4727,N_4591,N_4561);
and U4728 (N_4728,N_4505,N_4510);
xor U4729 (N_4729,N_4546,N_4503);
and U4730 (N_4730,N_4466,N_4403);
nand U4731 (N_4731,N_4579,N_4523);
and U4732 (N_4732,N_4497,N_4550);
and U4733 (N_4733,N_4404,N_4412);
or U4734 (N_4734,N_4563,N_4532);
or U4735 (N_4735,N_4526,N_4409);
or U4736 (N_4736,N_4522,N_4450);
or U4737 (N_4737,N_4400,N_4435);
and U4738 (N_4738,N_4596,N_4542);
nand U4739 (N_4739,N_4574,N_4541);
nor U4740 (N_4740,N_4475,N_4587);
xor U4741 (N_4741,N_4420,N_4530);
xor U4742 (N_4742,N_4558,N_4524);
and U4743 (N_4743,N_4586,N_4449);
nor U4744 (N_4744,N_4457,N_4406);
nor U4745 (N_4745,N_4408,N_4451);
nand U4746 (N_4746,N_4491,N_4469);
or U4747 (N_4747,N_4513,N_4538);
nor U4748 (N_4748,N_4514,N_4415);
or U4749 (N_4749,N_4536,N_4413);
xor U4750 (N_4750,N_4408,N_4596);
nor U4751 (N_4751,N_4464,N_4587);
and U4752 (N_4752,N_4584,N_4595);
xnor U4753 (N_4753,N_4572,N_4480);
xor U4754 (N_4754,N_4464,N_4582);
nand U4755 (N_4755,N_4472,N_4532);
nand U4756 (N_4756,N_4425,N_4559);
and U4757 (N_4757,N_4514,N_4465);
and U4758 (N_4758,N_4564,N_4527);
or U4759 (N_4759,N_4560,N_4571);
xnor U4760 (N_4760,N_4589,N_4445);
nor U4761 (N_4761,N_4487,N_4458);
or U4762 (N_4762,N_4425,N_4464);
nor U4763 (N_4763,N_4552,N_4461);
or U4764 (N_4764,N_4499,N_4475);
and U4765 (N_4765,N_4439,N_4575);
or U4766 (N_4766,N_4467,N_4437);
and U4767 (N_4767,N_4531,N_4521);
and U4768 (N_4768,N_4492,N_4563);
xor U4769 (N_4769,N_4461,N_4403);
and U4770 (N_4770,N_4550,N_4568);
and U4771 (N_4771,N_4583,N_4432);
nand U4772 (N_4772,N_4598,N_4572);
nand U4773 (N_4773,N_4481,N_4450);
and U4774 (N_4774,N_4544,N_4493);
or U4775 (N_4775,N_4449,N_4582);
and U4776 (N_4776,N_4567,N_4448);
nand U4777 (N_4777,N_4539,N_4485);
nand U4778 (N_4778,N_4506,N_4493);
xnor U4779 (N_4779,N_4520,N_4529);
or U4780 (N_4780,N_4585,N_4414);
nand U4781 (N_4781,N_4517,N_4530);
or U4782 (N_4782,N_4445,N_4446);
or U4783 (N_4783,N_4419,N_4479);
xnor U4784 (N_4784,N_4542,N_4574);
and U4785 (N_4785,N_4420,N_4443);
or U4786 (N_4786,N_4477,N_4452);
nor U4787 (N_4787,N_4440,N_4552);
nor U4788 (N_4788,N_4475,N_4471);
nand U4789 (N_4789,N_4586,N_4548);
nand U4790 (N_4790,N_4443,N_4570);
or U4791 (N_4791,N_4460,N_4481);
or U4792 (N_4792,N_4471,N_4419);
and U4793 (N_4793,N_4542,N_4450);
nor U4794 (N_4794,N_4555,N_4422);
or U4795 (N_4795,N_4557,N_4473);
nor U4796 (N_4796,N_4571,N_4454);
xor U4797 (N_4797,N_4535,N_4460);
xor U4798 (N_4798,N_4469,N_4447);
or U4799 (N_4799,N_4590,N_4437);
nor U4800 (N_4800,N_4625,N_4605);
and U4801 (N_4801,N_4709,N_4696);
nand U4802 (N_4802,N_4679,N_4737);
or U4803 (N_4803,N_4618,N_4763);
or U4804 (N_4804,N_4684,N_4769);
xor U4805 (N_4805,N_4771,N_4687);
and U4806 (N_4806,N_4702,N_4753);
and U4807 (N_4807,N_4607,N_4766);
nor U4808 (N_4808,N_4700,N_4776);
and U4809 (N_4809,N_4757,N_4641);
or U4810 (N_4810,N_4786,N_4671);
xnor U4811 (N_4811,N_4756,N_4619);
nand U4812 (N_4812,N_4646,N_4699);
or U4813 (N_4813,N_4785,N_4723);
nand U4814 (N_4814,N_4715,N_4666);
xnor U4815 (N_4815,N_4683,N_4634);
xnor U4816 (N_4816,N_4726,N_4639);
or U4817 (N_4817,N_4773,N_4676);
nor U4818 (N_4818,N_4620,N_4770);
and U4819 (N_4819,N_4677,N_4790);
nor U4820 (N_4820,N_4775,N_4791);
nor U4821 (N_4821,N_4701,N_4638);
nand U4822 (N_4822,N_4787,N_4716);
or U4823 (N_4823,N_4792,N_4688);
nand U4824 (N_4824,N_4720,N_4717);
nor U4825 (N_4825,N_4632,N_4784);
or U4826 (N_4826,N_4767,N_4635);
and U4827 (N_4827,N_4602,N_4662);
xnor U4828 (N_4828,N_4779,N_4747);
or U4829 (N_4829,N_4758,N_4660);
and U4830 (N_4830,N_4722,N_4669);
nor U4831 (N_4831,N_4780,N_4690);
or U4832 (N_4832,N_4736,N_4612);
nor U4833 (N_4833,N_4604,N_4713);
nand U4834 (N_4834,N_4682,N_4712);
xnor U4835 (N_4835,N_4661,N_4627);
xor U4836 (N_4836,N_4673,N_4686);
or U4837 (N_4837,N_4628,N_4631);
xnor U4838 (N_4838,N_4630,N_4610);
xor U4839 (N_4839,N_4755,N_4760);
nor U4840 (N_4840,N_4616,N_4796);
xor U4841 (N_4841,N_4691,N_4603);
nor U4842 (N_4842,N_4765,N_4651);
or U4843 (N_4843,N_4733,N_4652);
nand U4844 (N_4844,N_4793,N_4629);
or U4845 (N_4845,N_4740,N_4613);
or U4846 (N_4846,N_4749,N_4768);
and U4847 (N_4847,N_4744,N_4725);
nor U4848 (N_4848,N_4727,N_4781);
xnor U4849 (N_4849,N_4695,N_4729);
nand U4850 (N_4850,N_4777,N_4622);
xnor U4851 (N_4851,N_4647,N_4788);
or U4852 (N_4852,N_4611,N_4642);
nor U4853 (N_4853,N_4693,N_4643);
or U4854 (N_4854,N_4680,N_4746);
nor U4855 (N_4855,N_4694,N_4617);
or U4856 (N_4856,N_4672,N_4658);
nor U4857 (N_4857,N_4745,N_4640);
and U4858 (N_4858,N_4670,N_4730);
or U4859 (N_4859,N_4657,N_4728);
xor U4860 (N_4860,N_4734,N_4752);
nor U4861 (N_4861,N_4664,N_4789);
nor U4862 (N_4862,N_4681,N_4795);
xnor U4863 (N_4863,N_4759,N_4704);
nand U4864 (N_4864,N_4764,N_4719);
nor U4865 (N_4865,N_4678,N_4626);
and U4866 (N_4866,N_4762,N_4637);
or U4867 (N_4867,N_4708,N_4703);
nand U4868 (N_4868,N_4761,N_4675);
nor U4869 (N_4869,N_4606,N_4724);
and U4870 (N_4870,N_4794,N_4706);
and U4871 (N_4871,N_4659,N_4615);
xnor U4872 (N_4872,N_4692,N_4601);
nor U4873 (N_4873,N_4649,N_4707);
nor U4874 (N_4874,N_4689,N_4799);
or U4875 (N_4875,N_4674,N_4624);
and U4876 (N_4876,N_4645,N_4621);
xor U4877 (N_4877,N_4735,N_4668);
nand U4878 (N_4878,N_4714,N_4705);
and U4879 (N_4879,N_4665,N_4623);
and U4880 (N_4880,N_4772,N_4798);
or U4881 (N_4881,N_4663,N_4782);
nand U4882 (N_4882,N_4697,N_4754);
nand U4883 (N_4883,N_4721,N_4711);
and U4884 (N_4884,N_4710,N_4653);
xnor U4885 (N_4885,N_4778,N_4609);
xnor U4886 (N_4886,N_4654,N_4656);
and U4887 (N_4887,N_4614,N_4600);
nor U4888 (N_4888,N_4655,N_4667);
xor U4889 (N_4889,N_4650,N_4742);
xor U4890 (N_4890,N_4774,N_4743);
or U4891 (N_4891,N_4633,N_4718);
xor U4892 (N_4892,N_4783,N_4751);
nor U4893 (N_4893,N_4739,N_4750);
xnor U4894 (N_4894,N_4748,N_4797);
or U4895 (N_4895,N_4698,N_4648);
nand U4896 (N_4896,N_4732,N_4731);
nor U4897 (N_4897,N_4741,N_4644);
or U4898 (N_4898,N_4636,N_4685);
and U4899 (N_4899,N_4608,N_4738);
or U4900 (N_4900,N_4795,N_4642);
and U4901 (N_4901,N_4770,N_4736);
or U4902 (N_4902,N_4684,N_4716);
and U4903 (N_4903,N_4692,N_4714);
nor U4904 (N_4904,N_4726,N_4794);
and U4905 (N_4905,N_4723,N_4763);
xnor U4906 (N_4906,N_4651,N_4638);
or U4907 (N_4907,N_4664,N_4721);
nand U4908 (N_4908,N_4741,N_4713);
and U4909 (N_4909,N_4717,N_4780);
xnor U4910 (N_4910,N_4766,N_4731);
nor U4911 (N_4911,N_4770,N_4779);
nor U4912 (N_4912,N_4756,N_4609);
xnor U4913 (N_4913,N_4792,N_4631);
and U4914 (N_4914,N_4781,N_4701);
nand U4915 (N_4915,N_4670,N_4776);
nand U4916 (N_4916,N_4684,N_4607);
nor U4917 (N_4917,N_4676,N_4691);
or U4918 (N_4918,N_4638,N_4698);
and U4919 (N_4919,N_4663,N_4618);
xor U4920 (N_4920,N_4783,N_4654);
nand U4921 (N_4921,N_4745,N_4646);
or U4922 (N_4922,N_4757,N_4606);
or U4923 (N_4923,N_4653,N_4728);
or U4924 (N_4924,N_4651,N_4647);
xor U4925 (N_4925,N_4736,N_4646);
or U4926 (N_4926,N_4699,N_4727);
nand U4927 (N_4927,N_4705,N_4610);
or U4928 (N_4928,N_4749,N_4662);
xnor U4929 (N_4929,N_4777,N_4665);
xnor U4930 (N_4930,N_4670,N_4794);
or U4931 (N_4931,N_4617,N_4634);
xor U4932 (N_4932,N_4714,N_4611);
xor U4933 (N_4933,N_4676,N_4614);
nand U4934 (N_4934,N_4791,N_4663);
or U4935 (N_4935,N_4684,N_4794);
or U4936 (N_4936,N_4620,N_4690);
nor U4937 (N_4937,N_4798,N_4677);
nand U4938 (N_4938,N_4751,N_4660);
xnor U4939 (N_4939,N_4745,N_4705);
or U4940 (N_4940,N_4743,N_4788);
nor U4941 (N_4941,N_4622,N_4623);
xnor U4942 (N_4942,N_4685,N_4755);
nor U4943 (N_4943,N_4674,N_4604);
nor U4944 (N_4944,N_4613,N_4725);
xor U4945 (N_4945,N_4694,N_4660);
nor U4946 (N_4946,N_4715,N_4744);
nand U4947 (N_4947,N_4737,N_4610);
or U4948 (N_4948,N_4684,N_4646);
xnor U4949 (N_4949,N_4733,N_4708);
nand U4950 (N_4950,N_4657,N_4674);
nand U4951 (N_4951,N_4630,N_4725);
or U4952 (N_4952,N_4783,N_4622);
or U4953 (N_4953,N_4770,N_4782);
nor U4954 (N_4954,N_4758,N_4724);
or U4955 (N_4955,N_4730,N_4659);
and U4956 (N_4956,N_4778,N_4747);
nand U4957 (N_4957,N_4635,N_4734);
nor U4958 (N_4958,N_4760,N_4730);
xnor U4959 (N_4959,N_4604,N_4680);
and U4960 (N_4960,N_4630,N_4711);
xnor U4961 (N_4961,N_4782,N_4740);
nand U4962 (N_4962,N_4748,N_4659);
xnor U4963 (N_4963,N_4613,N_4664);
xnor U4964 (N_4964,N_4622,N_4724);
xor U4965 (N_4965,N_4704,N_4755);
or U4966 (N_4966,N_4624,N_4681);
or U4967 (N_4967,N_4747,N_4662);
xor U4968 (N_4968,N_4617,N_4740);
and U4969 (N_4969,N_4637,N_4710);
nor U4970 (N_4970,N_4770,N_4662);
or U4971 (N_4971,N_4741,N_4682);
nand U4972 (N_4972,N_4619,N_4654);
nor U4973 (N_4973,N_4752,N_4650);
and U4974 (N_4974,N_4726,N_4714);
nand U4975 (N_4975,N_4776,N_4778);
nand U4976 (N_4976,N_4695,N_4763);
nand U4977 (N_4977,N_4778,N_4696);
and U4978 (N_4978,N_4711,N_4708);
xor U4979 (N_4979,N_4619,N_4611);
nand U4980 (N_4980,N_4786,N_4718);
and U4981 (N_4981,N_4736,N_4643);
and U4982 (N_4982,N_4600,N_4719);
or U4983 (N_4983,N_4712,N_4630);
nor U4984 (N_4984,N_4723,N_4783);
or U4985 (N_4985,N_4787,N_4717);
nor U4986 (N_4986,N_4751,N_4611);
and U4987 (N_4987,N_4656,N_4721);
nor U4988 (N_4988,N_4764,N_4689);
nand U4989 (N_4989,N_4725,N_4676);
nand U4990 (N_4990,N_4607,N_4774);
nor U4991 (N_4991,N_4740,N_4756);
or U4992 (N_4992,N_4764,N_4766);
and U4993 (N_4993,N_4738,N_4790);
nor U4994 (N_4994,N_4785,N_4657);
nor U4995 (N_4995,N_4751,N_4659);
and U4996 (N_4996,N_4624,N_4703);
nor U4997 (N_4997,N_4771,N_4712);
or U4998 (N_4998,N_4660,N_4739);
nand U4999 (N_4999,N_4723,N_4778);
and U5000 (N_5000,N_4954,N_4911);
or U5001 (N_5001,N_4938,N_4965);
nand U5002 (N_5002,N_4835,N_4800);
and U5003 (N_5003,N_4993,N_4940);
or U5004 (N_5004,N_4959,N_4841);
or U5005 (N_5005,N_4801,N_4931);
nor U5006 (N_5006,N_4817,N_4848);
and U5007 (N_5007,N_4810,N_4857);
or U5008 (N_5008,N_4869,N_4888);
or U5009 (N_5009,N_4831,N_4949);
nor U5010 (N_5010,N_4815,N_4821);
nand U5011 (N_5011,N_4834,N_4813);
xor U5012 (N_5012,N_4960,N_4845);
nor U5013 (N_5013,N_4896,N_4832);
or U5014 (N_5014,N_4871,N_4865);
xnor U5015 (N_5015,N_4805,N_4804);
and U5016 (N_5016,N_4880,N_4825);
or U5017 (N_5017,N_4983,N_4967);
nor U5018 (N_5018,N_4926,N_4933);
or U5019 (N_5019,N_4973,N_4890);
or U5020 (N_5020,N_4830,N_4893);
nand U5021 (N_5021,N_4898,N_4945);
nor U5022 (N_5022,N_4878,N_4979);
or U5023 (N_5023,N_4870,N_4908);
or U5024 (N_5024,N_4846,N_4950);
xor U5025 (N_5025,N_4970,N_4854);
xor U5026 (N_5026,N_4808,N_4824);
and U5027 (N_5027,N_4877,N_4910);
nand U5028 (N_5028,N_4930,N_4892);
or U5029 (N_5029,N_4838,N_4944);
and U5030 (N_5030,N_4975,N_4873);
nor U5031 (N_5031,N_4914,N_4939);
nand U5032 (N_5032,N_4929,N_4925);
and U5033 (N_5033,N_4946,N_4943);
xnor U5034 (N_5034,N_4852,N_4936);
nor U5035 (N_5035,N_4992,N_4836);
nand U5036 (N_5036,N_4998,N_4995);
nor U5037 (N_5037,N_4912,N_4903);
nand U5038 (N_5038,N_4863,N_4875);
nand U5039 (N_5039,N_4828,N_4806);
nor U5040 (N_5040,N_4840,N_4897);
xor U5041 (N_5041,N_4809,N_4844);
nand U5042 (N_5042,N_4884,N_4847);
or U5043 (N_5043,N_4972,N_4851);
nor U5044 (N_5044,N_4937,N_4891);
nor U5045 (N_5045,N_4966,N_4924);
nor U5046 (N_5046,N_4905,N_4902);
nor U5047 (N_5047,N_4822,N_4881);
xnor U5048 (N_5048,N_4802,N_4920);
and U5049 (N_5049,N_4961,N_4989);
and U5050 (N_5050,N_4963,N_4853);
or U5051 (N_5051,N_4874,N_4872);
nor U5052 (N_5052,N_4819,N_4866);
xnor U5053 (N_5053,N_4919,N_4957);
nand U5054 (N_5054,N_4867,N_4969);
nand U5055 (N_5055,N_4952,N_4895);
or U5056 (N_5056,N_4827,N_4850);
or U5057 (N_5057,N_4837,N_4971);
xor U5058 (N_5058,N_4807,N_4826);
nor U5059 (N_5059,N_4861,N_4814);
xor U5060 (N_5060,N_4996,N_4981);
or U5061 (N_5061,N_4923,N_4849);
or U5062 (N_5062,N_4916,N_4951);
and U5063 (N_5063,N_4907,N_4956);
nor U5064 (N_5064,N_4859,N_4883);
nor U5065 (N_5065,N_4986,N_4823);
nor U5066 (N_5066,N_4934,N_4894);
and U5067 (N_5067,N_4889,N_4921);
nor U5068 (N_5068,N_4860,N_4990);
nor U5069 (N_5069,N_4999,N_4977);
or U5070 (N_5070,N_4811,N_4928);
xnor U5071 (N_5071,N_4886,N_4917);
nand U5072 (N_5072,N_4829,N_4879);
nor U5073 (N_5073,N_4976,N_4842);
xnor U5074 (N_5074,N_4958,N_4978);
nor U5075 (N_5075,N_4988,N_4913);
xor U5076 (N_5076,N_4868,N_4812);
or U5077 (N_5077,N_4816,N_4955);
nand U5078 (N_5078,N_4904,N_4953);
nor U5079 (N_5079,N_4882,N_4906);
nor U5080 (N_5080,N_4818,N_4974);
xnor U5081 (N_5081,N_4968,N_4987);
nand U5082 (N_5082,N_4901,N_4932);
nor U5083 (N_5083,N_4985,N_4991);
nor U5084 (N_5084,N_4885,N_4856);
or U5085 (N_5085,N_4935,N_4962);
xor U5086 (N_5086,N_4942,N_4864);
or U5087 (N_5087,N_4964,N_4915);
and U5088 (N_5088,N_4909,N_4839);
xor U5089 (N_5089,N_4900,N_4855);
nand U5090 (N_5090,N_4927,N_4997);
nor U5091 (N_5091,N_4899,N_4858);
or U5092 (N_5092,N_4876,N_4862);
xnor U5093 (N_5093,N_4947,N_4994);
nor U5094 (N_5094,N_4948,N_4887);
nor U5095 (N_5095,N_4982,N_4833);
nor U5096 (N_5096,N_4984,N_4803);
or U5097 (N_5097,N_4820,N_4980);
xnor U5098 (N_5098,N_4918,N_4941);
and U5099 (N_5099,N_4922,N_4843);
nand U5100 (N_5100,N_4882,N_4943);
xor U5101 (N_5101,N_4961,N_4972);
and U5102 (N_5102,N_4977,N_4854);
xnor U5103 (N_5103,N_4850,N_4814);
xor U5104 (N_5104,N_4837,N_4968);
xnor U5105 (N_5105,N_4868,N_4929);
nor U5106 (N_5106,N_4945,N_4926);
nor U5107 (N_5107,N_4963,N_4851);
nand U5108 (N_5108,N_4952,N_4989);
or U5109 (N_5109,N_4936,N_4993);
nand U5110 (N_5110,N_4987,N_4919);
nor U5111 (N_5111,N_4951,N_4978);
nor U5112 (N_5112,N_4881,N_4832);
or U5113 (N_5113,N_4914,N_4845);
and U5114 (N_5114,N_4936,N_4847);
xnor U5115 (N_5115,N_4984,N_4892);
nand U5116 (N_5116,N_4874,N_4979);
nor U5117 (N_5117,N_4880,N_4943);
or U5118 (N_5118,N_4999,N_4937);
nor U5119 (N_5119,N_4907,N_4818);
nand U5120 (N_5120,N_4934,N_4983);
nand U5121 (N_5121,N_4972,N_4860);
nand U5122 (N_5122,N_4949,N_4850);
or U5123 (N_5123,N_4844,N_4896);
nand U5124 (N_5124,N_4929,N_4906);
nand U5125 (N_5125,N_4850,N_4877);
xnor U5126 (N_5126,N_4986,N_4899);
nand U5127 (N_5127,N_4934,N_4900);
xor U5128 (N_5128,N_4806,N_4948);
and U5129 (N_5129,N_4896,N_4819);
nand U5130 (N_5130,N_4839,N_4865);
and U5131 (N_5131,N_4972,N_4897);
and U5132 (N_5132,N_4935,N_4950);
nor U5133 (N_5133,N_4951,N_4994);
and U5134 (N_5134,N_4853,N_4852);
or U5135 (N_5135,N_4956,N_4844);
and U5136 (N_5136,N_4875,N_4825);
nand U5137 (N_5137,N_4984,N_4819);
and U5138 (N_5138,N_4820,N_4908);
or U5139 (N_5139,N_4840,N_4875);
nor U5140 (N_5140,N_4937,N_4831);
or U5141 (N_5141,N_4826,N_4891);
and U5142 (N_5142,N_4827,N_4973);
and U5143 (N_5143,N_4813,N_4996);
xor U5144 (N_5144,N_4828,N_4985);
and U5145 (N_5145,N_4844,N_4964);
nand U5146 (N_5146,N_4933,N_4837);
xor U5147 (N_5147,N_4907,N_4920);
nor U5148 (N_5148,N_4955,N_4968);
and U5149 (N_5149,N_4848,N_4918);
and U5150 (N_5150,N_4966,N_4818);
or U5151 (N_5151,N_4926,N_4863);
and U5152 (N_5152,N_4847,N_4839);
nor U5153 (N_5153,N_4949,N_4971);
xnor U5154 (N_5154,N_4941,N_4933);
nand U5155 (N_5155,N_4911,N_4823);
and U5156 (N_5156,N_4945,N_4800);
or U5157 (N_5157,N_4859,N_4945);
xor U5158 (N_5158,N_4940,N_4928);
nand U5159 (N_5159,N_4873,N_4852);
nor U5160 (N_5160,N_4833,N_4850);
xnor U5161 (N_5161,N_4865,N_4894);
xor U5162 (N_5162,N_4993,N_4911);
nand U5163 (N_5163,N_4949,N_4886);
xor U5164 (N_5164,N_4968,N_4847);
nor U5165 (N_5165,N_4892,N_4949);
xor U5166 (N_5166,N_4921,N_4977);
or U5167 (N_5167,N_4955,N_4983);
nand U5168 (N_5168,N_4927,N_4808);
xnor U5169 (N_5169,N_4808,N_4911);
xor U5170 (N_5170,N_4866,N_4935);
nand U5171 (N_5171,N_4945,N_4963);
nand U5172 (N_5172,N_4980,N_4912);
xnor U5173 (N_5173,N_4965,N_4997);
nor U5174 (N_5174,N_4815,N_4924);
nor U5175 (N_5175,N_4873,N_4931);
xor U5176 (N_5176,N_4905,N_4929);
nor U5177 (N_5177,N_4846,N_4825);
xnor U5178 (N_5178,N_4975,N_4844);
or U5179 (N_5179,N_4974,N_4969);
and U5180 (N_5180,N_4842,N_4821);
xnor U5181 (N_5181,N_4982,N_4871);
nor U5182 (N_5182,N_4922,N_4813);
nand U5183 (N_5183,N_4951,N_4983);
and U5184 (N_5184,N_4875,N_4821);
nor U5185 (N_5185,N_4811,N_4951);
or U5186 (N_5186,N_4906,N_4941);
xnor U5187 (N_5187,N_4923,N_4890);
nand U5188 (N_5188,N_4890,N_4850);
or U5189 (N_5189,N_4860,N_4888);
nor U5190 (N_5190,N_4918,N_4876);
and U5191 (N_5191,N_4840,N_4953);
nor U5192 (N_5192,N_4978,N_4864);
and U5193 (N_5193,N_4828,N_4864);
and U5194 (N_5194,N_4978,N_4903);
or U5195 (N_5195,N_4819,N_4933);
nor U5196 (N_5196,N_4818,N_4829);
nor U5197 (N_5197,N_4981,N_4891);
and U5198 (N_5198,N_4830,N_4904);
or U5199 (N_5199,N_4866,N_4851);
or U5200 (N_5200,N_5057,N_5119);
xor U5201 (N_5201,N_5193,N_5049);
or U5202 (N_5202,N_5148,N_5006);
and U5203 (N_5203,N_5018,N_5113);
or U5204 (N_5204,N_5188,N_5104);
nor U5205 (N_5205,N_5091,N_5074);
or U5206 (N_5206,N_5121,N_5122);
and U5207 (N_5207,N_5003,N_5157);
and U5208 (N_5208,N_5128,N_5098);
nand U5209 (N_5209,N_5085,N_5025);
and U5210 (N_5210,N_5096,N_5064);
and U5211 (N_5211,N_5007,N_5095);
nor U5212 (N_5212,N_5165,N_5183);
or U5213 (N_5213,N_5195,N_5029);
nor U5214 (N_5214,N_5196,N_5069);
nor U5215 (N_5215,N_5154,N_5024);
nand U5216 (N_5216,N_5130,N_5134);
nor U5217 (N_5217,N_5033,N_5194);
or U5218 (N_5218,N_5042,N_5050);
nand U5219 (N_5219,N_5010,N_5186);
xnor U5220 (N_5220,N_5117,N_5079);
nor U5221 (N_5221,N_5144,N_5060);
nand U5222 (N_5222,N_5184,N_5116);
nor U5223 (N_5223,N_5170,N_5012);
nand U5224 (N_5224,N_5112,N_5129);
or U5225 (N_5225,N_5051,N_5123);
xor U5226 (N_5226,N_5089,N_5125);
xor U5227 (N_5227,N_5043,N_5027);
xnor U5228 (N_5228,N_5030,N_5011);
nand U5229 (N_5229,N_5002,N_5107);
xnor U5230 (N_5230,N_5093,N_5164);
or U5231 (N_5231,N_5044,N_5178);
nand U5232 (N_5232,N_5000,N_5180);
or U5233 (N_5233,N_5199,N_5082);
nand U5234 (N_5234,N_5040,N_5108);
xor U5235 (N_5235,N_5181,N_5143);
nand U5236 (N_5236,N_5090,N_5167);
xor U5237 (N_5237,N_5155,N_5073);
nor U5238 (N_5238,N_5031,N_5022);
nor U5239 (N_5239,N_5126,N_5072);
and U5240 (N_5240,N_5026,N_5156);
and U5241 (N_5241,N_5146,N_5099);
nand U5242 (N_5242,N_5190,N_5092);
and U5243 (N_5243,N_5133,N_5150);
xor U5244 (N_5244,N_5061,N_5087);
and U5245 (N_5245,N_5136,N_5004);
or U5246 (N_5246,N_5048,N_5198);
nor U5247 (N_5247,N_5109,N_5086);
nor U5248 (N_5248,N_5177,N_5052);
xor U5249 (N_5249,N_5127,N_5078);
xor U5250 (N_5250,N_5065,N_5021);
or U5251 (N_5251,N_5151,N_5187);
nor U5252 (N_5252,N_5118,N_5075);
or U5253 (N_5253,N_5034,N_5139);
nand U5254 (N_5254,N_5160,N_5088);
xor U5255 (N_5255,N_5019,N_5163);
and U5256 (N_5256,N_5077,N_5142);
nor U5257 (N_5257,N_5192,N_5162);
nor U5258 (N_5258,N_5032,N_5041);
nand U5259 (N_5259,N_5056,N_5101);
nor U5260 (N_5260,N_5046,N_5138);
xnor U5261 (N_5261,N_5014,N_5054);
nor U5262 (N_5262,N_5141,N_5047);
nand U5263 (N_5263,N_5053,N_5103);
nand U5264 (N_5264,N_5110,N_5037);
or U5265 (N_5265,N_5100,N_5023);
and U5266 (N_5266,N_5102,N_5070);
nor U5267 (N_5267,N_5179,N_5058);
or U5268 (N_5268,N_5115,N_5166);
and U5269 (N_5269,N_5016,N_5076);
and U5270 (N_5270,N_5038,N_5071);
and U5271 (N_5271,N_5137,N_5045);
nand U5272 (N_5272,N_5197,N_5124);
nand U5273 (N_5273,N_5158,N_5036);
nand U5274 (N_5274,N_5013,N_5120);
nor U5275 (N_5275,N_5055,N_5017);
or U5276 (N_5276,N_5001,N_5084);
or U5277 (N_5277,N_5111,N_5094);
or U5278 (N_5278,N_5097,N_5171);
xnor U5279 (N_5279,N_5009,N_5149);
or U5280 (N_5280,N_5174,N_5059);
or U5281 (N_5281,N_5114,N_5080);
nand U5282 (N_5282,N_5189,N_5182);
or U5283 (N_5283,N_5066,N_5185);
and U5284 (N_5284,N_5140,N_5039);
and U5285 (N_5285,N_5005,N_5176);
nand U5286 (N_5286,N_5105,N_5063);
and U5287 (N_5287,N_5131,N_5020);
nand U5288 (N_5288,N_5168,N_5062);
nor U5289 (N_5289,N_5135,N_5083);
nand U5290 (N_5290,N_5145,N_5067);
or U5291 (N_5291,N_5172,N_5132);
nor U5292 (N_5292,N_5147,N_5153);
and U5293 (N_5293,N_5169,N_5008);
or U5294 (N_5294,N_5173,N_5175);
or U5295 (N_5295,N_5068,N_5191);
nand U5296 (N_5296,N_5161,N_5152);
and U5297 (N_5297,N_5015,N_5028);
nor U5298 (N_5298,N_5106,N_5035);
nor U5299 (N_5299,N_5159,N_5081);
xor U5300 (N_5300,N_5040,N_5009);
nor U5301 (N_5301,N_5060,N_5066);
xnor U5302 (N_5302,N_5039,N_5059);
or U5303 (N_5303,N_5099,N_5115);
nor U5304 (N_5304,N_5029,N_5153);
xnor U5305 (N_5305,N_5180,N_5147);
nor U5306 (N_5306,N_5166,N_5170);
and U5307 (N_5307,N_5099,N_5043);
nand U5308 (N_5308,N_5050,N_5169);
nand U5309 (N_5309,N_5006,N_5143);
xor U5310 (N_5310,N_5096,N_5058);
and U5311 (N_5311,N_5004,N_5142);
nor U5312 (N_5312,N_5083,N_5110);
nand U5313 (N_5313,N_5165,N_5185);
xnor U5314 (N_5314,N_5107,N_5183);
nand U5315 (N_5315,N_5041,N_5084);
or U5316 (N_5316,N_5005,N_5009);
or U5317 (N_5317,N_5177,N_5049);
nor U5318 (N_5318,N_5060,N_5149);
nand U5319 (N_5319,N_5154,N_5092);
nand U5320 (N_5320,N_5164,N_5038);
or U5321 (N_5321,N_5047,N_5087);
and U5322 (N_5322,N_5003,N_5151);
nand U5323 (N_5323,N_5155,N_5074);
or U5324 (N_5324,N_5075,N_5186);
or U5325 (N_5325,N_5094,N_5179);
nor U5326 (N_5326,N_5181,N_5109);
xnor U5327 (N_5327,N_5094,N_5032);
xnor U5328 (N_5328,N_5154,N_5164);
and U5329 (N_5329,N_5091,N_5101);
nand U5330 (N_5330,N_5107,N_5185);
xor U5331 (N_5331,N_5096,N_5007);
and U5332 (N_5332,N_5056,N_5117);
or U5333 (N_5333,N_5111,N_5011);
nand U5334 (N_5334,N_5145,N_5037);
nor U5335 (N_5335,N_5162,N_5035);
nand U5336 (N_5336,N_5147,N_5181);
xnor U5337 (N_5337,N_5124,N_5091);
or U5338 (N_5338,N_5046,N_5128);
nand U5339 (N_5339,N_5108,N_5073);
nand U5340 (N_5340,N_5094,N_5190);
xor U5341 (N_5341,N_5008,N_5139);
nand U5342 (N_5342,N_5042,N_5165);
nand U5343 (N_5343,N_5134,N_5089);
xor U5344 (N_5344,N_5133,N_5140);
or U5345 (N_5345,N_5146,N_5105);
nand U5346 (N_5346,N_5036,N_5049);
nor U5347 (N_5347,N_5064,N_5020);
nor U5348 (N_5348,N_5114,N_5006);
and U5349 (N_5349,N_5061,N_5083);
and U5350 (N_5350,N_5103,N_5182);
xor U5351 (N_5351,N_5108,N_5121);
or U5352 (N_5352,N_5161,N_5110);
nor U5353 (N_5353,N_5180,N_5054);
nand U5354 (N_5354,N_5148,N_5017);
and U5355 (N_5355,N_5048,N_5097);
xnor U5356 (N_5356,N_5009,N_5100);
or U5357 (N_5357,N_5053,N_5041);
nand U5358 (N_5358,N_5185,N_5173);
and U5359 (N_5359,N_5181,N_5018);
or U5360 (N_5360,N_5082,N_5053);
xnor U5361 (N_5361,N_5152,N_5009);
nor U5362 (N_5362,N_5091,N_5108);
nand U5363 (N_5363,N_5025,N_5164);
or U5364 (N_5364,N_5037,N_5199);
xnor U5365 (N_5365,N_5015,N_5168);
nand U5366 (N_5366,N_5045,N_5059);
nand U5367 (N_5367,N_5181,N_5001);
nor U5368 (N_5368,N_5121,N_5020);
and U5369 (N_5369,N_5051,N_5017);
xnor U5370 (N_5370,N_5122,N_5086);
and U5371 (N_5371,N_5082,N_5097);
and U5372 (N_5372,N_5016,N_5137);
nand U5373 (N_5373,N_5109,N_5056);
xor U5374 (N_5374,N_5067,N_5175);
nor U5375 (N_5375,N_5174,N_5194);
or U5376 (N_5376,N_5031,N_5162);
and U5377 (N_5377,N_5106,N_5038);
or U5378 (N_5378,N_5160,N_5030);
nand U5379 (N_5379,N_5028,N_5018);
xor U5380 (N_5380,N_5105,N_5143);
or U5381 (N_5381,N_5024,N_5072);
nand U5382 (N_5382,N_5116,N_5109);
nor U5383 (N_5383,N_5102,N_5095);
xnor U5384 (N_5384,N_5194,N_5188);
or U5385 (N_5385,N_5178,N_5020);
nor U5386 (N_5386,N_5083,N_5190);
nor U5387 (N_5387,N_5027,N_5165);
xnor U5388 (N_5388,N_5146,N_5170);
nor U5389 (N_5389,N_5136,N_5129);
nand U5390 (N_5390,N_5188,N_5128);
or U5391 (N_5391,N_5042,N_5178);
nor U5392 (N_5392,N_5012,N_5053);
and U5393 (N_5393,N_5087,N_5103);
and U5394 (N_5394,N_5193,N_5042);
nand U5395 (N_5395,N_5165,N_5003);
xnor U5396 (N_5396,N_5177,N_5061);
nand U5397 (N_5397,N_5098,N_5080);
or U5398 (N_5398,N_5193,N_5198);
nor U5399 (N_5399,N_5166,N_5142);
xnor U5400 (N_5400,N_5380,N_5375);
nor U5401 (N_5401,N_5287,N_5290);
xor U5402 (N_5402,N_5376,N_5389);
or U5403 (N_5403,N_5286,N_5243);
xor U5404 (N_5404,N_5354,N_5264);
or U5405 (N_5405,N_5236,N_5350);
nor U5406 (N_5406,N_5232,N_5211);
and U5407 (N_5407,N_5285,N_5229);
xnor U5408 (N_5408,N_5320,N_5218);
nand U5409 (N_5409,N_5328,N_5395);
nand U5410 (N_5410,N_5318,N_5242);
nand U5411 (N_5411,N_5291,N_5215);
nor U5412 (N_5412,N_5269,N_5208);
nand U5413 (N_5413,N_5321,N_5273);
or U5414 (N_5414,N_5388,N_5222);
or U5415 (N_5415,N_5301,N_5268);
xnor U5416 (N_5416,N_5345,N_5314);
nand U5417 (N_5417,N_5246,N_5326);
xnor U5418 (N_5418,N_5295,N_5270);
nand U5419 (N_5419,N_5245,N_5393);
or U5420 (N_5420,N_5378,N_5343);
nor U5421 (N_5421,N_5374,N_5384);
or U5422 (N_5422,N_5260,N_5340);
or U5423 (N_5423,N_5262,N_5338);
nor U5424 (N_5424,N_5255,N_5294);
nor U5425 (N_5425,N_5308,N_5348);
or U5426 (N_5426,N_5382,N_5250);
or U5427 (N_5427,N_5339,N_5271);
nand U5428 (N_5428,N_5240,N_5239);
or U5429 (N_5429,N_5281,N_5275);
nor U5430 (N_5430,N_5233,N_5399);
xnor U5431 (N_5431,N_5228,N_5247);
and U5432 (N_5432,N_5324,N_5235);
nor U5433 (N_5433,N_5204,N_5333);
and U5434 (N_5434,N_5357,N_5227);
and U5435 (N_5435,N_5279,N_5372);
and U5436 (N_5436,N_5307,N_5312);
and U5437 (N_5437,N_5244,N_5309);
nand U5438 (N_5438,N_5306,N_5266);
nor U5439 (N_5439,N_5216,N_5254);
or U5440 (N_5440,N_5369,N_5371);
and U5441 (N_5441,N_5353,N_5203);
or U5442 (N_5442,N_5362,N_5379);
or U5443 (N_5443,N_5230,N_5282);
or U5444 (N_5444,N_5366,N_5315);
xor U5445 (N_5445,N_5323,N_5258);
and U5446 (N_5446,N_5319,N_5283);
or U5447 (N_5447,N_5390,N_5241);
and U5448 (N_5448,N_5207,N_5322);
xnor U5449 (N_5449,N_5261,N_5313);
nor U5450 (N_5450,N_5212,N_5223);
nand U5451 (N_5451,N_5302,N_5289);
and U5452 (N_5452,N_5359,N_5332);
and U5453 (N_5453,N_5385,N_5298);
nand U5454 (N_5454,N_5327,N_5202);
nor U5455 (N_5455,N_5391,N_5231);
nand U5456 (N_5456,N_5311,N_5297);
nor U5457 (N_5457,N_5252,N_5325);
xor U5458 (N_5458,N_5304,N_5381);
or U5459 (N_5459,N_5394,N_5364);
nor U5460 (N_5460,N_5387,N_5392);
nand U5461 (N_5461,N_5317,N_5248);
and U5462 (N_5462,N_5249,N_5300);
xor U5463 (N_5463,N_5288,N_5272);
nor U5464 (N_5464,N_5370,N_5274);
xor U5465 (N_5465,N_5259,N_5373);
xor U5466 (N_5466,N_5201,N_5200);
nand U5467 (N_5467,N_5347,N_5299);
xor U5468 (N_5468,N_5293,N_5377);
or U5469 (N_5469,N_5267,N_5253);
or U5470 (N_5470,N_5349,N_5226);
or U5471 (N_5471,N_5292,N_5346);
nor U5472 (N_5472,N_5303,N_5276);
and U5473 (N_5473,N_5217,N_5237);
and U5474 (N_5474,N_5310,N_5234);
nand U5475 (N_5475,N_5221,N_5238);
nand U5476 (N_5476,N_5219,N_5342);
and U5477 (N_5477,N_5257,N_5210);
or U5478 (N_5478,N_5365,N_5398);
nand U5479 (N_5479,N_5251,N_5209);
or U5480 (N_5480,N_5205,N_5344);
nor U5481 (N_5481,N_5305,N_5337);
or U5482 (N_5482,N_5225,N_5278);
xnor U5483 (N_5483,N_5280,N_5341);
or U5484 (N_5484,N_5284,N_5296);
or U5485 (N_5485,N_5386,N_5265);
nand U5486 (N_5486,N_5397,N_5363);
and U5487 (N_5487,N_5368,N_5383);
xor U5488 (N_5488,N_5330,N_5361);
nand U5489 (N_5489,N_5206,N_5396);
xor U5490 (N_5490,N_5224,N_5356);
nand U5491 (N_5491,N_5331,N_5316);
nor U5492 (N_5492,N_5336,N_5334);
and U5493 (N_5493,N_5367,N_5355);
or U5494 (N_5494,N_5351,N_5220);
and U5495 (N_5495,N_5360,N_5263);
nand U5496 (N_5496,N_5358,N_5277);
or U5497 (N_5497,N_5352,N_5256);
nand U5498 (N_5498,N_5329,N_5213);
xnor U5499 (N_5499,N_5214,N_5335);
or U5500 (N_5500,N_5217,N_5398);
nor U5501 (N_5501,N_5346,N_5207);
nand U5502 (N_5502,N_5350,N_5228);
nand U5503 (N_5503,N_5284,N_5241);
nand U5504 (N_5504,N_5248,N_5345);
nor U5505 (N_5505,N_5249,N_5232);
nor U5506 (N_5506,N_5364,N_5348);
or U5507 (N_5507,N_5351,N_5383);
nor U5508 (N_5508,N_5346,N_5389);
nor U5509 (N_5509,N_5396,N_5366);
or U5510 (N_5510,N_5314,N_5245);
and U5511 (N_5511,N_5235,N_5387);
or U5512 (N_5512,N_5343,N_5364);
nor U5513 (N_5513,N_5277,N_5292);
nor U5514 (N_5514,N_5326,N_5397);
nand U5515 (N_5515,N_5338,N_5255);
or U5516 (N_5516,N_5371,N_5300);
or U5517 (N_5517,N_5215,N_5225);
nor U5518 (N_5518,N_5282,N_5336);
and U5519 (N_5519,N_5241,N_5347);
xor U5520 (N_5520,N_5398,N_5375);
nand U5521 (N_5521,N_5352,N_5264);
and U5522 (N_5522,N_5357,N_5350);
xor U5523 (N_5523,N_5382,N_5278);
nand U5524 (N_5524,N_5212,N_5372);
nor U5525 (N_5525,N_5266,N_5309);
or U5526 (N_5526,N_5232,N_5304);
nand U5527 (N_5527,N_5263,N_5340);
nand U5528 (N_5528,N_5296,N_5298);
xor U5529 (N_5529,N_5250,N_5295);
nor U5530 (N_5530,N_5273,N_5225);
nor U5531 (N_5531,N_5288,N_5229);
and U5532 (N_5532,N_5213,N_5299);
and U5533 (N_5533,N_5271,N_5248);
nor U5534 (N_5534,N_5330,N_5367);
nand U5535 (N_5535,N_5211,N_5334);
or U5536 (N_5536,N_5314,N_5366);
and U5537 (N_5537,N_5325,N_5282);
or U5538 (N_5538,N_5235,N_5261);
nor U5539 (N_5539,N_5252,N_5251);
nand U5540 (N_5540,N_5331,N_5213);
nand U5541 (N_5541,N_5399,N_5262);
or U5542 (N_5542,N_5205,N_5211);
nand U5543 (N_5543,N_5296,N_5307);
and U5544 (N_5544,N_5386,N_5330);
nand U5545 (N_5545,N_5322,N_5316);
xor U5546 (N_5546,N_5318,N_5321);
nor U5547 (N_5547,N_5391,N_5359);
nand U5548 (N_5548,N_5354,N_5387);
nor U5549 (N_5549,N_5224,N_5215);
and U5550 (N_5550,N_5344,N_5245);
xnor U5551 (N_5551,N_5393,N_5216);
nand U5552 (N_5552,N_5214,N_5260);
and U5553 (N_5553,N_5333,N_5305);
or U5554 (N_5554,N_5303,N_5310);
and U5555 (N_5555,N_5208,N_5234);
nor U5556 (N_5556,N_5366,N_5278);
nand U5557 (N_5557,N_5388,N_5311);
xor U5558 (N_5558,N_5363,N_5336);
xor U5559 (N_5559,N_5290,N_5362);
nand U5560 (N_5560,N_5363,N_5222);
nand U5561 (N_5561,N_5345,N_5337);
or U5562 (N_5562,N_5283,N_5396);
xor U5563 (N_5563,N_5267,N_5254);
xor U5564 (N_5564,N_5390,N_5267);
nor U5565 (N_5565,N_5274,N_5396);
or U5566 (N_5566,N_5322,N_5388);
or U5567 (N_5567,N_5322,N_5200);
or U5568 (N_5568,N_5216,N_5236);
or U5569 (N_5569,N_5228,N_5315);
and U5570 (N_5570,N_5224,N_5335);
nor U5571 (N_5571,N_5369,N_5394);
xnor U5572 (N_5572,N_5245,N_5280);
and U5573 (N_5573,N_5309,N_5360);
nand U5574 (N_5574,N_5371,N_5238);
nand U5575 (N_5575,N_5353,N_5372);
and U5576 (N_5576,N_5383,N_5220);
nand U5577 (N_5577,N_5217,N_5301);
nor U5578 (N_5578,N_5316,N_5345);
and U5579 (N_5579,N_5257,N_5305);
and U5580 (N_5580,N_5248,N_5213);
and U5581 (N_5581,N_5319,N_5372);
nor U5582 (N_5582,N_5382,N_5291);
xnor U5583 (N_5583,N_5242,N_5223);
or U5584 (N_5584,N_5396,N_5346);
xnor U5585 (N_5585,N_5309,N_5241);
and U5586 (N_5586,N_5398,N_5333);
nand U5587 (N_5587,N_5320,N_5301);
nand U5588 (N_5588,N_5378,N_5290);
nand U5589 (N_5589,N_5222,N_5281);
nor U5590 (N_5590,N_5237,N_5313);
xnor U5591 (N_5591,N_5207,N_5224);
nor U5592 (N_5592,N_5233,N_5257);
nand U5593 (N_5593,N_5320,N_5298);
xor U5594 (N_5594,N_5254,N_5228);
nand U5595 (N_5595,N_5265,N_5220);
and U5596 (N_5596,N_5202,N_5277);
or U5597 (N_5597,N_5245,N_5281);
xor U5598 (N_5598,N_5343,N_5213);
nand U5599 (N_5599,N_5230,N_5380);
nor U5600 (N_5600,N_5435,N_5597);
xor U5601 (N_5601,N_5450,N_5537);
nand U5602 (N_5602,N_5506,N_5404);
or U5603 (N_5603,N_5587,N_5425);
or U5604 (N_5604,N_5589,N_5459);
xnor U5605 (N_5605,N_5498,N_5484);
or U5606 (N_5606,N_5451,N_5517);
xnor U5607 (N_5607,N_5493,N_5562);
xor U5608 (N_5608,N_5447,N_5488);
nor U5609 (N_5609,N_5532,N_5586);
xnor U5610 (N_5610,N_5553,N_5476);
and U5611 (N_5611,N_5556,N_5565);
xor U5612 (N_5612,N_5531,N_5555);
and U5613 (N_5613,N_5462,N_5591);
nor U5614 (N_5614,N_5489,N_5465);
nor U5615 (N_5615,N_5473,N_5432);
nor U5616 (N_5616,N_5558,N_5544);
nor U5617 (N_5617,N_5491,N_5442);
nor U5618 (N_5618,N_5509,N_5570);
and U5619 (N_5619,N_5411,N_5436);
and U5620 (N_5620,N_5480,N_5594);
nand U5621 (N_5621,N_5566,N_5449);
nand U5622 (N_5622,N_5464,N_5426);
xnor U5623 (N_5623,N_5495,N_5487);
xor U5624 (N_5624,N_5401,N_5581);
and U5625 (N_5625,N_5576,N_5513);
and U5626 (N_5626,N_5413,N_5481);
xnor U5627 (N_5627,N_5472,N_5564);
xnor U5628 (N_5628,N_5524,N_5504);
nand U5629 (N_5629,N_5547,N_5560);
or U5630 (N_5630,N_5535,N_5529);
nand U5631 (N_5631,N_5474,N_5567);
xor U5632 (N_5632,N_5595,N_5554);
or U5633 (N_5633,N_5423,N_5519);
xor U5634 (N_5634,N_5541,N_5503);
and U5635 (N_5635,N_5416,N_5407);
and U5636 (N_5636,N_5499,N_5482);
nand U5637 (N_5637,N_5578,N_5420);
and U5638 (N_5638,N_5526,N_5461);
nand U5639 (N_5639,N_5458,N_5417);
nor U5640 (N_5640,N_5477,N_5421);
nor U5641 (N_5641,N_5453,N_5582);
xnor U5642 (N_5642,N_5405,N_5580);
nand U5643 (N_5643,N_5414,N_5505);
nand U5644 (N_5644,N_5551,N_5409);
nand U5645 (N_5645,N_5585,N_5475);
or U5646 (N_5646,N_5550,N_5527);
nand U5647 (N_5647,N_5559,N_5511);
and U5648 (N_5648,N_5466,N_5533);
nand U5649 (N_5649,N_5463,N_5599);
nand U5650 (N_5650,N_5557,N_5437);
or U5651 (N_5651,N_5440,N_5485);
and U5652 (N_5652,N_5561,N_5446);
nor U5653 (N_5653,N_5479,N_5523);
xor U5654 (N_5654,N_5443,N_5593);
nand U5655 (N_5655,N_5444,N_5448);
nor U5656 (N_5656,N_5402,N_5584);
nand U5657 (N_5657,N_5500,N_5486);
and U5658 (N_5658,N_5483,N_5540);
and U5659 (N_5659,N_5467,N_5563);
xor U5660 (N_5660,N_5536,N_5548);
and U5661 (N_5661,N_5471,N_5521);
and U5662 (N_5662,N_5433,N_5431);
xor U5663 (N_5663,N_5510,N_5516);
or U5664 (N_5664,N_5574,N_5590);
nor U5665 (N_5665,N_5592,N_5469);
nor U5666 (N_5666,N_5460,N_5429);
and U5667 (N_5667,N_5434,N_5525);
nor U5668 (N_5668,N_5512,N_5456);
nor U5669 (N_5669,N_5497,N_5400);
nand U5670 (N_5670,N_5445,N_5549);
or U5671 (N_5671,N_5427,N_5573);
or U5672 (N_5672,N_5412,N_5494);
and U5673 (N_5673,N_5569,N_5568);
or U5674 (N_5674,N_5542,N_5518);
or U5675 (N_5675,N_5408,N_5530);
or U5676 (N_5676,N_5545,N_5428);
xnor U5677 (N_5677,N_5514,N_5468);
and U5678 (N_5678,N_5454,N_5539);
and U5679 (N_5679,N_5528,N_5577);
nor U5680 (N_5680,N_5522,N_5579);
or U5681 (N_5681,N_5430,N_5515);
nor U5682 (N_5682,N_5410,N_5415);
or U5683 (N_5683,N_5508,N_5438);
xnor U5684 (N_5684,N_5507,N_5583);
xor U5685 (N_5685,N_5470,N_5441);
xnor U5686 (N_5686,N_5552,N_5543);
nor U5687 (N_5687,N_5457,N_5439);
or U5688 (N_5688,N_5452,N_5588);
or U5689 (N_5689,N_5403,N_5422);
nor U5690 (N_5690,N_5546,N_5598);
nor U5691 (N_5691,N_5520,N_5418);
nor U5692 (N_5692,N_5534,N_5596);
or U5693 (N_5693,N_5455,N_5478);
nor U5694 (N_5694,N_5575,N_5502);
nand U5695 (N_5695,N_5496,N_5492);
and U5696 (N_5696,N_5572,N_5406);
nor U5697 (N_5697,N_5538,N_5424);
or U5698 (N_5698,N_5419,N_5490);
or U5699 (N_5699,N_5501,N_5571);
nor U5700 (N_5700,N_5527,N_5503);
or U5701 (N_5701,N_5416,N_5505);
and U5702 (N_5702,N_5573,N_5533);
xor U5703 (N_5703,N_5434,N_5530);
nor U5704 (N_5704,N_5588,N_5454);
and U5705 (N_5705,N_5482,N_5512);
and U5706 (N_5706,N_5538,N_5498);
or U5707 (N_5707,N_5481,N_5455);
or U5708 (N_5708,N_5476,N_5408);
nand U5709 (N_5709,N_5424,N_5500);
or U5710 (N_5710,N_5437,N_5538);
nor U5711 (N_5711,N_5479,N_5435);
xnor U5712 (N_5712,N_5473,N_5483);
or U5713 (N_5713,N_5549,N_5468);
xor U5714 (N_5714,N_5510,N_5430);
and U5715 (N_5715,N_5443,N_5414);
or U5716 (N_5716,N_5489,N_5564);
nand U5717 (N_5717,N_5414,N_5598);
or U5718 (N_5718,N_5498,N_5499);
and U5719 (N_5719,N_5525,N_5549);
xor U5720 (N_5720,N_5470,N_5524);
xnor U5721 (N_5721,N_5439,N_5528);
xnor U5722 (N_5722,N_5488,N_5419);
xnor U5723 (N_5723,N_5526,N_5492);
nor U5724 (N_5724,N_5577,N_5544);
xor U5725 (N_5725,N_5417,N_5470);
or U5726 (N_5726,N_5433,N_5425);
and U5727 (N_5727,N_5589,N_5425);
or U5728 (N_5728,N_5497,N_5597);
xnor U5729 (N_5729,N_5429,N_5401);
xnor U5730 (N_5730,N_5441,N_5535);
nand U5731 (N_5731,N_5450,N_5455);
nor U5732 (N_5732,N_5431,N_5535);
nor U5733 (N_5733,N_5576,N_5452);
xor U5734 (N_5734,N_5540,N_5529);
and U5735 (N_5735,N_5430,N_5422);
nor U5736 (N_5736,N_5404,N_5468);
or U5737 (N_5737,N_5503,N_5484);
and U5738 (N_5738,N_5501,N_5561);
nor U5739 (N_5739,N_5543,N_5473);
or U5740 (N_5740,N_5504,N_5519);
or U5741 (N_5741,N_5426,N_5588);
or U5742 (N_5742,N_5436,N_5517);
nor U5743 (N_5743,N_5469,N_5565);
xnor U5744 (N_5744,N_5476,N_5539);
nand U5745 (N_5745,N_5566,N_5412);
and U5746 (N_5746,N_5459,N_5533);
and U5747 (N_5747,N_5404,N_5416);
nor U5748 (N_5748,N_5558,N_5473);
and U5749 (N_5749,N_5405,N_5436);
nand U5750 (N_5750,N_5484,N_5432);
xor U5751 (N_5751,N_5498,N_5434);
or U5752 (N_5752,N_5573,N_5489);
xor U5753 (N_5753,N_5420,N_5424);
and U5754 (N_5754,N_5557,N_5596);
nand U5755 (N_5755,N_5482,N_5549);
nand U5756 (N_5756,N_5506,N_5588);
nor U5757 (N_5757,N_5442,N_5451);
nand U5758 (N_5758,N_5493,N_5430);
or U5759 (N_5759,N_5472,N_5484);
or U5760 (N_5760,N_5581,N_5418);
or U5761 (N_5761,N_5506,N_5452);
nand U5762 (N_5762,N_5407,N_5448);
and U5763 (N_5763,N_5452,N_5404);
nor U5764 (N_5764,N_5485,N_5400);
nor U5765 (N_5765,N_5449,N_5580);
xnor U5766 (N_5766,N_5506,N_5501);
nand U5767 (N_5767,N_5562,N_5541);
xnor U5768 (N_5768,N_5563,N_5572);
and U5769 (N_5769,N_5581,N_5544);
or U5770 (N_5770,N_5430,N_5562);
or U5771 (N_5771,N_5478,N_5522);
xor U5772 (N_5772,N_5467,N_5436);
or U5773 (N_5773,N_5545,N_5593);
and U5774 (N_5774,N_5588,N_5440);
or U5775 (N_5775,N_5438,N_5556);
nor U5776 (N_5776,N_5494,N_5593);
nor U5777 (N_5777,N_5547,N_5448);
nor U5778 (N_5778,N_5436,N_5569);
nand U5779 (N_5779,N_5572,N_5584);
nand U5780 (N_5780,N_5494,N_5517);
xnor U5781 (N_5781,N_5583,N_5526);
nor U5782 (N_5782,N_5418,N_5590);
nor U5783 (N_5783,N_5573,N_5400);
nor U5784 (N_5784,N_5437,N_5591);
nor U5785 (N_5785,N_5536,N_5539);
nand U5786 (N_5786,N_5435,N_5594);
and U5787 (N_5787,N_5488,N_5497);
and U5788 (N_5788,N_5512,N_5416);
or U5789 (N_5789,N_5490,N_5594);
nand U5790 (N_5790,N_5496,N_5431);
or U5791 (N_5791,N_5516,N_5564);
or U5792 (N_5792,N_5598,N_5513);
xnor U5793 (N_5793,N_5568,N_5591);
nor U5794 (N_5794,N_5413,N_5514);
nor U5795 (N_5795,N_5455,N_5440);
xnor U5796 (N_5796,N_5575,N_5516);
and U5797 (N_5797,N_5410,N_5434);
or U5798 (N_5798,N_5552,N_5432);
nand U5799 (N_5799,N_5556,N_5597);
and U5800 (N_5800,N_5702,N_5726);
xnor U5801 (N_5801,N_5656,N_5774);
and U5802 (N_5802,N_5618,N_5758);
or U5803 (N_5803,N_5783,N_5780);
xnor U5804 (N_5804,N_5744,N_5708);
or U5805 (N_5805,N_5766,N_5692);
or U5806 (N_5806,N_5749,N_5799);
nor U5807 (N_5807,N_5771,N_5621);
and U5808 (N_5808,N_5717,N_5678);
or U5809 (N_5809,N_5677,N_5777);
nand U5810 (N_5810,N_5691,N_5690);
nand U5811 (N_5811,N_5666,N_5721);
or U5812 (N_5812,N_5657,N_5668);
or U5813 (N_5813,N_5623,N_5785);
and U5814 (N_5814,N_5698,N_5757);
or U5815 (N_5815,N_5626,N_5792);
and U5816 (N_5816,N_5743,N_5671);
nor U5817 (N_5817,N_5738,N_5741);
and U5818 (N_5818,N_5659,N_5700);
and U5819 (N_5819,N_5636,N_5706);
nor U5820 (N_5820,N_5759,N_5781);
nand U5821 (N_5821,N_5739,N_5663);
xor U5822 (N_5822,N_5712,N_5673);
nor U5823 (N_5823,N_5797,N_5796);
and U5824 (N_5824,N_5633,N_5609);
nor U5825 (N_5825,N_5630,N_5687);
nor U5826 (N_5826,N_5790,N_5769);
nand U5827 (N_5827,N_5763,N_5787);
or U5828 (N_5828,N_5637,N_5729);
nand U5829 (N_5829,N_5788,N_5751);
and U5830 (N_5830,N_5746,N_5620);
nand U5831 (N_5831,N_5639,N_5709);
and U5832 (N_5832,N_5635,N_5755);
xnor U5833 (N_5833,N_5638,N_5754);
or U5834 (N_5834,N_5778,N_5683);
nor U5835 (N_5835,N_5697,N_5694);
xnor U5836 (N_5836,N_5646,N_5719);
nor U5837 (N_5837,N_5629,N_5725);
nor U5838 (N_5838,N_5670,N_5756);
nor U5839 (N_5839,N_5684,N_5776);
or U5840 (N_5840,N_5614,N_5718);
or U5841 (N_5841,N_5791,N_5723);
or U5842 (N_5842,N_5710,N_5612);
xnor U5843 (N_5843,N_5768,N_5649);
nor U5844 (N_5844,N_5602,N_5604);
nand U5845 (N_5845,N_5640,N_5658);
and U5846 (N_5846,N_5617,N_5679);
and U5847 (N_5847,N_5753,N_5632);
or U5848 (N_5848,N_5793,N_5610);
nand U5849 (N_5849,N_5681,N_5760);
nand U5850 (N_5850,N_5740,N_5795);
xnor U5851 (N_5851,N_5724,N_5752);
nand U5852 (N_5852,N_5607,N_5601);
or U5853 (N_5853,N_5653,N_5733);
and U5854 (N_5854,N_5643,N_5619);
or U5855 (N_5855,N_5603,N_5714);
or U5856 (N_5856,N_5655,N_5622);
or U5857 (N_5857,N_5789,N_5644);
nand U5858 (N_5858,N_5716,N_5693);
nor U5859 (N_5859,N_5695,N_5642);
nand U5860 (N_5860,N_5705,N_5625);
or U5861 (N_5861,N_5711,N_5775);
and U5862 (N_5862,N_5742,N_5722);
or U5863 (N_5863,N_5680,N_5765);
nand U5864 (N_5864,N_5664,N_5786);
xor U5865 (N_5865,N_5682,N_5665);
or U5866 (N_5866,N_5732,N_5675);
and U5867 (N_5867,N_5660,N_5767);
and U5868 (N_5868,N_5779,N_5696);
or U5869 (N_5869,N_5662,N_5608);
nor U5870 (N_5870,N_5699,N_5600);
nor U5871 (N_5871,N_5661,N_5667);
and U5872 (N_5872,N_5772,N_5615);
xor U5873 (N_5873,N_5731,N_5648);
or U5874 (N_5874,N_5707,N_5761);
nor U5875 (N_5875,N_5686,N_5727);
or U5876 (N_5876,N_5764,N_5688);
or U5877 (N_5877,N_5782,N_5650);
nand U5878 (N_5878,N_5773,N_5701);
or U5879 (N_5879,N_5703,N_5627);
xnor U5880 (N_5880,N_5794,N_5720);
and U5881 (N_5881,N_5611,N_5641);
nor U5882 (N_5882,N_5605,N_5713);
xor U5883 (N_5883,N_5669,N_5736);
nor U5884 (N_5884,N_5735,N_5730);
xor U5885 (N_5885,N_5798,N_5770);
xor U5886 (N_5886,N_5628,N_5651);
nor U5887 (N_5887,N_5676,N_5654);
xor U5888 (N_5888,N_5734,N_5613);
and U5889 (N_5889,N_5647,N_5624);
and U5890 (N_5890,N_5704,N_5737);
or U5891 (N_5891,N_5616,N_5745);
and U5892 (N_5892,N_5631,N_5674);
nor U5893 (N_5893,N_5762,N_5645);
nand U5894 (N_5894,N_5728,N_5715);
or U5895 (N_5895,N_5652,N_5606);
nand U5896 (N_5896,N_5634,N_5685);
and U5897 (N_5897,N_5747,N_5689);
nand U5898 (N_5898,N_5784,N_5748);
nor U5899 (N_5899,N_5672,N_5750);
and U5900 (N_5900,N_5610,N_5788);
nor U5901 (N_5901,N_5742,N_5629);
or U5902 (N_5902,N_5646,N_5768);
nand U5903 (N_5903,N_5742,N_5643);
nor U5904 (N_5904,N_5781,N_5754);
and U5905 (N_5905,N_5770,N_5719);
nor U5906 (N_5906,N_5733,N_5677);
and U5907 (N_5907,N_5663,N_5727);
or U5908 (N_5908,N_5791,N_5680);
nand U5909 (N_5909,N_5799,N_5692);
xor U5910 (N_5910,N_5699,N_5728);
or U5911 (N_5911,N_5638,N_5623);
and U5912 (N_5912,N_5631,N_5671);
nand U5913 (N_5913,N_5601,N_5685);
nand U5914 (N_5914,N_5634,N_5770);
nand U5915 (N_5915,N_5630,N_5692);
nand U5916 (N_5916,N_5651,N_5674);
nand U5917 (N_5917,N_5721,N_5745);
and U5918 (N_5918,N_5760,N_5632);
and U5919 (N_5919,N_5730,N_5690);
nand U5920 (N_5920,N_5677,N_5793);
or U5921 (N_5921,N_5776,N_5743);
and U5922 (N_5922,N_5767,N_5621);
nand U5923 (N_5923,N_5709,N_5735);
nor U5924 (N_5924,N_5663,N_5710);
nor U5925 (N_5925,N_5703,N_5615);
and U5926 (N_5926,N_5797,N_5673);
nor U5927 (N_5927,N_5770,N_5797);
and U5928 (N_5928,N_5701,N_5712);
and U5929 (N_5929,N_5726,N_5643);
xnor U5930 (N_5930,N_5614,N_5655);
or U5931 (N_5931,N_5667,N_5624);
nor U5932 (N_5932,N_5771,N_5618);
nor U5933 (N_5933,N_5706,N_5663);
or U5934 (N_5934,N_5695,N_5667);
or U5935 (N_5935,N_5736,N_5631);
and U5936 (N_5936,N_5737,N_5620);
and U5937 (N_5937,N_5606,N_5771);
or U5938 (N_5938,N_5689,N_5786);
xor U5939 (N_5939,N_5744,N_5734);
or U5940 (N_5940,N_5755,N_5717);
and U5941 (N_5941,N_5758,N_5628);
xor U5942 (N_5942,N_5686,N_5736);
xnor U5943 (N_5943,N_5604,N_5720);
xor U5944 (N_5944,N_5651,N_5625);
nor U5945 (N_5945,N_5689,N_5712);
nand U5946 (N_5946,N_5778,N_5793);
nor U5947 (N_5947,N_5796,N_5682);
xor U5948 (N_5948,N_5789,N_5636);
or U5949 (N_5949,N_5741,N_5625);
nand U5950 (N_5950,N_5719,N_5789);
and U5951 (N_5951,N_5669,N_5745);
nor U5952 (N_5952,N_5798,N_5607);
nor U5953 (N_5953,N_5726,N_5778);
and U5954 (N_5954,N_5667,N_5607);
xor U5955 (N_5955,N_5612,N_5770);
nand U5956 (N_5956,N_5655,N_5674);
or U5957 (N_5957,N_5698,N_5787);
nand U5958 (N_5958,N_5683,N_5764);
nand U5959 (N_5959,N_5656,N_5686);
nor U5960 (N_5960,N_5697,N_5799);
xor U5961 (N_5961,N_5639,N_5667);
and U5962 (N_5962,N_5611,N_5787);
xor U5963 (N_5963,N_5632,N_5620);
nor U5964 (N_5964,N_5690,N_5696);
nor U5965 (N_5965,N_5756,N_5782);
nand U5966 (N_5966,N_5671,N_5728);
or U5967 (N_5967,N_5645,N_5629);
and U5968 (N_5968,N_5622,N_5725);
or U5969 (N_5969,N_5633,N_5730);
xnor U5970 (N_5970,N_5747,N_5707);
and U5971 (N_5971,N_5766,N_5628);
xor U5972 (N_5972,N_5605,N_5783);
nor U5973 (N_5973,N_5691,N_5612);
xor U5974 (N_5974,N_5614,N_5784);
xor U5975 (N_5975,N_5658,N_5679);
nor U5976 (N_5976,N_5694,N_5776);
and U5977 (N_5977,N_5706,N_5602);
nor U5978 (N_5978,N_5723,N_5637);
or U5979 (N_5979,N_5626,N_5734);
nand U5980 (N_5980,N_5776,N_5772);
or U5981 (N_5981,N_5689,N_5642);
xor U5982 (N_5982,N_5643,N_5719);
or U5983 (N_5983,N_5762,N_5633);
or U5984 (N_5984,N_5639,N_5797);
nand U5985 (N_5985,N_5794,N_5663);
xnor U5986 (N_5986,N_5661,N_5638);
or U5987 (N_5987,N_5712,N_5731);
xor U5988 (N_5988,N_5745,N_5612);
nor U5989 (N_5989,N_5669,N_5755);
and U5990 (N_5990,N_5627,N_5795);
nor U5991 (N_5991,N_5602,N_5708);
or U5992 (N_5992,N_5623,N_5695);
nand U5993 (N_5993,N_5661,N_5692);
and U5994 (N_5994,N_5768,N_5770);
or U5995 (N_5995,N_5769,N_5642);
nand U5996 (N_5996,N_5727,N_5601);
and U5997 (N_5997,N_5656,N_5639);
nor U5998 (N_5998,N_5645,N_5615);
or U5999 (N_5999,N_5674,N_5798);
xnor U6000 (N_6000,N_5800,N_5861);
xnor U6001 (N_6001,N_5806,N_5980);
nand U6002 (N_6002,N_5839,N_5901);
xnor U6003 (N_6003,N_5906,N_5949);
nor U6004 (N_6004,N_5928,N_5903);
nand U6005 (N_6005,N_5878,N_5993);
or U6006 (N_6006,N_5907,N_5852);
nand U6007 (N_6007,N_5879,N_5837);
and U6008 (N_6008,N_5963,N_5825);
or U6009 (N_6009,N_5977,N_5909);
nor U6010 (N_6010,N_5941,N_5944);
xor U6011 (N_6011,N_5926,N_5898);
nand U6012 (N_6012,N_5889,N_5845);
and U6013 (N_6013,N_5976,N_5814);
nor U6014 (N_6014,N_5885,N_5816);
nand U6015 (N_6015,N_5994,N_5959);
and U6016 (N_6016,N_5831,N_5841);
and U6017 (N_6017,N_5855,N_5829);
xnor U6018 (N_6018,N_5821,N_5844);
or U6019 (N_6019,N_5988,N_5848);
and U6020 (N_6020,N_5914,N_5937);
nand U6021 (N_6021,N_5948,N_5896);
xnor U6022 (N_6022,N_5902,N_5953);
or U6023 (N_6023,N_5972,N_5862);
or U6024 (N_6024,N_5875,N_5849);
and U6025 (N_6025,N_5812,N_5854);
nand U6026 (N_6026,N_5983,N_5815);
and U6027 (N_6027,N_5888,N_5882);
or U6028 (N_6028,N_5807,N_5874);
nor U6029 (N_6029,N_5921,N_5964);
nand U6030 (N_6030,N_5801,N_5883);
nand U6031 (N_6031,N_5984,N_5819);
nor U6032 (N_6032,N_5927,N_5917);
xor U6033 (N_6033,N_5895,N_5833);
or U6034 (N_6034,N_5870,N_5938);
nand U6035 (N_6035,N_5804,N_5967);
and U6036 (N_6036,N_5891,N_5805);
xor U6037 (N_6037,N_5824,N_5872);
and U6038 (N_6038,N_5823,N_5956);
nor U6039 (N_6039,N_5913,N_5915);
or U6040 (N_6040,N_5960,N_5982);
and U6041 (N_6041,N_5985,N_5971);
nor U6042 (N_6042,N_5951,N_5857);
nor U6043 (N_6043,N_5865,N_5905);
or U6044 (N_6044,N_5850,N_5822);
and U6045 (N_6045,N_5899,N_5999);
and U6046 (N_6046,N_5890,N_5990);
nand U6047 (N_6047,N_5893,N_5920);
or U6048 (N_6048,N_5897,N_5877);
nor U6049 (N_6049,N_5908,N_5876);
and U6050 (N_6050,N_5946,N_5832);
or U6051 (N_6051,N_5974,N_5813);
nand U6052 (N_6052,N_5863,N_5945);
or U6053 (N_6053,N_5916,N_5842);
and U6054 (N_6054,N_5970,N_5978);
or U6055 (N_6055,N_5904,N_5851);
nand U6056 (N_6056,N_5900,N_5838);
or U6057 (N_6057,N_5931,N_5886);
nor U6058 (N_6058,N_5939,N_5818);
nor U6059 (N_6059,N_5968,N_5962);
xnor U6060 (N_6060,N_5830,N_5979);
nor U6061 (N_6061,N_5986,N_5910);
nor U6062 (N_6062,N_5933,N_5894);
xnor U6063 (N_6063,N_5892,N_5998);
xor U6064 (N_6064,N_5820,N_5932);
xor U6065 (N_6065,N_5943,N_5924);
nand U6066 (N_6066,N_5961,N_5834);
xor U6067 (N_6067,N_5952,N_5836);
nand U6068 (N_6068,N_5973,N_5846);
xor U6069 (N_6069,N_5940,N_5930);
nand U6070 (N_6070,N_5992,N_5811);
or U6071 (N_6071,N_5826,N_5969);
xor U6072 (N_6072,N_5867,N_5955);
nand U6073 (N_6073,N_5802,N_5966);
nand U6074 (N_6074,N_5869,N_5871);
nor U6075 (N_6075,N_5942,N_5873);
and U6076 (N_6076,N_5996,N_5843);
nand U6077 (N_6077,N_5860,N_5840);
or U6078 (N_6078,N_5981,N_5936);
nor U6079 (N_6079,N_5997,N_5958);
xor U6080 (N_6080,N_5950,N_5864);
nand U6081 (N_6081,N_5995,N_5817);
xnor U6082 (N_6082,N_5853,N_5957);
xnor U6083 (N_6083,N_5856,N_5919);
nand U6084 (N_6084,N_5847,N_5918);
nor U6085 (N_6085,N_5954,N_5868);
or U6086 (N_6086,N_5935,N_5987);
xnor U6087 (N_6087,N_5881,N_5827);
nand U6088 (N_6088,N_5912,N_5934);
and U6089 (N_6089,N_5929,N_5947);
and U6090 (N_6090,N_5925,N_5880);
or U6091 (N_6091,N_5866,N_5835);
and U6092 (N_6092,N_5989,N_5803);
xnor U6093 (N_6093,N_5828,N_5975);
nor U6094 (N_6094,N_5858,N_5808);
nor U6095 (N_6095,N_5922,N_5991);
nor U6096 (N_6096,N_5884,N_5859);
nor U6097 (N_6097,N_5887,N_5923);
nor U6098 (N_6098,N_5965,N_5810);
xnor U6099 (N_6099,N_5911,N_5809);
and U6100 (N_6100,N_5927,N_5947);
xnor U6101 (N_6101,N_5867,N_5835);
xor U6102 (N_6102,N_5922,N_5810);
nand U6103 (N_6103,N_5868,N_5901);
and U6104 (N_6104,N_5930,N_5889);
nor U6105 (N_6105,N_5999,N_5893);
nor U6106 (N_6106,N_5991,N_5906);
nand U6107 (N_6107,N_5897,N_5874);
nor U6108 (N_6108,N_5888,N_5859);
nor U6109 (N_6109,N_5928,N_5827);
nand U6110 (N_6110,N_5981,N_5939);
or U6111 (N_6111,N_5800,N_5888);
nand U6112 (N_6112,N_5859,N_5957);
nor U6113 (N_6113,N_5949,N_5856);
or U6114 (N_6114,N_5860,N_5915);
or U6115 (N_6115,N_5816,N_5964);
or U6116 (N_6116,N_5981,N_5883);
nand U6117 (N_6117,N_5958,N_5919);
nand U6118 (N_6118,N_5975,N_5841);
xor U6119 (N_6119,N_5839,N_5990);
nor U6120 (N_6120,N_5913,N_5834);
nand U6121 (N_6121,N_5881,N_5987);
and U6122 (N_6122,N_5920,N_5888);
and U6123 (N_6123,N_5987,N_5969);
nand U6124 (N_6124,N_5972,N_5904);
nand U6125 (N_6125,N_5847,N_5858);
xor U6126 (N_6126,N_5876,N_5868);
or U6127 (N_6127,N_5868,N_5926);
nor U6128 (N_6128,N_5808,N_5902);
nand U6129 (N_6129,N_5815,N_5860);
and U6130 (N_6130,N_5897,N_5928);
or U6131 (N_6131,N_5909,N_5913);
xor U6132 (N_6132,N_5826,N_5860);
nand U6133 (N_6133,N_5836,N_5972);
xor U6134 (N_6134,N_5834,N_5969);
and U6135 (N_6135,N_5973,N_5929);
nand U6136 (N_6136,N_5925,N_5931);
or U6137 (N_6137,N_5970,N_5894);
or U6138 (N_6138,N_5882,N_5904);
nand U6139 (N_6139,N_5852,N_5859);
nand U6140 (N_6140,N_5916,N_5823);
nand U6141 (N_6141,N_5808,N_5911);
or U6142 (N_6142,N_5904,N_5891);
xor U6143 (N_6143,N_5818,N_5839);
nand U6144 (N_6144,N_5917,N_5959);
or U6145 (N_6145,N_5988,N_5887);
nor U6146 (N_6146,N_5816,N_5878);
nand U6147 (N_6147,N_5995,N_5868);
nor U6148 (N_6148,N_5823,N_5806);
nor U6149 (N_6149,N_5937,N_5904);
and U6150 (N_6150,N_5960,N_5965);
or U6151 (N_6151,N_5920,N_5830);
and U6152 (N_6152,N_5999,N_5990);
xnor U6153 (N_6153,N_5932,N_5908);
xor U6154 (N_6154,N_5835,N_5889);
nor U6155 (N_6155,N_5828,N_5963);
and U6156 (N_6156,N_5999,N_5866);
nor U6157 (N_6157,N_5840,N_5886);
nor U6158 (N_6158,N_5820,N_5988);
or U6159 (N_6159,N_5810,N_5951);
nor U6160 (N_6160,N_5984,N_5976);
nand U6161 (N_6161,N_5966,N_5805);
xnor U6162 (N_6162,N_5933,N_5966);
and U6163 (N_6163,N_5959,N_5987);
xor U6164 (N_6164,N_5969,N_5802);
and U6165 (N_6165,N_5806,N_5863);
nor U6166 (N_6166,N_5974,N_5987);
nand U6167 (N_6167,N_5849,N_5861);
xor U6168 (N_6168,N_5825,N_5934);
or U6169 (N_6169,N_5982,N_5802);
xnor U6170 (N_6170,N_5900,N_5906);
xor U6171 (N_6171,N_5961,N_5832);
nand U6172 (N_6172,N_5901,N_5894);
and U6173 (N_6173,N_5911,N_5928);
nand U6174 (N_6174,N_5890,N_5913);
or U6175 (N_6175,N_5896,N_5976);
nor U6176 (N_6176,N_5885,N_5913);
or U6177 (N_6177,N_5912,N_5991);
xor U6178 (N_6178,N_5986,N_5800);
or U6179 (N_6179,N_5846,N_5963);
and U6180 (N_6180,N_5950,N_5828);
xor U6181 (N_6181,N_5955,N_5886);
nor U6182 (N_6182,N_5922,N_5893);
and U6183 (N_6183,N_5958,N_5841);
nand U6184 (N_6184,N_5925,N_5917);
nand U6185 (N_6185,N_5967,N_5893);
or U6186 (N_6186,N_5940,N_5907);
or U6187 (N_6187,N_5884,N_5951);
xor U6188 (N_6188,N_5853,N_5877);
or U6189 (N_6189,N_5962,N_5983);
and U6190 (N_6190,N_5928,N_5991);
or U6191 (N_6191,N_5813,N_5902);
nand U6192 (N_6192,N_5894,N_5815);
nand U6193 (N_6193,N_5966,N_5857);
or U6194 (N_6194,N_5926,N_5932);
and U6195 (N_6195,N_5993,N_5985);
nor U6196 (N_6196,N_5874,N_5811);
and U6197 (N_6197,N_5922,N_5939);
and U6198 (N_6198,N_5858,N_5981);
or U6199 (N_6199,N_5862,N_5926);
nand U6200 (N_6200,N_6101,N_6197);
and U6201 (N_6201,N_6105,N_6170);
nand U6202 (N_6202,N_6097,N_6060);
nand U6203 (N_6203,N_6146,N_6087);
nor U6204 (N_6204,N_6137,N_6028);
nor U6205 (N_6205,N_6190,N_6051);
or U6206 (N_6206,N_6021,N_6042);
and U6207 (N_6207,N_6127,N_6052);
nor U6208 (N_6208,N_6158,N_6120);
and U6209 (N_6209,N_6050,N_6187);
or U6210 (N_6210,N_6186,N_6129);
or U6211 (N_6211,N_6126,N_6020);
and U6212 (N_6212,N_6108,N_6037);
nand U6213 (N_6213,N_6139,N_6025);
nand U6214 (N_6214,N_6176,N_6059);
nor U6215 (N_6215,N_6089,N_6111);
or U6216 (N_6216,N_6093,N_6068);
or U6217 (N_6217,N_6173,N_6065);
and U6218 (N_6218,N_6143,N_6110);
xnor U6219 (N_6219,N_6177,N_6026);
xnor U6220 (N_6220,N_6081,N_6144);
nor U6221 (N_6221,N_6077,N_6045);
and U6222 (N_6222,N_6189,N_6011);
and U6223 (N_6223,N_6024,N_6083);
nand U6224 (N_6224,N_6073,N_6099);
nor U6225 (N_6225,N_6191,N_6049);
nor U6226 (N_6226,N_6172,N_6138);
nor U6227 (N_6227,N_6062,N_6182);
and U6228 (N_6228,N_6032,N_6174);
and U6229 (N_6229,N_6076,N_6074);
or U6230 (N_6230,N_6167,N_6088);
and U6231 (N_6231,N_6107,N_6160);
nor U6232 (N_6232,N_6000,N_6057);
nand U6233 (N_6233,N_6161,N_6184);
xnor U6234 (N_6234,N_6165,N_6078);
nor U6235 (N_6235,N_6071,N_6112);
xnor U6236 (N_6236,N_6022,N_6106);
xnor U6237 (N_6237,N_6153,N_6118);
nor U6238 (N_6238,N_6154,N_6156);
or U6239 (N_6239,N_6103,N_6179);
xnor U6240 (N_6240,N_6023,N_6019);
and U6241 (N_6241,N_6058,N_6027);
nand U6242 (N_6242,N_6113,N_6157);
and U6243 (N_6243,N_6013,N_6125);
and U6244 (N_6244,N_6193,N_6055);
or U6245 (N_6245,N_6016,N_6119);
nor U6246 (N_6246,N_6043,N_6085);
and U6247 (N_6247,N_6151,N_6034);
xor U6248 (N_6248,N_6199,N_6084);
nand U6249 (N_6249,N_6039,N_6009);
nand U6250 (N_6250,N_6183,N_6185);
nand U6251 (N_6251,N_6123,N_6079);
nor U6252 (N_6252,N_6140,N_6192);
nor U6253 (N_6253,N_6072,N_6168);
and U6254 (N_6254,N_6116,N_6069);
xor U6255 (N_6255,N_6132,N_6117);
nor U6256 (N_6256,N_6086,N_6018);
nor U6257 (N_6257,N_6029,N_6122);
and U6258 (N_6258,N_6036,N_6030);
and U6259 (N_6259,N_6003,N_6198);
xnor U6260 (N_6260,N_6100,N_6135);
nor U6261 (N_6261,N_6195,N_6096);
nand U6262 (N_6262,N_6038,N_6128);
xnor U6263 (N_6263,N_6005,N_6004);
and U6264 (N_6264,N_6066,N_6180);
or U6265 (N_6265,N_6044,N_6053);
or U6266 (N_6266,N_6136,N_6114);
nand U6267 (N_6267,N_6090,N_6035);
or U6268 (N_6268,N_6075,N_6142);
nand U6269 (N_6269,N_6147,N_6082);
nor U6270 (N_6270,N_6002,N_6010);
nor U6271 (N_6271,N_6054,N_6094);
nand U6272 (N_6272,N_6041,N_6091);
nand U6273 (N_6273,N_6063,N_6092);
nand U6274 (N_6274,N_6015,N_6007);
xnor U6275 (N_6275,N_6056,N_6001);
nor U6276 (N_6276,N_6163,N_6064);
nor U6277 (N_6277,N_6150,N_6171);
and U6278 (N_6278,N_6169,N_6115);
xor U6279 (N_6279,N_6012,N_6008);
or U6280 (N_6280,N_6188,N_6006);
xor U6281 (N_6281,N_6134,N_6148);
and U6282 (N_6282,N_6155,N_6047);
or U6283 (N_6283,N_6162,N_6124);
or U6284 (N_6284,N_6067,N_6133);
or U6285 (N_6285,N_6102,N_6061);
xnor U6286 (N_6286,N_6194,N_6178);
xor U6287 (N_6287,N_6164,N_6130);
nor U6288 (N_6288,N_6181,N_6080);
nor U6289 (N_6289,N_6109,N_6046);
nor U6290 (N_6290,N_6014,N_6196);
and U6291 (N_6291,N_6149,N_6095);
xor U6292 (N_6292,N_6098,N_6104);
nor U6293 (N_6293,N_6131,N_6017);
nor U6294 (N_6294,N_6033,N_6152);
and U6295 (N_6295,N_6031,N_6048);
nor U6296 (N_6296,N_6159,N_6040);
xnor U6297 (N_6297,N_6166,N_6141);
nor U6298 (N_6298,N_6070,N_6121);
xnor U6299 (N_6299,N_6145,N_6175);
or U6300 (N_6300,N_6157,N_6154);
nor U6301 (N_6301,N_6019,N_6135);
or U6302 (N_6302,N_6069,N_6130);
nand U6303 (N_6303,N_6195,N_6170);
and U6304 (N_6304,N_6079,N_6133);
or U6305 (N_6305,N_6032,N_6177);
xor U6306 (N_6306,N_6132,N_6080);
nor U6307 (N_6307,N_6075,N_6125);
nor U6308 (N_6308,N_6132,N_6021);
and U6309 (N_6309,N_6004,N_6100);
and U6310 (N_6310,N_6172,N_6068);
xor U6311 (N_6311,N_6065,N_6137);
xor U6312 (N_6312,N_6091,N_6184);
xor U6313 (N_6313,N_6171,N_6106);
or U6314 (N_6314,N_6130,N_6178);
nor U6315 (N_6315,N_6167,N_6132);
xor U6316 (N_6316,N_6021,N_6030);
nand U6317 (N_6317,N_6014,N_6053);
xnor U6318 (N_6318,N_6166,N_6022);
xor U6319 (N_6319,N_6045,N_6032);
nand U6320 (N_6320,N_6180,N_6012);
nor U6321 (N_6321,N_6103,N_6065);
and U6322 (N_6322,N_6183,N_6081);
nor U6323 (N_6323,N_6197,N_6070);
xnor U6324 (N_6324,N_6128,N_6049);
nor U6325 (N_6325,N_6142,N_6194);
and U6326 (N_6326,N_6000,N_6042);
xor U6327 (N_6327,N_6150,N_6027);
nand U6328 (N_6328,N_6123,N_6140);
and U6329 (N_6329,N_6153,N_6091);
and U6330 (N_6330,N_6015,N_6129);
xnor U6331 (N_6331,N_6146,N_6075);
or U6332 (N_6332,N_6143,N_6080);
nand U6333 (N_6333,N_6146,N_6106);
xor U6334 (N_6334,N_6049,N_6148);
or U6335 (N_6335,N_6056,N_6080);
nand U6336 (N_6336,N_6067,N_6174);
and U6337 (N_6337,N_6123,N_6194);
nor U6338 (N_6338,N_6043,N_6151);
nor U6339 (N_6339,N_6026,N_6024);
xor U6340 (N_6340,N_6101,N_6069);
xor U6341 (N_6341,N_6130,N_6076);
or U6342 (N_6342,N_6160,N_6192);
nor U6343 (N_6343,N_6128,N_6178);
or U6344 (N_6344,N_6049,N_6077);
nor U6345 (N_6345,N_6061,N_6004);
nand U6346 (N_6346,N_6161,N_6172);
nor U6347 (N_6347,N_6079,N_6002);
or U6348 (N_6348,N_6063,N_6059);
nor U6349 (N_6349,N_6076,N_6174);
xnor U6350 (N_6350,N_6136,N_6169);
and U6351 (N_6351,N_6168,N_6186);
nor U6352 (N_6352,N_6004,N_6060);
and U6353 (N_6353,N_6045,N_6074);
nor U6354 (N_6354,N_6118,N_6012);
and U6355 (N_6355,N_6009,N_6189);
and U6356 (N_6356,N_6094,N_6184);
xnor U6357 (N_6357,N_6036,N_6184);
nor U6358 (N_6358,N_6181,N_6143);
and U6359 (N_6359,N_6192,N_6128);
or U6360 (N_6360,N_6036,N_6092);
xnor U6361 (N_6361,N_6133,N_6139);
and U6362 (N_6362,N_6178,N_6150);
or U6363 (N_6363,N_6010,N_6143);
nand U6364 (N_6364,N_6001,N_6077);
xnor U6365 (N_6365,N_6070,N_6013);
xnor U6366 (N_6366,N_6082,N_6104);
nand U6367 (N_6367,N_6141,N_6111);
and U6368 (N_6368,N_6199,N_6154);
nand U6369 (N_6369,N_6088,N_6180);
nor U6370 (N_6370,N_6044,N_6039);
or U6371 (N_6371,N_6118,N_6182);
or U6372 (N_6372,N_6154,N_6134);
nand U6373 (N_6373,N_6015,N_6035);
or U6374 (N_6374,N_6034,N_6035);
xnor U6375 (N_6375,N_6184,N_6122);
nor U6376 (N_6376,N_6093,N_6065);
and U6377 (N_6377,N_6107,N_6172);
xnor U6378 (N_6378,N_6020,N_6047);
and U6379 (N_6379,N_6066,N_6156);
nor U6380 (N_6380,N_6154,N_6123);
and U6381 (N_6381,N_6014,N_6127);
or U6382 (N_6382,N_6106,N_6017);
nor U6383 (N_6383,N_6139,N_6033);
xor U6384 (N_6384,N_6188,N_6031);
nor U6385 (N_6385,N_6140,N_6119);
nand U6386 (N_6386,N_6082,N_6178);
and U6387 (N_6387,N_6093,N_6092);
or U6388 (N_6388,N_6188,N_6152);
or U6389 (N_6389,N_6166,N_6077);
xnor U6390 (N_6390,N_6064,N_6099);
or U6391 (N_6391,N_6185,N_6087);
nor U6392 (N_6392,N_6052,N_6145);
xnor U6393 (N_6393,N_6134,N_6114);
and U6394 (N_6394,N_6030,N_6073);
or U6395 (N_6395,N_6187,N_6062);
or U6396 (N_6396,N_6078,N_6115);
xor U6397 (N_6397,N_6094,N_6157);
nor U6398 (N_6398,N_6084,N_6014);
nand U6399 (N_6399,N_6087,N_6077);
or U6400 (N_6400,N_6277,N_6302);
and U6401 (N_6401,N_6237,N_6337);
nand U6402 (N_6402,N_6306,N_6280);
and U6403 (N_6403,N_6398,N_6228);
and U6404 (N_6404,N_6342,N_6386);
nor U6405 (N_6405,N_6311,N_6396);
nand U6406 (N_6406,N_6221,N_6326);
and U6407 (N_6407,N_6297,N_6270);
xor U6408 (N_6408,N_6225,N_6314);
nor U6409 (N_6409,N_6364,N_6298);
xnor U6410 (N_6410,N_6262,N_6344);
nor U6411 (N_6411,N_6282,N_6211);
xor U6412 (N_6412,N_6365,N_6208);
nor U6413 (N_6413,N_6328,N_6230);
nand U6414 (N_6414,N_6254,N_6369);
or U6415 (N_6415,N_6374,N_6336);
or U6416 (N_6416,N_6257,N_6261);
or U6417 (N_6417,N_6216,N_6347);
and U6418 (N_6418,N_6331,N_6395);
and U6419 (N_6419,N_6391,N_6332);
nor U6420 (N_6420,N_6379,N_6383);
or U6421 (N_6421,N_6264,N_6368);
nand U6422 (N_6422,N_6291,N_6233);
and U6423 (N_6423,N_6327,N_6317);
nand U6424 (N_6424,N_6325,N_6222);
or U6425 (N_6425,N_6318,N_6371);
nand U6426 (N_6426,N_6350,N_6323);
xnor U6427 (N_6427,N_6312,N_6346);
nor U6428 (N_6428,N_6219,N_6355);
xnor U6429 (N_6429,N_6360,N_6266);
nand U6430 (N_6430,N_6315,N_6235);
or U6431 (N_6431,N_6263,N_6210);
nor U6432 (N_6432,N_6231,N_6308);
xor U6433 (N_6433,N_6265,N_6375);
or U6434 (N_6434,N_6259,N_6351);
nand U6435 (N_6435,N_6304,N_6349);
or U6436 (N_6436,N_6240,N_6388);
or U6437 (N_6437,N_6394,N_6341);
nand U6438 (N_6438,N_6376,N_6275);
and U6439 (N_6439,N_6258,N_6253);
nor U6440 (N_6440,N_6358,N_6252);
xor U6441 (N_6441,N_6356,N_6373);
nand U6442 (N_6442,N_6378,N_6239);
nor U6443 (N_6443,N_6289,N_6354);
xor U6444 (N_6444,N_6370,N_6305);
nand U6445 (N_6445,N_6292,N_6392);
xor U6446 (N_6446,N_6256,N_6202);
nand U6447 (N_6447,N_6301,N_6322);
and U6448 (N_6448,N_6321,N_6307);
or U6449 (N_6449,N_6242,N_6377);
or U6450 (N_6450,N_6381,N_6224);
nand U6451 (N_6451,N_6284,N_6296);
nor U6452 (N_6452,N_6330,N_6212);
xor U6453 (N_6453,N_6313,N_6290);
xnor U6454 (N_6454,N_6207,N_6385);
nand U6455 (N_6455,N_6293,N_6361);
nor U6456 (N_6456,N_6299,N_6203);
or U6457 (N_6457,N_6279,N_6229);
xnor U6458 (N_6458,N_6272,N_6324);
nor U6459 (N_6459,N_6226,N_6362);
nor U6460 (N_6460,N_6204,N_6287);
nor U6461 (N_6461,N_6363,N_6393);
nand U6462 (N_6462,N_6281,N_6294);
xnor U6463 (N_6463,N_6276,N_6340);
xor U6464 (N_6464,N_6345,N_6335);
nor U6465 (N_6465,N_6223,N_6251);
nand U6466 (N_6466,N_6234,N_6397);
nand U6467 (N_6467,N_6384,N_6329);
nor U6468 (N_6468,N_6288,N_6300);
nor U6469 (N_6469,N_6260,N_6250);
and U6470 (N_6470,N_6205,N_6236);
or U6471 (N_6471,N_6241,N_6320);
and U6472 (N_6472,N_6334,N_6227);
or U6473 (N_6473,N_6246,N_6389);
nor U6474 (N_6474,N_6244,N_6285);
nor U6475 (N_6475,N_6303,N_6218);
nor U6476 (N_6476,N_6399,N_6215);
and U6477 (N_6477,N_6209,N_6338);
nand U6478 (N_6478,N_6201,N_6232);
nand U6479 (N_6479,N_6309,N_6238);
and U6480 (N_6480,N_6206,N_6372);
and U6481 (N_6481,N_6255,N_6357);
xnor U6482 (N_6482,N_6367,N_6359);
nor U6483 (N_6483,N_6353,N_6286);
nor U6484 (N_6484,N_6248,N_6352);
or U6485 (N_6485,N_6339,N_6333);
or U6486 (N_6486,N_6214,N_6278);
nand U6487 (N_6487,N_6343,N_6213);
nand U6488 (N_6488,N_6319,N_6366);
nand U6489 (N_6489,N_6268,N_6271);
nand U6490 (N_6490,N_6382,N_6295);
nand U6491 (N_6491,N_6310,N_6217);
nor U6492 (N_6492,N_6249,N_6274);
and U6493 (N_6493,N_6387,N_6220);
or U6494 (N_6494,N_6243,N_6267);
and U6495 (N_6495,N_6273,N_6269);
nor U6496 (N_6496,N_6316,N_6348);
nor U6497 (N_6497,N_6380,N_6245);
xor U6498 (N_6498,N_6247,N_6283);
xor U6499 (N_6499,N_6390,N_6200);
xnor U6500 (N_6500,N_6224,N_6371);
and U6501 (N_6501,N_6249,N_6336);
and U6502 (N_6502,N_6268,N_6284);
nand U6503 (N_6503,N_6337,N_6311);
xnor U6504 (N_6504,N_6320,N_6290);
and U6505 (N_6505,N_6232,N_6351);
nor U6506 (N_6506,N_6312,N_6294);
nor U6507 (N_6507,N_6337,N_6382);
and U6508 (N_6508,N_6364,N_6279);
nor U6509 (N_6509,N_6238,N_6342);
xor U6510 (N_6510,N_6239,N_6210);
or U6511 (N_6511,N_6212,N_6225);
xnor U6512 (N_6512,N_6356,N_6371);
nor U6513 (N_6513,N_6328,N_6211);
nand U6514 (N_6514,N_6377,N_6369);
and U6515 (N_6515,N_6235,N_6381);
nor U6516 (N_6516,N_6327,N_6353);
and U6517 (N_6517,N_6310,N_6360);
nor U6518 (N_6518,N_6311,N_6257);
nor U6519 (N_6519,N_6245,N_6314);
and U6520 (N_6520,N_6388,N_6202);
xor U6521 (N_6521,N_6370,N_6265);
nor U6522 (N_6522,N_6310,N_6328);
or U6523 (N_6523,N_6314,N_6328);
xor U6524 (N_6524,N_6235,N_6307);
or U6525 (N_6525,N_6285,N_6286);
and U6526 (N_6526,N_6299,N_6265);
xnor U6527 (N_6527,N_6249,N_6388);
nor U6528 (N_6528,N_6208,N_6239);
nand U6529 (N_6529,N_6369,N_6268);
nor U6530 (N_6530,N_6295,N_6224);
xor U6531 (N_6531,N_6316,N_6272);
and U6532 (N_6532,N_6302,N_6235);
and U6533 (N_6533,N_6223,N_6395);
or U6534 (N_6534,N_6372,N_6239);
xor U6535 (N_6535,N_6222,N_6225);
nand U6536 (N_6536,N_6370,N_6383);
or U6537 (N_6537,N_6363,N_6299);
nor U6538 (N_6538,N_6337,N_6350);
and U6539 (N_6539,N_6285,N_6304);
nand U6540 (N_6540,N_6330,N_6215);
xor U6541 (N_6541,N_6241,N_6238);
or U6542 (N_6542,N_6342,N_6282);
or U6543 (N_6543,N_6391,N_6379);
nand U6544 (N_6544,N_6346,N_6288);
nand U6545 (N_6545,N_6280,N_6358);
nor U6546 (N_6546,N_6320,N_6231);
xnor U6547 (N_6547,N_6387,N_6200);
xor U6548 (N_6548,N_6216,N_6305);
xor U6549 (N_6549,N_6202,N_6350);
or U6550 (N_6550,N_6247,N_6302);
or U6551 (N_6551,N_6355,N_6267);
nor U6552 (N_6552,N_6253,N_6371);
xnor U6553 (N_6553,N_6300,N_6298);
and U6554 (N_6554,N_6289,N_6378);
xnor U6555 (N_6555,N_6287,N_6260);
and U6556 (N_6556,N_6344,N_6275);
or U6557 (N_6557,N_6305,N_6210);
and U6558 (N_6558,N_6391,N_6259);
nor U6559 (N_6559,N_6264,N_6270);
or U6560 (N_6560,N_6207,N_6342);
and U6561 (N_6561,N_6253,N_6296);
xor U6562 (N_6562,N_6311,N_6274);
xnor U6563 (N_6563,N_6329,N_6372);
and U6564 (N_6564,N_6379,N_6249);
or U6565 (N_6565,N_6253,N_6271);
and U6566 (N_6566,N_6390,N_6286);
nand U6567 (N_6567,N_6326,N_6232);
nor U6568 (N_6568,N_6318,N_6327);
and U6569 (N_6569,N_6337,N_6293);
or U6570 (N_6570,N_6280,N_6354);
nand U6571 (N_6571,N_6204,N_6208);
nand U6572 (N_6572,N_6333,N_6337);
and U6573 (N_6573,N_6219,N_6314);
and U6574 (N_6574,N_6223,N_6291);
nand U6575 (N_6575,N_6253,N_6306);
xnor U6576 (N_6576,N_6227,N_6207);
nor U6577 (N_6577,N_6215,N_6230);
and U6578 (N_6578,N_6327,N_6264);
and U6579 (N_6579,N_6319,N_6297);
and U6580 (N_6580,N_6339,N_6245);
or U6581 (N_6581,N_6210,N_6260);
or U6582 (N_6582,N_6383,N_6279);
nand U6583 (N_6583,N_6300,N_6343);
xnor U6584 (N_6584,N_6215,N_6326);
and U6585 (N_6585,N_6237,N_6365);
nand U6586 (N_6586,N_6264,N_6329);
xnor U6587 (N_6587,N_6254,N_6379);
or U6588 (N_6588,N_6275,N_6268);
nand U6589 (N_6589,N_6393,N_6203);
or U6590 (N_6590,N_6360,N_6209);
xnor U6591 (N_6591,N_6209,N_6224);
and U6592 (N_6592,N_6217,N_6224);
nand U6593 (N_6593,N_6294,N_6379);
xor U6594 (N_6594,N_6326,N_6302);
nand U6595 (N_6595,N_6367,N_6355);
nor U6596 (N_6596,N_6384,N_6313);
and U6597 (N_6597,N_6284,N_6281);
nand U6598 (N_6598,N_6395,N_6314);
or U6599 (N_6599,N_6357,N_6353);
xnor U6600 (N_6600,N_6464,N_6560);
nand U6601 (N_6601,N_6438,N_6584);
or U6602 (N_6602,N_6477,N_6463);
nand U6603 (N_6603,N_6567,N_6515);
nand U6604 (N_6604,N_6586,N_6530);
or U6605 (N_6605,N_6525,N_6471);
or U6606 (N_6606,N_6565,N_6541);
xor U6607 (N_6607,N_6483,N_6572);
nand U6608 (N_6608,N_6418,N_6454);
nor U6609 (N_6609,N_6547,N_6408);
nor U6610 (N_6610,N_6439,N_6594);
nor U6611 (N_6611,N_6577,N_6410);
xor U6612 (N_6612,N_6513,N_6435);
and U6613 (N_6613,N_6568,N_6516);
nor U6614 (N_6614,N_6589,N_6544);
nor U6615 (N_6615,N_6585,N_6531);
xnor U6616 (N_6616,N_6412,N_6534);
xor U6617 (N_6617,N_6543,N_6593);
or U6618 (N_6618,N_6555,N_6432);
and U6619 (N_6619,N_6479,N_6413);
nor U6620 (N_6620,N_6521,N_6490);
nand U6621 (N_6621,N_6448,N_6427);
or U6622 (N_6622,N_6480,N_6474);
and U6623 (N_6623,N_6491,N_6403);
nor U6624 (N_6624,N_6506,N_6465);
nand U6625 (N_6625,N_6424,N_6468);
xor U6626 (N_6626,N_6504,N_6536);
xor U6627 (N_6627,N_6466,N_6523);
xor U6628 (N_6628,N_6422,N_6539);
or U6629 (N_6629,N_6545,N_6533);
xnor U6630 (N_6630,N_6417,N_6467);
nor U6631 (N_6631,N_6546,N_6590);
and U6632 (N_6632,N_6538,N_6442);
and U6633 (N_6633,N_6542,N_6524);
nand U6634 (N_6634,N_6475,N_6420);
xnor U6635 (N_6635,N_6532,N_6401);
nor U6636 (N_6636,N_6592,N_6486);
and U6637 (N_6637,N_6429,N_6453);
xnor U6638 (N_6638,N_6574,N_6457);
and U6639 (N_6639,N_6423,N_6558);
nor U6640 (N_6640,N_6469,N_6409);
and U6641 (N_6641,N_6591,N_6582);
nand U6642 (N_6642,N_6443,N_6596);
nand U6643 (N_6643,N_6455,N_6562);
xnor U6644 (N_6644,N_6495,N_6419);
nor U6645 (N_6645,N_6487,N_6581);
nor U6646 (N_6646,N_6499,N_6470);
and U6647 (N_6647,N_6415,N_6440);
nor U6648 (N_6648,N_6407,N_6500);
nand U6649 (N_6649,N_6445,N_6484);
or U6650 (N_6650,N_6595,N_6553);
nor U6651 (N_6651,N_6598,N_6599);
or U6652 (N_6652,N_6450,N_6433);
xnor U6653 (N_6653,N_6497,N_6434);
and U6654 (N_6654,N_6489,N_6557);
nor U6655 (N_6655,N_6404,N_6556);
nor U6656 (N_6656,N_6402,N_6566);
nand U6657 (N_6657,N_6451,N_6548);
or U6658 (N_6658,N_6576,N_6520);
or U6659 (N_6659,N_6462,N_6549);
xnor U6660 (N_6660,N_6551,N_6405);
nand U6661 (N_6661,N_6570,N_6554);
nand U6662 (N_6662,N_6501,N_6441);
xnor U6663 (N_6663,N_6421,N_6411);
or U6664 (N_6664,N_6588,N_6456);
nand U6665 (N_6665,N_6571,N_6436);
and U6666 (N_6666,N_6459,N_6444);
xnor U6667 (N_6667,N_6452,N_6476);
nand U6668 (N_6668,N_6498,N_6587);
or U6669 (N_6669,N_6569,N_6430);
xor U6670 (N_6670,N_6488,N_6406);
nor U6671 (N_6671,N_6461,N_6561);
nand U6672 (N_6672,N_6496,N_6529);
xnor U6673 (N_6673,N_6522,N_6578);
or U6674 (N_6674,N_6507,N_6473);
nand U6675 (N_6675,N_6514,N_6519);
or U6676 (N_6676,N_6416,N_6447);
nand U6677 (N_6677,N_6400,N_6552);
nor U6678 (N_6678,N_6505,N_6414);
nor U6679 (N_6679,N_6425,N_6493);
xor U6680 (N_6680,N_6503,N_6509);
nor U6681 (N_6681,N_6472,N_6485);
nand U6682 (N_6682,N_6426,N_6460);
and U6683 (N_6683,N_6494,N_6437);
and U6684 (N_6684,N_6597,N_6540);
and U6685 (N_6685,N_6579,N_6550);
xnor U6686 (N_6686,N_6580,N_6446);
nand U6687 (N_6687,N_6478,N_6510);
xnor U6688 (N_6688,N_6583,N_6458);
and U6689 (N_6689,N_6575,N_6518);
or U6690 (N_6690,N_6428,N_6431);
nor U6691 (N_6691,N_6511,N_6492);
nor U6692 (N_6692,N_6481,N_6573);
xor U6693 (N_6693,N_6528,N_6559);
nand U6694 (N_6694,N_6526,N_6502);
nor U6695 (N_6695,N_6512,N_6537);
and U6696 (N_6696,N_6535,N_6508);
and U6697 (N_6697,N_6517,N_6527);
or U6698 (N_6698,N_6482,N_6563);
nor U6699 (N_6699,N_6564,N_6449);
or U6700 (N_6700,N_6546,N_6580);
or U6701 (N_6701,N_6537,N_6579);
nor U6702 (N_6702,N_6423,N_6549);
xor U6703 (N_6703,N_6585,N_6589);
nand U6704 (N_6704,N_6422,N_6508);
nor U6705 (N_6705,N_6427,N_6562);
and U6706 (N_6706,N_6523,N_6454);
and U6707 (N_6707,N_6585,N_6580);
and U6708 (N_6708,N_6451,N_6565);
nand U6709 (N_6709,N_6591,N_6463);
nor U6710 (N_6710,N_6426,N_6468);
and U6711 (N_6711,N_6478,N_6443);
xnor U6712 (N_6712,N_6424,N_6472);
xor U6713 (N_6713,N_6582,N_6588);
and U6714 (N_6714,N_6408,N_6481);
nor U6715 (N_6715,N_6403,N_6510);
and U6716 (N_6716,N_6465,N_6407);
and U6717 (N_6717,N_6481,N_6544);
xnor U6718 (N_6718,N_6483,N_6422);
nand U6719 (N_6719,N_6473,N_6597);
nand U6720 (N_6720,N_6418,N_6440);
and U6721 (N_6721,N_6518,N_6583);
or U6722 (N_6722,N_6461,N_6422);
xor U6723 (N_6723,N_6429,N_6566);
and U6724 (N_6724,N_6452,N_6426);
or U6725 (N_6725,N_6408,N_6508);
or U6726 (N_6726,N_6524,N_6513);
or U6727 (N_6727,N_6524,N_6451);
or U6728 (N_6728,N_6511,N_6552);
or U6729 (N_6729,N_6543,N_6471);
nor U6730 (N_6730,N_6552,N_6473);
or U6731 (N_6731,N_6534,N_6509);
nand U6732 (N_6732,N_6504,N_6596);
nor U6733 (N_6733,N_6531,N_6440);
and U6734 (N_6734,N_6563,N_6560);
xor U6735 (N_6735,N_6497,N_6408);
or U6736 (N_6736,N_6584,N_6455);
nor U6737 (N_6737,N_6479,N_6566);
and U6738 (N_6738,N_6434,N_6491);
nand U6739 (N_6739,N_6497,N_6459);
xor U6740 (N_6740,N_6530,N_6527);
or U6741 (N_6741,N_6587,N_6546);
or U6742 (N_6742,N_6521,N_6401);
nor U6743 (N_6743,N_6471,N_6446);
nor U6744 (N_6744,N_6547,N_6566);
nor U6745 (N_6745,N_6441,N_6411);
and U6746 (N_6746,N_6429,N_6569);
or U6747 (N_6747,N_6564,N_6548);
xnor U6748 (N_6748,N_6525,N_6408);
and U6749 (N_6749,N_6554,N_6473);
nand U6750 (N_6750,N_6511,N_6476);
nand U6751 (N_6751,N_6530,N_6468);
nor U6752 (N_6752,N_6551,N_6482);
nand U6753 (N_6753,N_6414,N_6520);
nor U6754 (N_6754,N_6481,N_6587);
xnor U6755 (N_6755,N_6453,N_6504);
nor U6756 (N_6756,N_6513,N_6585);
or U6757 (N_6757,N_6560,N_6403);
and U6758 (N_6758,N_6527,N_6474);
xor U6759 (N_6759,N_6422,N_6453);
nand U6760 (N_6760,N_6502,N_6505);
nor U6761 (N_6761,N_6581,N_6401);
or U6762 (N_6762,N_6463,N_6531);
nor U6763 (N_6763,N_6583,N_6568);
and U6764 (N_6764,N_6526,N_6447);
nand U6765 (N_6765,N_6482,N_6431);
and U6766 (N_6766,N_6577,N_6516);
or U6767 (N_6767,N_6441,N_6583);
nand U6768 (N_6768,N_6577,N_6568);
nand U6769 (N_6769,N_6439,N_6589);
nand U6770 (N_6770,N_6468,N_6459);
or U6771 (N_6771,N_6570,N_6432);
or U6772 (N_6772,N_6470,N_6588);
or U6773 (N_6773,N_6564,N_6412);
xnor U6774 (N_6774,N_6544,N_6426);
nor U6775 (N_6775,N_6474,N_6574);
nor U6776 (N_6776,N_6551,N_6564);
xnor U6777 (N_6777,N_6525,N_6436);
or U6778 (N_6778,N_6464,N_6582);
nand U6779 (N_6779,N_6435,N_6455);
or U6780 (N_6780,N_6571,N_6496);
nor U6781 (N_6781,N_6519,N_6549);
and U6782 (N_6782,N_6547,N_6507);
or U6783 (N_6783,N_6504,N_6490);
and U6784 (N_6784,N_6443,N_6539);
nand U6785 (N_6785,N_6507,N_6421);
nor U6786 (N_6786,N_6468,N_6404);
nand U6787 (N_6787,N_6585,N_6469);
or U6788 (N_6788,N_6471,N_6486);
and U6789 (N_6789,N_6493,N_6464);
or U6790 (N_6790,N_6563,N_6483);
or U6791 (N_6791,N_6489,N_6435);
nor U6792 (N_6792,N_6488,N_6490);
xor U6793 (N_6793,N_6430,N_6493);
xnor U6794 (N_6794,N_6426,N_6506);
nand U6795 (N_6795,N_6551,N_6529);
or U6796 (N_6796,N_6514,N_6468);
or U6797 (N_6797,N_6480,N_6517);
and U6798 (N_6798,N_6568,N_6541);
nand U6799 (N_6799,N_6464,N_6408);
or U6800 (N_6800,N_6788,N_6704);
nor U6801 (N_6801,N_6794,N_6737);
and U6802 (N_6802,N_6630,N_6757);
nand U6803 (N_6803,N_6735,N_6694);
and U6804 (N_6804,N_6612,N_6642);
nor U6805 (N_6805,N_6623,N_6751);
xnor U6806 (N_6806,N_6667,N_6746);
and U6807 (N_6807,N_6654,N_6635);
nor U6808 (N_6808,N_6738,N_6701);
nor U6809 (N_6809,N_6613,N_6793);
xnor U6810 (N_6810,N_6616,N_6674);
xor U6811 (N_6811,N_6703,N_6618);
nand U6812 (N_6812,N_6656,N_6740);
and U6813 (N_6813,N_6759,N_6789);
xnor U6814 (N_6814,N_6648,N_6784);
and U6815 (N_6815,N_6773,N_6614);
xor U6816 (N_6816,N_6795,N_6649);
nor U6817 (N_6817,N_6756,N_6763);
nor U6818 (N_6818,N_6710,N_6750);
or U6819 (N_6819,N_6605,N_6693);
and U6820 (N_6820,N_6624,N_6779);
nor U6821 (N_6821,N_6675,N_6657);
xnor U6822 (N_6822,N_6691,N_6732);
xnor U6823 (N_6823,N_6764,N_6603);
xor U6824 (N_6824,N_6730,N_6781);
and U6825 (N_6825,N_6765,N_6775);
nand U6826 (N_6826,N_6660,N_6606);
xor U6827 (N_6827,N_6709,N_6692);
or U6828 (N_6828,N_6714,N_6638);
xor U6829 (N_6829,N_6622,N_6698);
and U6830 (N_6830,N_6601,N_6680);
and U6831 (N_6831,N_6723,N_6604);
xnor U6832 (N_6832,N_6628,N_6672);
nand U6833 (N_6833,N_6625,N_6729);
or U6834 (N_6834,N_6780,N_6627);
or U6835 (N_6835,N_6719,N_6760);
xor U6836 (N_6836,N_6713,N_6762);
xor U6837 (N_6837,N_6696,N_6647);
and U6838 (N_6838,N_6676,N_6689);
xnor U6839 (N_6839,N_6639,N_6753);
nand U6840 (N_6840,N_6652,N_6786);
xor U6841 (N_6841,N_6743,N_6636);
nand U6842 (N_6842,N_6679,N_6705);
nand U6843 (N_6843,N_6621,N_6697);
nor U6844 (N_6844,N_6708,N_6699);
or U6845 (N_6845,N_6734,N_6620);
nand U6846 (N_6846,N_6783,N_6727);
nand U6847 (N_6847,N_6655,N_6641);
or U6848 (N_6848,N_6690,N_6798);
and U6849 (N_6849,N_6646,N_6758);
and U6850 (N_6850,N_6742,N_6650);
or U6851 (N_6851,N_6768,N_6711);
or U6852 (N_6852,N_6643,N_6683);
nand U6853 (N_6853,N_6633,N_6653);
and U6854 (N_6854,N_6769,N_6637);
nor U6855 (N_6855,N_6778,N_6761);
or U6856 (N_6856,N_6670,N_6748);
and U6857 (N_6857,N_6640,N_6752);
xnor U6858 (N_6858,N_6610,N_6695);
xor U6859 (N_6859,N_6725,N_6682);
nor U6860 (N_6860,N_6700,N_6722);
nand U6861 (N_6861,N_6777,N_6629);
nor U6862 (N_6862,N_6745,N_6688);
or U6863 (N_6863,N_6754,N_6790);
nand U6864 (N_6864,N_6792,N_6776);
or U6865 (N_6865,N_6669,N_6767);
nor U6866 (N_6866,N_6617,N_6717);
xor U6867 (N_6867,N_6782,N_6706);
or U6868 (N_6868,N_6681,N_6720);
and U6869 (N_6869,N_6771,N_6662);
xor U6870 (N_6870,N_6744,N_6685);
nand U6871 (N_6871,N_6770,N_6666);
nand U6872 (N_6872,N_6651,N_6600);
and U6873 (N_6873,N_6626,N_6684);
or U6874 (N_6874,N_6749,N_6772);
nand U6875 (N_6875,N_6632,N_6645);
and U6876 (N_6876,N_6728,N_6615);
nor U6877 (N_6877,N_6712,N_6671);
nor U6878 (N_6878,N_6631,N_6733);
or U6879 (N_6879,N_6668,N_6687);
nand U6880 (N_6880,N_6787,N_6707);
and U6881 (N_6881,N_6611,N_6608);
or U6882 (N_6882,N_6785,N_6673);
or U6883 (N_6883,N_6724,N_6796);
nor U6884 (N_6884,N_6659,N_6799);
nor U6885 (N_6885,N_6665,N_6686);
xnor U6886 (N_6886,N_6644,N_6774);
or U6887 (N_6887,N_6766,N_6741);
and U6888 (N_6888,N_6663,N_6678);
nor U6889 (N_6889,N_6661,N_6739);
xor U6890 (N_6890,N_6716,N_6602);
and U6891 (N_6891,N_6736,N_6791);
nand U6892 (N_6892,N_6634,N_6702);
nand U6893 (N_6893,N_6677,N_6731);
nand U6894 (N_6894,N_6755,N_6658);
xor U6895 (N_6895,N_6718,N_6607);
nand U6896 (N_6896,N_6747,N_6664);
xor U6897 (N_6897,N_6619,N_6797);
nor U6898 (N_6898,N_6726,N_6721);
and U6899 (N_6899,N_6609,N_6715);
nand U6900 (N_6900,N_6796,N_6721);
nand U6901 (N_6901,N_6646,N_6702);
and U6902 (N_6902,N_6756,N_6737);
xor U6903 (N_6903,N_6730,N_6680);
nor U6904 (N_6904,N_6723,N_6608);
nor U6905 (N_6905,N_6665,N_6716);
nand U6906 (N_6906,N_6794,N_6602);
xnor U6907 (N_6907,N_6788,N_6676);
nand U6908 (N_6908,N_6622,N_6741);
and U6909 (N_6909,N_6687,N_6616);
or U6910 (N_6910,N_6732,N_6638);
nand U6911 (N_6911,N_6639,N_6767);
nand U6912 (N_6912,N_6602,N_6766);
xnor U6913 (N_6913,N_6622,N_6670);
xnor U6914 (N_6914,N_6777,N_6670);
nand U6915 (N_6915,N_6638,N_6763);
xor U6916 (N_6916,N_6668,N_6768);
or U6917 (N_6917,N_6779,N_6722);
xnor U6918 (N_6918,N_6749,N_6618);
or U6919 (N_6919,N_6702,N_6686);
nor U6920 (N_6920,N_6621,N_6662);
xor U6921 (N_6921,N_6619,N_6708);
xor U6922 (N_6922,N_6640,N_6602);
or U6923 (N_6923,N_6761,N_6713);
or U6924 (N_6924,N_6654,N_6611);
nor U6925 (N_6925,N_6661,N_6680);
nor U6926 (N_6926,N_6682,N_6744);
nor U6927 (N_6927,N_6635,N_6639);
or U6928 (N_6928,N_6716,N_6727);
nor U6929 (N_6929,N_6759,N_6784);
and U6930 (N_6930,N_6717,N_6716);
or U6931 (N_6931,N_6712,N_6744);
nand U6932 (N_6932,N_6669,N_6664);
xnor U6933 (N_6933,N_6755,N_6696);
and U6934 (N_6934,N_6681,N_6609);
nor U6935 (N_6935,N_6773,N_6672);
or U6936 (N_6936,N_6623,N_6670);
nand U6937 (N_6937,N_6642,N_6741);
nand U6938 (N_6938,N_6746,N_6611);
nor U6939 (N_6939,N_6677,N_6729);
or U6940 (N_6940,N_6715,N_6797);
nor U6941 (N_6941,N_6776,N_6659);
or U6942 (N_6942,N_6632,N_6732);
nand U6943 (N_6943,N_6731,N_6626);
nor U6944 (N_6944,N_6752,N_6732);
or U6945 (N_6945,N_6667,N_6734);
or U6946 (N_6946,N_6624,N_6632);
or U6947 (N_6947,N_6781,N_6786);
nand U6948 (N_6948,N_6730,N_6776);
xnor U6949 (N_6949,N_6789,N_6742);
nand U6950 (N_6950,N_6651,N_6798);
and U6951 (N_6951,N_6736,N_6789);
and U6952 (N_6952,N_6721,N_6606);
xor U6953 (N_6953,N_6661,N_6662);
nor U6954 (N_6954,N_6669,N_6777);
xnor U6955 (N_6955,N_6798,N_6667);
nor U6956 (N_6956,N_6653,N_6688);
nand U6957 (N_6957,N_6661,N_6644);
or U6958 (N_6958,N_6647,N_6658);
nor U6959 (N_6959,N_6623,N_6713);
xnor U6960 (N_6960,N_6632,N_6699);
and U6961 (N_6961,N_6607,N_6757);
nand U6962 (N_6962,N_6657,N_6780);
nor U6963 (N_6963,N_6628,N_6717);
nand U6964 (N_6964,N_6649,N_6771);
or U6965 (N_6965,N_6726,N_6792);
or U6966 (N_6966,N_6709,N_6636);
xnor U6967 (N_6967,N_6773,N_6699);
nand U6968 (N_6968,N_6714,N_6667);
nand U6969 (N_6969,N_6749,N_6764);
xnor U6970 (N_6970,N_6626,N_6633);
nand U6971 (N_6971,N_6663,N_6789);
nand U6972 (N_6972,N_6750,N_6635);
nor U6973 (N_6973,N_6759,N_6630);
nand U6974 (N_6974,N_6722,N_6703);
and U6975 (N_6975,N_6614,N_6634);
and U6976 (N_6976,N_6697,N_6603);
xnor U6977 (N_6977,N_6790,N_6682);
xor U6978 (N_6978,N_6697,N_6751);
and U6979 (N_6979,N_6753,N_6698);
xnor U6980 (N_6980,N_6739,N_6638);
and U6981 (N_6981,N_6770,N_6610);
xor U6982 (N_6982,N_6631,N_6620);
and U6983 (N_6983,N_6758,N_6628);
or U6984 (N_6984,N_6635,N_6798);
nand U6985 (N_6985,N_6687,N_6703);
xnor U6986 (N_6986,N_6683,N_6701);
xor U6987 (N_6987,N_6760,N_6716);
or U6988 (N_6988,N_6752,N_6602);
xor U6989 (N_6989,N_6791,N_6665);
nor U6990 (N_6990,N_6696,N_6648);
and U6991 (N_6991,N_6692,N_6606);
or U6992 (N_6992,N_6739,N_6780);
nand U6993 (N_6993,N_6724,N_6698);
nor U6994 (N_6994,N_6704,N_6722);
or U6995 (N_6995,N_6600,N_6736);
or U6996 (N_6996,N_6617,N_6697);
and U6997 (N_6997,N_6711,N_6710);
nand U6998 (N_6998,N_6746,N_6776);
nand U6999 (N_6999,N_6629,N_6634);
nand U7000 (N_7000,N_6808,N_6855);
and U7001 (N_7001,N_6862,N_6887);
nand U7002 (N_7002,N_6900,N_6915);
and U7003 (N_7003,N_6916,N_6985);
xnor U7004 (N_7004,N_6801,N_6810);
xor U7005 (N_7005,N_6852,N_6920);
or U7006 (N_7006,N_6983,N_6835);
or U7007 (N_7007,N_6807,N_6950);
or U7008 (N_7008,N_6904,N_6940);
nand U7009 (N_7009,N_6890,N_6935);
nor U7010 (N_7010,N_6944,N_6806);
or U7011 (N_7011,N_6824,N_6878);
nand U7012 (N_7012,N_6838,N_6814);
and U7013 (N_7013,N_6948,N_6811);
xor U7014 (N_7014,N_6926,N_6883);
nor U7015 (N_7015,N_6974,N_6831);
and U7016 (N_7016,N_6909,N_6991);
and U7017 (N_7017,N_6975,N_6962);
or U7018 (N_7018,N_6825,N_6861);
or U7019 (N_7019,N_6860,N_6999);
and U7020 (N_7020,N_6871,N_6843);
nor U7021 (N_7021,N_6864,N_6911);
nand U7022 (N_7022,N_6874,N_6973);
nand U7023 (N_7023,N_6943,N_6817);
nand U7024 (N_7024,N_6869,N_6823);
xor U7025 (N_7025,N_6839,N_6936);
nand U7026 (N_7026,N_6967,N_6851);
or U7027 (N_7027,N_6829,N_6856);
and U7028 (N_7028,N_6834,N_6875);
nor U7029 (N_7029,N_6939,N_6894);
xnor U7030 (N_7030,N_6859,N_6832);
nand U7031 (N_7031,N_6917,N_6809);
or U7032 (N_7032,N_6946,N_6921);
and U7033 (N_7033,N_6820,N_6906);
xor U7034 (N_7034,N_6930,N_6961);
and U7035 (N_7035,N_6879,N_6932);
nor U7036 (N_7036,N_6980,N_6964);
nor U7037 (N_7037,N_6903,N_6853);
and U7038 (N_7038,N_6959,N_6866);
xnor U7039 (N_7039,N_6818,N_6901);
nor U7040 (N_7040,N_6858,N_6989);
xnor U7041 (N_7041,N_6847,N_6837);
and U7042 (N_7042,N_6927,N_6951);
xor U7043 (N_7043,N_6919,N_6937);
nor U7044 (N_7044,N_6997,N_6842);
nand U7045 (N_7045,N_6868,N_6992);
and U7046 (N_7046,N_6914,N_6830);
nand U7047 (N_7047,N_6912,N_6925);
nand U7048 (N_7048,N_6895,N_6945);
xor U7049 (N_7049,N_6836,N_6876);
xor U7050 (N_7050,N_6978,N_6918);
xor U7051 (N_7051,N_6970,N_6952);
xnor U7052 (N_7052,N_6899,N_6913);
nor U7053 (N_7053,N_6965,N_6984);
xor U7054 (N_7054,N_6891,N_6947);
and U7055 (N_7055,N_6816,N_6953);
nor U7056 (N_7056,N_6854,N_6888);
nand U7057 (N_7057,N_6885,N_6845);
nor U7058 (N_7058,N_6833,N_6922);
or U7059 (N_7059,N_6907,N_6982);
xor U7060 (N_7060,N_6872,N_6934);
nor U7061 (N_7061,N_6979,N_6955);
and U7062 (N_7062,N_6998,N_6923);
nand U7063 (N_7063,N_6828,N_6902);
xor U7064 (N_7064,N_6928,N_6821);
and U7065 (N_7065,N_6969,N_6849);
or U7066 (N_7066,N_6819,N_6993);
xor U7067 (N_7067,N_6897,N_6933);
or U7068 (N_7068,N_6877,N_6822);
and U7069 (N_7069,N_6898,N_6882);
or U7070 (N_7070,N_6960,N_6813);
xnor U7071 (N_7071,N_6977,N_6886);
nand U7072 (N_7072,N_6880,N_6841);
xor U7073 (N_7073,N_6971,N_6949);
xnor U7074 (N_7074,N_6805,N_6929);
xnor U7075 (N_7075,N_6802,N_6931);
nand U7076 (N_7076,N_6892,N_6867);
nor U7077 (N_7077,N_6924,N_6968);
and U7078 (N_7078,N_6800,N_6910);
xor U7079 (N_7079,N_6994,N_6815);
xor U7080 (N_7080,N_6938,N_6976);
and U7081 (N_7081,N_6996,N_6826);
xnor U7082 (N_7082,N_6956,N_6942);
and U7083 (N_7083,N_6987,N_6840);
or U7084 (N_7084,N_6850,N_6846);
nor U7085 (N_7085,N_6889,N_6908);
and U7086 (N_7086,N_6966,N_6958);
and U7087 (N_7087,N_6865,N_6827);
nand U7088 (N_7088,N_6954,N_6848);
nor U7089 (N_7089,N_6905,N_6995);
and U7090 (N_7090,N_6896,N_6941);
nor U7091 (N_7091,N_6963,N_6870);
and U7092 (N_7092,N_6986,N_6812);
nand U7093 (N_7093,N_6884,N_6972);
xnor U7094 (N_7094,N_6863,N_6803);
xor U7095 (N_7095,N_6804,N_6957);
nand U7096 (N_7096,N_6990,N_6981);
nor U7097 (N_7097,N_6844,N_6881);
nand U7098 (N_7098,N_6988,N_6857);
nor U7099 (N_7099,N_6873,N_6893);
xor U7100 (N_7100,N_6848,N_6845);
xnor U7101 (N_7101,N_6981,N_6991);
and U7102 (N_7102,N_6897,N_6840);
xor U7103 (N_7103,N_6881,N_6858);
nand U7104 (N_7104,N_6802,N_6879);
and U7105 (N_7105,N_6892,N_6829);
or U7106 (N_7106,N_6822,N_6894);
xor U7107 (N_7107,N_6987,N_6951);
or U7108 (N_7108,N_6899,N_6829);
or U7109 (N_7109,N_6921,N_6808);
xnor U7110 (N_7110,N_6922,N_6942);
nor U7111 (N_7111,N_6830,N_6802);
nand U7112 (N_7112,N_6927,N_6806);
and U7113 (N_7113,N_6845,N_6947);
nand U7114 (N_7114,N_6996,N_6922);
nor U7115 (N_7115,N_6891,N_6876);
and U7116 (N_7116,N_6944,N_6971);
or U7117 (N_7117,N_6871,N_6986);
nor U7118 (N_7118,N_6926,N_6877);
nand U7119 (N_7119,N_6964,N_6935);
and U7120 (N_7120,N_6992,N_6901);
and U7121 (N_7121,N_6931,N_6923);
xor U7122 (N_7122,N_6914,N_6854);
nand U7123 (N_7123,N_6896,N_6973);
xnor U7124 (N_7124,N_6837,N_6928);
nor U7125 (N_7125,N_6880,N_6864);
nand U7126 (N_7126,N_6959,N_6801);
and U7127 (N_7127,N_6974,N_6847);
or U7128 (N_7128,N_6904,N_6902);
nand U7129 (N_7129,N_6804,N_6991);
and U7130 (N_7130,N_6928,N_6942);
or U7131 (N_7131,N_6899,N_6953);
or U7132 (N_7132,N_6928,N_6956);
nor U7133 (N_7133,N_6935,N_6877);
or U7134 (N_7134,N_6811,N_6998);
nor U7135 (N_7135,N_6953,N_6922);
nand U7136 (N_7136,N_6850,N_6814);
or U7137 (N_7137,N_6986,N_6846);
and U7138 (N_7138,N_6808,N_6866);
nor U7139 (N_7139,N_6955,N_6931);
nand U7140 (N_7140,N_6885,N_6923);
nor U7141 (N_7141,N_6951,N_6999);
and U7142 (N_7142,N_6972,N_6849);
or U7143 (N_7143,N_6866,N_6941);
or U7144 (N_7144,N_6898,N_6853);
nor U7145 (N_7145,N_6900,N_6972);
or U7146 (N_7146,N_6837,N_6849);
or U7147 (N_7147,N_6898,N_6924);
xnor U7148 (N_7148,N_6871,N_6878);
or U7149 (N_7149,N_6835,N_6865);
xor U7150 (N_7150,N_6885,N_6948);
xor U7151 (N_7151,N_6931,N_6842);
xor U7152 (N_7152,N_6921,N_6993);
or U7153 (N_7153,N_6983,N_6981);
and U7154 (N_7154,N_6889,N_6944);
or U7155 (N_7155,N_6964,N_6936);
or U7156 (N_7156,N_6893,N_6888);
nor U7157 (N_7157,N_6935,N_6829);
or U7158 (N_7158,N_6895,N_6960);
xor U7159 (N_7159,N_6871,N_6902);
or U7160 (N_7160,N_6956,N_6826);
xor U7161 (N_7161,N_6968,N_6865);
or U7162 (N_7162,N_6960,N_6879);
nor U7163 (N_7163,N_6816,N_6846);
nand U7164 (N_7164,N_6956,N_6966);
and U7165 (N_7165,N_6928,N_6957);
and U7166 (N_7166,N_6883,N_6818);
nor U7167 (N_7167,N_6834,N_6872);
or U7168 (N_7168,N_6831,N_6909);
xor U7169 (N_7169,N_6820,N_6844);
nor U7170 (N_7170,N_6975,N_6932);
and U7171 (N_7171,N_6848,N_6859);
or U7172 (N_7172,N_6908,N_6903);
xor U7173 (N_7173,N_6843,N_6887);
nand U7174 (N_7174,N_6939,N_6827);
and U7175 (N_7175,N_6880,N_6995);
nand U7176 (N_7176,N_6827,N_6821);
nor U7177 (N_7177,N_6925,N_6851);
nor U7178 (N_7178,N_6938,N_6885);
or U7179 (N_7179,N_6870,N_6891);
or U7180 (N_7180,N_6830,N_6927);
and U7181 (N_7181,N_6820,N_6955);
xor U7182 (N_7182,N_6880,N_6927);
nor U7183 (N_7183,N_6912,N_6815);
xnor U7184 (N_7184,N_6863,N_6988);
or U7185 (N_7185,N_6819,N_6909);
nor U7186 (N_7186,N_6952,N_6995);
nand U7187 (N_7187,N_6952,N_6837);
or U7188 (N_7188,N_6860,N_6863);
or U7189 (N_7189,N_6850,N_6822);
or U7190 (N_7190,N_6828,N_6953);
nor U7191 (N_7191,N_6993,N_6886);
or U7192 (N_7192,N_6827,N_6914);
and U7193 (N_7193,N_6984,N_6956);
and U7194 (N_7194,N_6880,N_6918);
nor U7195 (N_7195,N_6929,N_6956);
xor U7196 (N_7196,N_6957,N_6812);
nor U7197 (N_7197,N_6882,N_6997);
or U7198 (N_7198,N_6996,N_6885);
xnor U7199 (N_7199,N_6961,N_6866);
xnor U7200 (N_7200,N_7076,N_7184);
nand U7201 (N_7201,N_7099,N_7124);
and U7202 (N_7202,N_7082,N_7090);
nor U7203 (N_7203,N_7079,N_7033);
xnor U7204 (N_7204,N_7046,N_7009);
and U7205 (N_7205,N_7186,N_7064);
xor U7206 (N_7206,N_7161,N_7032);
and U7207 (N_7207,N_7195,N_7061);
xor U7208 (N_7208,N_7140,N_7085);
and U7209 (N_7209,N_7190,N_7163);
nor U7210 (N_7210,N_7146,N_7013);
xor U7211 (N_7211,N_7056,N_7088);
or U7212 (N_7212,N_7156,N_7011);
or U7213 (N_7213,N_7074,N_7096);
nand U7214 (N_7214,N_7168,N_7104);
or U7215 (N_7215,N_7150,N_7160);
nand U7216 (N_7216,N_7182,N_7050);
and U7217 (N_7217,N_7114,N_7149);
and U7218 (N_7218,N_7093,N_7008);
xnor U7219 (N_7219,N_7002,N_7128);
nor U7220 (N_7220,N_7192,N_7087);
or U7221 (N_7221,N_7034,N_7139);
nor U7222 (N_7222,N_7131,N_7118);
or U7223 (N_7223,N_7062,N_7047);
and U7224 (N_7224,N_7059,N_7018);
or U7225 (N_7225,N_7169,N_7045);
and U7226 (N_7226,N_7196,N_7081);
and U7227 (N_7227,N_7148,N_7084);
xnor U7228 (N_7228,N_7103,N_7051);
and U7229 (N_7229,N_7158,N_7028);
nor U7230 (N_7230,N_7198,N_7017);
nand U7231 (N_7231,N_7107,N_7119);
nor U7232 (N_7232,N_7180,N_7029);
nor U7233 (N_7233,N_7170,N_7199);
or U7234 (N_7234,N_7066,N_7166);
or U7235 (N_7235,N_7055,N_7157);
nor U7236 (N_7236,N_7016,N_7007);
nand U7237 (N_7237,N_7134,N_7015);
nand U7238 (N_7238,N_7174,N_7136);
and U7239 (N_7239,N_7181,N_7031);
nand U7240 (N_7240,N_7164,N_7072);
nor U7241 (N_7241,N_7154,N_7135);
and U7242 (N_7242,N_7121,N_7142);
nand U7243 (N_7243,N_7069,N_7075);
and U7244 (N_7244,N_7035,N_7147);
nand U7245 (N_7245,N_7073,N_7126);
nor U7246 (N_7246,N_7165,N_7153);
xor U7247 (N_7247,N_7141,N_7193);
xnor U7248 (N_7248,N_7191,N_7130);
or U7249 (N_7249,N_7178,N_7097);
and U7250 (N_7250,N_7167,N_7098);
or U7251 (N_7251,N_7176,N_7083);
or U7252 (N_7252,N_7110,N_7172);
or U7253 (N_7253,N_7039,N_7127);
xnor U7254 (N_7254,N_7125,N_7122);
or U7255 (N_7255,N_7057,N_7042);
nor U7256 (N_7256,N_7094,N_7113);
nor U7257 (N_7257,N_7111,N_7038);
and U7258 (N_7258,N_7068,N_7185);
nand U7259 (N_7259,N_7189,N_7106);
nor U7260 (N_7260,N_7115,N_7120);
and U7261 (N_7261,N_7112,N_7105);
and U7262 (N_7262,N_7022,N_7040);
xnor U7263 (N_7263,N_7027,N_7137);
and U7264 (N_7264,N_7023,N_7052);
or U7265 (N_7265,N_7151,N_7067);
nor U7266 (N_7266,N_7025,N_7021);
xnor U7267 (N_7267,N_7177,N_7019);
nand U7268 (N_7268,N_7014,N_7162);
and U7269 (N_7269,N_7030,N_7077);
xnor U7270 (N_7270,N_7058,N_7116);
nor U7271 (N_7271,N_7005,N_7036);
xnor U7272 (N_7272,N_7070,N_7003);
nand U7273 (N_7273,N_7092,N_7071);
xnor U7274 (N_7274,N_7100,N_7091);
xnor U7275 (N_7275,N_7173,N_7159);
or U7276 (N_7276,N_7175,N_7026);
or U7277 (N_7277,N_7108,N_7044);
and U7278 (N_7278,N_7152,N_7004);
nand U7279 (N_7279,N_7109,N_7024);
or U7280 (N_7280,N_7138,N_7194);
xnor U7281 (N_7281,N_7183,N_7048);
or U7282 (N_7282,N_7197,N_7123);
xor U7283 (N_7283,N_7133,N_7000);
nor U7284 (N_7284,N_7020,N_7080);
or U7285 (N_7285,N_7012,N_7006);
nand U7286 (N_7286,N_7155,N_7132);
xor U7287 (N_7287,N_7102,N_7188);
and U7288 (N_7288,N_7187,N_7037);
and U7289 (N_7289,N_7065,N_7145);
nand U7290 (N_7290,N_7063,N_7060);
or U7291 (N_7291,N_7001,N_7095);
or U7292 (N_7292,N_7179,N_7053);
and U7293 (N_7293,N_7171,N_7129);
nand U7294 (N_7294,N_7101,N_7089);
or U7295 (N_7295,N_7010,N_7143);
and U7296 (N_7296,N_7117,N_7041);
xnor U7297 (N_7297,N_7049,N_7043);
xnor U7298 (N_7298,N_7054,N_7144);
nand U7299 (N_7299,N_7078,N_7086);
nand U7300 (N_7300,N_7030,N_7047);
and U7301 (N_7301,N_7001,N_7048);
and U7302 (N_7302,N_7056,N_7136);
or U7303 (N_7303,N_7011,N_7105);
xor U7304 (N_7304,N_7112,N_7126);
xor U7305 (N_7305,N_7051,N_7157);
xnor U7306 (N_7306,N_7176,N_7195);
or U7307 (N_7307,N_7012,N_7162);
xnor U7308 (N_7308,N_7117,N_7015);
xnor U7309 (N_7309,N_7125,N_7140);
or U7310 (N_7310,N_7168,N_7150);
nor U7311 (N_7311,N_7198,N_7188);
nand U7312 (N_7312,N_7149,N_7003);
and U7313 (N_7313,N_7058,N_7086);
and U7314 (N_7314,N_7145,N_7134);
and U7315 (N_7315,N_7046,N_7010);
nor U7316 (N_7316,N_7190,N_7146);
nand U7317 (N_7317,N_7196,N_7186);
nor U7318 (N_7318,N_7144,N_7035);
or U7319 (N_7319,N_7161,N_7010);
xnor U7320 (N_7320,N_7118,N_7034);
nor U7321 (N_7321,N_7023,N_7105);
or U7322 (N_7322,N_7104,N_7144);
xor U7323 (N_7323,N_7051,N_7030);
nor U7324 (N_7324,N_7016,N_7097);
nand U7325 (N_7325,N_7051,N_7115);
nand U7326 (N_7326,N_7000,N_7013);
or U7327 (N_7327,N_7146,N_7108);
and U7328 (N_7328,N_7059,N_7101);
xnor U7329 (N_7329,N_7073,N_7046);
nor U7330 (N_7330,N_7187,N_7197);
xor U7331 (N_7331,N_7005,N_7100);
or U7332 (N_7332,N_7038,N_7071);
nand U7333 (N_7333,N_7029,N_7114);
nor U7334 (N_7334,N_7102,N_7185);
and U7335 (N_7335,N_7199,N_7109);
xnor U7336 (N_7336,N_7108,N_7007);
xnor U7337 (N_7337,N_7122,N_7050);
and U7338 (N_7338,N_7081,N_7029);
nor U7339 (N_7339,N_7128,N_7144);
and U7340 (N_7340,N_7108,N_7028);
nor U7341 (N_7341,N_7010,N_7196);
and U7342 (N_7342,N_7025,N_7028);
nor U7343 (N_7343,N_7087,N_7096);
xnor U7344 (N_7344,N_7054,N_7146);
nand U7345 (N_7345,N_7195,N_7107);
or U7346 (N_7346,N_7096,N_7080);
nand U7347 (N_7347,N_7150,N_7142);
and U7348 (N_7348,N_7184,N_7118);
nor U7349 (N_7349,N_7165,N_7084);
and U7350 (N_7350,N_7092,N_7125);
nand U7351 (N_7351,N_7009,N_7110);
nand U7352 (N_7352,N_7167,N_7146);
and U7353 (N_7353,N_7119,N_7019);
or U7354 (N_7354,N_7104,N_7109);
and U7355 (N_7355,N_7000,N_7171);
xor U7356 (N_7356,N_7112,N_7005);
xor U7357 (N_7357,N_7077,N_7031);
and U7358 (N_7358,N_7163,N_7161);
nand U7359 (N_7359,N_7146,N_7041);
nor U7360 (N_7360,N_7020,N_7151);
or U7361 (N_7361,N_7058,N_7024);
or U7362 (N_7362,N_7075,N_7032);
and U7363 (N_7363,N_7041,N_7053);
nand U7364 (N_7364,N_7009,N_7192);
xnor U7365 (N_7365,N_7027,N_7131);
or U7366 (N_7366,N_7033,N_7153);
or U7367 (N_7367,N_7000,N_7050);
or U7368 (N_7368,N_7107,N_7095);
nand U7369 (N_7369,N_7162,N_7114);
or U7370 (N_7370,N_7100,N_7120);
nand U7371 (N_7371,N_7022,N_7052);
xnor U7372 (N_7372,N_7137,N_7031);
nor U7373 (N_7373,N_7030,N_7137);
or U7374 (N_7374,N_7045,N_7148);
nor U7375 (N_7375,N_7124,N_7014);
or U7376 (N_7376,N_7160,N_7019);
nor U7377 (N_7377,N_7061,N_7039);
and U7378 (N_7378,N_7194,N_7000);
and U7379 (N_7379,N_7138,N_7002);
nand U7380 (N_7380,N_7191,N_7152);
and U7381 (N_7381,N_7048,N_7160);
nand U7382 (N_7382,N_7087,N_7005);
or U7383 (N_7383,N_7146,N_7086);
nor U7384 (N_7384,N_7142,N_7047);
nor U7385 (N_7385,N_7198,N_7163);
xor U7386 (N_7386,N_7098,N_7102);
nor U7387 (N_7387,N_7033,N_7057);
or U7388 (N_7388,N_7024,N_7098);
nor U7389 (N_7389,N_7056,N_7181);
xnor U7390 (N_7390,N_7121,N_7005);
xnor U7391 (N_7391,N_7046,N_7126);
and U7392 (N_7392,N_7082,N_7091);
nand U7393 (N_7393,N_7142,N_7077);
nand U7394 (N_7394,N_7104,N_7110);
nand U7395 (N_7395,N_7194,N_7175);
and U7396 (N_7396,N_7047,N_7165);
nand U7397 (N_7397,N_7139,N_7112);
nand U7398 (N_7398,N_7053,N_7100);
and U7399 (N_7399,N_7038,N_7164);
and U7400 (N_7400,N_7247,N_7227);
xor U7401 (N_7401,N_7342,N_7258);
or U7402 (N_7402,N_7210,N_7351);
xnor U7403 (N_7403,N_7330,N_7283);
xor U7404 (N_7404,N_7314,N_7349);
xnor U7405 (N_7405,N_7339,N_7297);
or U7406 (N_7406,N_7315,N_7320);
nor U7407 (N_7407,N_7251,N_7368);
nand U7408 (N_7408,N_7213,N_7359);
or U7409 (N_7409,N_7310,N_7252);
nand U7410 (N_7410,N_7305,N_7375);
and U7411 (N_7411,N_7290,N_7353);
nor U7412 (N_7412,N_7214,N_7201);
nor U7413 (N_7413,N_7321,N_7222);
nand U7414 (N_7414,N_7340,N_7396);
or U7415 (N_7415,N_7218,N_7240);
xor U7416 (N_7416,N_7219,N_7386);
or U7417 (N_7417,N_7387,N_7331);
nand U7418 (N_7418,N_7298,N_7385);
nor U7419 (N_7419,N_7301,N_7394);
nor U7420 (N_7420,N_7371,N_7278);
nor U7421 (N_7421,N_7206,N_7395);
nand U7422 (N_7422,N_7273,N_7265);
nor U7423 (N_7423,N_7398,N_7236);
and U7424 (N_7424,N_7391,N_7355);
nand U7425 (N_7425,N_7317,N_7257);
nor U7426 (N_7426,N_7309,N_7380);
and U7427 (N_7427,N_7281,N_7350);
xor U7428 (N_7428,N_7231,N_7284);
xnor U7429 (N_7429,N_7261,N_7361);
or U7430 (N_7430,N_7303,N_7296);
xnor U7431 (N_7431,N_7319,N_7279);
nand U7432 (N_7432,N_7239,N_7203);
xnor U7433 (N_7433,N_7260,N_7332);
and U7434 (N_7434,N_7366,N_7267);
nor U7435 (N_7435,N_7243,N_7277);
nor U7436 (N_7436,N_7338,N_7250);
xor U7437 (N_7437,N_7274,N_7217);
xnor U7438 (N_7438,N_7244,N_7376);
or U7439 (N_7439,N_7256,N_7208);
or U7440 (N_7440,N_7364,N_7367);
and U7441 (N_7441,N_7271,N_7343);
nor U7442 (N_7442,N_7381,N_7226);
or U7443 (N_7443,N_7334,N_7245);
xnor U7444 (N_7444,N_7288,N_7254);
xor U7445 (N_7445,N_7242,N_7299);
or U7446 (N_7446,N_7204,N_7282);
xnor U7447 (N_7447,N_7392,N_7223);
nand U7448 (N_7448,N_7289,N_7313);
xnor U7449 (N_7449,N_7293,N_7358);
and U7450 (N_7450,N_7360,N_7246);
xor U7451 (N_7451,N_7200,N_7229);
or U7452 (N_7452,N_7341,N_7354);
nand U7453 (N_7453,N_7312,N_7294);
nand U7454 (N_7454,N_7324,N_7225);
nand U7455 (N_7455,N_7233,N_7378);
and U7456 (N_7456,N_7291,N_7221);
nand U7457 (N_7457,N_7234,N_7295);
nor U7458 (N_7458,N_7308,N_7325);
and U7459 (N_7459,N_7264,N_7307);
nor U7460 (N_7460,N_7232,N_7302);
nand U7461 (N_7461,N_7263,N_7292);
nor U7462 (N_7462,N_7382,N_7357);
nor U7463 (N_7463,N_7270,N_7345);
nor U7464 (N_7464,N_7397,N_7370);
or U7465 (N_7465,N_7209,N_7369);
nand U7466 (N_7466,N_7272,N_7215);
nand U7467 (N_7467,N_7248,N_7390);
nand U7468 (N_7468,N_7336,N_7379);
nor U7469 (N_7469,N_7318,N_7399);
nand U7470 (N_7470,N_7322,N_7304);
nor U7471 (N_7471,N_7216,N_7326);
nand U7472 (N_7472,N_7306,N_7280);
and U7473 (N_7473,N_7202,N_7333);
xor U7474 (N_7474,N_7346,N_7327);
and U7475 (N_7475,N_7275,N_7228);
and U7476 (N_7476,N_7235,N_7316);
or U7477 (N_7477,N_7205,N_7347);
nor U7478 (N_7478,N_7286,N_7328);
nand U7479 (N_7479,N_7363,N_7335);
nand U7480 (N_7480,N_7384,N_7323);
or U7481 (N_7481,N_7212,N_7269);
nor U7482 (N_7482,N_7262,N_7276);
nand U7483 (N_7483,N_7300,N_7237);
xnor U7484 (N_7484,N_7207,N_7388);
xnor U7485 (N_7485,N_7372,N_7337);
and U7486 (N_7486,N_7224,N_7344);
or U7487 (N_7487,N_7389,N_7352);
or U7488 (N_7488,N_7362,N_7285);
xnor U7489 (N_7489,N_7238,N_7241);
nor U7490 (N_7490,N_7393,N_7377);
or U7491 (N_7491,N_7253,N_7348);
xor U7492 (N_7492,N_7249,N_7220);
nor U7493 (N_7493,N_7329,N_7287);
nand U7494 (N_7494,N_7356,N_7311);
and U7495 (N_7495,N_7266,N_7255);
nand U7496 (N_7496,N_7374,N_7259);
or U7497 (N_7497,N_7373,N_7383);
or U7498 (N_7498,N_7230,N_7211);
nand U7499 (N_7499,N_7268,N_7365);
nand U7500 (N_7500,N_7398,N_7354);
nand U7501 (N_7501,N_7260,N_7209);
nor U7502 (N_7502,N_7349,N_7382);
and U7503 (N_7503,N_7294,N_7365);
nor U7504 (N_7504,N_7344,N_7201);
xor U7505 (N_7505,N_7273,N_7309);
nand U7506 (N_7506,N_7390,N_7249);
nor U7507 (N_7507,N_7351,N_7231);
xnor U7508 (N_7508,N_7341,N_7295);
xnor U7509 (N_7509,N_7358,N_7349);
xor U7510 (N_7510,N_7235,N_7346);
xnor U7511 (N_7511,N_7253,N_7381);
nor U7512 (N_7512,N_7217,N_7201);
or U7513 (N_7513,N_7287,N_7333);
nand U7514 (N_7514,N_7382,N_7337);
or U7515 (N_7515,N_7234,N_7300);
and U7516 (N_7516,N_7227,N_7374);
xor U7517 (N_7517,N_7338,N_7322);
nand U7518 (N_7518,N_7230,N_7269);
and U7519 (N_7519,N_7215,N_7251);
nor U7520 (N_7520,N_7345,N_7369);
nor U7521 (N_7521,N_7208,N_7242);
nand U7522 (N_7522,N_7398,N_7355);
nand U7523 (N_7523,N_7274,N_7218);
xnor U7524 (N_7524,N_7332,N_7279);
xor U7525 (N_7525,N_7242,N_7228);
nor U7526 (N_7526,N_7216,N_7377);
or U7527 (N_7527,N_7208,N_7255);
or U7528 (N_7528,N_7241,N_7242);
and U7529 (N_7529,N_7335,N_7251);
nor U7530 (N_7530,N_7371,N_7340);
and U7531 (N_7531,N_7226,N_7216);
nand U7532 (N_7532,N_7267,N_7347);
or U7533 (N_7533,N_7334,N_7338);
and U7534 (N_7534,N_7382,N_7363);
xnor U7535 (N_7535,N_7381,N_7272);
nor U7536 (N_7536,N_7319,N_7354);
and U7537 (N_7537,N_7300,N_7326);
nand U7538 (N_7538,N_7270,N_7370);
xor U7539 (N_7539,N_7282,N_7243);
nand U7540 (N_7540,N_7398,N_7293);
nor U7541 (N_7541,N_7297,N_7344);
xnor U7542 (N_7542,N_7244,N_7363);
or U7543 (N_7543,N_7343,N_7275);
or U7544 (N_7544,N_7282,N_7285);
nor U7545 (N_7545,N_7320,N_7229);
nand U7546 (N_7546,N_7213,N_7217);
or U7547 (N_7547,N_7397,N_7378);
nand U7548 (N_7548,N_7337,N_7218);
and U7549 (N_7549,N_7366,N_7207);
nand U7550 (N_7550,N_7393,N_7212);
and U7551 (N_7551,N_7315,N_7274);
nor U7552 (N_7552,N_7291,N_7392);
or U7553 (N_7553,N_7207,N_7365);
or U7554 (N_7554,N_7341,N_7361);
and U7555 (N_7555,N_7218,N_7313);
and U7556 (N_7556,N_7251,N_7210);
nand U7557 (N_7557,N_7261,N_7293);
nor U7558 (N_7558,N_7310,N_7309);
and U7559 (N_7559,N_7300,N_7390);
or U7560 (N_7560,N_7356,N_7226);
xor U7561 (N_7561,N_7248,N_7371);
or U7562 (N_7562,N_7329,N_7341);
nor U7563 (N_7563,N_7317,N_7378);
nor U7564 (N_7564,N_7224,N_7314);
and U7565 (N_7565,N_7309,N_7370);
nand U7566 (N_7566,N_7269,N_7372);
and U7567 (N_7567,N_7273,N_7307);
nand U7568 (N_7568,N_7220,N_7386);
nand U7569 (N_7569,N_7363,N_7259);
or U7570 (N_7570,N_7297,N_7211);
or U7571 (N_7571,N_7271,N_7296);
xor U7572 (N_7572,N_7268,N_7252);
xnor U7573 (N_7573,N_7234,N_7337);
or U7574 (N_7574,N_7349,N_7345);
nor U7575 (N_7575,N_7358,N_7394);
and U7576 (N_7576,N_7357,N_7325);
xnor U7577 (N_7577,N_7319,N_7263);
nor U7578 (N_7578,N_7207,N_7262);
and U7579 (N_7579,N_7308,N_7374);
and U7580 (N_7580,N_7345,N_7207);
xor U7581 (N_7581,N_7247,N_7256);
and U7582 (N_7582,N_7201,N_7334);
nand U7583 (N_7583,N_7262,N_7329);
and U7584 (N_7584,N_7272,N_7366);
or U7585 (N_7585,N_7383,N_7228);
nand U7586 (N_7586,N_7290,N_7304);
xnor U7587 (N_7587,N_7322,N_7283);
nor U7588 (N_7588,N_7363,N_7209);
and U7589 (N_7589,N_7367,N_7282);
nand U7590 (N_7590,N_7367,N_7270);
xnor U7591 (N_7591,N_7296,N_7254);
xor U7592 (N_7592,N_7273,N_7378);
xnor U7593 (N_7593,N_7320,N_7331);
nand U7594 (N_7594,N_7349,N_7377);
and U7595 (N_7595,N_7219,N_7294);
xor U7596 (N_7596,N_7259,N_7212);
and U7597 (N_7597,N_7314,N_7218);
nand U7598 (N_7598,N_7386,N_7303);
and U7599 (N_7599,N_7304,N_7399);
xnor U7600 (N_7600,N_7551,N_7537);
nor U7601 (N_7601,N_7594,N_7575);
and U7602 (N_7602,N_7426,N_7564);
or U7603 (N_7603,N_7457,N_7417);
nand U7604 (N_7604,N_7413,N_7508);
xnor U7605 (N_7605,N_7574,N_7448);
and U7606 (N_7606,N_7556,N_7506);
nor U7607 (N_7607,N_7495,N_7431);
nor U7608 (N_7608,N_7521,N_7467);
or U7609 (N_7609,N_7509,N_7470);
and U7610 (N_7610,N_7445,N_7582);
nand U7611 (N_7611,N_7450,N_7485);
or U7612 (N_7612,N_7444,N_7419);
xor U7613 (N_7613,N_7486,N_7539);
nor U7614 (N_7614,N_7436,N_7500);
nor U7615 (N_7615,N_7472,N_7475);
nor U7616 (N_7616,N_7547,N_7473);
or U7617 (N_7617,N_7573,N_7523);
or U7618 (N_7618,N_7548,N_7498);
xor U7619 (N_7619,N_7410,N_7449);
or U7620 (N_7620,N_7528,N_7578);
or U7621 (N_7621,N_7412,N_7598);
nand U7622 (N_7622,N_7595,N_7593);
xnor U7623 (N_7623,N_7532,N_7512);
and U7624 (N_7624,N_7519,N_7502);
nand U7625 (N_7625,N_7568,N_7458);
xor U7626 (N_7626,N_7554,N_7433);
or U7627 (N_7627,N_7443,N_7538);
nand U7628 (N_7628,N_7442,N_7405);
and U7629 (N_7629,N_7513,N_7488);
xor U7630 (N_7630,N_7460,N_7526);
nand U7631 (N_7631,N_7453,N_7507);
xnor U7632 (N_7632,N_7452,N_7558);
nand U7633 (N_7633,N_7557,N_7477);
and U7634 (N_7634,N_7424,N_7409);
or U7635 (N_7635,N_7536,N_7591);
nand U7636 (N_7636,N_7516,N_7446);
and U7637 (N_7637,N_7461,N_7511);
and U7638 (N_7638,N_7561,N_7441);
xnor U7639 (N_7639,N_7514,N_7510);
or U7640 (N_7640,N_7503,N_7476);
xnor U7641 (N_7641,N_7418,N_7560);
nand U7642 (N_7642,N_7541,N_7530);
nand U7643 (N_7643,N_7543,N_7484);
and U7644 (N_7644,N_7435,N_7430);
xnor U7645 (N_7645,N_7469,N_7553);
nor U7646 (N_7646,N_7403,N_7583);
and U7647 (N_7647,N_7524,N_7559);
and U7648 (N_7648,N_7459,N_7563);
nor U7649 (N_7649,N_7534,N_7479);
or U7650 (N_7650,N_7599,N_7487);
or U7651 (N_7651,N_7581,N_7542);
or U7652 (N_7652,N_7566,N_7439);
or U7653 (N_7653,N_7569,N_7429);
nor U7654 (N_7654,N_7520,N_7579);
or U7655 (N_7655,N_7465,N_7555);
or U7656 (N_7656,N_7466,N_7474);
and U7657 (N_7657,N_7404,N_7496);
and U7658 (N_7658,N_7590,N_7489);
and U7659 (N_7659,N_7483,N_7428);
nand U7660 (N_7660,N_7592,N_7464);
or U7661 (N_7661,N_7468,N_7411);
xnor U7662 (N_7662,N_7501,N_7425);
or U7663 (N_7663,N_7490,N_7401);
nor U7664 (N_7664,N_7423,N_7420);
and U7665 (N_7665,N_7492,N_7427);
and U7666 (N_7666,N_7584,N_7505);
and U7667 (N_7667,N_7545,N_7462);
nand U7668 (N_7668,N_7565,N_7454);
nor U7669 (N_7669,N_7432,N_7549);
nand U7670 (N_7670,N_7589,N_7572);
or U7671 (N_7671,N_7463,N_7451);
nor U7672 (N_7672,N_7525,N_7407);
nand U7673 (N_7673,N_7531,N_7434);
nand U7674 (N_7674,N_7540,N_7517);
and U7675 (N_7675,N_7518,N_7567);
or U7676 (N_7676,N_7535,N_7406);
xor U7677 (N_7677,N_7408,N_7447);
or U7678 (N_7678,N_7552,N_7493);
xor U7679 (N_7679,N_7456,N_7497);
xor U7680 (N_7680,N_7546,N_7587);
nand U7681 (N_7681,N_7416,N_7533);
and U7682 (N_7682,N_7402,N_7491);
nand U7683 (N_7683,N_7596,N_7544);
or U7684 (N_7684,N_7422,N_7415);
and U7685 (N_7685,N_7597,N_7571);
nand U7686 (N_7686,N_7585,N_7440);
and U7687 (N_7687,N_7515,N_7400);
nand U7688 (N_7688,N_7421,N_7414);
and U7689 (N_7689,N_7494,N_7580);
or U7690 (N_7690,N_7576,N_7455);
and U7691 (N_7691,N_7577,N_7438);
or U7692 (N_7692,N_7478,N_7562);
or U7693 (N_7693,N_7527,N_7482);
and U7694 (N_7694,N_7437,N_7570);
or U7695 (N_7695,N_7588,N_7586);
nand U7696 (N_7696,N_7499,N_7529);
xor U7697 (N_7697,N_7471,N_7522);
xor U7698 (N_7698,N_7504,N_7550);
or U7699 (N_7699,N_7481,N_7480);
or U7700 (N_7700,N_7572,N_7421);
or U7701 (N_7701,N_7545,N_7490);
nand U7702 (N_7702,N_7576,N_7425);
xor U7703 (N_7703,N_7543,N_7512);
or U7704 (N_7704,N_7465,N_7422);
or U7705 (N_7705,N_7575,N_7507);
nor U7706 (N_7706,N_7421,N_7558);
and U7707 (N_7707,N_7427,N_7490);
nand U7708 (N_7708,N_7498,N_7507);
or U7709 (N_7709,N_7582,N_7578);
nand U7710 (N_7710,N_7433,N_7480);
nand U7711 (N_7711,N_7418,N_7477);
nor U7712 (N_7712,N_7572,N_7567);
xor U7713 (N_7713,N_7549,N_7585);
nand U7714 (N_7714,N_7528,N_7593);
and U7715 (N_7715,N_7400,N_7411);
nor U7716 (N_7716,N_7487,N_7549);
nand U7717 (N_7717,N_7526,N_7415);
nand U7718 (N_7718,N_7466,N_7568);
nor U7719 (N_7719,N_7592,N_7576);
nor U7720 (N_7720,N_7545,N_7442);
and U7721 (N_7721,N_7551,N_7593);
nand U7722 (N_7722,N_7597,N_7577);
or U7723 (N_7723,N_7493,N_7463);
nor U7724 (N_7724,N_7510,N_7409);
or U7725 (N_7725,N_7422,N_7519);
nor U7726 (N_7726,N_7465,N_7570);
and U7727 (N_7727,N_7551,N_7428);
xor U7728 (N_7728,N_7521,N_7417);
or U7729 (N_7729,N_7553,N_7439);
xnor U7730 (N_7730,N_7457,N_7588);
xnor U7731 (N_7731,N_7403,N_7456);
and U7732 (N_7732,N_7454,N_7529);
or U7733 (N_7733,N_7532,N_7480);
and U7734 (N_7734,N_7466,N_7436);
nand U7735 (N_7735,N_7564,N_7505);
or U7736 (N_7736,N_7590,N_7436);
or U7737 (N_7737,N_7495,N_7594);
or U7738 (N_7738,N_7579,N_7435);
nor U7739 (N_7739,N_7573,N_7469);
nor U7740 (N_7740,N_7477,N_7552);
nor U7741 (N_7741,N_7430,N_7537);
xnor U7742 (N_7742,N_7520,N_7486);
nor U7743 (N_7743,N_7567,N_7504);
nor U7744 (N_7744,N_7587,N_7599);
xnor U7745 (N_7745,N_7579,N_7400);
and U7746 (N_7746,N_7469,N_7406);
or U7747 (N_7747,N_7474,N_7403);
nor U7748 (N_7748,N_7528,N_7494);
or U7749 (N_7749,N_7489,N_7528);
xor U7750 (N_7750,N_7413,N_7406);
xnor U7751 (N_7751,N_7519,N_7484);
nor U7752 (N_7752,N_7567,N_7441);
xor U7753 (N_7753,N_7584,N_7508);
nor U7754 (N_7754,N_7519,N_7577);
nand U7755 (N_7755,N_7468,N_7572);
and U7756 (N_7756,N_7533,N_7419);
xor U7757 (N_7757,N_7528,N_7539);
xnor U7758 (N_7758,N_7471,N_7441);
and U7759 (N_7759,N_7409,N_7573);
xor U7760 (N_7760,N_7463,N_7465);
nor U7761 (N_7761,N_7529,N_7543);
and U7762 (N_7762,N_7581,N_7404);
nor U7763 (N_7763,N_7436,N_7423);
xnor U7764 (N_7764,N_7542,N_7474);
or U7765 (N_7765,N_7444,N_7410);
or U7766 (N_7766,N_7487,N_7581);
nand U7767 (N_7767,N_7523,N_7436);
xnor U7768 (N_7768,N_7536,N_7483);
or U7769 (N_7769,N_7595,N_7493);
and U7770 (N_7770,N_7505,N_7592);
or U7771 (N_7771,N_7402,N_7435);
or U7772 (N_7772,N_7548,N_7440);
xnor U7773 (N_7773,N_7490,N_7549);
nor U7774 (N_7774,N_7450,N_7506);
nor U7775 (N_7775,N_7442,N_7563);
nor U7776 (N_7776,N_7477,N_7440);
xor U7777 (N_7777,N_7403,N_7475);
or U7778 (N_7778,N_7576,N_7538);
nand U7779 (N_7779,N_7555,N_7422);
nand U7780 (N_7780,N_7592,N_7591);
nor U7781 (N_7781,N_7410,N_7564);
nor U7782 (N_7782,N_7513,N_7568);
nand U7783 (N_7783,N_7477,N_7423);
xnor U7784 (N_7784,N_7421,N_7509);
nor U7785 (N_7785,N_7565,N_7508);
nor U7786 (N_7786,N_7585,N_7569);
xnor U7787 (N_7787,N_7463,N_7551);
nand U7788 (N_7788,N_7590,N_7484);
xor U7789 (N_7789,N_7454,N_7525);
or U7790 (N_7790,N_7513,N_7539);
xor U7791 (N_7791,N_7586,N_7403);
nand U7792 (N_7792,N_7451,N_7461);
nor U7793 (N_7793,N_7569,N_7479);
or U7794 (N_7794,N_7467,N_7595);
and U7795 (N_7795,N_7500,N_7598);
nor U7796 (N_7796,N_7581,N_7529);
xor U7797 (N_7797,N_7514,N_7519);
xnor U7798 (N_7798,N_7430,N_7509);
and U7799 (N_7799,N_7481,N_7584);
nand U7800 (N_7800,N_7717,N_7601);
xor U7801 (N_7801,N_7622,N_7626);
xnor U7802 (N_7802,N_7708,N_7731);
nor U7803 (N_7803,N_7666,N_7652);
xor U7804 (N_7804,N_7640,N_7675);
nor U7805 (N_7805,N_7605,N_7781);
and U7806 (N_7806,N_7662,N_7677);
and U7807 (N_7807,N_7710,N_7639);
nand U7808 (N_7808,N_7686,N_7676);
nor U7809 (N_7809,N_7793,N_7608);
and U7810 (N_7810,N_7768,N_7611);
nand U7811 (N_7811,N_7619,N_7769);
nor U7812 (N_7812,N_7607,N_7715);
and U7813 (N_7813,N_7689,N_7798);
and U7814 (N_7814,N_7737,N_7694);
and U7815 (N_7815,N_7774,N_7760);
nor U7816 (N_7816,N_7748,N_7782);
nand U7817 (N_7817,N_7645,N_7751);
or U7818 (N_7818,N_7763,N_7623);
nor U7819 (N_7819,N_7691,N_7706);
or U7820 (N_7820,N_7722,N_7704);
xor U7821 (N_7821,N_7682,N_7721);
and U7822 (N_7822,N_7628,N_7606);
or U7823 (N_7823,N_7655,N_7674);
and U7824 (N_7824,N_7787,N_7610);
xor U7825 (N_7825,N_7600,N_7612);
nand U7826 (N_7826,N_7716,N_7744);
or U7827 (N_7827,N_7685,N_7777);
and U7828 (N_7828,N_7669,N_7688);
and U7829 (N_7829,N_7651,N_7732);
or U7830 (N_7830,N_7735,N_7758);
xnor U7831 (N_7831,N_7698,N_7630);
and U7832 (N_7832,N_7711,N_7753);
and U7833 (N_7833,N_7773,N_7673);
xnor U7834 (N_7834,N_7743,N_7799);
xnor U7835 (N_7835,N_7778,N_7775);
and U7836 (N_7836,N_7684,N_7700);
xor U7837 (N_7837,N_7614,N_7667);
xnor U7838 (N_7838,N_7767,N_7747);
nor U7839 (N_7839,N_7720,N_7620);
nor U7840 (N_7840,N_7795,N_7770);
nand U7841 (N_7841,N_7784,N_7702);
and U7842 (N_7842,N_7757,N_7602);
nand U7843 (N_7843,N_7734,N_7738);
or U7844 (N_7844,N_7796,N_7638);
nand U7845 (N_7845,N_7692,N_7794);
xor U7846 (N_7846,N_7671,N_7730);
or U7847 (N_7847,N_7739,N_7797);
or U7848 (N_7848,N_7723,N_7643);
xor U7849 (N_7849,N_7785,N_7615);
xnor U7850 (N_7850,N_7786,N_7665);
nor U7851 (N_7851,N_7648,N_7696);
nand U7852 (N_7852,N_7650,N_7742);
or U7853 (N_7853,N_7637,N_7772);
nand U7854 (N_7854,N_7727,N_7729);
and U7855 (N_7855,N_7765,N_7707);
or U7856 (N_7856,N_7679,N_7693);
or U7857 (N_7857,N_7646,N_7695);
xnor U7858 (N_7858,N_7624,N_7701);
or U7859 (N_7859,N_7613,N_7604);
nand U7860 (N_7860,N_7766,N_7644);
or U7861 (N_7861,N_7641,N_7703);
and U7862 (N_7862,N_7746,N_7776);
xor U7863 (N_7863,N_7661,N_7647);
nand U7864 (N_7864,N_7736,N_7752);
nor U7865 (N_7865,N_7713,N_7690);
nand U7866 (N_7866,N_7792,N_7714);
nand U7867 (N_7867,N_7719,N_7663);
or U7868 (N_7868,N_7718,N_7625);
and U7869 (N_7869,N_7632,N_7764);
nor U7870 (N_7870,N_7779,N_7726);
nand U7871 (N_7871,N_7780,N_7697);
xnor U7872 (N_7872,N_7633,N_7728);
xnor U7873 (N_7873,N_7683,N_7627);
or U7874 (N_7874,N_7788,N_7634);
and U7875 (N_7875,N_7660,N_7759);
xor U7876 (N_7876,N_7664,N_7653);
and U7877 (N_7877,N_7712,N_7745);
nor U7878 (N_7878,N_7678,N_7670);
or U7879 (N_7879,N_7649,N_7672);
or U7880 (N_7880,N_7790,N_7617);
nand U7881 (N_7881,N_7635,N_7629);
xnor U7882 (N_7882,N_7699,N_7783);
xor U7883 (N_7883,N_7705,N_7750);
or U7884 (N_7884,N_7754,N_7618);
and U7885 (N_7885,N_7636,N_7642);
xor U7886 (N_7886,N_7733,N_7621);
nand U7887 (N_7887,N_7791,N_7725);
and U7888 (N_7888,N_7755,N_7609);
and U7889 (N_7889,N_7656,N_7709);
nand U7890 (N_7890,N_7741,N_7681);
nand U7891 (N_7891,N_7616,N_7756);
and U7892 (N_7892,N_7724,N_7740);
nor U7893 (N_7893,N_7658,N_7659);
nand U7894 (N_7894,N_7749,N_7762);
nor U7895 (N_7895,N_7761,N_7654);
nor U7896 (N_7896,N_7771,N_7631);
xnor U7897 (N_7897,N_7603,N_7668);
xnor U7898 (N_7898,N_7789,N_7680);
nand U7899 (N_7899,N_7657,N_7687);
nand U7900 (N_7900,N_7621,N_7717);
and U7901 (N_7901,N_7647,N_7618);
xor U7902 (N_7902,N_7711,N_7658);
nor U7903 (N_7903,N_7790,N_7750);
nand U7904 (N_7904,N_7741,N_7604);
xnor U7905 (N_7905,N_7727,N_7602);
and U7906 (N_7906,N_7691,N_7620);
nor U7907 (N_7907,N_7750,N_7726);
nor U7908 (N_7908,N_7755,N_7727);
and U7909 (N_7909,N_7710,N_7788);
xor U7910 (N_7910,N_7641,N_7785);
or U7911 (N_7911,N_7629,N_7670);
or U7912 (N_7912,N_7611,N_7799);
and U7913 (N_7913,N_7702,N_7751);
nand U7914 (N_7914,N_7702,N_7661);
nor U7915 (N_7915,N_7601,N_7710);
and U7916 (N_7916,N_7735,N_7660);
or U7917 (N_7917,N_7633,N_7643);
nand U7918 (N_7918,N_7609,N_7733);
nand U7919 (N_7919,N_7754,N_7753);
or U7920 (N_7920,N_7619,N_7712);
and U7921 (N_7921,N_7673,N_7663);
nor U7922 (N_7922,N_7634,N_7670);
xnor U7923 (N_7923,N_7790,N_7736);
xnor U7924 (N_7924,N_7630,N_7794);
nor U7925 (N_7925,N_7757,N_7704);
or U7926 (N_7926,N_7660,N_7797);
nor U7927 (N_7927,N_7717,N_7668);
nand U7928 (N_7928,N_7789,N_7797);
or U7929 (N_7929,N_7678,N_7748);
xnor U7930 (N_7930,N_7694,N_7791);
xor U7931 (N_7931,N_7627,N_7616);
nor U7932 (N_7932,N_7774,N_7651);
xnor U7933 (N_7933,N_7783,N_7690);
nand U7934 (N_7934,N_7746,N_7706);
xor U7935 (N_7935,N_7790,N_7698);
or U7936 (N_7936,N_7662,N_7621);
or U7937 (N_7937,N_7655,N_7704);
or U7938 (N_7938,N_7721,N_7720);
nand U7939 (N_7939,N_7600,N_7722);
or U7940 (N_7940,N_7614,N_7749);
and U7941 (N_7941,N_7674,N_7694);
or U7942 (N_7942,N_7706,N_7743);
or U7943 (N_7943,N_7654,N_7643);
nand U7944 (N_7944,N_7750,N_7696);
or U7945 (N_7945,N_7702,N_7725);
nor U7946 (N_7946,N_7760,N_7792);
xnor U7947 (N_7947,N_7687,N_7764);
nand U7948 (N_7948,N_7730,N_7728);
nand U7949 (N_7949,N_7638,N_7651);
xor U7950 (N_7950,N_7703,N_7697);
nand U7951 (N_7951,N_7653,N_7739);
nand U7952 (N_7952,N_7600,N_7603);
nand U7953 (N_7953,N_7791,N_7772);
or U7954 (N_7954,N_7787,N_7704);
or U7955 (N_7955,N_7734,N_7708);
or U7956 (N_7956,N_7727,N_7687);
nor U7957 (N_7957,N_7719,N_7776);
nand U7958 (N_7958,N_7778,N_7613);
nor U7959 (N_7959,N_7645,N_7730);
xnor U7960 (N_7960,N_7660,N_7662);
xor U7961 (N_7961,N_7771,N_7679);
nand U7962 (N_7962,N_7651,N_7696);
or U7963 (N_7963,N_7755,N_7717);
nor U7964 (N_7964,N_7659,N_7657);
xor U7965 (N_7965,N_7712,N_7738);
nor U7966 (N_7966,N_7650,N_7653);
or U7967 (N_7967,N_7733,N_7788);
or U7968 (N_7968,N_7700,N_7653);
xnor U7969 (N_7969,N_7711,N_7613);
and U7970 (N_7970,N_7643,N_7744);
nand U7971 (N_7971,N_7764,N_7780);
xnor U7972 (N_7972,N_7729,N_7616);
or U7973 (N_7973,N_7628,N_7739);
nand U7974 (N_7974,N_7674,N_7714);
or U7975 (N_7975,N_7656,N_7631);
xor U7976 (N_7976,N_7637,N_7730);
nand U7977 (N_7977,N_7760,N_7710);
xor U7978 (N_7978,N_7612,N_7716);
or U7979 (N_7979,N_7682,N_7603);
nand U7980 (N_7980,N_7633,N_7688);
and U7981 (N_7981,N_7781,N_7730);
nor U7982 (N_7982,N_7771,N_7633);
nor U7983 (N_7983,N_7747,N_7613);
or U7984 (N_7984,N_7646,N_7622);
and U7985 (N_7985,N_7769,N_7736);
nand U7986 (N_7986,N_7631,N_7750);
or U7987 (N_7987,N_7756,N_7712);
nor U7988 (N_7988,N_7703,N_7761);
nor U7989 (N_7989,N_7601,N_7693);
xor U7990 (N_7990,N_7786,N_7719);
nor U7991 (N_7991,N_7761,N_7661);
or U7992 (N_7992,N_7606,N_7736);
xnor U7993 (N_7993,N_7742,N_7643);
xnor U7994 (N_7994,N_7669,N_7674);
xor U7995 (N_7995,N_7791,N_7786);
nand U7996 (N_7996,N_7725,N_7771);
nand U7997 (N_7997,N_7788,N_7625);
nand U7998 (N_7998,N_7679,N_7703);
nand U7999 (N_7999,N_7772,N_7611);
nand U8000 (N_8000,N_7936,N_7940);
xnor U8001 (N_8001,N_7976,N_7861);
nor U8002 (N_8002,N_7832,N_7876);
or U8003 (N_8003,N_7895,N_7883);
and U8004 (N_8004,N_7965,N_7875);
and U8005 (N_8005,N_7927,N_7970);
or U8006 (N_8006,N_7975,N_7887);
nor U8007 (N_8007,N_7801,N_7998);
nor U8008 (N_8008,N_7826,N_7972);
or U8009 (N_8009,N_7837,N_7921);
xnor U8010 (N_8010,N_7977,N_7920);
xnor U8011 (N_8011,N_7850,N_7834);
or U8012 (N_8012,N_7820,N_7866);
or U8013 (N_8013,N_7821,N_7918);
xnor U8014 (N_8014,N_7819,N_7848);
xnor U8015 (N_8015,N_7956,N_7962);
nor U8016 (N_8016,N_7852,N_7950);
and U8017 (N_8017,N_7890,N_7860);
and U8018 (N_8018,N_7828,N_7856);
nor U8019 (N_8019,N_7853,N_7893);
and U8020 (N_8020,N_7859,N_7989);
nand U8021 (N_8021,N_7857,N_7872);
and U8022 (N_8022,N_7966,N_7910);
and U8023 (N_8023,N_7879,N_7980);
or U8024 (N_8024,N_7984,N_7825);
nand U8025 (N_8025,N_7897,N_7934);
xor U8026 (N_8026,N_7961,N_7891);
or U8027 (N_8027,N_7948,N_7968);
nand U8028 (N_8028,N_7967,N_7881);
and U8029 (N_8029,N_7952,N_7835);
nand U8030 (N_8030,N_7963,N_7959);
nor U8031 (N_8031,N_7924,N_7844);
and U8032 (N_8032,N_7878,N_7877);
and U8033 (N_8033,N_7944,N_7886);
or U8034 (N_8034,N_7811,N_7986);
or U8035 (N_8035,N_7930,N_7933);
and U8036 (N_8036,N_7917,N_7817);
nand U8037 (N_8037,N_7949,N_7939);
nor U8038 (N_8038,N_7882,N_7869);
and U8039 (N_8039,N_7903,N_7809);
nand U8040 (N_8040,N_7922,N_7923);
xnor U8041 (N_8041,N_7988,N_7831);
or U8042 (N_8042,N_7957,N_7953);
nor U8043 (N_8043,N_7854,N_7843);
and U8044 (N_8044,N_7894,N_7845);
or U8045 (N_8045,N_7937,N_7816);
or U8046 (N_8046,N_7992,N_7812);
and U8047 (N_8047,N_7946,N_7991);
nand U8048 (N_8048,N_7870,N_7805);
or U8049 (N_8049,N_7942,N_7987);
and U8050 (N_8050,N_7912,N_7873);
nand U8051 (N_8051,N_7838,N_7855);
and U8052 (N_8052,N_7981,N_7849);
nand U8053 (N_8053,N_7983,N_7806);
or U8054 (N_8054,N_7911,N_7851);
xnor U8055 (N_8055,N_7935,N_7958);
nand U8056 (N_8056,N_7964,N_7863);
xnor U8057 (N_8057,N_7889,N_7867);
nor U8058 (N_8058,N_7931,N_7808);
and U8059 (N_8059,N_7804,N_7892);
xor U8060 (N_8060,N_7824,N_7978);
nand U8061 (N_8061,N_7836,N_7990);
nand U8062 (N_8062,N_7862,N_7994);
or U8063 (N_8063,N_7902,N_7830);
and U8064 (N_8064,N_7943,N_7960);
nor U8065 (N_8065,N_7840,N_7813);
or U8066 (N_8066,N_7904,N_7995);
xnor U8067 (N_8067,N_7880,N_7916);
or U8068 (N_8068,N_7802,N_7979);
xor U8069 (N_8069,N_7929,N_7913);
nand U8070 (N_8070,N_7818,N_7919);
nand U8071 (N_8071,N_7810,N_7847);
nor U8072 (N_8072,N_7971,N_7996);
xnor U8073 (N_8073,N_7846,N_7815);
nor U8074 (N_8074,N_7868,N_7908);
nor U8075 (N_8075,N_7803,N_7814);
or U8076 (N_8076,N_7999,N_7951);
nor U8077 (N_8077,N_7907,N_7969);
xor U8078 (N_8078,N_7829,N_7898);
or U8079 (N_8079,N_7841,N_7865);
xnor U8080 (N_8080,N_7871,N_7874);
nand U8081 (N_8081,N_7982,N_7928);
nor U8082 (N_8082,N_7858,N_7906);
nand U8083 (N_8083,N_7842,N_7823);
xor U8084 (N_8084,N_7833,N_7974);
xnor U8085 (N_8085,N_7941,N_7926);
nand U8086 (N_8086,N_7925,N_7884);
and U8087 (N_8087,N_7899,N_7955);
nand U8088 (N_8088,N_7885,N_7947);
nor U8089 (N_8089,N_7896,N_7905);
nor U8090 (N_8090,N_7938,N_7864);
nor U8091 (N_8091,N_7993,N_7822);
xnor U8092 (N_8092,N_7915,N_7954);
nor U8093 (N_8093,N_7945,N_7914);
nor U8094 (N_8094,N_7932,N_7901);
and U8095 (N_8095,N_7827,N_7888);
nor U8096 (N_8096,N_7839,N_7985);
nand U8097 (N_8097,N_7909,N_7973);
xor U8098 (N_8098,N_7997,N_7807);
xnor U8099 (N_8099,N_7800,N_7900);
xor U8100 (N_8100,N_7830,N_7804);
or U8101 (N_8101,N_7869,N_7990);
or U8102 (N_8102,N_7950,N_7875);
and U8103 (N_8103,N_7873,N_7973);
and U8104 (N_8104,N_7911,N_7893);
and U8105 (N_8105,N_7805,N_7865);
nor U8106 (N_8106,N_7946,N_7954);
or U8107 (N_8107,N_7851,N_7800);
or U8108 (N_8108,N_7887,N_7915);
or U8109 (N_8109,N_7809,N_7894);
nor U8110 (N_8110,N_7901,N_7876);
and U8111 (N_8111,N_7902,N_7964);
nor U8112 (N_8112,N_7937,N_7889);
nor U8113 (N_8113,N_7839,N_7983);
or U8114 (N_8114,N_7988,N_7996);
xnor U8115 (N_8115,N_7815,N_7834);
nor U8116 (N_8116,N_7967,N_7959);
or U8117 (N_8117,N_7825,N_7811);
nand U8118 (N_8118,N_7980,N_7939);
nand U8119 (N_8119,N_7817,N_7898);
xor U8120 (N_8120,N_7873,N_7899);
nor U8121 (N_8121,N_7888,N_7863);
nand U8122 (N_8122,N_7852,N_7888);
or U8123 (N_8123,N_7870,N_7987);
and U8124 (N_8124,N_7970,N_7845);
nor U8125 (N_8125,N_7933,N_7897);
and U8126 (N_8126,N_7860,N_7958);
and U8127 (N_8127,N_7909,N_7998);
xnor U8128 (N_8128,N_7940,N_7834);
nand U8129 (N_8129,N_7962,N_7963);
xor U8130 (N_8130,N_7917,N_7923);
nor U8131 (N_8131,N_7989,N_7875);
or U8132 (N_8132,N_7956,N_7995);
or U8133 (N_8133,N_7888,N_7948);
nand U8134 (N_8134,N_7952,N_7946);
nor U8135 (N_8135,N_7922,N_7829);
and U8136 (N_8136,N_7951,N_7940);
and U8137 (N_8137,N_7932,N_7962);
xor U8138 (N_8138,N_7902,N_7844);
nor U8139 (N_8139,N_7979,N_7900);
and U8140 (N_8140,N_7916,N_7910);
nor U8141 (N_8141,N_7943,N_7807);
or U8142 (N_8142,N_7911,N_7818);
and U8143 (N_8143,N_7890,N_7807);
or U8144 (N_8144,N_7874,N_7869);
or U8145 (N_8145,N_7954,N_7962);
or U8146 (N_8146,N_7917,N_7826);
nor U8147 (N_8147,N_7926,N_7878);
nand U8148 (N_8148,N_7968,N_7853);
xnor U8149 (N_8149,N_7980,N_7906);
nor U8150 (N_8150,N_7880,N_7896);
and U8151 (N_8151,N_7947,N_7938);
or U8152 (N_8152,N_7808,N_7888);
or U8153 (N_8153,N_7925,N_7997);
xnor U8154 (N_8154,N_7839,N_7996);
nand U8155 (N_8155,N_7959,N_7928);
and U8156 (N_8156,N_7871,N_7906);
and U8157 (N_8157,N_7882,N_7881);
xor U8158 (N_8158,N_7946,N_7867);
xnor U8159 (N_8159,N_7999,N_7978);
nand U8160 (N_8160,N_7813,N_7883);
xnor U8161 (N_8161,N_7972,N_7910);
xor U8162 (N_8162,N_7905,N_7898);
nor U8163 (N_8163,N_7863,N_7937);
or U8164 (N_8164,N_7865,N_7908);
or U8165 (N_8165,N_7862,N_7802);
and U8166 (N_8166,N_7867,N_7829);
nand U8167 (N_8167,N_7973,N_7947);
nor U8168 (N_8168,N_7984,N_7978);
and U8169 (N_8169,N_7960,N_7837);
xor U8170 (N_8170,N_7923,N_7935);
or U8171 (N_8171,N_7924,N_7823);
xnor U8172 (N_8172,N_7943,N_7909);
nor U8173 (N_8173,N_7940,N_7865);
and U8174 (N_8174,N_7810,N_7972);
nand U8175 (N_8175,N_7945,N_7988);
and U8176 (N_8176,N_7963,N_7823);
nor U8177 (N_8177,N_7887,N_7936);
or U8178 (N_8178,N_7983,N_7969);
or U8179 (N_8179,N_7808,N_7819);
nand U8180 (N_8180,N_7856,N_7923);
xor U8181 (N_8181,N_7879,N_7903);
or U8182 (N_8182,N_7870,N_7929);
nor U8183 (N_8183,N_7916,N_7816);
or U8184 (N_8184,N_7881,N_7898);
and U8185 (N_8185,N_7873,N_7876);
nor U8186 (N_8186,N_7809,N_7806);
xnor U8187 (N_8187,N_7901,N_7890);
or U8188 (N_8188,N_7952,N_7988);
nand U8189 (N_8189,N_7919,N_7897);
or U8190 (N_8190,N_7911,N_7821);
nand U8191 (N_8191,N_7806,N_7917);
nor U8192 (N_8192,N_7910,N_7873);
xnor U8193 (N_8193,N_7823,N_7848);
or U8194 (N_8194,N_7832,N_7812);
xnor U8195 (N_8195,N_7977,N_7948);
nand U8196 (N_8196,N_7868,N_7947);
and U8197 (N_8197,N_7965,N_7872);
nor U8198 (N_8198,N_7993,N_7987);
nand U8199 (N_8199,N_7868,N_7995);
nor U8200 (N_8200,N_8134,N_8082);
xor U8201 (N_8201,N_8081,N_8197);
or U8202 (N_8202,N_8014,N_8133);
nor U8203 (N_8203,N_8145,N_8062);
or U8204 (N_8204,N_8075,N_8066);
xor U8205 (N_8205,N_8119,N_8091);
nand U8206 (N_8206,N_8144,N_8138);
nor U8207 (N_8207,N_8123,N_8137);
and U8208 (N_8208,N_8087,N_8195);
nor U8209 (N_8209,N_8131,N_8189);
or U8210 (N_8210,N_8140,N_8172);
xor U8211 (N_8211,N_8065,N_8152);
or U8212 (N_8212,N_8072,N_8028);
or U8213 (N_8213,N_8070,N_8151);
nand U8214 (N_8214,N_8034,N_8074);
or U8215 (N_8215,N_8157,N_8049);
xnor U8216 (N_8216,N_8167,N_8135);
xor U8217 (N_8217,N_8009,N_8054);
nand U8218 (N_8218,N_8090,N_8098);
xnor U8219 (N_8219,N_8035,N_8171);
xnor U8220 (N_8220,N_8043,N_8084);
and U8221 (N_8221,N_8122,N_8096);
nand U8222 (N_8222,N_8024,N_8060);
xnor U8223 (N_8223,N_8143,N_8190);
nand U8224 (N_8224,N_8017,N_8030);
nor U8225 (N_8225,N_8177,N_8033);
or U8226 (N_8226,N_8183,N_8176);
nor U8227 (N_8227,N_8088,N_8046);
nor U8228 (N_8228,N_8185,N_8184);
nand U8229 (N_8229,N_8044,N_8001);
xnor U8230 (N_8230,N_8108,N_8048);
nor U8231 (N_8231,N_8050,N_8022);
nand U8232 (N_8232,N_8042,N_8051);
nor U8233 (N_8233,N_8193,N_8003);
xor U8234 (N_8234,N_8079,N_8045);
or U8235 (N_8235,N_8162,N_8194);
xnor U8236 (N_8236,N_8002,N_8076);
nor U8237 (N_8237,N_8187,N_8013);
nand U8238 (N_8238,N_8118,N_8020);
or U8239 (N_8239,N_8186,N_8016);
or U8240 (N_8240,N_8164,N_8080);
nor U8241 (N_8241,N_8121,N_8114);
xnor U8242 (N_8242,N_8097,N_8041);
or U8243 (N_8243,N_8115,N_8125);
or U8244 (N_8244,N_8095,N_8175);
or U8245 (N_8245,N_8163,N_8104);
nor U8246 (N_8246,N_8169,N_8128);
and U8247 (N_8247,N_8061,N_8165);
nor U8248 (N_8248,N_8141,N_8099);
nand U8249 (N_8249,N_8139,N_8101);
nor U8250 (N_8250,N_8126,N_8094);
nor U8251 (N_8251,N_8181,N_8153);
xnor U8252 (N_8252,N_8158,N_8058);
and U8253 (N_8253,N_8083,N_8064);
or U8254 (N_8254,N_8120,N_8111);
and U8255 (N_8255,N_8092,N_8019);
and U8256 (N_8256,N_8178,N_8170);
xnor U8257 (N_8257,N_8124,N_8107);
nand U8258 (N_8258,N_8057,N_8007);
nor U8259 (N_8259,N_8155,N_8038);
or U8260 (N_8260,N_8148,N_8156);
xnor U8261 (N_8261,N_8027,N_8173);
or U8262 (N_8262,N_8063,N_8086);
and U8263 (N_8263,N_8168,N_8150);
nor U8264 (N_8264,N_8077,N_8093);
nor U8265 (N_8265,N_8010,N_8073);
or U8266 (N_8266,N_8021,N_8032);
nand U8267 (N_8267,N_8085,N_8110);
nand U8268 (N_8268,N_8161,N_8117);
nor U8269 (N_8269,N_8102,N_8089);
xor U8270 (N_8270,N_8040,N_8182);
nor U8271 (N_8271,N_8059,N_8067);
nand U8272 (N_8272,N_8037,N_8047);
nand U8273 (N_8273,N_8023,N_8069);
xnor U8274 (N_8274,N_8174,N_8198);
xor U8275 (N_8275,N_8116,N_8191);
xor U8276 (N_8276,N_8029,N_8113);
and U8277 (N_8277,N_8000,N_8100);
xnor U8278 (N_8278,N_8142,N_8056);
and U8279 (N_8279,N_8106,N_8192);
xnor U8280 (N_8280,N_8136,N_8159);
or U8281 (N_8281,N_8103,N_8053);
xor U8282 (N_8282,N_8078,N_8004);
nand U8283 (N_8283,N_8071,N_8129);
nand U8284 (N_8284,N_8011,N_8132);
xnor U8285 (N_8285,N_8052,N_8068);
nand U8286 (N_8286,N_8008,N_8026);
nor U8287 (N_8287,N_8146,N_8166);
nor U8288 (N_8288,N_8055,N_8031);
and U8289 (N_8289,N_8039,N_8025);
or U8290 (N_8290,N_8180,N_8006);
nand U8291 (N_8291,N_8012,N_8005);
or U8292 (N_8292,N_8188,N_8154);
xor U8293 (N_8293,N_8109,N_8036);
xnor U8294 (N_8294,N_8147,N_8112);
nand U8295 (N_8295,N_8179,N_8199);
and U8296 (N_8296,N_8105,N_8196);
and U8297 (N_8297,N_8015,N_8018);
nor U8298 (N_8298,N_8127,N_8149);
and U8299 (N_8299,N_8160,N_8130);
xnor U8300 (N_8300,N_8073,N_8051);
and U8301 (N_8301,N_8010,N_8040);
nor U8302 (N_8302,N_8142,N_8170);
or U8303 (N_8303,N_8072,N_8113);
nor U8304 (N_8304,N_8195,N_8151);
nor U8305 (N_8305,N_8178,N_8198);
and U8306 (N_8306,N_8129,N_8002);
xor U8307 (N_8307,N_8141,N_8131);
nor U8308 (N_8308,N_8022,N_8095);
and U8309 (N_8309,N_8081,N_8052);
and U8310 (N_8310,N_8123,N_8070);
nand U8311 (N_8311,N_8027,N_8059);
and U8312 (N_8312,N_8188,N_8075);
xnor U8313 (N_8313,N_8152,N_8175);
xnor U8314 (N_8314,N_8117,N_8094);
xor U8315 (N_8315,N_8125,N_8000);
and U8316 (N_8316,N_8148,N_8081);
and U8317 (N_8317,N_8172,N_8160);
or U8318 (N_8318,N_8174,N_8133);
nand U8319 (N_8319,N_8037,N_8082);
nand U8320 (N_8320,N_8024,N_8068);
nor U8321 (N_8321,N_8082,N_8006);
nand U8322 (N_8322,N_8099,N_8061);
xor U8323 (N_8323,N_8075,N_8113);
xnor U8324 (N_8324,N_8075,N_8175);
nor U8325 (N_8325,N_8072,N_8173);
nor U8326 (N_8326,N_8016,N_8185);
xnor U8327 (N_8327,N_8083,N_8198);
nor U8328 (N_8328,N_8002,N_8124);
nand U8329 (N_8329,N_8009,N_8097);
and U8330 (N_8330,N_8031,N_8097);
or U8331 (N_8331,N_8084,N_8146);
or U8332 (N_8332,N_8149,N_8154);
and U8333 (N_8333,N_8085,N_8099);
xnor U8334 (N_8334,N_8097,N_8050);
or U8335 (N_8335,N_8033,N_8034);
and U8336 (N_8336,N_8162,N_8058);
and U8337 (N_8337,N_8014,N_8150);
nand U8338 (N_8338,N_8058,N_8069);
nand U8339 (N_8339,N_8105,N_8007);
xnor U8340 (N_8340,N_8109,N_8179);
and U8341 (N_8341,N_8034,N_8119);
nand U8342 (N_8342,N_8042,N_8086);
nor U8343 (N_8343,N_8028,N_8157);
and U8344 (N_8344,N_8056,N_8187);
or U8345 (N_8345,N_8006,N_8044);
or U8346 (N_8346,N_8111,N_8006);
and U8347 (N_8347,N_8127,N_8176);
nand U8348 (N_8348,N_8117,N_8111);
or U8349 (N_8349,N_8100,N_8089);
nor U8350 (N_8350,N_8143,N_8109);
nor U8351 (N_8351,N_8160,N_8111);
nand U8352 (N_8352,N_8140,N_8162);
nand U8353 (N_8353,N_8061,N_8104);
or U8354 (N_8354,N_8087,N_8069);
nand U8355 (N_8355,N_8038,N_8067);
xor U8356 (N_8356,N_8086,N_8058);
xor U8357 (N_8357,N_8102,N_8158);
or U8358 (N_8358,N_8175,N_8023);
nor U8359 (N_8359,N_8052,N_8025);
or U8360 (N_8360,N_8143,N_8031);
nand U8361 (N_8361,N_8073,N_8093);
and U8362 (N_8362,N_8133,N_8024);
and U8363 (N_8363,N_8109,N_8063);
and U8364 (N_8364,N_8194,N_8016);
xnor U8365 (N_8365,N_8051,N_8116);
or U8366 (N_8366,N_8081,N_8138);
xor U8367 (N_8367,N_8060,N_8134);
or U8368 (N_8368,N_8111,N_8056);
xor U8369 (N_8369,N_8043,N_8034);
or U8370 (N_8370,N_8178,N_8071);
and U8371 (N_8371,N_8082,N_8123);
nor U8372 (N_8372,N_8108,N_8179);
nand U8373 (N_8373,N_8004,N_8172);
or U8374 (N_8374,N_8114,N_8101);
and U8375 (N_8375,N_8143,N_8104);
nand U8376 (N_8376,N_8143,N_8111);
or U8377 (N_8377,N_8148,N_8001);
and U8378 (N_8378,N_8080,N_8154);
or U8379 (N_8379,N_8045,N_8141);
nand U8380 (N_8380,N_8126,N_8180);
or U8381 (N_8381,N_8199,N_8046);
and U8382 (N_8382,N_8167,N_8136);
or U8383 (N_8383,N_8139,N_8170);
nand U8384 (N_8384,N_8196,N_8095);
xor U8385 (N_8385,N_8011,N_8007);
xnor U8386 (N_8386,N_8171,N_8027);
xnor U8387 (N_8387,N_8123,N_8093);
and U8388 (N_8388,N_8182,N_8076);
and U8389 (N_8389,N_8130,N_8124);
nand U8390 (N_8390,N_8196,N_8187);
xnor U8391 (N_8391,N_8177,N_8027);
or U8392 (N_8392,N_8171,N_8170);
xnor U8393 (N_8393,N_8166,N_8022);
nor U8394 (N_8394,N_8088,N_8000);
xor U8395 (N_8395,N_8100,N_8091);
or U8396 (N_8396,N_8178,N_8144);
nand U8397 (N_8397,N_8128,N_8156);
nor U8398 (N_8398,N_8014,N_8091);
or U8399 (N_8399,N_8068,N_8154);
nor U8400 (N_8400,N_8340,N_8378);
and U8401 (N_8401,N_8370,N_8246);
or U8402 (N_8402,N_8341,N_8372);
and U8403 (N_8403,N_8350,N_8365);
and U8404 (N_8404,N_8251,N_8247);
nor U8405 (N_8405,N_8376,N_8267);
nand U8406 (N_8406,N_8225,N_8294);
nand U8407 (N_8407,N_8362,N_8269);
and U8408 (N_8408,N_8345,N_8383);
nand U8409 (N_8409,N_8399,N_8289);
xnor U8410 (N_8410,N_8297,N_8238);
nor U8411 (N_8411,N_8302,N_8286);
nor U8412 (N_8412,N_8306,N_8321);
or U8413 (N_8413,N_8208,N_8346);
nand U8414 (N_8414,N_8356,N_8369);
nor U8415 (N_8415,N_8351,N_8298);
nor U8416 (N_8416,N_8311,N_8248);
xnor U8417 (N_8417,N_8388,N_8256);
or U8418 (N_8418,N_8393,N_8221);
or U8419 (N_8419,N_8352,N_8366);
nand U8420 (N_8420,N_8230,N_8257);
and U8421 (N_8421,N_8210,N_8397);
and U8422 (N_8422,N_8308,N_8220);
and U8423 (N_8423,N_8342,N_8389);
nand U8424 (N_8424,N_8374,N_8395);
nand U8425 (N_8425,N_8327,N_8270);
or U8426 (N_8426,N_8272,N_8285);
nand U8427 (N_8427,N_8275,N_8283);
and U8428 (N_8428,N_8320,N_8343);
nor U8429 (N_8429,N_8240,N_8266);
nor U8430 (N_8430,N_8313,N_8245);
or U8431 (N_8431,N_8203,N_8334);
nand U8432 (N_8432,N_8337,N_8277);
and U8433 (N_8433,N_8265,N_8358);
nor U8434 (N_8434,N_8259,N_8328);
xor U8435 (N_8435,N_8214,N_8202);
nand U8436 (N_8436,N_8258,N_8296);
or U8437 (N_8437,N_8288,N_8200);
nor U8438 (N_8438,N_8386,N_8316);
and U8439 (N_8439,N_8304,N_8241);
and U8440 (N_8440,N_8305,N_8355);
nand U8441 (N_8441,N_8254,N_8377);
xor U8442 (N_8442,N_8209,N_8293);
nand U8443 (N_8443,N_8219,N_8222);
nor U8444 (N_8444,N_8236,N_8260);
nor U8445 (N_8445,N_8391,N_8398);
xor U8446 (N_8446,N_8216,N_8299);
or U8447 (N_8447,N_8335,N_8368);
nand U8448 (N_8448,N_8255,N_8371);
or U8449 (N_8449,N_8344,N_8367);
nor U8450 (N_8450,N_8326,N_8339);
xnor U8451 (N_8451,N_8360,N_8291);
or U8452 (N_8452,N_8348,N_8315);
and U8453 (N_8453,N_8295,N_8274);
xor U8454 (N_8454,N_8310,N_8354);
and U8455 (N_8455,N_8278,N_8234);
xor U8456 (N_8456,N_8264,N_8357);
nand U8457 (N_8457,N_8280,N_8282);
xor U8458 (N_8458,N_8330,N_8281);
xor U8459 (N_8459,N_8307,N_8211);
and U8460 (N_8460,N_8381,N_8226);
nor U8461 (N_8461,N_8396,N_8217);
nor U8462 (N_8462,N_8215,N_8213);
or U8463 (N_8463,N_8359,N_8392);
or U8464 (N_8464,N_8323,N_8224);
or U8465 (N_8465,N_8312,N_8394);
and U8466 (N_8466,N_8232,N_8290);
nand U8467 (N_8467,N_8375,N_8300);
nor U8468 (N_8468,N_8336,N_8218);
nor U8469 (N_8469,N_8373,N_8233);
or U8470 (N_8470,N_8324,N_8271);
xor U8471 (N_8471,N_8204,N_8364);
nand U8472 (N_8472,N_8262,N_8244);
nor U8473 (N_8473,N_8287,N_8338);
nand U8474 (N_8474,N_8279,N_8361);
and U8475 (N_8475,N_8273,N_8243);
and U8476 (N_8476,N_8318,N_8363);
nand U8477 (N_8477,N_8390,N_8303);
nor U8478 (N_8478,N_8201,N_8206);
nor U8479 (N_8479,N_8237,N_8332);
xnor U8480 (N_8480,N_8347,N_8231);
nor U8481 (N_8481,N_8252,N_8239);
or U8482 (N_8482,N_8387,N_8207);
or U8483 (N_8483,N_8379,N_8212);
or U8484 (N_8484,N_8382,N_8268);
xor U8485 (N_8485,N_8253,N_8380);
or U8486 (N_8486,N_8250,N_8263);
or U8487 (N_8487,N_8317,N_8325);
or U8488 (N_8488,N_8276,N_8322);
nand U8489 (N_8489,N_8249,N_8331);
or U8490 (N_8490,N_8385,N_8349);
nor U8491 (N_8491,N_8261,N_8284);
nor U8492 (N_8492,N_8301,N_8309);
nand U8493 (N_8493,N_8329,N_8235);
or U8494 (N_8494,N_8292,N_8223);
and U8495 (N_8495,N_8384,N_8319);
or U8496 (N_8496,N_8314,N_8227);
or U8497 (N_8497,N_8228,N_8333);
and U8498 (N_8498,N_8353,N_8205);
nand U8499 (N_8499,N_8229,N_8242);
and U8500 (N_8500,N_8277,N_8338);
nand U8501 (N_8501,N_8355,N_8286);
nor U8502 (N_8502,N_8301,N_8395);
nor U8503 (N_8503,N_8304,N_8281);
xnor U8504 (N_8504,N_8250,N_8254);
nor U8505 (N_8505,N_8305,N_8379);
xnor U8506 (N_8506,N_8217,N_8391);
nor U8507 (N_8507,N_8392,N_8280);
nand U8508 (N_8508,N_8288,N_8285);
nand U8509 (N_8509,N_8375,N_8391);
xnor U8510 (N_8510,N_8365,N_8221);
nand U8511 (N_8511,N_8365,N_8245);
xnor U8512 (N_8512,N_8252,N_8308);
nor U8513 (N_8513,N_8395,N_8273);
or U8514 (N_8514,N_8375,N_8396);
or U8515 (N_8515,N_8245,N_8299);
xor U8516 (N_8516,N_8240,N_8331);
nand U8517 (N_8517,N_8233,N_8214);
xnor U8518 (N_8518,N_8247,N_8344);
and U8519 (N_8519,N_8264,N_8349);
and U8520 (N_8520,N_8245,N_8308);
or U8521 (N_8521,N_8300,N_8395);
and U8522 (N_8522,N_8372,N_8353);
and U8523 (N_8523,N_8231,N_8395);
xnor U8524 (N_8524,N_8369,N_8352);
and U8525 (N_8525,N_8307,N_8305);
nand U8526 (N_8526,N_8294,N_8359);
nor U8527 (N_8527,N_8268,N_8319);
or U8528 (N_8528,N_8275,N_8344);
or U8529 (N_8529,N_8293,N_8341);
nor U8530 (N_8530,N_8299,N_8266);
and U8531 (N_8531,N_8207,N_8378);
nor U8532 (N_8532,N_8393,N_8282);
xor U8533 (N_8533,N_8341,N_8395);
nand U8534 (N_8534,N_8371,N_8204);
nor U8535 (N_8535,N_8221,N_8358);
and U8536 (N_8536,N_8327,N_8271);
or U8537 (N_8537,N_8261,N_8214);
xor U8538 (N_8538,N_8207,N_8251);
nor U8539 (N_8539,N_8337,N_8346);
or U8540 (N_8540,N_8375,N_8367);
xnor U8541 (N_8541,N_8304,N_8209);
xor U8542 (N_8542,N_8206,N_8213);
nand U8543 (N_8543,N_8300,N_8352);
or U8544 (N_8544,N_8305,N_8252);
nor U8545 (N_8545,N_8379,N_8326);
nor U8546 (N_8546,N_8260,N_8252);
nor U8547 (N_8547,N_8297,N_8273);
nor U8548 (N_8548,N_8367,N_8391);
xor U8549 (N_8549,N_8235,N_8300);
or U8550 (N_8550,N_8392,N_8278);
nand U8551 (N_8551,N_8295,N_8299);
nand U8552 (N_8552,N_8314,N_8274);
xnor U8553 (N_8553,N_8263,N_8251);
xnor U8554 (N_8554,N_8296,N_8238);
nand U8555 (N_8555,N_8223,N_8344);
nand U8556 (N_8556,N_8277,N_8254);
xor U8557 (N_8557,N_8220,N_8248);
nor U8558 (N_8558,N_8257,N_8351);
or U8559 (N_8559,N_8307,N_8364);
nor U8560 (N_8560,N_8255,N_8217);
xnor U8561 (N_8561,N_8258,N_8394);
xor U8562 (N_8562,N_8328,N_8238);
nand U8563 (N_8563,N_8308,N_8250);
or U8564 (N_8564,N_8253,N_8358);
nand U8565 (N_8565,N_8386,N_8250);
or U8566 (N_8566,N_8214,N_8270);
nor U8567 (N_8567,N_8395,N_8311);
or U8568 (N_8568,N_8289,N_8326);
nor U8569 (N_8569,N_8211,N_8372);
nor U8570 (N_8570,N_8312,N_8351);
or U8571 (N_8571,N_8210,N_8366);
and U8572 (N_8572,N_8315,N_8359);
or U8573 (N_8573,N_8288,N_8397);
xnor U8574 (N_8574,N_8236,N_8297);
and U8575 (N_8575,N_8339,N_8275);
xor U8576 (N_8576,N_8379,N_8291);
nor U8577 (N_8577,N_8204,N_8229);
or U8578 (N_8578,N_8329,N_8231);
or U8579 (N_8579,N_8307,N_8266);
nor U8580 (N_8580,N_8283,N_8346);
xnor U8581 (N_8581,N_8237,N_8390);
and U8582 (N_8582,N_8298,N_8320);
xnor U8583 (N_8583,N_8229,N_8282);
and U8584 (N_8584,N_8267,N_8316);
nor U8585 (N_8585,N_8342,N_8208);
nor U8586 (N_8586,N_8297,N_8394);
nand U8587 (N_8587,N_8208,N_8249);
or U8588 (N_8588,N_8326,N_8262);
nor U8589 (N_8589,N_8265,N_8204);
xor U8590 (N_8590,N_8214,N_8361);
xnor U8591 (N_8591,N_8396,N_8248);
xor U8592 (N_8592,N_8256,N_8211);
nand U8593 (N_8593,N_8377,N_8323);
nand U8594 (N_8594,N_8252,N_8264);
nor U8595 (N_8595,N_8364,N_8286);
and U8596 (N_8596,N_8375,N_8227);
nand U8597 (N_8597,N_8315,N_8258);
and U8598 (N_8598,N_8295,N_8372);
nand U8599 (N_8599,N_8255,N_8380);
xor U8600 (N_8600,N_8560,N_8454);
nand U8601 (N_8601,N_8557,N_8462);
nand U8602 (N_8602,N_8504,N_8412);
nor U8603 (N_8603,N_8401,N_8516);
nor U8604 (N_8604,N_8506,N_8427);
nor U8605 (N_8605,N_8419,N_8459);
or U8606 (N_8606,N_8501,N_8574);
nor U8607 (N_8607,N_8542,N_8416);
nand U8608 (N_8608,N_8596,N_8407);
xor U8609 (N_8609,N_8476,N_8442);
xnor U8610 (N_8610,N_8447,N_8452);
xor U8611 (N_8611,N_8472,N_8525);
xnor U8612 (N_8612,N_8543,N_8505);
xnor U8613 (N_8613,N_8541,N_8456);
nand U8614 (N_8614,N_8530,N_8413);
xor U8615 (N_8615,N_8575,N_8555);
nand U8616 (N_8616,N_8517,N_8518);
xnor U8617 (N_8617,N_8545,N_8551);
xnor U8618 (N_8618,N_8582,N_8550);
nor U8619 (N_8619,N_8467,N_8532);
xor U8620 (N_8620,N_8562,N_8586);
or U8621 (N_8621,N_8421,N_8563);
xor U8622 (N_8622,N_8438,N_8593);
nor U8623 (N_8623,N_8410,N_8417);
nand U8624 (N_8624,N_8439,N_8430);
nand U8625 (N_8625,N_8585,N_8415);
or U8626 (N_8626,N_8468,N_8507);
and U8627 (N_8627,N_8423,N_8595);
nand U8628 (N_8628,N_8564,N_8526);
nor U8629 (N_8629,N_8475,N_8571);
nor U8630 (N_8630,N_8524,N_8469);
nor U8631 (N_8631,N_8455,N_8435);
or U8632 (N_8632,N_8559,N_8436);
or U8633 (N_8633,N_8514,N_8498);
nor U8634 (N_8634,N_8408,N_8466);
nor U8635 (N_8635,N_8544,N_8553);
nand U8636 (N_8636,N_8428,N_8448);
or U8637 (N_8637,N_8493,N_8481);
nand U8638 (N_8638,N_8426,N_8473);
and U8639 (N_8639,N_8495,N_8418);
xnor U8640 (N_8640,N_8597,N_8443);
xnor U8641 (N_8641,N_8536,N_8533);
xor U8642 (N_8642,N_8433,N_8569);
nand U8643 (N_8643,N_8486,N_8519);
nor U8644 (N_8644,N_8441,N_8568);
xor U8645 (N_8645,N_8485,N_8409);
nor U8646 (N_8646,N_8405,N_8477);
and U8647 (N_8647,N_8509,N_8592);
and U8648 (N_8648,N_8583,N_8523);
xor U8649 (N_8649,N_8515,N_8449);
nand U8650 (N_8650,N_8487,N_8591);
xnor U8651 (N_8651,N_8598,N_8502);
or U8652 (N_8652,N_8414,N_8589);
nor U8653 (N_8653,N_8579,N_8461);
nand U8654 (N_8654,N_8534,N_8552);
or U8655 (N_8655,N_8482,N_8402);
or U8656 (N_8656,N_8520,N_8494);
nand U8657 (N_8657,N_8500,N_8577);
or U8658 (N_8658,N_8599,N_8513);
and U8659 (N_8659,N_8471,N_8573);
and U8660 (N_8660,N_8445,N_8465);
nor U8661 (N_8661,N_8411,N_8479);
xnor U8662 (N_8662,N_8420,N_8588);
and U8663 (N_8663,N_8554,N_8444);
nand U8664 (N_8664,N_8440,N_8457);
xor U8665 (N_8665,N_8546,N_8572);
nand U8666 (N_8666,N_8522,N_8531);
or U8667 (N_8667,N_8499,N_8431);
and U8668 (N_8668,N_8529,N_8460);
xor U8669 (N_8669,N_8537,N_8483);
nor U8670 (N_8670,N_8450,N_8581);
and U8671 (N_8671,N_8566,N_8548);
nand U8672 (N_8672,N_8510,N_8496);
xnor U8673 (N_8673,N_8474,N_8549);
and U8674 (N_8674,N_8511,N_8434);
or U8675 (N_8675,N_8538,N_8490);
and U8676 (N_8676,N_8429,N_8503);
xnor U8677 (N_8677,N_8578,N_8489);
and U8678 (N_8678,N_8446,N_8508);
and U8679 (N_8679,N_8587,N_8478);
nand U8680 (N_8680,N_8463,N_8540);
nor U8681 (N_8681,N_8512,N_8521);
nand U8682 (N_8682,N_8451,N_8484);
or U8683 (N_8683,N_8565,N_8422);
xor U8684 (N_8684,N_8437,N_8480);
and U8685 (N_8685,N_8528,N_8567);
or U8686 (N_8686,N_8406,N_8590);
nand U8687 (N_8687,N_8558,N_8539);
nor U8688 (N_8688,N_8453,N_8570);
and U8689 (N_8689,N_8580,N_8424);
xnor U8690 (N_8690,N_8584,N_8470);
and U8691 (N_8691,N_8464,N_8547);
and U8692 (N_8692,N_8432,N_8400);
and U8693 (N_8693,N_8404,N_8492);
nand U8694 (N_8694,N_8535,N_8556);
and U8695 (N_8695,N_8576,N_8497);
or U8696 (N_8696,N_8527,N_8458);
nor U8697 (N_8697,N_8488,N_8403);
and U8698 (N_8698,N_8425,N_8491);
nand U8699 (N_8699,N_8561,N_8594);
and U8700 (N_8700,N_8543,N_8482);
xor U8701 (N_8701,N_8520,N_8497);
or U8702 (N_8702,N_8586,N_8457);
nor U8703 (N_8703,N_8410,N_8519);
nor U8704 (N_8704,N_8414,N_8431);
nand U8705 (N_8705,N_8479,N_8430);
and U8706 (N_8706,N_8432,N_8560);
or U8707 (N_8707,N_8567,N_8583);
or U8708 (N_8708,N_8574,N_8427);
nor U8709 (N_8709,N_8431,N_8467);
or U8710 (N_8710,N_8561,N_8513);
xor U8711 (N_8711,N_8570,N_8477);
nor U8712 (N_8712,N_8411,N_8427);
and U8713 (N_8713,N_8582,N_8564);
nor U8714 (N_8714,N_8563,N_8427);
and U8715 (N_8715,N_8447,N_8423);
or U8716 (N_8716,N_8584,N_8409);
xnor U8717 (N_8717,N_8518,N_8410);
and U8718 (N_8718,N_8485,N_8418);
nor U8719 (N_8719,N_8421,N_8489);
xor U8720 (N_8720,N_8508,N_8463);
xnor U8721 (N_8721,N_8421,N_8418);
nand U8722 (N_8722,N_8545,N_8534);
or U8723 (N_8723,N_8412,N_8578);
and U8724 (N_8724,N_8418,N_8490);
nand U8725 (N_8725,N_8403,N_8587);
xnor U8726 (N_8726,N_8554,N_8595);
and U8727 (N_8727,N_8556,N_8448);
and U8728 (N_8728,N_8511,N_8557);
xor U8729 (N_8729,N_8455,N_8432);
nand U8730 (N_8730,N_8576,N_8437);
xor U8731 (N_8731,N_8544,N_8477);
and U8732 (N_8732,N_8454,N_8540);
nor U8733 (N_8733,N_8581,N_8542);
nor U8734 (N_8734,N_8591,N_8544);
xor U8735 (N_8735,N_8538,N_8574);
nor U8736 (N_8736,N_8421,N_8582);
nor U8737 (N_8737,N_8585,N_8470);
nand U8738 (N_8738,N_8591,N_8418);
xnor U8739 (N_8739,N_8493,N_8579);
nor U8740 (N_8740,N_8471,N_8579);
or U8741 (N_8741,N_8576,N_8454);
nor U8742 (N_8742,N_8567,N_8429);
nor U8743 (N_8743,N_8407,N_8588);
and U8744 (N_8744,N_8458,N_8489);
or U8745 (N_8745,N_8596,N_8411);
nand U8746 (N_8746,N_8403,N_8443);
xnor U8747 (N_8747,N_8494,N_8576);
nand U8748 (N_8748,N_8417,N_8567);
nand U8749 (N_8749,N_8550,N_8519);
and U8750 (N_8750,N_8590,N_8435);
xor U8751 (N_8751,N_8594,N_8411);
nand U8752 (N_8752,N_8430,N_8526);
or U8753 (N_8753,N_8478,N_8512);
nor U8754 (N_8754,N_8471,N_8529);
nor U8755 (N_8755,N_8519,N_8490);
nand U8756 (N_8756,N_8574,N_8592);
xor U8757 (N_8757,N_8454,N_8414);
nor U8758 (N_8758,N_8539,N_8424);
nand U8759 (N_8759,N_8434,N_8487);
nand U8760 (N_8760,N_8497,N_8592);
nand U8761 (N_8761,N_8435,N_8464);
and U8762 (N_8762,N_8521,N_8568);
nand U8763 (N_8763,N_8417,N_8497);
nand U8764 (N_8764,N_8581,N_8595);
and U8765 (N_8765,N_8459,N_8426);
nor U8766 (N_8766,N_8586,N_8452);
nand U8767 (N_8767,N_8482,N_8562);
xnor U8768 (N_8768,N_8466,N_8539);
nand U8769 (N_8769,N_8559,N_8404);
and U8770 (N_8770,N_8418,N_8584);
nor U8771 (N_8771,N_8584,N_8533);
or U8772 (N_8772,N_8446,N_8502);
and U8773 (N_8773,N_8493,N_8553);
and U8774 (N_8774,N_8507,N_8502);
xor U8775 (N_8775,N_8449,N_8408);
nor U8776 (N_8776,N_8517,N_8459);
nor U8777 (N_8777,N_8448,N_8469);
nand U8778 (N_8778,N_8492,N_8461);
nand U8779 (N_8779,N_8502,N_8528);
and U8780 (N_8780,N_8557,N_8402);
nand U8781 (N_8781,N_8491,N_8501);
or U8782 (N_8782,N_8484,N_8434);
or U8783 (N_8783,N_8449,N_8486);
or U8784 (N_8784,N_8506,N_8406);
and U8785 (N_8785,N_8408,N_8486);
nand U8786 (N_8786,N_8512,N_8544);
nor U8787 (N_8787,N_8582,N_8579);
nand U8788 (N_8788,N_8594,N_8532);
nand U8789 (N_8789,N_8497,N_8594);
nand U8790 (N_8790,N_8518,N_8438);
xnor U8791 (N_8791,N_8472,N_8409);
nand U8792 (N_8792,N_8573,N_8587);
nor U8793 (N_8793,N_8597,N_8401);
and U8794 (N_8794,N_8545,N_8441);
and U8795 (N_8795,N_8430,N_8413);
or U8796 (N_8796,N_8572,N_8413);
and U8797 (N_8797,N_8423,N_8433);
and U8798 (N_8798,N_8542,N_8550);
xnor U8799 (N_8799,N_8483,N_8432);
xor U8800 (N_8800,N_8725,N_8644);
xnor U8801 (N_8801,N_8692,N_8791);
nor U8802 (N_8802,N_8659,N_8719);
nand U8803 (N_8803,N_8765,N_8636);
nand U8804 (N_8804,N_8735,N_8766);
nor U8805 (N_8805,N_8618,N_8738);
nand U8806 (N_8806,N_8747,N_8761);
and U8807 (N_8807,N_8709,N_8693);
xor U8808 (N_8808,N_8619,N_8694);
and U8809 (N_8809,N_8617,N_8634);
and U8810 (N_8810,N_8625,N_8751);
and U8811 (N_8811,N_8600,N_8796);
and U8812 (N_8812,N_8641,N_8744);
or U8813 (N_8813,N_8767,N_8718);
xnor U8814 (N_8814,N_8724,N_8611);
xor U8815 (N_8815,N_8760,N_8605);
or U8816 (N_8816,N_8731,N_8601);
or U8817 (N_8817,N_8717,N_8670);
nand U8818 (N_8818,N_8784,N_8739);
nor U8819 (N_8819,N_8777,N_8632);
nor U8820 (N_8820,N_8713,N_8716);
nor U8821 (N_8821,N_8736,N_8706);
nor U8822 (N_8822,N_8762,N_8745);
nor U8823 (N_8823,N_8781,N_8633);
nand U8824 (N_8824,N_8612,N_8666);
and U8825 (N_8825,N_8780,N_8771);
nor U8826 (N_8826,N_8732,N_8671);
nor U8827 (N_8827,N_8770,N_8646);
and U8828 (N_8828,N_8668,N_8654);
xor U8829 (N_8829,N_8757,N_8728);
and U8830 (N_8830,N_8793,N_8642);
xnor U8831 (N_8831,N_8686,N_8613);
and U8832 (N_8832,N_8789,N_8710);
and U8833 (N_8833,N_8622,N_8786);
nor U8834 (N_8834,N_8750,N_8741);
and U8835 (N_8835,N_8701,N_8697);
nor U8836 (N_8836,N_8788,N_8655);
and U8837 (N_8837,N_8626,N_8620);
nand U8838 (N_8838,N_8779,N_8755);
and U8839 (N_8839,N_8608,N_8743);
nand U8840 (N_8840,N_8683,N_8763);
and U8841 (N_8841,N_8638,N_8690);
nand U8842 (N_8842,N_8773,N_8794);
nor U8843 (N_8843,N_8695,N_8676);
nand U8844 (N_8844,N_8774,N_8639);
or U8845 (N_8845,N_8722,N_8696);
nand U8846 (N_8846,N_8698,N_8720);
or U8847 (N_8847,N_8687,N_8606);
nand U8848 (N_8848,N_8652,N_8792);
or U8849 (N_8849,N_8680,N_8637);
xnor U8850 (N_8850,N_8707,N_8653);
nand U8851 (N_8851,N_8658,N_8663);
nor U8852 (N_8852,N_8799,N_8688);
nor U8853 (N_8853,N_8685,N_8700);
and U8854 (N_8854,N_8629,N_8769);
or U8855 (N_8855,N_8754,N_8705);
or U8856 (N_8856,N_8649,N_8785);
nand U8857 (N_8857,N_8733,N_8616);
or U8858 (N_8858,N_8702,N_8635);
xor U8859 (N_8859,N_8778,N_8651);
or U8860 (N_8860,N_8602,N_8787);
and U8861 (N_8861,N_8795,N_8630);
or U8862 (N_8862,N_8758,N_8782);
nand U8863 (N_8863,N_8662,N_8624);
nand U8864 (N_8864,N_8689,N_8740);
xor U8865 (N_8865,N_8684,N_8703);
and U8866 (N_8866,N_8746,N_8631);
nand U8867 (N_8867,N_8628,N_8607);
nor U8868 (N_8868,N_8772,N_8661);
nor U8869 (N_8869,N_8749,N_8621);
and U8870 (N_8870,N_8603,N_8678);
nor U8871 (N_8871,N_8648,N_8764);
nor U8872 (N_8872,N_8759,N_8726);
xnor U8873 (N_8873,N_8610,N_8776);
and U8874 (N_8874,N_8708,N_8756);
nor U8875 (N_8875,N_8714,N_8650);
xnor U8876 (N_8876,N_8730,N_8729);
nor U8877 (N_8877,N_8677,N_8669);
nor U8878 (N_8878,N_8615,N_8775);
or U8879 (N_8879,N_8748,N_8704);
or U8880 (N_8880,N_8643,N_8627);
or U8881 (N_8881,N_8604,N_8674);
xor U8882 (N_8882,N_8656,N_8711);
and U8883 (N_8883,N_8673,N_8797);
nand U8884 (N_8884,N_8691,N_8681);
nand U8885 (N_8885,N_8679,N_8667);
xnor U8886 (N_8886,N_8609,N_8721);
nor U8887 (N_8887,N_8672,N_8734);
or U8888 (N_8888,N_8712,N_8742);
and U8889 (N_8889,N_8664,N_8753);
nand U8890 (N_8890,N_8647,N_8665);
and U8891 (N_8891,N_8660,N_8783);
xnor U8892 (N_8892,N_8623,N_8614);
xnor U8893 (N_8893,N_8640,N_8657);
xnor U8894 (N_8894,N_8682,N_8723);
or U8895 (N_8895,N_8798,N_8768);
or U8896 (N_8896,N_8737,N_8645);
or U8897 (N_8897,N_8715,N_8752);
nand U8898 (N_8898,N_8675,N_8699);
nor U8899 (N_8899,N_8727,N_8790);
nand U8900 (N_8900,N_8722,N_8788);
xnor U8901 (N_8901,N_8731,N_8614);
and U8902 (N_8902,N_8694,N_8766);
nand U8903 (N_8903,N_8677,N_8706);
or U8904 (N_8904,N_8711,N_8763);
nor U8905 (N_8905,N_8773,N_8612);
nor U8906 (N_8906,N_8682,N_8738);
or U8907 (N_8907,N_8676,N_8773);
and U8908 (N_8908,N_8735,N_8760);
xnor U8909 (N_8909,N_8607,N_8675);
and U8910 (N_8910,N_8794,N_8795);
nand U8911 (N_8911,N_8636,N_8762);
nor U8912 (N_8912,N_8786,N_8683);
xor U8913 (N_8913,N_8699,N_8697);
nor U8914 (N_8914,N_8773,N_8626);
and U8915 (N_8915,N_8798,N_8748);
xor U8916 (N_8916,N_8613,N_8798);
and U8917 (N_8917,N_8643,N_8608);
and U8918 (N_8918,N_8742,N_8616);
and U8919 (N_8919,N_8623,N_8726);
or U8920 (N_8920,N_8781,N_8625);
or U8921 (N_8921,N_8719,N_8711);
nor U8922 (N_8922,N_8722,N_8683);
or U8923 (N_8923,N_8744,N_8687);
xnor U8924 (N_8924,N_8630,N_8738);
and U8925 (N_8925,N_8677,N_8656);
nor U8926 (N_8926,N_8768,N_8670);
nor U8927 (N_8927,N_8742,N_8624);
xnor U8928 (N_8928,N_8788,N_8669);
xnor U8929 (N_8929,N_8727,N_8766);
xor U8930 (N_8930,N_8730,N_8799);
xnor U8931 (N_8931,N_8759,N_8750);
and U8932 (N_8932,N_8629,N_8669);
and U8933 (N_8933,N_8691,N_8716);
nand U8934 (N_8934,N_8712,N_8641);
or U8935 (N_8935,N_8601,N_8754);
nor U8936 (N_8936,N_8771,N_8795);
or U8937 (N_8937,N_8637,N_8763);
xor U8938 (N_8938,N_8732,N_8712);
and U8939 (N_8939,N_8640,N_8631);
xnor U8940 (N_8940,N_8725,N_8778);
nand U8941 (N_8941,N_8715,N_8659);
xnor U8942 (N_8942,N_8724,N_8768);
nand U8943 (N_8943,N_8726,N_8777);
or U8944 (N_8944,N_8707,N_8654);
and U8945 (N_8945,N_8793,N_8795);
or U8946 (N_8946,N_8692,N_8738);
or U8947 (N_8947,N_8794,N_8732);
xnor U8948 (N_8948,N_8670,N_8735);
or U8949 (N_8949,N_8625,N_8782);
or U8950 (N_8950,N_8712,N_8688);
or U8951 (N_8951,N_8610,N_8622);
nor U8952 (N_8952,N_8684,N_8731);
nand U8953 (N_8953,N_8637,N_8665);
and U8954 (N_8954,N_8772,N_8656);
or U8955 (N_8955,N_8762,N_8665);
nand U8956 (N_8956,N_8643,N_8796);
nand U8957 (N_8957,N_8687,N_8726);
or U8958 (N_8958,N_8624,N_8725);
and U8959 (N_8959,N_8653,N_8741);
nand U8960 (N_8960,N_8739,N_8674);
xnor U8961 (N_8961,N_8720,N_8633);
nor U8962 (N_8962,N_8616,N_8697);
and U8963 (N_8963,N_8695,N_8667);
xnor U8964 (N_8964,N_8664,N_8738);
and U8965 (N_8965,N_8681,N_8737);
nor U8966 (N_8966,N_8780,N_8680);
nor U8967 (N_8967,N_8712,N_8647);
or U8968 (N_8968,N_8661,N_8655);
xor U8969 (N_8969,N_8707,N_8784);
xor U8970 (N_8970,N_8719,N_8716);
or U8971 (N_8971,N_8608,N_8738);
xnor U8972 (N_8972,N_8678,N_8665);
nand U8973 (N_8973,N_8600,N_8699);
xnor U8974 (N_8974,N_8633,N_8615);
and U8975 (N_8975,N_8767,N_8711);
and U8976 (N_8976,N_8694,N_8639);
or U8977 (N_8977,N_8775,N_8636);
xor U8978 (N_8978,N_8728,N_8655);
and U8979 (N_8979,N_8605,N_8771);
and U8980 (N_8980,N_8635,N_8632);
xnor U8981 (N_8981,N_8757,N_8628);
nor U8982 (N_8982,N_8732,N_8658);
or U8983 (N_8983,N_8653,N_8750);
xor U8984 (N_8984,N_8613,N_8743);
and U8985 (N_8985,N_8617,N_8654);
nor U8986 (N_8986,N_8628,N_8688);
xnor U8987 (N_8987,N_8777,N_8660);
xor U8988 (N_8988,N_8790,N_8714);
nand U8989 (N_8989,N_8712,N_8708);
and U8990 (N_8990,N_8772,N_8782);
and U8991 (N_8991,N_8798,N_8632);
nor U8992 (N_8992,N_8685,N_8697);
xnor U8993 (N_8993,N_8734,N_8669);
or U8994 (N_8994,N_8773,N_8724);
xor U8995 (N_8995,N_8672,N_8759);
or U8996 (N_8996,N_8754,N_8704);
nand U8997 (N_8997,N_8700,N_8722);
nand U8998 (N_8998,N_8747,N_8621);
xor U8999 (N_8999,N_8730,N_8626);
nand U9000 (N_9000,N_8994,N_8914);
nand U9001 (N_9001,N_8941,N_8852);
nor U9002 (N_9002,N_8935,N_8943);
xor U9003 (N_9003,N_8979,N_8853);
xor U9004 (N_9004,N_8868,N_8865);
or U9005 (N_9005,N_8855,N_8981);
or U9006 (N_9006,N_8802,N_8910);
or U9007 (N_9007,N_8880,N_8919);
or U9008 (N_9008,N_8801,N_8832);
or U9009 (N_9009,N_8825,N_8982);
nor U9010 (N_9010,N_8997,N_8907);
xor U9011 (N_9011,N_8992,N_8893);
and U9012 (N_9012,N_8987,N_8975);
and U9013 (N_9013,N_8995,N_8999);
nand U9014 (N_9014,N_8898,N_8953);
xor U9015 (N_9015,N_8835,N_8831);
and U9016 (N_9016,N_8937,N_8805);
nand U9017 (N_9017,N_8978,N_8957);
nor U9018 (N_9018,N_8856,N_8846);
nand U9019 (N_9019,N_8811,N_8922);
nor U9020 (N_9020,N_8845,N_8921);
and U9021 (N_9021,N_8905,N_8955);
xor U9022 (N_9022,N_8810,N_8862);
and U9023 (N_9023,N_8918,N_8840);
or U9024 (N_9024,N_8900,N_8912);
or U9025 (N_9025,N_8808,N_8988);
or U9026 (N_9026,N_8903,N_8806);
nand U9027 (N_9027,N_8863,N_8895);
nand U9028 (N_9028,N_8986,N_8976);
or U9029 (N_9029,N_8933,N_8977);
or U9030 (N_9030,N_8822,N_8944);
and U9031 (N_9031,N_8817,N_8843);
and U9032 (N_9032,N_8938,N_8899);
xnor U9033 (N_9033,N_8815,N_8948);
xor U9034 (N_9034,N_8872,N_8967);
nand U9035 (N_9035,N_8980,N_8915);
nor U9036 (N_9036,N_8871,N_8854);
or U9037 (N_9037,N_8858,N_8881);
nor U9038 (N_9038,N_8886,N_8913);
nand U9039 (N_9039,N_8823,N_8932);
nand U9040 (N_9040,N_8807,N_8896);
or U9041 (N_9041,N_8925,N_8884);
nor U9042 (N_9042,N_8973,N_8991);
and U9043 (N_9043,N_8926,N_8816);
and U9044 (N_9044,N_8847,N_8839);
nor U9045 (N_9045,N_8949,N_8965);
and U9046 (N_9046,N_8833,N_8826);
or U9047 (N_9047,N_8993,N_8878);
or U9048 (N_9048,N_8809,N_8963);
nor U9049 (N_9049,N_8964,N_8813);
or U9050 (N_9050,N_8836,N_8962);
nor U9051 (N_9051,N_8947,N_8984);
and U9052 (N_9052,N_8902,N_8950);
nor U9053 (N_9053,N_8959,N_8876);
nor U9054 (N_9054,N_8861,N_8850);
or U9055 (N_9055,N_8904,N_8911);
xnor U9056 (N_9056,N_8800,N_8875);
nor U9057 (N_9057,N_8824,N_8877);
and U9058 (N_9058,N_8945,N_8985);
xor U9059 (N_9059,N_8859,N_8972);
nand U9060 (N_9060,N_8917,N_8939);
nand U9061 (N_9061,N_8934,N_8803);
and U9062 (N_9062,N_8866,N_8916);
nand U9063 (N_9063,N_8827,N_8942);
nor U9064 (N_9064,N_8990,N_8838);
xor U9065 (N_9065,N_8829,N_8974);
or U9066 (N_9066,N_8901,N_8819);
and U9067 (N_9067,N_8882,N_8956);
nand U9068 (N_9068,N_8966,N_8830);
nand U9069 (N_9069,N_8834,N_8958);
xor U9070 (N_9070,N_8996,N_8879);
or U9071 (N_9071,N_8931,N_8844);
nor U9072 (N_9072,N_8969,N_8820);
xor U9073 (N_9073,N_8971,N_8954);
nand U9074 (N_9074,N_8883,N_8940);
and U9075 (N_9075,N_8849,N_8857);
nor U9076 (N_9076,N_8909,N_8860);
and U9077 (N_9077,N_8814,N_8891);
nand U9078 (N_9078,N_8930,N_8989);
and U9079 (N_9079,N_8894,N_8864);
xnor U9080 (N_9080,N_8848,N_8961);
xor U9081 (N_9081,N_8870,N_8983);
and U9082 (N_9082,N_8867,N_8890);
and U9083 (N_9083,N_8892,N_8887);
or U9084 (N_9084,N_8821,N_8924);
nor U9085 (N_9085,N_8968,N_8828);
and U9086 (N_9086,N_8946,N_8812);
nand U9087 (N_9087,N_8841,N_8874);
nand U9088 (N_9088,N_8929,N_8936);
nand U9089 (N_9089,N_8897,N_8818);
xnor U9090 (N_9090,N_8906,N_8923);
xnor U9091 (N_9091,N_8873,N_8889);
and U9092 (N_9092,N_8804,N_8952);
nor U9093 (N_9093,N_8888,N_8920);
and U9094 (N_9094,N_8869,N_8927);
or U9095 (N_9095,N_8851,N_8837);
and U9096 (N_9096,N_8885,N_8908);
nor U9097 (N_9097,N_8998,N_8928);
and U9098 (N_9098,N_8960,N_8951);
nor U9099 (N_9099,N_8842,N_8970);
and U9100 (N_9100,N_8977,N_8812);
nand U9101 (N_9101,N_8802,N_8985);
and U9102 (N_9102,N_8890,N_8889);
nor U9103 (N_9103,N_8997,N_8854);
and U9104 (N_9104,N_8800,N_8930);
nand U9105 (N_9105,N_8962,N_8887);
and U9106 (N_9106,N_8892,N_8942);
or U9107 (N_9107,N_8837,N_8962);
nand U9108 (N_9108,N_8835,N_8919);
xor U9109 (N_9109,N_8929,N_8801);
or U9110 (N_9110,N_8915,N_8935);
nand U9111 (N_9111,N_8930,N_8868);
nand U9112 (N_9112,N_8824,N_8947);
xnor U9113 (N_9113,N_8848,N_8821);
or U9114 (N_9114,N_8874,N_8930);
xor U9115 (N_9115,N_8972,N_8871);
and U9116 (N_9116,N_8993,N_8890);
xor U9117 (N_9117,N_8832,N_8987);
nor U9118 (N_9118,N_8821,N_8926);
and U9119 (N_9119,N_8976,N_8873);
nand U9120 (N_9120,N_8805,N_8832);
or U9121 (N_9121,N_8817,N_8895);
nor U9122 (N_9122,N_8851,N_8862);
or U9123 (N_9123,N_8823,N_8928);
xnor U9124 (N_9124,N_8807,N_8838);
xnor U9125 (N_9125,N_8822,N_8995);
or U9126 (N_9126,N_8943,N_8863);
and U9127 (N_9127,N_8980,N_8942);
nand U9128 (N_9128,N_8869,N_8889);
nand U9129 (N_9129,N_8914,N_8812);
nand U9130 (N_9130,N_8927,N_8944);
xnor U9131 (N_9131,N_8841,N_8988);
nand U9132 (N_9132,N_8924,N_8813);
nor U9133 (N_9133,N_8939,N_8963);
or U9134 (N_9134,N_8945,N_8858);
nand U9135 (N_9135,N_8845,N_8868);
nand U9136 (N_9136,N_8905,N_8945);
nand U9137 (N_9137,N_8891,N_8867);
xor U9138 (N_9138,N_8937,N_8874);
nand U9139 (N_9139,N_8890,N_8989);
xnor U9140 (N_9140,N_8956,N_8856);
nor U9141 (N_9141,N_8926,N_8872);
nand U9142 (N_9142,N_8932,N_8867);
or U9143 (N_9143,N_8807,N_8806);
nor U9144 (N_9144,N_8826,N_8925);
and U9145 (N_9145,N_8993,N_8873);
and U9146 (N_9146,N_8994,N_8834);
nand U9147 (N_9147,N_8891,N_8940);
nor U9148 (N_9148,N_8933,N_8956);
nor U9149 (N_9149,N_8824,N_8942);
and U9150 (N_9150,N_8937,N_8868);
nand U9151 (N_9151,N_8992,N_8872);
xnor U9152 (N_9152,N_8839,N_8886);
nand U9153 (N_9153,N_8922,N_8960);
xnor U9154 (N_9154,N_8984,N_8811);
or U9155 (N_9155,N_8973,N_8875);
nand U9156 (N_9156,N_8958,N_8910);
and U9157 (N_9157,N_8945,N_8937);
nor U9158 (N_9158,N_8934,N_8894);
nand U9159 (N_9159,N_8807,N_8882);
nor U9160 (N_9160,N_8822,N_8976);
and U9161 (N_9161,N_8907,N_8948);
and U9162 (N_9162,N_8850,N_8965);
and U9163 (N_9163,N_8902,N_8843);
and U9164 (N_9164,N_8859,N_8879);
and U9165 (N_9165,N_8848,N_8843);
nand U9166 (N_9166,N_8931,N_8836);
xor U9167 (N_9167,N_8865,N_8816);
nand U9168 (N_9168,N_8972,N_8867);
and U9169 (N_9169,N_8842,N_8923);
or U9170 (N_9170,N_8863,N_8930);
xnor U9171 (N_9171,N_8975,N_8985);
or U9172 (N_9172,N_8812,N_8968);
and U9173 (N_9173,N_8970,N_8992);
xnor U9174 (N_9174,N_8862,N_8869);
nand U9175 (N_9175,N_8926,N_8995);
or U9176 (N_9176,N_8875,N_8922);
or U9177 (N_9177,N_8848,N_8908);
xor U9178 (N_9178,N_8991,N_8877);
nand U9179 (N_9179,N_8855,N_8859);
xor U9180 (N_9180,N_8966,N_8995);
or U9181 (N_9181,N_8977,N_8921);
nor U9182 (N_9182,N_8878,N_8954);
nand U9183 (N_9183,N_8827,N_8807);
nor U9184 (N_9184,N_8985,N_8818);
nand U9185 (N_9185,N_8972,N_8878);
nand U9186 (N_9186,N_8967,N_8837);
or U9187 (N_9187,N_8980,N_8866);
nor U9188 (N_9188,N_8905,N_8826);
nor U9189 (N_9189,N_8815,N_8976);
or U9190 (N_9190,N_8985,N_8955);
nor U9191 (N_9191,N_8819,N_8894);
nand U9192 (N_9192,N_8966,N_8888);
and U9193 (N_9193,N_8999,N_8803);
and U9194 (N_9194,N_8824,N_8820);
or U9195 (N_9195,N_8910,N_8979);
and U9196 (N_9196,N_8883,N_8996);
nand U9197 (N_9197,N_8895,N_8988);
nand U9198 (N_9198,N_8852,N_8880);
or U9199 (N_9199,N_8899,N_8998);
nand U9200 (N_9200,N_9012,N_9077);
nand U9201 (N_9201,N_9122,N_9156);
nand U9202 (N_9202,N_9191,N_9041);
xor U9203 (N_9203,N_9151,N_9010);
or U9204 (N_9204,N_9032,N_9022);
xor U9205 (N_9205,N_9044,N_9131);
xor U9206 (N_9206,N_9154,N_9005);
and U9207 (N_9207,N_9070,N_9106);
nand U9208 (N_9208,N_9027,N_9061);
nand U9209 (N_9209,N_9132,N_9148);
or U9210 (N_9210,N_9052,N_9187);
nor U9211 (N_9211,N_9031,N_9082);
xor U9212 (N_9212,N_9109,N_9084);
xor U9213 (N_9213,N_9184,N_9193);
and U9214 (N_9214,N_9124,N_9197);
xnor U9215 (N_9215,N_9086,N_9118);
or U9216 (N_9216,N_9180,N_9046);
and U9217 (N_9217,N_9006,N_9091);
or U9218 (N_9218,N_9126,N_9105);
nand U9219 (N_9219,N_9176,N_9099);
nand U9220 (N_9220,N_9108,N_9030);
xnor U9221 (N_9221,N_9094,N_9163);
nor U9222 (N_9222,N_9165,N_9004);
nor U9223 (N_9223,N_9016,N_9159);
and U9224 (N_9224,N_9085,N_9121);
nand U9225 (N_9225,N_9059,N_9034);
nor U9226 (N_9226,N_9018,N_9185);
or U9227 (N_9227,N_9097,N_9160);
or U9228 (N_9228,N_9134,N_9172);
or U9229 (N_9229,N_9025,N_9115);
nor U9230 (N_9230,N_9069,N_9179);
nor U9231 (N_9231,N_9001,N_9083);
and U9232 (N_9232,N_9095,N_9068);
nor U9233 (N_9233,N_9064,N_9143);
and U9234 (N_9234,N_9033,N_9063);
or U9235 (N_9235,N_9152,N_9073);
nor U9236 (N_9236,N_9186,N_9168);
xor U9237 (N_9237,N_9190,N_9139);
and U9238 (N_9238,N_9011,N_9150);
or U9239 (N_9239,N_9050,N_9111);
nand U9240 (N_9240,N_9072,N_9040);
nor U9241 (N_9241,N_9123,N_9024);
or U9242 (N_9242,N_9021,N_9053);
nor U9243 (N_9243,N_9065,N_9098);
nor U9244 (N_9244,N_9110,N_9107);
or U9245 (N_9245,N_9141,N_9096);
nor U9246 (N_9246,N_9007,N_9177);
nand U9247 (N_9247,N_9116,N_9170);
nand U9248 (N_9248,N_9199,N_9000);
nor U9249 (N_9249,N_9142,N_9067);
and U9250 (N_9250,N_9146,N_9079);
xor U9251 (N_9251,N_9056,N_9066);
nand U9252 (N_9252,N_9162,N_9137);
nor U9253 (N_9253,N_9173,N_9057);
nor U9254 (N_9254,N_9092,N_9049);
nand U9255 (N_9255,N_9045,N_9080);
xnor U9256 (N_9256,N_9051,N_9003);
and U9257 (N_9257,N_9117,N_9171);
or U9258 (N_9258,N_9189,N_9135);
xor U9259 (N_9259,N_9138,N_9178);
xnor U9260 (N_9260,N_9075,N_9074);
nor U9261 (N_9261,N_9062,N_9013);
nor U9262 (N_9262,N_9039,N_9113);
and U9263 (N_9263,N_9104,N_9158);
xor U9264 (N_9264,N_9008,N_9015);
xor U9265 (N_9265,N_9153,N_9054);
nor U9266 (N_9266,N_9198,N_9164);
and U9267 (N_9267,N_9145,N_9119);
xnor U9268 (N_9268,N_9103,N_9002);
and U9269 (N_9269,N_9023,N_9081);
nor U9270 (N_9270,N_9130,N_9060);
and U9271 (N_9271,N_9088,N_9020);
nand U9272 (N_9272,N_9129,N_9161);
xor U9273 (N_9273,N_9155,N_9035);
or U9274 (N_9274,N_9102,N_9090);
and U9275 (N_9275,N_9026,N_9038);
and U9276 (N_9276,N_9157,N_9144);
nand U9277 (N_9277,N_9042,N_9112);
xor U9278 (N_9278,N_9125,N_9188);
xnor U9279 (N_9279,N_9017,N_9037);
or U9280 (N_9280,N_9166,N_9140);
or U9281 (N_9281,N_9183,N_9128);
nand U9282 (N_9282,N_9029,N_9089);
xor U9283 (N_9283,N_9133,N_9120);
and U9284 (N_9284,N_9048,N_9195);
and U9285 (N_9285,N_9181,N_9087);
nor U9286 (N_9286,N_9194,N_9071);
xnor U9287 (N_9287,N_9078,N_9147);
nand U9288 (N_9288,N_9014,N_9028);
nor U9289 (N_9289,N_9196,N_9009);
and U9290 (N_9290,N_9182,N_9127);
and U9291 (N_9291,N_9076,N_9093);
nand U9292 (N_9292,N_9058,N_9055);
xnor U9293 (N_9293,N_9100,N_9167);
xnor U9294 (N_9294,N_9101,N_9175);
or U9295 (N_9295,N_9169,N_9043);
xnor U9296 (N_9296,N_9192,N_9047);
nand U9297 (N_9297,N_9174,N_9149);
nand U9298 (N_9298,N_9136,N_9036);
xor U9299 (N_9299,N_9019,N_9114);
or U9300 (N_9300,N_9041,N_9113);
nor U9301 (N_9301,N_9151,N_9046);
and U9302 (N_9302,N_9098,N_9180);
or U9303 (N_9303,N_9022,N_9006);
nor U9304 (N_9304,N_9166,N_9078);
nand U9305 (N_9305,N_9173,N_9071);
nor U9306 (N_9306,N_9039,N_9103);
xor U9307 (N_9307,N_9062,N_9127);
xnor U9308 (N_9308,N_9084,N_9171);
nor U9309 (N_9309,N_9159,N_9186);
or U9310 (N_9310,N_9033,N_9101);
xnor U9311 (N_9311,N_9153,N_9050);
nand U9312 (N_9312,N_9038,N_9034);
nor U9313 (N_9313,N_9088,N_9159);
xor U9314 (N_9314,N_9062,N_9098);
and U9315 (N_9315,N_9054,N_9050);
nor U9316 (N_9316,N_9073,N_9197);
nor U9317 (N_9317,N_9073,N_9052);
nor U9318 (N_9318,N_9081,N_9006);
and U9319 (N_9319,N_9094,N_9060);
nand U9320 (N_9320,N_9164,N_9158);
nand U9321 (N_9321,N_9097,N_9142);
nand U9322 (N_9322,N_9030,N_9126);
and U9323 (N_9323,N_9091,N_9041);
or U9324 (N_9324,N_9015,N_9032);
and U9325 (N_9325,N_9056,N_9033);
nand U9326 (N_9326,N_9061,N_9025);
nor U9327 (N_9327,N_9135,N_9095);
and U9328 (N_9328,N_9157,N_9029);
xor U9329 (N_9329,N_9031,N_9033);
nor U9330 (N_9330,N_9130,N_9074);
nor U9331 (N_9331,N_9117,N_9053);
nand U9332 (N_9332,N_9075,N_9116);
nor U9333 (N_9333,N_9070,N_9123);
nand U9334 (N_9334,N_9086,N_9133);
xor U9335 (N_9335,N_9121,N_9046);
nor U9336 (N_9336,N_9104,N_9083);
or U9337 (N_9337,N_9093,N_9149);
or U9338 (N_9338,N_9184,N_9062);
nand U9339 (N_9339,N_9111,N_9044);
xor U9340 (N_9340,N_9149,N_9177);
nor U9341 (N_9341,N_9151,N_9033);
xnor U9342 (N_9342,N_9164,N_9115);
nand U9343 (N_9343,N_9048,N_9188);
nand U9344 (N_9344,N_9133,N_9022);
nand U9345 (N_9345,N_9173,N_9036);
nand U9346 (N_9346,N_9147,N_9069);
nor U9347 (N_9347,N_9052,N_9017);
nor U9348 (N_9348,N_9171,N_9125);
nor U9349 (N_9349,N_9169,N_9158);
and U9350 (N_9350,N_9002,N_9189);
xnor U9351 (N_9351,N_9163,N_9085);
or U9352 (N_9352,N_9085,N_9081);
nand U9353 (N_9353,N_9108,N_9029);
nand U9354 (N_9354,N_9052,N_9004);
xor U9355 (N_9355,N_9029,N_9033);
or U9356 (N_9356,N_9077,N_9144);
and U9357 (N_9357,N_9085,N_9009);
nor U9358 (N_9358,N_9186,N_9141);
or U9359 (N_9359,N_9166,N_9191);
and U9360 (N_9360,N_9012,N_9133);
nor U9361 (N_9361,N_9110,N_9129);
nor U9362 (N_9362,N_9147,N_9033);
nor U9363 (N_9363,N_9172,N_9024);
xnor U9364 (N_9364,N_9016,N_9107);
or U9365 (N_9365,N_9038,N_9010);
nand U9366 (N_9366,N_9153,N_9029);
and U9367 (N_9367,N_9168,N_9090);
or U9368 (N_9368,N_9021,N_9061);
and U9369 (N_9369,N_9141,N_9017);
nor U9370 (N_9370,N_9006,N_9178);
or U9371 (N_9371,N_9065,N_9165);
or U9372 (N_9372,N_9166,N_9018);
nor U9373 (N_9373,N_9029,N_9183);
and U9374 (N_9374,N_9085,N_9183);
or U9375 (N_9375,N_9079,N_9148);
or U9376 (N_9376,N_9091,N_9161);
or U9377 (N_9377,N_9036,N_9147);
nor U9378 (N_9378,N_9087,N_9129);
or U9379 (N_9379,N_9085,N_9089);
nand U9380 (N_9380,N_9166,N_9146);
nand U9381 (N_9381,N_9179,N_9131);
nor U9382 (N_9382,N_9122,N_9014);
xor U9383 (N_9383,N_9108,N_9177);
and U9384 (N_9384,N_9133,N_9130);
and U9385 (N_9385,N_9184,N_9056);
xor U9386 (N_9386,N_9063,N_9023);
and U9387 (N_9387,N_9006,N_9130);
nor U9388 (N_9388,N_9161,N_9158);
xnor U9389 (N_9389,N_9187,N_9118);
nor U9390 (N_9390,N_9165,N_9103);
and U9391 (N_9391,N_9103,N_9014);
xor U9392 (N_9392,N_9178,N_9073);
nor U9393 (N_9393,N_9126,N_9165);
nor U9394 (N_9394,N_9077,N_9016);
or U9395 (N_9395,N_9192,N_9054);
nand U9396 (N_9396,N_9108,N_9003);
or U9397 (N_9397,N_9080,N_9114);
nor U9398 (N_9398,N_9062,N_9088);
and U9399 (N_9399,N_9034,N_9014);
xnor U9400 (N_9400,N_9291,N_9226);
and U9401 (N_9401,N_9247,N_9217);
or U9402 (N_9402,N_9285,N_9273);
nand U9403 (N_9403,N_9346,N_9286);
or U9404 (N_9404,N_9296,N_9207);
nor U9405 (N_9405,N_9342,N_9210);
nor U9406 (N_9406,N_9324,N_9330);
xor U9407 (N_9407,N_9303,N_9382);
xor U9408 (N_9408,N_9201,N_9253);
nor U9409 (N_9409,N_9227,N_9368);
and U9410 (N_9410,N_9350,N_9343);
or U9411 (N_9411,N_9397,N_9388);
and U9412 (N_9412,N_9381,N_9352);
or U9413 (N_9413,N_9244,N_9275);
xnor U9414 (N_9414,N_9386,N_9311);
nand U9415 (N_9415,N_9357,N_9264);
xnor U9416 (N_9416,N_9345,N_9336);
or U9417 (N_9417,N_9220,N_9265);
nor U9418 (N_9418,N_9304,N_9281);
nor U9419 (N_9419,N_9295,N_9231);
xor U9420 (N_9420,N_9234,N_9325);
xnor U9421 (N_9421,N_9338,N_9351);
and U9422 (N_9422,N_9211,N_9334);
nand U9423 (N_9423,N_9242,N_9322);
nor U9424 (N_9424,N_9384,N_9378);
or U9425 (N_9425,N_9307,N_9259);
nand U9426 (N_9426,N_9312,N_9288);
nor U9427 (N_9427,N_9235,N_9233);
xnor U9428 (N_9428,N_9380,N_9299);
and U9429 (N_9429,N_9245,N_9329);
nor U9430 (N_9430,N_9251,N_9208);
and U9431 (N_9431,N_9365,N_9374);
xor U9432 (N_9432,N_9373,N_9387);
or U9433 (N_9433,N_9315,N_9331);
nand U9434 (N_9434,N_9375,N_9367);
xnor U9435 (N_9435,N_9349,N_9268);
nand U9436 (N_9436,N_9277,N_9212);
xor U9437 (N_9437,N_9279,N_9293);
or U9438 (N_9438,N_9354,N_9284);
xor U9439 (N_9439,N_9355,N_9290);
and U9440 (N_9440,N_9202,N_9358);
nor U9441 (N_9441,N_9361,N_9250);
and U9442 (N_9442,N_9280,N_9230);
or U9443 (N_9443,N_9321,N_9326);
xnor U9444 (N_9444,N_9269,N_9252);
or U9445 (N_9445,N_9218,N_9364);
nor U9446 (N_9446,N_9258,N_9309);
nand U9447 (N_9447,N_9310,N_9240);
nand U9448 (N_9448,N_9254,N_9228);
and U9449 (N_9449,N_9359,N_9369);
xnor U9450 (N_9450,N_9289,N_9256);
nor U9451 (N_9451,N_9371,N_9300);
nand U9452 (N_9452,N_9249,N_9395);
or U9453 (N_9453,N_9393,N_9278);
xnor U9454 (N_9454,N_9389,N_9215);
nand U9455 (N_9455,N_9261,N_9313);
xor U9456 (N_9456,N_9246,N_9385);
nand U9457 (N_9457,N_9363,N_9379);
and U9458 (N_9458,N_9391,N_9248);
and U9459 (N_9459,N_9206,N_9216);
and U9460 (N_9460,N_9219,N_9333);
or U9461 (N_9461,N_9292,N_9238);
nor U9462 (N_9462,N_9287,N_9337);
and U9463 (N_9463,N_9276,N_9270);
xnor U9464 (N_9464,N_9294,N_9257);
and U9465 (N_9465,N_9229,N_9318);
xor U9466 (N_9466,N_9319,N_9362);
nor U9467 (N_9467,N_9377,N_9370);
xor U9468 (N_9468,N_9327,N_9271);
and U9469 (N_9469,N_9272,N_9347);
and U9470 (N_9470,N_9396,N_9306);
and U9471 (N_9471,N_9221,N_9283);
nand U9472 (N_9472,N_9232,N_9320);
or U9473 (N_9473,N_9340,N_9398);
and U9474 (N_9474,N_9353,N_9243);
or U9475 (N_9475,N_9314,N_9222);
xor U9476 (N_9476,N_9344,N_9204);
nand U9477 (N_9477,N_9332,N_9394);
or U9478 (N_9478,N_9203,N_9376);
xnor U9479 (N_9479,N_9282,N_9267);
xnor U9480 (N_9480,N_9262,N_9214);
nand U9481 (N_9481,N_9360,N_9328);
xnor U9482 (N_9482,N_9241,N_9348);
and U9483 (N_9483,N_9390,N_9225);
and U9484 (N_9484,N_9399,N_9366);
xnor U9485 (N_9485,N_9316,N_9209);
xor U9486 (N_9486,N_9213,N_9301);
xor U9487 (N_9487,N_9305,N_9205);
xnor U9488 (N_9488,N_9335,N_9274);
nand U9489 (N_9489,N_9239,N_9263);
nand U9490 (N_9490,N_9392,N_9341);
nor U9491 (N_9491,N_9308,N_9323);
xor U9492 (N_9492,N_9200,N_9237);
nor U9493 (N_9493,N_9224,N_9317);
nand U9494 (N_9494,N_9236,N_9255);
nand U9495 (N_9495,N_9223,N_9298);
or U9496 (N_9496,N_9383,N_9297);
xnor U9497 (N_9497,N_9372,N_9266);
nor U9498 (N_9498,N_9339,N_9302);
or U9499 (N_9499,N_9356,N_9260);
xor U9500 (N_9500,N_9345,N_9357);
and U9501 (N_9501,N_9254,N_9294);
xor U9502 (N_9502,N_9365,N_9380);
nor U9503 (N_9503,N_9383,N_9382);
and U9504 (N_9504,N_9250,N_9389);
nor U9505 (N_9505,N_9320,N_9362);
xnor U9506 (N_9506,N_9242,N_9365);
or U9507 (N_9507,N_9282,N_9322);
or U9508 (N_9508,N_9314,N_9385);
and U9509 (N_9509,N_9230,N_9363);
nor U9510 (N_9510,N_9333,N_9302);
nand U9511 (N_9511,N_9360,N_9247);
or U9512 (N_9512,N_9312,N_9320);
xor U9513 (N_9513,N_9267,N_9297);
and U9514 (N_9514,N_9237,N_9202);
nor U9515 (N_9515,N_9328,N_9366);
nor U9516 (N_9516,N_9396,N_9282);
or U9517 (N_9517,N_9225,N_9350);
or U9518 (N_9518,N_9217,N_9316);
nor U9519 (N_9519,N_9220,N_9300);
xor U9520 (N_9520,N_9317,N_9296);
or U9521 (N_9521,N_9237,N_9270);
or U9522 (N_9522,N_9374,N_9273);
or U9523 (N_9523,N_9346,N_9326);
nor U9524 (N_9524,N_9378,N_9203);
nor U9525 (N_9525,N_9321,N_9350);
and U9526 (N_9526,N_9352,N_9380);
nand U9527 (N_9527,N_9232,N_9205);
and U9528 (N_9528,N_9245,N_9234);
nor U9529 (N_9529,N_9217,N_9255);
nor U9530 (N_9530,N_9219,N_9340);
or U9531 (N_9531,N_9228,N_9286);
and U9532 (N_9532,N_9201,N_9234);
xor U9533 (N_9533,N_9352,N_9204);
xnor U9534 (N_9534,N_9223,N_9388);
nor U9535 (N_9535,N_9309,N_9268);
xor U9536 (N_9536,N_9361,N_9220);
nor U9537 (N_9537,N_9328,N_9321);
nand U9538 (N_9538,N_9355,N_9367);
nand U9539 (N_9539,N_9240,N_9387);
xor U9540 (N_9540,N_9236,N_9269);
nand U9541 (N_9541,N_9357,N_9243);
nor U9542 (N_9542,N_9231,N_9366);
and U9543 (N_9543,N_9284,N_9280);
or U9544 (N_9544,N_9257,N_9377);
xor U9545 (N_9545,N_9273,N_9279);
and U9546 (N_9546,N_9282,N_9299);
nor U9547 (N_9547,N_9325,N_9360);
or U9548 (N_9548,N_9352,N_9252);
nor U9549 (N_9549,N_9392,N_9229);
nand U9550 (N_9550,N_9270,N_9201);
nor U9551 (N_9551,N_9388,N_9254);
and U9552 (N_9552,N_9353,N_9312);
xor U9553 (N_9553,N_9278,N_9220);
nor U9554 (N_9554,N_9398,N_9217);
nand U9555 (N_9555,N_9336,N_9379);
nor U9556 (N_9556,N_9387,N_9316);
nor U9557 (N_9557,N_9210,N_9348);
nand U9558 (N_9558,N_9304,N_9211);
xor U9559 (N_9559,N_9263,N_9212);
nor U9560 (N_9560,N_9297,N_9351);
and U9561 (N_9561,N_9251,N_9264);
and U9562 (N_9562,N_9369,N_9373);
and U9563 (N_9563,N_9292,N_9370);
nand U9564 (N_9564,N_9379,N_9350);
or U9565 (N_9565,N_9208,N_9338);
xor U9566 (N_9566,N_9373,N_9379);
and U9567 (N_9567,N_9309,N_9284);
and U9568 (N_9568,N_9363,N_9318);
xor U9569 (N_9569,N_9265,N_9353);
xor U9570 (N_9570,N_9287,N_9309);
nor U9571 (N_9571,N_9306,N_9307);
nand U9572 (N_9572,N_9222,N_9302);
nand U9573 (N_9573,N_9334,N_9269);
and U9574 (N_9574,N_9241,N_9261);
and U9575 (N_9575,N_9272,N_9226);
xnor U9576 (N_9576,N_9317,N_9227);
and U9577 (N_9577,N_9306,N_9249);
xor U9578 (N_9578,N_9277,N_9395);
and U9579 (N_9579,N_9267,N_9235);
or U9580 (N_9580,N_9342,N_9366);
xnor U9581 (N_9581,N_9391,N_9312);
xnor U9582 (N_9582,N_9247,N_9313);
and U9583 (N_9583,N_9337,N_9261);
nor U9584 (N_9584,N_9217,N_9236);
and U9585 (N_9585,N_9387,N_9243);
and U9586 (N_9586,N_9308,N_9367);
xnor U9587 (N_9587,N_9266,N_9327);
nor U9588 (N_9588,N_9242,N_9205);
and U9589 (N_9589,N_9347,N_9262);
nand U9590 (N_9590,N_9308,N_9327);
xor U9591 (N_9591,N_9217,N_9328);
or U9592 (N_9592,N_9264,N_9383);
xnor U9593 (N_9593,N_9323,N_9225);
nor U9594 (N_9594,N_9224,N_9215);
nand U9595 (N_9595,N_9374,N_9280);
nor U9596 (N_9596,N_9250,N_9332);
nand U9597 (N_9597,N_9264,N_9387);
nor U9598 (N_9598,N_9394,N_9259);
and U9599 (N_9599,N_9311,N_9313);
or U9600 (N_9600,N_9550,N_9444);
xor U9601 (N_9601,N_9582,N_9518);
or U9602 (N_9602,N_9571,N_9457);
xnor U9603 (N_9603,N_9408,N_9525);
nand U9604 (N_9604,N_9509,N_9505);
nand U9605 (N_9605,N_9415,N_9545);
or U9606 (N_9606,N_9535,N_9506);
nor U9607 (N_9607,N_9581,N_9529);
or U9608 (N_9608,N_9416,N_9587);
nand U9609 (N_9609,N_9460,N_9423);
or U9610 (N_9610,N_9401,N_9442);
and U9611 (N_9611,N_9520,N_9407);
or U9612 (N_9612,N_9494,N_9438);
nand U9613 (N_9613,N_9548,N_9501);
nor U9614 (N_9614,N_9595,N_9483);
or U9615 (N_9615,N_9482,N_9499);
nor U9616 (N_9616,N_9452,N_9523);
and U9617 (N_9617,N_9448,N_9593);
nor U9618 (N_9618,N_9431,N_9569);
nand U9619 (N_9619,N_9576,N_9459);
xnor U9620 (N_9620,N_9488,N_9403);
or U9621 (N_9621,N_9544,N_9447);
and U9622 (N_9622,N_9429,N_9566);
nor U9623 (N_9623,N_9589,N_9539);
nor U9624 (N_9624,N_9543,N_9413);
xnor U9625 (N_9625,N_9532,N_9495);
or U9626 (N_9626,N_9585,N_9421);
and U9627 (N_9627,N_9469,N_9489);
or U9628 (N_9628,N_9575,N_9422);
xnor U9629 (N_9629,N_9528,N_9480);
and U9630 (N_9630,N_9561,N_9552);
xor U9631 (N_9631,N_9443,N_9455);
nand U9632 (N_9632,N_9484,N_9433);
nor U9633 (N_9633,N_9511,N_9445);
or U9634 (N_9634,N_9573,N_9590);
nand U9635 (N_9635,N_9538,N_9531);
xor U9636 (N_9636,N_9490,N_9425);
and U9637 (N_9637,N_9504,N_9540);
nand U9638 (N_9638,N_9512,N_9434);
nor U9639 (N_9639,N_9567,N_9412);
or U9640 (N_9640,N_9430,N_9492);
xnor U9641 (N_9641,N_9414,N_9417);
nor U9642 (N_9642,N_9473,N_9436);
nor U9643 (N_9643,N_9592,N_9537);
nand U9644 (N_9644,N_9519,N_9449);
or U9645 (N_9645,N_9534,N_9580);
or U9646 (N_9646,N_9424,N_9551);
or U9647 (N_9647,N_9405,N_9549);
xor U9648 (N_9648,N_9502,N_9439);
xnor U9649 (N_9649,N_9476,N_9564);
or U9650 (N_9650,N_9527,N_9542);
xnor U9651 (N_9651,N_9487,N_9458);
xor U9652 (N_9652,N_9541,N_9406);
and U9653 (N_9653,N_9441,N_9546);
nor U9654 (N_9654,N_9510,N_9598);
nand U9655 (N_9655,N_9554,N_9450);
xor U9656 (N_9656,N_9479,N_9594);
xor U9657 (N_9657,N_9474,N_9461);
xor U9658 (N_9658,N_9462,N_9516);
or U9659 (N_9659,N_9517,N_9464);
xnor U9660 (N_9660,N_9477,N_9420);
and U9661 (N_9661,N_9586,N_9486);
or U9662 (N_9662,N_9596,N_9463);
xor U9663 (N_9663,N_9556,N_9579);
nor U9664 (N_9664,N_9565,N_9454);
nand U9665 (N_9665,N_9418,N_9524);
xor U9666 (N_9666,N_9599,N_9426);
xor U9667 (N_9667,N_9451,N_9456);
nand U9668 (N_9668,N_9428,N_9491);
xnor U9669 (N_9669,N_9478,N_9533);
or U9670 (N_9670,N_9470,N_9446);
nor U9671 (N_9671,N_9588,N_9526);
or U9672 (N_9672,N_9513,N_9583);
nand U9673 (N_9673,N_9467,N_9570);
or U9674 (N_9674,N_9591,N_9568);
or U9675 (N_9675,N_9503,N_9555);
and U9676 (N_9676,N_9496,N_9562);
xor U9677 (N_9677,N_9522,N_9572);
nor U9678 (N_9678,N_9559,N_9465);
nor U9679 (N_9679,N_9475,N_9497);
nand U9680 (N_9680,N_9507,N_9500);
or U9681 (N_9681,N_9493,N_9563);
nand U9682 (N_9682,N_9560,N_9409);
nor U9683 (N_9683,N_9410,N_9597);
or U9684 (N_9684,N_9419,N_9547);
or U9685 (N_9685,N_9558,N_9432);
nor U9686 (N_9686,N_9481,N_9468);
and U9687 (N_9687,N_9440,N_9577);
nor U9688 (N_9688,N_9435,N_9485);
nand U9689 (N_9689,N_9536,N_9530);
and U9690 (N_9690,N_9521,N_9578);
nand U9691 (N_9691,N_9553,N_9400);
xor U9692 (N_9692,N_9472,N_9466);
and U9693 (N_9693,N_9471,N_9515);
and U9694 (N_9694,N_9514,N_9498);
nor U9695 (N_9695,N_9574,N_9584);
xor U9696 (N_9696,N_9411,N_9453);
or U9697 (N_9697,N_9437,N_9557);
nor U9698 (N_9698,N_9404,N_9508);
xor U9699 (N_9699,N_9427,N_9402);
or U9700 (N_9700,N_9538,N_9444);
nand U9701 (N_9701,N_9424,N_9514);
xnor U9702 (N_9702,N_9499,N_9587);
xor U9703 (N_9703,N_9552,N_9472);
and U9704 (N_9704,N_9539,N_9408);
nor U9705 (N_9705,N_9533,N_9474);
or U9706 (N_9706,N_9587,N_9590);
or U9707 (N_9707,N_9570,N_9517);
xor U9708 (N_9708,N_9494,N_9470);
nand U9709 (N_9709,N_9565,N_9420);
xor U9710 (N_9710,N_9568,N_9546);
xor U9711 (N_9711,N_9515,N_9484);
or U9712 (N_9712,N_9464,N_9571);
and U9713 (N_9713,N_9454,N_9564);
nand U9714 (N_9714,N_9439,N_9550);
nand U9715 (N_9715,N_9457,N_9533);
nand U9716 (N_9716,N_9519,N_9566);
or U9717 (N_9717,N_9493,N_9515);
nor U9718 (N_9718,N_9598,N_9579);
and U9719 (N_9719,N_9502,N_9464);
and U9720 (N_9720,N_9588,N_9540);
xor U9721 (N_9721,N_9521,N_9510);
and U9722 (N_9722,N_9424,N_9491);
xnor U9723 (N_9723,N_9460,N_9455);
or U9724 (N_9724,N_9538,N_9518);
xor U9725 (N_9725,N_9555,N_9435);
xor U9726 (N_9726,N_9471,N_9582);
nor U9727 (N_9727,N_9563,N_9593);
xor U9728 (N_9728,N_9420,N_9460);
and U9729 (N_9729,N_9541,N_9559);
and U9730 (N_9730,N_9596,N_9598);
and U9731 (N_9731,N_9495,N_9401);
or U9732 (N_9732,N_9496,N_9449);
or U9733 (N_9733,N_9553,N_9430);
and U9734 (N_9734,N_9494,N_9479);
and U9735 (N_9735,N_9455,N_9478);
nand U9736 (N_9736,N_9587,N_9476);
and U9737 (N_9737,N_9501,N_9566);
and U9738 (N_9738,N_9420,N_9436);
and U9739 (N_9739,N_9443,N_9417);
nand U9740 (N_9740,N_9446,N_9406);
and U9741 (N_9741,N_9415,N_9553);
and U9742 (N_9742,N_9548,N_9566);
nand U9743 (N_9743,N_9547,N_9450);
and U9744 (N_9744,N_9465,N_9484);
and U9745 (N_9745,N_9436,N_9490);
and U9746 (N_9746,N_9507,N_9497);
xor U9747 (N_9747,N_9597,N_9599);
nor U9748 (N_9748,N_9586,N_9545);
or U9749 (N_9749,N_9512,N_9440);
nor U9750 (N_9750,N_9440,N_9528);
nor U9751 (N_9751,N_9465,N_9418);
or U9752 (N_9752,N_9576,N_9550);
nor U9753 (N_9753,N_9467,N_9535);
nor U9754 (N_9754,N_9431,N_9415);
and U9755 (N_9755,N_9407,N_9550);
and U9756 (N_9756,N_9451,N_9426);
nand U9757 (N_9757,N_9554,N_9503);
nor U9758 (N_9758,N_9480,N_9518);
xor U9759 (N_9759,N_9415,N_9493);
nor U9760 (N_9760,N_9507,N_9572);
and U9761 (N_9761,N_9504,N_9572);
nand U9762 (N_9762,N_9489,N_9455);
xnor U9763 (N_9763,N_9407,N_9439);
nand U9764 (N_9764,N_9561,N_9521);
nor U9765 (N_9765,N_9560,N_9452);
xor U9766 (N_9766,N_9592,N_9443);
nor U9767 (N_9767,N_9452,N_9591);
nor U9768 (N_9768,N_9400,N_9417);
nor U9769 (N_9769,N_9555,N_9408);
and U9770 (N_9770,N_9512,N_9511);
nor U9771 (N_9771,N_9596,N_9486);
xnor U9772 (N_9772,N_9459,N_9454);
and U9773 (N_9773,N_9466,N_9521);
or U9774 (N_9774,N_9535,N_9438);
nand U9775 (N_9775,N_9524,N_9498);
xnor U9776 (N_9776,N_9484,N_9532);
and U9777 (N_9777,N_9589,N_9576);
nor U9778 (N_9778,N_9511,N_9531);
or U9779 (N_9779,N_9553,N_9404);
or U9780 (N_9780,N_9409,N_9479);
xnor U9781 (N_9781,N_9511,N_9488);
nand U9782 (N_9782,N_9523,N_9543);
and U9783 (N_9783,N_9547,N_9519);
xor U9784 (N_9784,N_9493,N_9492);
and U9785 (N_9785,N_9535,N_9574);
and U9786 (N_9786,N_9404,N_9535);
and U9787 (N_9787,N_9486,N_9434);
nor U9788 (N_9788,N_9507,N_9416);
nor U9789 (N_9789,N_9444,N_9592);
nand U9790 (N_9790,N_9579,N_9471);
xnor U9791 (N_9791,N_9568,N_9421);
xor U9792 (N_9792,N_9416,N_9464);
or U9793 (N_9793,N_9591,N_9558);
and U9794 (N_9794,N_9466,N_9523);
xnor U9795 (N_9795,N_9585,N_9482);
xor U9796 (N_9796,N_9545,N_9576);
or U9797 (N_9797,N_9425,N_9450);
or U9798 (N_9798,N_9445,N_9489);
nor U9799 (N_9799,N_9425,N_9512);
or U9800 (N_9800,N_9620,N_9713);
xnor U9801 (N_9801,N_9730,N_9787);
nand U9802 (N_9802,N_9652,N_9641);
xor U9803 (N_9803,N_9741,N_9695);
and U9804 (N_9804,N_9720,N_9698);
or U9805 (N_9805,N_9607,N_9601);
or U9806 (N_9806,N_9674,N_9666);
nand U9807 (N_9807,N_9765,N_9625);
xor U9808 (N_9808,N_9746,N_9776);
xor U9809 (N_9809,N_9661,N_9703);
nor U9810 (N_9810,N_9604,N_9690);
or U9811 (N_9811,N_9667,N_9657);
nor U9812 (N_9812,N_9788,N_9617);
or U9813 (N_9813,N_9634,N_9760);
xnor U9814 (N_9814,N_9767,N_9649);
xnor U9815 (N_9815,N_9688,N_9736);
nand U9816 (N_9816,N_9626,N_9790);
nor U9817 (N_9817,N_9792,N_9648);
or U9818 (N_9818,N_9615,N_9753);
nor U9819 (N_9819,N_9723,N_9785);
nand U9820 (N_9820,N_9750,N_9619);
nand U9821 (N_9821,N_9766,N_9752);
and U9822 (N_9822,N_9778,N_9722);
xnor U9823 (N_9823,N_9799,N_9739);
nand U9824 (N_9824,N_9731,N_9671);
xnor U9825 (N_9825,N_9654,N_9629);
nand U9826 (N_9826,N_9784,N_9635);
and U9827 (N_9827,N_9623,N_9775);
nor U9828 (N_9828,N_9795,N_9691);
nor U9829 (N_9829,N_9611,N_9725);
or U9830 (N_9830,N_9718,N_9763);
and U9831 (N_9831,N_9793,N_9791);
xnor U9832 (N_9832,N_9737,N_9719);
nor U9833 (N_9833,N_9733,N_9678);
and U9834 (N_9834,N_9675,N_9662);
nand U9835 (N_9835,N_9773,N_9774);
xor U9836 (N_9836,N_9780,N_9747);
and U9837 (N_9837,N_9697,N_9624);
xor U9838 (N_9838,N_9660,N_9743);
xnor U9839 (N_9839,N_9646,N_9779);
or U9840 (N_9840,N_9632,N_9764);
and U9841 (N_9841,N_9679,N_9770);
nor U9842 (N_9842,N_9762,N_9717);
and U9843 (N_9843,N_9603,N_9644);
and U9844 (N_9844,N_9769,N_9682);
or U9845 (N_9845,N_9658,N_9714);
nor U9846 (N_9846,N_9702,N_9668);
nand U9847 (N_9847,N_9716,N_9721);
nand U9848 (N_9848,N_9692,N_9751);
and U9849 (N_9849,N_9676,N_9664);
nor U9850 (N_9850,N_9724,N_9732);
xnor U9851 (N_9851,N_9712,N_9687);
or U9852 (N_9852,N_9602,N_9783);
and U9853 (N_9853,N_9758,N_9735);
or U9854 (N_9854,N_9655,N_9631);
and U9855 (N_9855,N_9663,N_9689);
and U9856 (N_9856,N_9618,N_9748);
nand U9857 (N_9857,N_9630,N_9777);
or U9858 (N_9858,N_9613,N_9772);
xor U9859 (N_9859,N_9627,N_9707);
nand U9860 (N_9860,N_9606,N_9786);
nand U9861 (N_9861,N_9756,N_9693);
or U9862 (N_9862,N_9709,N_9705);
nand U9863 (N_9863,N_9636,N_9706);
nor U9864 (N_9864,N_9639,N_9609);
xor U9865 (N_9865,N_9757,N_9659);
or U9866 (N_9866,N_9768,N_9734);
nor U9867 (N_9867,N_9794,N_9789);
nand U9868 (N_9868,N_9740,N_9638);
xor U9869 (N_9869,N_9651,N_9650);
nand U9870 (N_9870,N_9621,N_9643);
nor U9871 (N_9871,N_9642,N_9633);
nor U9872 (N_9872,N_9686,N_9680);
nor U9873 (N_9873,N_9653,N_9749);
nor U9874 (N_9874,N_9665,N_9628);
and U9875 (N_9875,N_9670,N_9610);
nor U9876 (N_9876,N_9711,N_9685);
nand U9877 (N_9877,N_9781,N_9647);
nor U9878 (N_9878,N_9672,N_9726);
nand U9879 (N_9879,N_9605,N_9640);
nor U9880 (N_9880,N_9738,N_9656);
nand U9881 (N_9881,N_9759,N_9754);
xor U9882 (N_9882,N_9699,N_9616);
xor U9883 (N_9883,N_9798,N_9694);
and U9884 (N_9884,N_9710,N_9600);
or U9885 (N_9885,N_9701,N_9745);
and U9886 (N_9886,N_9728,N_9727);
and U9887 (N_9887,N_9622,N_9700);
or U9888 (N_9888,N_9797,N_9771);
nand U9889 (N_9889,N_9729,N_9608);
and U9890 (N_9890,N_9673,N_9645);
or U9891 (N_9891,N_9612,N_9696);
or U9892 (N_9892,N_9782,N_9708);
xnor U9893 (N_9893,N_9683,N_9744);
nor U9894 (N_9894,N_9677,N_9614);
nand U9895 (N_9895,N_9796,N_9755);
nor U9896 (N_9896,N_9704,N_9684);
xnor U9897 (N_9897,N_9742,N_9637);
xor U9898 (N_9898,N_9669,N_9681);
nor U9899 (N_9899,N_9715,N_9761);
xnor U9900 (N_9900,N_9728,N_9760);
or U9901 (N_9901,N_9795,N_9792);
xor U9902 (N_9902,N_9782,N_9704);
nor U9903 (N_9903,N_9793,N_9708);
or U9904 (N_9904,N_9730,N_9611);
and U9905 (N_9905,N_9664,N_9756);
or U9906 (N_9906,N_9710,N_9790);
and U9907 (N_9907,N_9649,N_9790);
or U9908 (N_9908,N_9631,N_9729);
and U9909 (N_9909,N_9687,N_9731);
or U9910 (N_9910,N_9710,N_9777);
nand U9911 (N_9911,N_9764,N_9661);
nand U9912 (N_9912,N_9767,N_9786);
nand U9913 (N_9913,N_9749,N_9752);
nand U9914 (N_9914,N_9736,N_9713);
and U9915 (N_9915,N_9793,N_9674);
or U9916 (N_9916,N_9707,N_9613);
and U9917 (N_9917,N_9739,N_9753);
and U9918 (N_9918,N_9605,N_9728);
nor U9919 (N_9919,N_9698,N_9675);
xor U9920 (N_9920,N_9618,N_9658);
nor U9921 (N_9921,N_9653,N_9704);
xnor U9922 (N_9922,N_9775,N_9705);
and U9923 (N_9923,N_9697,N_9705);
nand U9924 (N_9924,N_9777,N_9644);
nor U9925 (N_9925,N_9646,N_9756);
nand U9926 (N_9926,N_9747,N_9711);
nor U9927 (N_9927,N_9645,N_9717);
or U9928 (N_9928,N_9653,N_9606);
xor U9929 (N_9929,N_9679,N_9749);
xnor U9930 (N_9930,N_9670,N_9673);
nand U9931 (N_9931,N_9705,N_9778);
or U9932 (N_9932,N_9657,N_9709);
nor U9933 (N_9933,N_9784,N_9659);
and U9934 (N_9934,N_9759,N_9725);
xnor U9935 (N_9935,N_9685,N_9668);
or U9936 (N_9936,N_9637,N_9641);
or U9937 (N_9937,N_9739,N_9622);
nand U9938 (N_9938,N_9737,N_9672);
nor U9939 (N_9939,N_9791,N_9677);
and U9940 (N_9940,N_9619,N_9602);
nand U9941 (N_9941,N_9688,N_9649);
or U9942 (N_9942,N_9603,N_9627);
nor U9943 (N_9943,N_9757,N_9619);
nand U9944 (N_9944,N_9677,N_9698);
nor U9945 (N_9945,N_9623,N_9648);
xor U9946 (N_9946,N_9659,N_9652);
xnor U9947 (N_9947,N_9732,N_9606);
xnor U9948 (N_9948,N_9678,N_9601);
xor U9949 (N_9949,N_9717,N_9625);
nor U9950 (N_9950,N_9785,N_9614);
or U9951 (N_9951,N_9748,N_9729);
xnor U9952 (N_9952,N_9779,N_9760);
xor U9953 (N_9953,N_9604,N_9686);
and U9954 (N_9954,N_9694,N_9642);
or U9955 (N_9955,N_9634,N_9618);
nor U9956 (N_9956,N_9610,N_9611);
nor U9957 (N_9957,N_9718,N_9656);
and U9958 (N_9958,N_9779,N_9690);
nand U9959 (N_9959,N_9731,N_9666);
xor U9960 (N_9960,N_9736,N_9768);
nand U9961 (N_9961,N_9732,N_9665);
and U9962 (N_9962,N_9693,N_9645);
xnor U9963 (N_9963,N_9680,N_9720);
and U9964 (N_9964,N_9706,N_9769);
xnor U9965 (N_9965,N_9612,N_9734);
xor U9966 (N_9966,N_9658,N_9764);
and U9967 (N_9967,N_9755,N_9683);
and U9968 (N_9968,N_9730,N_9623);
or U9969 (N_9969,N_9736,N_9694);
and U9970 (N_9970,N_9660,N_9731);
nand U9971 (N_9971,N_9776,N_9781);
and U9972 (N_9972,N_9767,N_9741);
and U9973 (N_9973,N_9638,N_9610);
xor U9974 (N_9974,N_9717,N_9679);
xor U9975 (N_9975,N_9775,N_9659);
xnor U9976 (N_9976,N_9699,N_9745);
and U9977 (N_9977,N_9675,N_9712);
or U9978 (N_9978,N_9703,N_9744);
nor U9979 (N_9979,N_9646,N_9715);
or U9980 (N_9980,N_9724,N_9664);
nor U9981 (N_9981,N_9783,N_9611);
or U9982 (N_9982,N_9792,N_9757);
and U9983 (N_9983,N_9783,N_9799);
and U9984 (N_9984,N_9754,N_9718);
xnor U9985 (N_9985,N_9685,N_9655);
nor U9986 (N_9986,N_9641,N_9666);
nand U9987 (N_9987,N_9618,N_9734);
and U9988 (N_9988,N_9771,N_9620);
or U9989 (N_9989,N_9660,N_9777);
and U9990 (N_9990,N_9748,N_9755);
nand U9991 (N_9991,N_9649,N_9709);
and U9992 (N_9992,N_9743,N_9670);
or U9993 (N_9993,N_9600,N_9661);
and U9994 (N_9994,N_9662,N_9786);
or U9995 (N_9995,N_9622,N_9788);
nor U9996 (N_9996,N_9698,N_9628);
and U9997 (N_9997,N_9603,N_9657);
and U9998 (N_9998,N_9633,N_9767);
and U9999 (N_9999,N_9773,N_9678);
xor U10000 (N_10000,N_9921,N_9954);
nand U10001 (N_10001,N_9953,N_9805);
xor U10002 (N_10002,N_9996,N_9935);
and U10003 (N_10003,N_9880,N_9861);
or U10004 (N_10004,N_9997,N_9899);
nor U10005 (N_10005,N_9906,N_9922);
and U10006 (N_10006,N_9867,N_9943);
xor U10007 (N_10007,N_9856,N_9853);
or U10008 (N_10008,N_9901,N_9854);
nand U10009 (N_10009,N_9957,N_9893);
nor U10010 (N_10010,N_9987,N_9814);
and U10011 (N_10011,N_9855,N_9982);
nand U10012 (N_10012,N_9864,N_9990);
and U10013 (N_10013,N_9846,N_9995);
and U10014 (N_10014,N_9972,N_9938);
and U10015 (N_10015,N_9986,N_9916);
or U10016 (N_10016,N_9947,N_9807);
xnor U10017 (N_10017,N_9844,N_9877);
or U10018 (N_10018,N_9845,N_9925);
and U10019 (N_10019,N_9840,N_9847);
nand U10020 (N_10020,N_9865,N_9993);
xnor U10021 (N_10021,N_9822,N_9800);
nor U10022 (N_10022,N_9891,N_9961);
nand U10023 (N_10023,N_9904,N_9929);
nor U10024 (N_10024,N_9831,N_9971);
xnor U10025 (N_10025,N_9875,N_9905);
nor U10026 (N_10026,N_9923,N_9978);
xnor U10027 (N_10027,N_9991,N_9803);
or U10028 (N_10028,N_9888,N_9895);
and U10029 (N_10029,N_9983,N_9956);
nor U10030 (N_10030,N_9999,N_9825);
nand U10031 (N_10031,N_9886,N_9898);
nor U10032 (N_10032,N_9850,N_9866);
xor U10033 (N_10033,N_9962,N_9900);
nor U10034 (N_10034,N_9832,N_9911);
or U10035 (N_10035,N_9830,N_9964);
and U10036 (N_10036,N_9824,N_9835);
nand U10037 (N_10037,N_9812,N_9909);
or U10038 (N_10038,N_9931,N_9810);
nand U10039 (N_10039,N_9811,N_9950);
or U10040 (N_10040,N_9939,N_9809);
xnor U10041 (N_10041,N_9903,N_9843);
or U10042 (N_10042,N_9801,N_9963);
nand U10043 (N_10043,N_9883,N_9976);
nor U10044 (N_10044,N_9827,N_9873);
nor U10045 (N_10045,N_9839,N_9979);
nand U10046 (N_10046,N_9826,N_9858);
or U10047 (N_10047,N_9970,N_9913);
and U10048 (N_10048,N_9896,N_9892);
or U10049 (N_10049,N_9946,N_9992);
xor U10050 (N_10050,N_9889,N_9940);
nor U10051 (N_10051,N_9818,N_9802);
nand U10052 (N_10052,N_9879,N_9980);
or U10053 (N_10053,N_9823,N_9942);
xor U10054 (N_10054,N_9819,N_9887);
or U10055 (N_10055,N_9915,N_9908);
xor U10056 (N_10056,N_9833,N_9977);
or U10057 (N_10057,N_9876,N_9828);
xor U10058 (N_10058,N_9981,N_9933);
and U10059 (N_10059,N_9842,N_9816);
xnor U10060 (N_10060,N_9837,N_9907);
or U10061 (N_10061,N_9967,N_9872);
and U10062 (N_10062,N_9984,N_9804);
and U10063 (N_10063,N_9949,N_9863);
xor U10064 (N_10064,N_9817,N_9930);
nand U10065 (N_10065,N_9926,N_9958);
xnor U10066 (N_10066,N_9945,N_9838);
nand U10067 (N_10067,N_9918,N_9894);
xnor U10068 (N_10068,N_9955,N_9815);
nand U10069 (N_10069,N_9914,N_9968);
nand U10070 (N_10070,N_9820,N_9937);
or U10071 (N_10071,N_9920,N_9927);
or U10072 (N_10072,N_9897,N_9878);
and U10073 (N_10073,N_9944,N_9951);
xnor U10074 (N_10074,N_9910,N_9969);
nand U10075 (N_10075,N_9989,N_9821);
or U10076 (N_10076,N_9934,N_9870);
xor U10077 (N_10077,N_9860,N_9902);
or U10078 (N_10078,N_9912,N_9919);
or U10079 (N_10079,N_9834,N_9868);
xnor U10080 (N_10080,N_9885,N_9952);
nand U10081 (N_10081,N_9924,N_9973);
and U10082 (N_10082,N_9917,N_9975);
and U10083 (N_10083,N_9859,N_9932);
or U10084 (N_10084,N_9848,N_9959);
xor U10085 (N_10085,N_9974,N_9836);
or U10086 (N_10086,N_9849,N_9985);
nand U10087 (N_10087,N_9936,N_9882);
or U10088 (N_10088,N_9881,N_9806);
xor U10089 (N_10089,N_9994,N_9808);
nor U10090 (N_10090,N_9890,N_9948);
nor U10091 (N_10091,N_9965,N_9871);
or U10092 (N_10092,N_9998,N_9852);
xor U10093 (N_10093,N_9884,N_9960);
xor U10094 (N_10094,N_9857,N_9851);
xnor U10095 (N_10095,N_9869,N_9829);
and U10096 (N_10096,N_9941,N_9928);
nor U10097 (N_10097,N_9862,N_9966);
nor U10098 (N_10098,N_9988,N_9874);
nor U10099 (N_10099,N_9841,N_9813);
xor U10100 (N_10100,N_9847,N_9994);
or U10101 (N_10101,N_9964,N_9844);
or U10102 (N_10102,N_9924,N_9813);
xnor U10103 (N_10103,N_9944,N_9960);
nand U10104 (N_10104,N_9964,N_9961);
nor U10105 (N_10105,N_9963,N_9879);
and U10106 (N_10106,N_9893,N_9917);
or U10107 (N_10107,N_9896,N_9936);
or U10108 (N_10108,N_9856,N_9958);
xnor U10109 (N_10109,N_9872,N_9886);
or U10110 (N_10110,N_9915,N_9828);
nor U10111 (N_10111,N_9946,N_9808);
or U10112 (N_10112,N_9816,N_9904);
and U10113 (N_10113,N_9889,N_9914);
and U10114 (N_10114,N_9838,N_9997);
nor U10115 (N_10115,N_9889,N_9920);
or U10116 (N_10116,N_9955,N_9981);
or U10117 (N_10117,N_9861,N_9866);
or U10118 (N_10118,N_9971,N_9984);
xnor U10119 (N_10119,N_9872,N_9800);
nand U10120 (N_10120,N_9915,N_9963);
or U10121 (N_10121,N_9843,N_9874);
or U10122 (N_10122,N_9829,N_9940);
nor U10123 (N_10123,N_9935,N_9933);
nand U10124 (N_10124,N_9953,N_9906);
and U10125 (N_10125,N_9954,N_9891);
or U10126 (N_10126,N_9897,N_9882);
nand U10127 (N_10127,N_9851,N_9916);
nand U10128 (N_10128,N_9983,N_9905);
nand U10129 (N_10129,N_9955,N_9836);
or U10130 (N_10130,N_9869,N_9958);
nor U10131 (N_10131,N_9920,N_9804);
xnor U10132 (N_10132,N_9923,N_9980);
nor U10133 (N_10133,N_9963,N_9893);
nor U10134 (N_10134,N_9986,N_9998);
nand U10135 (N_10135,N_9891,N_9955);
xnor U10136 (N_10136,N_9985,N_9923);
nand U10137 (N_10137,N_9971,N_9847);
and U10138 (N_10138,N_9866,N_9999);
or U10139 (N_10139,N_9884,N_9849);
or U10140 (N_10140,N_9962,N_9803);
nor U10141 (N_10141,N_9868,N_9923);
or U10142 (N_10142,N_9937,N_9914);
xor U10143 (N_10143,N_9832,N_9863);
and U10144 (N_10144,N_9847,N_9997);
or U10145 (N_10145,N_9907,N_9872);
nand U10146 (N_10146,N_9859,N_9987);
or U10147 (N_10147,N_9988,N_9916);
or U10148 (N_10148,N_9959,N_9860);
nor U10149 (N_10149,N_9955,N_9870);
and U10150 (N_10150,N_9835,N_9906);
xor U10151 (N_10151,N_9959,N_9881);
or U10152 (N_10152,N_9936,N_9814);
or U10153 (N_10153,N_9808,N_9913);
nand U10154 (N_10154,N_9950,N_9915);
and U10155 (N_10155,N_9890,N_9862);
and U10156 (N_10156,N_9945,N_9903);
or U10157 (N_10157,N_9809,N_9865);
or U10158 (N_10158,N_9992,N_9897);
xnor U10159 (N_10159,N_9891,N_9830);
xnor U10160 (N_10160,N_9935,N_9877);
or U10161 (N_10161,N_9920,N_9850);
nor U10162 (N_10162,N_9952,N_9930);
and U10163 (N_10163,N_9881,N_9997);
nand U10164 (N_10164,N_9902,N_9873);
xnor U10165 (N_10165,N_9927,N_9939);
nand U10166 (N_10166,N_9930,N_9920);
nand U10167 (N_10167,N_9895,N_9948);
nand U10168 (N_10168,N_9964,N_9962);
nor U10169 (N_10169,N_9868,N_9969);
and U10170 (N_10170,N_9863,N_9973);
and U10171 (N_10171,N_9968,N_9943);
and U10172 (N_10172,N_9911,N_9970);
nand U10173 (N_10173,N_9897,N_9956);
nor U10174 (N_10174,N_9804,N_9827);
xor U10175 (N_10175,N_9858,N_9879);
or U10176 (N_10176,N_9935,N_9896);
nand U10177 (N_10177,N_9971,N_9989);
and U10178 (N_10178,N_9926,N_9940);
nor U10179 (N_10179,N_9984,N_9836);
nand U10180 (N_10180,N_9917,N_9964);
nor U10181 (N_10181,N_9827,N_9930);
nor U10182 (N_10182,N_9895,N_9954);
nand U10183 (N_10183,N_9931,N_9981);
and U10184 (N_10184,N_9905,N_9991);
or U10185 (N_10185,N_9887,N_9962);
nand U10186 (N_10186,N_9831,N_9870);
nand U10187 (N_10187,N_9940,N_9840);
nand U10188 (N_10188,N_9908,N_9961);
or U10189 (N_10189,N_9983,N_9927);
xor U10190 (N_10190,N_9845,N_9995);
or U10191 (N_10191,N_9890,N_9922);
or U10192 (N_10192,N_9869,N_9907);
xnor U10193 (N_10193,N_9832,N_9889);
nand U10194 (N_10194,N_9849,N_9811);
nor U10195 (N_10195,N_9853,N_9871);
and U10196 (N_10196,N_9866,N_9944);
nand U10197 (N_10197,N_9962,N_9999);
xnor U10198 (N_10198,N_9842,N_9991);
nor U10199 (N_10199,N_9815,N_9894);
or U10200 (N_10200,N_10095,N_10115);
xor U10201 (N_10201,N_10059,N_10133);
nor U10202 (N_10202,N_10039,N_10035);
nand U10203 (N_10203,N_10036,N_10171);
and U10204 (N_10204,N_10021,N_10192);
nand U10205 (N_10205,N_10110,N_10048);
and U10206 (N_10206,N_10143,N_10196);
xor U10207 (N_10207,N_10189,N_10122);
or U10208 (N_10208,N_10161,N_10108);
or U10209 (N_10209,N_10132,N_10188);
xnor U10210 (N_10210,N_10026,N_10060);
xor U10211 (N_10211,N_10064,N_10128);
or U10212 (N_10212,N_10118,N_10051);
or U10213 (N_10213,N_10104,N_10075);
nand U10214 (N_10214,N_10100,N_10163);
or U10215 (N_10215,N_10136,N_10015);
xor U10216 (N_10216,N_10151,N_10056);
xor U10217 (N_10217,N_10050,N_10065);
and U10218 (N_10218,N_10199,N_10005);
or U10219 (N_10219,N_10014,N_10010);
and U10220 (N_10220,N_10067,N_10099);
nand U10221 (N_10221,N_10022,N_10028);
nor U10222 (N_10222,N_10093,N_10089);
and U10223 (N_10223,N_10000,N_10183);
or U10224 (N_10224,N_10123,N_10125);
xor U10225 (N_10225,N_10024,N_10107);
xnor U10226 (N_10226,N_10029,N_10081);
nor U10227 (N_10227,N_10079,N_10044);
xor U10228 (N_10228,N_10087,N_10038);
or U10229 (N_10229,N_10086,N_10130);
xnor U10230 (N_10230,N_10076,N_10013);
xnor U10231 (N_10231,N_10185,N_10102);
or U10232 (N_10232,N_10194,N_10043);
xnor U10233 (N_10233,N_10154,N_10114);
xnor U10234 (N_10234,N_10146,N_10063);
nor U10235 (N_10235,N_10047,N_10178);
and U10236 (N_10236,N_10167,N_10016);
xnor U10237 (N_10237,N_10106,N_10160);
xor U10238 (N_10238,N_10082,N_10072);
nand U10239 (N_10239,N_10131,N_10141);
xnor U10240 (N_10240,N_10138,N_10037);
and U10241 (N_10241,N_10165,N_10155);
or U10242 (N_10242,N_10070,N_10144);
nor U10243 (N_10243,N_10034,N_10190);
nor U10244 (N_10244,N_10055,N_10158);
and U10245 (N_10245,N_10053,N_10049);
and U10246 (N_10246,N_10008,N_10139);
and U10247 (N_10247,N_10174,N_10083);
nor U10248 (N_10248,N_10181,N_10195);
nor U10249 (N_10249,N_10045,N_10121);
nand U10250 (N_10250,N_10069,N_10074);
xor U10251 (N_10251,N_10135,N_10071);
xnor U10252 (N_10252,N_10054,N_10162);
nor U10253 (N_10253,N_10127,N_10091);
nand U10254 (N_10254,N_10124,N_10197);
nand U10255 (N_10255,N_10169,N_10159);
nand U10256 (N_10256,N_10041,N_10078);
or U10257 (N_10257,N_10166,N_10172);
nor U10258 (N_10258,N_10182,N_10103);
xor U10259 (N_10259,N_10180,N_10033);
nand U10260 (N_10260,N_10198,N_10168);
xnor U10261 (N_10261,N_10061,N_10119);
or U10262 (N_10262,N_10134,N_10175);
nor U10263 (N_10263,N_10164,N_10062);
nand U10264 (N_10264,N_10109,N_10177);
xor U10265 (N_10265,N_10052,N_10023);
and U10266 (N_10266,N_10046,N_10187);
and U10267 (N_10267,N_10073,N_10027);
nor U10268 (N_10268,N_10006,N_10191);
xor U10269 (N_10269,N_10153,N_10184);
xnor U10270 (N_10270,N_10157,N_10032);
and U10271 (N_10271,N_10003,N_10096);
nor U10272 (N_10272,N_10085,N_10018);
or U10273 (N_10273,N_10030,N_10170);
and U10274 (N_10274,N_10092,N_10145);
and U10275 (N_10275,N_10019,N_10176);
nor U10276 (N_10276,N_10137,N_10031);
nand U10277 (N_10277,N_10001,N_10193);
and U10278 (N_10278,N_10068,N_10101);
xnor U10279 (N_10279,N_10148,N_10126);
nand U10280 (N_10280,N_10012,N_10150);
and U10281 (N_10281,N_10149,N_10088);
nand U10282 (N_10282,N_10007,N_10142);
and U10283 (N_10283,N_10097,N_10094);
or U10284 (N_10284,N_10129,N_10113);
nor U10285 (N_10285,N_10173,N_10084);
nor U10286 (N_10286,N_10098,N_10058);
xor U10287 (N_10287,N_10009,N_10042);
nand U10288 (N_10288,N_10186,N_10020);
and U10289 (N_10289,N_10117,N_10112);
and U10290 (N_10290,N_10140,N_10011);
and U10291 (N_10291,N_10057,N_10179);
nand U10292 (N_10292,N_10017,N_10120);
nor U10293 (N_10293,N_10040,N_10066);
nor U10294 (N_10294,N_10025,N_10156);
xor U10295 (N_10295,N_10147,N_10152);
xor U10296 (N_10296,N_10004,N_10080);
and U10297 (N_10297,N_10077,N_10111);
or U10298 (N_10298,N_10090,N_10002);
and U10299 (N_10299,N_10105,N_10116);
nor U10300 (N_10300,N_10004,N_10066);
or U10301 (N_10301,N_10071,N_10048);
xor U10302 (N_10302,N_10075,N_10100);
nand U10303 (N_10303,N_10143,N_10156);
nor U10304 (N_10304,N_10053,N_10008);
and U10305 (N_10305,N_10135,N_10092);
nand U10306 (N_10306,N_10063,N_10029);
xnor U10307 (N_10307,N_10095,N_10057);
nor U10308 (N_10308,N_10088,N_10005);
nand U10309 (N_10309,N_10157,N_10038);
nor U10310 (N_10310,N_10153,N_10059);
nand U10311 (N_10311,N_10054,N_10112);
nor U10312 (N_10312,N_10009,N_10169);
and U10313 (N_10313,N_10085,N_10047);
xor U10314 (N_10314,N_10026,N_10130);
nand U10315 (N_10315,N_10146,N_10021);
or U10316 (N_10316,N_10116,N_10126);
nand U10317 (N_10317,N_10028,N_10189);
nand U10318 (N_10318,N_10081,N_10052);
or U10319 (N_10319,N_10130,N_10150);
and U10320 (N_10320,N_10148,N_10099);
xnor U10321 (N_10321,N_10156,N_10089);
xor U10322 (N_10322,N_10065,N_10076);
and U10323 (N_10323,N_10092,N_10082);
and U10324 (N_10324,N_10123,N_10158);
nand U10325 (N_10325,N_10060,N_10126);
or U10326 (N_10326,N_10041,N_10008);
or U10327 (N_10327,N_10186,N_10057);
or U10328 (N_10328,N_10173,N_10184);
or U10329 (N_10329,N_10154,N_10118);
nor U10330 (N_10330,N_10051,N_10122);
nor U10331 (N_10331,N_10025,N_10068);
or U10332 (N_10332,N_10113,N_10167);
nand U10333 (N_10333,N_10074,N_10158);
nor U10334 (N_10334,N_10173,N_10090);
xor U10335 (N_10335,N_10160,N_10002);
xnor U10336 (N_10336,N_10147,N_10130);
nand U10337 (N_10337,N_10144,N_10078);
nor U10338 (N_10338,N_10025,N_10053);
nor U10339 (N_10339,N_10068,N_10112);
and U10340 (N_10340,N_10025,N_10166);
and U10341 (N_10341,N_10050,N_10168);
xor U10342 (N_10342,N_10130,N_10188);
and U10343 (N_10343,N_10171,N_10098);
and U10344 (N_10344,N_10068,N_10178);
nand U10345 (N_10345,N_10137,N_10168);
nor U10346 (N_10346,N_10013,N_10163);
xnor U10347 (N_10347,N_10180,N_10178);
xnor U10348 (N_10348,N_10106,N_10107);
nor U10349 (N_10349,N_10052,N_10180);
or U10350 (N_10350,N_10115,N_10107);
or U10351 (N_10351,N_10136,N_10135);
and U10352 (N_10352,N_10009,N_10015);
or U10353 (N_10353,N_10067,N_10183);
and U10354 (N_10354,N_10103,N_10155);
and U10355 (N_10355,N_10009,N_10183);
and U10356 (N_10356,N_10069,N_10130);
or U10357 (N_10357,N_10096,N_10121);
and U10358 (N_10358,N_10039,N_10079);
or U10359 (N_10359,N_10081,N_10103);
or U10360 (N_10360,N_10042,N_10196);
nand U10361 (N_10361,N_10017,N_10117);
nor U10362 (N_10362,N_10033,N_10053);
nor U10363 (N_10363,N_10081,N_10099);
nand U10364 (N_10364,N_10160,N_10183);
nand U10365 (N_10365,N_10167,N_10150);
nor U10366 (N_10366,N_10198,N_10152);
nor U10367 (N_10367,N_10145,N_10098);
nor U10368 (N_10368,N_10086,N_10016);
xnor U10369 (N_10369,N_10182,N_10099);
xor U10370 (N_10370,N_10107,N_10005);
nor U10371 (N_10371,N_10109,N_10143);
and U10372 (N_10372,N_10199,N_10168);
or U10373 (N_10373,N_10130,N_10035);
and U10374 (N_10374,N_10095,N_10060);
or U10375 (N_10375,N_10136,N_10081);
xor U10376 (N_10376,N_10005,N_10153);
xnor U10377 (N_10377,N_10035,N_10099);
and U10378 (N_10378,N_10045,N_10120);
nor U10379 (N_10379,N_10039,N_10136);
and U10380 (N_10380,N_10142,N_10073);
or U10381 (N_10381,N_10129,N_10091);
xor U10382 (N_10382,N_10122,N_10026);
xor U10383 (N_10383,N_10103,N_10102);
and U10384 (N_10384,N_10005,N_10029);
and U10385 (N_10385,N_10084,N_10190);
or U10386 (N_10386,N_10085,N_10067);
and U10387 (N_10387,N_10082,N_10111);
and U10388 (N_10388,N_10044,N_10180);
nand U10389 (N_10389,N_10034,N_10024);
nand U10390 (N_10390,N_10176,N_10077);
and U10391 (N_10391,N_10105,N_10049);
nand U10392 (N_10392,N_10148,N_10004);
and U10393 (N_10393,N_10065,N_10166);
nor U10394 (N_10394,N_10123,N_10131);
or U10395 (N_10395,N_10036,N_10119);
xnor U10396 (N_10396,N_10004,N_10160);
and U10397 (N_10397,N_10040,N_10195);
nand U10398 (N_10398,N_10196,N_10127);
or U10399 (N_10399,N_10083,N_10149);
and U10400 (N_10400,N_10258,N_10318);
nor U10401 (N_10401,N_10380,N_10296);
nand U10402 (N_10402,N_10328,N_10275);
nor U10403 (N_10403,N_10280,N_10322);
nand U10404 (N_10404,N_10357,N_10289);
or U10405 (N_10405,N_10383,N_10387);
or U10406 (N_10406,N_10259,N_10268);
nand U10407 (N_10407,N_10202,N_10292);
nand U10408 (N_10408,N_10338,N_10270);
and U10409 (N_10409,N_10320,N_10364);
and U10410 (N_10410,N_10267,N_10245);
and U10411 (N_10411,N_10260,N_10234);
and U10412 (N_10412,N_10251,N_10290);
or U10413 (N_10413,N_10395,N_10355);
xor U10414 (N_10414,N_10365,N_10264);
nand U10415 (N_10415,N_10212,N_10216);
nor U10416 (N_10416,N_10236,N_10210);
or U10417 (N_10417,N_10237,N_10229);
nand U10418 (N_10418,N_10315,N_10223);
nand U10419 (N_10419,N_10266,N_10217);
nand U10420 (N_10420,N_10325,N_10220);
and U10421 (N_10421,N_10363,N_10324);
nand U10422 (N_10422,N_10254,N_10329);
or U10423 (N_10423,N_10358,N_10333);
and U10424 (N_10424,N_10398,N_10389);
nand U10425 (N_10425,N_10359,N_10263);
nor U10426 (N_10426,N_10386,N_10310);
and U10427 (N_10427,N_10213,N_10265);
nand U10428 (N_10428,N_10271,N_10201);
or U10429 (N_10429,N_10283,N_10313);
xor U10430 (N_10430,N_10255,N_10397);
nand U10431 (N_10431,N_10346,N_10238);
xor U10432 (N_10432,N_10285,N_10227);
nand U10433 (N_10433,N_10391,N_10312);
nor U10434 (N_10434,N_10208,N_10399);
nor U10435 (N_10435,N_10350,N_10360);
xor U10436 (N_10436,N_10301,N_10392);
nor U10437 (N_10437,N_10240,N_10294);
or U10438 (N_10438,N_10337,N_10252);
or U10439 (N_10439,N_10330,N_10393);
and U10440 (N_10440,N_10343,N_10345);
xnor U10441 (N_10441,N_10336,N_10394);
nand U10442 (N_10442,N_10204,N_10390);
or U10443 (N_10443,N_10256,N_10369);
and U10444 (N_10444,N_10250,N_10308);
or U10445 (N_10445,N_10287,N_10299);
xor U10446 (N_10446,N_10249,N_10306);
nor U10447 (N_10447,N_10243,N_10278);
nand U10448 (N_10448,N_10311,N_10370);
or U10449 (N_10449,N_10262,N_10281);
and U10450 (N_10450,N_10362,N_10206);
and U10451 (N_10451,N_10203,N_10261);
xnor U10452 (N_10452,N_10317,N_10348);
nor U10453 (N_10453,N_10344,N_10339);
and U10454 (N_10454,N_10366,N_10335);
nor U10455 (N_10455,N_10309,N_10274);
and U10456 (N_10456,N_10342,N_10307);
nand U10457 (N_10457,N_10233,N_10209);
nor U10458 (N_10458,N_10303,N_10298);
or U10459 (N_10459,N_10372,N_10305);
and U10460 (N_10460,N_10327,N_10211);
nor U10461 (N_10461,N_10205,N_10269);
xnor U10462 (N_10462,N_10291,N_10257);
nor U10463 (N_10463,N_10377,N_10323);
nand U10464 (N_10464,N_10378,N_10331);
nor U10465 (N_10465,N_10297,N_10379);
nor U10466 (N_10466,N_10279,N_10215);
xor U10467 (N_10467,N_10207,N_10241);
xor U10468 (N_10468,N_10321,N_10341);
xnor U10469 (N_10469,N_10288,N_10225);
and U10470 (N_10470,N_10230,N_10224);
nand U10471 (N_10471,N_10352,N_10218);
xnor U10472 (N_10472,N_10228,N_10214);
nand U10473 (N_10473,N_10239,N_10248);
nand U10474 (N_10474,N_10232,N_10367);
and U10475 (N_10475,N_10226,N_10242);
and U10476 (N_10476,N_10276,N_10382);
or U10477 (N_10477,N_10200,N_10361);
and U10478 (N_10478,N_10231,N_10347);
nor U10479 (N_10479,N_10374,N_10284);
and U10480 (N_10480,N_10272,N_10385);
nor U10481 (N_10481,N_10277,N_10273);
xnor U10482 (N_10482,N_10302,N_10247);
xor U10483 (N_10483,N_10396,N_10221);
xnor U10484 (N_10484,N_10295,N_10246);
nor U10485 (N_10485,N_10326,N_10222);
nor U10486 (N_10486,N_10381,N_10219);
or U10487 (N_10487,N_10253,N_10244);
nor U10488 (N_10488,N_10368,N_10353);
nand U10489 (N_10489,N_10384,N_10373);
and U10490 (N_10490,N_10332,N_10235);
and U10491 (N_10491,N_10340,N_10351);
nor U10492 (N_10492,N_10376,N_10349);
and U10493 (N_10493,N_10388,N_10356);
and U10494 (N_10494,N_10282,N_10286);
nand U10495 (N_10495,N_10319,N_10300);
xnor U10496 (N_10496,N_10375,N_10314);
nor U10497 (N_10497,N_10293,N_10316);
nor U10498 (N_10498,N_10304,N_10354);
or U10499 (N_10499,N_10371,N_10334);
nand U10500 (N_10500,N_10326,N_10383);
nand U10501 (N_10501,N_10355,N_10383);
nor U10502 (N_10502,N_10210,N_10320);
xnor U10503 (N_10503,N_10392,N_10276);
nand U10504 (N_10504,N_10349,N_10358);
nand U10505 (N_10505,N_10273,N_10358);
or U10506 (N_10506,N_10231,N_10250);
or U10507 (N_10507,N_10243,N_10372);
and U10508 (N_10508,N_10315,N_10217);
xor U10509 (N_10509,N_10383,N_10200);
and U10510 (N_10510,N_10204,N_10229);
or U10511 (N_10511,N_10302,N_10255);
and U10512 (N_10512,N_10328,N_10288);
or U10513 (N_10513,N_10221,N_10227);
nor U10514 (N_10514,N_10208,N_10271);
nand U10515 (N_10515,N_10378,N_10367);
xor U10516 (N_10516,N_10381,N_10358);
nand U10517 (N_10517,N_10358,N_10306);
nand U10518 (N_10518,N_10300,N_10213);
and U10519 (N_10519,N_10376,N_10273);
xnor U10520 (N_10520,N_10243,N_10399);
and U10521 (N_10521,N_10302,N_10385);
and U10522 (N_10522,N_10308,N_10278);
xor U10523 (N_10523,N_10347,N_10249);
or U10524 (N_10524,N_10203,N_10240);
or U10525 (N_10525,N_10372,N_10212);
nor U10526 (N_10526,N_10200,N_10229);
or U10527 (N_10527,N_10244,N_10389);
nor U10528 (N_10528,N_10294,N_10236);
nor U10529 (N_10529,N_10262,N_10309);
or U10530 (N_10530,N_10206,N_10263);
or U10531 (N_10531,N_10274,N_10268);
nor U10532 (N_10532,N_10397,N_10291);
nand U10533 (N_10533,N_10269,N_10232);
nand U10534 (N_10534,N_10365,N_10284);
or U10535 (N_10535,N_10383,N_10251);
and U10536 (N_10536,N_10262,N_10392);
or U10537 (N_10537,N_10351,N_10232);
and U10538 (N_10538,N_10328,N_10268);
or U10539 (N_10539,N_10388,N_10391);
and U10540 (N_10540,N_10350,N_10295);
xnor U10541 (N_10541,N_10207,N_10324);
and U10542 (N_10542,N_10307,N_10388);
or U10543 (N_10543,N_10244,N_10321);
xor U10544 (N_10544,N_10344,N_10362);
and U10545 (N_10545,N_10396,N_10295);
and U10546 (N_10546,N_10262,N_10269);
or U10547 (N_10547,N_10297,N_10281);
or U10548 (N_10548,N_10391,N_10313);
nor U10549 (N_10549,N_10200,N_10367);
xor U10550 (N_10550,N_10223,N_10367);
and U10551 (N_10551,N_10285,N_10228);
nor U10552 (N_10552,N_10284,N_10305);
and U10553 (N_10553,N_10341,N_10291);
nand U10554 (N_10554,N_10261,N_10213);
and U10555 (N_10555,N_10346,N_10383);
nor U10556 (N_10556,N_10287,N_10282);
or U10557 (N_10557,N_10357,N_10310);
and U10558 (N_10558,N_10356,N_10289);
xnor U10559 (N_10559,N_10230,N_10258);
or U10560 (N_10560,N_10242,N_10299);
or U10561 (N_10561,N_10391,N_10375);
nor U10562 (N_10562,N_10394,N_10288);
or U10563 (N_10563,N_10368,N_10286);
or U10564 (N_10564,N_10259,N_10314);
nor U10565 (N_10565,N_10323,N_10260);
nand U10566 (N_10566,N_10321,N_10357);
nor U10567 (N_10567,N_10315,N_10285);
or U10568 (N_10568,N_10279,N_10336);
and U10569 (N_10569,N_10229,N_10399);
nand U10570 (N_10570,N_10274,N_10371);
nor U10571 (N_10571,N_10244,N_10366);
or U10572 (N_10572,N_10252,N_10277);
and U10573 (N_10573,N_10331,N_10338);
xor U10574 (N_10574,N_10368,N_10271);
nor U10575 (N_10575,N_10301,N_10344);
nand U10576 (N_10576,N_10301,N_10378);
nand U10577 (N_10577,N_10242,N_10370);
and U10578 (N_10578,N_10394,N_10254);
nor U10579 (N_10579,N_10334,N_10221);
nand U10580 (N_10580,N_10319,N_10399);
nand U10581 (N_10581,N_10270,N_10388);
xor U10582 (N_10582,N_10290,N_10237);
nand U10583 (N_10583,N_10292,N_10301);
nand U10584 (N_10584,N_10345,N_10210);
and U10585 (N_10585,N_10362,N_10254);
nor U10586 (N_10586,N_10398,N_10255);
and U10587 (N_10587,N_10200,N_10321);
nand U10588 (N_10588,N_10398,N_10223);
nor U10589 (N_10589,N_10341,N_10252);
or U10590 (N_10590,N_10388,N_10232);
xor U10591 (N_10591,N_10219,N_10276);
nand U10592 (N_10592,N_10360,N_10261);
and U10593 (N_10593,N_10246,N_10328);
nor U10594 (N_10594,N_10258,N_10382);
or U10595 (N_10595,N_10376,N_10259);
and U10596 (N_10596,N_10308,N_10206);
or U10597 (N_10597,N_10244,N_10281);
xor U10598 (N_10598,N_10353,N_10232);
or U10599 (N_10599,N_10369,N_10376);
nand U10600 (N_10600,N_10522,N_10415);
and U10601 (N_10601,N_10488,N_10597);
or U10602 (N_10602,N_10479,N_10412);
or U10603 (N_10603,N_10506,N_10583);
xor U10604 (N_10604,N_10407,N_10552);
nor U10605 (N_10605,N_10465,N_10564);
xor U10606 (N_10606,N_10416,N_10551);
xor U10607 (N_10607,N_10433,N_10524);
nor U10608 (N_10608,N_10484,N_10428);
nor U10609 (N_10609,N_10430,N_10408);
nor U10610 (N_10610,N_10444,N_10409);
xnor U10611 (N_10611,N_10449,N_10451);
and U10612 (N_10612,N_10491,N_10487);
or U10613 (N_10613,N_10505,N_10553);
nor U10614 (N_10614,N_10545,N_10585);
nand U10615 (N_10615,N_10565,N_10536);
nand U10616 (N_10616,N_10533,N_10581);
and U10617 (N_10617,N_10466,N_10475);
or U10618 (N_10618,N_10427,N_10578);
xnor U10619 (N_10619,N_10418,N_10434);
or U10620 (N_10620,N_10580,N_10582);
nor U10621 (N_10621,N_10405,N_10579);
xor U10622 (N_10622,N_10435,N_10489);
or U10623 (N_10623,N_10439,N_10547);
nand U10624 (N_10624,N_10598,N_10570);
nor U10625 (N_10625,N_10515,N_10520);
nand U10626 (N_10626,N_10414,N_10561);
and U10627 (N_10627,N_10503,N_10425);
nor U10628 (N_10628,N_10442,N_10459);
or U10629 (N_10629,N_10542,N_10483);
nand U10630 (N_10630,N_10508,N_10539);
nor U10631 (N_10631,N_10555,N_10420);
or U10632 (N_10632,N_10504,N_10422);
or U10633 (N_10633,N_10431,N_10461);
nor U10634 (N_10634,N_10535,N_10467);
nand U10635 (N_10635,N_10492,N_10440);
or U10636 (N_10636,N_10519,N_10485);
xor U10637 (N_10637,N_10472,N_10493);
and U10638 (N_10638,N_10443,N_10562);
or U10639 (N_10639,N_10588,N_10474);
nand U10640 (N_10640,N_10595,N_10497);
xor U10641 (N_10641,N_10432,N_10557);
xor U10642 (N_10642,N_10586,N_10452);
and U10643 (N_10643,N_10401,N_10404);
xnor U10644 (N_10644,N_10511,N_10546);
nor U10645 (N_10645,N_10478,N_10512);
nand U10646 (N_10646,N_10453,N_10464);
nand U10647 (N_10647,N_10406,N_10584);
or U10648 (N_10648,N_10460,N_10436);
xor U10649 (N_10649,N_10556,N_10498);
xor U10650 (N_10650,N_10476,N_10523);
xnor U10651 (N_10651,N_10458,N_10501);
or U10652 (N_10652,N_10576,N_10477);
nor U10653 (N_10653,N_10530,N_10468);
and U10654 (N_10654,N_10531,N_10575);
nand U10655 (N_10655,N_10470,N_10499);
and U10656 (N_10656,N_10446,N_10509);
xor U10657 (N_10657,N_10495,N_10599);
xor U10658 (N_10658,N_10541,N_10481);
xnor U10659 (N_10659,N_10456,N_10590);
or U10660 (N_10660,N_10423,N_10527);
and U10661 (N_10661,N_10571,N_10486);
xnor U10662 (N_10662,N_10592,N_10514);
nand U10663 (N_10663,N_10573,N_10560);
nand U10664 (N_10664,N_10574,N_10502);
and U10665 (N_10665,N_10594,N_10426);
nand U10666 (N_10666,N_10596,N_10550);
nand U10667 (N_10667,N_10455,N_10532);
nor U10668 (N_10668,N_10589,N_10462);
nor U10669 (N_10669,N_10463,N_10513);
or U10670 (N_10670,N_10510,N_10438);
and U10671 (N_10671,N_10450,N_10419);
and U10672 (N_10672,N_10447,N_10525);
xor U10673 (N_10673,N_10469,N_10402);
nand U10674 (N_10674,N_10448,N_10548);
nand U10675 (N_10675,N_10569,N_10558);
xnor U10676 (N_10676,N_10566,N_10457);
nor U10677 (N_10677,N_10410,N_10494);
nor U10678 (N_10678,N_10526,N_10441);
or U10679 (N_10679,N_10413,N_10538);
and U10680 (N_10680,N_10437,N_10537);
nand U10681 (N_10681,N_10500,N_10549);
nor U10682 (N_10682,N_10593,N_10517);
nand U10683 (N_10683,N_10482,N_10403);
nor U10684 (N_10684,N_10516,N_10587);
xnor U10685 (N_10685,N_10572,N_10567);
nand U10686 (N_10686,N_10490,N_10454);
nand U10687 (N_10687,N_10471,N_10473);
xnor U10688 (N_10688,N_10421,N_10429);
or U10689 (N_10689,N_10554,N_10540);
nor U10690 (N_10690,N_10445,N_10507);
or U10691 (N_10691,N_10544,N_10563);
nor U10692 (N_10692,N_10400,N_10496);
nand U10693 (N_10693,N_10424,N_10577);
xor U10694 (N_10694,N_10411,N_10518);
or U10695 (N_10695,N_10543,N_10559);
xnor U10696 (N_10696,N_10534,N_10591);
xnor U10697 (N_10697,N_10417,N_10521);
nand U10698 (N_10698,N_10529,N_10480);
xnor U10699 (N_10699,N_10568,N_10528);
nor U10700 (N_10700,N_10420,N_10492);
or U10701 (N_10701,N_10471,N_10457);
nand U10702 (N_10702,N_10401,N_10483);
nor U10703 (N_10703,N_10475,N_10411);
nand U10704 (N_10704,N_10477,N_10587);
xor U10705 (N_10705,N_10514,N_10407);
or U10706 (N_10706,N_10544,N_10582);
nor U10707 (N_10707,N_10510,N_10458);
xor U10708 (N_10708,N_10509,N_10422);
nand U10709 (N_10709,N_10498,N_10403);
or U10710 (N_10710,N_10510,N_10533);
nand U10711 (N_10711,N_10589,N_10537);
xnor U10712 (N_10712,N_10540,N_10506);
and U10713 (N_10713,N_10417,N_10562);
xor U10714 (N_10714,N_10457,N_10523);
and U10715 (N_10715,N_10426,N_10412);
xnor U10716 (N_10716,N_10421,N_10406);
and U10717 (N_10717,N_10492,N_10570);
and U10718 (N_10718,N_10486,N_10587);
and U10719 (N_10719,N_10572,N_10540);
or U10720 (N_10720,N_10426,N_10547);
nor U10721 (N_10721,N_10590,N_10415);
and U10722 (N_10722,N_10597,N_10450);
nor U10723 (N_10723,N_10531,N_10434);
or U10724 (N_10724,N_10494,N_10559);
nand U10725 (N_10725,N_10479,N_10540);
and U10726 (N_10726,N_10418,N_10414);
xor U10727 (N_10727,N_10420,N_10499);
xor U10728 (N_10728,N_10483,N_10415);
nor U10729 (N_10729,N_10427,N_10489);
or U10730 (N_10730,N_10488,N_10416);
nor U10731 (N_10731,N_10559,N_10496);
nand U10732 (N_10732,N_10441,N_10426);
and U10733 (N_10733,N_10568,N_10593);
nand U10734 (N_10734,N_10404,N_10495);
and U10735 (N_10735,N_10444,N_10565);
nor U10736 (N_10736,N_10485,N_10427);
xnor U10737 (N_10737,N_10541,N_10574);
nand U10738 (N_10738,N_10574,N_10519);
nor U10739 (N_10739,N_10510,N_10482);
or U10740 (N_10740,N_10497,N_10494);
xor U10741 (N_10741,N_10443,N_10522);
or U10742 (N_10742,N_10590,N_10541);
or U10743 (N_10743,N_10538,N_10490);
or U10744 (N_10744,N_10579,N_10476);
and U10745 (N_10745,N_10539,N_10456);
nor U10746 (N_10746,N_10560,N_10418);
nand U10747 (N_10747,N_10505,N_10537);
or U10748 (N_10748,N_10453,N_10443);
nor U10749 (N_10749,N_10418,N_10466);
xnor U10750 (N_10750,N_10524,N_10585);
xnor U10751 (N_10751,N_10503,N_10445);
nand U10752 (N_10752,N_10502,N_10403);
or U10753 (N_10753,N_10518,N_10462);
or U10754 (N_10754,N_10581,N_10560);
and U10755 (N_10755,N_10481,N_10528);
and U10756 (N_10756,N_10481,N_10413);
xor U10757 (N_10757,N_10427,N_10460);
nand U10758 (N_10758,N_10523,N_10531);
nor U10759 (N_10759,N_10449,N_10563);
and U10760 (N_10760,N_10415,N_10420);
nor U10761 (N_10761,N_10508,N_10518);
and U10762 (N_10762,N_10517,N_10467);
or U10763 (N_10763,N_10596,N_10459);
xor U10764 (N_10764,N_10418,N_10544);
and U10765 (N_10765,N_10522,N_10499);
nand U10766 (N_10766,N_10461,N_10588);
nand U10767 (N_10767,N_10428,N_10576);
or U10768 (N_10768,N_10575,N_10592);
and U10769 (N_10769,N_10506,N_10501);
xnor U10770 (N_10770,N_10444,N_10426);
or U10771 (N_10771,N_10570,N_10450);
and U10772 (N_10772,N_10507,N_10509);
and U10773 (N_10773,N_10584,N_10576);
and U10774 (N_10774,N_10475,N_10599);
xor U10775 (N_10775,N_10407,N_10494);
and U10776 (N_10776,N_10532,N_10482);
nor U10777 (N_10777,N_10499,N_10416);
or U10778 (N_10778,N_10578,N_10583);
xor U10779 (N_10779,N_10494,N_10550);
nand U10780 (N_10780,N_10538,N_10454);
xnor U10781 (N_10781,N_10474,N_10561);
nand U10782 (N_10782,N_10558,N_10535);
or U10783 (N_10783,N_10463,N_10595);
nand U10784 (N_10784,N_10524,N_10419);
nand U10785 (N_10785,N_10517,N_10546);
or U10786 (N_10786,N_10557,N_10591);
nor U10787 (N_10787,N_10427,N_10501);
nor U10788 (N_10788,N_10472,N_10547);
nor U10789 (N_10789,N_10438,N_10439);
nand U10790 (N_10790,N_10483,N_10597);
nor U10791 (N_10791,N_10497,N_10433);
and U10792 (N_10792,N_10507,N_10532);
nor U10793 (N_10793,N_10449,N_10458);
nand U10794 (N_10794,N_10516,N_10422);
or U10795 (N_10795,N_10540,N_10442);
xnor U10796 (N_10796,N_10578,N_10576);
nor U10797 (N_10797,N_10464,N_10491);
and U10798 (N_10798,N_10553,N_10522);
nand U10799 (N_10799,N_10501,N_10560);
and U10800 (N_10800,N_10652,N_10795);
xor U10801 (N_10801,N_10655,N_10695);
xor U10802 (N_10802,N_10794,N_10797);
and U10803 (N_10803,N_10714,N_10705);
nor U10804 (N_10804,N_10673,N_10757);
xnor U10805 (N_10805,N_10611,N_10639);
nor U10806 (N_10806,N_10798,N_10656);
or U10807 (N_10807,N_10783,N_10684);
nor U10808 (N_10808,N_10632,N_10614);
xor U10809 (N_10809,N_10734,N_10644);
or U10810 (N_10810,N_10762,N_10676);
nand U10811 (N_10811,N_10666,N_10775);
nor U10812 (N_10812,N_10670,N_10698);
and U10813 (N_10813,N_10788,N_10736);
xor U10814 (N_10814,N_10659,N_10615);
and U10815 (N_10815,N_10715,N_10761);
or U10816 (N_10816,N_10612,N_10607);
nor U10817 (N_10817,N_10694,N_10763);
or U10818 (N_10818,N_10702,N_10687);
xor U10819 (N_10819,N_10648,N_10746);
and U10820 (N_10820,N_10600,N_10786);
xnor U10821 (N_10821,N_10679,N_10704);
and U10822 (N_10822,N_10789,N_10641);
nand U10823 (N_10823,N_10647,N_10770);
xor U10824 (N_10824,N_10646,N_10608);
nand U10825 (N_10825,N_10706,N_10766);
nand U10826 (N_10826,N_10785,N_10660);
xnor U10827 (N_10827,N_10773,N_10633);
and U10828 (N_10828,N_10737,N_10604);
xor U10829 (N_10829,N_10752,N_10740);
nor U10830 (N_10830,N_10793,N_10719);
xnor U10831 (N_10831,N_10732,N_10758);
nand U10832 (N_10832,N_10617,N_10663);
nor U10833 (N_10833,N_10693,N_10686);
and U10834 (N_10834,N_10651,N_10631);
and U10835 (N_10835,N_10602,N_10721);
nor U10836 (N_10836,N_10662,N_10699);
or U10837 (N_10837,N_10603,N_10689);
or U10838 (N_10838,N_10674,N_10735);
and U10839 (N_10839,N_10791,N_10707);
xor U10840 (N_10840,N_10754,N_10624);
or U10841 (N_10841,N_10671,N_10759);
nor U10842 (N_10842,N_10653,N_10755);
xnor U10843 (N_10843,N_10657,N_10729);
and U10844 (N_10844,N_10627,N_10700);
nor U10845 (N_10845,N_10621,N_10756);
or U10846 (N_10846,N_10629,N_10726);
nor U10847 (N_10847,N_10716,N_10744);
xnor U10848 (N_10848,N_10749,N_10605);
nor U10849 (N_10849,N_10696,N_10668);
or U10850 (N_10850,N_10690,N_10799);
and U10851 (N_10851,N_10709,N_10664);
nor U10852 (N_10852,N_10654,N_10796);
xnor U10853 (N_10853,N_10681,N_10661);
nand U10854 (N_10854,N_10748,N_10622);
nand U10855 (N_10855,N_10634,N_10645);
xnor U10856 (N_10856,N_10723,N_10730);
nand U10857 (N_10857,N_10677,N_10711);
and U10858 (N_10858,N_10768,N_10692);
xnor U10859 (N_10859,N_10739,N_10609);
nand U10860 (N_10860,N_10792,N_10787);
xor U10861 (N_10861,N_10720,N_10742);
and U10862 (N_10862,N_10642,N_10623);
or U10863 (N_10863,N_10697,N_10767);
xnor U10864 (N_10864,N_10727,N_10669);
or U10865 (N_10865,N_10665,N_10683);
or U10866 (N_10866,N_10765,N_10640);
or U10867 (N_10867,N_10731,N_10643);
or U10868 (N_10868,N_10710,N_10712);
xor U10869 (N_10869,N_10658,N_10784);
nand U10870 (N_10870,N_10636,N_10717);
nor U10871 (N_10871,N_10672,N_10619);
and U10872 (N_10872,N_10625,N_10667);
and U10873 (N_10873,N_10713,N_10628);
nand U10874 (N_10874,N_10774,N_10637);
nand U10875 (N_10875,N_10777,N_10747);
nand U10876 (N_10876,N_10620,N_10685);
or U10877 (N_10877,N_10701,N_10728);
nand U10878 (N_10878,N_10764,N_10678);
and U10879 (N_10879,N_10741,N_10616);
nor U10880 (N_10880,N_10776,N_10691);
or U10881 (N_10881,N_10610,N_10778);
and U10882 (N_10882,N_10772,N_10618);
xor U10883 (N_10883,N_10743,N_10724);
nor U10884 (N_10884,N_10649,N_10606);
or U10885 (N_10885,N_10638,N_10760);
xnor U10886 (N_10886,N_10626,N_10769);
or U10887 (N_10887,N_10722,N_10680);
nand U10888 (N_10888,N_10708,N_10753);
and U10889 (N_10889,N_10630,N_10688);
and U10890 (N_10890,N_10725,N_10790);
nor U10891 (N_10891,N_10751,N_10675);
nor U10892 (N_10892,N_10771,N_10781);
xnor U10893 (N_10893,N_10745,N_10738);
xnor U10894 (N_10894,N_10779,N_10733);
nor U10895 (N_10895,N_10601,N_10613);
or U10896 (N_10896,N_10750,N_10650);
nor U10897 (N_10897,N_10718,N_10682);
nor U10898 (N_10898,N_10703,N_10780);
or U10899 (N_10899,N_10782,N_10635);
nor U10900 (N_10900,N_10778,N_10731);
nor U10901 (N_10901,N_10786,N_10723);
or U10902 (N_10902,N_10732,N_10635);
nand U10903 (N_10903,N_10743,N_10770);
xnor U10904 (N_10904,N_10728,N_10706);
or U10905 (N_10905,N_10674,N_10658);
and U10906 (N_10906,N_10641,N_10731);
and U10907 (N_10907,N_10631,N_10618);
nand U10908 (N_10908,N_10688,N_10784);
nand U10909 (N_10909,N_10694,N_10705);
nor U10910 (N_10910,N_10704,N_10698);
and U10911 (N_10911,N_10669,N_10628);
and U10912 (N_10912,N_10643,N_10631);
or U10913 (N_10913,N_10748,N_10769);
nand U10914 (N_10914,N_10713,N_10663);
and U10915 (N_10915,N_10607,N_10646);
nand U10916 (N_10916,N_10714,N_10758);
and U10917 (N_10917,N_10782,N_10760);
xor U10918 (N_10918,N_10605,N_10614);
nor U10919 (N_10919,N_10751,N_10760);
nand U10920 (N_10920,N_10682,N_10631);
or U10921 (N_10921,N_10737,N_10721);
or U10922 (N_10922,N_10725,N_10697);
xor U10923 (N_10923,N_10733,N_10766);
or U10924 (N_10924,N_10640,N_10600);
nand U10925 (N_10925,N_10663,N_10762);
xnor U10926 (N_10926,N_10611,N_10601);
or U10927 (N_10927,N_10699,N_10638);
nor U10928 (N_10928,N_10644,N_10661);
nand U10929 (N_10929,N_10772,N_10607);
or U10930 (N_10930,N_10664,N_10744);
nand U10931 (N_10931,N_10605,N_10782);
or U10932 (N_10932,N_10775,N_10644);
xor U10933 (N_10933,N_10691,N_10727);
and U10934 (N_10934,N_10711,N_10700);
xor U10935 (N_10935,N_10721,N_10736);
nor U10936 (N_10936,N_10680,N_10770);
and U10937 (N_10937,N_10604,N_10658);
nand U10938 (N_10938,N_10763,N_10766);
nand U10939 (N_10939,N_10759,N_10795);
nand U10940 (N_10940,N_10778,N_10656);
or U10941 (N_10941,N_10774,N_10751);
or U10942 (N_10942,N_10614,N_10740);
and U10943 (N_10943,N_10665,N_10751);
or U10944 (N_10944,N_10658,N_10688);
or U10945 (N_10945,N_10799,N_10600);
and U10946 (N_10946,N_10727,N_10763);
and U10947 (N_10947,N_10647,N_10786);
nand U10948 (N_10948,N_10628,N_10721);
nor U10949 (N_10949,N_10625,N_10661);
or U10950 (N_10950,N_10620,N_10611);
nor U10951 (N_10951,N_10784,N_10601);
xnor U10952 (N_10952,N_10751,N_10715);
nand U10953 (N_10953,N_10684,N_10629);
xor U10954 (N_10954,N_10611,N_10706);
xnor U10955 (N_10955,N_10643,N_10682);
nor U10956 (N_10956,N_10753,N_10770);
xor U10957 (N_10957,N_10725,N_10696);
xnor U10958 (N_10958,N_10663,N_10725);
xor U10959 (N_10959,N_10685,N_10712);
xnor U10960 (N_10960,N_10772,N_10606);
nand U10961 (N_10961,N_10770,N_10659);
and U10962 (N_10962,N_10652,N_10616);
xor U10963 (N_10963,N_10711,N_10640);
and U10964 (N_10964,N_10658,N_10777);
nand U10965 (N_10965,N_10771,N_10718);
xnor U10966 (N_10966,N_10696,N_10799);
and U10967 (N_10967,N_10754,N_10764);
and U10968 (N_10968,N_10728,N_10694);
nand U10969 (N_10969,N_10644,N_10762);
xor U10970 (N_10970,N_10705,N_10667);
nand U10971 (N_10971,N_10766,N_10658);
nand U10972 (N_10972,N_10761,N_10757);
and U10973 (N_10973,N_10722,N_10660);
nand U10974 (N_10974,N_10672,N_10789);
nor U10975 (N_10975,N_10674,N_10799);
xnor U10976 (N_10976,N_10692,N_10684);
nor U10977 (N_10977,N_10617,N_10619);
nor U10978 (N_10978,N_10605,N_10756);
or U10979 (N_10979,N_10679,N_10744);
nand U10980 (N_10980,N_10672,N_10604);
nand U10981 (N_10981,N_10741,N_10617);
nand U10982 (N_10982,N_10750,N_10745);
and U10983 (N_10983,N_10671,N_10617);
xor U10984 (N_10984,N_10702,N_10783);
and U10985 (N_10985,N_10709,N_10632);
nand U10986 (N_10986,N_10767,N_10616);
and U10987 (N_10987,N_10738,N_10656);
nor U10988 (N_10988,N_10617,N_10677);
and U10989 (N_10989,N_10611,N_10665);
xor U10990 (N_10990,N_10732,N_10771);
or U10991 (N_10991,N_10791,N_10789);
xor U10992 (N_10992,N_10607,N_10687);
nand U10993 (N_10993,N_10664,N_10656);
and U10994 (N_10994,N_10640,N_10634);
xor U10995 (N_10995,N_10630,N_10757);
and U10996 (N_10996,N_10776,N_10674);
nor U10997 (N_10997,N_10749,N_10660);
nand U10998 (N_10998,N_10658,N_10689);
nor U10999 (N_10999,N_10786,N_10748);
xor U11000 (N_11000,N_10896,N_10908);
nand U11001 (N_11001,N_10860,N_10808);
nor U11002 (N_11002,N_10809,N_10961);
nand U11003 (N_11003,N_10870,N_10943);
nor U11004 (N_11004,N_10812,N_10970);
xnor U11005 (N_11005,N_10933,N_10982);
xnor U11006 (N_11006,N_10810,N_10911);
xor U11007 (N_11007,N_10851,N_10892);
nand U11008 (N_11008,N_10996,N_10955);
or U11009 (N_11009,N_10873,N_10947);
xor U11010 (N_11010,N_10887,N_10975);
nand U11011 (N_11011,N_10838,N_10979);
xnor U11012 (N_11012,N_10994,N_10874);
and U11013 (N_11013,N_10925,N_10803);
nor U11014 (N_11014,N_10937,N_10928);
nor U11015 (N_11015,N_10916,N_10846);
nand U11016 (N_11016,N_10964,N_10879);
or U11017 (N_11017,N_10912,N_10847);
xnor U11018 (N_11018,N_10944,N_10826);
xor U11019 (N_11019,N_10800,N_10835);
or U11020 (N_11020,N_10841,N_10929);
xor U11021 (N_11021,N_10959,N_10967);
nor U11022 (N_11022,N_10830,N_10872);
and U11023 (N_11023,N_10981,N_10844);
nor U11024 (N_11024,N_10932,N_10913);
nand U11025 (N_11025,N_10958,N_10877);
xnor U11026 (N_11026,N_10968,N_10865);
xor U11027 (N_11027,N_10997,N_10920);
or U11028 (N_11028,N_10998,N_10934);
or U11029 (N_11029,N_10811,N_10890);
or U11030 (N_11030,N_10884,N_10923);
or U11031 (N_11031,N_10829,N_10856);
nand U11032 (N_11032,N_10918,N_10946);
nor U11033 (N_11033,N_10899,N_10802);
xor U11034 (N_11034,N_10985,N_10906);
nor U11035 (N_11035,N_10969,N_10858);
or U11036 (N_11036,N_10840,N_10903);
or U11037 (N_11037,N_10861,N_10930);
and U11038 (N_11038,N_10882,N_10945);
or U11039 (N_11039,N_10924,N_10842);
and U11040 (N_11040,N_10907,N_10845);
xor U11041 (N_11041,N_10986,N_10902);
and U11042 (N_11042,N_10950,N_10813);
or U11043 (N_11043,N_10876,N_10926);
and U11044 (N_11044,N_10833,N_10956);
or U11045 (N_11045,N_10854,N_10839);
nand U11046 (N_11046,N_10965,N_10817);
and U11047 (N_11047,N_10921,N_10991);
nor U11048 (N_11048,N_10867,N_10836);
and U11049 (N_11049,N_10960,N_10825);
nor U11050 (N_11050,N_10935,N_10855);
xor U11051 (N_11051,N_10992,N_10818);
nor U11052 (N_11052,N_10828,N_10862);
nor U11053 (N_11053,N_10821,N_10922);
or U11054 (N_11054,N_10848,N_10939);
nor U11055 (N_11055,N_10832,N_10931);
and U11056 (N_11056,N_10966,N_10962);
nor U11057 (N_11057,N_10852,N_10941);
xor U11058 (N_11058,N_10927,N_10919);
and U11059 (N_11059,N_10990,N_10837);
xnor U11060 (N_11060,N_10973,N_10987);
and U11061 (N_11061,N_10963,N_10976);
nand U11062 (N_11062,N_10831,N_10875);
nand U11063 (N_11063,N_10823,N_10901);
xor U11064 (N_11064,N_10843,N_10910);
nor U11065 (N_11065,N_10864,N_10834);
xor U11066 (N_11066,N_10816,N_10989);
nor U11067 (N_11067,N_10999,N_10894);
nor U11068 (N_11068,N_10983,N_10978);
or U11069 (N_11069,N_10801,N_10914);
nand U11070 (N_11070,N_10988,N_10980);
nand U11071 (N_11071,N_10878,N_10805);
nor U11072 (N_11072,N_10885,N_10971);
or U11073 (N_11073,N_10820,N_10897);
xor U11074 (N_11074,N_10917,N_10806);
xnor U11075 (N_11075,N_10900,N_10868);
nand U11076 (N_11076,N_10880,N_10889);
nor U11077 (N_11077,N_10822,N_10957);
nand U11078 (N_11078,N_10948,N_10871);
nor U11079 (N_11079,N_10905,N_10850);
and U11080 (N_11080,N_10993,N_10883);
or U11081 (N_11081,N_10891,N_10974);
or U11082 (N_11082,N_10824,N_10881);
xnor U11083 (N_11083,N_10815,N_10951);
and U11084 (N_11084,N_10807,N_10866);
and U11085 (N_11085,N_10853,N_10904);
and U11086 (N_11086,N_10952,N_10804);
nand U11087 (N_11087,N_10995,N_10940);
nor U11088 (N_11088,N_10972,N_10893);
nor U11089 (N_11089,N_10886,N_10814);
nand U11090 (N_11090,N_10915,N_10857);
nand U11091 (N_11091,N_10869,N_10819);
nor U11092 (N_11092,N_10977,N_10938);
and U11093 (N_11093,N_10863,N_10849);
and U11094 (N_11094,N_10984,N_10936);
or U11095 (N_11095,N_10859,N_10895);
nor U11096 (N_11096,N_10898,N_10942);
nor U11097 (N_11097,N_10827,N_10909);
or U11098 (N_11098,N_10949,N_10954);
nand U11099 (N_11099,N_10888,N_10953);
nor U11100 (N_11100,N_10800,N_10997);
xnor U11101 (N_11101,N_10835,N_10943);
and U11102 (N_11102,N_10991,N_10886);
nand U11103 (N_11103,N_10964,N_10897);
and U11104 (N_11104,N_10804,N_10975);
and U11105 (N_11105,N_10909,N_10832);
or U11106 (N_11106,N_10813,N_10986);
and U11107 (N_11107,N_10845,N_10843);
nand U11108 (N_11108,N_10943,N_10840);
nand U11109 (N_11109,N_10948,N_10887);
nor U11110 (N_11110,N_10999,N_10860);
or U11111 (N_11111,N_10808,N_10897);
xnor U11112 (N_11112,N_10934,N_10812);
and U11113 (N_11113,N_10933,N_10844);
and U11114 (N_11114,N_10982,N_10914);
nand U11115 (N_11115,N_10823,N_10940);
and U11116 (N_11116,N_10935,N_10991);
xnor U11117 (N_11117,N_10917,N_10947);
nand U11118 (N_11118,N_10969,N_10896);
nand U11119 (N_11119,N_10993,N_10898);
and U11120 (N_11120,N_10947,N_10828);
xnor U11121 (N_11121,N_10927,N_10813);
and U11122 (N_11122,N_10975,N_10984);
xnor U11123 (N_11123,N_10963,N_10857);
xnor U11124 (N_11124,N_10891,N_10852);
xor U11125 (N_11125,N_10861,N_10821);
and U11126 (N_11126,N_10965,N_10945);
nand U11127 (N_11127,N_10806,N_10997);
or U11128 (N_11128,N_10926,N_10928);
and U11129 (N_11129,N_10848,N_10885);
nand U11130 (N_11130,N_10925,N_10846);
nor U11131 (N_11131,N_10879,N_10858);
nand U11132 (N_11132,N_10816,N_10902);
or U11133 (N_11133,N_10866,N_10990);
xor U11134 (N_11134,N_10843,N_10915);
and U11135 (N_11135,N_10858,N_10890);
and U11136 (N_11136,N_10918,N_10865);
nand U11137 (N_11137,N_10818,N_10887);
and U11138 (N_11138,N_10951,N_10999);
or U11139 (N_11139,N_10891,N_10992);
xor U11140 (N_11140,N_10951,N_10816);
nand U11141 (N_11141,N_10941,N_10897);
xnor U11142 (N_11142,N_10894,N_10988);
or U11143 (N_11143,N_10855,N_10933);
nand U11144 (N_11144,N_10971,N_10991);
xor U11145 (N_11145,N_10964,N_10874);
and U11146 (N_11146,N_10996,N_10957);
nor U11147 (N_11147,N_10842,N_10966);
xnor U11148 (N_11148,N_10869,N_10925);
or U11149 (N_11149,N_10914,N_10903);
nor U11150 (N_11150,N_10945,N_10821);
or U11151 (N_11151,N_10922,N_10996);
or U11152 (N_11152,N_10846,N_10804);
or U11153 (N_11153,N_10833,N_10995);
xor U11154 (N_11154,N_10882,N_10865);
or U11155 (N_11155,N_10952,N_10880);
or U11156 (N_11156,N_10893,N_10945);
and U11157 (N_11157,N_10925,N_10809);
nor U11158 (N_11158,N_10858,N_10876);
nor U11159 (N_11159,N_10831,N_10942);
nor U11160 (N_11160,N_10861,N_10954);
or U11161 (N_11161,N_10802,N_10876);
nor U11162 (N_11162,N_10816,N_10858);
and U11163 (N_11163,N_10817,N_10963);
xnor U11164 (N_11164,N_10801,N_10939);
or U11165 (N_11165,N_10881,N_10952);
xnor U11166 (N_11166,N_10953,N_10900);
xor U11167 (N_11167,N_10813,N_10867);
nor U11168 (N_11168,N_10808,N_10963);
nand U11169 (N_11169,N_10989,N_10863);
xnor U11170 (N_11170,N_10994,N_10951);
nand U11171 (N_11171,N_10867,N_10846);
and U11172 (N_11172,N_10976,N_10980);
xnor U11173 (N_11173,N_10890,N_10885);
nand U11174 (N_11174,N_10849,N_10985);
nand U11175 (N_11175,N_10994,N_10964);
and U11176 (N_11176,N_10973,N_10816);
xor U11177 (N_11177,N_10941,N_10942);
nand U11178 (N_11178,N_10910,N_10942);
xnor U11179 (N_11179,N_10971,N_10967);
nor U11180 (N_11180,N_10806,N_10807);
nor U11181 (N_11181,N_10960,N_10933);
or U11182 (N_11182,N_10915,N_10887);
xnor U11183 (N_11183,N_10995,N_10848);
and U11184 (N_11184,N_10937,N_10864);
nor U11185 (N_11185,N_10995,N_10858);
or U11186 (N_11186,N_10938,N_10873);
nor U11187 (N_11187,N_10878,N_10980);
or U11188 (N_11188,N_10960,N_10838);
xor U11189 (N_11189,N_10953,N_10913);
xnor U11190 (N_11190,N_10928,N_10840);
nor U11191 (N_11191,N_10955,N_10929);
and U11192 (N_11192,N_10851,N_10895);
nor U11193 (N_11193,N_10960,N_10957);
nor U11194 (N_11194,N_10883,N_10900);
or U11195 (N_11195,N_10964,N_10871);
nand U11196 (N_11196,N_10971,N_10866);
xnor U11197 (N_11197,N_10975,N_10946);
or U11198 (N_11198,N_10824,N_10836);
and U11199 (N_11199,N_10907,N_10996);
nand U11200 (N_11200,N_11013,N_11077);
nand U11201 (N_11201,N_11005,N_11044);
nand U11202 (N_11202,N_11041,N_11063);
or U11203 (N_11203,N_11034,N_11178);
nor U11204 (N_11204,N_11169,N_11152);
or U11205 (N_11205,N_11084,N_11174);
nand U11206 (N_11206,N_11004,N_11031);
xnor U11207 (N_11207,N_11131,N_11050);
xor U11208 (N_11208,N_11097,N_11166);
nor U11209 (N_11209,N_11007,N_11072);
nand U11210 (N_11210,N_11130,N_11183);
or U11211 (N_11211,N_11060,N_11001);
nor U11212 (N_11212,N_11135,N_11008);
nor U11213 (N_11213,N_11116,N_11117);
nor U11214 (N_11214,N_11104,N_11101);
or U11215 (N_11215,N_11188,N_11002);
xor U11216 (N_11216,N_11168,N_11124);
or U11217 (N_11217,N_11125,N_11153);
nand U11218 (N_11218,N_11122,N_11054);
nand U11219 (N_11219,N_11038,N_11182);
nor U11220 (N_11220,N_11134,N_11139);
nor U11221 (N_11221,N_11155,N_11069);
nor U11222 (N_11222,N_11156,N_11190);
or U11223 (N_11223,N_11137,N_11067);
nand U11224 (N_11224,N_11017,N_11193);
or U11225 (N_11225,N_11076,N_11073);
nand U11226 (N_11226,N_11048,N_11138);
and U11227 (N_11227,N_11146,N_11033);
or U11228 (N_11228,N_11098,N_11100);
and U11229 (N_11229,N_11071,N_11059);
xor U11230 (N_11230,N_11023,N_11057);
or U11231 (N_11231,N_11037,N_11012);
and U11232 (N_11232,N_11114,N_11172);
xor U11233 (N_11233,N_11070,N_11159);
and U11234 (N_11234,N_11011,N_11016);
or U11235 (N_11235,N_11180,N_11092);
or U11236 (N_11236,N_11160,N_11085);
xor U11237 (N_11237,N_11019,N_11158);
xor U11238 (N_11238,N_11091,N_11068);
xnor U11239 (N_11239,N_11024,N_11093);
or U11240 (N_11240,N_11043,N_11052);
nand U11241 (N_11241,N_11195,N_11095);
or U11242 (N_11242,N_11119,N_11000);
or U11243 (N_11243,N_11140,N_11022);
xnor U11244 (N_11244,N_11086,N_11055);
nand U11245 (N_11245,N_11027,N_11157);
xnor U11246 (N_11246,N_11147,N_11025);
xor U11247 (N_11247,N_11197,N_11187);
or U11248 (N_11248,N_11003,N_11039);
nand U11249 (N_11249,N_11075,N_11026);
or U11250 (N_11250,N_11148,N_11082);
xor U11251 (N_11251,N_11032,N_11189);
or U11252 (N_11252,N_11066,N_11170);
xnor U11253 (N_11253,N_11128,N_11106);
nand U11254 (N_11254,N_11030,N_11141);
or U11255 (N_11255,N_11181,N_11192);
and U11256 (N_11256,N_11145,N_11133);
or U11257 (N_11257,N_11103,N_11121);
nor U11258 (N_11258,N_11020,N_11087);
xor U11259 (N_11259,N_11080,N_11171);
xnor U11260 (N_11260,N_11015,N_11053);
nor U11261 (N_11261,N_11061,N_11079);
and U11262 (N_11262,N_11163,N_11173);
or U11263 (N_11263,N_11149,N_11143);
xnor U11264 (N_11264,N_11040,N_11162);
and U11265 (N_11265,N_11136,N_11047);
xnor U11266 (N_11266,N_11109,N_11110);
nor U11267 (N_11267,N_11045,N_11089);
nand U11268 (N_11268,N_11028,N_11126);
or U11269 (N_11269,N_11132,N_11167);
nor U11270 (N_11270,N_11185,N_11018);
nor U11271 (N_11271,N_11049,N_11165);
nor U11272 (N_11272,N_11111,N_11083);
xor U11273 (N_11273,N_11029,N_11081);
nor U11274 (N_11274,N_11035,N_11058);
xnor U11275 (N_11275,N_11056,N_11113);
or U11276 (N_11276,N_11199,N_11065);
or U11277 (N_11277,N_11078,N_11064);
nor U11278 (N_11278,N_11151,N_11176);
nand U11279 (N_11279,N_11115,N_11129);
nand U11280 (N_11280,N_11051,N_11107);
or U11281 (N_11281,N_11074,N_11123);
or U11282 (N_11282,N_11042,N_11036);
nor U11283 (N_11283,N_11105,N_11194);
nand U11284 (N_11284,N_11021,N_11161);
nand U11285 (N_11285,N_11088,N_11099);
or U11286 (N_11286,N_11009,N_11198);
or U11287 (N_11287,N_11186,N_11127);
nor U11288 (N_11288,N_11118,N_11094);
nor U11289 (N_11289,N_11006,N_11154);
or U11290 (N_11290,N_11112,N_11177);
nand U11291 (N_11291,N_11062,N_11164);
or U11292 (N_11292,N_11179,N_11108);
nand U11293 (N_11293,N_11196,N_11142);
xnor U11294 (N_11294,N_11191,N_11184);
and U11295 (N_11295,N_11096,N_11150);
xor U11296 (N_11296,N_11175,N_11102);
nor U11297 (N_11297,N_11014,N_11144);
or U11298 (N_11298,N_11090,N_11046);
nor U11299 (N_11299,N_11010,N_11120);
or U11300 (N_11300,N_11017,N_11121);
and U11301 (N_11301,N_11185,N_11160);
or U11302 (N_11302,N_11107,N_11021);
xnor U11303 (N_11303,N_11124,N_11108);
and U11304 (N_11304,N_11062,N_11137);
and U11305 (N_11305,N_11058,N_11157);
and U11306 (N_11306,N_11148,N_11158);
xor U11307 (N_11307,N_11101,N_11003);
xor U11308 (N_11308,N_11070,N_11022);
and U11309 (N_11309,N_11054,N_11080);
nor U11310 (N_11310,N_11061,N_11053);
and U11311 (N_11311,N_11100,N_11042);
and U11312 (N_11312,N_11050,N_11121);
nand U11313 (N_11313,N_11192,N_11141);
nand U11314 (N_11314,N_11162,N_11148);
or U11315 (N_11315,N_11060,N_11040);
and U11316 (N_11316,N_11118,N_11172);
nand U11317 (N_11317,N_11130,N_11126);
nand U11318 (N_11318,N_11069,N_11197);
and U11319 (N_11319,N_11170,N_11132);
nor U11320 (N_11320,N_11005,N_11104);
nand U11321 (N_11321,N_11009,N_11185);
nor U11322 (N_11322,N_11122,N_11031);
nand U11323 (N_11323,N_11110,N_11059);
and U11324 (N_11324,N_11108,N_11019);
and U11325 (N_11325,N_11054,N_11043);
or U11326 (N_11326,N_11092,N_11134);
nor U11327 (N_11327,N_11103,N_11041);
and U11328 (N_11328,N_11012,N_11035);
nor U11329 (N_11329,N_11100,N_11082);
and U11330 (N_11330,N_11075,N_11165);
xor U11331 (N_11331,N_11132,N_11165);
nor U11332 (N_11332,N_11119,N_11111);
nand U11333 (N_11333,N_11102,N_11049);
or U11334 (N_11334,N_11143,N_11160);
or U11335 (N_11335,N_11095,N_11071);
or U11336 (N_11336,N_11065,N_11162);
or U11337 (N_11337,N_11020,N_11064);
nand U11338 (N_11338,N_11011,N_11072);
or U11339 (N_11339,N_11005,N_11190);
or U11340 (N_11340,N_11065,N_11117);
or U11341 (N_11341,N_11029,N_11026);
and U11342 (N_11342,N_11063,N_11106);
xnor U11343 (N_11343,N_11150,N_11060);
and U11344 (N_11344,N_11089,N_11083);
and U11345 (N_11345,N_11127,N_11021);
or U11346 (N_11346,N_11119,N_11101);
and U11347 (N_11347,N_11169,N_11147);
nor U11348 (N_11348,N_11089,N_11086);
nand U11349 (N_11349,N_11106,N_11062);
nand U11350 (N_11350,N_11034,N_11101);
and U11351 (N_11351,N_11085,N_11190);
xor U11352 (N_11352,N_11049,N_11017);
nor U11353 (N_11353,N_11171,N_11161);
nand U11354 (N_11354,N_11063,N_11077);
xor U11355 (N_11355,N_11055,N_11129);
or U11356 (N_11356,N_11186,N_11117);
xor U11357 (N_11357,N_11032,N_11168);
nor U11358 (N_11358,N_11093,N_11156);
nand U11359 (N_11359,N_11067,N_11194);
nand U11360 (N_11360,N_11076,N_11004);
and U11361 (N_11361,N_11054,N_11033);
nand U11362 (N_11362,N_11054,N_11023);
nand U11363 (N_11363,N_11077,N_11140);
nand U11364 (N_11364,N_11136,N_11096);
nor U11365 (N_11365,N_11139,N_11050);
nand U11366 (N_11366,N_11173,N_11090);
and U11367 (N_11367,N_11164,N_11018);
xor U11368 (N_11368,N_11152,N_11023);
xnor U11369 (N_11369,N_11112,N_11196);
xor U11370 (N_11370,N_11022,N_11007);
or U11371 (N_11371,N_11151,N_11029);
nor U11372 (N_11372,N_11055,N_11143);
and U11373 (N_11373,N_11062,N_11084);
or U11374 (N_11374,N_11091,N_11113);
xor U11375 (N_11375,N_11097,N_11081);
nand U11376 (N_11376,N_11013,N_11113);
nor U11377 (N_11377,N_11125,N_11115);
and U11378 (N_11378,N_11181,N_11103);
nor U11379 (N_11379,N_11076,N_11119);
nor U11380 (N_11380,N_11175,N_11149);
nor U11381 (N_11381,N_11185,N_11015);
nor U11382 (N_11382,N_11020,N_11074);
and U11383 (N_11383,N_11127,N_11105);
or U11384 (N_11384,N_11047,N_11041);
or U11385 (N_11385,N_11074,N_11007);
nand U11386 (N_11386,N_11180,N_11100);
and U11387 (N_11387,N_11092,N_11032);
nor U11388 (N_11388,N_11034,N_11121);
xor U11389 (N_11389,N_11060,N_11002);
nand U11390 (N_11390,N_11131,N_11024);
or U11391 (N_11391,N_11129,N_11157);
or U11392 (N_11392,N_11044,N_11056);
or U11393 (N_11393,N_11089,N_11043);
nor U11394 (N_11394,N_11091,N_11002);
and U11395 (N_11395,N_11076,N_11160);
or U11396 (N_11396,N_11126,N_11006);
and U11397 (N_11397,N_11074,N_11066);
and U11398 (N_11398,N_11079,N_11015);
and U11399 (N_11399,N_11160,N_11186);
nor U11400 (N_11400,N_11399,N_11308);
nand U11401 (N_11401,N_11281,N_11317);
nand U11402 (N_11402,N_11213,N_11359);
or U11403 (N_11403,N_11348,N_11276);
and U11404 (N_11404,N_11202,N_11298);
xor U11405 (N_11405,N_11309,N_11294);
nand U11406 (N_11406,N_11268,N_11284);
xor U11407 (N_11407,N_11349,N_11303);
or U11408 (N_11408,N_11285,N_11218);
nand U11409 (N_11409,N_11283,N_11367);
xor U11410 (N_11410,N_11203,N_11265);
xnor U11411 (N_11411,N_11327,N_11331);
nand U11412 (N_11412,N_11352,N_11251);
and U11413 (N_11413,N_11393,N_11205);
nor U11414 (N_11414,N_11235,N_11320);
nand U11415 (N_11415,N_11237,N_11244);
or U11416 (N_11416,N_11270,N_11330);
and U11417 (N_11417,N_11259,N_11217);
nand U11418 (N_11418,N_11373,N_11200);
xor U11419 (N_11419,N_11390,N_11333);
nor U11420 (N_11420,N_11275,N_11232);
and U11421 (N_11421,N_11324,N_11292);
nand U11422 (N_11422,N_11382,N_11347);
or U11423 (N_11423,N_11274,N_11304);
nand U11424 (N_11424,N_11338,N_11351);
and U11425 (N_11425,N_11344,N_11346);
and U11426 (N_11426,N_11295,N_11266);
nand U11427 (N_11427,N_11236,N_11239);
and U11428 (N_11428,N_11245,N_11378);
nand U11429 (N_11429,N_11358,N_11247);
and U11430 (N_11430,N_11354,N_11287);
nor U11431 (N_11431,N_11350,N_11326);
or U11432 (N_11432,N_11353,N_11246);
nand U11433 (N_11433,N_11211,N_11214);
nor U11434 (N_11434,N_11343,N_11278);
and U11435 (N_11435,N_11241,N_11248);
xor U11436 (N_11436,N_11238,N_11206);
nand U11437 (N_11437,N_11249,N_11291);
nand U11438 (N_11438,N_11225,N_11250);
or U11439 (N_11439,N_11254,N_11384);
or U11440 (N_11440,N_11222,N_11311);
and U11441 (N_11441,N_11356,N_11305);
and U11442 (N_11442,N_11307,N_11253);
xor U11443 (N_11443,N_11328,N_11362);
or U11444 (N_11444,N_11374,N_11323);
or U11445 (N_11445,N_11372,N_11306);
and U11446 (N_11446,N_11369,N_11234);
or U11447 (N_11447,N_11355,N_11260);
xor U11448 (N_11448,N_11263,N_11375);
xnor U11449 (N_11449,N_11243,N_11256);
and U11450 (N_11450,N_11314,N_11345);
or U11451 (N_11451,N_11386,N_11231);
or U11452 (N_11452,N_11230,N_11376);
nor U11453 (N_11453,N_11233,N_11242);
nor U11454 (N_11454,N_11336,N_11267);
nor U11455 (N_11455,N_11312,N_11370);
xor U11456 (N_11456,N_11209,N_11318);
nor U11457 (N_11457,N_11365,N_11357);
nand U11458 (N_11458,N_11315,N_11223);
nor U11459 (N_11459,N_11216,N_11368);
nor U11460 (N_11460,N_11334,N_11394);
xnor U11461 (N_11461,N_11271,N_11221);
and U11462 (N_11462,N_11322,N_11341);
nand U11463 (N_11463,N_11293,N_11364);
or U11464 (N_11464,N_11340,N_11360);
nor U11465 (N_11465,N_11302,N_11337);
or U11466 (N_11466,N_11299,N_11383);
or U11467 (N_11467,N_11389,N_11286);
xor U11468 (N_11468,N_11325,N_11224);
nand U11469 (N_11469,N_11379,N_11319);
or U11470 (N_11470,N_11339,N_11329);
nor U11471 (N_11471,N_11332,N_11220);
or U11472 (N_11472,N_11363,N_11228);
xnor U11473 (N_11473,N_11366,N_11255);
and U11474 (N_11474,N_11371,N_11289);
nor U11475 (N_11475,N_11396,N_11321);
and U11476 (N_11476,N_11226,N_11279);
and U11477 (N_11477,N_11258,N_11277);
nand U11478 (N_11478,N_11300,N_11316);
nand U11479 (N_11479,N_11342,N_11229);
xor U11480 (N_11480,N_11210,N_11273);
xor U11481 (N_11481,N_11392,N_11257);
nand U11482 (N_11482,N_11201,N_11313);
nor U11483 (N_11483,N_11272,N_11215);
or U11484 (N_11484,N_11377,N_11385);
nand U11485 (N_11485,N_11208,N_11288);
nor U11486 (N_11486,N_11301,N_11204);
and U11487 (N_11487,N_11240,N_11212);
nand U11488 (N_11488,N_11395,N_11387);
xor U11489 (N_11489,N_11380,N_11391);
xnor U11490 (N_11490,N_11269,N_11261);
xnor U11491 (N_11491,N_11219,N_11297);
or U11492 (N_11492,N_11335,N_11227);
nand U11493 (N_11493,N_11262,N_11388);
xor U11494 (N_11494,N_11252,N_11207);
xnor U11495 (N_11495,N_11280,N_11290);
nor U11496 (N_11496,N_11310,N_11264);
and U11497 (N_11497,N_11361,N_11398);
xor U11498 (N_11498,N_11296,N_11397);
nand U11499 (N_11499,N_11282,N_11381);
xnor U11500 (N_11500,N_11235,N_11257);
and U11501 (N_11501,N_11315,N_11399);
nand U11502 (N_11502,N_11203,N_11275);
and U11503 (N_11503,N_11359,N_11399);
and U11504 (N_11504,N_11367,N_11320);
and U11505 (N_11505,N_11263,N_11384);
xnor U11506 (N_11506,N_11226,N_11264);
or U11507 (N_11507,N_11258,N_11371);
xor U11508 (N_11508,N_11207,N_11262);
xnor U11509 (N_11509,N_11370,N_11336);
nor U11510 (N_11510,N_11381,N_11203);
and U11511 (N_11511,N_11305,N_11256);
nand U11512 (N_11512,N_11373,N_11366);
nor U11513 (N_11513,N_11219,N_11356);
xnor U11514 (N_11514,N_11203,N_11260);
xor U11515 (N_11515,N_11283,N_11391);
xor U11516 (N_11516,N_11351,N_11243);
nor U11517 (N_11517,N_11233,N_11258);
xor U11518 (N_11518,N_11258,N_11244);
or U11519 (N_11519,N_11212,N_11251);
nor U11520 (N_11520,N_11275,N_11295);
nor U11521 (N_11521,N_11360,N_11229);
nor U11522 (N_11522,N_11235,N_11364);
and U11523 (N_11523,N_11384,N_11322);
xnor U11524 (N_11524,N_11323,N_11224);
and U11525 (N_11525,N_11302,N_11276);
nor U11526 (N_11526,N_11325,N_11351);
nand U11527 (N_11527,N_11277,N_11378);
xor U11528 (N_11528,N_11313,N_11356);
nor U11529 (N_11529,N_11220,N_11202);
or U11530 (N_11530,N_11372,N_11219);
nand U11531 (N_11531,N_11371,N_11370);
and U11532 (N_11532,N_11398,N_11237);
xnor U11533 (N_11533,N_11245,N_11356);
nor U11534 (N_11534,N_11232,N_11336);
nand U11535 (N_11535,N_11371,N_11360);
nand U11536 (N_11536,N_11256,N_11320);
nor U11537 (N_11537,N_11209,N_11242);
xor U11538 (N_11538,N_11396,N_11375);
xnor U11539 (N_11539,N_11309,N_11233);
or U11540 (N_11540,N_11297,N_11366);
nor U11541 (N_11541,N_11231,N_11395);
or U11542 (N_11542,N_11381,N_11356);
nand U11543 (N_11543,N_11284,N_11233);
xor U11544 (N_11544,N_11274,N_11265);
nor U11545 (N_11545,N_11229,N_11292);
and U11546 (N_11546,N_11282,N_11396);
and U11547 (N_11547,N_11378,N_11257);
nor U11548 (N_11548,N_11237,N_11277);
or U11549 (N_11549,N_11350,N_11266);
nor U11550 (N_11550,N_11355,N_11380);
and U11551 (N_11551,N_11247,N_11339);
nand U11552 (N_11552,N_11223,N_11347);
or U11553 (N_11553,N_11329,N_11240);
xor U11554 (N_11554,N_11248,N_11221);
nand U11555 (N_11555,N_11230,N_11373);
nand U11556 (N_11556,N_11207,N_11261);
and U11557 (N_11557,N_11389,N_11298);
or U11558 (N_11558,N_11223,N_11282);
or U11559 (N_11559,N_11340,N_11229);
nand U11560 (N_11560,N_11269,N_11380);
nand U11561 (N_11561,N_11222,N_11246);
xor U11562 (N_11562,N_11336,N_11274);
and U11563 (N_11563,N_11234,N_11278);
or U11564 (N_11564,N_11392,N_11239);
nand U11565 (N_11565,N_11285,N_11262);
nand U11566 (N_11566,N_11242,N_11218);
xor U11567 (N_11567,N_11280,N_11225);
xnor U11568 (N_11568,N_11208,N_11378);
and U11569 (N_11569,N_11372,N_11246);
and U11570 (N_11570,N_11389,N_11270);
xnor U11571 (N_11571,N_11307,N_11261);
and U11572 (N_11572,N_11351,N_11398);
nor U11573 (N_11573,N_11287,N_11386);
nor U11574 (N_11574,N_11231,N_11299);
xnor U11575 (N_11575,N_11387,N_11285);
nand U11576 (N_11576,N_11335,N_11270);
nor U11577 (N_11577,N_11374,N_11218);
nor U11578 (N_11578,N_11242,N_11267);
nor U11579 (N_11579,N_11202,N_11263);
or U11580 (N_11580,N_11232,N_11297);
nand U11581 (N_11581,N_11284,N_11256);
nor U11582 (N_11582,N_11294,N_11329);
or U11583 (N_11583,N_11219,N_11374);
or U11584 (N_11584,N_11294,N_11272);
nand U11585 (N_11585,N_11245,N_11233);
nand U11586 (N_11586,N_11372,N_11352);
xor U11587 (N_11587,N_11355,N_11381);
nand U11588 (N_11588,N_11322,N_11378);
nand U11589 (N_11589,N_11254,N_11390);
nor U11590 (N_11590,N_11261,N_11363);
xor U11591 (N_11591,N_11222,N_11336);
nand U11592 (N_11592,N_11273,N_11322);
xnor U11593 (N_11593,N_11204,N_11307);
nand U11594 (N_11594,N_11319,N_11310);
nor U11595 (N_11595,N_11314,N_11204);
xnor U11596 (N_11596,N_11289,N_11347);
nand U11597 (N_11597,N_11362,N_11266);
xnor U11598 (N_11598,N_11257,N_11329);
nor U11599 (N_11599,N_11364,N_11367);
xnor U11600 (N_11600,N_11548,N_11456);
or U11601 (N_11601,N_11416,N_11406);
or U11602 (N_11602,N_11586,N_11594);
and U11603 (N_11603,N_11486,N_11582);
and U11604 (N_11604,N_11419,N_11570);
xnor U11605 (N_11605,N_11501,N_11423);
or U11606 (N_11606,N_11543,N_11408);
nor U11607 (N_11607,N_11430,N_11588);
nand U11608 (N_11608,N_11529,N_11526);
nand U11609 (N_11609,N_11410,N_11415);
nor U11610 (N_11610,N_11592,N_11412);
nand U11611 (N_11611,N_11540,N_11461);
nand U11612 (N_11612,N_11434,N_11433);
nand U11613 (N_11613,N_11523,N_11496);
nand U11614 (N_11614,N_11598,N_11489);
xor U11615 (N_11615,N_11530,N_11542);
or U11616 (N_11616,N_11466,N_11517);
and U11617 (N_11617,N_11591,N_11509);
xor U11618 (N_11618,N_11477,N_11485);
nand U11619 (N_11619,N_11567,N_11450);
or U11620 (N_11620,N_11413,N_11460);
nand U11621 (N_11621,N_11505,N_11455);
and U11622 (N_11622,N_11537,N_11403);
or U11623 (N_11623,N_11472,N_11584);
xor U11624 (N_11624,N_11476,N_11404);
or U11625 (N_11625,N_11470,N_11506);
and U11626 (N_11626,N_11568,N_11418);
xor U11627 (N_11627,N_11411,N_11562);
xor U11628 (N_11628,N_11578,N_11405);
and U11629 (N_11629,N_11561,N_11475);
xnor U11630 (N_11630,N_11432,N_11481);
and U11631 (N_11631,N_11576,N_11593);
nor U11632 (N_11632,N_11532,N_11555);
nor U11633 (N_11633,N_11452,N_11417);
nand U11634 (N_11634,N_11577,N_11585);
nand U11635 (N_11635,N_11428,N_11484);
nor U11636 (N_11636,N_11550,N_11563);
and U11637 (N_11637,N_11522,N_11448);
or U11638 (N_11638,N_11508,N_11512);
and U11639 (N_11639,N_11597,N_11422);
xor U11640 (N_11640,N_11515,N_11587);
nor U11641 (N_11641,N_11497,N_11534);
nor U11642 (N_11642,N_11491,N_11465);
nand U11643 (N_11643,N_11440,N_11554);
and U11644 (N_11644,N_11414,N_11462);
nand U11645 (N_11645,N_11431,N_11574);
nor U11646 (N_11646,N_11493,N_11590);
nor U11647 (N_11647,N_11559,N_11494);
or U11648 (N_11648,N_11488,N_11420);
and U11649 (N_11649,N_11518,N_11579);
and U11650 (N_11650,N_11513,N_11467);
nand U11651 (N_11651,N_11546,N_11459);
nor U11652 (N_11652,N_11492,N_11596);
nand U11653 (N_11653,N_11464,N_11407);
or U11654 (N_11654,N_11444,N_11478);
and U11655 (N_11655,N_11575,N_11564);
or U11656 (N_11656,N_11439,N_11566);
nor U11657 (N_11657,N_11580,N_11401);
xor U11658 (N_11658,N_11502,N_11572);
nor U11659 (N_11659,N_11453,N_11551);
xor U11660 (N_11660,N_11435,N_11507);
and U11661 (N_11661,N_11521,N_11544);
or U11662 (N_11662,N_11511,N_11442);
and U11663 (N_11663,N_11516,N_11528);
or U11664 (N_11664,N_11498,N_11451);
or U11665 (N_11665,N_11429,N_11569);
nor U11666 (N_11666,N_11531,N_11473);
xor U11667 (N_11667,N_11487,N_11463);
nor U11668 (N_11668,N_11443,N_11557);
nand U11669 (N_11669,N_11527,N_11524);
nor U11670 (N_11670,N_11457,N_11454);
nor U11671 (N_11671,N_11549,N_11482);
and U11672 (N_11672,N_11589,N_11556);
or U11673 (N_11673,N_11445,N_11533);
or U11674 (N_11674,N_11565,N_11599);
xor U11675 (N_11675,N_11545,N_11421);
nor U11676 (N_11676,N_11541,N_11427);
and U11677 (N_11677,N_11538,N_11471);
xor U11678 (N_11678,N_11446,N_11535);
nor U11679 (N_11679,N_11500,N_11525);
or U11680 (N_11680,N_11436,N_11480);
nor U11681 (N_11681,N_11595,N_11539);
nand U11682 (N_11682,N_11474,N_11583);
xnor U11683 (N_11683,N_11479,N_11402);
xnor U11684 (N_11684,N_11400,N_11425);
and U11685 (N_11685,N_11458,N_11495);
nand U11686 (N_11686,N_11553,N_11483);
or U11687 (N_11687,N_11499,N_11409);
or U11688 (N_11688,N_11504,N_11424);
or U11689 (N_11689,N_11581,N_11520);
xnor U11690 (N_11690,N_11510,N_11503);
and U11691 (N_11691,N_11438,N_11552);
nor U11692 (N_11692,N_11437,N_11573);
and U11693 (N_11693,N_11447,N_11547);
nand U11694 (N_11694,N_11514,N_11558);
or U11695 (N_11695,N_11490,N_11441);
or U11696 (N_11696,N_11571,N_11426);
nor U11697 (N_11697,N_11469,N_11449);
xnor U11698 (N_11698,N_11468,N_11560);
or U11699 (N_11699,N_11536,N_11519);
xnor U11700 (N_11700,N_11452,N_11492);
nor U11701 (N_11701,N_11403,N_11441);
or U11702 (N_11702,N_11460,N_11489);
nor U11703 (N_11703,N_11495,N_11598);
xor U11704 (N_11704,N_11437,N_11469);
or U11705 (N_11705,N_11521,N_11428);
nand U11706 (N_11706,N_11595,N_11532);
nand U11707 (N_11707,N_11571,N_11558);
and U11708 (N_11708,N_11409,N_11576);
and U11709 (N_11709,N_11578,N_11563);
or U11710 (N_11710,N_11404,N_11538);
nand U11711 (N_11711,N_11486,N_11550);
nor U11712 (N_11712,N_11460,N_11580);
or U11713 (N_11713,N_11548,N_11524);
or U11714 (N_11714,N_11465,N_11526);
nand U11715 (N_11715,N_11412,N_11457);
and U11716 (N_11716,N_11545,N_11550);
nand U11717 (N_11717,N_11494,N_11578);
or U11718 (N_11718,N_11441,N_11508);
and U11719 (N_11719,N_11598,N_11478);
xor U11720 (N_11720,N_11535,N_11528);
nand U11721 (N_11721,N_11459,N_11502);
and U11722 (N_11722,N_11446,N_11529);
or U11723 (N_11723,N_11480,N_11592);
nor U11724 (N_11724,N_11544,N_11501);
and U11725 (N_11725,N_11419,N_11503);
or U11726 (N_11726,N_11494,N_11584);
nor U11727 (N_11727,N_11562,N_11522);
nor U11728 (N_11728,N_11526,N_11454);
xnor U11729 (N_11729,N_11478,N_11532);
nand U11730 (N_11730,N_11583,N_11411);
nor U11731 (N_11731,N_11542,N_11436);
or U11732 (N_11732,N_11416,N_11414);
nand U11733 (N_11733,N_11507,N_11475);
xor U11734 (N_11734,N_11595,N_11525);
and U11735 (N_11735,N_11458,N_11425);
xnor U11736 (N_11736,N_11560,N_11405);
and U11737 (N_11737,N_11413,N_11458);
and U11738 (N_11738,N_11415,N_11539);
nor U11739 (N_11739,N_11573,N_11583);
nor U11740 (N_11740,N_11503,N_11526);
xnor U11741 (N_11741,N_11555,N_11586);
nand U11742 (N_11742,N_11499,N_11407);
or U11743 (N_11743,N_11460,N_11497);
nor U11744 (N_11744,N_11570,N_11579);
xor U11745 (N_11745,N_11581,N_11553);
nor U11746 (N_11746,N_11549,N_11535);
or U11747 (N_11747,N_11586,N_11472);
nor U11748 (N_11748,N_11532,N_11516);
or U11749 (N_11749,N_11484,N_11493);
xnor U11750 (N_11750,N_11465,N_11501);
nand U11751 (N_11751,N_11476,N_11579);
and U11752 (N_11752,N_11522,N_11518);
or U11753 (N_11753,N_11547,N_11542);
nor U11754 (N_11754,N_11432,N_11474);
nand U11755 (N_11755,N_11468,N_11558);
and U11756 (N_11756,N_11412,N_11445);
xnor U11757 (N_11757,N_11450,N_11443);
and U11758 (N_11758,N_11538,N_11484);
nand U11759 (N_11759,N_11577,N_11546);
and U11760 (N_11760,N_11475,N_11538);
and U11761 (N_11761,N_11527,N_11406);
xnor U11762 (N_11762,N_11583,N_11542);
nand U11763 (N_11763,N_11598,N_11536);
and U11764 (N_11764,N_11516,N_11445);
and U11765 (N_11765,N_11491,N_11402);
xnor U11766 (N_11766,N_11415,N_11528);
xor U11767 (N_11767,N_11508,N_11577);
or U11768 (N_11768,N_11589,N_11484);
nor U11769 (N_11769,N_11562,N_11478);
and U11770 (N_11770,N_11466,N_11587);
nand U11771 (N_11771,N_11582,N_11574);
nor U11772 (N_11772,N_11560,N_11438);
nor U11773 (N_11773,N_11580,N_11451);
or U11774 (N_11774,N_11464,N_11548);
xor U11775 (N_11775,N_11459,N_11576);
nor U11776 (N_11776,N_11432,N_11579);
nor U11777 (N_11777,N_11440,N_11514);
and U11778 (N_11778,N_11485,N_11543);
nor U11779 (N_11779,N_11484,N_11520);
or U11780 (N_11780,N_11454,N_11550);
or U11781 (N_11781,N_11524,N_11439);
xor U11782 (N_11782,N_11556,N_11533);
nor U11783 (N_11783,N_11475,N_11430);
or U11784 (N_11784,N_11545,N_11415);
and U11785 (N_11785,N_11462,N_11569);
xnor U11786 (N_11786,N_11548,N_11410);
and U11787 (N_11787,N_11427,N_11415);
xnor U11788 (N_11788,N_11577,N_11595);
or U11789 (N_11789,N_11504,N_11459);
and U11790 (N_11790,N_11535,N_11445);
or U11791 (N_11791,N_11526,N_11459);
xor U11792 (N_11792,N_11458,N_11510);
nand U11793 (N_11793,N_11420,N_11409);
nor U11794 (N_11794,N_11457,N_11476);
nand U11795 (N_11795,N_11417,N_11532);
and U11796 (N_11796,N_11495,N_11472);
nand U11797 (N_11797,N_11525,N_11564);
nand U11798 (N_11798,N_11548,N_11433);
nand U11799 (N_11799,N_11484,N_11463);
nand U11800 (N_11800,N_11669,N_11717);
nand U11801 (N_11801,N_11763,N_11658);
xor U11802 (N_11802,N_11682,N_11655);
and U11803 (N_11803,N_11633,N_11759);
and U11804 (N_11804,N_11611,N_11775);
nor U11805 (N_11805,N_11687,N_11753);
and U11806 (N_11806,N_11751,N_11784);
nor U11807 (N_11807,N_11649,N_11607);
nand U11808 (N_11808,N_11632,N_11690);
nand U11809 (N_11809,N_11680,N_11664);
xnor U11810 (N_11810,N_11740,N_11748);
nor U11811 (N_11811,N_11625,N_11760);
or U11812 (N_11812,N_11743,N_11711);
and U11813 (N_11813,N_11615,N_11641);
xor U11814 (N_11814,N_11644,N_11779);
xnor U11815 (N_11815,N_11755,N_11667);
and U11816 (N_11816,N_11624,N_11745);
nand U11817 (N_11817,N_11636,N_11684);
xor U11818 (N_11818,N_11764,N_11742);
xnor U11819 (N_11819,N_11731,N_11673);
xor U11820 (N_11820,N_11694,N_11696);
and U11821 (N_11821,N_11640,N_11612);
and U11822 (N_11822,N_11787,N_11729);
nor U11823 (N_11823,N_11702,N_11650);
nand U11824 (N_11824,N_11668,N_11710);
xnor U11825 (N_11825,N_11619,N_11785);
nor U11826 (N_11826,N_11705,N_11732);
xor U11827 (N_11827,N_11704,N_11693);
xnor U11828 (N_11828,N_11662,N_11620);
nand U11829 (N_11829,N_11602,N_11677);
nand U11830 (N_11830,N_11609,N_11689);
xnor U11831 (N_11831,N_11697,N_11638);
xnor U11832 (N_11832,N_11622,N_11700);
and U11833 (N_11833,N_11651,N_11648);
xor U11834 (N_11834,N_11772,N_11600);
or U11835 (N_11835,N_11623,N_11777);
and U11836 (N_11836,N_11618,N_11781);
or U11837 (N_11837,N_11707,N_11774);
nand U11838 (N_11838,N_11652,N_11726);
and U11839 (N_11839,N_11765,N_11631);
xnor U11840 (N_11840,N_11686,N_11685);
and U11841 (N_11841,N_11637,N_11725);
nand U11842 (N_11842,N_11790,N_11661);
and U11843 (N_11843,N_11756,N_11703);
and U11844 (N_11844,N_11776,N_11646);
xor U11845 (N_11845,N_11714,N_11752);
or U11846 (N_11846,N_11741,N_11749);
and U11847 (N_11847,N_11718,N_11750);
or U11848 (N_11848,N_11653,N_11746);
or U11849 (N_11849,N_11713,N_11616);
xnor U11850 (N_11850,N_11758,N_11681);
nand U11851 (N_11851,N_11642,N_11692);
nand U11852 (N_11852,N_11773,N_11698);
and U11853 (N_11853,N_11720,N_11724);
nand U11854 (N_11854,N_11783,N_11671);
xor U11855 (N_11855,N_11709,N_11603);
xor U11856 (N_11856,N_11782,N_11723);
xnor U11857 (N_11857,N_11792,N_11791);
or U11858 (N_11858,N_11701,N_11706);
xor U11859 (N_11859,N_11736,N_11639);
nand U11860 (N_11860,N_11617,N_11730);
nor U11861 (N_11861,N_11794,N_11762);
xnor U11862 (N_11862,N_11606,N_11647);
and U11863 (N_11863,N_11770,N_11665);
or U11864 (N_11864,N_11610,N_11739);
or U11865 (N_11865,N_11675,N_11799);
or U11866 (N_11866,N_11767,N_11728);
and U11867 (N_11867,N_11663,N_11735);
nor U11868 (N_11868,N_11712,N_11768);
nand U11869 (N_11869,N_11757,N_11786);
xor U11870 (N_11870,N_11771,N_11766);
or U11871 (N_11871,N_11659,N_11747);
and U11872 (N_11872,N_11715,N_11676);
nand U11873 (N_11873,N_11734,N_11634);
nor U11874 (N_11874,N_11716,N_11629);
nor U11875 (N_11875,N_11727,N_11635);
or U11876 (N_11876,N_11601,N_11780);
nor U11877 (N_11877,N_11795,N_11626);
nand U11878 (N_11878,N_11744,N_11793);
or U11879 (N_11879,N_11695,N_11688);
nor U11880 (N_11880,N_11654,N_11737);
nor U11881 (N_11881,N_11719,N_11670);
nor U11882 (N_11882,N_11604,N_11613);
or U11883 (N_11883,N_11778,N_11660);
or U11884 (N_11884,N_11630,N_11733);
or U11885 (N_11885,N_11678,N_11643);
nor U11886 (N_11886,N_11754,N_11657);
xor U11887 (N_11887,N_11679,N_11788);
nand U11888 (N_11888,N_11656,N_11628);
xnor U11889 (N_11889,N_11769,N_11796);
and U11890 (N_11890,N_11708,N_11627);
and U11891 (N_11891,N_11738,N_11672);
nor U11892 (N_11892,N_11798,N_11605);
and U11893 (N_11893,N_11674,N_11691);
nor U11894 (N_11894,N_11608,N_11621);
or U11895 (N_11895,N_11761,N_11699);
xnor U11896 (N_11896,N_11645,N_11722);
xor U11897 (N_11897,N_11797,N_11789);
nand U11898 (N_11898,N_11683,N_11666);
and U11899 (N_11899,N_11614,N_11721);
and U11900 (N_11900,N_11744,N_11644);
or U11901 (N_11901,N_11625,N_11776);
or U11902 (N_11902,N_11720,N_11734);
nand U11903 (N_11903,N_11753,N_11697);
nor U11904 (N_11904,N_11723,N_11668);
or U11905 (N_11905,N_11664,N_11603);
and U11906 (N_11906,N_11796,N_11785);
and U11907 (N_11907,N_11769,N_11749);
or U11908 (N_11908,N_11799,N_11784);
xnor U11909 (N_11909,N_11607,N_11625);
or U11910 (N_11910,N_11702,N_11785);
nor U11911 (N_11911,N_11772,N_11665);
xor U11912 (N_11912,N_11730,N_11600);
and U11913 (N_11913,N_11654,N_11616);
nand U11914 (N_11914,N_11617,N_11674);
nand U11915 (N_11915,N_11605,N_11744);
and U11916 (N_11916,N_11614,N_11643);
or U11917 (N_11917,N_11682,N_11649);
and U11918 (N_11918,N_11714,N_11729);
or U11919 (N_11919,N_11723,N_11705);
xor U11920 (N_11920,N_11643,N_11773);
and U11921 (N_11921,N_11633,N_11613);
and U11922 (N_11922,N_11737,N_11601);
nand U11923 (N_11923,N_11759,N_11766);
nor U11924 (N_11924,N_11759,N_11796);
nor U11925 (N_11925,N_11613,N_11625);
nor U11926 (N_11926,N_11771,N_11658);
and U11927 (N_11927,N_11600,N_11666);
and U11928 (N_11928,N_11627,N_11671);
and U11929 (N_11929,N_11623,N_11722);
nor U11930 (N_11930,N_11743,N_11796);
or U11931 (N_11931,N_11779,N_11707);
and U11932 (N_11932,N_11633,N_11672);
nor U11933 (N_11933,N_11713,N_11775);
and U11934 (N_11934,N_11738,N_11773);
xor U11935 (N_11935,N_11648,N_11708);
xor U11936 (N_11936,N_11621,N_11620);
xor U11937 (N_11937,N_11728,N_11646);
and U11938 (N_11938,N_11659,N_11729);
xor U11939 (N_11939,N_11660,N_11618);
nor U11940 (N_11940,N_11649,N_11601);
nor U11941 (N_11941,N_11664,N_11717);
xnor U11942 (N_11942,N_11776,N_11705);
nand U11943 (N_11943,N_11714,N_11663);
nor U11944 (N_11944,N_11713,N_11785);
or U11945 (N_11945,N_11755,N_11600);
nor U11946 (N_11946,N_11690,N_11648);
or U11947 (N_11947,N_11789,N_11679);
or U11948 (N_11948,N_11655,N_11706);
xnor U11949 (N_11949,N_11718,N_11639);
xnor U11950 (N_11950,N_11669,N_11693);
and U11951 (N_11951,N_11796,N_11737);
or U11952 (N_11952,N_11728,N_11750);
nand U11953 (N_11953,N_11771,N_11625);
and U11954 (N_11954,N_11649,N_11628);
xnor U11955 (N_11955,N_11765,N_11708);
xnor U11956 (N_11956,N_11740,N_11710);
and U11957 (N_11957,N_11605,N_11623);
and U11958 (N_11958,N_11600,N_11635);
and U11959 (N_11959,N_11708,N_11698);
and U11960 (N_11960,N_11673,N_11661);
or U11961 (N_11961,N_11764,N_11757);
nor U11962 (N_11962,N_11710,N_11635);
nand U11963 (N_11963,N_11707,N_11786);
xor U11964 (N_11964,N_11790,N_11798);
xor U11965 (N_11965,N_11653,N_11644);
nor U11966 (N_11966,N_11662,N_11728);
or U11967 (N_11967,N_11794,N_11706);
and U11968 (N_11968,N_11626,N_11629);
xnor U11969 (N_11969,N_11661,N_11671);
and U11970 (N_11970,N_11766,N_11608);
nand U11971 (N_11971,N_11630,N_11646);
or U11972 (N_11972,N_11750,N_11715);
xor U11973 (N_11973,N_11748,N_11716);
nor U11974 (N_11974,N_11740,N_11700);
and U11975 (N_11975,N_11799,N_11641);
nand U11976 (N_11976,N_11701,N_11728);
nor U11977 (N_11977,N_11722,N_11689);
nand U11978 (N_11978,N_11661,N_11788);
nand U11979 (N_11979,N_11721,N_11744);
or U11980 (N_11980,N_11771,N_11707);
or U11981 (N_11981,N_11722,N_11644);
and U11982 (N_11982,N_11753,N_11696);
or U11983 (N_11983,N_11792,N_11616);
nor U11984 (N_11984,N_11752,N_11680);
or U11985 (N_11985,N_11652,N_11683);
nor U11986 (N_11986,N_11746,N_11719);
or U11987 (N_11987,N_11709,N_11602);
nor U11988 (N_11988,N_11768,N_11765);
and U11989 (N_11989,N_11618,N_11736);
nor U11990 (N_11990,N_11659,N_11796);
xor U11991 (N_11991,N_11746,N_11678);
or U11992 (N_11992,N_11746,N_11705);
nor U11993 (N_11993,N_11798,N_11643);
and U11994 (N_11994,N_11714,N_11765);
and U11995 (N_11995,N_11782,N_11607);
xor U11996 (N_11996,N_11766,N_11698);
xor U11997 (N_11997,N_11645,N_11774);
xnor U11998 (N_11998,N_11761,N_11734);
nand U11999 (N_11999,N_11670,N_11678);
or U12000 (N_12000,N_11953,N_11908);
or U12001 (N_12001,N_11950,N_11892);
nand U12002 (N_12002,N_11921,N_11850);
xor U12003 (N_12003,N_11825,N_11926);
nand U12004 (N_12004,N_11972,N_11981);
nand U12005 (N_12005,N_11896,N_11983);
nand U12006 (N_12006,N_11846,N_11862);
or U12007 (N_12007,N_11873,N_11871);
or U12008 (N_12008,N_11868,N_11909);
xnor U12009 (N_12009,N_11945,N_11931);
nand U12010 (N_12010,N_11867,N_11821);
nand U12011 (N_12011,N_11823,N_11923);
or U12012 (N_12012,N_11853,N_11958);
xor U12013 (N_12013,N_11857,N_11841);
nand U12014 (N_12014,N_11939,N_11886);
nor U12015 (N_12015,N_11959,N_11837);
nor U12016 (N_12016,N_11883,N_11954);
nor U12017 (N_12017,N_11810,N_11885);
nor U12018 (N_12018,N_11806,N_11961);
and U12019 (N_12019,N_11912,N_11832);
xnor U12020 (N_12020,N_11803,N_11922);
xnor U12021 (N_12021,N_11955,N_11811);
and U12022 (N_12022,N_11845,N_11976);
and U12023 (N_12023,N_11947,N_11990);
and U12024 (N_12024,N_11944,N_11942);
nor U12025 (N_12025,N_11865,N_11970);
nor U12026 (N_12026,N_11924,N_11993);
nor U12027 (N_12027,N_11992,N_11969);
nand U12028 (N_12028,N_11989,N_11848);
nor U12029 (N_12029,N_11964,N_11965);
and U12030 (N_12030,N_11902,N_11874);
nand U12031 (N_12031,N_11987,N_11877);
nand U12032 (N_12032,N_11834,N_11984);
nand U12033 (N_12033,N_11804,N_11977);
nor U12034 (N_12034,N_11920,N_11980);
nand U12035 (N_12035,N_11893,N_11826);
nand U12036 (N_12036,N_11836,N_11847);
and U12037 (N_12037,N_11808,N_11991);
nor U12038 (N_12038,N_11956,N_11890);
and U12039 (N_12039,N_11986,N_11824);
nor U12040 (N_12040,N_11988,N_11929);
nor U12041 (N_12041,N_11996,N_11899);
or U12042 (N_12042,N_11975,N_11861);
nand U12043 (N_12043,N_11974,N_11916);
nor U12044 (N_12044,N_11919,N_11872);
nor U12045 (N_12045,N_11835,N_11895);
xnor U12046 (N_12046,N_11968,N_11875);
and U12047 (N_12047,N_11948,N_11888);
nand U12048 (N_12048,N_11928,N_11915);
nor U12049 (N_12049,N_11998,N_11805);
and U12050 (N_12050,N_11960,N_11833);
and U12051 (N_12051,N_11809,N_11820);
nand U12052 (N_12052,N_11973,N_11844);
and U12053 (N_12053,N_11876,N_11822);
and U12054 (N_12054,N_11938,N_11897);
nor U12055 (N_12055,N_11930,N_11949);
xnor U12056 (N_12056,N_11831,N_11830);
nand U12057 (N_12057,N_11863,N_11935);
nand U12058 (N_12058,N_11843,N_11901);
xor U12059 (N_12059,N_11851,N_11952);
and U12060 (N_12060,N_11828,N_11997);
nand U12061 (N_12061,N_11894,N_11891);
or U12062 (N_12062,N_11913,N_11906);
or U12063 (N_12063,N_11904,N_11827);
or U12064 (N_12064,N_11860,N_11817);
nand U12065 (N_12065,N_11936,N_11917);
or U12066 (N_12066,N_11887,N_11802);
xor U12067 (N_12067,N_11957,N_11979);
xor U12068 (N_12068,N_11814,N_11941);
and U12069 (N_12069,N_11878,N_11829);
nand U12070 (N_12070,N_11978,N_11816);
or U12071 (N_12071,N_11927,N_11925);
xnor U12072 (N_12072,N_11967,N_11943);
xor U12073 (N_12073,N_11866,N_11880);
or U12074 (N_12074,N_11994,N_11813);
or U12075 (N_12075,N_11918,N_11858);
xnor U12076 (N_12076,N_11963,N_11881);
nor U12077 (N_12077,N_11999,N_11898);
or U12078 (N_12078,N_11849,N_11995);
and U12079 (N_12079,N_11838,N_11937);
xnor U12080 (N_12080,N_11884,N_11842);
or U12081 (N_12081,N_11934,N_11801);
and U12082 (N_12082,N_11852,N_11900);
and U12083 (N_12083,N_11985,N_11932);
and U12084 (N_12084,N_11911,N_11819);
xor U12085 (N_12085,N_11951,N_11812);
nand U12086 (N_12086,N_11940,N_11870);
xnor U12087 (N_12087,N_11815,N_11982);
nor U12088 (N_12088,N_11966,N_11882);
xor U12089 (N_12089,N_11855,N_11818);
xor U12090 (N_12090,N_11859,N_11879);
nor U12091 (N_12091,N_11800,N_11807);
nor U12092 (N_12092,N_11869,N_11910);
and U12093 (N_12093,N_11933,N_11946);
xor U12094 (N_12094,N_11905,N_11839);
and U12095 (N_12095,N_11856,N_11914);
or U12096 (N_12096,N_11889,N_11962);
nand U12097 (N_12097,N_11840,N_11907);
and U12098 (N_12098,N_11971,N_11903);
xnor U12099 (N_12099,N_11864,N_11854);
or U12100 (N_12100,N_11811,N_11888);
or U12101 (N_12101,N_11821,N_11986);
nand U12102 (N_12102,N_11856,N_11837);
nor U12103 (N_12103,N_11919,N_11865);
and U12104 (N_12104,N_11899,N_11944);
xor U12105 (N_12105,N_11837,N_11961);
and U12106 (N_12106,N_11908,N_11932);
xnor U12107 (N_12107,N_11834,N_11899);
nand U12108 (N_12108,N_11821,N_11990);
and U12109 (N_12109,N_11832,N_11840);
nand U12110 (N_12110,N_11825,N_11806);
nand U12111 (N_12111,N_11938,N_11914);
and U12112 (N_12112,N_11848,N_11809);
nor U12113 (N_12113,N_11955,N_11977);
and U12114 (N_12114,N_11991,N_11970);
xnor U12115 (N_12115,N_11970,N_11937);
nand U12116 (N_12116,N_11899,N_11838);
nor U12117 (N_12117,N_11850,N_11980);
and U12118 (N_12118,N_11845,N_11915);
nor U12119 (N_12119,N_11955,N_11936);
xor U12120 (N_12120,N_11926,N_11857);
nor U12121 (N_12121,N_11958,N_11994);
and U12122 (N_12122,N_11934,N_11861);
nor U12123 (N_12123,N_11860,N_11811);
or U12124 (N_12124,N_11846,N_11896);
or U12125 (N_12125,N_11843,N_11965);
or U12126 (N_12126,N_11884,N_11915);
nor U12127 (N_12127,N_11976,N_11879);
nand U12128 (N_12128,N_11858,N_11881);
nand U12129 (N_12129,N_11816,N_11865);
or U12130 (N_12130,N_11983,N_11830);
nand U12131 (N_12131,N_11870,N_11852);
nor U12132 (N_12132,N_11885,N_11897);
nand U12133 (N_12133,N_11870,N_11990);
xnor U12134 (N_12134,N_11930,N_11857);
or U12135 (N_12135,N_11932,N_11865);
nand U12136 (N_12136,N_11828,N_11979);
xnor U12137 (N_12137,N_11918,N_11830);
nor U12138 (N_12138,N_11927,N_11816);
nand U12139 (N_12139,N_11991,N_11803);
nand U12140 (N_12140,N_11896,N_11841);
xor U12141 (N_12141,N_11896,N_11905);
nand U12142 (N_12142,N_11811,N_11838);
xnor U12143 (N_12143,N_11869,N_11959);
nand U12144 (N_12144,N_11915,N_11864);
and U12145 (N_12145,N_11809,N_11965);
nand U12146 (N_12146,N_11925,N_11959);
xnor U12147 (N_12147,N_11922,N_11992);
nand U12148 (N_12148,N_11967,N_11805);
xnor U12149 (N_12149,N_11932,N_11830);
nor U12150 (N_12150,N_11957,N_11953);
xor U12151 (N_12151,N_11819,N_11828);
or U12152 (N_12152,N_11901,N_11803);
and U12153 (N_12153,N_11958,N_11831);
xor U12154 (N_12154,N_11962,N_11911);
or U12155 (N_12155,N_11885,N_11942);
and U12156 (N_12156,N_11922,N_11876);
or U12157 (N_12157,N_11870,N_11869);
and U12158 (N_12158,N_11896,N_11853);
nor U12159 (N_12159,N_11861,N_11814);
nand U12160 (N_12160,N_11806,N_11948);
and U12161 (N_12161,N_11918,N_11912);
and U12162 (N_12162,N_11831,N_11931);
xor U12163 (N_12163,N_11927,N_11823);
nor U12164 (N_12164,N_11919,N_11819);
nor U12165 (N_12165,N_11857,N_11828);
nand U12166 (N_12166,N_11880,N_11935);
nor U12167 (N_12167,N_11916,N_11966);
and U12168 (N_12168,N_11896,N_11909);
xnor U12169 (N_12169,N_11836,N_11861);
nor U12170 (N_12170,N_11964,N_11975);
nor U12171 (N_12171,N_11955,N_11971);
nand U12172 (N_12172,N_11899,N_11858);
nand U12173 (N_12173,N_11924,N_11860);
nand U12174 (N_12174,N_11852,N_11968);
xor U12175 (N_12175,N_11997,N_11923);
nand U12176 (N_12176,N_11802,N_11973);
and U12177 (N_12177,N_11994,N_11943);
or U12178 (N_12178,N_11998,N_11862);
or U12179 (N_12179,N_11945,N_11963);
nor U12180 (N_12180,N_11940,N_11895);
nand U12181 (N_12181,N_11958,N_11916);
nor U12182 (N_12182,N_11814,N_11887);
nand U12183 (N_12183,N_11900,N_11951);
nand U12184 (N_12184,N_11844,N_11934);
or U12185 (N_12185,N_11870,N_11845);
and U12186 (N_12186,N_11974,N_11825);
nand U12187 (N_12187,N_11948,N_11939);
nand U12188 (N_12188,N_11922,N_11841);
nand U12189 (N_12189,N_11998,N_11844);
or U12190 (N_12190,N_11940,N_11802);
nor U12191 (N_12191,N_11950,N_11877);
and U12192 (N_12192,N_11824,N_11979);
or U12193 (N_12193,N_11877,N_11870);
or U12194 (N_12194,N_11887,N_11822);
and U12195 (N_12195,N_11910,N_11934);
nor U12196 (N_12196,N_11823,N_11847);
nand U12197 (N_12197,N_11957,N_11977);
or U12198 (N_12198,N_11964,N_11962);
nor U12199 (N_12199,N_11961,N_11882);
nor U12200 (N_12200,N_12008,N_12128);
nand U12201 (N_12201,N_12173,N_12024);
or U12202 (N_12202,N_12193,N_12012);
and U12203 (N_12203,N_12121,N_12070);
or U12204 (N_12204,N_12107,N_12146);
nand U12205 (N_12205,N_12112,N_12068);
nand U12206 (N_12206,N_12100,N_12035);
xor U12207 (N_12207,N_12002,N_12021);
and U12208 (N_12208,N_12114,N_12136);
or U12209 (N_12209,N_12110,N_12033);
nor U12210 (N_12210,N_12025,N_12057);
xnor U12211 (N_12211,N_12199,N_12054);
nor U12212 (N_12212,N_12122,N_12067);
and U12213 (N_12213,N_12142,N_12196);
and U12214 (N_12214,N_12034,N_12190);
and U12215 (N_12215,N_12032,N_12064);
nor U12216 (N_12216,N_12195,N_12104);
and U12217 (N_12217,N_12073,N_12105);
nor U12218 (N_12218,N_12094,N_12078);
or U12219 (N_12219,N_12076,N_12144);
nand U12220 (N_12220,N_12086,N_12171);
xnor U12221 (N_12221,N_12091,N_12179);
xor U12222 (N_12222,N_12069,N_12071);
nand U12223 (N_12223,N_12113,N_12041);
and U12224 (N_12224,N_12124,N_12188);
nand U12225 (N_12225,N_12162,N_12053);
xnor U12226 (N_12226,N_12186,N_12158);
or U12227 (N_12227,N_12184,N_12149);
nand U12228 (N_12228,N_12116,N_12049);
and U12229 (N_12229,N_12020,N_12165);
and U12230 (N_12230,N_12017,N_12000);
or U12231 (N_12231,N_12077,N_12085);
xor U12232 (N_12232,N_12151,N_12159);
nor U12233 (N_12233,N_12132,N_12138);
nand U12234 (N_12234,N_12014,N_12103);
or U12235 (N_12235,N_12191,N_12084);
xor U12236 (N_12236,N_12029,N_12163);
or U12237 (N_12237,N_12045,N_12013);
nand U12238 (N_12238,N_12123,N_12197);
or U12239 (N_12239,N_12133,N_12063);
xnor U12240 (N_12240,N_12050,N_12130);
nor U12241 (N_12241,N_12182,N_12161);
or U12242 (N_12242,N_12001,N_12023);
or U12243 (N_12243,N_12044,N_12031);
xor U12244 (N_12244,N_12090,N_12175);
and U12245 (N_12245,N_12119,N_12164);
or U12246 (N_12246,N_12028,N_12066);
xor U12247 (N_12247,N_12027,N_12139);
and U12248 (N_12248,N_12111,N_12183);
nand U12249 (N_12249,N_12172,N_12009);
nand U12250 (N_12250,N_12087,N_12106);
xnor U12251 (N_12251,N_12074,N_12192);
and U12252 (N_12252,N_12180,N_12169);
nor U12253 (N_12253,N_12048,N_12040);
and U12254 (N_12254,N_12148,N_12055);
nor U12255 (N_12255,N_12155,N_12176);
or U12256 (N_12256,N_12082,N_12152);
nand U12257 (N_12257,N_12089,N_12059);
nor U12258 (N_12258,N_12154,N_12194);
or U12259 (N_12259,N_12102,N_12178);
xnor U12260 (N_12260,N_12125,N_12185);
xor U12261 (N_12261,N_12051,N_12093);
nand U12262 (N_12262,N_12126,N_12039);
nand U12263 (N_12263,N_12150,N_12056);
nand U12264 (N_12264,N_12010,N_12062);
nor U12265 (N_12265,N_12147,N_12166);
xor U12266 (N_12266,N_12109,N_12092);
and U12267 (N_12267,N_12134,N_12037);
or U12268 (N_12268,N_12079,N_12108);
and U12269 (N_12269,N_12047,N_12038);
or U12270 (N_12270,N_12004,N_12120);
nor U12271 (N_12271,N_12088,N_12043);
and U12272 (N_12272,N_12016,N_12006);
or U12273 (N_12273,N_12030,N_12083);
and U12274 (N_12274,N_12117,N_12036);
or U12275 (N_12275,N_12167,N_12095);
and U12276 (N_12276,N_12018,N_12046);
nor U12277 (N_12277,N_12052,N_12072);
and U12278 (N_12278,N_12131,N_12075);
xnor U12279 (N_12279,N_12168,N_12098);
and U12280 (N_12280,N_12189,N_12140);
nor U12281 (N_12281,N_12181,N_12022);
xnor U12282 (N_12282,N_12061,N_12015);
nand U12283 (N_12283,N_12118,N_12160);
and U12284 (N_12284,N_12127,N_12141);
xnor U12285 (N_12285,N_12177,N_12081);
xor U12286 (N_12286,N_12153,N_12065);
xnor U12287 (N_12287,N_12099,N_12003);
xnor U12288 (N_12288,N_12157,N_12137);
nand U12289 (N_12289,N_12097,N_12096);
nand U12290 (N_12290,N_12101,N_12019);
or U12291 (N_12291,N_12005,N_12042);
nor U12292 (N_12292,N_12060,N_12170);
nand U12293 (N_12293,N_12135,N_12187);
xnor U12294 (N_12294,N_12143,N_12115);
and U12295 (N_12295,N_12145,N_12129);
xnor U12296 (N_12296,N_12011,N_12080);
nand U12297 (N_12297,N_12007,N_12174);
or U12298 (N_12298,N_12026,N_12156);
or U12299 (N_12299,N_12058,N_12198);
nor U12300 (N_12300,N_12027,N_12054);
xor U12301 (N_12301,N_12069,N_12052);
and U12302 (N_12302,N_12137,N_12099);
nor U12303 (N_12303,N_12024,N_12020);
nand U12304 (N_12304,N_12067,N_12130);
or U12305 (N_12305,N_12002,N_12036);
or U12306 (N_12306,N_12089,N_12100);
nor U12307 (N_12307,N_12081,N_12001);
nand U12308 (N_12308,N_12178,N_12117);
xnor U12309 (N_12309,N_12127,N_12040);
nor U12310 (N_12310,N_12033,N_12165);
and U12311 (N_12311,N_12037,N_12162);
xor U12312 (N_12312,N_12116,N_12006);
nand U12313 (N_12313,N_12187,N_12176);
nand U12314 (N_12314,N_12051,N_12078);
nor U12315 (N_12315,N_12019,N_12179);
or U12316 (N_12316,N_12143,N_12061);
and U12317 (N_12317,N_12158,N_12049);
and U12318 (N_12318,N_12156,N_12076);
or U12319 (N_12319,N_12067,N_12006);
or U12320 (N_12320,N_12119,N_12054);
nor U12321 (N_12321,N_12033,N_12076);
nor U12322 (N_12322,N_12126,N_12167);
nand U12323 (N_12323,N_12113,N_12180);
and U12324 (N_12324,N_12015,N_12171);
or U12325 (N_12325,N_12154,N_12067);
or U12326 (N_12326,N_12159,N_12120);
and U12327 (N_12327,N_12157,N_12134);
xor U12328 (N_12328,N_12172,N_12075);
xnor U12329 (N_12329,N_12047,N_12085);
or U12330 (N_12330,N_12178,N_12172);
and U12331 (N_12331,N_12104,N_12018);
and U12332 (N_12332,N_12167,N_12145);
and U12333 (N_12333,N_12114,N_12127);
or U12334 (N_12334,N_12001,N_12130);
or U12335 (N_12335,N_12003,N_12145);
or U12336 (N_12336,N_12189,N_12161);
and U12337 (N_12337,N_12171,N_12019);
nand U12338 (N_12338,N_12040,N_12154);
and U12339 (N_12339,N_12065,N_12096);
xor U12340 (N_12340,N_12092,N_12197);
or U12341 (N_12341,N_12195,N_12198);
and U12342 (N_12342,N_12113,N_12073);
or U12343 (N_12343,N_12054,N_12017);
nor U12344 (N_12344,N_12087,N_12124);
nor U12345 (N_12345,N_12132,N_12064);
nand U12346 (N_12346,N_12003,N_12044);
and U12347 (N_12347,N_12156,N_12080);
nor U12348 (N_12348,N_12148,N_12073);
nor U12349 (N_12349,N_12177,N_12039);
nand U12350 (N_12350,N_12015,N_12000);
nor U12351 (N_12351,N_12084,N_12135);
nand U12352 (N_12352,N_12123,N_12171);
or U12353 (N_12353,N_12173,N_12150);
and U12354 (N_12354,N_12177,N_12149);
xor U12355 (N_12355,N_12175,N_12163);
nor U12356 (N_12356,N_12143,N_12102);
xnor U12357 (N_12357,N_12010,N_12168);
xor U12358 (N_12358,N_12028,N_12111);
and U12359 (N_12359,N_12098,N_12081);
and U12360 (N_12360,N_12148,N_12120);
xor U12361 (N_12361,N_12050,N_12014);
nand U12362 (N_12362,N_12046,N_12066);
and U12363 (N_12363,N_12184,N_12039);
xor U12364 (N_12364,N_12096,N_12095);
or U12365 (N_12365,N_12076,N_12163);
xor U12366 (N_12366,N_12176,N_12034);
nor U12367 (N_12367,N_12040,N_12159);
nor U12368 (N_12368,N_12101,N_12100);
and U12369 (N_12369,N_12120,N_12023);
nand U12370 (N_12370,N_12132,N_12165);
nand U12371 (N_12371,N_12028,N_12007);
nor U12372 (N_12372,N_12071,N_12035);
or U12373 (N_12373,N_12093,N_12126);
nor U12374 (N_12374,N_12034,N_12123);
and U12375 (N_12375,N_12029,N_12009);
xor U12376 (N_12376,N_12093,N_12085);
nand U12377 (N_12377,N_12055,N_12144);
nor U12378 (N_12378,N_12168,N_12028);
and U12379 (N_12379,N_12166,N_12104);
xnor U12380 (N_12380,N_12060,N_12105);
nor U12381 (N_12381,N_12030,N_12079);
or U12382 (N_12382,N_12099,N_12064);
nand U12383 (N_12383,N_12132,N_12105);
and U12384 (N_12384,N_12178,N_12110);
nand U12385 (N_12385,N_12048,N_12123);
and U12386 (N_12386,N_12024,N_12176);
xnor U12387 (N_12387,N_12120,N_12189);
xor U12388 (N_12388,N_12188,N_12039);
nand U12389 (N_12389,N_12015,N_12149);
and U12390 (N_12390,N_12001,N_12162);
or U12391 (N_12391,N_12073,N_12075);
or U12392 (N_12392,N_12134,N_12061);
or U12393 (N_12393,N_12094,N_12036);
xnor U12394 (N_12394,N_12071,N_12150);
xnor U12395 (N_12395,N_12081,N_12040);
xnor U12396 (N_12396,N_12156,N_12085);
and U12397 (N_12397,N_12018,N_12191);
and U12398 (N_12398,N_12194,N_12083);
and U12399 (N_12399,N_12185,N_12004);
and U12400 (N_12400,N_12347,N_12204);
or U12401 (N_12401,N_12328,N_12276);
or U12402 (N_12402,N_12249,N_12238);
and U12403 (N_12403,N_12302,N_12319);
nand U12404 (N_12404,N_12248,N_12368);
nand U12405 (N_12405,N_12270,N_12338);
and U12406 (N_12406,N_12366,N_12350);
or U12407 (N_12407,N_12371,N_12246);
nand U12408 (N_12408,N_12278,N_12221);
nor U12409 (N_12409,N_12341,N_12218);
or U12410 (N_12410,N_12277,N_12339);
and U12411 (N_12411,N_12318,N_12200);
nand U12412 (N_12412,N_12256,N_12356);
xor U12413 (N_12413,N_12201,N_12247);
xor U12414 (N_12414,N_12299,N_12300);
or U12415 (N_12415,N_12229,N_12304);
nor U12416 (N_12416,N_12337,N_12205);
or U12417 (N_12417,N_12367,N_12202);
and U12418 (N_12418,N_12351,N_12352);
nand U12419 (N_12419,N_12281,N_12364);
or U12420 (N_12420,N_12309,N_12237);
nor U12421 (N_12421,N_12267,N_12254);
and U12422 (N_12422,N_12324,N_12297);
or U12423 (N_12423,N_12264,N_12245);
xor U12424 (N_12424,N_12291,N_12227);
xnor U12425 (N_12425,N_12342,N_12209);
nor U12426 (N_12426,N_12308,N_12288);
nand U12427 (N_12427,N_12388,N_12212);
nor U12428 (N_12428,N_12322,N_12327);
and U12429 (N_12429,N_12244,N_12354);
xnor U12430 (N_12430,N_12259,N_12386);
xor U12431 (N_12431,N_12359,N_12358);
and U12432 (N_12432,N_12286,N_12280);
nor U12433 (N_12433,N_12207,N_12384);
nand U12434 (N_12434,N_12253,N_12226);
nand U12435 (N_12435,N_12306,N_12345);
nor U12436 (N_12436,N_12239,N_12320);
nand U12437 (N_12437,N_12290,N_12349);
xnor U12438 (N_12438,N_12283,N_12310);
nor U12439 (N_12439,N_12363,N_12233);
nor U12440 (N_12440,N_12343,N_12295);
xnor U12441 (N_12441,N_12214,N_12383);
nand U12442 (N_12442,N_12390,N_12379);
or U12443 (N_12443,N_12323,N_12369);
nand U12444 (N_12444,N_12397,N_12334);
nor U12445 (N_12445,N_12287,N_12274);
nand U12446 (N_12446,N_12216,N_12213);
or U12447 (N_12447,N_12292,N_12375);
and U12448 (N_12448,N_12321,N_12241);
xnor U12449 (N_12449,N_12335,N_12385);
and U12450 (N_12450,N_12340,N_12217);
xnor U12451 (N_12451,N_12316,N_12333);
nor U12452 (N_12452,N_12398,N_12305);
nor U12453 (N_12453,N_12263,N_12353);
and U12454 (N_12454,N_12208,N_12266);
nand U12455 (N_12455,N_12243,N_12370);
or U12456 (N_12456,N_12326,N_12377);
nor U12457 (N_12457,N_12220,N_12381);
or U12458 (N_12458,N_12225,N_12240);
nand U12459 (N_12459,N_12275,N_12273);
nand U12460 (N_12460,N_12374,N_12293);
and U12461 (N_12461,N_12357,N_12389);
nor U12462 (N_12462,N_12344,N_12311);
and U12463 (N_12463,N_12250,N_12255);
xnor U12464 (N_12464,N_12392,N_12269);
nor U12465 (N_12465,N_12394,N_12234);
and U12466 (N_12466,N_12313,N_12317);
xnor U12467 (N_12467,N_12257,N_12296);
nor U12468 (N_12468,N_12399,N_12391);
or U12469 (N_12469,N_12230,N_12312);
and U12470 (N_12470,N_12382,N_12372);
and U12471 (N_12471,N_12262,N_12271);
nor U12472 (N_12472,N_12303,N_12348);
or U12473 (N_12473,N_12332,N_12223);
and U12474 (N_12474,N_12251,N_12285);
or U12475 (N_12475,N_12331,N_12294);
or U12476 (N_12476,N_12307,N_12282);
nor U12477 (N_12477,N_12376,N_12361);
and U12478 (N_12478,N_12329,N_12330);
xnor U12479 (N_12479,N_12268,N_12206);
nor U12480 (N_12480,N_12365,N_12396);
and U12481 (N_12481,N_12235,N_12346);
nor U12482 (N_12482,N_12236,N_12362);
xor U12483 (N_12483,N_12279,N_12325);
nor U12484 (N_12484,N_12315,N_12284);
or U12485 (N_12485,N_12219,N_12222);
xnor U12486 (N_12486,N_12336,N_12298);
nand U12487 (N_12487,N_12265,N_12210);
nand U12488 (N_12488,N_12387,N_12393);
nor U12489 (N_12489,N_12242,N_12355);
xnor U12490 (N_12490,N_12395,N_12301);
or U12491 (N_12491,N_12203,N_12228);
or U12492 (N_12492,N_12373,N_12272);
nor U12493 (N_12493,N_12252,N_12232);
nor U12494 (N_12494,N_12224,N_12378);
or U12495 (N_12495,N_12261,N_12360);
xnor U12496 (N_12496,N_12215,N_12289);
nand U12497 (N_12497,N_12260,N_12314);
or U12498 (N_12498,N_12380,N_12211);
nand U12499 (N_12499,N_12231,N_12258);
xor U12500 (N_12500,N_12399,N_12270);
and U12501 (N_12501,N_12225,N_12219);
or U12502 (N_12502,N_12332,N_12345);
nand U12503 (N_12503,N_12364,N_12304);
nor U12504 (N_12504,N_12280,N_12259);
or U12505 (N_12505,N_12369,N_12209);
or U12506 (N_12506,N_12349,N_12280);
nand U12507 (N_12507,N_12269,N_12375);
and U12508 (N_12508,N_12236,N_12209);
or U12509 (N_12509,N_12344,N_12325);
xnor U12510 (N_12510,N_12224,N_12295);
xor U12511 (N_12511,N_12340,N_12292);
nor U12512 (N_12512,N_12313,N_12232);
nor U12513 (N_12513,N_12239,N_12304);
xor U12514 (N_12514,N_12328,N_12348);
or U12515 (N_12515,N_12229,N_12378);
and U12516 (N_12516,N_12262,N_12336);
nor U12517 (N_12517,N_12392,N_12289);
or U12518 (N_12518,N_12215,N_12243);
xnor U12519 (N_12519,N_12221,N_12337);
nor U12520 (N_12520,N_12382,N_12346);
xnor U12521 (N_12521,N_12229,N_12265);
xnor U12522 (N_12522,N_12332,N_12356);
xnor U12523 (N_12523,N_12384,N_12281);
nand U12524 (N_12524,N_12315,N_12277);
or U12525 (N_12525,N_12397,N_12314);
xor U12526 (N_12526,N_12234,N_12262);
or U12527 (N_12527,N_12230,N_12383);
nand U12528 (N_12528,N_12348,N_12292);
nand U12529 (N_12529,N_12331,N_12369);
or U12530 (N_12530,N_12217,N_12319);
xor U12531 (N_12531,N_12220,N_12268);
and U12532 (N_12532,N_12277,N_12335);
and U12533 (N_12533,N_12306,N_12383);
and U12534 (N_12534,N_12220,N_12343);
nand U12535 (N_12535,N_12392,N_12255);
or U12536 (N_12536,N_12278,N_12366);
or U12537 (N_12537,N_12327,N_12203);
xnor U12538 (N_12538,N_12375,N_12276);
and U12539 (N_12539,N_12252,N_12355);
nand U12540 (N_12540,N_12393,N_12289);
and U12541 (N_12541,N_12268,N_12349);
nor U12542 (N_12542,N_12357,N_12216);
nand U12543 (N_12543,N_12356,N_12377);
or U12544 (N_12544,N_12273,N_12364);
or U12545 (N_12545,N_12331,N_12213);
nor U12546 (N_12546,N_12248,N_12397);
xor U12547 (N_12547,N_12391,N_12307);
xnor U12548 (N_12548,N_12211,N_12252);
or U12549 (N_12549,N_12252,N_12334);
xnor U12550 (N_12550,N_12366,N_12208);
or U12551 (N_12551,N_12216,N_12375);
nor U12552 (N_12552,N_12311,N_12317);
or U12553 (N_12553,N_12300,N_12337);
and U12554 (N_12554,N_12305,N_12220);
xnor U12555 (N_12555,N_12381,N_12306);
and U12556 (N_12556,N_12302,N_12291);
and U12557 (N_12557,N_12365,N_12252);
and U12558 (N_12558,N_12248,N_12262);
and U12559 (N_12559,N_12268,N_12299);
and U12560 (N_12560,N_12287,N_12248);
nand U12561 (N_12561,N_12224,N_12389);
or U12562 (N_12562,N_12399,N_12243);
and U12563 (N_12563,N_12368,N_12245);
or U12564 (N_12564,N_12357,N_12272);
or U12565 (N_12565,N_12398,N_12272);
and U12566 (N_12566,N_12356,N_12329);
nand U12567 (N_12567,N_12228,N_12250);
or U12568 (N_12568,N_12331,N_12279);
or U12569 (N_12569,N_12363,N_12291);
nand U12570 (N_12570,N_12213,N_12207);
and U12571 (N_12571,N_12244,N_12263);
and U12572 (N_12572,N_12219,N_12275);
nor U12573 (N_12573,N_12355,N_12396);
nor U12574 (N_12574,N_12363,N_12229);
or U12575 (N_12575,N_12295,N_12225);
nor U12576 (N_12576,N_12203,N_12394);
nand U12577 (N_12577,N_12221,N_12370);
xnor U12578 (N_12578,N_12286,N_12393);
nor U12579 (N_12579,N_12221,N_12358);
or U12580 (N_12580,N_12291,N_12287);
nor U12581 (N_12581,N_12288,N_12362);
nand U12582 (N_12582,N_12297,N_12283);
and U12583 (N_12583,N_12315,N_12291);
nor U12584 (N_12584,N_12368,N_12335);
xnor U12585 (N_12585,N_12364,N_12382);
or U12586 (N_12586,N_12322,N_12316);
and U12587 (N_12587,N_12320,N_12381);
and U12588 (N_12588,N_12279,N_12333);
nand U12589 (N_12589,N_12360,N_12286);
and U12590 (N_12590,N_12204,N_12210);
xnor U12591 (N_12591,N_12339,N_12203);
and U12592 (N_12592,N_12289,N_12394);
or U12593 (N_12593,N_12221,N_12213);
xnor U12594 (N_12594,N_12388,N_12217);
or U12595 (N_12595,N_12298,N_12221);
or U12596 (N_12596,N_12320,N_12337);
and U12597 (N_12597,N_12264,N_12261);
nor U12598 (N_12598,N_12365,N_12394);
or U12599 (N_12599,N_12368,N_12364);
and U12600 (N_12600,N_12492,N_12500);
nand U12601 (N_12601,N_12583,N_12430);
xnor U12602 (N_12602,N_12584,N_12465);
or U12603 (N_12603,N_12532,N_12576);
and U12604 (N_12604,N_12569,N_12435);
nand U12605 (N_12605,N_12514,N_12407);
and U12606 (N_12606,N_12516,N_12457);
nor U12607 (N_12607,N_12416,N_12597);
nor U12608 (N_12608,N_12505,N_12421);
nand U12609 (N_12609,N_12444,N_12535);
and U12610 (N_12610,N_12491,N_12429);
nand U12611 (N_12611,N_12408,N_12469);
xnor U12612 (N_12612,N_12404,N_12446);
xor U12613 (N_12613,N_12451,N_12463);
nand U12614 (N_12614,N_12533,N_12536);
or U12615 (N_12615,N_12562,N_12439);
or U12616 (N_12616,N_12461,N_12493);
and U12617 (N_12617,N_12587,N_12401);
or U12618 (N_12618,N_12534,N_12511);
or U12619 (N_12619,N_12415,N_12464);
and U12620 (N_12620,N_12594,N_12485);
nor U12621 (N_12621,N_12510,N_12557);
or U12622 (N_12622,N_12445,N_12427);
nand U12623 (N_12623,N_12498,N_12437);
and U12624 (N_12624,N_12580,N_12555);
nand U12625 (N_12625,N_12410,N_12522);
nor U12626 (N_12626,N_12566,N_12554);
xor U12627 (N_12627,N_12443,N_12547);
and U12628 (N_12628,N_12561,N_12552);
xor U12629 (N_12629,N_12486,N_12470);
nor U12630 (N_12630,N_12543,N_12438);
nor U12631 (N_12631,N_12546,N_12577);
or U12632 (N_12632,N_12468,N_12459);
nor U12633 (N_12633,N_12565,N_12483);
or U12634 (N_12634,N_12524,N_12455);
xor U12635 (N_12635,N_12507,N_12527);
nand U12636 (N_12636,N_12556,N_12509);
or U12637 (N_12637,N_12454,N_12409);
nor U12638 (N_12638,N_12403,N_12472);
xor U12639 (N_12639,N_12520,N_12489);
xor U12640 (N_12640,N_12585,N_12542);
and U12641 (N_12641,N_12538,N_12578);
and U12642 (N_12642,N_12448,N_12423);
nor U12643 (N_12643,N_12517,N_12406);
xor U12644 (N_12644,N_12539,N_12420);
or U12645 (N_12645,N_12418,N_12523);
or U12646 (N_12646,N_12467,N_12508);
nand U12647 (N_12647,N_12490,N_12590);
xor U12648 (N_12648,N_12519,N_12440);
nor U12649 (N_12649,N_12503,N_12488);
and U12650 (N_12650,N_12480,N_12458);
xnor U12651 (N_12651,N_12419,N_12521);
and U12652 (N_12652,N_12400,N_12506);
nand U12653 (N_12653,N_12413,N_12579);
nor U12654 (N_12654,N_12598,N_12518);
nand U12655 (N_12655,N_12482,N_12481);
xnor U12656 (N_12656,N_12499,N_12588);
nand U12657 (N_12657,N_12550,N_12572);
nand U12658 (N_12658,N_12487,N_12479);
nand U12659 (N_12659,N_12450,N_12412);
and U12660 (N_12660,N_12582,N_12586);
nand U12661 (N_12661,N_12405,N_12563);
and U12662 (N_12662,N_12417,N_12466);
nand U12663 (N_12663,N_12564,N_12537);
nor U12664 (N_12664,N_12548,N_12570);
nand U12665 (N_12665,N_12471,N_12425);
nor U12666 (N_12666,N_12558,N_12595);
and U12667 (N_12667,N_12593,N_12599);
xor U12668 (N_12668,N_12559,N_12402);
nand U12669 (N_12669,N_12477,N_12540);
nand U12670 (N_12670,N_12447,N_12453);
and U12671 (N_12671,N_12411,N_12592);
nand U12672 (N_12672,N_12449,N_12530);
nor U12673 (N_12673,N_12441,N_12544);
xnor U12674 (N_12674,N_12553,N_12526);
nand U12675 (N_12675,N_12529,N_12478);
or U12676 (N_12676,N_12575,N_12424);
and U12677 (N_12677,N_12571,N_12502);
nand U12678 (N_12678,N_12474,N_12591);
or U12679 (N_12679,N_12496,N_12560);
nand U12680 (N_12680,N_12442,N_12501);
or U12681 (N_12681,N_12568,N_12436);
xnor U12682 (N_12682,N_12432,N_12431);
nor U12683 (N_12683,N_12495,N_12574);
nor U12684 (N_12684,N_12497,N_12513);
and U12685 (N_12685,N_12573,N_12452);
and U12686 (N_12686,N_12484,N_12515);
nor U12687 (N_12687,N_12549,N_12473);
xor U12688 (N_12688,N_12525,N_12504);
xnor U12689 (N_12689,N_12428,N_12414);
xnor U12690 (N_12690,N_12422,N_12541);
xor U12691 (N_12691,N_12434,N_12476);
nor U12692 (N_12692,N_12581,N_12494);
and U12693 (N_12693,N_12460,N_12456);
and U12694 (N_12694,N_12433,N_12545);
nand U12695 (N_12695,N_12528,N_12551);
and U12696 (N_12696,N_12567,N_12531);
nor U12697 (N_12697,N_12426,N_12512);
nand U12698 (N_12698,N_12462,N_12475);
and U12699 (N_12699,N_12589,N_12596);
nand U12700 (N_12700,N_12410,N_12484);
nor U12701 (N_12701,N_12580,N_12594);
nor U12702 (N_12702,N_12599,N_12542);
or U12703 (N_12703,N_12504,N_12522);
and U12704 (N_12704,N_12534,N_12504);
nor U12705 (N_12705,N_12550,N_12573);
nor U12706 (N_12706,N_12577,N_12568);
nor U12707 (N_12707,N_12432,N_12599);
xnor U12708 (N_12708,N_12593,N_12519);
or U12709 (N_12709,N_12454,N_12443);
nand U12710 (N_12710,N_12538,N_12453);
xnor U12711 (N_12711,N_12581,N_12446);
xnor U12712 (N_12712,N_12507,N_12535);
nand U12713 (N_12713,N_12414,N_12582);
nand U12714 (N_12714,N_12532,N_12410);
and U12715 (N_12715,N_12504,N_12440);
nor U12716 (N_12716,N_12406,N_12433);
nor U12717 (N_12717,N_12526,N_12409);
nor U12718 (N_12718,N_12465,N_12543);
nand U12719 (N_12719,N_12590,N_12517);
xnor U12720 (N_12720,N_12402,N_12557);
xor U12721 (N_12721,N_12578,N_12417);
xor U12722 (N_12722,N_12590,N_12417);
xnor U12723 (N_12723,N_12471,N_12415);
or U12724 (N_12724,N_12586,N_12508);
and U12725 (N_12725,N_12435,N_12436);
and U12726 (N_12726,N_12462,N_12434);
xnor U12727 (N_12727,N_12583,N_12553);
and U12728 (N_12728,N_12584,N_12468);
nand U12729 (N_12729,N_12533,N_12489);
nor U12730 (N_12730,N_12573,N_12592);
nand U12731 (N_12731,N_12473,N_12408);
and U12732 (N_12732,N_12592,N_12401);
nor U12733 (N_12733,N_12500,N_12512);
xor U12734 (N_12734,N_12460,N_12454);
xor U12735 (N_12735,N_12571,N_12417);
and U12736 (N_12736,N_12475,N_12470);
nand U12737 (N_12737,N_12585,N_12441);
nand U12738 (N_12738,N_12465,N_12558);
and U12739 (N_12739,N_12545,N_12484);
nor U12740 (N_12740,N_12505,N_12407);
nand U12741 (N_12741,N_12586,N_12452);
nor U12742 (N_12742,N_12515,N_12440);
xor U12743 (N_12743,N_12569,N_12546);
xnor U12744 (N_12744,N_12439,N_12564);
or U12745 (N_12745,N_12453,N_12462);
xor U12746 (N_12746,N_12428,N_12579);
or U12747 (N_12747,N_12404,N_12429);
nand U12748 (N_12748,N_12500,N_12567);
or U12749 (N_12749,N_12411,N_12588);
nand U12750 (N_12750,N_12566,N_12548);
nor U12751 (N_12751,N_12470,N_12493);
or U12752 (N_12752,N_12533,N_12555);
or U12753 (N_12753,N_12419,N_12414);
nor U12754 (N_12754,N_12588,N_12558);
nand U12755 (N_12755,N_12487,N_12589);
or U12756 (N_12756,N_12559,N_12456);
nand U12757 (N_12757,N_12450,N_12501);
or U12758 (N_12758,N_12510,N_12473);
or U12759 (N_12759,N_12576,N_12539);
or U12760 (N_12760,N_12500,N_12422);
nand U12761 (N_12761,N_12445,N_12502);
or U12762 (N_12762,N_12430,N_12460);
nand U12763 (N_12763,N_12439,N_12581);
xor U12764 (N_12764,N_12475,N_12455);
or U12765 (N_12765,N_12435,N_12429);
and U12766 (N_12766,N_12424,N_12531);
and U12767 (N_12767,N_12531,N_12457);
nand U12768 (N_12768,N_12560,N_12577);
nor U12769 (N_12769,N_12501,N_12505);
or U12770 (N_12770,N_12410,N_12510);
nand U12771 (N_12771,N_12441,N_12410);
and U12772 (N_12772,N_12576,N_12515);
nand U12773 (N_12773,N_12591,N_12559);
nand U12774 (N_12774,N_12577,N_12474);
nand U12775 (N_12775,N_12454,N_12479);
xor U12776 (N_12776,N_12574,N_12518);
nand U12777 (N_12777,N_12544,N_12541);
nor U12778 (N_12778,N_12537,N_12417);
nor U12779 (N_12779,N_12468,N_12594);
or U12780 (N_12780,N_12452,N_12414);
nor U12781 (N_12781,N_12510,N_12448);
nand U12782 (N_12782,N_12522,N_12441);
and U12783 (N_12783,N_12438,N_12452);
xor U12784 (N_12784,N_12528,N_12425);
or U12785 (N_12785,N_12404,N_12497);
or U12786 (N_12786,N_12560,N_12595);
nor U12787 (N_12787,N_12570,N_12451);
or U12788 (N_12788,N_12422,N_12543);
xor U12789 (N_12789,N_12569,N_12493);
and U12790 (N_12790,N_12552,N_12432);
and U12791 (N_12791,N_12526,N_12522);
nand U12792 (N_12792,N_12401,N_12574);
nand U12793 (N_12793,N_12461,N_12582);
nor U12794 (N_12794,N_12442,N_12557);
nor U12795 (N_12795,N_12432,N_12511);
nand U12796 (N_12796,N_12539,N_12481);
nor U12797 (N_12797,N_12587,N_12512);
nor U12798 (N_12798,N_12527,N_12544);
nand U12799 (N_12799,N_12410,N_12538);
and U12800 (N_12800,N_12751,N_12610);
and U12801 (N_12801,N_12739,N_12716);
and U12802 (N_12802,N_12607,N_12679);
nor U12803 (N_12803,N_12733,N_12783);
or U12804 (N_12804,N_12726,N_12602);
nand U12805 (N_12805,N_12772,N_12795);
or U12806 (N_12806,N_12673,N_12680);
nand U12807 (N_12807,N_12682,N_12600);
or U12808 (N_12808,N_12691,N_12638);
and U12809 (N_12809,N_12753,N_12755);
nand U12810 (N_12810,N_12737,N_12654);
or U12811 (N_12811,N_12765,N_12613);
or U12812 (N_12812,N_12653,N_12674);
and U12813 (N_12813,N_12721,N_12760);
nand U12814 (N_12814,N_12616,N_12605);
nor U12815 (N_12815,N_12759,N_12723);
nand U12816 (N_12816,N_12782,N_12722);
or U12817 (N_12817,N_12685,N_12784);
nand U12818 (N_12818,N_12729,N_12746);
and U12819 (N_12819,N_12786,N_12608);
nor U12820 (N_12820,N_12693,N_12697);
and U12821 (N_12821,N_12659,N_12713);
or U12822 (N_12822,N_12668,N_12719);
or U12823 (N_12823,N_12624,N_12611);
nand U12824 (N_12824,N_12766,N_12769);
nor U12825 (N_12825,N_12735,N_12627);
nor U12826 (N_12826,N_12690,N_12656);
nand U12827 (N_12827,N_12606,N_12628);
nor U12828 (N_12828,N_12789,N_12650);
nand U12829 (N_12829,N_12618,N_12712);
nand U12830 (N_12830,N_12762,N_12764);
and U12831 (N_12831,N_12730,N_12745);
nand U12832 (N_12832,N_12662,N_12792);
nand U12833 (N_12833,N_12672,N_12647);
nor U12834 (N_12834,N_12695,N_12698);
or U12835 (N_12835,N_12774,N_12666);
xor U12836 (N_12836,N_12617,N_12796);
nor U12837 (N_12837,N_12683,N_12758);
xnor U12838 (N_12838,N_12700,N_12715);
or U12839 (N_12839,N_12655,N_12775);
and U12840 (N_12840,N_12787,N_12625);
and U12841 (N_12841,N_12641,N_12614);
or U12842 (N_12842,N_12699,N_12752);
and U12843 (N_12843,N_12703,N_12687);
or U12844 (N_12844,N_12718,N_12701);
and U12845 (N_12845,N_12645,N_12731);
xnor U12846 (N_12846,N_12757,N_12619);
and U12847 (N_12847,N_12648,N_12770);
nand U12848 (N_12848,N_12761,N_12704);
and U12849 (N_12849,N_12709,N_12660);
xor U12850 (N_12850,N_12675,N_12686);
nand U12851 (N_12851,N_12747,N_12740);
xnor U12852 (N_12852,N_12707,N_12652);
xnor U12853 (N_12853,N_12702,N_12741);
xnor U12854 (N_12854,N_12754,N_12706);
or U12855 (N_12855,N_12630,N_12724);
or U12856 (N_12856,N_12620,N_12738);
or U12857 (N_12857,N_12615,N_12657);
nand U12858 (N_12858,N_12636,N_12736);
xnor U12859 (N_12859,N_12694,N_12670);
nand U12860 (N_12860,N_12776,N_12678);
nand U12861 (N_12861,N_12637,N_12643);
and U12862 (N_12862,N_12728,N_12788);
nand U12863 (N_12863,N_12669,N_12767);
xor U12864 (N_12864,N_12734,N_12661);
xor U12865 (N_12865,N_12646,N_12640);
and U12866 (N_12866,N_12604,N_12744);
or U12867 (N_12867,N_12711,N_12609);
or U12868 (N_12868,N_12612,N_12742);
and U12869 (N_12869,N_12756,N_12785);
nand U12870 (N_12870,N_12749,N_12658);
nand U12871 (N_12871,N_12797,N_12631);
nand U12872 (N_12872,N_12748,N_12671);
nand U12873 (N_12873,N_12603,N_12720);
and U12874 (N_12874,N_12644,N_12681);
and U12875 (N_12875,N_12750,N_12705);
nand U12876 (N_12876,N_12692,N_12773);
xnor U12877 (N_12877,N_12793,N_12663);
and U12878 (N_12878,N_12725,N_12689);
nand U12879 (N_12879,N_12777,N_12635);
nor U12880 (N_12880,N_12779,N_12714);
and U12881 (N_12881,N_12629,N_12732);
nor U12882 (N_12882,N_12778,N_12622);
nand U12883 (N_12883,N_12623,N_12667);
or U12884 (N_12884,N_12649,N_12688);
or U12885 (N_12885,N_12708,N_12790);
xnor U12886 (N_12886,N_12634,N_12639);
nand U12887 (N_12887,N_12771,N_12684);
or U12888 (N_12888,N_12664,N_12696);
nor U12889 (N_12889,N_12763,N_12781);
nand U12890 (N_12890,N_12717,N_12799);
and U12891 (N_12891,N_12626,N_12727);
nor U12892 (N_12892,N_12601,N_12676);
nor U12893 (N_12893,N_12677,N_12651);
and U12894 (N_12894,N_12794,N_12743);
nand U12895 (N_12895,N_12791,N_12632);
and U12896 (N_12896,N_12665,N_12642);
nand U12897 (N_12897,N_12798,N_12710);
and U12898 (N_12898,N_12780,N_12621);
or U12899 (N_12899,N_12633,N_12768);
nor U12900 (N_12900,N_12781,N_12665);
nand U12901 (N_12901,N_12713,N_12763);
nor U12902 (N_12902,N_12699,N_12668);
or U12903 (N_12903,N_12645,N_12726);
nor U12904 (N_12904,N_12726,N_12754);
or U12905 (N_12905,N_12644,N_12607);
nor U12906 (N_12906,N_12788,N_12608);
nor U12907 (N_12907,N_12656,N_12720);
or U12908 (N_12908,N_12743,N_12739);
nand U12909 (N_12909,N_12655,N_12714);
and U12910 (N_12910,N_12740,N_12683);
or U12911 (N_12911,N_12672,N_12654);
xor U12912 (N_12912,N_12615,N_12669);
nand U12913 (N_12913,N_12774,N_12703);
nand U12914 (N_12914,N_12714,N_12664);
nor U12915 (N_12915,N_12661,N_12626);
xnor U12916 (N_12916,N_12776,N_12756);
xor U12917 (N_12917,N_12767,N_12693);
nor U12918 (N_12918,N_12792,N_12735);
nor U12919 (N_12919,N_12758,N_12737);
nand U12920 (N_12920,N_12733,N_12689);
xnor U12921 (N_12921,N_12778,N_12605);
xnor U12922 (N_12922,N_12622,N_12641);
nor U12923 (N_12923,N_12646,N_12760);
nor U12924 (N_12924,N_12618,N_12773);
xnor U12925 (N_12925,N_12723,N_12621);
nor U12926 (N_12926,N_12675,N_12711);
xor U12927 (N_12927,N_12748,N_12664);
xnor U12928 (N_12928,N_12721,N_12731);
and U12929 (N_12929,N_12773,N_12766);
or U12930 (N_12930,N_12792,N_12720);
or U12931 (N_12931,N_12744,N_12789);
and U12932 (N_12932,N_12616,N_12645);
and U12933 (N_12933,N_12791,N_12634);
nor U12934 (N_12934,N_12637,N_12611);
or U12935 (N_12935,N_12610,N_12791);
xor U12936 (N_12936,N_12726,N_12710);
and U12937 (N_12937,N_12792,N_12769);
and U12938 (N_12938,N_12705,N_12706);
nand U12939 (N_12939,N_12720,N_12722);
nor U12940 (N_12940,N_12661,N_12611);
nand U12941 (N_12941,N_12691,N_12686);
xnor U12942 (N_12942,N_12767,N_12739);
xor U12943 (N_12943,N_12630,N_12659);
xnor U12944 (N_12944,N_12659,N_12749);
nor U12945 (N_12945,N_12601,N_12700);
and U12946 (N_12946,N_12704,N_12689);
nor U12947 (N_12947,N_12650,N_12615);
nand U12948 (N_12948,N_12724,N_12645);
xnor U12949 (N_12949,N_12735,N_12785);
xnor U12950 (N_12950,N_12680,N_12645);
xor U12951 (N_12951,N_12787,N_12732);
and U12952 (N_12952,N_12712,N_12684);
nor U12953 (N_12953,N_12684,N_12734);
or U12954 (N_12954,N_12764,N_12707);
or U12955 (N_12955,N_12740,N_12787);
and U12956 (N_12956,N_12749,N_12734);
and U12957 (N_12957,N_12683,N_12714);
nand U12958 (N_12958,N_12689,N_12645);
xor U12959 (N_12959,N_12629,N_12640);
and U12960 (N_12960,N_12684,N_12644);
and U12961 (N_12961,N_12696,N_12752);
or U12962 (N_12962,N_12780,N_12741);
or U12963 (N_12963,N_12614,N_12765);
or U12964 (N_12964,N_12709,N_12607);
and U12965 (N_12965,N_12719,N_12692);
xor U12966 (N_12966,N_12736,N_12734);
and U12967 (N_12967,N_12761,N_12702);
nor U12968 (N_12968,N_12609,N_12639);
and U12969 (N_12969,N_12710,N_12763);
nand U12970 (N_12970,N_12683,N_12743);
nor U12971 (N_12971,N_12799,N_12735);
or U12972 (N_12972,N_12679,N_12701);
nand U12973 (N_12973,N_12763,N_12705);
xnor U12974 (N_12974,N_12698,N_12779);
xor U12975 (N_12975,N_12697,N_12796);
and U12976 (N_12976,N_12602,N_12720);
and U12977 (N_12977,N_12708,N_12669);
nand U12978 (N_12978,N_12792,N_12699);
xor U12979 (N_12979,N_12692,N_12622);
nor U12980 (N_12980,N_12749,N_12660);
nor U12981 (N_12981,N_12617,N_12658);
nand U12982 (N_12982,N_12628,N_12758);
xnor U12983 (N_12983,N_12661,N_12750);
nor U12984 (N_12984,N_12735,N_12753);
and U12985 (N_12985,N_12673,N_12700);
xor U12986 (N_12986,N_12641,N_12748);
nand U12987 (N_12987,N_12603,N_12791);
or U12988 (N_12988,N_12680,N_12745);
nor U12989 (N_12989,N_12614,N_12704);
xor U12990 (N_12990,N_12630,N_12763);
and U12991 (N_12991,N_12691,N_12705);
and U12992 (N_12992,N_12788,N_12777);
nand U12993 (N_12993,N_12692,N_12713);
xor U12994 (N_12994,N_12736,N_12775);
and U12995 (N_12995,N_12727,N_12729);
and U12996 (N_12996,N_12717,N_12610);
nor U12997 (N_12997,N_12758,N_12763);
nand U12998 (N_12998,N_12723,N_12643);
xnor U12999 (N_12999,N_12638,N_12607);
xnor U13000 (N_13000,N_12923,N_12914);
nor U13001 (N_13001,N_12938,N_12954);
nand U13002 (N_13002,N_12837,N_12859);
or U13003 (N_13003,N_12806,N_12835);
xnor U13004 (N_13004,N_12838,N_12944);
or U13005 (N_13005,N_12941,N_12811);
nor U13006 (N_13006,N_12945,N_12857);
and U13007 (N_13007,N_12893,N_12829);
nor U13008 (N_13008,N_12860,N_12831);
or U13009 (N_13009,N_12836,N_12872);
nand U13010 (N_13010,N_12854,N_12992);
nor U13011 (N_13011,N_12973,N_12863);
and U13012 (N_13012,N_12826,N_12972);
nor U13013 (N_13013,N_12980,N_12902);
and U13014 (N_13014,N_12959,N_12886);
xnor U13015 (N_13015,N_12927,N_12918);
and U13016 (N_13016,N_12996,N_12804);
nand U13017 (N_13017,N_12948,N_12809);
or U13018 (N_13018,N_12897,N_12853);
nand U13019 (N_13019,N_12883,N_12916);
xor U13020 (N_13020,N_12984,N_12906);
and U13021 (N_13021,N_12917,N_12919);
or U13022 (N_13022,N_12908,N_12977);
xnor U13023 (N_13023,N_12818,N_12899);
nor U13024 (N_13024,N_12841,N_12869);
xnor U13025 (N_13025,N_12852,N_12820);
nand U13026 (N_13026,N_12929,N_12957);
nor U13027 (N_13027,N_12981,N_12817);
nand U13028 (N_13028,N_12849,N_12861);
or U13029 (N_13029,N_12952,N_12892);
and U13030 (N_13030,N_12879,N_12928);
xor U13031 (N_13031,N_12898,N_12813);
nor U13032 (N_13032,N_12846,N_12987);
or U13033 (N_13033,N_12878,N_12909);
and U13034 (N_13034,N_12800,N_12876);
or U13035 (N_13035,N_12905,N_12896);
or U13036 (N_13036,N_12833,N_12913);
nor U13037 (N_13037,N_12915,N_12974);
nor U13038 (N_13038,N_12966,N_12976);
or U13039 (N_13039,N_12866,N_12979);
nand U13040 (N_13040,N_12888,N_12868);
and U13041 (N_13041,N_12807,N_12900);
nand U13042 (N_13042,N_12812,N_12814);
and U13043 (N_13043,N_12985,N_12951);
xnor U13044 (N_13044,N_12873,N_12856);
and U13045 (N_13045,N_12930,N_12884);
or U13046 (N_13046,N_12848,N_12998);
nor U13047 (N_13047,N_12825,N_12864);
nor U13048 (N_13048,N_12978,N_12983);
xnor U13049 (N_13049,N_12842,N_12895);
nor U13050 (N_13050,N_12969,N_12982);
xor U13051 (N_13051,N_12991,N_12988);
nand U13052 (N_13052,N_12815,N_12964);
or U13053 (N_13053,N_12845,N_12931);
nor U13054 (N_13054,N_12862,N_12953);
or U13055 (N_13055,N_12828,N_12962);
xor U13056 (N_13056,N_12882,N_12949);
nand U13057 (N_13057,N_12801,N_12858);
nor U13058 (N_13058,N_12875,N_12989);
xnor U13059 (N_13059,N_12885,N_12874);
xor U13060 (N_13060,N_12901,N_12922);
and U13061 (N_13061,N_12986,N_12822);
nor U13062 (N_13062,N_12926,N_12939);
xnor U13063 (N_13063,N_12955,N_12890);
xnor U13064 (N_13064,N_12993,N_12990);
nor U13065 (N_13065,N_12850,N_12925);
nand U13066 (N_13066,N_12865,N_12963);
nand U13067 (N_13067,N_12910,N_12970);
nor U13068 (N_13068,N_12840,N_12903);
nor U13069 (N_13069,N_12997,N_12946);
xor U13070 (N_13070,N_12867,N_12994);
nor U13071 (N_13071,N_12940,N_12880);
nand U13072 (N_13072,N_12847,N_12832);
nand U13073 (N_13073,N_12961,N_12808);
nand U13074 (N_13074,N_12839,N_12843);
nand U13075 (N_13075,N_12891,N_12934);
nand U13076 (N_13076,N_12920,N_12947);
xor U13077 (N_13077,N_12819,N_12937);
nand U13078 (N_13078,N_12889,N_12821);
or U13079 (N_13079,N_12834,N_12971);
or U13080 (N_13080,N_12968,N_12887);
nand U13081 (N_13081,N_12975,N_12871);
nand U13082 (N_13082,N_12870,N_12823);
nor U13083 (N_13083,N_12936,N_12932);
and U13084 (N_13084,N_12995,N_12999);
and U13085 (N_13085,N_12912,N_12907);
or U13086 (N_13086,N_12958,N_12802);
nand U13087 (N_13087,N_12816,N_12924);
nor U13088 (N_13088,N_12830,N_12956);
or U13089 (N_13089,N_12942,N_12827);
xor U13090 (N_13090,N_12824,N_12881);
nand U13091 (N_13091,N_12810,N_12933);
or U13092 (N_13092,N_12851,N_12965);
xor U13093 (N_13093,N_12904,N_12950);
xnor U13094 (N_13094,N_12935,N_12894);
or U13095 (N_13095,N_12877,N_12911);
and U13096 (N_13096,N_12921,N_12967);
and U13097 (N_13097,N_12803,N_12805);
xor U13098 (N_13098,N_12855,N_12960);
or U13099 (N_13099,N_12943,N_12844);
or U13100 (N_13100,N_12877,N_12837);
or U13101 (N_13101,N_12871,N_12812);
and U13102 (N_13102,N_12835,N_12896);
xor U13103 (N_13103,N_12827,N_12839);
xor U13104 (N_13104,N_12995,N_12818);
nand U13105 (N_13105,N_12865,N_12854);
nor U13106 (N_13106,N_12948,N_12879);
nor U13107 (N_13107,N_12840,N_12824);
xor U13108 (N_13108,N_12839,N_12950);
or U13109 (N_13109,N_12901,N_12935);
xnor U13110 (N_13110,N_12871,N_12832);
and U13111 (N_13111,N_12807,N_12881);
or U13112 (N_13112,N_12889,N_12962);
nor U13113 (N_13113,N_12863,N_12875);
xnor U13114 (N_13114,N_12956,N_12843);
xnor U13115 (N_13115,N_12889,N_12960);
xor U13116 (N_13116,N_12918,N_12946);
xor U13117 (N_13117,N_12904,N_12858);
nand U13118 (N_13118,N_12899,N_12991);
nand U13119 (N_13119,N_12865,N_12927);
xor U13120 (N_13120,N_12850,N_12881);
xor U13121 (N_13121,N_12976,N_12969);
nor U13122 (N_13122,N_12812,N_12948);
and U13123 (N_13123,N_12917,N_12857);
and U13124 (N_13124,N_12924,N_12845);
nand U13125 (N_13125,N_12957,N_12845);
nor U13126 (N_13126,N_12861,N_12824);
xor U13127 (N_13127,N_12832,N_12977);
or U13128 (N_13128,N_12891,N_12829);
xnor U13129 (N_13129,N_12815,N_12831);
nand U13130 (N_13130,N_12955,N_12944);
nor U13131 (N_13131,N_12976,N_12907);
xnor U13132 (N_13132,N_12937,N_12942);
nor U13133 (N_13133,N_12849,N_12954);
nor U13134 (N_13134,N_12984,N_12971);
nor U13135 (N_13135,N_12957,N_12921);
xnor U13136 (N_13136,N_12978,N_12846);
nand U13137 (N_13137,N_12884,N_12941);
nor U13138 (N_13138,N_12878,N_12984);
or U13139 (N_13139,N_12871,N_12823);
or U13140 (N_13140,N_12905,N_12879);
nand U13141 (N_13141,N_12961,N_12903);
and U13142 (N_13142,N_12963,N_12938);
and U13143 (N_13143,N_12876,N_12830);
nor U13144 (N_13144,N_12822,N_12977);
or U13145 (N_13145,N_12937,N_12838);
and U13146 (N_13146,N_12886,N_12813);
nand U13147 (N_13147,N_12958,N_12993);
nor U13148 (N_13148,N_12957,N_12964);
nor U13149 (N_13149,N_12941,N_12874);
and U13150 (N_13150,N_12963,N_12983);
and U13151 (N_13151,N_12936,N_12868);
xnor U13152 (N_13152,N_12863,N_12900);
and U13153 (N_13153,N_12859,N_12886);
nand U13154 (N_13154,N_12906,N_12958);
nor U13155 (N_13155,N_12887,N_12933);
xnor U13156 (N_13156,N_12887,N_12873);
xor U13157 (N_13157,N_12975,N_12913);
xor U13158 (N_13158,N_12894,N_12855);
xor U13159 (N_13159,N_12955,N_12885);
and U13160 (N_13160,N_12805,N_12915);
or U13161 (N_13161,N_12930,N_12894);
nor U13162 (N_13162,N_12817,N_12957);
nor U13163 (N_13163,N_12854,N_12993);
nor U13164 (N_13164,N_12886,N_12984);
nand U13165 (N_13165,N_12802,N_12986);
nor U13166 (N_13166,N_12964,N_12855);
nand U13167 (N_13167,N_12871,N_12923);
or U13168 (N_13168,N_12813,N_12958);
and U13169 (N_13169,N_12949,N_12894);
xnor U13170 (N_13170,N_12926,N_12885);
nand U13171 (N_13171,N_12843,N_12878);
or U13172 (N_13172,N_12909,N_12948);
xnor U13173 (N_13173,N_12844,N_12849);
nand U13174 (N_13174,N_12919,N_12871);
nor U13175 (N_13175,N_12948,N_12848);
nor U13176 (N_13176,N_12916,N_12939);
or U13177 (N_13177,N_12995,N_12966);
nor U13178 (N_13178,N_12960,N_12832);
and U13179 (N_13179,N_12831,N_12872);
xnor U13180 (N_13180,N_12909,N_12967);
or U13181 (N_13181,N_12837,N_12811);
nor U13182 (N_13182,N_12820,N_12825);
xnor U13183 (N_13183,N_12862,N_12955);
xnor U13184 (N_13184,N_12946,N_12994);
or U13185 (N_13185,N_12842,N_12810);
or U13186 (N_13186,N_12860,N_12813);
xnor U13187 (N_13187,N_12906,N_12887);
nand U13188 (N_13188,N_12896,N_12852);
and U13189 (N_13189,N_12841,N_12931);
nand U13190 (N_13190,N_12815,N_12892);
or U13191 (N_13191,N_12980,N_12895);
nor U13192 (N_13192,N_12954,N_12953);
nor U13193 (N_13193,N_12869,N_12963);
xnor U13194 (N_13194,N_12857,N_12979);
nand U13195 (N_13195,N_12905,N_12988);
nand U13196 (N_13196,N_12953,N_12869);
nand U13197 (N_13197,N_12953,N_12854);
nand U13198 (N_13198,N_12849,N_12986);
nor U13199 (N_13199,N_12880,N_12861);
and U13200 (N_13200,N_13107,N_13009);
nand U13201 (N_13201,N_13152,N_13025);
nor U13202 (N_13202,N_13189,N_13002);
nand U13203 (N_13203,N_13068,N_13190);
nor U13204 (N_13204,N_13125,N_13140);
nor U13205 (N_13205,N_13003,N_13163);
or U13206 (N_13206,N_13134,N_13011);
xnor U13207 (N_13207,N_13085,N_13071);
and U13208 (N_13208,N_13067,N_13102);
nand U13209 (N_13209,N_13058,N_13130);
and U13210 (N_13210,N_13162,N_13165);
or U13211 (N_13211,N_13166,N_13147);
nand U13212 (N_13212,N_13059,N_13041);
xnor U13213 (N_13213,N_13031,N_13176);
and U13214 (N_13214,N_13052,N_13061);
or U13215 (N_13215,N_13108,N_13132);
nand U13216 (N_13216,N_13048,N_13167);
or U13217 (N_13217,N_13157,N_13136);
nand U13218 (N_13218,N_13191,N_13019);
or U13219 (N_13219,N_13083,N_13184);
and U13220 (N_13220,N_13076,N_13032);
or U13221 (N_13221,N_13103,N_13001);
or U13222 (N_13222,N_13013,N_13036);
or U13223 (N_13223,N_13123,N_13151);
nor U13224 (N_13224,N_13155,N_13110);
nor U13225 (N_13225,N_13017,N_13042);
and U13226 (N_13226,N_13137,N_13075);
or U13227 (N_13227,N_13006,N_13100);
nand U13228 (N_13228,N_13038,N_13033);
or U13229 (N_13229,N_13084,N_13158);
nor U13230 (N_13230,N_13012,N_13142);
nor U13231 (N_13231,N_13092,N_13024);
xor U13232 (N_13232,N_13004,N_13112);
nor U13233 (N_13233,N_13069,N_13007);
and U13234 (N_13234,N_13104,N_13049);
nor U13235 (N_13235,N_13192,N_13141);
nor U13236 (N_13236,N_13156,N_13015);
nor U13237 (N_13237,N_13118,N_13060);
and U13238 (N_13238,N_13078,N_13050);
nor U13239 (N_13239,N_13139,N_13154);
nor U13240 (N_13240,N_13077,N_13131);
nor U13241 (N_13241,N_13037,N_13129);
xor U13242 (N_13242,N_13095,N_13128);
or U13243 (N_13243,N_13117,N_13090);
and U13244 (N_13244,N_13010,N_13040);
or U13245 (N_13245,N_13096,N_13093);
nor U13246 (N_13246,N_13105,N_13080);
or U13247 (N_13247,N_13113,N_13046);
xor U13248 (N_13248,N_13020,N_13047);
xnor U13249 (N_13249,N_13063,N_13028);
or U13250 (N_13250,N_13062,N_13044);
xnor U13251 (N_13251,N_13122,N_13175);
nand U13252 (N_13252,N_13111,N_13149);
or U13253 (N_13253,N_13144,N_13014);
and U13254 (N_13254,N_13022,N_13053);
nor U13255 (N_13255,N_13194,N_13043);
or U13256 (N_13256,N_13146,N_13180);
xnor U13257 (N_13257,N_13164,N_13109);
xnor U13258 (N_13258,N_13018,N_13055);
xor U13259 (N_13259,N_13121,N_13196);
nand U13260 (N_13260,N_13116,N_13072);
and U13261 (N_13261,N_13161,N_13101);
nand U13262 (N_13262,N_13150,N_13115);
nand U13263 (N_13263,N_13119,N_13021);
nand U13264 (N_13264,N_13073,N_13000);
or U13265 (N_13265,N_13098,N_13120);
nor U13266 (N_13266,N_13088,N_13126);
or U13267 (N_13267,N_13057,N_13193);
nand U13268 (N_13268,N_13135,N_13099);
xor U13269 (N_13269,N_13133,N_13185);
nand U13270 (N_13270,N_13081,N_13169);
nand U13271 (N_13271,N_13064,N_13181);
or U13272 (N_13272,N_13089,N_13039);
or U13273 (N_13273,N_13074,N_13198);
and U13274 (N_13274,N_13091,N_13186);
and U13275 (N_13275,N_13160,N_13127);
or U13276 (N_13276,N_13082,N_13051);
or U13277 (N_13277,N_13029,N_13183);
nor U13278 (N_13278,N_13056,N_13023);
or U13279 (N_13279,N_13027,N_13035);
xnor U13280 (N_13280,N_13177,N_13016);
nor U13281 (N_13281,N_13026,N_13030);
xor U13282 (N_13282,N_13079,N_13195);
and U13283 (N_13283,N_13173,N_13045);
or U13284 (N_13284,N_13106,N_13066);
nand U13285 (N_13285,N_13187,N_13086);
and U13286 (N_13286,N_13065,N_13178);
nor U13287 (N_13287,N_13168,N_13199);
and U13288 (N_13288,N_13145,N_13174);
or U13289 (N_13289,N_13124,N_13170);
xnor U13290 (N_13290,N_13172,N_13054);
or U13291 (N_13291,N_13094,N_13034);
and U13292 (N_13292,N_13008,N_13159);
xnor U13293 (N_13293,N_13097,N_13143);
and U13294 (N_13294,N_13114,N_13197);
nand U13295 (N_13295,N_13182,N_13188);
nand U13296 (N_13296,N_13005,N_13070);
xnor U13297 (N_13297,N_13138,N_13148);
xor U13298 (N_13298,N_13153,N_13087);
and U13299 (N_13299,N_13171,N_13179);
nor U13300 (N_13300,N_13131,N_13027);
and U13301 (N_13301,N_13115,N_13157);
xnor U13302 (N_13302,N_13087,N_13139);
xor U13303 (N_13303,N_13004,N_13186);
and U13304 (N_13304,N_13024,N_13043);
or U13305 (N_13305,N_13118,N_13088);
nor U13306 (N_13306,N_13071,N_13161);
xnor U13307 (N_13307,N_13136,N_13127);
nand U13308 (N_13308,N_13181,N_13066);
or U13309 (N_13309,N_13044,N_13054);
xnor U13310 (N_13310,N_13048,N_13150);
xor U13311 (N_13311,N_13016,N_13050);
or U13312 (N_13312,N_13161,N_13018);
or U13313 (N_13313,N_13140,N_13022);
nand U13314 (N_13314,N_13062,N_13101);
nor U13315 (N_13315,N_13080,N_13037);
nor U13316 (N_13316,N_13095,N_13048);
nor U13317 (N_13317,N_13062,N_13060);
nand U13318 (N_13318,N_13006,N_13108);
or U13319 (N_13319,N_13131,N_13148);
nand U13320 (N_13320,N_13154,N_13103);
nor U13321 (N_13321,N_13139,N_13014);
nor U13322 (N_13322,N_13004,N_13095);
xor U13323 (N_13323,N_13056,N_13048);
xor U13324 (N_13324,N_13061,N_13119);
nor U13325 (N_13325,N_13177,N_13068);
or U13326 (N_13326,N_13050,N_13091);
and U13327 (N_13327,N_13065,N_13016);
nand U13328 (N_13328,N_13165,N_13031);
nor U13329 (N_13329,N_13049,N_13178);
nor U13330 (N_13330,N_13021,N_13054);
nand U13331 (N_13331,N_13169,N_13125);
and U13332 (N_13332,N_13161,N_13140);
nand U13333 (N_13333,N_13066,N_13198);
nand U13334 (N_13334,N_13122,N_13193);
xor U13335 (N_13335,N_13019,N_13158);
or U13336 (N_13336,N_13166,N_13131);
xor U13337 (N_13337,N_13037,N_13178);
and U13338 (N_13338,N_13141,N_13081);
nand U13339 (N_13339,N_13109,N_13137);
and U13340 (N_13340,N_13064,N_13161);
or U13341 (N_13341,N_13167,N_13182);
or U13342 (N_13342,N_13106,N_13176);
nand U13343 (N_13343,N_13187,N_13199);
xnor U13344 (N_13344,N_13183,N_13005);
and U13345 (N_13345,N_13034,N_13192);
or U13346 (N_13346,N_13196,N_13093);
nor U13347 (N_13347,N_13057,N_13067);
and U13348 (N_13348,N_13105,N_13040);
xnor U13349 (N_13349,N_13088,N_13170);
or U13350 (N_13350,N_13087,N_13137);
nand U13351 (N_13351,N_13110,N_13003);
xor U13352 (N_13352,N_13153,N_13174);
nor U13353 (N_13353,N_13168,N_13072);
nor U13354 (N_13354,N_13120,N_13058);
or U13355 (N_13355,N_13132,N_13067);
nor U13356 (N_13356,N_13081,N_13048);
xnor U13357 (N_13357,N_13138,N_13069);
and U13358 (N_13358,N_13120,N_13087);
nor U13359 (N_13359,N_13099,N_13012);
nor U13360 (N_13360,N_13015,N_13031);
and U13361 (N_13361,N_13074,N_13195);
or U13362 (N_13362,N_13149,N_13092);
or U13363 (N_13363,N_13074,N_13090);
or U13364 (N_13364,N_13128,N_13065);
and U13365 (N_13365,N_13132,N_13002);
xnor U13366 (N_13366,N_13182,N_13053);
and U13367 (N_13367,N_13028,N_13048);
nor U13368 (N_13368,N_13190,N_13121);
and U13369 (N_13369,N_13129,N_13067);
nand U13370 (N_13370,N_13188,N_13022);
nor U13371 (N_13371,N_13075,N_13045);
xor U13372 (N_13372,N_13157,N_13001);
nand U13373 (N_13373,N_13071,N_13107);
or U13374 (N_13374,N_13197,N_13055);
xor U13375 (N_13375,N_13102,N_13025);
or U13376 (N_13376,N_13067,N_13177);
and U13377 (N_13377,N_13001,N_13197);
or U13378 (N_13378,N_13142,N_13019);
nand U13379 (N_13379,N_13189,N_13060);
or U13380 (N_13380,N_13042,N_13108);
or U13381 (N_13381,N_13144,N_13012);
nand U13382 (N_13382,N_13159,N_13011);
nor U13383 (N_13383,N_13070,N_13051);
xor U13384 (N_13384,N_13060,N_13031);
nor U13385 (N_13385,N_13020,N_13011);
and U13386 (N_13386,N_13119,N_13095);
and U13387 (N_13387,N_13067,N_13133);
and U13388 (N_13388,N_13170,N_13110);
or U13389 (N_13389,N_13121,N_13092);
and U13390 (N_13390,N_13065,N_13022);
xor U13391 (N_13391,N_13181,N_13012);
or U13392 (N_13392,N_13145,N_13025);
nor U13393 (N_13393,N_13040,N_13057);
nor U13394 (N_13394,N_13040,N_13115);
nand U13395 (N_13395,N_13176,N_13042);
xor U13396 (N_13396,N_13023,N_13126);
nand U13397 (N_13397,N_13051,N_13100);
or U13398 (N_13398,N_13043,N_13087);
nor U13399 (N_13399,N_13120,N_13036);
or U13400 (N_13400,N_13393,N_13271);
nor U13401 (N_13401,N_13363,N_13315);
nor U13402 (N_13402,N_13298,N_13341);
or U13403 (N_13403,N_13381,N_13370);
nor U13404 (N_13404,N_13226,N_13246);
nand U13405 (N_13405,N_13277,N_13361);
nor U13406 (N_13406,N_13220,N_13203);
or U13407 (N_13407,N_13338,N_13222);
xor U13408 (N_13408,N_13373,N_13229);
nor U13409 (N_13409,N_13334,N_13335);
nand U13410 (N_13410,N_13319,N_13254);
and U13411 (N_13411,N_13245,N_13325);
xnor U13412 (N_13412,N_13297,N_13251);
or U13413 (N_13413,N_13336,N_13244);
and U13414 (N_13414,N_13202,N_13378);
nor U13415 (N_13415,N_13322,N_13377);
xor U13416 (N_13416,N_13265,N_13279);
xnor U13417 (N_13417,N_13309,N_13206);
xnor U13418 (N_13418,N_13369,N_13347);
xnor U13419 (N_13419,N_13293,N_13337);
nor U13420 (N_13420,N_13273,N_13362);
xor U13421 (N_13421,N_13349,N_13212);
nand U13422 (N_13422,N_13204,N_13283);
xnor U13423 (N_13423,N_13234,N_13323);
nand U13424 (N_13424,N_13224,N_13300);
and U13425 (N_13425,N_13238,N_13386);
xor U13426 (N_13426,N_13215,N_13385);
xor U13427 (N_13427,N_13372,N_13270);
and U13428 (N_13428,N_13321,N_13328);
and U13429 (N_13429,N_13258,N_13289);
and U13430 (N_13430,N_13342,N_13213);
nand U13431 (N_13431,N_13272,N_13307);
xnor U13432 (N_13432,N_13350,N_13292);
nor U13433 (N_13433,N_13299,N_13324);
or U13434 (N_13434,N_13313,N_13312);
or U13435 (N_13435,N_13262,N_13382);
nand U13436 (N_13436,N_13329,N_13353);
or U13437 (N_13437,N_13388,N_13276);
nand U13438 (N_13438,N_13242,N_13354);
xor U13439 (N_13439,N_13290,N_13318);
or U13440 (N_13440,N_13291,N_13376);
or U13441 (N_13441,N_13383,N_13201);
xnor U13442 (N_13442,N_13379,N_13239);
xnor U13443 (N_13443,N_13394,N_13264);
xor U13444 (N_13444,N_13227,N_13331);
and U13445 (N_13445,N_13345,N_13305);
nand U13446 (N_13446,N_13384,N_13282);
xnor U13447 (N_13447,N_13236,N_13285);
nand U13448 (N_13448,N_13301,N_13281);
and U13449 (N_13449,N_13266,N_13374);
and U13450 (N_13450,N_13219,N_13340);
or U13451 (N_13451,N_13274,N_13294);
nand U13452 (N_13452,N_13397,N_13314);
and U13453 (N_13453,N_13303,N_13233);
or U13454 (N_13454,N_13398,N_13320);
or U13455 (N_13455,N_13333,N_13352);
and U13456 (N_13456,N_13280,N_13359);
and U13457 (N_13457,N_13356,N_13217);
and U13458 (N_13458,N_13228,N_13232);
xnor U13459 (N_13459,N_13267,N_13390);
xor U13460 (N_13460,N_13387,N_13216);
xnor U13461 (N_13461,N_13346,N_13344);
nor U13462 (N_13462,N_13207,N_13278);
nor U13463 (N_13463,N_13210,N_13259);
nor U13464 (N_13464,N_13371,N_13308);
and U13465 (N_13465,N_13235,N_13286);
and U13466 (N_13466,N_13360,N_13358);
nor U13467 (N_13467,N_13348,N_13256);
and U13468 (N_13468,N_13351,N_13392);
or U13469 (N_13469,N_13316,N_13296);
xnor U13470 (N_13470,N_13241,N_13218);
nor U13471 (N_13471,N_13339,N_13306);
nor U13472 (N_13472,N_13399,N_13368);
xnor U13473 (N_13473,N_13330,N_13249);
nand U13474 (N_13474,N_13243,N_13260);
and U13475 (N_13475,N_13357,N_13327);
or U13476 (N_13476,N_13275,N_13302);
nor U13477 (N_13477,N_13326,N_13252);
or U13478 (N_13478,N_13288,N_13223);
or U13479 (N_13479,N_13311,N_13263);
or U13480 (N_13480,N_13211,N_13250);
or U13481 (N_13481,N_13284,N_13389);
nor U13482 (N_13482,N_13221,N_13255);
nor U13483 (N_13483,N_13209,N_13230);
nand U13484 (N_13484,N_13332,N_13317);
xnor U13485 (N_13485,N_13231,N_13364);
nand U13486 (N_13486,N_13240,N_13375);
or U13487 (N_13487,N_13205,N_13380);
or U13488 (N_13488,N_13365,N_13225);
or U13489 (N_13489,N_13257,N_13391);
nand U13490 (N_13490,N_13304,N_13367);
nand U13491 (N_13491,N_13310,N_13268);
xor U13492 (N_13492,N_13237,N_13287);
xor U13493 (N_13493,N_13247,N_13261);
or U13494 (N_13494,N_13366,N_13396);
nand U13495 (N_13495,N_13200,N_13208);
nor U13496 (N_13496,N_13355,N_13248);
and U13497 (N_13497,N_13343,N_13395);
and U13498 (N_13498,N_13214,N_13253);
or U13499 (N_13499,N_13269,N_13295);
or U13500 (N_13500,N_13270,N_13295);
xor U13501 (N_13501,N_13290,N_13356);
nor U13502 (N_13502,N_13337,N_13363);
xor U13503 (N_13503,N_13277,N_13390);
and U13504 (N_13504,N_13238,N_13381);
nand U13505 (N_13505,N_13296,N_13267);
nor U13506 (N_13506,N_13342,N_13230);
nand U13507 (N_13507,N_13356,N_13264);
nor U13508 (N_13508,N_13372,N_13319);
nand U13509 (N_13509,N_13321,N_13327);
nor U13510 (N_13510,N_13321,N_13315);
xnor U13511 (N_13511,N_13341,N_13229);
and U13512 (N_13512,N_13228,N_13373);
nor U13513 (N_13513,N_13206,N_13222);
xnor U13514 (N_13514,N_13396,N_13387);
and U13515 (N_13515,N_13346,N_13298);
or U13516 (N_13516,N_13314,N_13368);
or U13517 (N_13517,N_13250,N_13322);
or U13518 (N_13518,N_13399,N_13210);
and U13519 (N_13519,N_13297,N_13373);
or U13520 (N_13520,N_13365,N_13236);
or U13521 (N_13521,N_13264,N_13204);
and U13522 (N_13522,N_13278,N_13393);
xor U13523 (N_13523,N_13318,N_13283);
xor U13524 (N_13524,N_13340,N_13210);
nand U13525 (N_13525,N_13329,N_13338);
xor U13526 (N_13526,N_13367,N_13313);
or U13527 (N_13527,N_13399,N_13357);
xnor U13528 (N_13528,N_13256,N_13231);
or U13529 (N_13529,N_13206,N_13331);
nand U13530 (N_13530,N_13364,N_13368);
nor U13531 (N_13531,N_13287,N_13289);
nor U13532 (N_13532,N_13244,N_13206);
or U13533 (N_13533,N_13200,N_13243);
xor U13534 (N_13534,N_13377,N_13357);
or U13535 (N_13535,N_13323,N_13207);
xor U13536 (N_13536,N_13298,N_13260);
nor U13537 (N_13537,N_13240,N_13350);
xor U13538 (N_13538,N_13228,N_13387);
nand U13539 (N_13539,N_13250,N_13348);
and U13540 (N_13540,N_13234,N_13364);
and U13541 (N_13541,N_13385,N_13332);
and U13542 (N_13542,N_13397,N_13234);
nand U13543 (N_13543,N_13266,N_13384);
or U13544 (N_13544,N_13365,N_13268);
or U13545 (N_13545,N_13307,N_13212);
and U13546 (N_13546,N_13353,N_13393);
xor U13547 (N_13547,N_13249,N_13329);
nand U13548 (N_13548,N_13354,N_13308);
xor U13549 (N_13549,N_13307,N_13331);
nand U13550 (N_13550,N_13377,N_13361);
xor U13551 (N_13551,N_13364,N_13251);
and U13552 (N_13552,N_13237,N_13278);
or U13553 (N_13553,N_13218,N_13237);
nand U13554 (N_13554,N_13360,N_13274);
and U13555 (N_13555,N_13303,N_13240);
and U13556 (N_13556,N_13221,N_13323);
or U13557 (N_13557,N_13250,N_13390);
and U13558 (N_13558,N_13207,N_13287);
and U13559 (N_13559,N_13286,N_13227);
or U13560 (N_13560,N_13395,N_13227);
xor U13561 (N_13561,N_13208,N_13278);
or U13562 (N_13562,N_13305,N_13244);
xnor U13563 (N_13563,N_13222,N_13269);
xnor U13564 (N_13564,N_13232,N_13376);
nand U13565 (N_13565,N_13292,N_13331);
nand U13566 (N_13566,N_13242,N_13303);
nor U13567 (N_13567,N_13364,N_13221);
nand U13568 (N_13568,N_13345,N_13331);
nand U13569 (N_13569,N_13258,N_13343);
or U13570 (N_13570,N_13399,N_13244);
or U13571 (N_13571,N_13392,N_13357);
nand U13572 (N_13572,N_13300,N_13231);
or U13573 (N_13573,N_13218,N_13355);
and U13574 (N_13574,N_13312,N_13291);
or U13575 (N_13575,N_13307,N_13260);
nand U13576 (N_13576,N_13383,N_13392);
or U13577 (N_13577,N_13375,N_13282);
or U13578 (N_13578,N_13383,N_13239);
and U13579 (N_13579,N_13398,N_13326);
xor U13580 (N_13580,N_13390,N_13330);
or U13581 (N_13581,N_13381,N_13274);
and U13582 (N_13582,N_13343,N_13312);
nand U13583 (N_13583,N_13297,N_13212);
and U13584 (N_13584,N_13257,N_13221);
or U13585 (N_13585,N_13234,N_13367);
nand U13586 (N_13586,N_13326,N_13298);
nand U13587 (N_13587,N_13373,N_13342);
or U13588 (N_13588,N_13359,N_13252);
or U13589 (N_13589,N_13298,N_13217);
nand U13590 (N_13590,N_13357,N_13207);
nand U13591 (N_13591,N_13321,N_13284);
and U13592 (N_13592,N_13389,N_13323);
nor U13593 (N_13593,N_13305,N_13384);
xnor U13594 (N_13594,N_13392,N_13269);
xnor U13595 (N_13595,N_13355,N_13212);
xnor U13596 (N_13596,N_13205,N_13213);
nor U13597 (N_13597,N_13235,N_13370);
nand U13598 (N_13598,N_13348,N_13325);
or U13599 (N_13599,N_13367,N_13350);
xnor U13600 (N_13600,N_13545,N_13471);
nand U13601 (N_13601,N_13590,N_13580);
or U13602 (N_13602,N_13475,N_13510);
and U13603 (N_13603,N_13542,N_13478);
xor U13604 (N_13604,N_13522,N_13430);
xnor U13605 (N_13605,N_13455,N_13581);
and U13606 (N_13606,N_13418,N_13578);
xor U13607 (N_13607,N_13498,N_13408);
xnor U13608 (N_13608,N_13440,N_13537);
nand U13609 (N_13609,N_13520,N_13548);
and U13610 (N_13610,N_13555,N_13492);
and U13611 (N_13611,N_13579,N_13420);
xor U13612 (N_13612,N_13469,N_13525);
nor U13613 (N_13613,N_13495,N_13532);
and U13614 (N_13614,N_13444,N_13477);
and U13615 (N_13615,N_13423,N_13547);
nor U13616 (N_13616,N_13415,N_13509);
and U13617 (N_13617,N_13587,N_13527);
nor U13618 (N_13618,N_13445,N_13557);
or U13619 (N_13619,N_13493,N_13565);
xnor U13620 (N_13620,N_13464,N_13480);
nand U13621 (N_13621,N_13403,N_13530);
and U13622 (N_13622,N_13436,N_13531);
nand U13623 (N_13623,N_13550,N_13459);
nor U13624 (N_13624,N_13597,N_13570);
and U13625 (N_13625,N_13473,N_13448);
xor U13626 (N_13626,N_13504,N_13465);
and U13627 (N_13627,N_13515,N_13472);
nand U13628 (N_13628,N_13512,N_13529);
and U13629 (N_13629,N_13558,N_13588);
nor U13630 (N_13630,N_13425,N_13576);
xnor U13631 (N_13631,N_13567,N_13483);
xor U13632 (N_13632,N_13589,N_13407);
nand U13633 (N_13633,N_13596,N_13563);
or U13634 (N_13634,N_13461,N_13466);
and U13635 (N_13635,N_13595,N_13534);
nand U13636 (N_13636,N_13426,N_13553);
or U13637 (N_13637,N_13442,N_13546);
and U13638 (N_13638,N_13412,N_13541);
or U13639 (N_13639,N_13583,N_13561);
nor U13640 (N_13640,N_13457,N_13552);
or U13641 (N_13641,N_13574,N_13406);
and U13642 (N_13642,N_13454,N_13584);
or U13643 (N_13643,N_13593,N_13462);
or U13644 (N_13644,N_13439,N_13599);
or U13645 (N_13645,N_13435,N_13433);
nor U13646 (N_13646,N_13488,N_13421);
xor U13647 (N_13647,N_13571,N_13463);
or U13648 (N_13648,N_13487,N_13416);
xor U13649 (N_13649,N_13559,N_13564);
xnor U13650 (N_13650,N_13479,N_13538);
nand U13651 (N_13651,N_13575,N_13400);
nand U13652 (N_13652,N_13511,N_13517);
and U13653 (N_13653,N_13404,N_13486);
and U13654 (N_13654,N_13437,N_13535);
and U13655 (N_13655,N_13566,N_13491);
or U13656 (N_13656,N_13401,N_13447);
nand U13657 (N_13657,N_13499,N_13544);
xnor U13658 (N_13658,N_13526,N_13503);
nand U13659 (N_13659,N_13524,N_13470);
xnor U13660 (N_13660,N_13556,N_13539);
xnor U13661 (N_13661,N_13452,N_13568);
nand U13662 (N_13662,N_13496,N_13409);
nand U13663 (N_13663,N_13540,N_13536);
xnor U13664 (N_13664,N_13573,N_13419);
nor U13665 (N_13665,N_13572,N_13598);
nand U13666 (N_13666,N_13582,N_13489);
nand U13667 (N_13667,N_13577,N_13482);
nor U13668 (N_13668,N_13458,N_13521);
nor U13669 (N_13669,N_13446,N_13453);
nor U13670 (N_13670,N_13451,N_13481);
nand U13671 (N_13671,N_13560,N_13506);
and U13672 (N_13672,N_13410,N_13424);
and U13673 (N_13673,N_13497,N_13562);
or U13674 (N_13674,N_13502,N_13476);
nand U13675 (N_13675,N_13591,N_13594);
nand U13676 (N_13676,N_13468,N_13438);
xor U13677 (N_13677,N_13528,N_13449);
nand U13678 (N_13678,N_13441,N_13405);
or U13679 (N_13679,N_13585,N_13514);
or U13680 (N_13680,N_13413,N_13427);
nand U13681 (N_13681,N_13505,N_13474);
and U13682 (N_13682,N_13516,N_13428);
nor U13683 (N_13683,N_13569,N_13443);
nand U13684 (N_13684,N_13519,N_13414);
or U13685 (N_13685,N_13543,N_13554);
and U13686 (N_13686,N_13485,N_13508);
or U13687 (N_13687,N_13500,N_13484);
xnor U13688 (N_13688,N_13429,N_13586);
and U13689 (N_13689,N_13551,N_13494);
or U13690 (N_13690,N_13450,N_13507);
and U13691 (N_13691,N_13592,N_13411);
nor U13692 (N_13692,N_13518,N_13467);
xnor U13693 (N_13693,N_13456,N_13490);
or U13694 (N_13694,N_13431,N_13402);
nor U13695 (N_13695,N_13523,N_13501);
xor U13696 (N_13696,N_13422,N_13549);
or U13697 (N_13697,N_13417,N_13460);
nand U13698 (N_13698,N_13533,N_13513);
nor U13699 (N_13699,N_13434,N_13432);
nor U13700 (N_13700,N_13412,N_13451);
and U13701 (N_13701,N_13510,N_13598);
or U13702 (N_13702,N_13566,N_13404);
nor U13703 (N_13703,N_13549,N_13520);
nor U13704 (N_13704,N_13580,N_13519);
xor U13705 (N_13705,N_13461,N_13511);
or U13706 (N_13706,N_13591,N_13412);
and U13707 (N_13707,N_13410,N_13544);
and U13708 (N_13708,N_13554,N_13545);
xor U13709 (N_13709,N_13422,N_13560);
nor U13710 (N_13710,N_13428,N_13434);
xnor U13711 (N_13711,N_13578,N_13564);
nor U13712 (N_13712,N_13468,N_13515);
nand U13713 (N_13713,N_13514,N_13538);
xnor U13714 (N_13714,N_13599,N_13558);
nand U13715 (N_13715,N_13582,N_13421);
nand U13716 (N_13716,N_13571,N_13451);
nand U13717 (N_13717,N_13490,N_13459);
xor U13718 (N_13718,N_13551,N_13418);
xnor U13719 (N_13719,N_13403,N_13505);
nor U13720 (N_13720,N_13546,N_13429);
nor U13721 (N_13721,N_13595,N_13540);
or U13722 (N_13722,N_13426,N_13472);
xor U13723 (N_13723,N_13422,N_13500);
nor U13724 (N_13724,N_13537,N_13582);
and U13725 (N_13725,N_13553,N_13412);
nor U13726 (N_13726,N_13573,N_13556);
or U13727 (N_13727,N_13526,N_13420);
nand U13728 (N_13728,N_13557,N_13564);
and U13729 (N_13729,N_13497,N_13551);
nor U13730 (N_13730,N_13516,N_13421);
or U13731 (N_13731,N_13588,N_13586);
nor U13732 (N_13732,N_13501,N_13582);
or U13733 (N_13733,N_13596,N_13529);
nand U13734 (N_13734,N_13532,N_13482);
or U13735 (N_13735,N_13432,N_13467);
nor U13736 (N_13736,N_13411,N_13523);
xor U13737 (N_13737,N_13566,N_13591);
or U13738 (N_13738,N_13511,N_13541);
xor U13739 (N_13739,N_13490,N_13486);
and U13740 (N_13740,N_13439,N_13498);
or U13741 (N_13741,N_13419,N_13436);
nand U13742 (N_13742,N_13559,N_13586);
nor U13743 (N_13743,N_13424,N_13580);
nand U13744 (N_13744,N_13441,N_13410);
nor U13745 (N_13745,N_13592,N_13414);
nor U13746 (N_13746,N_13460,N_13554);
nand U13747 (N_13747,N_13596,N_13454);
nand U13748 (N_13748,N_13548,N_13523);
or U13749 (N_13749,N_13504,N_13493);
and U13750 (N_13750,N_13499,N_13537);
nand U13751 (N_13751,N_13485,N_13589);
xor U13752 (N_13752,N_13440,N_13437);
or U13753 (N_13753,N_13449,N_13520);
and U13754 (N_13754,N_13580,N_13531);
nor U13755 (N_13755,N_13479,N_13562);
and U13756 (N_13756,N_13582,N_13483);
nor U13757 (N_13757,N_13516,N_13508);
nor U13758 (N_13758,N_13415,N_13488);
and U13759 (N_13759,N_13494,N_13540);
or U13760 (N_13760,N_13585,N_13401);
or U13761 (N_13761,N_13573,N_13442);
nor U13762 (N_13762,N_13472,N_13516);
nand U13763 (N_13763,N_13578,N_13536);
xnor U13764 (N_13764,N_13517,N_13477);
nor U13765 (N_13765,N_13547,N_13450);
nand U13766 (N_13766,N_13503,N_13465);
xnor U13767 (N_13767,N_13593,N_13428);
xor U13768 (N_13768,N_13599,N_13446);
or U13769 (N_13769,N_13448,N_13518);
xor U13770 (N_13770,N_13585,N_13573);
or U13771 (N_13771,N_13508,N_13496);
and U13772 (N_13772,N_13479,N_13480);
nor U13773 (N_13773,N_13565,N_13445);
or U13774 (N_13774,N_13574,N_13499);
nor U13775 (N_13775,N_13597,N_13557);
xor U13776 (N_13776,N_13553,N_13551);
xnor U13777 (N_13777,N_13479,N_13543);
xnor U13778 (N_13778,N_13417,N_13598);
nand U13779 (N_13779,N_13432,N_13429);
and U13780 (N_13780,N_13528,N_13509);
nor U13781 (N_13781,N_13401,N_13421);
nand U13782 (N_13782,N_13411,N_13567);
and U13783 (N_13783,N_13560,N_13595);
xor U13784 (N_13784,N_13548,N_13410);
nand U13785 (N_13785,N_13402,N_13586);
nand U13786 (N_13786,N_13581,N_13410);
and U13787 (N_13787,N_13443,N_13417);
nand U13788 (N_13788,N_13544,N_13479);
and U13789 (N_13789,N_13448,N_13587);
nor U13790 (N_13790,N_13574,N_13562);
xnor U13791 (N_13791,N_13558,N_13426);
and U13792 (N_13792,N_13476,N_13478);
and U13793 (N_13793,N_13406,N_13579);
or U13794 (N_13794,N_13544,N_13553);
xor U13795 (N_13795,N_13443,N_13511);
and U13796 (N_13796,N_13579,N_13584);
nand U13797 (N_13797,N_13543,N_13478);
and U13798 (N_13798,N_13516,N_13519);
xor U13799 (N_13799,N_13593,N_13401);
or U13800 (N_13800,N_13661,N_13796);
and U13801 (N_13801,N_13617,N_13656);
and U13802 (N_13802,N_13709,N_13645);
or U13803 (N_13803,N_13689,N_13730);
nor U13804 (N_13804,N_13662,N_13680);
nor U13805 (N_13805,N_13708,N_13748);
nand U13806 (N_13806,N_13749,N_13695);
and U13807 (N_13807,N_13732,N_13764);
nand U13808 (N_13808,N_13757,N_13717);
and U13809 (N_13809,N_13774,N_13752);
nor U13810 (N_13810,N_13734,N_13690);
nor U13811 (N_13811,N_13642,N_13779);
or U13812 (N_13812,N_13616,N_13669);
and U13813 (N_13813,N_13753,N_13718);
and U13814 (N_13814,N_13737,N_13623);
xnor U13815 (N_13815,N_13784,N_13798);
and U13816 (N_13816,N_13769,N_13713);
or U13817 (N_13817,N_13776,N_13740);
nand U13818 (N_13818,N_13722,N_13791);
nor U13819 (N_13819,N_13610,N_13675);
nand U13820 (N_13820,N_13634,N_13787);
nand U13821 (N_13821,N_13723,N_13684);
xor U13822 (N_13822,N_13604,N_13668);
nor U13823 (N_13823,N_13758,N_13778);
nor U13824 (N_13824,N_13681,N_13697);
xor U13825 (N_13825,N_13724,N_13728);
xor U13826 (N_13826,N_13711,N_13712);
nand U13827 (N_13827,N_13636,N_13676);
xor U13828 (N_13828,N_13624,N_13739);
xnor U13829 (N_13829,N_13747,N_13630);
nand U13830 (N_13830,N_13729,N_13685);
or U13831 (N_13831,N_13647,N_13710);
xor U13832 (N_13832,N_13664,N_13614);
nand U13833 (N_13833,N_13750,N_13702);
nor U13834 (N_13834,N_13621,N_13657);
nor U13835 (N_13835,N_13782,N_13775);
nand U13836 (N_13836,N_13620,N_13666);
nand U13837 (N_13837,N_13738,N_13785);
nand U13838 (N_13838,N_13694,N_13635);
and U13839 (N_13839,N_13631,N_13673);
nor U13840 (N_13840,N_13660,N_13793);
and U13841 (N_13841,N_13726,N_13659);
and U13842 (N_13842,N_13772,N_13638);
nand U13843 (N_13843,N_13698,N_13742);
and U13844 (N_13844,N_13733,N_13612);
nand U13845 (N_13845,N_13692,N_13788);
nand U13846 (N_13846,N_13626,N_13688);
or U13847 (N_13847,N_13756,N_13780);
or U13848 (N_13848,N_13633,N_13672);
nor U13849 (N_13849,N_13651,N_13686);
or U13850 (N_13850,N_13608,N_13670);
nand U13851 (N_13851,N_13703,N_13767);
or U13852 (N_13852,N_13783,N_13683);
xnor U13853 (N_13853,N_13606,N_13605);
nor U13854 (N_13854,N_13607,N_13639);
xor U13855 (N_13855,N_13720,N_13637);
nand U13856 (N_13856,N_13762,N_13618);
nor U13857 (N_13857,N_13768,N_13601);
xnor U13858 (N_13858,N_13755,N_13736);
nand U13859 (N_13859,N_13705,N_13658);
nand U13860 (N_13860,N_13765,N_13627);
nor U13861 (N_13861,N_13629,N_13603);
and U13862 (N_13862,N_13699,N_13693);
or U13863 (N_13863,N_13632,N_13760);
nand U13864 (N_13864,N_13786,N_13679);
or U13865 (N_13865,N_13613,N_13719);
and U13866 (N_13866,N_13721,N_13714);
or U13867 (N_13867,N_13619,N_13687);
or U13868 (N_13868,N_13671,N_13770);
nand U13869 (N_13869,N_13655,N_13650);
xor U13870 (N_13870,N_13625,N_13715);
or U13871 (N_13871,N_13643,N_13746);
xnor U13872 (N_13872,N_13741,N_13761);
nand U13873 (N_13873,N_13790,N_13644);
and U13874 (N_13874,N_13701,N_13704);
nor U13875 (N_13875,N_13628,N_13797);
nand U13876 (N_13876,N_13794,N_13648);
nor U13877 (N_13877,N_13696,N_13600);
nor U13878 (N_13878,N_13789,N_13777);
and U13879 (N_13879,N_13743,N_13773);
or U13880 (N_13880,N_13640,N_13678);
and U13881 (N_13881,N_13727,N_13622);
and U13882 (N_13882,N_13799,N_13735);
xor U13883 (N_13883,N_13754,N_13763);
nor U13884 (N_13884,N_13665,N_13654);
or U13885 (N_13885,N_13667,N_13707);
xnor U13886 (N_13886,N_13652,N_13677);
nand U13887 (N_13887,N_13700,N_13649);
or U13888 (N_13888,N_13771,N_13716);
nor U13889 (N_13889,N_13792,N_13611);
and U13890 (N_13890,N_13766,N_13646);
and U13891 (N_13891,N_13641,N_13725);
nand U13892 (N_13892,N_13781,N_13744);
and U13893 (N_13893,N_13609,N_13653);
nand U13894 (N_13894,N_13615,N_13759);
or U13895 (N_13895,N_13731,N_13663);
nand U13896 (N_13896,N_13674,N_13795);
or U13897 (N_13897,N_13682,N_13602);
and U13898 (N_13898,N_13751,N_13691);
nor U13899 (N_13899,N_13706,N_13745);
nor U13900 (N_13900,N_13609,N_13648);
nand U13901 (N_13901,N_13674,N_13733);
xnor U13902 (N_13902,N_13731,N_13704);
nand U13903 (N_13903,N_13618,N_13633);
nand U13904 (N_13904,N_13748,N_13614);
nor U13905 (N_13905,N_13663,N_13622);
or U13906 (N_13906,N_13799,N_13710);
and U13907 (N_13907,N_13750,N_13672);
and U13908 (N_13908,N_13736,N_13671);
xor U13909 (N_13909,N_13667,N_13729);
or U13910 (N_13910,N_13693,N_13696);
nor U13911 (N_13911,N_13649,N_13617);
xnor U13912 (N_13912,N_13681,N_13637);
or U13913 (N_13913,N_13792,N_13625);
xor U13914 (N_13914,N_13767,N_13633);
nor U13915 (N_13915,N_13727,N_13680);
nor U13916 (N_13916,N_13794,N_13738);
or U13917 (N_13917,N_13692,N_13646);
nor U13918 (N_13918,N_13697,N_13793);
nand U13919 (N_13919,N_13752,N_13656);
nor U13920 (N_13920,N_13733,N_13799);
xor U13921 (N_13921,N_13657,N_13663);
and U13922 (N_13922,N_13769,N_13798);
nand U13923 (N_13923,N_13775,N_13653);
or U13924 (N_13924,N_13668,N_13778);
or U13925 (N_13925,N_13789,N_13669);
or U13926 (N_13926,N_13763,N_13784);
nor U13927 (N_13927,N_13656,N_13692);
nand U13928 (N_13928,N_13663,N_13613);
nand U13929 (N_13929,N_13692,N_13681);
nor U13930 (N_13930,N_13750,N_13617);
xnor U13931 (N_13931,N_13612,N_13716);
nor U13932 (N_13932,N_13752,N_13793);
nor U13933 (N_13933,N_13616,N_13692);
nor U13934 (N_13934,N_13793,N_13644);
and U13935 (N_13935,N_13728,N_13767);
nand U13936 (N_13936,N_13711,N_13749);
and U13937 (N_13937,N_13673,N_13677);
and U13938 (N_13938,N_13785,N_13715);
and U13939 (N_13939,N_13670,N_13677);
nand U13940 (N_13940,N_13760,N_13660);
nor U13941 (N_13941,N_13695,N_13776);
or U13942 (N_13942,N_13703,N_13750);
or U13943 (N_13943,N_13686,N_13791);
and U13944 (N_13944,N_13744,N_13668);
and U13945 (N_13945,N_13660,N_13736);
and U13946 (N_13946,N_13689,N_13734);
and U13947 (N_13947,N_13769,N_13638);
nand U13948 (N_13948,N_13639,N_13729);
or U13949 (N_13949,N_13658,N_13666);
nand U13950 (N_13950,N_13654,N_13725);
nand U13951 (N_13951,N_13602,N_13794);
nand U13952 (N_13952,N_13649,N_13659);
nor U13953 (N_13953,N_13718,N_13765);
xor U13954 (N_13954,N_13669,N_13700);
or U13955 (N_13955,N_13670,N_13785);
xnor U13956 (N_13956,N_13738,N_13694);
nand U13957 (N_13957,N_13648,N_13697);
and U13958 (N_13958,N_13701,N_13728);
nor U13959 (N_13959,N_13757,N_13650);
or U13960 (N_13960,N_13658,N_13745);
nor U13961 (N_13961,N_13685,N_13670);
nor U13962 (N_13962,N_13643,N_13760);
or U13963 (N_13963,N_13704,N_13792);
and U13964 (N_13964,N_13648,N_13693);
nor U13965 (N_13965,N_13768,N_13737);
or U13966 (N_13966,N_13623,N_13781);
xor U13967 (N_13967,N_13705,N_13686);
nand U13968 (N_13968,N_13740,N_13687);
nand U13969 (N_13969,N_13650,N_13624);
nor U13970 (N_13970,N_13640,N_13794);
or U13971 (N_13971,N_13780,N_13642);
nand U13972 (N_13972,N_13639,N_13630);
nor U13973 (N_13973,N_13640,N_13612);
nor U13974 (N_13974,N_13687,N_13714);
or U13975 (N_13975,N_13677,N_13623);
nand U13976 (N_13976,N_13783,N_13715);
or U13977 (N_13977,N_13798,N_13654);
xor U13978 (N_13978,N_13741,N_13699);
and U13979 (N_13979,N_13642,N_13649);
nor U13980 (N_13980,N_13750,N_13734);
nand U13981 (N_13981,N_13662,N_13740);
or U13982 (N_13982,N_13629,N_13652);
nand U13983 (N_13983,N_13739,N_13606);
nor U13984 (N_13984,N_13798,N_13699);
or U13985 (N_13985,N_13684,N_13608);
xnor U13986 (N_13986,N_13678,N_13777);
xor U13987 (N_13987,N_13766,N_13749);
or U13988 (N_13988,N_13647,N_13658);
nand U13989 (N_13989,N_13637,N_13653);
or U13990 (N_13990,N_13651,N_13739);
nor U13991 (N_13991,N_13682,N_13697);
nor U13992 (N_13992,N_13683,N_13781);
and U13993 (N_13993,N_13741,N_13626);
nand U13994 (N_13994,N_13683,N_13607);
and U13995 (N_13995,N_13784,N_13661);
or U13996 (N_13996,N_13652,N_13683);
and U13997 (N_13997,N_13728,N_13764);
and U13998 (N_13998,N_13709,N_13601);
nand U13999 (N_13999,N_13701,N_13621);
and U14000 (N_14000,N_13804,N_13811);
xor U14001 (N_14001,N_13845,N_13813);
nand U14002 (N_14002,N_13984,N_13989);
xnor U14003 (N_14003,N_13809,N_13821);
nand U14004 (N_14004,N_13935,N_13826);
and U14005 (N_14005,N_13893,N_13927);
xor U14006 (N_14006,N_13978,N_13922);
nor U14007 (N_14007,N_13894,N_13833);
xnor U14008 (N_14008,N_13936,N_13946);
and U14009 (N_14009,N_13921,N_13866);
nor U14010 (N_14010,N_13883,N_13876);
or U14011 (N_14011,N_13930,N_13871);
xnor U14012 (N_14012,N_13825,N_13998);
xnor U14013 (N_14013,N_13942,N_13881);
and U14014 (N_14014,N_13865,N_13939);
or U14015 (N_14015,N_13891,N_13975);
nand U14016 (N_14016,N_13806,N_13872);
and U14017 (N_14017,N_13933,N_13976);
nand U14018 (N_14018,N_13832,N_13870);
and U14019 (N_14019,N_13977,N_13948);
or U14020 (N_14020,N_13869,N_13915);
xor U14021 (N_14021,N_13817,N_13836);
or U14022 (N_14022,N_13960,N_13850);
xnor U14023 (N_14023,N_13898,N_13892);
nor U14024 (N_14024,N_13993,N_13816);
and U14025 (N_14025,N_13996,N_13991);
nand U14026 (N_14026,N_13916,N_13980);
or U14027 (N_14027,N_13957,N_13937);
xnor U14028 (N_14028,N_13967,N_13958);
nand U14029 (N_14029,N_13838,N_13801);
or U14030 (N_14030,N_13952,N_13940);
nor U14031 (N_14031,N_13995,N_13943);
xor U14032 (N_14032,N_13928,N_13912);
xor U14033 (N_14033,N_13822,N_13887);
nand U14034 (N_14034,N_13819,N_13824);
xnor U14035 (N_14035,N_13878,N_13924);
nor U14036 (N_14036,N_13886,N_13964);
and U14037 (N_14037,N_13963,N_13875);
or U14038 (N_14038,N_13884,N_13910);
nor U14039 (N_14039,N_13835,N_13810);
and U14040 (N_14040,N_13854,N_13805);
or U14041 (N_14041,N_13938,N_13808);
nor U14042 (N_14042,N_13955,N_13862);
or U14043 (N_14043,N_13888,N_13920);
or U14044 (N_14044,N_13983,N_13800);
xnor U14045 (N_14045,N_13839,N_13844);
nor U14046 (N_14046,N_13842,N_13944);
and U14047 (N_14047,N_13970,N_13831);
or U14048 (N_14048,N_13987,N_13851);
xnor U14049 (N_14049,N_13953,N_13981);
nand U14050 (N_14050,N_13904,N_13969);
and U14051 (N_14051,N_13945,N_13867);
and U14052 (N_14052,N_13907,N_13968);
and U14053 (N_14053,N_13855,N_13807);
nor U14054 (N_14054,N_13814,N_13973);
xnor U14055 (N_14055,N_13949,N_13997);
xnor U14056 (N_14056,N_13934,N_13914);
nor U14057 (N_14057,N_13919,N_13961);
xor U14058 (N_14058,N_13902,N_13897);
nand U14059 (N_14059,N_13923,N_13925);
and U14060 (N_14060,N_13812,N_13896);
or U14061 (N_14061,N_13909,N_13846);
nand U14062 (N_14062,N_13905,N_13827);
nand U14063 (N_14063,N_13834,N_13829);
xor U14064 (N_14064,N_13972,N_13947);
or U14065 (N_14065,N_13874,N_13841);
nor U14066 (N_14066,N_13848,N_13861);
or U14067 (N_14067,N_13956,N_13863);
or U14068 (N_14068,N_13950,N_13885);
or U14069 (N_14069,N_13830,N_13959);
and U14070 (N_14070,N_13818,N_13820);
or U14071 (N_14071,N_13908,N_13889);
nand U14072 (N_14072,N_13988,N_13873);
nand U14073 (N_14073,N_13917,N_13954);
nor U14074 (N_14074,N_13994,N_13900);
or U14075 (N_14075,N_13906,N_13895);
xnor U14076 (N_14076,N_13926,N_13890);
or U14077 (N_14077,N_13974,N_13966);
nor U14078 (N_14078,N_13932,N_13856);
nor U14079 (N_14079,N_13860,N_13931);
xnor U14080 (N_14080,N_13837,N_13858);
and U14081 (N_14081,N_13868,N_13979);
xnor U14082 (N_14082,N_13985,N_13843);
or U14083 (N_14083,N_13999,N_13929);
nand U14084 (N_14084,N_13913,N_13859);
nor U14085 (N_14085,N_13986,N_13951);
nand U14086 (N_14086,N_13941,N_13962);
nor U14087 (N_14087,N_13982,N_13853);
xor U14088 (N_14088,N_13992,N_13823);
and U14089 (N_14089,N_13857,N_13899);
nor U14090 (N_14090,N_13971,N_13879);
and U14091 (N_14091,N_13802,N_13864);
or U14092 (N_14092,N_13903,N_13911);
nand U14093 (N_14093,N_13852,N_13901);
xnor U14094 (N_14094,N_13918,N_13815);
xor U14095 (N_14095,N_13849,N_13965);
xnor U14096 (N_14096,N_13803,N_13990);
xor U14097 (N_14097,N_13877,N_13847);
nor U14098 (N_14098,N_13840,N_13828);
nand U14099 (N_14099,N_13882,N_13880);
xnor U14100 (N_14100,N_13822,N_13829);
xor U14101 (N_14101,N_13864,N_13828);
or U14102 (N_14102,N_13919,N_13921);
or U14103 (N_14103,N_13824,N_13884);
and U14104 (N_14104,N_13914,N_13907);
nor U14105 (N_14105,N_13889,N_13818);
xor U14106 (N_14106,N_13859,N_13826);
xnor U14107 (N_14107,N_13863,N_13925);
and U14108 (N_14108,N_13846,N_13848);
xor U14109 (N_14109,N_13836,N_13806);
nand U14110 (N_14110,N_13832,N_13966);
or U14111 (N_14111,N_13998,N_13951);
or U14112 (N_14112,N_13992,N_13962);
xor U14113 (N_14113,N_13888,N_13968);
nor U14114 (N_14114,N_13975,N_13896);
and U14115 (N_14115,N_13999,N_13823);
nor U14116 (N_14116,N_13989,N_13883);
nor U14117 (N_14117,N_13868,N_13917);
or U14118 (N_14118,N_13853,N_13944);
or U14119 (N_14119,N_13885,N_13927);
nor U14120 (N_14120,N_13887,N_13936);
or U14121 (N_14121,N_13881,N_13940);
or U14122 (N_14122,N_13907,N_13898);
nor U14123 (N_14123,N_13962,N_13843);
nand U14124 (N_14124,N_13860,N_13911);
and U14125 (N_14125,N_13991,N_13816);
nor U14126 (N_14126,N_13879,N_13984);
nor U14127 (N_14127,N_13937,N_13908);
xnor U14128 (N_14128,N_13815,N_13939);
xnor U14129 (N_14129,N_13875,N_13962);
xnor U14130 (N_14130,N_13931,N_13897);
nand U14131 (N_14131,N_13834,N_13933);
xnor U14132 (N_14132,N_13940,N_13814);
nand U14133 (N_14133,N_13904,N_13991);
nor U14134 (N_14134,N_13909,N_13809);
or U14135 (N_14135,N_13863,N_13813);
xor U14136 (N_14136,N_13920,N_13956);
nand U14137 (N_14137,N_13864,N_13880);
and U14138 (N_14138,N_13929,N_13934);
or U14139 (N_14139,N_13928,N_13925);
nor U14140 (N_14140,N_13941,N_13873);
nor U14141 (N_14141,N_13986,N_13892);
and U14142 (N_14142,N_13944,N_13880);
nor U14143 (N_14143,N_13855,N_13918);
and U14144 (N_14144,N_13846,N_13815);
nor U14145 (N_14145,N_13893,N_13842);
nor U14146 (N_14146,N_13949,N_13980);
or U14147 (N_14147,N_13849,N_13950);
xnor U14148 (N_14148,N_13829,N_13855);
nand U14149 (N_14149,N_13991,N_13841);
and U14150 (N_14150,N_13878,N_13905);
xnor U14151 (N_14151,N_13830,N_13851);
nor U14152 (N_14152,N_13954,N_13823);
and U14153 (N_14153,N_13831,N_13984);
xnor U14154 (N_14154,N_13937,N_13817);
nor U14155 (N_14155,N_13875,N_13948);
and U14156 (N_14156,N_13876,N_13961);
and U14157 (N_14157,N_13878,N_13940);
xnor U14158 (N_14158,N_13941,N_13929);
nor U14159 (N_14159,N_13859,N_13804);
nand U14160 (N_14160,N_13808,N_13926);
nand U14161 (N_14161,N_13825,N_13920);
nor U14162 (N_14162,N_13921,N_13864);
nor U14163 (N_14163,N_13951,N_13895);
and U14164 (N_14164,N_13934,N_13963);
or U14165 (N_14165,N_13901,N_13892);
nor U14166 (N_14166,N_13973,N_13835);
xor U14167 (N_14167,N_13857,N_13982);
or U14168 (N_14168,N_13856,N_13838);
and U14169 (N_14169,N_13838,N_13873);
nand U14170 (N_14170,N_13871,N_13845);
and U14171 (N_14171,N_13859,N_13839);
nor U14172 (N_14172,N_13802,N_13927);
nand U14173 (N_14173,N_13939,N_13901);
nand U14174 (N_14174,N_13818,N_13968);
or U14175 (N_14175,N_13918,N_13898);
nand U14176 (N_14176,N_13828,N_13983);
or U14177 (N_14177,N_13880,N_13907);
xor U14178 (N_14178,N_13962,N_13809);
or U14179 (N_14179,N_13929,N_13914);
xor U14180 (N_14180,N_13964,N_13830);
nand U14181 (N_14181,N_13877,N_13875);
and U14182 (N_14182,N_13892,N_13899);
or U14183 (N_14183,N_13921,N_13922);
or U14184 (N_14184,N_13922,N_13939);
nand U14185 (N_14185,N_13889,N_13836);
nor U14186 (N_14186,N_13940,N_13829);
nor U14187 (N_14187,N_13852,N_13913);
nand U14188 (N_14188,N_13885,N_13996);
or U14189 (N_14189,N_13984,N_13890);
xor U14190 (N_14190,N_13924,N_13898);
xor U14191 (N_14191,N_13947,N_13905);
and U14192 (N_14192,N_13938,N_13909);
and U14193 (N_14193,N_13869,N_13969);
nand U14194 (N_14194,N_13960,N_13963);
nor U14195 (N_14195,N_13905,N_13879);
and U14196 (N_14196,N_13958,N_13861);
xor U14197 (N_14197,N_13868,N_13815);
and U14198 (N_14198,N_13852,N_13986);
and U14199 (N_14199,N_13857,N_13881);
nor U14200 (N_14200,N_14059,N_14052);
or U14201 (N_14201,N_14038,N_14057);
and U14202 (N_14202,N_14169,N_14143);
nor U14203 (N_14203,N_14097,N_14082);
and U14204 (N_14204,N_14094,N_14083);
xor U14205 (N_14205,N_14120,N_14100);
or U14206 (N_14206,N_14027,N_14118);
and U14207 (N_14207,N_14049,N_14075);
and U14208 (N_14208,N_14163,N_14146);
or U14209 (N_14209,N_14117,N_14104);
or U14210 (N_14210,N_14155,N_14149);
and U14211 (N_14211,N_14159,N_14178);
nor U14212 (N_14212,N_14054,N_14095);
and U14213 (N_14213,N_14076,N_14172);
xnor U14214 (N_14214,N_14193,N_14047);
nor U14215 (N_14215,N_14115,N_14081);
nor U14216 (N_14216,N_14026,N_14074);
and U14217 (N_14217,N_14157,N_14086);
nor U14218 (N_14218,N_14060,N_14152);
nand U14219 (N_14219,N_14138,N_14062);
nand U14220 (N_14220,N_14108,N_14024);
xnor U14221 (N_14221,N_14184,N_14069);
nand U14222 (N_14222,N_14106,N_14014);
nor U14223 (N_14223,N_14170,N_14037);
nand U14224 (N_14224,N_14020,N_14031);
and U14225 (N_14225,N_14071,N_14063);
nand U14226 (N_14226,N_14122,N_14085);
nand U14227 (N_14227,N_14187,N_14003);
and U14228 (N_14228,N_14176,N_14045);
and U14229 (N_14229,N_14034,N_14180);
xor U14230 (N_14230,N_14015,N_14011);
xnor U14231 (N_14231,N_14191,N_14182);
nand U14232 (N_14232,N_14194,N_14098);
nand U14233 (N_14233,N_14046,N_14010);
nand U14234 (N_14234,N_14165,N_14017);
xor U14235 (N_14235,N_14002,N_14039);
nor U14236 (N_14236,N_14116,N_14036);
or U14237 (N_14237,N_14087,N_14160);
or U14238 (N_14238,N_14012,N_14001);
nand U14239 (N_14239,N_14177,N_14158);
nand U14240 (N_14240,N_14032,N_14053);
xor U14241 (N_14241,N_14064,N_14025);
nor U14242 (N_14242,N_14009,N_14192);
nand U14243 (N_14243,N_14199,N_14088);
or U14244 (N_14244,N_14140,N_14171);
or U14245 (N_14245,N_14105,N_14096);
or U14246 (N_14246,N_14173,N_14154);
or U14247 (N_14247,N_14078,N_14103);
or U14248 (N_14248,N_14127,N_14050);
nor U14249 (N_14249,N_14123,N_14041);
or U14250 (N_14250,N_14005,N_14040);
xnor U14251 (N_14251,N_14091,N_14109);
nor U14252 (N_14252,N_14153,N_14055);
and U14253 (N_14253,N_14196,N_14197);
xor U14254 (N_14254,N_14029,N_14084);
nand U14255 (N_14255,N_14164,N_14042);
nor U14256 (N_14256,N_14121,N_14189);
nand U14257 (N_14257,N_14133,N_14072);
nand U14258 (N_14258,N_14181,N_14114);
or U14259 (N_14259,N_14007,N_14134);
xnor U14260 (N_14260,N_14058,N_14043);
xnor U14261 (N_14261,N_14019,N_14061);
nor U14262 (N_14262,N_14119,N_14021);
or U14263 (N_14263,N_14156,N_14148);
nor U14264 (N_14264,N_14186,N_14000);
nor U14265 (N_14265,N_14090,N_14022);
or U14266 (N_14266,N_14068,N_14185);
or U14267 (N_14267,N_14179,N_14142);
nand U14268 (N_14268,N_14136,N_14093);
nand U14269 (N_14269,N_14150,N_14006);
nor U14270 (N_14270,N_14145,N_14188);
nand U14271 (N_14271,N_14137,N_14077);
or U14272 (N_14272,N_14129,N_14139);
nor U14273 (N_14273,N_14018,N_14013);
or U14274 (N_14274,N_14124,N_14089);
or U14275 (N_14275,N_14079,N_14195);
xor U14276 (N_14276,N_14099,N_14125);
or U14277 (N_14277,N_14112,N_14080);
nand U14278 (N_14278,N_14144,N_14147);
and U14279 (N_14279,N_14110,N_14131);
and U14280 (N_14280,N_14198,N_14048);
nor U14281 (N_14281,N_14033,N_14126);
nor U14282 (N_14282,N_14128,N_14151);
nor U14283 (N_14283,N_14130,N_14035);
xnor U14284 (N_14284,N_14183,N_14190);
nand U14285 (N_14285,N_14141,N_14073);
xor U14286 (N_14286,N_14016,N_14113);
xor U14287 (N_14287,N_14162,N_14067);
nor U14288 (N_14288,N_14030,N_14161);
nor U14289 (N_14289,N_14167,N_14111);
xor U14290 (N_14290,N_14102,N_14092);
or U14291 (N_14291,N_14066,N_14023);
or U14292 (N_14292,N_14008,N_14070);
and U14293 (N_14293,N_14065,N_14028);
xnor U14294 (N_14294,N_14101,N_14051);
or U14295 (N_14295,N_14107,N_14175);
or U14296 (N_14296,N_14056,N_14174);
xnor U14297 (N_14297,N_14004,N_14132);
xnor U14298 (N_14298,N_14166,N_14044);
nor U14299 (N_14299,N_14135,N_14168);
xor U14300 (N_14300,N_14169,N_14125);
and U14301 (N_14301,N_14088,N_14189);
or U14302 (N_14302,N_14059,N_14117);
or U14303 (N_14303,N_14102,N_14096);
xnor U14304 (N_14304,N_14176,N_14091);
or U14305 (N_14305,N_14037,N_14047);
xor U14306 (N_14306,N_14154,N_14007);
nand U14307 (N_14307,N_14067,N_14086);
nor U14308 (N_14308,N_14123,N_14091);
nor U14309 (N_14309,N_14117,N_14163);
nor U14310 (N_14310,N_14020,N_14187);
nor U14311 (N_14311,N_14011,N_14040);
or U14312 (N_14312,N_14175,N_14111);
and U14313 (N_14313,N_14175,N_14072);
nor U14314 (N_14314,N_14158,N_14086);
xor U14315 (N_14315,N_14066,N_14024);
nor U14316 (N_14316,N_14017,N_14109);
nand U14317 (N_14317,N_14186,N_14176);
and U14318 (N_14318,N_14188,N_14018);
and U14319 (N_14319,N_14011,N_14144);
and U14320 (N_14320,N_14174,N_14189);
and U14321 (N_14321,N_14075,N_14127);
or U14322 (N_14322,N_14088,N_14159);
nand U14323 (N_14323,N_14010,N_14061);
or U14324 (N_14324,N_14161,N_14046);
or U14325 (N_14325,N_14096,N_14160);
nor U14326 (N_14326,N_14014,N_14113);
and U14327 (N_14327,N_14184,N_14162);
xnor U14328 (N_14328,N_14016,N_14042);
nor U14329 (N_14329,N_14048,N_14143);
xor U14330 (N_14330,N_14150,N_14079);
nand U14331 (N_14331,N_14120,N_14187);
xnor U14332 (N_14332,N_14108,N_14113);
and U14333 (N_14333,N_14152,N_14002);
xnor U14334 (N_14334,N_14177,N_14075);
xor U14335 (N_14335,N_14071,N_14061);
nor U14336 (N_14336,N_14077,N_14088);
nor U14337 (N_14337,N_14009,N_14010);
nand U14338 (N_14338,N_14143,N_14073);
nor U14339 (N_14339,N_14075,N_14176);
and U14340 (N_14340,N_14003,N_14162);
nand U14341 (N_14341,N_14030,N_14010);
nand U14342 (N_14342,N_14043,N_14021);
nor U14343 (N_14343,N_14199,N_14084);
or U14344 (N_14344,N_14160,N_14114);
nor U14345 (N_14345,N_14180,N_14117);
nand U14346 (N_14346,N_14194,N_14141);
and U14347 (N_14347,N_14155,N_14046);
xnor U14348 (N_14348,N_14148,N_14093);
xor U14349 (N_14349,N_14040,N_14103);
xnor U14350 (N_14350,N_14129,N_14126);
nor U14351 (N_14351,N_14135,N_14162);
or U14352 (N_14352,N_14041,N_14081);
xnor U14353 (N_14353,N_14140,N_14036);
or U14354 (N_14354,N_14061,N_14013);
or U14355 (N_14355,N_14190,N_14159);
xnor U14356 (N_14356,N_14102,N_14173);
nor U14357 (N_14357,N_14059,N_14068);
nor U14358 (N_14358,N_14029,N_14021);
and U14359 (N_14359,N_14128,N_14087);
nor U14360 (N_14360,N_14011,N_14089);
nand U14361 (N_14361,N_14092,N_14139);
nor U14362 (N_14362,N_14146,N_14077);
or U14363 (N_14363,N_14027,N_14140);
nor U14364 (N_14364,N_14031,N_14156);
or U14365 (N_14365,N_14168,N_14093);
and U14366 (N_14366,N_14183,N_14122);
and U14367 (N_14367,N_14048,N_14101);
nor U14368 (N_14368,N_14119,N_14032);
nand U14369 (N_14369,N_14179,N_14154);
nor U14370 (N_14370,N_14023,N_14144);
and U14371 (N_14371,N_14160,N_14162);
nor U14372 (N_14372,N_14102,N_14003);
xnor U14373 (N_14373,N_14069,N_14185);
or U14374 (N_14374,N_14035,N_14142);
nor U14375 (N_14375,N_14098,N_14177);
xnor U14376 (N_14376,N_14039,N_14107);
and U14377 (N_14377,N_14062,N_14061);
or U14378 (N_14378,N_14053,N_14064);
xor U14379 (N_14379,N_14056,N_14013);
and U14380 (N_14380,N_14008,N_14099);
or U14381 (N_14381,N_14141,N_14027);
nand U14382 (N_14382,N_14018,N_14034);
or U14383 (N_14383,N_14131,N_14022);
xnor U14384 (N_14384,N_14039,N_14083);
xnor U14385 (N_14385,N_14172,N_14019);
or U14386 (N_14386,N_14169,N_14082);
and U14387 (N_14387,N_14138,N_14162);
xnor U14388 (N_14388,N_14077,N_14157);
nor U14389 (N_14389,N_14196,N_14139);
nor U14390 (N_14390,N_14041,N_14090);
nand U14391 (N_14391,N_14198,N_14100);
and U14392 (N_14392,N_14183,N_14166);
xnor U14393 (N_14393,N_14095,N_14069);
xor U14394 (N_14394,N_14165,N_14152);
nand U14395 (N_14395,N_14012,N_14016);
and U14396 (N_14396,N_14084,N_14003);
or U14397 (N_14397,N_14079,N_14038);
xnor U14398 (N_14398,N_14070,N_14051);
and U14399 (N_14399,N_14163,N_14134);
nand U14400 (N_14400,N_14396,N_14209);
and U14401 (N_14401,N_14245,N_14366);
nor U14402 (N_14402,N_14358,N_14363);
nand U14403 (N_14403,N_14397,N_14316);
nand U14404 (N_14404,N_14342,N_14341);
nor U14405 (N_14405,N_14332,N_14235);
xnor U14406 (N_14406,N_14354,N_14222);
xnor U14407 (N_14407,N_14214,N_14251);
xnor U14408 (N_14408,N_14355,N_14319);
xnor U14409 (N_14409,N_14345,N_14310);
xnor U14410 (N_14410,N_14280,N_14391);
and U14411 (N_14411,N_14320,N_14290);
and U14412 (N_14412,N_14385,N_14333);
xor U14413 (N_14413,N_14348,N_14381);
or U14414 (N_14414,N_14337,N_14211);
nand U14415 (N_14415,N_14263,N_14240);
nor U14416 (N_14416,N_14379,N_14206);
or U14417 (N_14417,N_14253,N_14228);
nor U14418 (N_14418,N_14302,N_14250);
nor U14419 (N_14419,N_14344,N_14288);
nand U14420 (N_14420,N_14356,N_14324);
xor U14421 (N_14421,N_14289,N_14393);
or U14422 (N_14422,N_14306,N_14234);
xnor U14423 (N_14423,N_14231,N_14340);
or U14424 (N_14424,N_14359,N_14338);
nand U14425 (N_14425,N_14361,N_14293);
nor U14426 (N_14426,N_14285,N_14339);
nand U14427 (N_14427,N_14230,N_14266);
nor U14428 (N_14428,N_14217,N_14346);
xnor U14429 (N_14429,N_14352,N_14399);
nand U14430 (N_14430,N_14225,N_14314);
nand U14431 (N_14431,N_14331,N_14264);
nand U14432 (N_14432,N_14223,N_14369);
nor U14433 (N_14433,N_14201,N_14281);
and U14434 (N_14434,N_14274,N_14334);
nor U14435 (N_14435,N_14260,N_14203);
nor U14436 (N_14436,N_14227,N_14249);
xor U14437 (N_14437,N_14258,N_14270);
nor U14438 (N_14438,N_14311,N_14398);
or U14439 (N_14439,N_14376,N_14325);
nor U14440 (N_14440,N_14278,N_14374);
nand U14441 (N_14441,N_14248,N_14275);
nand U14442 (N_14442,N_14343,N_14202);
and U14443 (N_14443,N_14387,N_14257);
or U14444 (N_14444,N_14277,N_14262);
xor U14445 (N_14445,N_14205,N_14254);
nor U14446 (N_14446,N_14208,N_14216);
and U14447 (N_14447,N_14283,N_14318);
xor U14448 (N_14448,N_14232,N_14242);
xnor U14449 (N_14449,N_14207,N_14347);
nand U14450 (N_14450,N_14243,N_14323);
nor U14451 (N_14451,N_14291,N_14353);
nand U14452 (N_14452,N_14238,N_14237);
nand U14453 (N_14453,N_14226,N_14351);
nand U14454 (N_14454,N_14279,N_14365);
nand U14455 (N_14455,N_14256,N_14236);
nand U14456 (N_14456,N_14317,N_14269);
or U14457 (N_14457,N_14218,N_14375);
xnor U14458 (N_14458,N_14330,N_14372);
or U14459 (N_14459,N_14305,N_14350);
nand U14460 (N_14460,N_14259,N_14377);
and U14461 (N_14461,N_14296,N_14247);
and U14462 (N_14462,N_14267,N_14367);
and U14463 (N_14463,N_14284,N_14255);
xor U14464 (N_14464,N_14307,N_14384);
xnor U14465 (N_14465,N_14360,N_14294);
nand U14466 (N_14466,N_14215,N_14252);
xnor U14467 (N_14467,N_14378,N_14392);
nor U14468 (N_14468,N_14357,N_14271);
xnor U14469 (N_14469,N_14389,N_14390);
or U14470 (N_14470,N_14301,N_14370);
nand U14471 (N_14471,N_14241,N_14335);
and U14472 (N_14472,N_14308,N_14239);
nand U14473 (N_14473,N_14304,N_14246);
xor U14474 (N_14474,N_14297,N_14329);
nand U14475 (N_14475,N_14282,N_14336);
and U14476 (N_14476,N_14265,N_14313);
and U14477 (N_14477,N_14220,N_14287);
and U14478 (N_14478,N_14382,N_14261);
xnor U14479 (N_14479,N_14292,N_14364);
nand U14480 (N_14480,N_14273,N_14272);
nand U14481 (N_14481,N_14373,N_14315);
xor U14482 (N_14482,N_14349,N_14327);
nand U14483 (N_14483,N_14326,N_14200);
nand U14484 (N_14484,N_14212,N_14312);
nand U14485 (N_14485,N_14204,N_14295);
xnor U14486 (N_14486,N_14268,N_14371);
nor U14487 (N_14487,N_14322,N_14210);
xnor U14488 (N_14488,N_14276,N_14383);
or U14489 (N_14489,N_14286,N_14368);
nand U14490 (N_14490,N_14386,N_14244);
and U14491 (N_14491,N_14299,N_14362);
xnor U14492 (N_14492,N_14395,N_14303);
and U14493 (N_14493,N_14328,N_14388);
or U14494 (N_14494,N_14224,N_14213);
nor U14495 (N_14495,N_14219,N_14380);
nor U14496 (N_14496,N_14221,N_14394);
nor U14497 (N_14497,N_14321,N_14309);
xnor U14498 (N_14498,N_14229,N_14298);
xor U14499 (N_14499,N_14300,N_14233);
nand U14500 (N_14500,N_14380,N_14391);
and U14501 (N_14501,N_14398,N_14268);
nand U14502 (N_14502,N_14354,N_14260);
xnor U14503 (N_14503,N_14307,N_14300);
xnor U14504 (N_14504,N_14392,N_14330);
or U14505 (N_14505,N_14373,N_14276);
xor U14506 (N_14506,N_14374,N_14383);
nand U14507 (N_14507,N_14271,N_14211);
and U14508 (N_14508,N_14350,N_14204);
or U14509 (N_14509,N_14336,N_14270);
xor U14510 (N_14510,N_14355,N_14363);
or U14511 (N_14511,N_14323,N_14215);
xor U14512 (N_14512,N_14397,N_14201);
and U14513 (N_14513,N_14359,N_14208);
nand U14514 (N_14514,N_14397,N_14375);
or U14515 (N_14515,N_14281,N_14325);
or U14516 (N_14516,N_14228,N_14268);
and U14517 (N_14517,N_14349,N_14315);
and U14518 (N_14518,N_14396,N_14264);
xor U14519 (N_14519,N_14305,N_14394);
nand U14520 (N_14520,N_14252,N_14209);
and U14521 (N_14521,N_14249,N_14216);
nand U14522 (N_14522,N_14229,N_14284);
or U14523 (N_14523,N_14344,N_14311);
or U14524 (N_14524,N_14249,N_14217);
nand U14525 (N_14525,N_14273,N_14367);
xnor U14526 (N_14526,N_14364,N_14242);
or U14527 (N_14527,N_14304,N_14243);
and U14528 (N_14528,N_14216,N_14399);
or U14529 (N_14529,N_14296,N_14218);
or U14530 (N_14530,N_14218,N_14297);
or U14531 (N_14531,N_14288,N_14267);
and U14532 (N_14532,N_14381,N_14389);
and U14533 (N_14533,N_14352,N_14365);
nand U14534 (N_14534,N_14352,N_14253);
nor U14535 (N_14535,N_14244,N_14397);
or U14536 (N_14536,N_14245,N_14289);
nor U14537 (N_14537,N_14302,N_14248);
nor U14538 (N_14538,N_14336,N_14214);
xor U14539 (N_14539,N_14329,N_14369);
nand U14540 (N_14540,N_14205,N_14238);
nor U14541 (N_14541,N_14356,N_14251);
nand U14542 (N_14542,N_14267,N_14250);
xor U14543 (N_14543,N_14201,N_14285);
xnor U14544 (N_14544,N_14266,N_14354);
nand U14545 (N_14545,N_14271,N_14301);
or U14546 (N_14546,N_14340,N_14354);
and U14547 (N_14547,N_14308,N_14389);
xnor U14548 (N_14548,N_14397,N_14222);
and U14549 (N_14549,N_14293,N_14385);
nand U14550 (N_14550,N_14291,N_14366);
nand U14551 (N_14551,N_14308,N_14285);
nand U14552 (N_14552,N_14361,N_14271);
and U14553 (N_14553,N_14370,N_14392);
nand U14554 (N_14554,N_14272,N_14260);
or U14555 (N_14555,N_14346,N_14367);
nor U14556 (N_14556,N_14239,N_14251);
xnor U14557 (N_14557,N_14370,N_14328);
xor U14558 (N_14558,N_14304,N_14213);
and U14559 (N_14559,N_14325,N_14354);
xnor U14560 (N_14560,N_14265,N_14332);
and U14561 (N_14561,N_14275,N_14386);
nand U14562 (N_14562,N_14313,N_14294);
nor U14563 (N_14563,N_14215,N_14376);
and U14564 (N_14564,N_14235,N_14257);
nand U14565 (N_14565,N_14245,N_14344);
or U14566 (N_14566,N_14214,N_14235);
xor U14567 (N_14567,N_14268,N_14341);
and U14568 (N_14568,N_14313,N_14268);
nor U14569 (N_14569,N_14349,N_14297);
xnor U14570 (N_14570,N_14333,N_14332);
nand U14571 (N_14571,N_14282,N_14250);
nor U14572 (N_14572,N_14276,N_14307);
nor U14573 (N_14573,N_14200,N_14346);
and U14574 (N_14574,N_14357,N_14277);
and U14575 (N_14575,N_14354,N_14295);
or U14576 (N_14576,N_14309,N_14386);
xor U14577 (N_14577,N_14227,N_14393);
and U14578 (N_14578,N_14246,N_14262);
and U14579 (N_14579,N_14221,N_14379);
or U14580 (N_14580,N_14353,N_14308);
nor U14581 (N_14581,N_14268,N_14349);
nand U14582 (N_14582,N_14231,N_14240);
nand U14583 (N_14583,N_14393,N_14330);
xnor U14584 (N_14584,N_14324,N_14352);
nor U14585 (N_14585,N_14276,N_14211);
or U14586 (N_14586,N_14288,N_14239);
xor U14587 (N_14587,N_14269,N_14202);
or U14588 (N_14588,N_14307,N_14210);
and U14589 (N_14589,N_14393,N_14364);
nand U14590 (N_14590,N_14375,N_14324);
or U14591 (N_14591,N_14277,N_14367);
xnor U14592 (N_14592,N_14390,N_14210);
or U14593 (N_14593,N_14211,N_14286);
nand U14594 (N_14594,N_14358,N_14369);
nand U14595 (N_14595,N_14241,N_14273);
xnor U14596 (N_14596,N_14335,N_14300);
and U14597 (N_14597,N_14278,N_14381);
xnor U14598 (N_14598,N_14302,N_14317);
xor U14599 (N_14599,N_14348,N_14344);
nor U14600 (N_14600,N_14596,N_14598);
and U14601 (N_14601,N_14520,N_14535);
or U14602 (N_14602,N_14486,N_14464);
and U14603 (N_14603,N_14558,N_14523);
xnor U14604 (N_14604,N_14524,N_14431);
xnor U14605 (N_14605,N_14414,N_14566);
nor U14606 (N_14606,N_14561,N_14421);
xor U14607 (N_14607,N_14449,N_14441);
nand U14608 (N_14608,N_14578,N_14501);
nor U14609 (N_14609,N_14545,N_14574);
xnor U14610 (N_14610,N_14497,N_14594);
and U14611 (N_14611,N_14567,N_14554);
or U14612 (N_14612,N_14490,N_14415);
and U14613 (N_14613,N_14476,N_14468);
nand U14614 (N_14614,N_14466,N_14427);
nand U14615 (N_14615,N_14469,N_14452);
or U14616 (N_14616,N_14515,N_14495);
or U14617 (N_14617,N_14511,N_14539);
nand U14618 (N_14618,N_14517,N_14573);
and U14619 (N_14619,N_14454,N_14478);
nand U14620 (N_14620,N_14577,N_14503);
nor U14621 (N_14621,N_14475,N_14496);
nand U14622 (N_14622,N_14420,N_14576);
or U14623 (N_14623,N_14417,N_14423);
and U14624 (N_14624,N_14440,N_14544);
or U14625 (N_14625,N_14550,N_14487);
xnor U14626 (N_14626,N_14547,N_14589);
nand U14627 (N_14627,N_14568,N_14500);
nor U14628 (N_14628,N_14473,N_14461);
or U14629 (N_14629,N_14489,N_14453);
and U14630 (N_14630,N_14467,N_14562);
or U14631 (N_14631,N_14530,N_14548);
nand U14632 (N_14632,N_14422,N_14525);
and U14633 (N_14633,N_14529,N_14590);
or U14634 (N_14634,N_14512,N_14409);
and U14635 (N_14635,N_14400,N_14563);
nand U14636 (N_14636,N_14460,N_14405);
or U14637 (N_14637,N_14436,N_14418);
nand U14638 (N_14638,N_14521,N_14446);
nand U14639 (N_14639,N_14408,N_14581);
nor U14640 (N_14640,N_14527,N_14508);
nor U14641 (N_14641,N_14555,N_14597);
or U14642 (N_14642,N_14488,N_14498);
nand U14643 (N_14643,N_14557,N_14481);
and U14644 (N_14644,N_14565,N_14599);
xor U14645 (N_14645,N_14439,N_14438);
and U14646 (N_14646,N_14458,N_14419);
or U14647 (N_14647,N_14401,N_14484);
xnor U14648 (N_14648,N_14447,N_14445);
or U14649 (N_14649,N_14571,N_14528);
xor U14650 (N_14650,N_14504,N_14428);
nor U14651 (N_14651,N_14472,N_14451);
and U14652 (N_14652,N_14410,N_14522);
nor U14653 (N_14653,N_14492,N_14549);
and U14654 (N_14654,N_14588,N_14494);
nand U14655 (N_14655,N_14437,N_14583);
and U14656 (N_14656,N_14536,N_14491);
nand U14657 (N_14657,N_14592,N_14404);
nor U14658 (N_14658,N_14514,N_14411);
or U14659 (N_14659,N_14552,N_14448);
or U14660 (N_14660,N_14587,N_14507);
nand U14661 (N_14661,N_14531,N_14493);
and U14662 (N_14662,N_14564,N_14506);
and U14663 (N_14663,N_14456,N_14406);
and U14664 (N_14664,N_14553,N_14559);
nand U14665 (N_14665,N_14537,N_14593);
nand U14666 (N_14666,N_14402,N_14569);
nand U14667 (N_14667,N_14502,N_14575);
and U14668 (N_14668,N_14435,N_14543);
nor U14669 (N_14669,N_14450,N_14570);
or U14670 (N_14670,N_14499,N_14533);
nor U14671 (N_14671,N_14579,N_14426);
and U14672 (N_14672,N_14534,N_14572);
xor U14673 (N_14673,N_14585,N_14485);
xnor U14674 (N_14674,N_14595,N_14425);
nand U14675 (N_14675,N_14471,N_14518);
or U14676 (N_14676,N_14546,N_14519);
nand U14677 (N_14677,N_14538,N_14470);
xor U14678 (N_14678,N_14424,N_14432);
or U14679 (N_14679,N_14413,N_14463);
nand U14680 (N_14680,N_14477,N_14580);
xor U14681 (N_14681,N_14444,N_14591);
nor U14682 (N_14682,N_14510,N_14443);
xor U14683 (N_14683,N_14532,N_14542);
nor U14684 (N_14684,N_14540,N_14513);
and U14685 (N_14685,N_14526,N_14433);
or U14686 (N_14686,N_14465,N_14584);
or U14687 (N_14687,N_14560,N_14462);
nand U14688 (N_14688,N_14457,N_14479);
and U14689 (N_14689,N_14480,N_14509);
or U14690 (N_14690,N_14556,N_14416);
or U14691 (N_14691,N_14483,N_14403);
and U14692 (N_14692,N_14442,N_14586);
nor U14693 (N_14693,N_14474,N_14429);
and U14694 (N_14694,N_14516,N_14430);
or U14695 (N_14695,N_14582,N_14551);
nand U14696 (N_14696,N_14412,N_14455);
nand U14697 (N_14697,N_14434,N_14541);
nor U14698 (N_14698,N_14407,N_14459);
nand U14699 (N_14699,N_14482,N_14505);
nor U14700 (N_14700,N_14597,N_14599);
nand U14701 (N_14701,N_14539,N_14558);
and U14702 (N_14702,N_14447,N_14512);
and U14703 (N_14703,N_14459,N_14470);
nor U14704 (N_14704,N_14432,N_14469);
nand U14705 (N_14705,N_14471,N_14492);
nand U14706 (N_14706,N_14492,N_14530);
xnor U14707 (N_14707,N_14423,N_14535);
xnor U14708 (N_14708,N_14451,N_14448);
nand U14709 (N_14709,N_14458,N_14546);
or U14710 (N_14710,N_14518,N_14414);
and U14711 (N_14711,N_14499,N_14443);
and U14712 (N_14712,N_14437,N_14545);
and U14713 (N_14713,N_14552,N_14517);
nor U14714 (N_14714,N_14516,N_14513);
and U14715 (N_14715,N_14478,N_14520);
xnor U14716 (N_14716,N_14457,N_14463);
xor U14717 (N_14717,N_14480,N_14526);
nand U14718 (N_14718,N_14519,N_14439);
xnor U14719 (N_14719,N_14586,N_14445);
or U14720 (N_14720,N_14451,N_14405);
or U14721 (N_14721,N_14585,N_14412);
nor U14722 (N_14722,N_14598,N_14510);
and U14723 (N_14723,N_14475,N_14556);
and U14724 (N_14724,N_14565,N_14463);
or U14725 (N_14725,N_14563,N_14463);
and U14726 (N_14726,N_14436,N_14515);
and U14727 (N_14727,N_14507,N_14469);
nand U14728 (N_14728,N_14483,N_14458);
xnor U14729 (N_14729,N_14442,N_14535);
nand U14730 (N_14730,N_14428,N_14442);
and U14731 (N_14731,N_14486,N_14536);
nor U14732 (N_14732,N_14437,N_14493);
or U14733 (N_14733,N_14518,N_14534);
nand U14734 (N_14734,N_14484,N_14567);
or U14735 (N_14735,N_14454,N_14452);
and U14736 (N_14736,N_14520,N_14554);
xor U14737 (N_14737,N_14489,N_14540);
nor U14738 (N_14738,N_14488,N_14452);
nor U14739 (N_14739,N_14463,N_14484);
and U14740 (N_14740,N_14412,N_14403);
nand U14741 (N_14741,N_14433,N_14413);
or U14742 (N_14742,N_14444,N_14518);
nand U14743 (N_14743,N_14597,N_14450);
or U14744 (N_14744,N_14485,N_14422);
xor U14745 (N_14745,N_14481,N_14594);
nor U14746 (N_14746,N_14482,N_14468);
and U14747 (N_14747,N_14420,N_14534);
xor U14748 (N_14748,N_14587,N_14479);
or U14749 (N_14749,N_14419,N_14450);
xnor U14750 (N_14750,N_14441,N_14523);
xnor U14751 (N_14751,N_14508,N_14526);
or U14752 (N_14752,N_14506,N_14535);
and U14753 (N_14753,N_14487,N_14463);
nor U14754 (N_14754,N_14548,N_14407);
and U14755 (N_14755,N_14462,N_14491);
or U14756 (N_14756,N_14584,N_14428);
xor U14757 (N_14757,N_14434,N_14406);
xor U14758 (N_14758,N_14453,N_14526);
and U14759 (N_14759,N_14591,N_14481);
and U14760 (N_14760,N_14440,N_14592);
nor U14761 (N_14761,N_14471,N_14419);
nor U14762 (N_14762,N_14464,N_14475);
nor U14763 (N_14763,N_14423,N_14593);
or U14764 (N_14764,N_14577,N_14521);
and U14765 (N_14765,N_14430,N_14407);
and U14766 (N_14766,N_14483,N_14423);
or U14767 (N_14767,N_14548,N_14522);
or U14768 (N_14768,N_14419,N_14404);
or U14769 (N_14769,N_14541,N_14485);
or U14770 (N_14770,N_14597,N_14440);
xnor U14771 (N_14771,N_14565,N_14551);
nand U14772 (N_14772,N_14530,N_14517);
and U14773 (N_14773,N_14465,N_14497);
and U14774 (N_14774,N_14544,N_14431);
xor U14775 (N_14775,N_14407,N_14528);
nand U14776 (N_14776,N_14559,N_14530);
xnor U14777 (N_14777,N_14443,N_14540);
nand U14778 (N_14778,N_14413,N_14477);
nor U14779 (N_14779,N_14469,N_14492);
nand U14780 (N_14780,N_14456,N_14577);
and U14781 (N_14781,N_14431,N_14429);
nand U14782 (N_14782,N_14566,N_14543);
nand U14783 (N_14783,N_14529,N_14573);
and U14784 (N_14784,N_14574,N_14479);
nand U14785 (N_14785,N_14565,N_14433);
nor U14786 (N_14786,N_14547,N_14509);
and U14787 (N_14787,N_14553,N_14479);
xor U14788 (N_14788,N_14587,N_14586);
or U14789 (N_14789,N_14540,N_14571);
xor U14790 (N_14790,N_14597,N_14549);
nand U14791 (N_14791,N_14423,N_14435);
and U14792 (N_14792,N_14458,N_14525);
xnor U14793 (N_14793,N_14558,N_14549);
nor U14794 (N_14794,N_14546,N_14451);
or U14795 (N_14795,N_14499,N_14429);
or U14796 (N_14796,N_14527,N_14580);
and U14797 (N_14797,N_14499,N_14446);
nor U14798 (N_14798,N_14504,N_14529);
nand U14799 (N_14799,N_14475,N_14469);
nor U14800 (N_14800,N_14664,N_14700);
nand U14801 (N_14801,N_14644,N_14675);
nor U14802 (N_14802,N_14659,N_14796);
nand U14803 (N_14803,N_14723,N_14647);
nor U14804 (N_14804,N_14688,N_14758);
nor U14805 (N_14805,N_14681,N_14703);
or U14806 (N_14806,N_14743,N_14634);
nor U14807 (N_14807,N_14661,N_14750);
nand U14808 (N_14808,N_14776,N_14683);
xnor U14809 (N_14809,N_14694,N_14605);
xnor U14810 (N_14810,N_14774,N_14756);
and U14811 (N_14811,N_14669,N_14779);
nand U14812 (N_14812,N_14639,N_14650);
and U14813 (N_14813,N_14754,N_14642);
and U14814 (N_14814,N_14620,N_14765);
nand U14815 (N_14815,N_14770,N_14737);
and U14816 (N_14816,N_14649,N_14612);
nand U14817 (N_14817,N_14792,N_14739);
nor U14818 (N_14818,N_14711,N_14720);
or U14819 (N_14819,N_14665,N_14657);
and U14820 (N_14820,N_14794,N_14706);
nor U14821 (N_14821,N_14631,N_14783);
and U14822 (N_14822,N_14712,N_14714);
nand U14823 (N_14823,N_14748,N_14677);
and U14824 (N_14824,N_14759,N_14658);
xor U14825 (N_14825,N_14680,N_14693);
and U14826 (N_14826,N_14798,N_14666);
and U14827 (N_14827,N_14751,N_14771);
xnor U14828 (N_14828,N_14640,N_14670);
and U14829 (N_14829,N_14616,N_14610);
nor U14830 (N_14830,N_14733,N_14791);
nor U14831 (N_14831,N_14704,N_14672);
xnor U14832 (N_14832,N_14614,N_14717);
nor U14833 (N_14833,N_14752,N_14780);
and U14834 (N_14834,N_14698,N_14790);
xor U14835 (N_14835,N_14732,N_14797);
nand U14836 (N_14836,N_14787,N_14789);
xor U14837 (N_14837,N_14731,N_14615);
or U14838 (N_14838,N_14676,N_14707);
nor U14839 (N_14839,N_14709,N_14611);
nor U14840 (N_14840,N_14696,N_14769);
xnor U14841 (N_14841,N_14726,N_14622);
xnor U14842 (N_14842,N_14786,N_14697);
xnor U14843 (N_14843,N_14708,N_14777);
or U14844 (N_14844,N_14713,N_14745);
xor U14845 (N_14845,N_14646,N_14645);
nor U14846 (N_14846,N_14662,N_14686);
nor U14847 (N_14847,N_14600,N_14747);
or U14848 (N_14848,N_14764,N_14788);
and U14849 (N_14849,N_14629,N_14721);
nor U14850 (N_14850,N_14668,N_14724);
and U14851 (N_14851,N_14702,N_14648);
xnor U14852 (N_14852,N_14643,N_14799);
nor U14853 (N_14853,N_14772,N_14617);
xnor U14854 (N_14854,N_14716,N_14741);
nor U14855 (N_14855,N_14744,N_14652);
xor U14856 (N_14856,N_14637,N_14684);
nand U14857 (N_14857,N_14762,N_14602);
and U14858 (N_14858,N_14767,N_14763);
and U14859 (N_14859,N_14736,N_14734);
nor U14860 (N_14860,N_14749,N_14742);
xor U14861 (N_14861,N_14626,N_14690);
or U14862 (N_14862,N_14687,N_14701);
and U14863 (N_14863,N_14671,N_14604);
or U14864 (N_14864,N_14785,N_14689);
nand U14865 (N_14865,N_14627,N_14729);
or U14866 (N_14866,N_14718,N_14725);
and U14867 (N_14867,N_14606,N_14655);
and U14868 (N_14868,N_14607,N_14603);
or U14869 (N_14869,N_14715,N_14746);
xor U14870 (N_14870,N_14621,N_14727);
and U14871 (N_14871,N_14795,N_14678);
nand U14872 (N_14872,N_14738,N_14628);
nor U14873 (N_14873,N_14653,N_14755);
xnor U14874 (N_14874,N_14784,N_14722);
and U14875 (N_14875,N_14674,N_14638);
xor U14876 (N_14876,N_14692,N_14760);
xor U14877 (N_14877,N_14630,N_14740);
xor U14878 (N_14878,N_14768,N_14633);
and U14879 (N_14879,N_14735,N_14793);
nor U14880 (N_14880,N_14753,N_14635);
and U14881 (N_14881,N_14781,N_14766);
nor U14882 (N_14882,N_14682,N_14705);
xor U14883 (N_14883,N_14618,N_14663);
nand U14884 (N_14884,N_14624,N_14632);
xor U14885 (N_14885,N_14609,N_14710);
or U14886 (N_14886,N_14730,N_14761);
xor U14887 (N_14887,N_14685,N_14673);
xnor U14888 (N_14888,N_14757,N_14773);
xor U14889 (N_14889,N_14613,N_14691);
xnor U14890 (N_14890,N_14695,N_14608);
and U14891 (N_14891,N_14699,N_14667);
nor U14892 (N_14892,N_14601,N_14636);
nor U14893 (N_14893,N_14656,N_14775);
nand U14894 (N_14894,N_14719,N_14660);
xnor U14895 (N_14895,N_14625,N_14782);
xor U14896 (N_14896,N_14654,N_14728);
nor U14897 (N_14897,N_14623,N_14651);
nor U14898 (N_14898,N_14778,N_14641);
and U14899 (N_14899,N_14679,N_14619);
nor U14900 (N_14900,N_14632,N_14662);
or U14901 (N_14901,N_14704,N_14752);
xnor U14902 (N_14902,N_14712,N_14748);
xnor U14903 (N_14903,N_14780,N_14617);
or U14904 (N_14904,N_14661,N_14744);
nand U14905 (N_14905,N_14752,N_14750);
xor U14906 (N_14906,N_14702,N_14772);
xor U14907 (N_14907,N_14614,N_14692);
xor U14908 (N_14908,N_14725,N_14643);
xnor U14909 (N_14909,N_14760,N_14653);
nand U14910 (N_14910,N_14621,N_14604);
nand U14911 (N_14911,N_14636,N_14696);
xnor U14912 (N_14912,N_14636,N_14690);
or U14913 (N_14913,N_14707,N_14701);
nor U14914 (N_14914,N_14683,N_14750);
xnor U14915 (N_14915,N_14771,N_14769);
nor U14916 (N_14916,N_14728,N_14621);
nand U14917 (N_14917,N_14629,N_14660);
nand U14918 (N_14918,N_14748,N_14773);
nor U14919 (N_14919,N_14680,N_14665);
xor U14920 (N_14920,N_14648,N_14637);
nor U14921 (N_14921,N_14602,N_14672);
and U14922 (N_14922,N_14768,N_14787);
and U14923 (N_14923,N_14692,N_14612);
and U14924 (N_14924,N_14632,N_14601);
and U14925 (N_14925,N_14682,N_14724);
nor U14926 (N_14926,N_14799,N_14768);
or U14927 (N_14927,N_14643,N_14685);
and U14928 (N_14928,N_14645,N_14647);
xnor U14929 (N_14929,N_14797,N_14711);
and U14930 (N_14930,N_14745,N_14607);
nor U14931 (N_14931,N_14706,N_14702);
xnor U14932 (N_14932,N_14772,N_14777);
nand U14933 (N_14933,N_14611,N_14745);
nor U14934 (N_14934,N_14770,N_14704);
or U14935 (N_14935,N_14605,N_14619);
nor U14936 (N_14936,N_14649,N_14621);
nor U14937 (N_14937,N_14671,N_14613);
or U14938 (N_14938,N_14733,N_14713);
and U14939 (N_14939,N_14746,N_14676);
and U14940 (N_14940,N_14658,N_14692);
xor U14941 (N_14941,N_14677,N_14616);
nor U14942 (N_14942,N_14709,N_14718);
or U14943 (N_14943,N_14758,N_14798);
nand U14944 (N_14944,N_14687,N_14781);
nand U14945 (N_14945,N_14614,N_14649);
and U14946 (N_14946,N_14718,N_14606);
xor U14947 (N_14947,N_14763,N_14759);
xnor U14948 (N_14948,N_14669,N_14678);
nand U14949 (N_14949,N_14635,N_14775);
and U14950 (N_14950,N_14762,N_14612);
nand U14951 (N_14951,N_14728,N_14774);
nand U14952 (N_14952,N_14605,N_14697);
nand U14953 (N_14953,N_14699,N_14622);
xnor U14954 (N_14954,N_14755,N_14726);
nand U14955 (N_14955,N_14756,N_14728);
nor U14956 (N_14956,N_14781,N_14764);
or U14957 (N_14957,N_14702,N_14671);
or U14958 (N_14958,N_14755,N_14672);
and U14959 (N_14959,N_14612,N_14737);
and U14960 (N_14960,N_14624,N_14797);
and U14961 (N_14961,N_14753,N_14724);
and U14962 (N_14962,N_14634,N_14713);
or U14963 (N_14963,N_14694,N_14702);
or U14964 (N_14964,N_14683,N_14775);
nor U14965 (N_14965,N_14630,N_14706);
nand U14966 (N_14966,N_14702,N_14744);
nand U14967 (N_14967,N_14725,N_14665);
nor U14968 (N_14968,N_14658,N_14702);
or U14969 (N_14969,N_14730,N_14712);
nor U14970 (N_14970,N_14655,N_14711);
nor U14971 (N_14971,N_14715,N_14738);
and U14972 (N_14972,N_14618,N_14689);
and U14973 (N_14973,N_14643,N_14703);
xnor U14974 (N_14974,N_14734,N_14621);
nand U14975 (N_14975,N_14741,N_14670);
xnor U14976 (N_14976,N_14637,N_14718);
nor U14977 (N_14977,N_14721,N_14715);
and U14978 (N_14978,N_14647,N_14738);
nand U14979 (N_14979,N_14761,N_14788);
nor U14980 (N_14980,N_14739,N_14743);
and U14981 (N_14981,N_14641,N_14660);
and U14982 (N_14982,N_14669,N_14640);
nand U14983 (N_14983,N_14728,N_14795);
nand U14984 (N_14984,N_14622,N_14631);
nand U14985 (N_14985,N_14712,N_14762);
xor U14986 (N_14986,N_14790,N_14765);
xnor U14987 (N_14987,N_14698,N_14620);
nor U14988 (N_14988,N_14633,N_14749);
and U14989 (N_14989,N_14795,N_14656);
nor U14990 (N_14990,N_14601,N_14666);
nand U14991 (N_14991,N_14749,N_14658);
xnor U14992 (N_14992,N_14684,N_14736);
nand U14993 (N_14993,N_14799,N_14792);
or U14994 (N_14994,N_14688,N_14610);
or U14995 (N_14995,N_14678,N_14655);
nand U14996 (N_14996,N_14664,N_14638);
xnor U14997 (N_14997,N_14751,N_14647);
and U14998 (N_14998,N_14766,N_14606);
and U14999 (N_14999,N_14772,N_14734);
xor U15000 (N_15000,N_14940,N_14881);
nor U15001 (N_15001,N_14834,N_14813);
or U15002 (N_15002,N_14959,N_14835);
nand U15003 (N_15003,N_14981,N_14846);
nor U15004 (N_15004,N_14971,N_14926);
nand U15005 (N_15005,N_14919,N_14840);
or U15006 (N_15006,N_14934,N_14836);
and U15007 (N_15007,N_14831,N_14848);
xor U15008 (N_15008,N_14823,N_14904);
and U15009 (N_15009,N_14833,N_14930);
and U15010 (N_15010,N_14884,N_14993);
and U15011 (N_15011,N_14973,N_14924);
and U15012 (N_15012,N_14824,N_14969);
or U15013 (N_15013,N_14898,N_14986);
nand U15014 (N_15014,N_14911,N_14918);
nor U15015 (N_15015,N_14978,N_14941);
nand U15016 (N_15016,N_14950,N_14912);
nand U15017 (N_15017,N_14989,N_14822);
nor U15018 (N_15018,N_14841,N_14885);
xnor U15019 (N_15019,N_14997,N_14827);
nand U15020 (N_15020,N_14920,N_14803);
and U15021 (N_15021,N_14817,N_14850);
xnor U15022 (N_15022,N_14802,N_14873);
and U15023 (N_15023,N_14857,N_14985);
or U15024 (N_15024,N_14999,N_14921);
nand U15025 (N_15025,N_14821,N_14874);
nand U15026 (N_15026,N_14838,N_14937);
nor U15027 (N_15027,N_14829,N_14843);
nor U15028 (N_15028,N_14809,N_14979);
and U15029 (N_15029,N_14892,N_14845);
and U15030 (N_15030,N_14878,N_14984);
nor U15031 (N_15031,N_14945,N_14807);
and U15032 (N_15032,N_14887,N_14805);
nand U15033 (N_15033,N_14909,N_14871);
and U15034 (N_15034,N_14965,N_14900);
nand U15035 (N_15035,N_14812,N_14820);
or U15036 (N_15036,N_14972,N_14907);
nand U15037 (N_15037,N_14991,N_14872);
and U15038 (N_15038,N_14890,N_14929);
and U15039 (N_15039,N_14957,N_14863);
and U15040 (N_15040,N_14992,N_14830);
nor U15041 (N_15041,N_14927,N_14886);
or U15042 (N_15042,N_14931,N_14851);
nor U15043 (N_15043,N_14966,N_14854);
nor U15044 (N_15044,N_14906,N_14865);
nand U15045 (N_15045,N_14867,N_14987);
xor U15046 (N_15046,N_14858,N_14896);
and U15047 (N_15047,N_14853,N_14808);
xnor U15048 (N_15048,N_14968,N_14925);
nor U15049 (N_15049,N_14928,N_14977);
or U15050 (N_15050,N_14958,N_14902);
nand U15051 (N_15051,N_14883,N_14839);
and U15052 (N_15052,N_14814,N_14894);
xor U15053 (N_15053,N_14888,N_14893);
and U15054 (N_15054,N_14905,N_14889);
and U15055 (N_15055,N_14870,N_14879);
nand U15056 (N_15056,N_14882,N_14951);
xnor U15057 (N_15057,N_14939,N_14856);
and U15058 (N_15058,N_14903,N_14864);
and U15059 (N_15059,N_14988,N_14914);
nor U15060 (N_15060,N_14946,N_14962);
and U15061 (N_15061,N_14936,N_14956);
or U15062 (N_15062,N_14899,N_14947);
nand U15063 (N_15063,N_14942,N_14983);
nor U15064 (N_15064,N_14818,N_14970);
xor U15065 (N_15065,N_14967,N_14815);
nand U15066 (N_15066,N_14897,N_14855);
xnor U15067 (N_15067,N_14908,N_14861);
nor U15068 (N_15068,N_14922,N_14825);
and U15069 (N_15069,N_14837,N_14826);
nand U15070 (N_15070,N_14955,N_14891);
nor U15071 (N_15071,N_14995,N_14868);
and U15072 (N_15072,N_14869,N_14953);
nand U15073 (N_15073,N_14806,N_14996);
nand U15074 (N_15074,N_14954,N_14923);
nand U15075 (N_15075,N_14933,N_14917);
xor U15076 (N_15076,N_14943,N_14810);
xnor U15077 (N_15077,N_14880,N_14982);
xnor U15078 (N_15078,N_14938,N_14866);
or U15079 (N_15079,N_14832,N_14944);
nand U15080 (N_15080,N_14862,N_14915);
nand U15081 (N_15081,N_14932,N_14828);
nor U15082 (N_15082,N_14816,N_14860);
nand U15083 (N_15083,N_14847,N_14842);
xnor U15084 (N_15084,N_14804,N_14819);
nor U15085 (N_15085,N_14960,N_14875);
nor U15086 (N_15086,N_14963,N_14948);
nor U15087 (N_15087,N_14949,N_14913);
xor U15088 (N_15088,N_14877,N_14994);
xnor U15089 (N_15089,N_14964,N_14976);
nand U15090 (N_15090,N_14852,N_14901);
nand U15091 (N_15091,N_14801,N_14800);
nor U15092 (N_15092,N_14916,N_14961);
nand U15093 (N_15093,N_14849,N_14876);
nor U15094 (N_15094,N_14980,N_14895);
nand U15095 (N_15095,N_14990,N_14935);
nor U15096 (N_15096,N_14844,N_14952);
xnor U15097 (N_15097,N_14910,N_14974);
and U15098 (N_15098,N_14998,N_14811);
or U15099 (N_15099,N_14975,N_14859);
nand U15100 (N_15100,N_14888,N_14941);
and U15101 (N_15101,N_14988,N_14906);
nor U15102 (N_15102,N_14805,N_14931);
and U15103 (N_15103,N_14900,N_14986);
nand U15104 (N_15104,N_14944,N_14950);
nor U15105 (N_15105,N_14951,N_14866);
nand U15106 (N_15106,N_14887,N_14936);
or U15107 (N_15107,N_14940,N_14808);
nand U15108 (N_15108,N_14978,N_14866);
and U15109 (N_15109,N_14934,N_14991);
and U15110 (N_15110,N_14988,N_14900);
nand U15111 (N_15111,N_14821,N_14851);
or U15112 (N_15112,N_14880,N_14838);
nand U15113 (N_15113,N_14953,N_14961);
xor U15114 (N_15114,N_14912,N_14805);
or U15115 (N_15115,N_14968,N_14910);
nor U15116 (N_15116,N_14832,N_14889);
or U15117 (N_15117,N_14839,N_14802);
xnor U15118 (N_15118,N_14867,N_14918);
xnor U15119 (N_15119,N_14933,N_14914);
xor U15120 (N_15120,N_14871,N_14921);
nor U15121 (N_15121,N_14861,N_14873);
xnor U15122 (N_15122,N_14849,N_14887);
and U15123 (N_15123,N_14941,N_14804);
nor U15124 (N_15124,N_14971,N_14829);
and U15125 (N_15125,N_14833,N_14864);
xnor U15126 (N_15126,N_14828,N_14942);
nand U15127 (N_15127,N_14853,N_14846);
nor U15128 (N_15128,N_14890,N_14870);
nor U15129 (N_15129,N_14807,N_14827);
xor U15130 (N_15130,N_14946,N_14882);
and U15131 (N_15131,N_14811,N_14963);
nand U15132 (N_15132,N_14962,N_14819);
xnor U15133 (N_15133,N_14912,N_14943);
or U15134 (N_15134,N_14870,N_14854);
nor U15135 (N_15135,N_14966,N_14882);
nand U15136 (N_15136,N_14871,N_14897);
nor U15137 (N_15137,N_14906,N_14946);
xor U15138 (N_15138,N_14809,N_14841);
nand U15139 (N_15139,N_14876,N_14948);
nor U15140 (N_15140,N_14957,N_14862);
xor U15141 (N_15141,N_14892,N_14857);
nor U15142 (N_15142,N_14977,N_14933);
nand U15143 (N_15143,N_14956,N_14949);
or U15144 (N_15144,N_14960,N_14852);
and U15145 (N_15145,N_14841,N_14846);
nor U15146 (N_15146,N_14844,N_14919);
nand U15147 (N_15147,N_14866,N_14903);
nand U15148 (N_15148,N_14828,N_14947);
nor U15149 (N_15149,N_14950,N_14871);
xnor U15150 (N_15150,N_14817,N_14996);
xor U15151 (N_15151,N_14909,N_14840);
and U15152 (N_15152,N_14902,N_14883);
nor U15153 (N_15153,N_14819,N_14908);
nor U15154 (N_15154,N_14897,N_14877);
or U15155 (N_15155,N_14851,N_14995);
or U15156 (N_15156,N_14943,N_14941);
xor U15157 (N_15157,N_14836,N_14927);
xor U15158 (N_15158,N_14952,N_14981);
nand U15159 (N_15159,N_14944,N_14925);
nor U15160 (N_15160,N_14844,N_14821);
nor U15161 (N_15161,N_14912,N_14860);
xnor U15162 (N_15162,N_14965,N_14988);
nand U15163 (N_15163,N_14937,N_14842);
nand U15164 (N_15164,N_14862,N_14951);
nand U15165 (N_15165,N_14837,N_14828);
xor U15166 (N_15166,N_14814,N_14991);
nor U15167 (N_15167,N_14943,N_14969);
and U15168 (N_15168,N_14818,N_14884);
and U15169 (N_15169,N_14972,N_14964);
or U15170 (N_15170,N_14822,N_14814);
nor U15171 (N_15171,N_14913,N_14923);
nand U15172 (N_15172,N_14912,N_14864);
nor U15173 (N_15173,N_14848,N_14981);
or U15174 (N_15174,N_14846,N_14851);
or U15175 (N_15175,N_14807,N_14896);
nor U15176 (N_15176,N_14981,N_14932);
nor U15177 (N_15177,N_14926,N_14827);
nor U15178 (N_15178,N_14951,N_14944);
nor U15179 (N_15179,N_14847,N_14871);
and U15180 (N_15180,N_14849,N_14943);
or U15181 (N_15181,N_14926,N_14917);
and U15182 (N_15182,N_14872,N_14849);
nor U15183 (N_15183,N_14843,N_14967);
xor U15184 (N_15184,N_14842,N_14802);
or U15185 (N_15185,N_14948,N_14997);
xnor U15186 (N_15186,N_14995,N_14908);
nand U15187 (N_15187,N_14914,N_14967);
nor U15188 (N_15188,N_14800,N_14839);
nor U15189 (N_15189,N_14908,N_14809);
nand U15190 (N_15190,N_14970,N_14905);
nand U15191 (N_15191,N_14875,N_14866);
or U15192 (N_15192,N_14930,N_14874);
nand U15193 (N_15193,N_14918,N_14894);
nor U15194 (N_15194,N_14976,N_14807);
and U15195 (N_15195,N_14939,N_14922);
and U15196 (N_15196,N_14957,N_14903);
nor U15197 (N_15197,N_14893,N_14897);
nand U15198 (N_15198,N_14843,N_14996);
nand U15199 (N_15199,N_14942,N_14875);
xnor U15200 (N_15200,N_15160,N_15057);
nand U15201 (N_15201,N_15159,N_15051);
nor U15202 (N_15202,N_15068,N_15154);
and U15203 (N_15203,N_15048,N_15029);
nor U15204 (N_15204,N_15071,N_15149);
or U15205 (N_15205,N_15104,N_15103);
nor U15206 (N_15206,N_15046,N_15012);
xor U15207 (N_15207,N_15123,N_15036);
xnor U15208 (N_15208,N_15096,N_15176);
nor U15209 (N_15209,N_15007,N_15117);
or U15210 (N_15210,N_15185,N_15078);
xor U15211 (N_15211,N_15132,N_15105);
or U15212 (N_15212,N_15082,N_15147);
xnor U15213 (N_15213,N_15014,N_15191);
nand U15214 (N_15214,N_15120,N_15075);
nor U15215 (N_15215,N_15086,N_15166);
or U15216 (N_15216,N_15087,N_15076);
nand U15217 (N_15217,N_15034,N_15010);
xnor U15218 (N_15218,N_15140,N_15153);
nor U15219 (N_15219,N_15139,N_15148);
xor U15220 (N_15220,N_15188,N_15027);
nand U15221 (N_15221,N_15035,N_15002);
xnor U15222 (N_15222,N_15001,N_15156);
nand U15223 (N_15223,N_15128,N_15137);
xnor U15224 (N_15224,N_15026,N_15006);
nand U15225 (N_15225,N_15170,N_15152);
nand U15226 (N_15226,N_15088,N_15031);
or U15227 (N_15227,N_15172,N_15066);
nor U15228 (N_15228,N_15171,N_15193);
nor U15229 (N_15229,N_15119,N_15025);
nand U15230 (N_15230,N_15008,N_15135);
or U15231 (N_15231,N_15095,N_15106);
nand U15232 (N_15232,N_15072,N_15009);
or U15233 (N_15233,N_15146,N_15126);
and U15234 (N_15234,N_15199,N_15158);
xnor U15235 (N_15235,N_15060,N_15004);
or U15236 (N_15236,N_15033,N_15097);
nor U15237 (N_15237,N_15041,N_15050);
nor U15238 (N_15238,N_15168,N_15080);
and U15239 (N_15239,N_15094,N_15114);
or U15240 (N_15240,N_15013,N_15196);
or U15241 (N_15241,N_15183,N_15059);
xor U15242 (N_15242,N_15067,N_15182);
and U15243 (N_15243,N_15047,N_15063);
and U15244 (N_15244,N_15024,N_15052);
xnor U15245 (N_15245,N_15092,N_15016);
and U15246 (N_15246,N_15110,N_15161);
xnor U15247 (N_15247,N_15023,N_15115);
nand U15248 (N_15248,N_15181,N_15125);
nand U15249 (N_15249,N_15157,N_15037);
or U15250 (N_15250,N_15020,N_15102);
nor U15251 (N_15251,N_15089,N_15058);
nand U15252 (N_15252,N_15073,N_15129);
nand U15253 (N_15253,N_15151,N_15111);
nand U15254 (N_15254,N_15098,N_15169);
nand U15255 (N_15255,N_15138,N_15091);
and U15256 (N_15256,N_15133,N_15043);
or U15257 (N_15257,N_15093,N_15040);
or U15258 (N_15258,N_15175,N_15134);
nand U15259 (N_15259,N_15085,N_15142);
nor U15260 (N_15260,N_15165,N_15017);
or U15261 (N_15261,N_15167,N_15022);
nand U15262 (N_15262,N_15042,N_15194);
xor U15263 (N_15263,N_15056,N_15011);
and U15264 (N_15264,N_15064,N_15179);
nand U15265 (N_15265,N_15124,N_15174);
nand U15266 (N_15266,N_15065,N_15053);
nor U15267 (N_15267,N_15186,N_15099);
xnor U15268 (N_15268,N_15187,N_15018);
and U15269 (N_15269,N_15044,N_15021);
xor U15270 (N_15270,N_15145,N_15101);
nand U15271 (N_15271,N_15000,N_15150);
nor U15272 (N_15272,N_15061,N_15030);
xor U15273 (N_15273,N_15107,N_15003);
or U15274 (N_15274,N_15131,N_15141);
and U15275 (N_15275,N_15109,N_15192);
xnor U15276 (N_15276,N_15162,N_15081);
and U15277 (N_15277,N_15070,N_15015);
xnor U15278 (N_15278,N_15077,N_15032);
or U15279 (N_15279,N_15164,N_15074);
and U15280 (N_15280,N_15144,N_15005);
or U15281 (N_15281,N_15127,N_15116);
or U15282 (N_15282,N_15195,N_15121);
nor U15283 (N_15283,N_15197,N_15069);
nand U15284 (N_15284,N_15039,N_15118);
or U15285 (N_15285,N_15143,N_15108);
nand U15286 (N_15286,N_15079,N_15184);
and U15287 (N_15287,N_15084,N_15100);
and U15288 (N_15288,N_15112,N_15054);
nand U15289 (N_15289,N_15062,N_15136);
or U15290 (N_15290,N_15049,N_15019);
or U15291 (N_15291,N_15045,N_15122);
xor U15292 (N_15292,N_15173,N_15038);
nand U15293 (N_15293,N_15189,N_15055);
nand U15294 (N_15294,N_15177,N_15028);
and U15295 (N_15295,N_15163,N_15198);
and U15296 (N_15296,N_15155,N_15083);
nand U15297 (N_15297,N_15113,N_15090);
nor U15298 (N_15298,N_15130,N_15178);
nand U15299 (N_15299,N_15190,N_15180);
and U15300 (N_15300,N_15148,N_15001);
nor U15301 (N_15301,N_15154,N_15138);
nand U15302 (N_15302,N_15006,N_15176);
nand U15303 (N_15303,N_15061,N_15115);
nor U15304 (N_15304,N_15183,N_15164);
and U15305 (N_15305,N_15184,N_15013);
and U15306 (N_15306,N_15070,N_15197);
or U15307 (N_15307,N_15183,N_15172);
and U15308 (N_15308,N_15182,N_15127);
nor U15309 (N_15309,N_15109,N_15032);
nor U15310 (N_15310,N_15068,N_15079);
and U15311 (N_15311,N_15031,N_15165);
nand U15312 (N_15312,N_15076,N_15044);
nand U15313 (N_15313,N_15055,N_15018);
xor U15314 (N_15314,N_15147,N_15047);
nor U15315 (N_15315,N_15052,N_15089);
nand U15316 (N_15316,N_15086,N_15172);
nor U15317 (N_15317,N_15097,N_15169);
and U15318 (N_15318,N_15124,N_15182);
nor U15319 (N_15319,N_15007,N_15020);
xor U15320 (N_15320,N_15141,N_15174);
nor U15321 (N_15321,N_15189,N_15195);
xor U15322 (N_15322,N_15116,N_15015);
nor U15323 (N_15323,N_15064,N_15111);
and U15324 (N_15324,N_15082,N_15194);
and U15325 (N_15325,N_15098,N_15018);
or U15326 (N_15326,N_15182,N_15195);
and U15327 (N_15327,N_15192,N_15153);
or U15328 (N_15328,N_15132,N_15119);
or U15329 (N_15329,N_15169,N_15091);
nor U15330 (N_15330,N_15135,N_15044);
xnor U15331 (N_15331,N_15172,N_15087);
or U15332 (N_15332,N_15193,N_15102);
xor U15333 (N_15333,N_15167,N_15124);
or U15334 (N_15334,N_15007,N_15161);
or U15335 (N_15335,N_15144,N_15083);
or U15336 (N_15336,N_15135,N_15188);
nor U15337 (N_15337,N_15089,N_15034);
nand U15338 (N_15338,N_15189,N_15171);
nand U15339 (N_15339,N_15072,N_15170);
or U15340 (N_15340,N_15186,N_15022);
nand U15341 (N_15341,N_15085,N_15028);
nor U15342 (N_15342,N_15076,N_15022);
xnor U15343 (N_15343,N_15001,N_15149);
or U15344 (N_15344,N_15099,N_15089);
or U15345 (N_15345,N_15072,N_15169);
and U15346 (N_15346,N_15055,N_15141);
or U15347 (N_15347,N_15184,N_15105);
or U15348 (N_15348,N_15029,N_15167);
xnor U15349 (N_15349,N_15166,N_15142);
xnor U15350 (N_15350,N_15182,N_15048);
xor U15351 (N_15351,N_15000,N_15085);
nor U15352 (N_15352,N_15038,N_15116);
nand U15353 (N_15353,N_15082,N_15101);
nand U15354 (N_15354,N_15118,N_15197);
nand U15355 (N_15355,N_15028,N_15120);
nor U15356 (N_15356,N_15062,N_15133);
nor U15357 (N_15357,N_15013,N_15191);
nor U15358 (N_15358,N_15004,N_15068);
or U15359 (N_15359,N_15146,N_15003);
and U15360 (N_15360,N_15105,N_15040);
nor U15361 (N_15361,N_15021,N_15031);
nor U15362 (N_15362,N_15023,N_15011);
xor U15363 (N_15363,N_15064,N_15143);
and U15364 (N_15364,N_15159,N_15026);
nand U15365 (N_15365,N_15117,N_15030);
nor U15366 (N_15366,N_15015,N_15137);
nand U15367 (N_15367,N_15099,N_15194);
xnor U15368 (N_15368,N_15106,N_15094);
nor U15369 (N_15369,N_15156,N_15048);
or U15370 (N_15370,N_15019,N_15193);
xor U15371 (N_15371,N_15002,N_15187);
and U15372 (N_15372,N_15121,N_15070);
and U15373 (N_15373,N_15193,N_15034);
xnor U15374 (N_15374,N_15101,N_15033);
and U15375 (N_15375,N_15114,N_15007);
nor U15376 (N_15376,N_15163,N_15013);
and U15377 (N_15377,N_15198,N_15000);
and U15378 (N_15378,N_15131,N_15161);
nor U15379 (N_15379,N_15075,N_15089);
or U15380 (N_15380,N_15002,N_15198);
nor U15381 (N_15381,N_15011,N_15139);
nand U15382 (N_15382,N_15023,N_15122);
nor U15383 (N_15383,N_15052,N_15157);
nand U15384 (N_15384,N_15095,N_15142);
nor U15385 (N_15385,N_15182,N_15186);
and U15386 (N_15386,N_15139,N_15003);
nor U15387 (N_15387,N_15153,N_15095);
nor U15388 (N_15388,N_15067,N_15074);
nor U15389 (N_15389,N_15155,N_15060);
nor U15390 (N_15390,N_15060,N_15154);
and U15391 (N_15391,N_15170,N_15124);
and U15392 (N_15392,N_15093,N_15181);
and U15393 (N_15393,N_15069,N_15140);
and U15394 (N_15394,N_15038,N_15111);
and U15395 (N_15395,N_15015,N_15098);
xnor U15396 (N_15396,N_15066,N_15188);
and U15397 (N_15397,N_15149,N_15110);
nor U15398 (N_15398,N_15050,N_15121);
or U15399 (N_15399,N_15136,N_15150);
nor U15400 (N_15400,N_15379,N_15389);
and U15401 (N_15401,N_15235,N_15260);
nor U15402 (N_15402,N_15208,N_15300);
or U15403 (N_15403,N_15291,N_15398);
xnor U15404 (N_15404,N_15223,N_15392);
or U15405 (N_15405,N_15391,N_15282);
nand U15406 (N_15406,N_15278,N_15355);
nand U15407 (N_15407,N_15242,N_15340);
or U15408 (N_15408,N_15368,N_15248);
nor U15409 (N_15409,N_15207,N_15285);
nand U15410 (N_15410,N_15352,N_15206);
nor U15411 (N_15411,N_15220,N_15262);
nor U15412 (N_15412,N_15396,N_15232);
nor U15413 (N_15413,N_15313,N_15289);
or U15414 (N_15414,N_15348,N_15323);
nand U15415 (N_15415,N_15341,N_15266);
and U15416 (N_15416,N_15339,N_15205);
or U15417 (N_15417,N_15252,N_15351);
or U15418 (N_15418,N_15336,N_15247);
nand U15419 (N_15419,N_15342,N_15297);
nand U15420 (N_15420,N_15337,N_15239);
nand U15421 (N_15421,N_15306,N_15274);
and U15422 (N_15422,N_15222,N_15269);
or U15423 (N_15423,N_15281,N_15203);
or U15424 (N_15424,N_15338,N_15317);
nor U15425 (N_15425,N_15374,N_15312);
xor U15426 (N_15426,N_15261,N_15387);
and U15427 (N_15427,N_15292,N_15377);
and U15428 (N_15428,N_15212,N_15303);
or U15429 (N_15429,N_15251,N_15267);
xor U15430 (N_15430,N_15202,N_15393);
xor U15431 (N_15431,N_15201,N_15354);
xor U15432 (N_15432,N_15372,N_15369);
or U15433 (N_15433,N_15390,N_15302);
nand U15434 (N_15434,N_15350,N_15326);
nor U15435 (N_15435,N_15211,N_15361);
nor U15436 (N_15436,N_15225,N_15386);
and U15437 (N_15437,N_15244,N_15305);
nand U15438 (N_15438,N_15365,N_15246);
xor U15439 (N_15439,N_15264,N_15334);
nor U15440 (N_15440,N_15200,N_15258);
xnor U15441 (N_15441,N_15324,N_15357);
nor U15442 (N_15442,N_15397,N_15359);
xor U15443 (N_15443,N_15241,N_15349);
nand U15444 (N_15444,N_15367,N_15318);
xnor U15445 (N_15445,N_15287,N_15347);
and U15446 (N_15446,N_15237,N_15279);
and U15447 (N_15447,N_15228,N_15353);
nor U15448 (N_15448,N_15322,N_15358);
or U15449 (N_15449,N_15362,N_15245);
nand U15450 (N_15450,N_15325,N_15301);
nand U15451 (N_15451,N_15366,N_15309);
xor U15452 (N_15452,N_15356,N_15376);
nand U15453 (N_15453,N_15388,N_15219);
xnor U15454 (N_15454,N_15360,N_15375);
and U15455 (N_15455,N_15363,N_15315);
xor U15456 (N_15456,N_15231,N_15328);
nor U15457 (N_15457,N_15370,N_15382);
or U15458 (N_15458,N_15335,N_15271);
and U15459 (N_15459,N_15385,N_15229);
or U15460 (N_15460,N_15394,N_15224);
nor U15461 (N_15461,N_15288,N_15236);
or U15462 (N_15462,N_15215,N_15230);
xnor U15463 (N_15463,N_15380,N_15399);
and U15464 (N_15464,N_15316,N_15364);
xnor U15465 (N_15465,N_15331,N_15332);
xnor U15466 (N_15466,N_15384,N_15214);
nor U15467 (N_15467,N_15343,N_15275);
nor U15468 (N_15468,N_15277,N_15270);
xor U15469 (N_15469,N_15254,N_15255);
nand U15470 (N_15470,N_15276,N_15273);
nand U15471 (N_15471,N_15283,N_15209);
nor U15472 (N_15472,N_15204,N_15321);
nand U15473 (N_15473,N_15243,N_15233);
nand U15474 (N_15474,N_15227,N_15320);
nor U15475 (N_15475,N_15311,N_15381);
xor U15476 (N_15476,N_15218,N_15257);
nand U15477 (N_15477,N_15272,N_15344);
or U15478 (N_15478,N_15253,N_15378);
nand U15479 (N_15479,N_15329,N_15319);
nor U15480 (N_15480,N_15210,N_15256);
xor U15481 (N_15481,N_15346,N_15265);
nor U15482 (N_15482,N_15298,N_15249);
and U15483 (N_15483,N_15290,N_15263);
nor U15484 (N_15484,N_15383,N_15216);
or U15485 (N_15485,N_15240,N_15371);
or U15486 (N_15486,N_15284,N_15333);
nand U15487 (N_15487,N_15286,N_15373);
nand U15488 (N_15488,N_15345,N_15314);
nor U15489 (N_15489,N_15395,N_15304);
or U15490 (N_15490,N_15310,N_15259);
and U15491 (N_15491,N_15250,N_15268);
or U15492 (N_15492,N_15307,N_15226);
or U15493 (N_15493,N_15217,N_15293);
or U15494 (N_15494,N_15296,N_15295);
nor U15495 (N_15495,N_15299,N_15221);
nor U15496 (N_15496,N_15280,N_15327);
or U15497 (N_15497,N_15213,N_15234);
nor U15498 (N_15498,N_15330,N_15238);
and U15499 (N_15499,N_15294,N_15308);
nand U15500 (N_15500,N_15362,N_15296);
nor U15501 (N_15501,N_15355,N_15331);
and U15502 (N_15502,N_15322,N_15393);
and U15503 (N_15503,N_15243,N_15366);
and U15504 (N_15504,N_15354,N_15219);
xor U15505 (N_15505,N_15387,N_15285);
xnor U15506 (N_15506,N_15251,N_15360);
and U15507 (N_15507,N_15200,N_15262);
or U15508 (N_15508,N_15299,N_15319);
nor U15509 (N_15509,N_15213,N_15374);
or U15510 (N_15510,N_15314,N_15297);
nand U15511 (N_15511,N_15351,N_15307);
or U15512 (N_15512,N_15231,N_15224);
nand U15513 (N_15513,N_15282,N_15256);
nor U15514 (N_15514,N_15323,N_15228);
xnor U15515 (N_15515,N_15266,N_15260);
or U15516 (N_15516,N_15281,N_15265);
or U15517 (N_15517,N_15286,N_15349);
xor U15518 (N_15518,N_15238,N_15396);
or U15519 (N_15519,N_15236,N_15367);
xor U15520 (N_15520,N_15203,N_15364);
or U15521 (N_15521,N_15222,N_15320);
nand U15522 (N_15522,N_15336,N_15271);
nand U15523 (N_15523,N_15363,N_15380);
nor U15524 (N_15524,N_15276,N_15262);
nand U15525 (N_15525,N_15390,N_15304);
xnor U15526 (N_15526,N_15352,N_15342);
nor U15527 (N_15527,N_15259,N_15397);
and U15528 (N_15528,N_15305,N_15293);
nor U15529 (N_15529,N_15346,N_15306);
nor U15530 (N_15530,N_15357,N_15375);
nor U15531 (N_15531,N_15283,N_15260);
xnor U15532 (N_15532,N_15378,N_15323);
nor U15533 (N_15533,N_15336,N_15395);
or U15534 (N_15534,N_15398,N_15320);
and U15535 (N_15535,N_15247,N_15302);
nand U15536 (N_15536,N_15232,N_15370);
and U15537 (N_15537,N_15392,N_15274);
nand U15538 (N_15538,N_15339,N_15388);
nor U15539 (N_15539,N_15352,N_15339);
nand U15540 (N_15540,N_15269,N_15321);
nor U15541 (N_15541,N_15355,N_15303);
or U15542 (N_15542,N_15277,N_15219);
nor U15543 (N_15543,N_15356,N_15251);
and U15544 (N_15544,N_15314,N_15330);
and U15545 (N_15545,N_15271,N_15235);
nor U15546 (N_15546,N_15369,N_15320);
and U15547 (N_15547,N_15393,N_15278);
xnor U15548 (N_15548,N_15214,N_15308);
or U15549 (N_15549,N_15379,N_15258);
nand U15550 (N_15550,N_15286,N_15207);
nand U15551 (N_15551,N_15389,N_15336);
nor U15552 (N_15552,N_15289,N_15371);
nand U15553 (N_15553,N_15271,N_15240);
and U15554 (N_15554,N_15357,N_15247);
nor U15555 (N_15555,N_15211,N_15209);
nand U15556 (N_15556,N_15269,N_15254);
xnor U15557 (N_15557,N_15325,N_15205);
nand U15558 (N_15558,N_15223,N_15297);
or U15559 (N_15559,N_15243,N_15253);
xor U15560 (N_15560,N_15325,N_15260);
nor U15561 (N_15561,N_15373,N_15317);
and U15562 (N_15562,N_15343,N_15207);
nand U15563 (N_15563,N_15282,N_15232);
nor U15564 (N_15564,N_15286,N_15330);
nand U15565 (N_15565,N_15333,N_15364);
and U15566 (N_15566,N_15300,N_15385);
nand U15567 (N_15567,N_15303,N_15241);
and U15568 (N_15568,N_15311,N_15302);
or U15569 (N_15569,N_15399,N_15257);
and U15570 (N_15570,N_15246,N_15272);
and U15571 (N_15571,N_15317,N_15363);
xor U15572 (N_15572,N_15205,N_15241);
or U15573 (N_15573,N_15271,N_15343);
and U15574 (N_15574,N_15227,N_15286);
or U15575 (N_15575,N_15383,N_15367);
or U15576 (N_15576,N_15375,N_15364);
or U15577 (N_15577,N_15277,N_15258);
and U15578 (N_15578,N_15317,N_15276);
nor U15579 (N_15579,N_15290,N_15333);
nand U15580 (N_15580,N_15319,N_15389);
or U15581 (N_15581,N_15336,N_15282);
and U15582 (N_15582,N_15394,N_15331);
xor U15583 (N_15583,N_15215,N_15319);
nor U15584 (N_15584,N_15376,N_15208);
nand U15585 (N_15585,N_15238,N_15241);
nand U15586 (N_15586,N_15363,N_15267);
nor U15587 (N_15587,N_15217,N_15383);
or U15588 (N_15588,N_15271,N_15248);
or U15589 (N_15589,N_15380,N_15276);
or U15590 (N_15590,N_15352,N_15202);
xnor U15591 (N_15591,N_15291,N_15258);
and U15592 (N_15592,N_15343,N_15229);
nand U15593 (N_15593,N_15276,N_15367);
and U15594 (N_15594,N_15212,N_15253);
or U15595 (N_15595,N_15213,N_15238);
xnor U15596 (N_15596,N_15350,N_15292);
or U15597 (N_15597,N_15394,N_15201);
or U15598 (N_15598,N_15396,N_15306);
xnor U15599 (N_15599,N_15289,N_15286);
nand U15600 (N_15600,N_15551,N_15427);
nor U15601 (N_15601,N_15580,N_15522);
nor U15602 (N_15602,N_15445,N_15530);
and U15603 (N_15603,N_15521,N_15447);
xnor U15604 (N_15604,N_15537,N_15555);
or U15605 (N_15605,N_15422,N_15554);
nand U15606 (N_15606,N_15564,N_15458);
nand U15607 (N_15607,N_15587,N_15579);
or U15608 (N_15608,N_15444,N_15485);
nor U15609 (N_15609,N_15431,N_15480);
xnor U15610 (N_15610,N_15596,N_15478);
nor U15611 (N_15611,N_15534,N_15471);
nand U15612 (N_15612,N_15411,N_15414);
nor U15613 (N_15613,N_15466,N_15585);
xor U15614 (N_15614,N_15540,N_15568);
nand U15615 (N_15615,N_15497,N_15509);
xor U15616 (N_15616,N_15461,N_15476);
nand U15617 (N_15617,N_15547,N_15409);
and U15618 (N_15618,N_15408,N_15533);
nor U15619 (N_15619,N_15529,N_15506);
nand U15620 (N_15620,N_15566,N_15453);
nand U15621 (N_15621,N_15516,N_15502);
nand U15622 (N_15622,N_15582,N_15570);
nor U15623 (N_15623,N_15573,N_15457);
or U15624 (N_15624,N_15459,N_15538);
xor U15625 (N_15625,N_15424,N_15452);
nor U15626 (N_15626,N_15558,N_15462);
nand U15627 (N_15627,N_15438,N_15430);
or U15628 (N_15628,N_15592,N_15565);
nor U15629 (N_15629,N_15561,N_15429);
or U15630 (N_15630,N_15496,N_15586);
nor U15631 (N_15631,N_15553,N_15559);
or U15632 (N_15632,N_15406,N_15489);
nand U15633 (N_15633,N_15400,N_15590);
nand U15634 (N_15634,N_15493,N_15451);
and U15635 (N_15635,N_15441,N_15546);
xnor U15636 (N_15636,N_15526,N_15539);
and U15637 (N_15637,N_15486,N_15487);
and U15638 (N_15638,N_15577,N_15482);
nand U15639 (N_15639,N_15563,N_15472);
nor U15640 (N_15640,N_15463,N_15569);
or U15641 (N_15641,N_15432,N_15575);
nand U15642 (N_15642,N_15571,N_15523);
xor U15643 (N_15643,N_15543,N_15528);
nand U15644 (N_15644,N_15507,N_15500);
and U15645 (N_15645,N_15420,N_15410);
xnor U15646 (N_15646,N_15455,N_15473);
xor U15647 (N_15647,N_15544,N_15419);
xnor U15648 (N_15648,N_15405,N_15518);
or U15649 (N_15649,N_15498,N_15456);
or U15650 (N_15650,N_15483,N_15599);
xnor U15651 (N_15651,N_15595,N_15415);
nand U15652 (N_15652,N_15494,N_15560);
xor U15653 (N_15653,N_15572,N_15517);
nor U15654 (N_15654,N_15401,N_15598);
nand U15655 (N_15655,N_15413,N_15481);
nor U15656 (N_15656,N_15421,N_15508);
nor U15657 (N_15657,N_15491,N_15474);
and U15658 (N_15658,N_15552,N_15511);
and U15659 (N_15659,N_15578,N_15484);
nand U15660 (N_15660,N_15425,N_15515);
or U15661 (N_15661,N_15576,N_15426);
xor U15662 (N_15662,N_15532,N_15597);
nand U15663 (N_15663,N_15514,N_15404);
and U15664 (N_15664,N_15541,N_15503);
nor U15665 (N_15665,N_15454,N_15536);
xor U15666 (N_15666,N_15435,N_15557);
nor U15667 (N_15667,N_15510,N_15535);
or U15668 (N_15668,N_15512,N_15465);
and U15669 (N_15669,N_15488,N_15556);
nor U15670 (N_15670,N_15524,N_15469);
nor U15671 (N_15671,N_15520,N_15450);
nor U15672 (N_15672,N_15449,N_15545);
nand U15673 (N_15673,N_15562,N_15423);
nand U15674 (N_15674,N_15495,N_15542);
nor U15675 (N_15675,N_15504,N_15468);
nand U15676 (N_15676,N_15479,N_15492);
and U15677 (N_15677,N_15594,N_15433);
and U15678 (N_15678,N_15464,N_15428);
nor U15679 (N_15679,N_15549,N_15475);
nor U15680 (N_15680,N_15584,N_15550);
nor U15681 (N_15681,N_15470,N_15440);
nand U15682 (N_15682,N_15416,N_15443);
or U15683 (N_15683,N_15588,N_15591);
xor U15684 (N_15684,N_15513,N_15501);
or U15685 (N_15685,N_15446,N_15593);
or U15686 (N_15686,N_15467,N_15527);
or U15687 (N_15687,N_15525,N_15434);
xor U15688 (N_15688,N_15418,N_15574);
or U15689 (N_15689,N_15460,N_15402);
nor U15690 (N_15690,N_15531,N_15499);
nand U15691 (N_15691,N_15490,N_15548);
and U15692 (N_15692,N_15567,N_15505);
and U15693 (N_15693,N_15417,N_15519);
nand U15694 (N_15694,N_15436,N_15412);
or U15695 (N_15695,N_15442,N_15581);
nand U15696 (N_15696,N_15589,N_15477);
nand U15697 (N_15697,N_15583,N_15448);
xor U15698 (N_15698,N_15439,N_15437);
nor U15699 (N_15699,N_15403,N_15407);
nand U15700 (N_15700,N_15499,N_15420);
and U15701 (N_15701,N_15464,N_15547);
nor U15702 (N_15702,N_15451,N_15516);
or U15703 (N_15703,N_15453,N_15411);
xor U15704 (N_15704,N_15411,N_15452);
or U15705 (N_15705,N_15405,N_15535);
xor U15706 (N_15706,N_15416,N_15468);
or U15707 (N_15707,N_15546,N_15543);
and U15708 (N_15708,N_15417,N_15528);
and U15709 (N_15709,N_15456,N_15524);
or U15710 (N_15710,N_15535,N_15558);
nand U15711 (N_15711,N_15412,N_15560);
or U15712 (N_15712,N_15464,N_15495);
xnor U15713 (N_15713,N_15422,N_15514);
or U15714 (N_15714,N_15552,N_15595);
nand U15715 (N_15715,N_15498,N_15503);
xor U15716 (N_15716,N_15597,N_15595);
nor U15717 (N_15717,N_15473,N_15413);
nand U15718 (N_15718,N_15551,N_15454);
nand U15719 (N_15719,N_15452,N_15536);
xnor U15720 (N_15720,N_15482,N_15555);
xnor U15721 (N_15721,N_15592,N_15542);
nor U15722 (N_15722,N_15595,N_15507);
xnor U15723 (N_15723,N_15435,N_15519);
or U15724 (N_15724,N_15498,N_15480);
nor U15725 (N_15725,N_15477,N_15485);
xor U15726 (N_15726,N_15464,N_15435);
and U15727 (N_15727,N_15489,N_15426);
or U15728 (N_15728,N_15469,N_15503);
nor U15729 (N_15729,N_15410,N_15480);
or U15730 (N_15730,N_15522,N_15401);
and U15731 (N_15731,N_15556,N_15451);
nor U15732 (N_15732,N_15489,N_15589);
nand U15733 (N_15733,N_15452,N_15576);
nand U15734 (N_15734,N_15488,N_15413);
xnor U15735 (N_15735,N_15584,N_15502);
or U15736 (N_15736,N_15558,N_15471);
and U15737 (N_15737,N_15499,N_15496);
nand U15738 (N_15738,N_15598,N_15437);
nor U15739 (N_15739,N_15509,N_15585);
or U15740 (N_15740,N_15527,N_15505);
or U15741 (N_15741,N_15431,N_15596);
and U15742 (N_15742,N_15540,N_15594);
nor U15743 (N_15743,N_15481,N_15459);
and U15744 (N_15744,N_15486,N_15546);
and U15745 (N_15745,N_15582,N_15466);
nand U15746 (N_15746,N_15461,N_15544);
and U15747 (N_15747,N_15464,N_15434);
nand U15748 (N_15748,N_15501,N_15574);
or U15749 (N_15749,N_15518,N_15433);
nand U15750 (N_15750,N_15555,N_15491);
nand U15751 (N_15751,N_15415,N_15511);
or U15752 (N_15752,N_15434,N_15479);
and U15753 (N_15753,N_15450,N_15534);
nand U15754 (N_15754,N_15538,N_15441);
xor U15755 (N_15755,N_15591,N_15592);
xnor U15756 (N_15756,N_15490,N_15442);
and U15757 (N_15757,N_15541,N_15454);
and U15758 (N_15758,N_15481,N_15544);
and U15759 (N_15759,N_15430,N_15513);
xor U15760 (N_15760,N_15564,N_15445);
and U15761 (N_15761,N_15538,N_15584);
nor U15762 (N_15762,N_15579,N_15513);
xnor U15763 (N_15763,N_15424,N_15563);
nor U15764 (N_15764,N_15566,N_15455);
nor U15765 (N_15765,N_15512,N_15423);
or U15766 (N_15766,N_15434,N_15548);
or U15767 (N_15767,N_15534,N_15586);
nor U15768 (N_15768,N_15559,N_15535);
and U15769 (N_15769,N_15410,N_15419);
xor U15770 (N_15770,N_15519,N_15560);
and U15771 (N_15771,N_15537,N_15549);
or U15772 (N_15772,N_15474,N_15557);
nand U15773 (N_15773,N_15528,N_15596);
xor U15774 (N_15774,N_15468,N_15545);
nand U15775 (N_15775,N_15409,N_15493);
xor U15776 (N_15776,N_15446,N_15567);
nor U15777 (N_15777,N_15540,N_15432);
nor U15778 (N_15778,N_15504,N_15554);
nand U15779 (N_15779,N_15441,N_15589);
xnor U15780 (N_15780,N_15471,N_15484);
nor U15781 (N_15781,N_15439,N_15428);
nand U15782 (N_15782,N_15509,N_15522);
and U15783 (N_15783,N_15483,N_15423);
and U15784 (N_15784,N_15430,N_15479);
xor U15785 (N_15785,N_15500,N_15469);
nor U15786 (N_15786,N_15528,N_15533);
or U15787 (N_15787,N_15534,N_15529);
nand U15788 (N_15788,N_15482,N_15516);
and U15789 (N_15789,N_15475,N_15497);
xor U15790 (N_15790,N_15548,N_15553);
nor U15791 (N_15791,N_15402,N_15506);
nand U15792 (N_15792,N_15448,N_15541);
nand U15793 (N_15793,N_15451,N_15474);
nand U15794 (N_15794,N_15477,N_15587);
nand U15795 (N_15795,N_15567,N_15513);
or U15796 (N_15796,N_15554,N_15410);
or U15797 (N_15797,N_15468,N_15593);
or U15798 (N_15798,N_15440,N_15575);
xor U15799 (N_15799,N_15405,N_15541);
and U15800 (N_15800,N_15667,N_15783);
nand U15801 (N_15801,N_15739,N_15621);
or U15802 (N_15802,N_15698,N_15776);
nand U15803 (N_15803,N_15614,N_15668);
and U15804 (N_15804,N_15789,N_15730);
or U15805 (N_15805,N_15695,N_15627);
xnor U15806 (N_15806,N_15705,N_15609);
xnor U15807 (N_15807,N_15674,N_15626);
nand U15808 (N_15808,N_15703,N_15729);
and U15809 (N_15809,N_15639,N_15671);
xor U15810 (N_15810,N_15625,N_15719);
nor U15811 (N_15811,N_15778,N_15612);
nor U15812 (N_15812,N_15752,N_15722);
nor U15813 (N_15813,N_15608,N_15724);
xnor U15814 (N_15814,N_15696,N_15746);
and U15815 (N_15815,N_15723,N_15602);
xor U15816 (N_15816,N_15755,N_15706);
and U15817 (N_15817,N_15782,N_15766);
nor U15818 (N_15818,N_15715,N_15613);
and U15819 (N_15819,N_15663,N_15619);
or U15820 (N_15820,N_15760,N_15700);
nand U15821 (N_15821,N_15734,N_15655);
nand U15822 (N_15822,N_15740,N_15728);
nor U15823 (N_15823,N_15630,N_15793);
and U15824 (N_15824,N_15680,N_15794);
and U15825 (N_15825,N_15676,N_15606);
nor U15826 (N_15826,N_15763,N_15745);
nand U15827 (N_15827,N_15649,N_15617);
nand U15828 (N_15828,N_15610,N_15797);
nand U15829 (N_15829,N_15768,N_15711);
and U15830 (N_15830,N_15708,N_15628);
and U15831 (N_15831,N_15647,N_15699);
xor U15832 (N_15832,N_15634,N_15772);
nor U15833 (N_15833,N_15743,N_15748);
xnor U15834 (N_15834,N_15759,N_15682);
and U15835 (N_15835,N_15732,N_15678);
or U15836 (N_15836,N_15756,N_15623);
nor U15837 (N_15837,N_15640,N_15687);
xor U15838 (N_15838,N_15721,N_15603);
nand U15839 (N_15839,N_15720,N_15707);
nand U15840 (N_15840,N_15781,N_15651);
nor U15841 (N_15841,N_15633,N_15769);
and U15842 (N_15842,N_15712,N_15774);
nor U15843 (N_15843,N_15675,N_15765);
and U15844 (N_15844,N_15615,N_15691);
or U15845 (N_15845,N_15741,N_15631);
nand U15846 (N_15846,N_15672,N_15644);
and U15847 (N_15847,N_15662,N_15679);
xor U15848 (N_15848,N_15790,N_15777);
nor U15849 (N_15849,N_15799,N_15657);
xor U15850 (N_15850,N_15636,N_15786);
and U15851 (N_15851,N_15689,N_15666);
or U15852 (N_15852,N_15725,N_15685);
nor U15853 (N_15853,N_15714,N_15648);
nand U15854 (N_15854,N_15673,N_15677);
nand U15855 (N_15855,N_15638,N_15762);
nand U15856 (N_15856,N_15758,N_15670);
nand U15857 (N_15857,N_15779,N_15664);
xnor U15858 (N_15858,N_15686,N_15737);
nand U15859 (N_15859,N_15738,N_15692);
and U15860 (N_15860,N_15771,N_15751);
nand U15861 (N_15861,N_15618,N_15694);
or U15862 (N_15862,N_15641,N_15605);
or U15863 (N_15863,N_15600,N_15716);
and U15864 (N_15864,N_15796,N_15693);
nor U15865 (N_15865,N_15749,N_15690);
nor U15866 (N_15866,N_15791,N_15611);
xor U15867 (N_15867,N_15731,N_15653);
nor U15868 (N_15868,N_15757,N_15642);
xnor U15869 (N_15869,N_15713,N_15637);
and U15870 (N_15870,N_15726,N_15697);
or U15871 (N_15871,N_15775,N_15624);
or U15872 (N_15872,N_15656,N_15709);
and U15873 (N_15873,N_15684,N_15604);
xnor U15874 (N_15874,N_15750,N_15650);
and U15875 (N_15875,N_15616,N_15784);
and U15876 (N_15876,N_15773,N_15658);
xnor U15877 (N_15877,N_15665,N_15753);
and U15878 (N_15878,N_15702,N_15727);
and U15879 (N_15879,N_15761,N_15622);
nand U15880 (N_15880,N_15733,N_15654);
nand U15881 (N_15881,N_15767,N_15792);
or U15882 (N_15882,N_15681,N_15744);
nor U15883 (N_15883,N_15747,N_15736);
or U15884 (N_15884,N_15683,N_15646);
and U15885 (N_15885,N_15704,N_15718);
nor U15886 (N_15886,N_15601,N_15688);
nor U15887 (N_15887,N_15645,N_15659);
nand U15888 (N_15888,N_15785,N_15717);
and U15889 (N_15889,N_15643,N_15635);
xnor U15890 (N_15890,N_15660,N_15607);
nand U15891 (N_15891,N_15780,N_15669);
nor U15892 (N_15892,N_15620,N_15701);
nor U15893 (N_15893,N_15735,N_15764);
nand U15894 (N_15894,N_15629,N_15742);
nand U15895 (N_15895,N_15798,N_15795);
nor U15896 (N_15896,N_15770,N_15710);
nor U15897 (N_15897,N_15788,N_15661);
nand U15898 (N_15898,N_15787,N_15632);
nor U15899 (N_15899,N_15754,N_15652);
nand U15900 (N_15900,N_15733,N_15744);
xnor U15901 (N_15901,N_15729,N_15708);
xor U15902 (N_15902,N_15653,N_15737);
nand U15903 (N_15903,N_15696,N_15628);
or U15904 (N_15904,N_15710,N_15700);
nand U15905 (N_15905,N_15763,N_15760);
and U15906 (N_15906,N_15717,N_15668);
and U15907 (N_15907,N_15762,N_15721);
nor U15908 (N_15908,N_15669,N_15656);
xnor U15909 (N_15909,N_15780,N_15604);
xnor U15910 (N_15910,N_15711,N_15664);
nand U15911 (N_15911,N_15741,N_15728);
and U15912 (N_15912,N_15719,N_15661);
nor U15913 (N_15913,N_15711,N_15698);
nand U15914 (N_15914,N_15728,N_15776);
or U15915 (N_15915,N_15685,N_15763);
or U15916 (N_15916,N_15687,N_15667);
xnor U15917 (N_15917,N_15686,N_15672);
xnor U15918 (N_15918,N_15725,N_15733);
nand U15919 (N_15919,N_15654,N_15700);
xor U15920 (N_15920,N_15673,N_15666);
nand U15921 (N_15921,N_15653,N_15649);
nand U15922 (N_15922,N_15730,N_15678);
and U15923 (N_15923,N_15756,N_15798);
or U15924 (N_15924,N_15649,N_15761);
nor U15925 (N_15925,N_15683,N_15699);
nand U15926 (N_15926,N_15750,N_15699);
xnor U15927 (N_15927,N_15607,N_15676);
nand U15928 (N_15928,N_15695,N_15755);
and U15929 (N_15929,N_15649,N_15744);
nor U15930 (N_15930,N_15632,N_15643);
nor U15931 (N_15931,N_15656,N_15776);
nand U15932 (N_15932,N_15738,N_15696);
and U15933 (N_15933,N_15654,N_15785);
or U15934 (N_15934,N_15741,N_15601);
or U15935 (N_15935,N_15638,N_15601);
nor U15936 (N_15936,N_15665,N_15796);
nor U15937 (N_15937,N_15740,N_15625);
nor U15938 (N_15938,N_15757,N_15780);
nor U15939 (N_15939,N_15614,N_15796);
xor U15940 (N_15940,N_15675,N_15734);
xor U15941 (N_15941,N_15713,N_15676);
or U15942 (N_15942,N_15622,N_15719);
nor U15943 (N_15943,N_15629,N_15718);
or U15944 (N_15944,N_15657,N_15780);
and U15945 (N_15945,N_15659,N_15641);
and U15946 (N_15946,N_15656,N_15607);
or U15947 (N_15947,N_15731,N_15791);
nor U15948 (N_15948,N_15777,N_15627);
xor U15949 (N_15949,N_15745,N_15756);
xor U15950 (N_15950,N_15629,N_15770);
nor U15951 (N_15951,N_15758,N_15765);
and U15952 (N_15952,N_15749,N_15673);
nor U15953 (N_15953,N_15789,N_15776);
nor U15954 (N_15954,N_15733,N_15625);
nand U15955 (N_15955,N_15652,N_15746);
nor U15956 (N_15956,N_15608,N_15694);
nand U15957 (N_15957,N_15743,N_15773);
nor U15958 (N_15958,N_15626,N_15744);
nand U15959 (N_15959,N_15700,N_15666);
and U15960 (N_15960,N_15762,N_15767);
nor U15961 (N_15961,N_15783,N_15645);
nor U15962 (N_15962,N_15651,N_15655);
or U15963 (N_15963,N_15628,N_15632);
nor U15964 (N_15964,N_15646,N_15775);
and U15965 (N_15965,N_15791,N_15705);
and U15966 (N_15966,N_15787,N_15685);
nand U15967 (N_15967,N_15692,N_15782);
xor U15968 (N_15968,N_15757,N_15646);
xnor U15969 (N_15969,N_15738,N_15633);
nor U15970 (N_15970,N_15727,N_15613);
xnor U15971 (N_15971,N_15763,N_15689);
and U15972 (N_15972,N_15632,N_15675);
or U15973 (N_15973,N_15704,N_15723);
xnor U15974 (N_15974,N_15693,N_15743);
xnor U15975 (N_15975,N_15681,N_15667);
or U15976 (N_15976,N_15639,N_15702);
nor U15977 (N_15977,N_15686,N_15706);
nand U15978 (N_15978,N_15695,N_15710);
nor U15979 (N_15979,N_15659,N_15654);
xor U15980 (N_15980,N_15696,N_15687);
or U15981 (N_15981,N_15732,N_15659);
or U15982 (N_15982,N_15772,N_15651);
nor U15983 (N_15983,N_15709,N_15669);
or U15984 (N_15984,N_15632,N_15613);
and U15985 (N_15985,N_15643,N_15607);
or U15986 (N_15986,N_15776,N_15685);
nand U15987 (N_15987,N_15699,N_15697);
nand U15988 (N_15988,N_15640,N_15762);
or U15989 (N_15989,N_15658,N_15623);
or U15990 (N_15990,N_15667,N_15620);
nand U15991 (N_15991,N_15637,N_15742);
or U15992 (N_15992,N_15644,N_15779);
and U15993 (N_15993,N_15794,N_15775);
and U15994 (N_15994,N_15738,N_15615);
or U15995 (N_15995,N_15660,N_15702);
xnor U15996 (N_15996,N_15640,N_15712);
xnor U15997 (N_15997,N_15605,N_15649);
and U15998 (N_15998,N_15643,N_15667);
nand U15999 (N_15999,N_15623,N_15786);
nand U16000 (N_16000,N_15816,N_15833);
xor U16001 (N_16001,N_15843,N_15993);
and U16002 (N_16002,N_15962,N_15908);
nand U16003 (N_16003,N_15865,N_15835);
or U16004 (N_16004,N_15851,N_15961);
or U16005 (N_16005,N_15874,N_15971);
nand U16006 (N_16006,N_15814,N_15911);
xnor U16007 (N_16007,N_15922,N_15978);
or U16008 (N_16008,N_15827,N_15854);
xor U16009 (N_16009,N_15974,N_15891);
or U16010 (N_16010,N_15925,N_15878);
nor U16011 (N_16011,N_15844,N_15889);
xor U16012 (N_16012,N_15886,N_15803);
and U16013 (N_16013,N_15999,N_15857);
or U16014 (N_16014,N_15919,N_15881);
nand U16015 (N_16015,N_15951,N_15855);
or U16016 (N_16016,N_15829,N_15984);
and U16017 (N_16017,N_15868,N_15997);
xor U16018 (N_16018,N_15991,N_15920);
nand U16019 (N_16019,N_15960,N_15895);
xor U16020 (N_16020,N_15907,N_15860);
or U16021 (N_16021,N_15910,N_15975);
xnor U16022 (N_16022,N_15972,N_15847);
and U16023 (N_16023,N_15936,N_15807);
nand U16024 (N_16024,N_15882,N_15846);
nand U16025 (N_16025,N_15893,N_15822);
nand U16026 (N_16026,N_15887,N_15976);
nand U16027 (N_16027,N_15856,N_15837);
and U16028 (N_16028,N_15858,N_15995);
or U16029 (N_16029,N_15823,N_15894);
nand U16030 (N_16030,N_15914,N_15985);
and U16031 (N_16031,N_15841,N_15956);
xor U16032 (N_16032,N_15811,N_15830);
and U16033 (N_16033,N_15973,N_15970);
and U16034 (N_16034,N_15957,N_15812);
nor U16035 (N_16035,N_15992,N_15953);
nand U16036 (N_16036,N_15958,N_15963);
xor U16037 (N_16037,N_15988,N_15873);
xnor U16038 (N_16038,N_15986,N_15818);
nand U16039 (N_16039,N_15998,N_15921);
xnor U16040 (N_16040,N_15923,N_15813);
xnor U16041 (N_16041,N_15896,N_15831);
xor U16042 (N_16042,N_15966,N_15864);
xnor U16043 (N_16043,N_15982,N_15915);
nor U16044 (N_16044,N_15996,N_15815);
xor U16045 (N_16045,N_15949,N_15802);
and U16046 (N_16046,N_15950,N_15934);
nand U16047 (N_16047,N_15849,N_15870);
or U16048 (N_16048,N_15862,N_15826);
or U16049 (N_16049,N_15905,N_15944);
nor U16050 (N_16050,N_15932,N_15926);
and U16051 (N_16051,N_15819,N_15883);
xor U16052 (N_16052,N_15933,N_15927);
nor U16053 (N_16053,N_15848,N_15913);
and U16054 (N_16054,N_15989,N_15924);
and U16055 (N_16055,N_15938,N_15828);
and U16056 (N_16056,N_15918,N_15810);
xnor U16057 (N_16057,N_15824,N_15877);
or U16058 (N_16058,N_15930,N_15845);
or U16059 (N_16059,N_15821,N_15850);
or U16060 (N_16060,N_15943,N_15832);
nor U16061 (N_16061,N_15861,N_15890);
and U16062 (N_16062,N_15929,N_15939);
nand U16063 (N_16063,N_15990,N_15872);
xnor U16064 (N_16064,N_15947,N_15806);
nor U16065 (N_16065,N_15880,N_15866);
or U16066 (N_16066,N_15900,N_15888);
or U16067 (N_16067,N_15903,N_15955);
and U16068 (N_16068,N_15899,N_15987);
or U16069 (N_16069,N_15838,N_15800);
or U16070 (N_16070,N_15935,N_15983);
nor U16071 (N_16071,N_15875,N_15809);
or U16072 (N_16072,N_15871,N_15968);
nand U16073 (N_16073,N_15981,N_15928);
xor U16074 (N_16074,N_15836,N_15979);
and U16075 (N_16075,N_15859,N_15853);
nand U16076 (N_16076,N_15902,N_15839);
or U16077 (N_16077,N_15959,N_15852);
nand U16078 (N_16078,N_15912,N_15884);
or U16079 (N_16079,N_15946,N_15901);
nand U16080 (N_16080,N_15892,N_15965);
nand U16081 (N_16081,N_15917,N_15994);
or U16082 (N_16082,N_15942,N_15825);
or U16083 (N_16083,N_15977,N_15967);
and U16084 (N_16084,N_15916,N_15863);
xnor U16085 (N_16085,N_15801,N_15945);
xnor U16086 (N_16086,N_15876,N_15842);
xor U16087 (N_16087,N_15948,N_15969);
nor U16088 (N_16088,N_15817,N_15805);
nor U16089 (N_16089,N_15964,N_15937);
and U16090 (N_16090,N_15840,N_15931);
nor U16091 (N_16091,N_15906,N_15879);
and U16092 (N_16092,N_15808,N_15885);
nor U16093 (N_16093,N_15804,N_15904);
xor U16094 (N_16094,N_15869,N_15897);
xnor U16095 (N_16095,N_15909,N_15940);
or U16096 (N_16096,N_15952,N_15941);
nand U16097 (N_16097,N_15834,N_15820);
and U16098 (N_16098,N_15898,N_15954);
xor U16099 (N_16099,N_15867,N_15980);
nand U16100 (N_16100,N_15946,N_15839);
nor U16101 (N_16101,N_15812,N_15846);
and U16102 (N_16102,N_15879,N_15827);
or U16103 (N_16103,N_15968,N_15802);
nand U16104 (N_16104,N_15850,N_15946);
or U16105 (N_16105,N_15966,N_15927);
nand U16106 (N_16106,N_15937,N_15913);
or U16107 (N_16107,N_15814,N_15930);
xor U16108 (N_16108,N_15828,N_15965);
and U16109 (N_16109,N_15953,N_15866);
or U16110 (N_16110,N_15846,N_15988);
and U16111 (N_16111,N_15930,N_15917);
and U16112 (N_16112,N_15949,N_15858);
nand U16113 (N_16113,N_15887,N_15861);
nand U16114 (N_16114,N_15965,N_15984);
or U16115 (N_16115,N_15920,N_15930);
and U16116 (N_16116,N_15836,N_15877);
nand U16117 (N_16117,N_15970,N_15992);
nor U16118 (N_16118,N_15833,N_15823);
xnor U16119 (N_16119,N_15823,N_15943);
xor U16120 (N_16120,N_15818,N_15844);
or U16121 (N_16121,N_15920,N_15935);
nand U16122 (N_16122,N_15836,N_15925);
nand U16123 (N_16123,N_15839,N_15865);
or U16124 (N_16124,N_15986,N_15961);
and U16125 (N_16125,N_15851,N_15999);
and U16126 (N_16126,N_15896,N_15949);
and U16127 (N_16127,N_15928,N_15844);
or U16128 (N_16128,N_15889,N_15957);
and U16129 (N_16129,N_15933,N_15944);
or U16130 (N_16130,N_15869,N_15953);
xor U16131 (N_16131,N_15983,N_15872);
xnor U16132 (N_16132,N_15876,N_15995);
and U16133 (N_16133,N_15990,N_15938);
xor U16134 (N_16134,N_15869,N_15983);
or U16135 (N_16135,N_15826,N_15944);
nor U16136 (N_16136,N_15894,N_15974);
and U16137 (N_16137,N_15909,N_15888);
xnor U16138 (N_16138,N_15825,N_15952);
xnor U16139 (N_16139,N_15996,N_15955);
nand U16140 (N_16140,N_15817,N_15854);
and U16141 (N_16141,N_15963,N_15883);
xnor U16142 (N_16142,N_15912,N_15821);
nor U16143 (N_16143,N_15895,N_15808);
nand U16144 (N_16144,N_15853,N_15865);
and U16145 (N_16145,N_15903,N_15908);
and U16146 (N_16146,N_15950,N_15814);
or U16147 (N_16147,N_15915,N_15944);
or U16148 (N_16148,N_15966,N_15865);
and U16149 (N_16149,N_15918,N_15871);
nand U16150 (N_16150,N_15937,N_15819);
xnor U16151 (N_16151,N_15949,N_15882);
nor U16152 (N_16152,N_15835,N_15958);
xor U16153 (N_16153,N_15966,N_15959);
nor U16154 (N_16154,N_15954,N_15907);
nor U16155 (N_16155,N_15906,N_15956);
or U16156 (N_16156,N_15822,N_15975);
or U16157 (N_16157,N_15863,N_15864);
or U16158 (N_16158,N_15806,N_15816);
nor U16159 (N_16159,N_15906,N_15851);
or U16160 (N_16160,N_15829,N_15921);
and U16161 (N_16161,N_15895,N_15846);
nor U16162 (N_16162,N_15897,N_15957);
nor U16163 (N_16163,N_15889,N_15940);
nand U16164 (N_16164,N_15856,N_15984);
nor U16165 (N_16165,N_15977,N_15931);
nand U16166 (N_16166,N_15988,N_15886);
and U16167 (N_16167,N_15987,N_15825);
and U16168 (N_16168,N_15914,N_15822);
xnor U16169 (N_16169,N_15928,N_15936);
nand U16170 (N_16170,N_15918,N_15898);
nor U16171 (N_16171,N_15832,N_15809);
nor U16172 (N_16172,N_15925,N_15920);
xor U16173 (N_16173,N_15922,N_15874);
nor U16174 (N_16174,N_15950,N_15969);
nand U16175 (N_16175,N_15971,N_15920);
nand U16176 (N_16176,N_15954,N_15816);
nand U16177 (N_16177,N_15979,N_15985);
nand U16178 (N_16178,N_15966,N_15813);
nor U16179 (N_16179,N_15944,N_15975);
nor U16180 (N_16180,N_15960,N_15866);
or U16181 (N_16181,N_15903,N_15928);
nand U16182 (N_16182,N_15854,N_15924);
xnor U16183 (N_16183,N_15831,N_15958);
xor U16184 (N_16184,N_15988,N_15971);
or U16185 (N_16185,N_15957,N_15886);
xor U16186 (N_16186,N_15982,N_15891);
and U16187 (N_16187,N_15827,N_15824);
nand U16188 (N_16188,N_15978,N_15846);
and U16189 (N_16189,N_15998,N_15963);
nand U16190 (N_16190,N_15999,N_15939);
xnor U16191 (N_16191,N_15989,N_15811);
xor U16192 (N_16192,N_15825,N_15980);
and U16193 (N_16193,N_15942,N_15801);
xor U16194 (N_16194,N_15816,N_15981);
nor U16195 (N_16195,N_15871,N_15927);
and U16196 (N_16196,N_15923,N_15825);
and U16197 (N_16197,N_15839,N_15879);
nand U16198 (N_16198,N_15886,N_15880);
nor U16199 (N_16199,N_15869,N_15919);
nand U16200 (N_16200,N_16194,N_16009);
nor U16201 (N_16201,N_16121,N_16115);
xor U16202 (N_16202,N_16178,N_16183);
and U16203 (N_16203,N_16109,N_16119);
xor U16204 (N_16204,N_16186,N_16047);
or U16205 (N_16205,N_16006,N_16122);
nor U16206 (N_16206,N_16001,N_16058);
nand U16207 (N_16207,N_16083,N_16181);
nor U16208 (N_16208,N_16180,N_16104);
and U16209 (N_16209,N_16024,N_16196);
nor U16210 (N_16210,N_16184,N_16116);
nand U16211 (N_16211,N_16039,N_16074);
and U16212 (N_16212,N_16100,N_16051);
and U16213 (N_16213,N_16018,N_16099);
or U16214 (N_16214,N_16152,N_16075);
xnor U16215 (N_16215,N_16089,N_16002);
and U16216 (N_16216,N_16195,N_16064);
xnor U16217 (N_16217,N_16090,N_16069);
xor U16218 (N_16218,N_16163,N_16003);
nand U16219 (N_16219,N_16017,N_16060);
nand U16220 (N_16220,N_16054,N_16188);
xor U16221 (N_16221,N_16052,N_16143);
and U16222 (N_16222,N_16120,N_16037);
xor U16223 (N_16223,N_16045,N_16136);
and U16224 (N_16224,N_16103,N_16125);
and U16225 (N_16225,N_16050,N_16063);
xnor U16226 (N_16226,N_16000,N_16016);
nand U16227 (N_16227,N_16112,N_16161);
xor U16228 (N_16228,N_16179,N_16044);
and U16229 (N_16229,N_16030,N_16142);
nor U16230 (N_16230,N_16148,N_16111);
nor U16231 (N_16231,N_16156,N_16019);
nand U16232 (N_16232,N_16010,N_16146);
nand U16233 (N_16233,N_16034,N_16190);
nand U16234 (N_16234,N_16081,N_16055);
and U16235 (N_16235,N_16154,N_16134);
nand U16236 (N_16236,N_16185,N_16098);
nor U16237 (N_16237,N_16021,N_16086);
and U16238 (N_16238,N_16084,N_16038);
nand U16239 (N_16239,N_16110,N_16144);
or U16240 (N_16240,N_16182,N_16068);
or U16241 (N_16241,N_16166,N_16062);
nand U16242 (N_16242,N_16151,N_16013);
nand U16243 (N_16243,N_16005,N_16071);
xnor U16244 (N_16244,N_16102,N_16139);
or U16245 (N_16245,N_16087,N_16096);
or U16246 (N_16246,N_16026,N_16076);
nand U16247 (N_16247,N_16041,N_16197);
and U16248 (N_16248,N_16168,N_16118);
nor U16249 (N_16249,N_16042,N_16135);
and U16250 (N_16250,N_16130,N_16191);
and U16251 (N_16251,N_16059,N_16127);
nor U16252 (N_16252,N_16169,N_16080);
nor U16253 (N_16253,N_16117,N_16105);
or U16254 (N_16254,N_16023,N_16175);
nor U16255 (N_16255,N_16049,N_16078);
nand U16256 (N_16256,N_16028,N_16061);
nor U16257 (N_16257,N_16198,N_16124);
nor U16258 (N_16258,N_16020,N_16160);
xnor U16259 (N_16259,N_16177,N_16046);
nand U16260 (N_16260,N_16048,N_16174);
or U16261 (N_16261,N_16145,N_16070);
nor U16262 (N_16262,N_16065,N_16132);
or U16263 (N_16263,N_16072,N_16097);
nor U16264 (N_16264,N_16040,N_16192);
and U16265 (N_16265,N_16033,N_16140);
nand U16266 (N_16266,N_16157,N_16101);
xor U16267 (N_16267,N_16106,N_16007);
xor U16268 (N_16268,N_16082,N_16189);
or U16269 (N_16269,N_16137,N_16027);
nor U16270 (N_16270,N_16176,N_16053);
nor U16271 (N_16271,N_16159,N_16164);
or U16272 (N_16272,N_16141,N_16131);
nor U16273 (N_16273,N_16150,N_16129);
or U16274 (N_16274,N_16025,N_16031);
nand U16275 (N_16275,N_16155,N_16032);
nor U16276 (N_16276,N_16077,N_16107);
or U16277 (N_16277,N_16153,N_16066);
xor U16278 (N_16278,N_16158,N_16092);
or U16279 (N_16279,N_16079,N_16056);
nor U16280 (N_16280,N_16193,N_16138);
and U16281 (N_16281,N_16029,N_16187);
xnor U16282 (N_16282,N_16091,N_16057);
xnor U16283 (N_16283,N_16167,N_16015);
xor U16284 (N_16284,N_16004,N_16173);
nor U16285 (N_16285,N_16011,N_16036);
and U16286 (N_16286,N_16012,N_16093);
nand U16287 (N_16287,N_16149,N_16095);
nand U16288 (N_16288,N_16022,N_16108);
nor U16289 (N_16289,N_16171,N_16094);
or U16290 (N_16290,N_16088,N_16172);
xor U16291 (N_16291,N_16199,N_16147);
or U16292 (N_16292,N_16133,N_16014);
or U16293 (N_16293,N_16073,N_16128);
or U16294 (N_16294,N_16114,N_16170);
and U16295 (N_16295,N_16165,N_16113);
or U16296 (N_16296,N_16126,N_16043);
or U16297 (N_16297,N_16067,N_16162);
and U16298 (N_16298,N_16008,N_16035);
nor U16299 (N_16299,N_16085,N_16123);
nor U16300 (N_16300,N_16031,N_16174);
nor U16301 (N_16301,N_16094,N_16166);
nor U16302 (N_16302,N_16003,N_16120);
nor U16303 (N_16303,N_16076,N_16198);
and U16304 (N_16304,N_16103,N_16023);
nand U16305 (N_16305,N_16179,N_16074);
nand U16306 (N_16306,N_16118,N_16084);
or U16307 (N_16307,N_16080,N_16142);
nand U16308 (N_16308,N_16191,N_16119);
or U16309 (N_16309,N_16054,N_16165);
nand U16310 (N_16310,N_16178,N_16038);
and U16311 (N_16311,N_16189,N_16086);
nor U16312 (N_16312,N_16061,N_16194);
nand U16313 (N_16313,N_16110,N_16115);
nand U16314 (N_16314,N_16178,N_16165);
or U16315 (N_16315,N_16152,N_16021);
and U16316 (N_16316,N_16038,N_16134);
nand U16317 (N_16317,N_16104,N_16023);
or U16318 (N_16318,N_16006,N_16163);
nor U16319 (N_16319,N_16140,N_16004);
nand U16320 (N_16320,N_16133,N_16105);
or U16321 (N_16321,N_16170,N_16048);
nand U16322 (N_16322,N_16187,N_16110);
nand U16323 (N_16323,N_16011,N_16181);
xor U16324 (N_16324,N_16083,N_16037);
and U16325 (N_16325,N_16144,N_16102);
or U16326 (N_16326,N_16103,N_16097);
nor U16327 (N_16327,N_16071,N_16043);
or U16328 (N_16328,N_16107,N_16090);
nor U16329 (N_16329,N_16076,N_16089);
xnor U16330 (N_16330,N_16028,N_16080);
xnor U16331 (N_16331,N_16110,N_16011);
nor U16332 (N_16332,N_16015,N_16187);
nand U16333 (N_16333,N_16117,N_16123);
and U16334 (N_16334,N_16028,N_16033);
xor U16335 (N_16335,N_16143,N_16168);
and U16336 (N_16336,N_16058,N_16145);
xnor U16337 (N_16337,N_16038,N_16173);
nor U16338 (N_16338,N_16053,N_16099);
or U16339 (N_16339,N_16192,N_16064);
or U16340 (N_16340,N_16005,N_16075);
nor U16341 (N_16341,N_16074,N_16172);
or U16342 (N_16342,N_16067,N_16033);
nor U16343 (N_16343,N_16189,N_16178);
nor U16344 (N_16344,N_16030,N_16043);
nand U16345 (N_16345,N_16015,N_16073);
and U16346 (N_16346,N_16123,N_16186);
or U16347 (N_16347,N_16139,N_16170);
nor U16348 (N_16348,N_16014,N_16064);
or U16349 (N_16349,N_16011,N_16084);
nand U16350 (N_16350,N_16010,N_16049);
and U16351 (N_16351,N_16142,N_16090);
nor U16352 (N_16352,N_16132,N_16174);
nor U16353 (N_16353,N_16194,N_16130);
or U16354 (N_16354,N_16026,N_16063);
nand U16355 (N_16355,N_16095,N_16062);
nor U16356 (N_16356,N_16068,N_16087);
nor U16357 (N_16357,N_16134,N_16064);
and U16358 (N_16358,N_16145,N_16108);
and U16359 (N_16359,N_16006,N_16051);
nor U16360 (N_16360,N_16061,N_16009);
xor U16361 (N_16361,N_16010,N_16020);
or U16362 (N_16362,N_16079,N_16142);
or U16363 (N_16363,N_16095,N_16132);
and U16364 (N_16364,N_16142,N_16055);
nor U16365 (N_16365,N_16030,N_16193);
or U16366 (N_16366,N_16052,N_16151);
nor U16367 (N_16367,N_16167,N_16121);
and U16368 (N_16368,N_16168,N_16026);
nor U16369 (N_16369,N_16099,N_16019);
and U16370 (N_16370,N_16071,N_16022);
xor U16371 (N_16371,N_16036,N_16034);
xor U16372 (N_16372,N_16082,N_16147);
and U16373 (N_16373,N_16014,N_16015);
and U16374 (N_16374,N_16114,N_16172);
and U16375 (N_16375,N_16157,N_16119);
xnor U16376 (N_16376,N_16178,N_16023);
and U16377 (N_16377,N_16021,N_16147);
nor U16378 (N_16378,N_16167,N_16087);
nor U16379 (N_16379,N_16130,N_16095);
and U16380 (N_16380,N_16199,N_16138);
and U16381 (N_16381,N_16109,N_16116);
nand U16382 (N_16382,N_16035,N_16055);
nand U16383 (N_16383,N_16022,N_16114);
or U16384 (N_16384,N_16003,N_16191);
xnor U16385 (N_16385,N_16049,N_16001);
xor U16386 (N_16386,N_16066,N_16191);
nor U16387 (N_16387,N_16014,N_16191);
xnor U16388 (N_16388,N_16005,N_16095);
nand U16389 (N_16389,N_16038,N_16050);
nor U16390 (N_16390,N_16165,N_16089);
nand U16391 (N_16391,N_16098,N_16033);
nor U16392 (N_16392,N_16160,N_16184);
xnor U16393 (N_16393,N_16199,N_16148);
nor U16394 (N_16394,N_16074,N_16147);
nand U16395 (N_16395,N_16094,N_16191);
nor U16396 (N_16396,N_16008,N_16067);
nand U16397 (N_16397,N_16048,N_16087);
or U16398 (N_16398,N_16008,N_16144);
nand U16399 (N_16399,N_16197,N_16100);
nand U16400 (N_16400,N_16339,N_16379);
or U16401 (N_16401,N_16356,N_16215);
xnor U16402 (N_16402,N_16207,N_16280);
or U16403 (N_16403,N_16206,N_16292);
nand U16404 (N_16404,N_16313,N_16335);
or U16405 (N_16405,N_16380,N_16390);
and U16406 (N_16406,N_16258,N_16216);
nand U16407 (N_16407,N_16349,N_16371);
and U16408 (N_16408,N_16366,N_16267);
nor U16409 (N_16409,N_16359,N_16248);
or U16410 (N_16410,N_16393,N_16361);
nor U16411 (N_16411,N_16365,N_16214);
nor U16412 (N_16412,N_16249,N_16245);
and U16413 (N_16413,N_16381,N_16370);
and U16414 (N_16414,N_16257,N_16293);
or U16415 (N_16415,N_16364,N_16276);
nor U16416 (N_16416,N_16277,N_16347);
and U16417 (N_16417,N_16259,N_16325);
and U16418 (N_16418,N_16221,N_16240);
and U16419 (N_16419,N_16340,N_16373);
or U16420 (N_16420,N_16243,N_16352);
nand U16421 (N_16421,N_16296,N_16360);
and U16422 (N_16422,N_16387,N_16272);
and U16423 (N_16423,N_16279,N_16253);
xor U16424 (N_16424,N_16354,N_16374);
xnor U16425 (N_16425,N_16266,N_16274);
nand U16426 (N_16426,N_16200,N_16388);
nor U16427 (N_16427,N_16326,N_16319);
and U16428 (N_16428,N_16315,N_16254);
and U16429 (N_16429,N_16369,N_16289);
nor U16430 (N_16430,N_16210,N_16362);
nand U16431 (N_16431,N_16343,N_16247);
or U16432 (N_16432,N_16208,N_16353);
xnor U16433 (N_16433,N_16383,N_16263);
xor U16434 (N_16434,N_16386,N_16202);
nor U16435 (N_16435,N_16384,N_16331);
or U16436 (N_16436,N_16282,N_16290);
nand U16437 (N_16437,N_16382,N_16376);
or U16438 (N_16438,N_16234,N_16281);
and U16439 (N_16439,N_16226,N_16273);
xnor U16440 (N_16440,N_16291,N_16268);
or U16441 (N_16441,N_16278,N_16399);
nor U16442 (N_16442,N_16322,N_16348);
nor U16443 (N_16443,N_16261,N_16218);
xnor U16444 (N_16444,N_16396,N_16222);
nor U16445 (N_16445,N_16203,N_16389);
or U16446 (N_16446,N_16333,N_16311);
and U16447 (N_16447,N_16205,N_16330);
and U16448 (N_16448,N_16264,N_16262);
nor U16449 (N_16449,N_16255,N_16246);
nand U16450 (N_16450,N_16213,N_16233);
nor U16451 (N_16451,N_16204,N_16355);
nand U16452 (N_16452,N_16334,N_16227);
xnor U16453 (N_16453,N_16299,N_16239);
and U16454 (N_16454,N_16312,N_16219);
nor U16455 (N_16455,N_16209,N_16305);
nor U16456 (N_16456,N_16341,N_16269);
xor U16457 (N_16457,N_16302,N_16345);
nand U16458 (N_16458,N_16316,N_16397);
xor U16459 (N_16459,N_16217,N_16375);
xor U16460 (N_16460,N_16327,N_16350);
nand U16461 (N_16461,N_16323,N_16351);
and U16462 (N_16462,N_16271,N_16309);
and U16463 (N_16463,N_16270,N_16320);
nor U16464 (N_16464,N_16244,N_16363);
xor U16465 (N_16465,N_16285,N_16328);
nand U16466 (N_16466,N_16256,N_16314);
or U16467 (N_16467,N_16306,N_16237);
and U16468 (N_16468,N_16336,N_16225);
xor U16469 (N_16469,N_16298,N_16236);
nand U16470 (N_16470,N_16391,N_16392);
or U16471 (N_16471,N_16308,N_16287);
xor U16472 (N_16472,N_16346,N_16385);
xor U16473 (N_16473,N_16223,N_16304);
or U16474 (N_16474,N_16220,N_16295);
nand U16475 (N_16475,N_16232,N_16238);
nor U16476 (N_16476,N_16394,N_16342);
nor U16477 (N_16477,N_16395,N_16301);
nor U16478 (N_16478,N_16303,N_16211);
and U16479 (N_16479,N_16321,N_16251);
nor U16480 (N_16480,N_16338,N_16329);
or U16481 (N_16481,N_16297,N_16230);
and U16482 (N_16482,N_16284,N_16286);
xnor U16483 (N_16483,N_16224,N_16241);
and U16484 (N_16484,N_16310,N_16212);
nand U16485 (N_16485,N_16260,N_16378);
nor U16486 (N_16486,N_16344,N_16288);
and U16487 (N_16487,N_16337,N_16372);
and U16488 (N_16488,N_16324,N_16307);
nor U16489 (N_16489,N_16252,N_16332);
nand U16490 (N_16490,N_16229,N_16300);
and U16491 (N_16491,N_16294,N_16398);
or U16492 (N_16492,N_16368,N_16242);
or U16493 (N_16493,N_16228,N_16357);
or U16494 (N_16494,N_16250,N_16317);
and U16495 (N_16495,N_16367,N_16231);
or U16496 (N_16496,N_16318,N_16275);
xor U16497 (N_16497,N_16283,N_16358);
or U16498 (N_16498,N_16235,N_16377);
or U16499 (N_16499,N_16201,N_16265);
or U16500 (N_16500,N_16257,N_16240);
nor U16501 (N_16501,N_16249,N_16205);
or U16502 (N_16502,N_16237,N_16323);
nand U16503 (N_16503,N_16384,N_16311);
or U16504 (N_16504,N_16308,N_16284);
nor U16505 (N_16505,N_16327,N_16205);
and U16506 (N_16506,N_16367,N_16301);
nand U16507 (N_16507,N_16204,N_16340);
xnor U16508 (N_16508,N_16263,N_16295);
nand U16509 (N_16509,N_16240,N_16293);
or U16510 (N_16510,N_16322,N_16269);
nor U16511 (N_16511,N_16372,N_16247);
nor U16512 (N_16512,N_16373,N_16216);
nor U16513 (N_16513,N_16322,N_16264);
xor U16514 (N_16514,N_16249,N_16353);
and U16515 (N_16515,N_16389,N_16313);
xnor U16516 (N_16516,N_16388,N_16313);
or U16517 (N_16517,N_16349,N_16389);
and U16518 (N_16518,N_16297,N_16286);
or U16519 (N_16519,N_16302,N_16347);
xnor U16520 (N_16520,N_16227,N_16347);
xor U16521 (N_16521,N_16379,N_16214);
xor U16522 (N_16522,N_16380,N_16330);
nor U16523 (N_16523,N_16352,N_16231);
nor U16524 (N_16524,N_16307,N_16342);
nor U16525 (N_16525,N_16303,N_16252);
and U16526 (N_16526,N_16233,N_16206);
nor U16527 (N_16527,N_16396,N_16261);
nor U16528 (N_16528,N_16272,N_16249);
xnor U16529 (N_16529,N_16232,N_16359);
xor U16530 (N_16530,N_16332,N_16233);
nor U16531 (N_16531,N_16230,N_16396);
xor U16532 (N_16532,N_16292,N_16283);
xor U16533 (N_16533,N_16375,N_16374);
nor U16534 (N_16534,N_16270,N_16279);
nor U16535 (N_16535,N_16203,N_16335);
and U16536 (N_16536,N_16287,N_16385);
nor U16537 (N_16537,N_16300,N_16358);
xor U16538 (N_16538,N_16235,N_16273);
or U16539 (N_16539,N_16295,N_16330);
nor U16540 (N_16540,N_16224,N_16335);
nor U16541 (N_16541,N_16260,N_16344);
xnor U16542 (N_16542,N_16342,N_16312);
xnor U16543 (N_16543,N_16334,N_16261);
and U16544 (N_16544,N_16362,N_16207);
and U16545 (N_16545,N_16229,N_16255);
nand U16546 (N_16546,N_16303,N_16379);
or U16547 (N_16547,N_16270,N_16356);
xnor U16548 (N_16548,N_16349,N_16255);
or U16549 (N_16549,N_16233,N_16237);
xor U16550 (N_16550,N_16238,N_16281);
xnor U16551 (N_16551,N_16200,N_16289);
xnor U16552 (N_16552,N_16216,N_16280);
and U16553 (N_16553,N_16386,N_16336);
nand U16554 (N_16554,N_16260,N_16367);
nor U16555 (N_16555,N_16223,N_16204);
xor U16556 (N_16556,N_16255,N_16336);
nand U16557 (N_16557,N_16372,N_16270);
or U16558 (N_16558,N_16331,N_16235);
or U16559 (N_16559,N_16360,N_16331);
and U16560 (N_16560,N_16387,N_16222);
nand U16561 (N_16561,N_16288,N_16245);
nand U16562 (N_16562,N_16242,N_16207);
or U16563 (N_16563,N_16269,N_16310);
nor U16564 (N_16564,N_16394,N_16237);
nor U16565 (N_16565,N_16334,N_16338);
xnor U16566 (N_16566,N_16385,N_16395);
nand U16567 (N_16567,N_16314,N_16344);
xor U16568 (N_16568,N_16346,N_16392);
or U16569 (N_16569,N_16265,N_16320);
or U16570 (N_16570,N_16332,N_16264);
or U16571 (N_16571,N_16215,N_16228);
and U16572 (N_16572,N_16345,N_16281);
nor U16573 (N_16573,N_16335,N_16368);
nand U16574 (N_16574,N_16258,N_16243);
and U16575 (N_16575,N_16326,N_16307);
nor U16576 (N_16576,N_16241,N_16351);
xor U16577 (N_16577,N_16225,N_16245);
and U16578 (N_16578,N_16224,N_16271);
nor U16579 (N_16579,N_16349,N_16348);
or U16580 (N_16580,N_16332,N_16347);
xor U16581 (N_16581,N_16239,N_16348);
or U16582 (N_16582,N_16374,N_16357);
or U16583 (N_16583,N_16353,N_16246);
nor U16584 (N_16584,N_16213,N_16259);
xnor U16585 (N_16585,N_16267,N_16368);
or U16586 (N_16586,N_16265,N_16328);
nand U16587 (N_16587,N_16259,N_16267);
xor U16588 (N_16588,N_16353,N_16334);
and U16589 (N_16589,N_16299,N_16200);
nor U16590 (N_16590,N_16292,N_16362);
or U16591 (N_16591,N_16354,N_16300);
nand U16592 (N_16592,N_16303,N_16220);
or U16593 (N_16593,N_16203,N_16223);
nor U16594 (N_16594,N_16386,N_16395);
nand U16595 (N_16595,N_16396,N_16348);
nand U16596 (N_16596,N_16220,N_16255);
nand U16597 (N_16597,N_16214,N_16373);
nand U16598 (N_16598,N_16272,N_16332);
and U16599 (N_16599,N_16371,N_16364);
nor U16600 (N_16600,N_16504,N_16471);
nor U16601 (N_16601,N_16540,N_16503);
nand U16602 (N_16602,N_16549,N_16455);
nand U16603 (N_16603,N_16562,N_16501);
nand U16604 (N_16604,N_16598,N_16533);
nor U16605 (N_16605,N_16415,N_16401);
or U16606 (N_16606,N_16443,N_16580);
or U16607 (N_16607,N_16595,N_16457);
nor U16608 (N_16608,N_16507,N_16553);
and U16609 (N_16609,N_16536,N_16441);
nor U16610 (N_16610,N_16557,N_16546);
nor U16611 (N_16611,N_16468,N_16506);
and U16612 (N_16612,N_16541,N_16558);
nor U16613 (N_16613,N_16411,N_16577);
and U16614 (N_16614,N_16593,N_16565);
nand U16615 (N_16615,N_16519,N_16538);
nand U16616 (N_16616,N_16413,N_16402);
or U16617 (N_16617,N_16516,N_16500);
or U16618 (N_16618,N_16496,N_16494);
nand U16619 (N_16619,N_16465,N_16452);
and U16620 (N_16620,N_16573,N_16450);
nor U16621 (N_16621,N_16493,N_16583);
and U16622 (N_16622,N_16424,N_16480);
or U16623 (N_16623,N_16582,N_16545);
and U16624 (N_16624,N_16425,N_16466);
or U16625 (N_16625,N_16490,N_16431);
xor U16626 (N_16626,N_16547,N_16429);
or U16627 (N_16627,N_16551,N_16556);
nor U16628 (N_16628,N_16529,N_16400);
nor U16629 (N_16629,N_16570,N_16454);
or U16630 (N_16630,N_16485,N_16448);
nand U16631 (N_16631,N_16491,N_16515);
nor U16632 (N_16632,N_16572,N_16505);
and U16633 (N_16633,N_16563,N_16403);
nor U16634 (N_16634,N_16476,N_16592);
nand U16635 (N_16635,N_16520,N_16484);
or U16636 (N_16636,N_16474,N_16467);
xor U16637 (N_16637,N_16559,N_16550);
and U16638 (N_16638,N_16451,N_16408);
nand U16639 (N_16639,N_16445,N_16409);
and U16640 (N_16640,N_16492,N_16463);
or U16641 (N_16641,N_16428,N_16596);
and U16642 (N_16642,N_16555,N_16571);
or U16643 (N_16643,N_16446,N_16487);
nand U16644 (N_16644,N_16433,N_16420);
nor U16645 (N_16645,N_16512,N_16535);
nand U16646 (N_16646,N_16578,N_16499);
nand U16647 (N_16647,N_16508,N_16498);
or U16648 (N_16648,N_16513,N_16434);
or U16649 (N_16649,N_16502,N_16543);
xnor U16650 (N_16650,N_16440,N_16437);
nand U16651 (N_16651,N_16436,N_16597);
nor U16652 (N_16652,N_16404,N_16586);
xor U16653 (N_16653,N_16554,N_16406);
nor U16654 (N_16654,N_16456,N_16472);
nor U16655 (N_16655,N_16528,N_16599);
or U16656 (N_16656,N_16418,N_16552);
or U16657 (N_16657,N_16589,N_16511);
xnor U16658 (N_16658,N_16534,N_16438);
and U16659 (N_16659,N_16458,N_16587);
nor U16660 (N_16660,N_16489,N_16444);
or U16661 (N_16661,N_16419,N_16426);
and U16662 (N_16662,N_16421,N_16473);
nand U16663 (N_16663,N_16405,N_16477);
and U16664 (N_16664,N_16588,N_16497);
nand U16665 (N_16665,N_16407,N_16575);
and U16666 (N_16666,N_16481,N_16525);
xor U16667 (N_16667,N_16470,N_16584);
xor U16668 (N_16668,N_16560,N_16532);
xnor U16669 (N_16669,N_16469,N_16461);
or U16670 (N_16670,N_16561,N_16585);
xnor U16671 (N_16671,N_16591,N_16464);
nor U16672 (N_16672,N_16518,N_16539);
nor U16673 (N_16673,N_16422,N_16488);
or U16674 (N_16674,N_16521,N_16432);
and U16675 (N_16675,N_16514,N_16447);
xnor U16676 (N_16676,N_16568,N_16412);
nand U16677 (N_16677,N_16530,N_16486);
xor U16678 (N_16678,N_16542,N_16537);
and U16679 (N_16679,N_16459,N_16462);
nand U16680 (N_16680,N_16449,N_16564);
nand U16681 (N_16681,N_16569,N_16423);
nor U16682 (N_16682,N_16517,N_16522);
and U16683 (N_16683,N_16509,N_16590);
xor U16684 (N_16684,N_16581,N_16430);
nand U16685 (N_16685,N_16524,N_16483);
nand U16686 (N_16686,N_16427,N_16576);
xor U16687 (N_16687,N_16478,N_16579);
nand U16688 (N_16688,N_16416,N_16567);
or U16689 (N_16689,N_16479,N_16526);
nand U16690 (N_16690,N_16482,N_16531);
or U16691 (N_16691,N_16594,N_16574);
and U16692 (N_16692,N_16435,N_16475);
nand U16693 (N_16693,N_16544,N_16439);
nand U16694 (N_16694,N_16523,N_16527);
nand U16695 (N_16695,N_16495,N_16442);
nor U16696 (N_16696,N_16548,N_16566);
or U16697 (N_16697,N_16414,N_16510);
or U16698 (N_16698,N_16460,N_16410);
xor U16699 (N_16699,N_16417,N_16453);
xnor U16700 (N_16700,N_16586,N_16435);
nand U16701 (N_16701,N_16403,N_16530);
nand U16702 (N_16702,N_16476,N_16569);
nor U16703 (N_16703,N_16464,N_16474);
and U16704 (N_16704,N_16420,N_16481);
or U16705 (N_16705,N_16523,N_16599);
nand U16706 (N_16706,N_16494,N_16566);
and U16707 (N_16707,N_16546,N_16424);
and U16708 (N_16708,N_16445,N_16491);
xor U16709 (N_16709,N_16518,N_16501);
xor U16710 (N_16710,N_16591,N_16546);
or U16711 (N_16711,N_16403,N_16448);
and U16712 (N_16712,N_16495,N_16464);
nor U16713 (N_16713,N_16570,N_16561);
nand U16714 (N_16714,N_16497,N_16592);
xor U16715 (N_16715,N_16425,N_16515);
and U16716 (N_16716,N_16578,N_16551);
nand U16717 (N_16717,N_16576,N_16459);
xnor U16718 (N_16718,N_16577,N_16551);
or U16719 (N_16719,N_16462,N_16578);
xor U16720 (N_16720,N_16480,N_16478);
and U16721 (N_16721,N_16558,N_16572);
nor U16722 (N_16722,N_16587,N_16472);
or U16723 (N_16723,N_16544,N_16456);
nand U16724 (N_16724,N_16549,N_16470);
nor U16725 (N_16725,N_16503,N_16418);
nor U16726 (N_16726,N_16575,N_16557);
xnor U16727 (N_16727,N_16506,N_16532);
or U16728 (N_16728,N_16433,N_16411);
nor U16729 (N_16729,N_16480,N_16408);
nand U16730 (N_16730,N_16539,N_16525);
and U16731 (N_16731,N_16594,N_16456);
xor U16732 (N_16732,N_16420,N_16506);
or U16733 (N_16733,N_16570,N_16586);
nand U16734 (N_16734,N_16478,N_16565);
nand U16735 (N_16735,N_16495,N_16469);
and U16736 (N_16736,N_16590,N_16440);
nand U16737 (N_16737,N_16417,N_16455);
xor U16738 (N_16738,N_16446,N_16498);
and U16739 (N_16739,N_16519,N_16417);
and U16740 (N_16740,N_16443,N_16456);
and U16741 (N_16741,N_16418,N_16464);
or U16742 (N_16742,N_16587,N_16401);
nand U16743 (N_16743,N_16513,N_16529);
nand U16744 (N_16744,N_16574,N_16513);
or U16745 (N_16745,N_16493,N_16454);
xor U16746 (N_16746,N_16557,N_16539);
and U16747 (N_16747,N_16527,N_16531);
nand U16748 (N_16748,N_16455,N_16571);
or U16749 (N_16749,N_16541,N_16441);
xor U16750 (N_16750,N_16599,N_16492);
xor U16751 (N_16751,N_16489,N_16590);
or U16752 (N_16752,N_16431,N_16413);
nand U16753 (N_16753,N_16458,N_16552);
or U16754 (N_16754,N_16594,N_16476);
and U16755 (N_16755,N_16471,N_16545);
and U16756 (N_16756,N_16490,N_16410);
or U16757 (N_16757,N_16541,N_16450);
and U16758 (N_16758,N_16571,N_16531);
nand U16759 (N_16759,N_16562,N_16495);
xnor U16760 (N_16760,N_16584,N_16461);
xor U16761 (N_16761,N_16519,N_16562);
xnor U16762 (N_16762,N_16492,N_16475);
nor U16763 (N_16763,N_16424,N_16449);
nor U16764 (N_16764,N_16480,N_16583);
or U16765 (N_16765,N_16421,N_16523);
or U16766 (N_16766,N_16429,N_16458);
nor U16767 (N_16767,N_16425,N_16428);
nor U16768 (N_16768,N_16438,N_16568);
and U16769 (N_16769,N_16522,N_16508);
nand U16770 (N_16770,N_16589,N_16506);
nor U16771 (N_16771,N_16435,N_16457);
nor U16772 (N_16772,N_16572,N_16541);
and U16773 (N_16773,N_16569,N_16402);
nand U16774 (N_16774,N_16465,N_16425);
xor U16775 (N_16775,N_16551,N_16520);
and U16776 (N_16776,N_16524,N_16511);
nor U16777 (N_16777,N_16442,N_16505);
or U16778 (N_16778,N_16506,N_16565);
or U16779 (N_16779,N_16447,N_16433);
nor U16780 (N_16780,N_16490,N_16411);
nor U16781 (N_16781,N_16483,N_16511);
xnor U16782 (N_16782,N_16441,N_16403);
nor U16783 (N_16783,N_16548,N_16511);
nor U16784 (N_16784,N_16593,N_16503);
nand U16785 (N_16785,N_16533,N_16512);
xnor U16786 (N_16786,N_16533,N_16547);
nor U16787 (N_16787,N_16595,N_16592);
or U16788 (N_16788,N_16509,N_16411);
or U16789 (N_16789,N_16516,N_16488);
xor U16790 (N_16790,N_16419,N_16472);
or U16791 (N_16791,N_16493,N_16424);
nor U16792 (N_16792,N_16573,N_16497);
or U16793 (N_16793,N_16508,N_16572);
xor U16794 (N_16794,N_16546,N_16495);
and U16795 (N_16795,N_16469,N_16493);
and U16796 (N_16796,N_16502,N_16503);
nor U16797 (N_16797,N_16404,N_16421);
xor U16798 (N_16798,N_16439,N_16450);
nor U16799 (N_16799,N_16518,N_16570);
nor U16800 (N_16800,N_16781,N_16789);
xnor U16801 (N_16801,N_16744,N_16757);
and U16802 (N_16802,N_16649,N_16774);
or U16803 (N_16803,N_16640,N_16720);
xnor U16804 (N_16804,N_16743,N_16714);
nor U16805 (N_16805,N_16642,N_16735);
and U16806 (N_16806,N_16636,N_16681);
nor U16807 (N_16807,N_16673,N_16776);
or U16808 (N_16808,N_16603,N_16739);
or U16809 (N_16809,N_16783,N_16741);
xnor U16810 (N_16810,N_16758,N_16660);
nand U16811 (N_16811,N_16613,N_16703);
nand U16812 (N_16812,N_16699,N_16606);
nand U16813 (N_16813,N_16676,N_16794);
xor U16814 (N_16814,N_16750,N_16644);
nor U16815 (N_16815,N_16679,N_16621);
or U16816 (N_16816,N_16659,N_16709);
nand U16817 (N_16817,N_16713,N_16656);
nand U16818 (N_16818,N_16650,N_16790);
nand U16819 (N_16819,N_16648,N_16638);
nand U16820 (N_16820,N_16753,N_16622);
nand U16821 (N_16821,N_16682,N_16764);
nand U16822 (N_16822,N_16772,N_16782);
nor U16823 (N_16823,N_16605,N_16675);
nand U16824 (N_16824,N_16639,N_16761);
nor U16825 (N_16825,N_16604,N_16726);
or U16826 (N_16826,N_16686,N_16601);
nand U16827 (N_16827,N_16722,N_16786);
or U16828 (N_16828,N_16626,N_16632);
or U16829 (N_16829,N_16637,N_16770);
nand U16830 (N_16830,N_16729,N_16748);
or U16831 (N_16831,N_16669,N_16683);
xnor U16832 (N_16832,N_16687,N_16734);
and U16833 (N_16833,N_16643,N_16738);
and U16834 (N_16834,N_16711,N_16658);
nor U16835 (N_16835,N_16795,N_16763);
and U16836 (N_16836,N_16665,N_16766);
nor U16837 (N_16837,N_16667,N_16725);
and U16838 (N_16838,N_16652,N_16704);
xor U16839 (N_16839,N_16654,N_16762);
or U16840 (N_16840,N_16773,N_16661);
nand U16841 (N_16841,N_16765,N_16629);
and U16842 (N_16842,N_16787,N_16688);
nand U16843 (N_16843,N_16662,N_16723);
nand U16844 (N_16844,N_16633,N_16731);
nor U16845 (N_16845,N_16740,N_16784);
and U16846 (N_16846,N_16747,N_16615);
nor U16847 (N_16847,N_16627,N_16727);
nor U16848 (N_16848,N_16690,N_16689);
xor U16849 (N_16849,N_16695,N_16693);
nand U16850 (N_16850,N_16717,N_16630);
xor U16851 (N_16851,N_16791,N_16691);
xnor U16852 (N_16852,N_16756,N_16760);
nor U16853 (N_16853,N_16792,N_16618);
xnor U16854 (N_16854,N_16706,N_16712);
and U16855 (N_16855,N_16692,N_16777);
and U16856 (N_16856,N_16742,N_16719);
nand U16857 (N_16857,N_16755,N_16768);
xor U16858 (N_16858,N_16678,N_16625);
nand U16859 (N_16859,N_16724,N_16628);
nand U16860 (N_16860,N_16620,N_16798);
and U16861 (N_16861,N_16796,N_16702);
and U16862 (N_16862,N_16700,N_16746);
xnor U16863 (N_16863,N_16698,N_16752);
and U16864 (N_16864,N_16732,N_16799);
and U16865 (N_16865,N_16666,N_16697);
or U16866 (N_16866,N_16672,N_16705);
and U16867 (N_16867,N_16600,N_16663);
or U16868 (N_16868,N_16611,N_16617);
nor U16869 (N_16869,N_16749,N_16635);
nand U16870 (N_16870,N_16609,N_16707);
xnor U16871 (N_16871,N_16769,N_16614);
or U16872 (N_16872,N_16653,N_16780);
xnor U16873 (N_16873,N_16701,N_16767);
nand U16874 (N_16874,N_16671,N_16771);
and U16875 (N_16875,N_16646,N_16728);
xnor U16876 (N_16876,N_16715,N_16797);
nand U16877 (N_16877,N_16694,N_16710);
xnor U16878 (N_16878,N_16616,N_16670);
nand U16879 (N_16879,N_16612,N_16608);
or U16880 (N_16880,N_16730,N_16779);
or U16881 (N_16881,N_16716,N_16775);
and U16882 (N_16882,N_16754,N_16657);
xnor U16883 (N_16883,N_16696,N_16788);
xor U16884 (N_16884,N_16685,N_16651);
or U16885 (N_16885,N_16623,N_16778);
xnor U16886 (N_16886,N_16624,N_16602);
and U16887 (N_16887,N_16793,N_16733);
and U16888 (N_16888,N_16751,N_16785);
xor U16889 (N_16889,N_16745,N_16718);
nand U16890 (N_16890,N_16674,N_16721);
xor U16891 (N_16891,N_16677,N_16607);
xnor U16892 (N_16892,N_16680,N_16736);
nor U16893 (N_16893,N_16664,N_16631);
nor U16894 (N_16894,N_16641,N_16610);
and U16895 (N_16895,N_16619,N_16634);
nor U16896 (N_16896,N_16684,N_16737);
xnor U16897 (N_16897,N_16655,N_16647);
xnor U16898 (N_16898,N_16708,N_16668);
or U16899 (N_16899,N_16759,N_16645);
and U16900 (N_16900,N_16699,N_16716);
or U16901 (N_16901,N_16662,N_16615);
or U16902 (N_16902,N_16652,N_16660);
or U16903 (N_16903,N_16728,N_16663);
xnor U16904 (N_16904,N_16796,N_16691);
nor U16905 (N_16905,N_16741,N_16620);
xor U16906 (N_16906,N_16680,N_16717);
and U16907 (N_16907,N_16728,N_16759);
or U16908 (N_16908,N_16635,N_16750);
xnor U16909 (N_16909,N_16794,N_16697);
nor U16910 (N_16910,N_16729,N_16759);
or U16911 (N_16911,N_16696,N_16647);
and U16912 (N_16912,N_16787,N_16642);
or U16913 (N_16913,N_16608,N_16611);
xnor U16914 (N_16914,N_16665,N_16715);
nor U16915 (N_16915,N_16772,N_16690);
xnor U16916 (N_16916,N_16740,N_16607);
nand U16917 (N_16917,N_16766,N_16782);
nand U16918 (N_16918,N_16778,N_16748);
nand U16919 (N_16919,N_16662,N_16621);
or U16920 (N_16920,N_16716,N_16774);
and U16921 (N_16921,N_16719,N_16780);
or U16922 (N_16922,N_16676,N_16750);
xor U16923 (N_16923,N_16604,N_16752);
xnor U16924 (N_16924,N_16699,N_16735);
and U16925 (N_16925,N_16773,N_16647);
or U16926 (N_16926,N_16796,N_16640);
nand U16927 (N_16927,N_16739,N_16650);
and U16928 (N_16928,N_16673,N_16608);
or U16929 (N_16929,N_16715,N_16709);
nand U16930 (N_16930,N_16685,N_16753);
xor U16931 (N_16931,N_16767,N_16651);
nor U16932 (N_16932,N_16684,N_16713);
and U16933 (N_16933,N_16775,N_16675);
or U16934 (N_16934,N_16795,N_16616);
nand U16935 (N_16935,N_16733,N_16682);
nor U16936 (N_16936,N_16671,N_16693);
and U16937 (N_16937,N_16764,N_16724);
nor U16938 (N_16938,N_16732,N_16618);
or U16939 (N_16939,N_16729,N_16607);
nand U16940 (N_16940,N_16601,N_16703);
or U16941 (N_16941,N_16652,N_16698);
nor U16942 (N_16942,N_16771,N_16786);
nand U16943 (N_16943,N_16770,N_16713);
or U16944 (N_16944,N_16733,N_16703);
and U16945 (N_16945,N_16748,N_16788);
nor U16946 (N_16946,N_16603,N_16785);
nand U16947 (N_16947,N_16755,N_16703);
nand U16948 (N_16948,N_16616,N_16737);
nor U16949 (N_16949,N_16776,N_16653);
or U16950 (N_16950,N_16682,N_16766);
or U16951 (N_16951,N_16603,N_16769);
xnor U16952 (N_16952,N_16702,N_16624);
and U16953 (N_16953,N_16777,N_16740);
xor U16954 (N_16954,N_16715,N_16684);
xor U16955 (N_16955,N_16682,N_16608);
nor U16956 (N_16956,N_16742,N_16617);
and U16957 (N_16957,N_16609,N_16702);
nand U16958 (N_16958,N_16651,N_16706);
nor U16959 (N_16959,N_16719,N_16705);
and U16960 (N_16960,N_16724,N_16606);
and U16961 (N_16961,N_16640,N_16681);
nand U16962 (N_16962,N_16604,N_16639);
and U16963 (N_16963,N_16785,N_16770);
xor U16964 (N_16964,N_16681,N_16784);
nand U16965 (N_16965,N_16687,N_16653);
xor U16966 (N_16966,N_16639,N_16608);
or U16967 (N_16967,N_16676,N_16607);
nor U16968 (N_16968,N_16637,N_16728);
nand U16969 (N_16969,N_16610,N_16613);
xnor U16970 (N_16970,N_16634,N_16772);
nand U16971 (N_16971,N_16768,N_16605);
xor U16972 (N_16972,N_16672,N_16739);
or U16973 (N_16973,N_16643,N_16687);
nand U16974 (N_16974,N_16759,N_16793);
nor U16975 (N_16975,N_16619,N_16772);
xnor U16976 (N_16976,N_16747,N_16768);
nor U16977 (N_16977,N_16683,N_16747);
or U16978 (N_16978,N_16635,N_16782);
and U16979 (N_16979,N_16629,N_16757);
nor U16980 (N_16980,N_16694,N_16754);
and U16981 (N_16981,N_16647,N_16774);
or U16982 (N_16982,N_16608,N_16644);
nand U16983 (N_16983,N_16737,N_16671);
or U16984 (N_16984,N_16793,N_16648);
or U16985 (N_16985,N_16628,N_16693);
or U16986 (N_16986,N_16602,N_16777);
nand U16987 (N_16987,N_16705,N_16613);
nor U16988 (N_16988,N_16642,N_16780);
nand U16989 (N_16989,N_16699,N_16639);
xor U16990 (N_16990,N_16680,N_16731);
xnor U16991 (N_16991,N_16683,N_16717);
nor U16992 (N_16992,N_16739,N_16742);
nand U16993 (N_16993,N_16659,N_16762);
or U16994 (N_16994,N_16796,N_16696);
and U16995 (N_16995,N_16606,N_16739);
xnor U16996 (N_16996,N_16621,N_16733);
nand U16997 (N_16997,N_16718,N_16679);
nand U16998 (N_16998,N_16635,N_16610);
and U16999 (N_16999,N_16751,N_16601);
xor U17000 (N_17000,N_16802,N_16803);
nand U17001 (N_17001,N_16938,N_16906);
or U17002 (N_17002,N_16879,N_16836);
or U17003 (N_17003,N_16812,N_16954);
xnor U17004 (N_17004,N_16916,N_16995);
nor U17005 (N_17005,N_16847,N_16829);
xnor U17006 (N_17006,N_16824,N_16977);
nor U17007 (N_17007,N_16868,N_16988);
xnor U17008 (N_17008,N_16861,N_16939);
nand U17009 (N_17009,N_16928,N_16865);
and U17010 (N_17010,N_16964,N_16905);
and U17011 (N_17011,N_16854,N_16986);
nand U17012 (N_17012,N_16930,N_16818);
xnor U17013 (N_17013,N_16904,N_16896);
and U17014 (N_17014,N_16892,N_16805);
nand U17015 (N_17015,N_16846,N_16858);
nor U17016 (N_17016,N_16979,N_16820);
xnor U17017 (N_17017,N_16937,N_16819);
xor U17018 (N_17018,N_16852,N_16958);
or U17019 (N_17019,N_16994,N_16929);
or U17020 (N_17020,N_16911,N_16924);
xnor U17021 (N_17021,N_16817,N_16907);
and U17022 (N_17022,N_16899,N_16869);
or U17023 (N_17023,N_16814,N_16926);
xnor U17024 (N_17024,N_16931,N_16801);
or U17025 (N_17025,N_16843,N_16970);
xor U17026 (N_17026,N_16932,N_16804);
or U17027 (N_17027,N_16908,N_16889);
xnor U17028 (N_17028,N_16910,N_16902);
and U17029 (N_17029,N_16921,N_16975);
nor U17030 (N_17030,N_16841,N_16893);
and U17031 (N_17031,N_16981,N_16948);
and U17032 (N_17032,N_16933,N_16971);
or U17033 (N_17033,N_16987,N_16955);
nand U17034 (N_17034,N_16885,N_16856);
or U17035 (N_17035,N_16807,N_16880);
and U17036 (N_17036,N_16922,N_16800);
or U17037 (N_17037,N_16822,N_16844);
and U17038 (N_17038,N_16864,N_16888);
nor U17039 (N_17039,N_16942,N_16870);
xnor U17040 (N_17040,N_16877,N_16881);
nor U17041 (N_17041,N_16997,N_16855);
xor U17042 (N_17042,N_16830,N_16874);
nor U17043 (N_17043,N_16973,N_16990);
xor U17044 (N_17044,N_16991,N_16873);
nor U17045 (N_17045,N_16913,N_16900);
xor U17046 (N_17046,N_16941,N_16835);
nor U17047 (N_17047,N_16884,N_16978);
xor U17048 (N_17048,N_16882,N_16837);
or U17049 (N_17049,N_16898,N_16834);
nand U17050 (N_17050,N_16967,N_16860);
nor U17051 (N_17051,N_16912,N_16949);
or U17052 (N_17052,N_16821,N_16920);
and U17053 (N_17053,N_16887,N_16963);
and U17054 (N_17054,N_16998,N_16883);
nor U17055 (N_17055,N_16940,N_16823);
or U17056 (N_17056,N_16833,N_16903);
nand U17057 (N_17057,N_16917,N_16828);
and U17058 (N_17058,N_16989,N_16809);
nor U17059 (N_17059,N_16857,N_16816);
and U17060 (N_17060,N_16863,N_16952);
and U17061 (N_17061,N_16859,N_16943);
and U17062 (N_17062,N_16845,N_16985);
and U17063 (N_17063,N_16825,N_16831);
xor U17064 (N_17064,N_16983,N_16919);
xor U17065 (N_17065,N_16935,N_16810);
nand U17066 (N_17066,N_16872,N_16951);
or U17067 (N_17067,N_16875,N_16984);
and U17068 (N_17068,N_16936,N_16853);
or U17069 (N_17069,N_16815,N_16909);
and U17070 (N_17070,N_16961,N_16840);
and U17071 (N_17071,N_16953,N_16862);
nand U17072 (N_17072,N_16976,N_16945);
xnor U17073 (N_17073,N_16886,N_16827);
or U17074 (N_17074,N_16915,N_16966);
nand U17075 (N_17075,N_16832,N_16982);
nor U17076 (N_17076,N_16927,N_16842);
or U17077 (N_17077,N_16934,N_16851);
nor U17078 (N_17078,N_16878,N_16866);
or U17079 (N_17079,N_16867,N_16996);
nor U17080 (N_17080,N_16999,N_16923);
xnor U17081 (N_17081,N_16811,N_16813);
or U17082 (N_17082,N_16925,N_16947);
and U17083 (N_17083,N_16897,N_16993);
xnor U17084 (N_17084,N_16969,N_16959);
or U17085 (N_17085,N_16871,N_16950);
and U17086 (N_17086,N_16944,N_16808);
or U17087 (N_17087,N_16806,N_16876);
nand U17088 (N_17088,N_16901,N_16850);
nor U17089 (N_17089,N_16839,N_16956);
xor U17090 (N_17090,N_16914,N_16965);
or U17091 (N_17091,N_16895,N_16974);
nand U17092 (N_17092,N_16946,N_16957);
nor U17093 (N_17093,N_16894,N_16972);
and U17094 (N_17094,N_16890,N_16918);
xnor U17095 (N_17095,N_16980,N_16960);
xor U17096 (N_17096,N_16838,N_16848);
or U17097 (N_17097,N_16826,N_16968);
nor U17098 (N_17098,N_16891,N_16849);
nor U17099 (N_17099,N_16992,N_16962);
or U17100 (N_17100,N_16906,N_16963);
xor U17101 (N_17101,N_16940,N_16815);
and U17102 (N_17102,N_16973,N_16832);
and U17103 (N_17103,N_16999,N_16869);
nand U17104 (N_17104,N_16888,N_16875);
or U17105 (N_17105,N_16857,N_16900);
nand U17106 (N_17106,N_16820,N_16948);
xor U17107 (N_17107,N_16987,N_16889);
xor U17108 (N_17108,N_16983,N_16998);
xor U17109 (N_17109,N_16975,N_16969);
or U17110 (N_17110,N_16830,N_16979);
nand U17111 (N_17111,N_16933,N_16958);
xor U17112 (N_17112,N_16882,N_16886);
nor U17113 (N_17113,N_16992,N_16966);
xor U17114 (N_17114,N_16806,N_16984);
nor U17115 (N_17115,N_16865,N_16988);
nor U17116 (N_17116,N_16983,N_16860);
nor U17117 (N_17117,N_16800,N_16875);
xor U17118 (N_17118,N_16952,N_16808);
nand U17119 (N_17119,N_16987,N_16917);
nand U17120 (N_17120,N_16881,N_16919);
or U17121 (N_17121,N_16938,N_16847);
or U17122 (N_17122,N_16839,N_16884);
nand U17123 (N_17123,N_16929,N_16920);
or U17124 (N_17124,N_16829,N_16932);
xor U17125 (N_17125,N_16863,N_16879);
nand U17126 (N_17126,N_16889,N_16811);
and U17127 (N_17127,N_16974,N_16819);
nand U17128 (N_17128,N_16848,N_16939);
nand U17129 (N_17129,N_16889,N_16838);
or U17130 (N_17130,N_16938,N_16861);
nor U17131 (N_17131,N_16885,N_16970);
xnor U17132 (N_17132,N_16948,N_16804);
or U17133 (N_17133,N_16883,N_16806);
and U17134 (N_17134,N_16945,N_16947);
or U17135 (N_17135,N_16905,N_16820);
nand U17136 (N_17136,N_16930,N_16868);
nor U17137 (N_17137,N_16813,N_16980);
nor U17138 (N_17138,N_16973,N_16989);
and U17139 (N_17139,N_16807,N_16893);
nand U17140 (N_17140,N_16936,N_16856);
xor U17141 (N_17141,N_16847,N_16882);
or U17142 (N_17142,N_16894,N_16854);
or U17143 (N_17143,N_16878,N_16912);
and U17144 (N_17144,N_16988,N_16947);
nand U17145 (N_17145,N_16842,N_16915);
nand U17146 (N_17146,N_16814,N_16815);
xnor U17147 (N_17147,N_16858,N_16856);
and U17148 (N_17148,N_16897,N_16912);
nand U17149 (N_17149,N_16930,N_16801);
nand U17150 (N_17150,N_16802,N_16932);
and U17151 (N_17151,N_16964,N_16822);
xnor U17152 (N_17152,N_16884,N_16841);
xor U17153 (N_17153,N_16993,N_16994);
nor U17154 (N_17154,N_16995,N_16899);
nand U17155 (N_17155,N_16823,N_16908);
or U17156 (N_17156,N_16843,N_16937);
xnor U17157 (N_17157,N_16849,N_16887);
xnor U17158 (N_17158,N_16916,N_16946);
xor U17159 (N_17159,N_16879,N_16811);
nor U17160 (N_17160,N_16818,N_16924);
nor U17161 (N_17161,N_16890,N_16952);
xor U17162 (N_17162,N_16875,N_16874);
xor U17163 (N_17163,N_16856,N_16950);
nor U17164 (N_17164,N_16937,N_16947);
and U17165 (N_17165,N_16969,N_16878);
nand U17166 (N_17166,N_16832,N_16895);
or U17167 (N_17167,N_16875,N_16961);
nor U17168 (N_17168,N_16921,N_16834);
nand U17169 (N_17169,N_16872,N_16911);
nand U17170 (N_17170,N_16839,N_16869);
and U17171 (N_17171,N_16898,N_16992);
xnor U17172 (N_17172,N_16874,N_16905);
and U17173 (N_17173,N_16940,N_16884);
and U17174 (N_17174,N_16947,N_16954);
nand U17175 (N_17175,N_16814,N_16889);
xor U17176 (N_17176,N_16981,N_16983);
nor U17177 (N_17177,N_16855,N_16885);
and U17178 (N_17178,N_16834,N_16901);
and U17179 (N_17179,N_16969,N_16995);
xnor U17180 (N_17180,N_16890,N_16959);
nand U17181 (N_17181,N_16976,N_16916);
and U17182 (N_17182,N_16839,N_16929);
xor U17183 (N_17183,N_16963,N_16878);
or U17184 (N_17184,N_16954,N_16850);
nand U17185 (N_17185,N_16852,N_16835);
xor U17186 (N_17186,N_16857,N_16871);
nand U17187 (N_17187,N_16963,N_16954);
or U17188 (N_17188,N_16918,N_16864);
nand U17189 (N_17189,N_16870,N_16895);
or U17190 (N_17190,N_16889,N_16832);
nand U17191 (N_17191,N_16857,N_16922);
and U17192 (N_17192,N_16853,N_16894);
or U17193 (N_17193,N_16935,N_16802);
nand U17194 (N_17194,N_16846,N_16867);
or U17195 (N_17195,N_16990,N_16962);
nand U17196 (N_17196,N_16955,N_16886);
xnor U17197 (N_17197,N_16883,N_16835);
or U17198 (N_17198,N_16820,N_16935);
nor U17199 (N_17199,N_16958,N_16895);
nand U17200 (N_17200,N_17198,N_17147);
or U17201 (N_17201,N_17044,N_17100);
and U17202 (N_17202,N_17159,N_17077);
or U17203 (N_17203,N_17196,N_17004);
nand U17204 (N_17204,N_17127,N_17035);
nor U17205 (N_17205,N_17086,N_17118);
nor U17206 (N_17206,N_17050,N_17194);
and U17207 (N_17207,N_17136,N_17146);
nand U17208 (N_17208,N_17122,N_17131);
xnor U17209 (N_17209,N_17087,N_17169);
or U17210 (N_17210,N_17015,N_17030);
nand U17211 (N_17211,N_17121,N_17083);
nand U17212 (N_17212,N_17180,N_17082);
and U17213 (N_17213,N_17174,N_17167);
and U17214 (N_17214,N_17056,N_17037);
nand U17215 (N_17215,N_17098,N_17193);
or U17216 (N_17216,N_17094,N_17089);
nand U17217 (N_17217,N_17023,N_17101);
xnor U17218 (N_17218,N_17048,N_17027);
nand U17219 (N_17219,N_17079,N_17024);
and U17220 (N_17220,N_17085,N_17115);
xnor U17221 (N_17221,N_17172,N_17117);
and U17222 (N_17222,N_17154,N_17081);
nand U17223 (N_17223,N_17133,N_17187);
xor U17224 (N_17224,N_17008,N_17171);
xor U17225 (N_17225,N_17190,N_17033);
nor U17226 (N_17226,N_17074,N_17195);
or U17227 (N_17227,N_17152,N_17150);
or U17228 (N_17228,N_17104,N_17051);
xor U17229 (N_17229,N_17062,N_17179);
nor U17230 (N_17230,N_17175,N_17067);
or U17231 (N_17231,N_17058,N_17130);
nor U17232 (N_17232,N_17092,N_17064);
or U17233 (N_17233,N_17078,N_17096);
or U17234 (N_17234,N_17017,N_17156);
or U17235 (N_17235,N_17158,N_17139);
nor U17236 (N_17236,N_17123,N_17028);
xnor U17237 (N_17237,N_17076,N_17162);
xor U17238 (N_17238,N_17042,N_17163);
and U17239 (N_17239,N_17119,N_17025);
xor U17240 (N_17240,N_17183,N_17001);
xor U17241 (N_17241,N_17049,N_17059);
and U17242 (N_17242,N_17186,N_17138);
and U17243 (N_17243,N_17080,N_17151);
or U17244 (N_17244,N_17053,N_17165);
and U17245 (N_17245,N_17132,N_17075);
or U17246 (N_17246,N_17148,N_17181);
nor U17247 (N_17247,N_17091,N_17168);
or U17248 (N_17248,N_17057,N_17149);
nor U17249 (N_17249,N_17197,N_17066);
nand U17250 (N_17250,N_17061,N_17071);
and U17251 (N_17251,N_17107,N_17088);
or U17252 (N_17252,N_17128,N_17185);
or U17253 (N_17253,N_17142,N_17173);
nor U17254 (N_17254,N_17102,N_17093);
or U17255 (N_17255,N_17012,N_17105);
and U17256 (N_17256,N_17007,N_17054);
or U17257 (N_17257,N_17003,N_17182);
nand U17258 (N_17258,N_17170,N_17144);
nand U17259 (N_17259,N_17177,N_17014);
nor U17260 (N_17260,N_17099,N_17002);
or U17261 (N_17261,N_17164,N_17109);
nand U17262 (N_17262,N_17019,N_17191);
or U17263 (N_17263,N_17072,N_17010);
or U17264 (N_17264,N_17120,N_17047);
and U17265 (N_17265,N_17060,N_17039);
nor U17266 (N_17266,N_17124,N_17199);
or U17267 (N_17267,N_17009,N_17106);
nor U17268 (N_17268,N_17129,N_17022);
nor U17269 (N_17269,N_17026,N_17112);
and U17270 (N_17270,N_17108,N_17097);
xor U17271 (N_17271,N_17111,N_17192);
nand U17272 (N_17272,N_17137,N_17038);
nand U17273 (N_17273,N_17032,N_17063);
nor U17274 (N_17274,N_17020,N_17161);
nor U17275 (N_17275,N_17103,N_17188);
and U17276 (N_17276,N_17176,N_17155);
xnor U17277 (N_17277,N_17021,N_17070);
and U17278 (N_17278,N_17189,N_17095);
nor U17279 (N_17279,N_17068,N_17126);
nand U17280 (N_17280,N_17184,N_17052);
nor U17281 (N_17281,N_17073,N_17114);
xor U17282 (N_17282,N_17018,N_17113);
and U17283 (N_17283,N_17090,N_17029);
or U17284 (N_17284,N_17140,N_17110);
xnor U17285 (N_17285,N_17036,N_17143);
nor U17286 (N_17286,N_17046,N_17005);
nor U17287 (N_17287,N_17145,N_17011);
and U17288 (N_17288,N_17134,N_17031);
nand U17289 (N_17289,N_17178,N_17125);
nand U17290 (N_17290,N_17084,N_17013);
or U17291 (N_17291,N_17055,N_17040);
or U17292 (N_17292,N_17065,N_17045);
and U17293 (N_17293,N_17043,N_17116);
or U17294 (N_17294,N_17157,N_17041);
and U17295 (N_17295,N_17160,N_17153);
nor U17296 (N_17296,N_17016,N_17006);
or U17297 (N_17297,N_17000,N_17034);
xor U17298 (N_17298,N_17141,N_17166);
and U17299 (N_17299,N_17135,N_17069);
nor U17300 (N_17300,N_17195,N_17053);
and U17301 (N_17301,N_17013,N_17093);
and U17302 (N_17302,N_17006,N_17031);
and U17303 (N_17303,N_17003,N_17144);
xnor U17304 (N_17304,N_17160,N_17197);
or U17305 (N_17305,N_17031,N_17086);
nor U17306 (N_17306,N_17019,N_17144);
and U17307 (N_17307,N_17043,N_17137);
and U17308 (N_17308,N_17067,N_17090);
or U17309 (N_17309,N_17097,N_17093);
nor U17310 (N_17310,N_17190,N_17094);
xor U17311 (N_17311,N_17113,N_17197);
xnor U17312 (N_17312,N_17024,N_17007);
xor U17313 (N_17313,N_17095,N_17106);
nor U17314 (N_17314,N_17022,N_17066);
or U17315 (N_17315,N_17165,N_17115);
xor U17316 (N_17316,N_17166,N_17156);
nand U17317 (N_17317,N_17119,N_17184);
nand U17318 (N_17318,N_17098,N_17195);
nor U17319 (N_17319,N_17120,N_17011);
or U17320 (N_17320,N_17108,N_17126);
nand U17321 (N_17321,N_17166,N_17056);
nand U17322 (N_17322,N_17038,N_17173);
nand U17323 (N_17323,N_17010,N_17156);
and U17324 (N_17324,N_17169,N_17162);
nand U17325 (N_17325,N_17182,N_17017);
nor U17326 (N_17326,N_17029,N_17121);
nand U17327 (N_17327,N_17051,N_17022);
or U17328 (N_17328,N_17064,N_17036);
nor U17329 (N_17329,N_17139,N_17104);
or U17330 (N_17330,N_17056,N_17093);
or U17331 (N_17331,N_17194,N_17103);
nand U17332 (N_17332,N_17061,N_17001);
xnor U17333 (N_17333,N_17065,N_17129);
or U17334 (N_17334,N_17101,N_17091);
and U17335 (N_17335,N_17012,N_17170);
nand U17336 (N_17336,N_17059,N_17107);
nand U17337 (N_17337,N_17042,N_17104);
or U17338 (N_17338,N_17163,N_17171);
xor U17339 (N_17339,N_17049,N_17102);
nand U17340 (N_17340,N_17106,N_17164);
and U17341 (N_17341,N_17075,N_17178);
nor U17342 (N_17342,N_17098,N_17003);
or U17343 (N_17343,N_17152,N_17077);
or U17344 (N_17344,N_17108,N_17027);
xnor U17345 (N_17345,N_17026,N_17053);
or U17346 (N_17346,N_17097,N_17020);
nor U17347 (N_17347,N_17037,N_17197);
nand U17348 (N_17348,N_17023,N_17152);
and U17349 (N_17349,N_17152,N_17060);
xor U17350 (N_17350,N_17092,N_17127);
and U17351 (N_17351,N_17016,N_17158);
or U17352 (N_17352,N_17037,N_17176);
or U17353 (N_17353,N_17176,N_17075);
nand U17354 (N_17354,N_17012,N_17005);
nor U17355 (N_17355,N_17077,N_17060);
and U17356 (N_17356,N_17147,N_17112);
and U17357 (N_17357,N_17030,N_17101);
or U17358 (N_17358,N_17022,N_17154);
xor U17359 (N_17359,N_17024,N_17058);
nor U17360 (N_17360,N_17005,N_17008);
nand U17361 (N_17361,N_17063,N_17098);
nand U17362 (N_17362,N_17081,N_17151);
and U17363 (N_17363,N_17040,N_17167);
nand U17364 (N_17364,N_17071,N_17073);
nand U17365 (N_17365,N_17113,N_17038);
and U17366 (N_17366,N_17073,N_17092);
xor U17367 (N_17367,N_17182,N_17024);
nor U17368 (N_17368,N_17179,N_17104);
and U17369 (N_17369,N_17005,N_17098);
nor U17370 (N_17370,N_17012,N_17021);
nand U17371 (N_17371,N_17019,N_17159);
nand U17372 (N_17372,N_17084,N_17112);
xnor U17373 (N_17373,N_17147,N_17074);
nand U17374 (N_17374,N_17048,N_17102);
xor U17375 (N_17375,N_17166,N_17124);
xor U17376 (N_17376,N_17042,N_17105);
nor U17377 (N_17377,N_17097,N_17022);
xor U17378 (N_17378,N_17129,N_17123);
nand U17379 (N_17379,N_17034,N_17098);
and U17380 (N_17380,N_17191,N_17129);
xor U17381 (N_17381,N_17164,N_17150);
nor U17382 (N_17382,N_17194,N_17109);
nand U17383 (N_17383,N_17086,N_17184);
or U17384 (N_17384,N_17173,N_17130);
xnor U17385 (N_17385,N_17115,N_17155);
xor U17386 (N_17386,N_17085,N_17157);
and U17387 (N_17387,N_17178,N_17127);
or U17388 (N_17388,N_17114,N_17050);
xor U17389 (N_17389,N_17145,N_17149);
nand U17390 (N_17390,N_17023,N_17126);
or U17391 (N_17391,N_17041,N_17049);
and U17392 (N_17392,N_17044,N_17144);
nor U17393 (N_17393,N_17110,N_17080);
and U17394 (N_17394,N_17087,N_17157);
nor U17395 (N_17395,N_17146,N_17195);
xnor U17396 (N_17396,N_17094,N_17092);
xnor U17397 (N_17397,N_17145,N_17162);
or U17398 (N_17398,N_17169,N_17132);
nand U17399 (N_17399,N_17164,N_17058);
xnor U17400 (N_17400,N_17280,N_17259);
and U17401 (N_17401,N_17336,N_17334);
or U17402 (N_17402,N_17298,N_17331);
nor U17403 (N_17403,N_17385,N_17307);
and U17404 (N_17404,N_17201,N_17284);
nor U17405 (N_17405,N_17384,N_17202);
or U17406 (N_17406,N_17268,N_17363);
or U17407 (N_17407,N_17226,N_17275);
nor U17408 (N_17408,N_17227,N_17300);
nand U17409 (N_17409,N_17208,N_17231);
nand U17410 (N_17410,N_17313,N_17326);
xor U17411 (N_17411,N_17377,N_17248);
nand U17412 (N_17412,N_17253,N_17262);
or U17413 (N_17413,N_17210,N_17368);
xnor U17414 (N_17414,N_17371,N_17256);
or U17415 (N_17415,N_17299,N_17249);
xor U17416 (N_17416,N_17347,N_17203);
nand U17417 (N_17417,N_17351,N_17391);
and U17418 (N_17418,N_17346,N_17367);
nor U17419 (N_17419,N_17213,N_17247);
xor U17420 (N_17420,N_17221,N_17293);
xnor U17421 (N_17421,N_17333,N_17392);
and U17422 (N_17422,N_17276,N_17328);
xor U17423 (N_17423,N_17321,N_17200);
and U17424 (N_17424,N_17270,N_17322);
xnor U17425 (N_17425,N_17358,N_17397);
nor U17426 (N_17426,N_17225,N_17278);
and U17427 (N_17427,N_17327,N_17297);
and U17428 (N_17428,N_17264,N_17265);
and U17429 (N_17429,N_17303,N_17244);
nand U17430 (N_17430,N_17219,N_17261);
or U17431 (N_17431,N_17266,N_17332);
nor U17432 (N_17432,N_17323,N_17250);
or U17433 (N_17433,N_17204,N_17273);
nor U17434 (N_17434,N_17315,N_17362);
and U17435 (N_17435,N_17209,N_17366);
xor U17436 (N_17436,N_17390,N_17240);
or U17437 (N_17437,N_17373,N_17364);
and U17438 (N_17438,N_17337,N_17387);
nor U17439 (N_17439,N_17343,N_17237);
or U17440 (N_17440,N_17330,N_17207);
or U17441 (N_17441,N_17286,N_17238);
and U17442 (N_17442,N_17229,N_17290);
nor U17443 (N_17443,N_17230,N_17251);
nand U17444 (N_17444,N_17232,N_17356);
and U17445 (N_17445,N_17301,N_17393);
nand U17446 (N_17446,N_17379,N_17214);
nand U17447 (N_17447,N_17394,N_17295);
nor U17448 (N_17448,N_17271,N_17254);
nor U17449 (N_17449,N_17381,N_17329);
or U17450 (N_17450,N_17352,N_17296);
xor U17451 (N_17451,N_17241,N_17269);
nor U17452 (N_17452,N_17292,N_17388);
and U17453 (N_17453,N_17376,N_17304);
nand U17454 (N_17454,N_17339,N_17340);
and U17455 (N_17455,N_17345,N_17324);
nor U17456 (N_17456,N_17236,N_17320);
or U17457 (N_17457,N_17342,N_17206);
or U17458 (N_17458,N_17257,N_17223);
nor U17459 (N_17459,N_17314,N_17220);
and U17460 (N_17460,N_17306,N_17309);
or U17461 (N_17461,N_17382,N_17370);
or U17462 (N_17462,N_17305,N_17216);
and U17463 (N_17463,N_17294,N_17258);
xor U17464 (N_17464,N_17234,N_17235);
nand U17465 (N_17465,N_17374,N_17360);
and U17466 (N_17466,N_17325,N_17383);
or U17467 (N_17467,N_17282,N_17375);
or U17468 (N_17468,N_17335,N_17398);
and U17469 (N_17469,N_17380,N_17310);
nor U17470 (N_17470,N_17277,N_17399);
and U17471 (N_17471,N_17218,N_17243);
and U17472 (N_17472,N_17378,N_17349);
xor U17473 (N_17473,N_17289,N_17372);
xor U17474 (N_17474,N_17267,N_17274);
or U17475 (N_17475,N_17212,N_17287);
nor U17476 (N_17476,N_17255,N_17386);
nor U17477 (N_17477,N_17361,N_17291);
nor U17478 (N_17478,N_17354,N_17283);
nand U17479 (N_17479,N_17228,N_17365);
and U17480 (N_17480,N_17355,N_17396);
nor U17481 (N_17481,N_17205,N_17350);
xor U17482 (N_17482,N_17308,N_17341);
nor U17483 (N_17483,N_17389,N_17288);
and U17484 (N_17484,N_17245,N_17312);
or U17485 (N_17485,N_17211,N_17222);
xnor U17486 (N_17486,N_17318,N_17395);
nand U17487 (N_17487,N_17316,N_17281);
nor U17488 (N_17488,N_17311,N_17246);
xor U17489 (N_17489,N_17302,N_17260);
xnor U17490 (N_17490,N_17357,N_17369);
or U17491 (N_17491,N_17272,N_17344);
and U17492 (N_17492,N_17359,N_17338);
and U17493 (N_17493,N_17348,N_17239);
nand U17494 (N_17494,N_17263,N_17242);
and U17495 (N_17495,N_17224,N_17217);
nor U17496 (N_17496,N_17353,N_17279);
and U17497 (N_17497,N_17233,N_17252);
or U17498 (N_17498,N_17319,N_17285);
or U17499 (N_17499,N_17317,N_17215);
xor U17500 (N_17500,N_17278,N_17216);
or U17501 (N_17501,N_17343,N_17301);
or U17502 (N_17502,N_17328,N_17278);
nor U17503 (N_17503,N_17266,N_17222);
nand U17504 (N_17504,N_17221,N_17226);
and U17505 (N_17505,N_17213,N_17319);
xnor U17506 (N_17506,N_17205,N_17374);
or U17507 (N_17507,N_17399,N_17320);
and U17508 (N_17508,N_17353,N_17395);
and U17509 (N_17509,N_17208,N_17301);
and U17510 (N_17510,N_17394,N_17203);
xnor U17511 (N_17511,N_17287,N_17363);
nand U17512 (N_17512,N_17254,N_17384);
nor U17513 (N_17513,N_17259,N_17367);
xnor U17514 (N_17514,N_17338,N_17355);
nor U17515 (N_17515,N_17227,N_17269);
or U17516 (N_17516,N_17398,N_17329);
or U17517 (N_17517,N_17336,N_17265);
or U17518 (N_17518,N_17316,N_17380);
and U17519 (N_17519,N_17203,N_17387);
nand U17520 (N_17520,N_17303,N_17377);
nor U17521 (N_17521,N_17282,N_17202);
nand U17522 (N_17522,N_17367,N_17204);
or U17523 (N_17523,N_17273,N_17201);
and U17524 (N_17524,N_17339,N_17360);
nor U17525 (N_17525,N_17304,N_17363);
nand U17526 (N_17526,N_17208,N_17360);
or U17527 (N_17527,N_17370,N_17373);
xor U17528 (N_17528,N_17270,N_17280);
and U17529 (N_17529,N_17366,N_17281);
and U17530 (N_17530,N_17365,N_17258);
nor U17531 (N_17531,N_17311,N_17294);
and U17532 (N_17532,N_17357,N_17283);
and U17533 (N_17533,N_17346,N_17359);
nand U17534 (N_17534,N_17255,N_17240);
xnor U17535 (N_17535,N_17294,N_17318);
nor U17536 (N_17536,N_17268,N_17244);
or U17537 (N_17537,N_17270,N_17388);
xor U17538 (N_17538,N_17284,N_17210);
nand U17539 (N_17539,N_17319,N_17346);
or U17540 (N_17540,N_17363,N_17270);
nand U17541 (N_17541,N_17389,N_17265);
or U17542 (N_17542,N_17271,N_17289);
nor U17543 (N_17543,N_17280,N_17352);
nand U17544 (N_17544,N_17382,N_17250);
xnor U17545 (N_17545,N_17376,N_17241);
nor U17546 (N_17546,N_17393,N_17311);
xnor U17547 (N_17547,N_17309,N_17281);
xnor U17548 (N_17548,N_17384,N_17272);
xor U17549 (N_17549,N_17285,N_17294);
xor U17550 (N_17550,N_17328,N_17263);
and U17551 (N_17551,N_17308,N_17291);
nand U17552 (N_17552,N_17339,N_17253);
or U17553 (N_17553,N_17273,N_17303);
nand U17554 (N_17554,N_17372,N_17249);
nor U17555 (N_17555,N_17259,N_17313);
nor U17556 (N_17556,N_17240,N_17378);
or U17557 (N_17557,N_17267,N_17219);
nand U17558 (N_17558,N_17209,N_17212);
and U17559 (N_17559,N_17374,N_17204);
nand U17560 (N_17560,N_17272,N_17287);
nor U17561 (N_17561,N_17369,N_17220);
and U17562 (N_17562,N_17250,N_17317);
nor U17563 (N_17563,N_17247,N_17260);
xor U17564 (N_17564,N_17205,N_17366);
nor U17565 (N_17565,N_17283,N_17293);
and U17566 (N_17566,N_17240,N_17374);
nor U17567 (N_17567,N_17260,N_17359);
or U17568 (N_17568,N_17320,N_17215);
nor U17569 (N_17569,N_17282,N_17277);
nand U17570 (N_17570,N_17293,N_17209);
nor U17571 (N_17571,N_17234,N_17347);
xor U17572 (N_17572,N_17394,N_17362);
nand U17573 (N_17573,N_17392,N_17385);
xnor U17574 (N_17574,N_17288,N_17337);
or U17575 (N_17575,N_17345,N_17267);
or U17576 (N_17576,N_17325,N_17304);
nor U17577 (N_17577,N_17224,N_17206);
xor U17578 (N_17578,N_17244,N_17254);
or U17579 (N_17579,N_17205,N_17299);
and U17580 (N_17580,N_17269,N_17207);
and U17581 (N_17581,N_17320,N_17304);
xor U17582 (N_17582,N_17356,N_17382);
xnor U17583 (N_17583,N_17206,N_17330);
xor U17584 (N_17584,N_17298,N_17318);
and U17585 (N_17585,N_17259,N_17281);
and U17586 (N_17586,N_17399,N_17296);
xnor U17587 (N_17587,N_17327,N_17241);
or U17588 (N_17588,N_17318,N_17367);
nand U17589 (N_17589,N_17350,N_17331);
or U17590 (N_17590,N_17389,N_17380);
or U17591 (N_17591,N_17242,N_17230);
xor U17592 (N_17592,N_17388,N_17355);
and U17593 (N_17593,N_17380,N_17268);
nor U17594 (N_17594,N_17296,N_17226);
nor U17595 (N_17595,N_17259,N_17334);
xnor U17596 (N_17596,N_17391,N_17361);
nand U17597 (N_17597,N_17276,N_17304);
and U17598 (N_17598,N_17262,N_17252);
nand U17599 (N_17599,N_17275,N_17316);
or U17600 (N_17600,N_17516,N_17521);
or U17601 (N_17601,N_17518,N_17592);
and U17602 (N_17602,N_17568,N_17599);
nor U17603 (N_17603,N_17407,N_17548);
nand U17604 (N_17604,N_17528,N_17536);
xor U17605 (N_17605,N_17429,N_17538);
or U17606 (N_17606,N_17559,N_17546);
nor U17607 (N_17607,N_17519,N_17491);
and U17608 (N_17608,N_17591,N_17442);
nand U17609 (N_17609,N_17486,N_17462);
nand U17610 (N_17610,N_17417,N_17569);
xor U17611 (N_17611,N_17514,N_17474);
xor U17612 (N_17612,N_17461,N_17595);
nor U17613 (N_17613,N_17499,N_17594);
nand U17614 (N_17614,N_17423,N_17476);
and U17615 (N_17615,N_17404,N_17481);
nand U17616 (N_17616,N_17531,N_17441);
xnor U17617 (N_17617,N_17574,N_17421);
and U17618 (N_17618,N_17490,N_17494);
or U17619 (N_17619,N_17576,N_17509);
xnor U17620 (N_17620,N_17480,N_17517);
or U17621 (N_17621,N_17470,N_17586);
nor U17622 (N_17622,N_17506,N_17411);
xor U17623 (N_17623,N_17500,N_17504);
or U17624 (N_17624,N_17415,N_17552);
or U17625 (N_17625,N_17467,N_17501);
nand U17626 (N_17626,N_17505,N_17414);
nand U17627 (N_17627,N_17428,N_17406);
or U17628 (N_17628,N_17572,N_17471);
and U17629 (N_17629,N_17450,N_17497);
or U17630 (N_17630,N_17543,N_17431);
xor U17631 (N_17631,N_17403,N_17444);
nand U17632 (N_17632,N_17535,N_17458);
and U17633 (N_17633,N_17520,N_17537);
and U17634 (N_17634,N_17453,N_17589);
nand U17635 (N_17635,N_17454,N_17426);
nor U17636 (N_17636,N_17580,N_17456);
nor U17637 (N_17637,N_17511,N_17405);
nand U17638 (N_17638,N_17451,N_17425);
and U17639 (N_17639,N_17579,N_17432);
nor U17640 (N_17640,N_17557,N_17547);
nor U17641 (N_17641,N_17402,N_17488);
nor U17642 (N_17642,N_17484,N_17408);
xor U17643 (N_17643,N_17460,N_17598);
nand U17644 (N_17644,N_17447,N_17584);
nand U17645 (N_17645,N_17560,N_17446);
nor U17646 (N_17646,N_17443,N_17472);
and U17647 (N_17647,N_17561,N_17544);
or U17648 (N_17648,N_17495,N_17455);
and U17649 (N_17649,N_17545,N_17555);
xor U17650 (N_17650,N_17427,N_17412);
nor U17651 (N_17651,N_17558,N_17597);
nand U17652 (N_17652,N_17507,N_17590);
nor U17653 (N_17653,N_17577,N_17524);
nor U17654 (N_17654,N_17430,N_17510);
nor U17655 (N_17655,N_17448,N_17593);
and U17656 (N_17656,N_17463,N_17573);
nor U17657 (N_17657,N_17554,N_17483);
nor U17658 (N_17658,N_17588,N_17475);
nand U17659 (N_17659,N_17469,N_17409);
and U17660 (N_17660,N_17473,N_17401);
or U17661 (N_17661,N_17416,N_17527);
xor U17662 (N_17662,N_17468,N_17479);
or U17663 (N_17663,N_17477,N_17542);
and U17664 (N_17664,N_17526,N_17457);
or U17665 (N_17665,N_17549,N_17419);
nand U17666 (N_17666,N_17541,N_17496);
or U17667 (N_17667,N_17512,N_17437);
and U17668 (N_17668,N_17533,N_17540);
and U17669 (N_17669,N_17478,N_17465);
nor U17670 (N_17670,N_17513,N_17581);
xnor U17671 (N_17671,N_17565,N_17485);
and U17672 (N_17672,N_17571,N_17413);
and U17673 (N_17673,N_17529,N_17436);
nand U17674 (N_17674,N_17566,N_17418);
or U17675 (N_17675,N_17439,N_17530);
nand U17676 (N_17676,N_17570,N_17424);
nand U17677 (N_17677,N_17582,N_17422);
xor U17678 (N_17678,N_17438,N_17452);
nand U17679 (N_17679,N_17587,N_17449);
nand U17680 (N_17680,N_17551,N_17532);
nor U17681 (N_17681,N_17585,N_17420);
nand U17682 (N_17682,N_17492,N_17522);
nor U17683 (N_17683,N_17482,N_17433);
and U17684 (N_17684,N_17575,N_17523);
xnor U17685 (N_17685,N_17550,N_17502);
xnor U17686 (N_17686,N_17578,N_17487);
xor U17687 (N_17687,N_17508,N_17466);
nand U17688 (N_17688,N_17539,N_17410);
or U17689 (N_17689,N_17445,N_17435);
and U17690 (N_17690,N_17556,N_17434);
nand U17691 (N_17691,N_17525,N_17567);
nor U17692 (N_17692,N_17440,N_17534);
and U17693 (N_17693,N_17596,N_17459);
or U17694 (N_17694,N_17400,N_17563);
or U17695 (N_17695,N_17489,N_17503);
xor U17696 (N_17696,N_17553,N_17498);
xor U17697 (N_17697,N_17464,N_17583);
nor U17698 (N_17698,N_17493,N_17564);
xnor U17699 (N_17699,N_17562,N_17515);
nand U17700 (N_17700,N_17517,N_17497);
and U17701 (N_17701,N_17420,N_17516);
xnor U17702 (N_17702,N_17444,N_17471);
nand U17703 (N_17703,N_17529,N_17566);
and U17704 (N_17704,N_17546,N_17496);
xor U17705 (N_17705,N_17411,N_17557);
nor U17706 (N_17706,N_17504,N_17581);
nand U17707 (N_17707,N_17439,N_17569);
nand U17708 (N_17708,N_17444,N_17530);
and U17709 (N_17709,N_17519,N_17422);
xnor U17710 (N_17710,N_17525,N_17501);
nand U17711 (N_17711,N_17461,N_17568);
xnor U17712 (N_17712,N_17487,N_17448);
or U17713 (N_17713,N_17453,N_17401);
xnor U17714 (N_17714,N_17477,N_17472);
nor U17715 (N_17715,N_17525,N_17471);
and U17716 (N_17716,N_17496,N_17436);
and U17717 (N_17717,N_17525,N_17570);
xnor U17718 (N_17718,N_17405,N_17541);
and U17719 (N_17719,N_17508,N_17476);
and U17720 (N_17720,N_17570,N_17471);
nor U17721 (N_17721,N_17418,N_17491);
or U17722 (N_17722,N_17569,N_17416);
and U17723 (N_17723,N_17503,N_17584);
xnor U17724 (N_17724,N_17547,N_17462);
or U17725 (N_17725,N_17493,N_17461);
nor U17726 (N_17726,N_17470,N_17439);
xnor U17727 (N_17727,N_17528,N_17495);
xnor U17728 (N_17728,N_17529,N_17446);
or U17729 (N_17729,N_17445,N_17578);
or U17730 (N_17730,N_17458,N_17402);
nor U17731 (N_17731,N_17523,N_17572);
nand U17732 (N_17732,N_17435,N_17488);
nand U17733 (N_17733,N_17574,N_17522);
or U17734 (N_17734,N_17575,N_17571);
and U17735 (N_17735,N_17431,N_17466);
and U17736 (N_17736,N_17440,N_17528);
nor U17737 (N_17737,N_17414,N_17401);
nand U17738 (N_17738,N_17480,N_17428);
xnor U17739 (N_17739,N_17437,N_17504);
and U17740 (N_17740,N_17487,N_17497);
and U17741 (N_17741,N_17596,N_17454);
or U17742 (N_17742,N_17547,N_17541);
nor U17743 (N_17743,N_17487,N_17522);
nand U17744 (N_17744,N_17518,N_17574);
and U17745 (N_17745,N_17424,N_17555);
or U17746 (N_17746,N_17436,N_17459);
xor U17747 (N_17747,N_17543,N_17573);
nand U17748 (N_17748,N_17459,N_17513);
xor U17749 (N_17749,N_17453,N_17555);
nand U17750 (N_17750,N_17463,N_17503);
nor U17751 (N_17751,N_17591,N_17560);
nor U17752 (N_17752,N_17410,N_17520);
and U17753 (N_17753,N_17432,N_17487);
or U17754 (N_17754,N_17501,N_17533);
nor U17755 (N_17755,N_17544,N_17457);
nor U17756 (N_17756,N_17485,N_17463);
and U17757 (N_17757,N_17594,N_17542);
nor U17758 (N_17758,N_17461,N_17491);
nor U17759 (N_17759,N_17533,N_17478);
or U17760 (N_17760,N_17552,N_17421);
nor U17761 (N_17761,N_17418,N_17411);
nor U17762 (N_17762,N_17547,N_17528);
nand U17763 (N_17763,N_17490,N_17423);
nand U17764 (N_17764,N_17555,N_17494);
and U17765 (N_17765,N_17531,N_17507);
xor U17766 (N_17766,N_17423,N_17596);
or U17767 (N_17767,N_17536,N_17507);
nor U17768 (N_17768,N_17562,N_17485);
and U17769 (N_17769,N_17541,N_17485);
xor U17770 (N_17770,N_17502,N_17404);
and U17771 (N_17771,N_17560,N_17542);
nor U17772 (N_17772,N_17529,N_17420);
and U17773 (N_17773,N_17570,N_17439);
nand U17774 (N_17774,N_17451,N_17426);
nor U17775 (N_17775,N_17507,N_17495);
xnor U17776 (N_17776,N_17544,N_17503);
nand U17777 (N_17777,N_17576,N_17408);
nor U17778 (N_17778,N_17544,N_17572);
or U17779 (N_17779,N_17438,N_17484);
nand U17780 (N_17780,N_17444,N_17526);
nor U17781 (N_17781,N_17474,N_17587);
xnor U17782 (N_17782,N_17468,N_17413);
or U17783 (N_17783,N_17501,N_17413);
and U17784 (N_17784,N_17584,N_17558);
xnor U17785 (N_17785,N_17563,N_17494);
or U17786 (N_17786,N_17581,N_17515);
nand U17787 (N_17787,N_17484,N_17459);
and U17788 (N_17788,N_17425,N_17429);
xor U17789 (N_17789,N_17400,N_17545);
nor U17790 (N_17790,N_17427,N_17441);
nor U17791 (N_17791,N_17598,N_17496);
or U17792 (N_17792,N_17549,N_17448);
nand U17793 (N_17793,N_17497,N_17562);
xor U17794 (N_17794,N_17565,N_17521);
and U17795 (N_17795,N_17584,N_17403);
nor U17796 (N_17796,N_17523,N_17513);
or U17797 (N_17797,N_17434,N_17466);
and U17798 (N_17798,N_17424,N_17511);
xor U17799 (N_17799,N_17515,N_17457);
or U17800 (N_17800,N_17744,N_17727);
and U17801 (N_17801,N_17639,N_17787);
and U17802 (N_17802,N_17795,N_17612);
xnor U17803 (N_17803,N_17672,N_17750);
nor U17804 (N_17804,N_17792,N_17660);
or U17805 (N_17805,N_17670,N_17609);
or U17806 (N_17806,N_17668,N_17725);
nor U17807 (N_17807,N_17752,N_17679);
xnor U17808 (N_17808,N_17721,N_17729);
nand U17809 (N_17809,N_17793,N_17755);
xnor U17810 (N_17810,N_17693,N_17602);
nor U17811 (N_17811,N_17673,N_17620);
nand U17812 (N_17812,N_17601,N_17610);
nor U17813 (N_17813,N_17734,N_17799);
and U17814 (N_17814,N_17694,N_17716);
xor U17815 (N_17815,N_17798,N_17748);
and U17816 (N_17816,N_17652,N_17768);
nand U17817 (N_17817,N_17707,N_17700);
and U17818 (N_17818,N_17736,N_17715);
and U17819 (N_17819,N_17739,N_17770);
nand U17820 (N_17820,N_17765,N_17681);
and U17821 (N_17821,N_17684,N_17796);
or U17822 (N_17822,N_17701,N_17780);
nand U17823 (N_17823,N_17733,N_17615);
or U17824 (N_17824,N_17758,N_17712);
or U17825 (N_17825,N_17636,N_17779);
nor U17826 (N_17826,N_17666,N_17608);
nand U17827 (N_17827,N_17731,N_17726);
and U17828 (N_17828,N_17753,N_17789);
nand U17829 (N_17829,N_17738,N_17746);
and U17830 (N_17830,N_17688,N_17754);
and U17831 (N_17831,N_17760,N_17641);
xnor U17832 (N_17832,N_17767,N_17719);
nor U17833 (N_17833,N_17689,N_17613);
and U17834 (N_17834,N_17686,N_17617);
nand U17835 (N_17835,N_17614,N_17711);
nor U17836 (N_17836,N_17654,N_17717);
nand U17837 (N_17837,N_17775,N_17647);
nor U17838 (N_17838,N_17674,N_17783);
xor U17839 (N_17839,N_17737,N_17691);
nor U17840 (N_17840,N_17687,N_17624);
or U17841 (N_17841,N_17713,N_17678);
xnor U17842 (N_17842,N_17642,N_17606);
nor U17843 (N_17843,N_17742,N_17600);
xnor U17844 (N_17844,N_17782,N_17784);
nor U17845 (N_17845,N_17762,N_17671);
or U17846 (N_17846,N_17619,N_17661);
or U17847 (N_17847,N_17720,N_17616);
or U17848 (N_17848,N_17658,N_17667);
and U17849 (N_17849,N_17773,N_17683);
xor U17850 (N_17850,N_17644,N_17643);
and U17851 (N_17851,N_17634,N_17766);
nand U17852 (N_17852,N_17776,N_17769);
nor U17853 (N_17853,N_17669,N_17645);
nand U17854 (N_17854,N_17622,N_17651);
nor U17855 (N_17855,N_17648,N_17743);
nor U17856 (N_17856,N_17698,N_17695);
nor U17857 (N_17857,N_17665,N_17618);
and U17858 (N_17858,N_17764,N_17611);
nand U17859 (N_17859,N_17625,N_17794);
nor U17860 (N_17860,N_17680,N_17649);
and U17861 (N_17861,N_17756,N_17763);
and U17862 (N_17862,N_17685,N_17692);
nand U17863 (N_17863,N_17722,N_17708);
xor U17864 (N_17864,N_17637,N_17677);
xnor U17865 (N_17865,N_17761,N_17697);
or U17866 (N_17866,N_17638,N_17718);
or U17867 (N_17867,N_17772,N_17771);
nor U17868 (N_17868,N_17633,N_17714);
and U17869 (N_17869,N_17745,N_17728);
xnor U17870 (N_17870,N_17788,N_17626);
nand U17871 (N_17871,N_17732,N_17740);
nor U17872 (N_17872,N_17646,N_17621);
or U17873 (N_17873,N_17604,N_17751);
nand U17874 (N_17874,N_17778,N_17741);
nor U17875 (N_17875,N_17749,N_17705);
nor U17876 (N_17876,N_17786,N_17735);
xnor U17877 (N_17877,N_17696,N_17659);
nor U17878 (N_17878,N_17797,N_17709);
and U17879 (N_17879,N_17629,N_17664);
nand U17880 (N_17880,N_17632,N_17747);
nand U17881 (N_17881,N_17650,N_17759);
xor U17882 (N_17882,N_17657,N_17623);
nor U17883 (N_17883,N_17628,N_17702);
and U17884 (N_17884,N_17730,N_17631);
nor U17885 (N_17885,N_17723,N_17785);
xor U17886 (N_17886,N_17655,N_17699);
xnor U17887 (N_17887,N_17710,N_17777);
xor U17888 (N_17888,N_17682,N_17690);
nand U17889 (N_17889,N_17653,N_17703);
nor U17890 (N_17890,N_17656,N_17724);
or U17891 (N_17891,N_17605,N_17774);
xor U17892 (N_17892,N_17757,N_17706);
xor U17893 (N_17893,N_17627,N_17790);
xor U17894 (N_17894,N_17635,N_17640);
nor U17895 (N_17895,N_17675,N_17791);
nor U17896 (N_17896,N_17663,N_17603);
nor U17897 (N_17897,N_17676,N_17630);
nor U17898 (N_17898,N_17704,N_17662);
and U17899 (N_17899,N_17781,N_17607);
nor U17900 (N_17900,N_17635,N_17629);
nand U17901 (N_17901,N_17696,N_17642);
or U17902 (N_17902,N_17629,N_17654);
xor U17903 (N_17903,N_17618,N_17663);
nor U17904 (N_17904,N_17665,N_17721);
and U17905 (N_17905,N_17663,N_17735);
nor U17906 (N_17906,N_17734,N_17604);
xnor U17907 (N_17907,N_17722,N_17755);
nand U17908 (N_17908,N_17718,N_17602);
and U17909 (N_17909,N_17685,N_17781);
or U17910 (N_17910,N_17750,N_17698);
nor U17911 (N_17911,N_17620,N_17720);
and U17912 (N_17912,N_17681,N_17691);
or U17913 (N_17913,N_17717,N_17662);
or U17914 (N_17914,N_17738,N_17651);
nor U17915 (N_17915,N_17637,N_17721);
and U17916 (N_17916,N_17710,N_17770);
and U17917 (N_17917,N_17658,N_17642);
and U17918 (N_17918,N_17627,N_17723);
nor U17919 (N_17919,N_17766,N_17627);
nand U17920 (N_17920,N_17638,N_17660);
nor U17921 (N_17921,N_17652,N_17740);
or U17922 (N_17922,N_17656,N_17631);
nor U17923 (N_17923,N_17766,N_17792);
nand U17924 (N_17924,N_17738,N_17794);
and U17925 (N_17925,N_17759,N_17685);
and U17926 (N_17926,N_17692,N_17630);
xnor U17927 (N_17927,N_17765,N_17686);
or U17928 (N_17928,N_17712,N_17793);
nand U17929 (N_17929,N_17664,N_17763);
nand U17930 (N_17930,N_17724,N_17647);
and U17931 (N_17931,N_17719,N_17772);
or U17932 (N_17932,N_17717,N_17719);
nand U17933 (N_17933,N_17776,N_17670);
or U17934 (N_17934,N_17757,N_17704);
xor U17935 (N_17935,N_17653,N_17624);
xor U17936 (N_17936,N_17656,N_17787);
nor U17937 (N_17937,N_17666,N_17673);
nand U17938 (N_17938,N_17672,N_17794);
xor U17939 (N_17939,N_17742,N_17691);
nor U17940 (N_17940,N_17605,N_17644);
nor U17941 (N_17941,N_17724,N_17616);
and U17942 (N_17942,N_17772,N_17652);
xor U17943 (N_17943,N_17662,N_17782);
or U17944 (N_17944,N_17766,N_17721);
or U17945 (N_17945,N_17714,N_17632);
and U17946 (N_17946,N_17612,N_17661);
and U17947 (N_17947,N_17751,N_17772);
nand U17948 (N_17948,N_17670,N_17687);
nand U17949 (N_17949,N_17790,N_17750);
or U17950 (N_17950,N_17731,N_17759);
xor U17951 (N_17951,N_17705,N_17758);
xor U17952 (N_17952,N_17652,N_17792);
and U17953 (N_17953,N_17746,N_17618);
and U17954 (N_17954,N_17669,N_17710);
xnor U17955 (N_17955,N_17776,N_17684);
nand U17956 (N_17956,N_17661,N_17764);
nand U17957 (N_17957,N_17751,N_17700);
or U17958 (N_17958,N_17742,N_17727);
nor U17959 (N_17959,N_17773,N_17731);
xnor U17960 (N_17960,N_17634,N_17604);
or U17961 (N_17961,N_17741,N_17662);
nor U17962 (N_17962,N_17732,N_17769);
nor U17963 (N_17963,N_17762,N_17672);
and U17964 (N_17964,N_17707,N_17642);
xor U17965 (N_17965,N_17698,N_17700);
or U17966 (N_17966,N_17709,N_17685);
xor U17967 (N_17967,N_17645,N_17759);
and U17968 (N_17968,N_17767,N_17643);
and U17969 (N_17969,N_17644,N_17764);
nand U17970 (N_17970,N_17758,N_17614);
xnor U17971 (N_17971,N_17632,N_17662);
nand U17972 (N_17972,N_17706,N_17775);
and U17973 (N_17973,N_17734,N_17736);
and U17974 (N_17974,N_17771,N_17796);
or U17975 (N_17975,N_17647,N_17743);
xnor U17976 (N_17976,N_17669,N_17766);
or U17977 (N_17977,N_17758,N_17647);
nand U17978 (N_17978,N_17719,N_17676);
xnor U17979 (N_17979,N_17714,N_17734);
xnor U17980 (N_17980,N_17693,N_17648);
and U17981 (N_17981,N_17614,N_17769);
nand U17982 (N_17982,N_17679,N_17714);
nand U17983 (N_17983,N_17771,N_17713);
nand U17984 (N_17984,N_17775,N_17795);
or U17985 (N_17985,N_17745,N_17774);
xor U17986 (N_17986,N_17766,N_17687);
or U17987 (N_17987,N_17677,N_17779);
or U17988 (N_17988,N_17743,N_17631);
and U17989 (N_17989,N_17661,N_17678);
xor U17990 (N_17990,N_17658,N_17753);
xor U17991 (N_17991,N_17782,N_17787);
and U17992 (N_17992,N_17759,N_17745);
nor U17993 (N_17993,N_17782,N_17670);
and U17994 (N_17994,N_17747,N_17738);
or U17995 (N_17995,N_17628,N_17714);
nand U17996 (N_17996,N_17689,N_17786);
or U17997 (N_17997,N_17693,N_17645);
or U17998 (N_17998,N_17745,N_17638);
nor U17999 (N_17999,N_17679,N_17603);
xor U18000 (N_18000,N_17802,N_17940);
xnor U18001 (N_18001,N_17918,N_17888);
and U18002 (N_18002,N_17810,N_17962);
nor U18003 (N_18003,N_17993,N_17873);
or U18004 (N_18004,N_17970,N_17818);
and U18005 (N_18005,N_17913,N_17956);
nor U18006 (N_18006,N_17891,N_17850);
nor U18007 (N_18007,N_17870,N_17821);
xnor U18008 (N_18008,N_17832,N_17834);
and U18009 (N_18009,N_17883,N_17966);
or U18010 (N_18010,N_17939,N_17841);
nor U18011 (N_18011,N_17866,N_17836);
nor U18012 (N_18012,N_17983,N_17936);
nand U18013 (N_18013,N_17923,N_17961);
or U18014 (N_18014,N_17897,N_17998);
xor U18015 (N_18015,N_17955,N_17909);
and U18016 (N_18016,N_17808,N_17875);
or U18017 (N_18017,N_17819,N_17953);
or U18018 (N_18018,N_17986,N_17858);
nor U18019 (N_18019,N_17839,N_17872);
xnor U18020 (N_18020,N_17964,N_17889);
xor U18021 (N_18021,N_17963,N_17859);
nand U18022 (N_18022,N_17845,N_17843);
and U18023 (N_18023,N_17932,N_17933);
nand U18024 (N_18024,N_17945,N_17924);
or U18025 (N_18025,N_17903,N_17974);
xnor U18026 (N_18026,N_17860,N_17868);
xnor U18027 (N_18027,N_17907,N_17838);
xnor U18028 (N_18028,N_17852,N_17806);
xor U18029 (N_18029,N_17926,N_17977);
nand U18030 (N_18030,N_17823,N_17885);
nand U18031 (N_18031,N_17824,N_17912);
nand U18032 (N_18032,N_17813,N_17865);
and U18033 (N_18033,N_17809,N_17878);
or U18034 (N_18034,N_17816,N_17867);
xnor U18035 (N_18035,N_17895,N_17954);
xor U18036 (N_18036,N_17908,N_17904);
or U18037 (N_18037,N_17893,N_17915);
or U18038 (N_18038,N_17985,N_17864);
nor U18039 (N_18039,N_17959,N_17947);
and U18040 (N_18040,N_17920,N_17944);
or U18041 (N_18041,N_17911,N_17862);
and U18042 (N_18042,N_17822,N_17922);
nand U18043 (N_18043,N_17937,N_17826);
xnor U18044 (N_18044,N_17914,N_17930);
and U18045 (N_18045,N_17842,N_17968);
nor U18046 (N_18046,N_17975,N_17861);
nand U18047 (N_18047,N_17999,N_17951);
and U18048 (N_18048,N_17950,N_17910);
nand U18049 (N_18049,N_17869,N_17890);
xnor U18050 (N_18050,N_17995,N_17902);
nor U18051 (N_18051,N_17887,N_17942);
and U18052 (N_18052,N_17886,N_17803);
or U18053 (N_18053,N_17820,N_17997);
xnor U18054 (N_18054,N_17892,N_17996);
or U18055 (N_18055,N_17840,N_17811);
xnor U18056 (N_18056,N_17805,N_17828);
or U18057 (N_18057,N_17894,N_17934);
nand U18058 (N_18058,N_17880,N_17851);
nand U18059 (N_18059,N_17898,N_17928);
or U18060 (N_18060,N_17978,N_17979);
or U18061 (N_18061,N_17812,N_17849);
nor U18062 (N_18062,N_17877,N_17844);
xnor U18063 (N_18063,N_17817,N_17814);
or U18064 (N_18064,N_17801,N_17971);
and U18065 (N_18065,N_17965,N_17906);
or U18066 (N_18066,N_17921,N_17879);
nand U18067 (N_18067,N_17929,N_17952);
nor U18068 (N_18068,N_17857,N_17871);
nand U18069 (N_18069,N_17854,N_17991);
and U18070 (N_18070,N_17848,N_17882);
nor U18071 (N_18071,N_17946,N_17990);
xnor U18072 (N_18072,N_17927,N_17815);
and U18073 (N_18073,N_17958,N_17896);
and U18074 (N_18074,N_17973,N_17943);
nor U18075 (N_18075,N_17881,N_17957);
nand U18076 (N_18076,N_17941,N_17831);
and U18077 (N_18077,N_17833,N_17960);
nor U18078 (N_18078,N_17948,N_17847);
nor U18079 (N_18079,N_17925,N_17935);
or U18080 (N_18080,N_17876,N_17856);
and U18081 (N_18081,N_17829,N_17807);
nand U18082 (N_18082,N_17835,N_17804);
and U18083 (N_18083,N_17900,N_17949);
or U18084 (N_18084,N_17987,N_17874);
nor U18085 (N_18085,N_17830,N_17931);
nand U18086 (N_18086,N_17899,N_17980);
and U18087 (N_18087,N_17938,N_17919);
or U18088 (N_18088,N_17825,N_17853);
nand U18089 (N_18089,N_17837,N_17901);
and U18090 (N_18090,N_17969,N_17984);
xnor U18091 (N_18091,N_17905,N_17981);
nor U18092 (N_18092,N_17972,N_17989);
nand U18093 (N_18093,N_17994,N_17846);
xor U18094 (N_18094,N_17827,N_17992);
and U18095 (N_18095,N_17976,N_17982);
nand U18096 (N_18096,N_17855,N_17967);
and U18097 (N_18097,N_17917,N_17988);
and U18098 (N_18098,N_17863,N_17916);
and U18099 (N_18099,N_17884,N_17800);
nor U18100 (N_18100,N_17927,N_17867);
xnor U18101 (N_18101,N_17936,N_17871);
xnor U18102 (N_18102,N_17871,N_17876);
or U18103 (N_18103,N_17844,N_17974);
and U18104 (N_18104,N_17933,N_17958);
or U18105 (N_18105,N_17813,N_17936);
and U18106 (N_18106,N_17841,N_17913);
or U18107 (N_18107,N_17984,N_17823);
xnor U18108 (N_18108,N_17820,N_17990);
nor U18109 (N_18109,N_17845,N_17899);
or U18110 (N_18110,N_17986,N_17921);
and U18111 (N_18111,N_17972,N_17817);
xnor U18112 (N_18112,N_17847,N_17995);
nand U18113 (N_18113,N_17882,N_17988);
xnor U18114 (N_18114,N_17881,N_17991);
xnor U18115 (N_18115,N_17900,N_17913);
or U18116 (N_18116,N_17849,N_17866);
and U18117 (N_18117,N_17880,N_17987);
and U18118 (N_18118,N_17803,N_17854);
and U18119 (N_18119,N_17923,N_17865);
and U18120 (N_18120,N_17944,N_17907);
nand U18121 (N_18121,N_17981,N_17976);
nor U18122 (N_18122,N_17896,N_17814);
nand U18123 (N_18123,N_17844,N_17999);
or U18124 (N_18124,N_17932,N_17864);
xnor U18125 (N_18125,N_17994,N_17914);
and U18126 (N_18126,N_17920,N_17800);
and U18127 (N_18127,N_17832,N_17876);
nor U18128 (N_18128,N_17926,N_17941);
xnor U18129 (N_18129,N_17998,N_17999);
and U18130 (N_18130,N_17800,N_17834);
nand U18131 (N_18131,N_17800,N_17885);
or U18132 (N_18132,N_17813,N_17814);
xnor U18133 (N_18133,N_17900,N_17932);
nor U18134 (N_18134,N_17903,N_17855);
xor U18135 (N_18135,N_17888,N_17811);
or U18136 (N_18136,N_17979,N_17838);
nor U18137 (N_18137,N_17840,N_17895);
and U18138 (N_18138,N_17880,N_17897);
xor U18139 (N_18139,N_17949,N_17921);
or U18140 (N_18140,N_17800,N_17973);
nand U18141 (N_18141,N_17948,N_17856);
nand U18142 (N_18142,N_17854,N_17870);
nor U18143 (N_18143,N_17969,N_17875);
and U18144 (N_18144,N_17867,N_17862);
nor U18145 (N_18145,N_17961,N_17990);
and U18146 (N_18146,N_17844,N_17813);
and U18147 (N_18147,N_17850,N_17926);
xnor U18148 (N_18148,N_17854,N_17822);
nand U18149 (N_18149,N_17899,N_17914);
nor U18150 (N_18150,N_17917,N_17848);
nand U18151 (N_18151,N_17865,N_17808);
nor U18152 (N_18152,N_17897,N_17938);
and U18153 (N_18153,N_17943,N_17829);
xnor U18154 (N_18154,N_17837,N_17864);
or U18155 (N_18155,N_17867,N_17814);
and U18156 (N_18156,N_17849,N_17801);
nor U18157 (N_18157,N_17974,N_17898);
xnor U18158 (N_18158,N_17950,N_17845);
nor U18159 (N_18159,N_17993,N_17870);
or U18160 (N_18160,N_17922,N_17950);
nand U18161 (N_18161,N_17851,N_17992);
nand U18162 (N_18162,N_17909,N_17946);
or U18163 (N_18163,N_17971,N_17986);
or U18164 (N_18164,N_17920,N_17975);
nor U18165 (N_18165,N_17969,N_17950);
or U18166 (N_18166,N_17898,N_17968);
nand U18167 (N_18167,N_17801,N_17802);
or U18168 (N_18168,N_17985,N_17999);
or U18169 (N_18169,N_17961,N_17941);
nand U18170 (N_18170,N_17928,N_17957);
nor U18171 (N_18171,N_17856,N_17988);
nor U18172 (N_18172,N_17999,N_17845);
nor U18173 (N_18173,N_17804,N_17803);
nor U18174 (N_18174,N_17938,N_17997);
xor U18175 (N_18175,N_17975,N_17930);
nand U18176 (N_18176,N_17933,N_17925);
and U18177 (N_18177,N_17916,N_17924);
nand U18178 (N_18178,N_17892,N_17891);
nor U18179 (N_18179,N_17976,N_17866);
and U18180 (N_18180,N_17861,N_17815);
or U18181 (N_18181,N_17916,N_17968);
nand U18182 (N_18182,N_17986,N_17938);
nor U18183 (N_18183,N_17877,N_17848);
and U18184 (N_18184,N_17911,N_17914);
and U18185 (N_18185,N_17825,N_17989);
and U18186 (N_18186,N_17881,N_17917);
nor U18187 (N_18187,N_17989,N_17814);
or U18188 (N_18188,N_17914,N_17838);
nor U18189 (N_18189,N_17812,N_17802);
nand U18190 (N_18190,N_17993,N_17932);
nor U18191 (N_18191,N_17984,N_17865);
and U18192 (N_18192,N_17895,N_17929);
or U18193 (N_18193,N_17842,N_17853);
nor U18194 (N_18194,N_17860,N_17869);
or U18195 (N_18195,N_17929,N_17955);
nand U18196 (N_18196,N_17973,N_17995);
and U18197 (N_18197,N_17852,N_17988);
nand U18198 (N_18198,N_17935,N_17955);
and U18199 (N_18199,N_17831,N_17838);
xor U18200 (N_18200,N_18178,N_18075);
nor U18201 (N_18201,N_18017,N_18080);
xor U18202 (N_18202,N_18066,N_18112);
xnor U18203 (N_18203,N_18060,N_18193);
and U18204 (N_18204,N_18123,N_18088);
and U18205 (N_18205,N_18105,N_18086);
and U18206 (N_18206,N_18111,N_18072);
nor U18207 (N_18207,N_18125,N_18037);
xor U18208 (N_18208,N_18108,N_18023);
or U18209 (N_18209,N_18167,N_18002);
xor U18210 (N_18210,N_18093,N_18115);
or U18211 (N_18211,N_18024,N_18149);
and U18212 (N_18212,N_18189,N_18163);
and U18213 (N_18213,N_18106,N_18188);
and U18214 (N_18214,N_18103,N_18031);
nand U18215 (N_18215,N_18034,N_18001);
nand U18216 (N_18216,N_18176,N_18052);
xor U18217 (N_18217,N_18197,N_18107);
or U18218 (N_18218,N_18099,N_18136);
nand U18219 (N_18219,N_18000,N_18113);
or U18220 (N_18220,N_18196,N_18055);
nand U18221 (N_18221,N_18148,N_18076);
nand U18222 (N_18222,N_18137,N_18069);
nor U18223 (N_18223,N_18168,N_18110);
and U18224 (N_18224,N_18121,N_18025);
and U18225 (N_18225,N_18158,N_18128);
xor U18226 (N_18226,N_18179,N_18068);
and U18227 (N_18227,N_18057,N_18170);
xnor U18228 (N_18228,N_18195,N_18028);
nor U18229 (N_18229,N_18180,N_18120);
and U18230 (N_18230,N_18053,N_18114);
and U18231 (N_18231,N_18102,N_18135);
nand U18232 (N_18232,N_18145,N_18150);
and U18233 (N_18233,N_18140,N_18181);
nor U18234 (N_18234,N_18119,N_18008);
xnor U18235 (N_18235,N_18022,N_18154);
nand U18236 (N_18236,N_18071,N_18146);
or U18237 (N_18237,N_18160,N_18094);
or U18238 (N_18238,N_18184,N_18032);
nor U18239 (N_18239,N_18087,N_18147);
and U18240 (N_18240,N_18073,N_18162);
nor U18241 (N_18241,N_18159,N_18046);
xor U18242 (N_18242,N_18132,N_18144);
and U18243 (N_18243,N_18074,N_18062);
xor U18244 (N_18244,N_18141,N_18077);
and U18245 (N_18245,N_18174,N_18139);
xor U18246 (N_18246,N_18127,N_18133);
nor U18247 (N_18247,N_18045,N_18166);
nor U18248 (N_18248,N_18153,N_18011);
nand U18249 (N_18249,N_18117,N_18143);
or U18250 (N_18250,N_18030,N_18157);
nor U18251 (N_18251,N_18047,N_18100);
or U18252 (N_18252,N_18064,N_18005);
or U18253 (N_18253,N_18118,N_18056);
or U18254 (N_18254,N_18039,N_18097);
xor U18255 (N_18255,N_18169,N_18089);
and U18256 (N_18256,N_18186,N_18165);
or U18257 (N_18257,N_18019,N_18182);
nor U18258 (N_18258,N_18003,N_18009);
nand U18259 (N_18259,N_18065,N_18083);
nor U18260 (N_18260,N_18044,N_18026);
nor U18261 (N_18261,N_18092,N_18051);
or U18262 (N_18262,N_18050,N_18126);
nand U18263 (N_18263,N_18177,N_18043);
and U18264 (N_18264,N_18142,N_18063);
nand U18265 (N_18265,N_18067,N_18061);
and U18266 (N_18266,N_18049,N_18035);
nor U18267 (N_18267,N_18007,N_18156);
nand U18268 (N_18268,N_18194,N_18042);
nor U18269 (N_18269,N_18091,N_18109);
nand U18270 (N_18270,N_18048,N_18164);
and U18271 (N_18271,N_18041,N_18172);
xnor U18272 (N_18272,N_18116,N_18014);
nor U18273 (N_18273,N_18015,N_18013);
and U18274 (N_18274,N_18155,N_18130);
nand U18275 (N_18275,N_18151,N_18078);
and U18276 (N_18276,N_18183,N_18198);
or U18277 (N_18277,N_18081,N_18016);
nor U18278 (N_18278,N_18038,N_18058);
nor U18279 (N_18279,N_18098,N_18152);
or U18280 (N_18280,N_18082,N_18090);
xnor U18281 (N_18281,N_18101,N_18079);
and U18282 (N_18282,N_18012,N_18185);
nand U18283 (N_18283,N_18006,N_18173);
nand U18284 (N_18284,N_18040,N_18199);
or U18285 (N_18285,N_18033,N_18054);
and U18286 (N_18286,N_18175,N_18018);
or U18287 (N_18287,N_18010,N_18192);
nand U18288 (N_18288,N_18059,N_18096);
and U18289 (N_18289,N_18191,N_18129);
and U18290 (N_18290,N_18134,N_18027);
nand U18291 (N_18291,N_18124,N_18004);
and U18292 (N_18292,N_18161,N_18095);
nand U18293 (N_18293,N_18122,N_18029);
and U18294 (N_18294,N_18190,N_18021);
nor U18295 (N_18295,N_18085,N_18171);
xnor U18296 (N_18296,N_18138,N_18187);
nor U18297 (N_18297,N_18070,N_18020);
and U18298 (N_18298,N_18036,N_18104);
and U18299 (N_18299,N_18131,N_18084);
or U18300 (N_18300,N_18039,N_18049);
nor U18301 (N_18301,N_18167,N_18175);
xor U18302 (N_18302,N_18041,N_18129);
and U18303 (N_18303,N_18080,N_18028);
xnor U18304 (N_18304,N_18160,N_18115);
nand U18305 (N_18305,N_18112,N_18025);
and U18306 (N_18306,N_18083,N_18148);
or U18307 (N_18307,N_18037,N_18112);
and U18308 (N_18308,N_18020,N_18115);
or U18309 (N_18309,N_18196,N_18164);
nand U18310 (N_18310,N_18005,N_18003);
nor U18311 (N_18311,N_18016,N_18017);
xor U18312 (N_18312,N_18194,N_18187);
nand U18313 (N_18313,N_18121,N_18103);
and U18314 (N_18314,N_18024,N_18121);
nor U18315 (N_18315,N_18064,N_18097);
and U18316 (N_18316,N_18045,N_18056);
nand U18317 (N_18317,N_18030,N_18099);
and U18318 (N_18318,N_18153,N_18064);
nand U18319 (N_18319,N_18015,N_18166);
or U18320 (N_18320,N_18079,N_18136);
nand U18321 (N_18321,N_18097,N_18114);
nor U18322 (N_18322,N_18072,N_18040);
nor U18323 (N_18323,N_18164,N_18096);
or U18324 (N_18324,N_18172,N_18137);
or U18325 (N_18325,N_18021,N_18044);
or U18326 (N_18326,N_18077,N_18086);
or U18327 (N_18327,N_18003,N_18094);
and U18328 (N_18328,N_18170,N_18149);
or U18329 (N_18329,N_18119,N_18006);
or U18330 (N_18330,N_18143,N_18199);
xnor U18331 (N_18331,N_18114,N_18025);
nand U18332 (N_18332,N_18187,N_18140);
nand U18333 (N_18333,N_18135,N_18126);
nand U18334 (N_18334,N_18048,N_18159);
xor U18335 (N_18335,N_18061,N_18154);
xor U18336 (N_18336,N_18123,N_18162);
nor U18337 (N_18337,N_18148,N_18135);
nand U18338 (N_18338,N_18001,N_18020);
or U18339 (N_18339,N_18144,N_18136);
and U18340 (N_18340,N_18075,N_18023);
nand U18341 (N_18341,N_18008,N_18129);
nor U18342 (N_18342,N_18185,N_18101);
or U18343 (N_18343,N_18044,N_18168);
nor U18344 (N_18344,N_18094,N_18146);
or U18345 (N_18345,N_18005,N_18039);
or U18346 (N_18346,N_18158,N_18056);
nor U18347 (N_18347,N_18121,N_18097);
nand U18348 (N_18348,N_18031,N_18122);
nor U18349 (N_18349,N_18120,N_18074);
and U18350 (N_18350,N_18005,N_18131);
or U18351 (N_18351,N_18025,N_18119);
and U18352 (N_18352,N_18071,N_18108);
nand U18353 (N_18353,N_18125,N_18199);
or U18354 (N_18354,N_18075,N_18027);
xor U18355 (N_18355,N_18072,N_18006);
or U18356 (N_18356,N_18177,N_18086);
nor U18357 (N_18357,N_18189,N_18161);
or U18358 (N_18358,N_18184,N_18013);
or U18359 (N_18359,N_18160,N_18025);
nand U18360 (N_18360,N_18080,N_18169);
nand U18361 (N_18361,N_18028,N_18085);
xor U18362 (N_18362,N_18007,N_18046);
nor U18363 (N_18363,N_18063,N_18041);
xnor U18364 (N_18364,N_18188,N_18193);
or U18365 (N_18365,N_18059,N_18035);
and U18366 (N_18366,N_18094,N_18035);
nor U18367 (N_18367,N_18024,N_18134);
xor U18368 (N_18368,N_18170,N_18063);
nor U18369 (N_18369,N_18049,N_18114);
nor U18370 (N_18370,N_18025,N_18188);
nand U18371 (N_18371,N_18160,N_18052);
and U18372 (N_18372,N_18056,N_18001);
and U18373 (N_18373,N_18091,N_18063);
nor U18374 (N_18374,N_18108,N_18073);
xor U18375 (N_18375,N_18128,N_18006);
xnor U18376 (N_18376,N_18086,N_18062);
or U18377 (N_18377,N_18106,N_18136);
nor U18378 (N_18378,N_18050,N_18132);
nor U18379 (N_18379,N_18180,N_18003);
xor U18380 (N_18380,N_18091,N_18115);
and U18381 (N_18381,N_18196,N_18129);
nand U18382 (N_18382,N_18045,N_18115);
nor U18383 (N_18383,N_18154,N_18015);
nor U18384 (N_18384,N_18013,N_18040);
xnor U18385 (N_18385,N_18067,N_18112);
xor U18386 (N_18386,N_18087,N_18002);
nor U18387 (N_18387,N_18124,N_18023);
nand U18388 (N_18388,N_18111,N_18003);
xor U18389 (N_18389,N_18013,N_18176);
xnor U18390 (N_18390,N_18154,N_18043);
or U18391 (N_18391,N_18132,N_18151);
xnor U18392 (N_18392,N_18192,N_18130);
or U18393 (N_18393,N_18147,N_18138);
nor U18394 (N_18394,N_18173,N_18093);
nand U18395 (N_18395,N_18026,N_18076);
nand U18396 (N_18396,N_18150,N_18110);
nand U18397 (N_18397,N_18066,N_18120);
or U18398 (N_18398,N_18100,N_18142);
or U18399 (N_18399,N_18177,N_18166);
nand U18400 (N_18400,N_18237,N_18343);
xnor U18401 (N_18401,N_18247,N_18380);
xor U18402 (N_18402,N_18381,N_18245);
nor U18403 (N_18403,N_18373,N_18383);
nor U18404 (N_18404,N_18352,N_18362);
nand U18405 (N_18405,N_18319,N_18349);
or U18406 (N_18406,N_18332,N_18372);
or U18407 (N_18407,N_18251,N_18266);
or U18408 (N_18408,N_18293,N_18217);
xnor U18409 (N_18409,N_18369,N_18321);
nand U18410 (N_18410,N_18287,N_18370);
or U18411 (N_18411,N_18272,N_18398);
xor U18412 (N_18412,N_18270,N_18258);
nand U18413 (N_18413,N_18225,N_18390);
and U18414 (N_18414,N_18345,N_18221);
nor U18415 (N_18415,N_18214,N_18296);
xnor U18416 (N_18416,N_18213,N_18357);
nor U18417 (N_18417,N_18222,N_18368);
nor U18418 (N_18418,N_18229,N_18291);
and U18419 (N_18419,N_18361,N_18322);
xor U18420 (N_18420,N_18382,N_18252);
xnor U18421 (N_18421,N_18302,N_18391);
and U18422 (N_18422,N_18355,N_18201);
nand U18423 (N_18423,N_18297,N_18348);
nor U18424 (N_18424,N_18277,N_18329);
nand U18425 (N_18425,N_18255,N_18212);
or U18426 (N_18426,N_18261,N_18309);
or U18427 (N_18427,N_18336,N_18315);
xnor U18428 (N_18428,N_18394,N_18310);
and U18429 (N_18429,N_18353,N_18283);
nor U18430 (N_18430,N_18367,N_18338);
or U18431 (N_18431,N_18320,N_18239);
or U18432 (N_18432,N_18275,N_18379);
nand U18433 (N_18433,N_18253,N_18303);
nand U18434 (N_18434,N_18219,N_18334);
nor U18435 (N_18435,N_18215,N_18356);
and U18436 (N_18436,N_18374,N_18265);
xor U18437 (N_18437,N_18350,N_18290);
or U18438 (N_18438,N_18281,N_18318);
and U18439 (N_18439,N_18210,N_18286);
xnor U18440 (N_18440,N_18386,N_18274);
nor U18441 (N_18441,N_18276,N_18347);
xor U18442 (N_18442,N_18388,N_18295);
nor U18443 (N_18443,N_18282,N_18378);
and U18444 (N_18444,N_18260,N_18346);
nor U18445 (N_18445,N_18311,N_18396);
or U18446 (N_18446,N_18335,N_18231);
or U18447 (N_18447,N_18227,N_18244);
nand U18448 (N_18448,N_18366,N_18327);
or U18449 (N_18449,N_18351,N_18220);
or U18450 (N_18450,N_18230,N_18259);
and U18451 (N_18451,N_18326,N_18224);
or U18452 (N_18452,N_18384,N_18228);
and U18453 (N_18453,N_18306,N_18299);
and U18454 (N_18454,N_18284,N_18393);
and U18455 (N_18455,N_18202,N_18337);
nand U18456 (N_18456,N_18360,N_18300);
and U18457 (N_18457,N_18267,N_18389);
xnor U18458 (N_18458,N_18397,N_18278);
and U18459 (N_18459,N_18339,N_18285);
and U18460 (N_18460,N_18371,N_18223);
and U18461 (N_18461,N_18288,N_18200);
and U18462 (N_18462,N_18233,N_18271);
xor U18463 (N_18463,N_18205,N_18387);
xor U18464 (N_18464,N_18280,N_18375);
or U18465 (N_18465,N_18241,N_18279);
nand U18466 (N_18466,N_18323,N_18392);
or U18467 (N_18467,N_18333,N_18257);
nand U18468 (N_18468,N_18208,N_18289);
and U18469 (N_18469,N_18317,N_18324);
or U18470 (N_18470,N_18211,N_18246);
and U18471 (N_18471,N_18363,N_18365);
nor U18472 (N_18472,N_18313,N_18305);
and U18473 (N_18473,N_18236,N_18364);
or U18474 (N_18474,N_18268,N_18294);
or U18475 (N_18475,N_18377,N_18235);
xor U18476 (N_18476,N_18340,N_18248);
and U18477 (N_18477,N_18376,N_18325);
nor U18478 (N_18478,N_18308,N_18312);
nor U18479 (N_18479,N_18354,N_18207);
xnor U18480 (N_18480,N_18232,N_18328);
xor U18481 (N_18481,N_18204,N_18359);
and U18482 (N_18482,N_18216,N_18385);
xnor U18483 (N_18483,N_18307,N_18341);
xnor U18484 (N_18484,N_18331,N_18358);
and U18485 (N_18485,N_18234,N_18330);
xnor U18486 (N_18486,N_18206,N_18395);
and U18487 (N_18487,N_18254,N_18262);
nor U18488 (N_18488,N_18240,N_18218);
nand U18489 (N_18489,N_18264,N_18203);
nand U18490 (N_18490,N_18249,N_18238);
nor U18491 (N_18491,N_18226,N_18304);
and U18492 (N_18492,N_18298,N_18273);
nand U18493 (N_18493,N_18256,N_18316);
xnor U18494 (N_18494,N_18269,N_18209);
nand U18495 (N_18495,N_18342,N_18242);
or U18496 (N_18496,N_18344,N_18263);
or U18497 (N_18497,N_18243,N_18250);
or U18498 (N_18498,N_18301,N_18399);
xor U18499 (N_18499,N_18314,N_18292);
nand U18500 (N_18500,N_18231,N_18207);
or U18501 (N_18501,N_18367,N_18246);
xor U18502 (N_18502,N_18389,N_18377);
xnor U18503 (N_18503,N_18321,N_18296);
and U18504 (N_18504,N_18213,N_18344);
nand U18505 (N_18505,N_18285,N_18212);
or U18506 (N_18506,N_18244,N_18373);
nand U18507 (N_18507,N_18362,N_18321);
nand U18508 (N_18508,N_18394,N_18313);
nor U18509 (N_18509,N_18252,N_18237);
nand U18510 (N_18510,N_18302,N_18394);
nand U18511 (N_18511,N_18223,N_18226);
nor U18512 (N_18512,N_18351,N_18385);
nand U18513 (N_18513,N_18313,N_18277);
nor U18514 (N_18514,N_18381,N_18285);
xnor U18515 (N_18515,N_18257,N_18244);
xor U18516 (N_18516,N_18331,N_18271);
xor U18517 (N_18517,N_18315,N_18318);
or U18518 (N_18518,N_18232,N_18215);
nand U18519 (N_18519,N_18349,N_18220);
and U18520 (N_18520,N_18394,N_18338);
nand U18521 (N_18521,N_18281,N_18388);
nand U18522 (N_18522,N_18316,N_18380);
or U18523 (N_18523,N_18360,N_18229);
nor U18524 (N_18524,N_18223,N_18356);
nand U18525 (N_18525,N_18247,N_18316);
xnor U18526 (N_18526,N_18344,N_18220);
nor U18527 (N_18527,N_18288,N_18380);
or U18528 (N_18528,N_18279,N_18354);
nand U18529 (N_18529,N_18379,N_18292);
nor U18530 (N_18530,N_18368,N_18376);
nor U18531 (N_18531,N_18277,N_18327);
nor U18532 (N_18532,N_18383,N_18371);
nor U18533 (N_18533,N_18334,N_18269);
or U18534 (N_18534,N_18247,N_18212);
nor U18535 (N_18535,N_18258,N_18335);
nand U18536 (N_18536,N_18334,N_18339);
nor U18537 (N_18537,N_18253,N_18206);
nand U18538 (N_18538,N_18369,N_18249);
nand U18539 (N_18539,N_18280,N_18392);
nand U18540 (N_18540,N_18205,N_18288);
nand U18541 (N_18541,N_18223,N_18296);
nand U18542 (N_18542,N_18373,N_18266);
and U18543 (N_18543,N_18318,N_18213);
and U18544 (N_18544,N_18396,N_18210);
or U18545 (N_18545,N_18331,N_18349);
nand U18546 (N_18546,N_18282,N_18239);
nor U18547 (N_18547,N_18351,N_18344);
and U18548 (N_18548,N_18260,N_18365);
or U18549 (N_18549,N_18329,N_18394);
and U18550 (N_18550,N_18312,N_18357);
or U18551 (N_18551,N_18389,N_18309);
nand U18552 (N_18552,N_18396,N_18381);
nor U18553 (N_18553,N_18287,N_18232);
xnor U18554 (N_18554,N_18373,N_18387);
and U18555 (N_18555,N_18390,N_18241);
or U18556 (N_18556,N_18218,N_18290);
nor U18557 (N_18557,N_18399,N_18308);
nand U18558 (N_18558,N_18225,N_18206);
nand U18559 (N_18559,N_18268,N_18290);
nor U18560 (N_18560,N_18342,N_18207);
nand U18561 (N_18561,N_18244,N_18251);
nand U18562 (N_18562,N_18377,N_18211);
nor U18563 (N_18563,N_18224,N_18225);
nor U18564 (N_18564,N_18372,N_18256);
xor U18565 (N_18565,N_18251,N_18221);
xnor U18566 (N_18566,N_18272,N_18311);
or U18567 (N_18567,N_18208,N_18344);
and U18568 (N_18568,N_18312,N_18258);
xnor U18569 (N_18569,N_18388,N_18245);
nor U18570 (N_18570,N_18227,N_18382);
nor U18571 (N_18571,N_18241,N_18225);
and U18572 (N_18572,N_18387,N_18320);
and U18573 (N_18573,N_18354,N_18305);
xor U18574 (N_18574,N_18315,N_18223);
nand U18575 (N_18575,N_18352,N_18348);
and U18576 (N_18576,N_18385,N_18271);
or U18577 (N_18577,N_18201,N_18367);
xnor U18578 (N_18578,N_18375,N_18349);
nand U18579 (N_18579,N_18327,N_18236);
xor U18580 (N_18580,N_18318,N_18329);
and U18581 (N_18581,N_18343,N_18313);
nor U18582 (N_18582,N_18341,N_18306);
or U18583 (N_18583,N_18201,N_18235);
nor U18584 (N_18584,N_18276,N_18250);
or U18585 (N_18585,N_18322,N_18300);
nand U18586 (N_18586,N_18380,N_18344);
or U18587 (N_18587,N_18280,N_18385);
or U18588 (N_18588,N_18209,N_18346);
nand U18589 (N_18589,N_18365,N_18353);
xnor U18590 (N_18590,N_18231,N_18319);
xor U18591 (N_18591,N_18320,N_18210);
nand U18592 (N_18592,N_18208,N_18395);
xnor U18593 (N_18593,N_18266,N_18378);
nor U18594 (N_18594,N_18321,N_18378);
nor U18595 (N_18595,N_18248,N_18225);
nand U18596 (N_18596,N_18342,N_18259);
or U18597 (N_18597,N_18288,N_18316);
xor U18598 (N_18598,N_18275,N_18340);
nand U18599 (N_18599,N_18285,N_18203);
and U18600 (N_18600,N_18563,N_18522);
xor U18601 (N_18601,N_18469,N_18453);
nor U18602 (N_18602,N_18535,N_18533);
nor U18603 (N_18603,N_18579,N_18582);
nor U18604 (N_18604,N_18449,N_18450);
xor U18605 (N_18605,N_18452,N_18519);
nor U18606 (N_18606,N_18425,N_18442);
xor U18607 (N_18607,N_18546,N_18521);
or U18608 (N_18608,N_18551,N_18571);
or U18609 (N_18609,N_18495,N_18426);
or U18610 (N_18610,N_18524,N_18544);
or U18611 (N_18611,N_18508,N_18494);
xor U18612 (N_18612,N_18467,N_18411);
nand U18613 (N_18613,N_18470,N_18481);
xnor U18614 (N_18614,N_18594,N_18417);
and U18615 (N_18615,N_18457,N_18593);
or U18616 (N_18616,N_18488,N_18576);
or U18617 (N_18617,N_18447,N_18473);
nand U18618 (N_18618,N_18413,N_18460);
or U18619 (N_18619,N_18486,N_18574);
nor U18620 (N_18620,N_18402,N_18439);
nor U18621 (N_18621,N_18503,N_18557);
and U18622 (N_18622,N_18572,N_18536);
xor U18623 (N_18623,N_18548,N_18419);
nor U18624 (N_18624,N_18479,N_18553);
nand U18625 (N_18625,N_18578,N_18584);
xor U18626 (N_18626,N_18545,N_18491);
xor U18627 (N_18627,N_18547,N_18566);
or U18628 (N_18628,N_18400,N_18554);
or U18629 (N_18629,N_18454,N_18527);
and U18630 (N_18630,N_18575,N_18513);
or U18631 (N_18631,N_18592,N_18543);
or U18632 (N_18632,N_18461,N_18430);
and U18633 (N_18633,N_18423,N_18562);
xnor U18634 (N_18634,N_18504,N_18529);
and U18635 (N_18635,N_18506,N_18583);
xnor U18636 (N_18636,N_18466,N_18534);
or U18637 (N_18637,N_18532,N_18525);
nor U18638 (N_18638,N_18483,N_18518);
and U18639 (N_18639,N_18478,N_18500);
and U18640 (N_18640,N_18586,N_18451);
or U18641 (N_18641,N_18496,N_18493);
and U18642 (N_18642,N_18565,N_18590);
nand U18643 (N_18643,N_18403,N_18597);
xnor U18644 (N_18644,N_18427,N_18437);
xor U18645 (N_18645,N_18404,N_18541);
or U18646 (N_18646,N_18502,N_18538);
nor U18647 (N_18647,N_18581,N_18591);
nor U18648 (N_18648,N_18509,N_18462);
and U18649 (N_18649,N_18421,N_18511);
xnor U18650 (N_18650,N_18596,N_18599);
or U18651 (N_18651,N_18580,N_18490);
nor U18652 (N_18652,N_18415,N_18589);
and U18653 (N_18653,N_18487,N_18418);
nor U18654 (N_18654,N_18409,N_18528);
or U18655 (N_18655,N_18540,N_18468);
xnor U18656 (N_18656,N_18505,N_18492);
nand U18657 (N_18657,N_18420,N_18514);
xor U18658 (N_18658,N_18595,N_18448);
or U18659 (N_18659,N_18577,N_18560);
and U18660 (N_18660,N_18407,N_18432);
xor U18661 (N_18661,N_18414,N_18559);
xnor U18662 (N_18662,N_18556,N_18550);
nand U18663 (N_18663,N_18598,N_18477);
xnor U18664 (N_18664,N_18520,N_18440);
and U18665 (N_18665,N_18446,N_18474);
or U18666 (N_18666,N_18498,N_18424);
or U18667 (N_18667,N_18489,N_18501);
nand U18668 (N_18668,N_18438,N_18515);
and U18669 (N_18669,N_18416,N_18433);
and U18670 (N_18670,N_18549,N_18537);
nor U18671 (N_18671,N_18441,N_18431);
xnor U18672 (N_18672,N_18434,N_18480);
xnor U18673 (N_18673,N_18526,N_18463);
nand U18674 (N_18674,N_18499,N_18435);
or U18675 (N_18675,N_18471,N_18507);
nor U18676 (N_18676,N_18482,N_18542);
nor U18677 (N_18677,N_18570,N_18476);
or U18678 (N_18678,N_18568,N_18401);
xnor U18679 (N_18679,N_18429,N_18485);
nand U18680 (N_18680,N_18475,N_18585);
xor U18681 (N_18681,N_18567,N_18444);
nor U18682 (N_18682,N_18558,N_18569);
xnor U18683 (N_18683,N_18465,N_18464);
nand U18684 (N_18684,N_18564,N_18408);
xnor U18685 (N_18685,N_18456,N_18587);
nor U18686 (N_18686,N_18517,N_18552);
or U18687 (N_18687,N_18561,N_18436);
and U18688 (N_18688,N_18539,N_18458);
nand U18689 (N_18689,N_18555,N_18588);
xnor U18690 (N_18690,N_18422,N_18405);
xnor U18691 (N_18691,N_18516,N_18530);
nand U18692 (N_18692,N_18573,N_18497);
and U18693 (N_18693,N_18428,N_18443);
nor U18694 (N_18694,N_18472,N_18523);
nand U18695 (N_18695,N_18531,N_18459);
xor U18696 (N_18696,N_18512,N_18412);
nor U18697 (N_18697,N_18455,N_18410);
or U18698 (N_18698,N_18484,N_18406);
nor U18699 (N_18699,N_18510,N_18445);
nand U18700 (N_18700,N_18582,N_18500);
nand U18701 (N_18701,N_18498,N_18479);
nand U18702 (N_18702,N_18455,N_18544);
or U18703 (N_18703,N_18434,N_18441);
nor U18704 (N_18704,N_18549,N_18433);
and U18705 (N_18705,N_18504,N_18448);
and U18706 (N_18706,N_18571,N_18567);
xor U18707 (N_18707,N_18473,N_18538);
nor U18708 (N_18708,N_18514,N_18423);
nand U18709 (N_18709,N_18492,N_18571);
or U18710 (N_18710,N_18448,N_18512);
nor U18711 (N_18711,N_18550,N_18511);
and U18712 (N_18712,N_18540,N_18450);
xnor U18713 (N_18713,N_18516,N_18559);
or U18714 (N_18714,N_18587,N_18534);
or U18715 (N_18715,N_18424,N_18428);
and U18716 (N_18716,N_18565,N_18406);
nor U18717 (N_18717,N_18567,N_18468);
nand U18718 (N_18718,N_18570,N_18506);
xor U18719 (N_18719,N_18440,N_18487);
xor U18720 (N_18720,N_18407,N_18557);
nand U18721 (N_18721,N_18419,N_18583);
and U18722 (N_18722,N_18458,N_18576);
xor U18723 (N_18723,N_18527,N_18445);
or U18724 (N_18724,N_18577,N_18599);
nor U18725 (N_18725,N_18590,N_18419);
xor U18726 (N_18726,N_18495,N_18550);
nor U18727 (N_18727,N_18527,N_18512);
and U18728 (N_18728,N_18410,N_18413);
or U18729 (N_18729,N_18585,N_18459);
nor U18730 (N_18730,N_18465,N_18400);
or U18731 (N_18731,N_18412,N_18555);
or U18732 (N_18732,N_18454,N_18531);
and U18733 (N_18733,N_18405,N_18548);
nand U18734 (N_18734,N_18474,N_18558);
and U18735 (N_18735,N_18417,N_18531);
xnor U18736 (N_18736,N_18540,N_18511);
and U18737 (N_18737,N_18464,N_18507);
and U18738 (N_18738,N_18556,N_18553);
or U18739 (N_18739,N_18576,N_18438);
nor U18740 (N_18740,N_18445,N_18438);
or U18741 (N_18741,N_18481,N_18450);
and U18742 (N_18742,N_18457,N_18486);
and U18743 (N_18743,N_18484,N_18530);
nand U18744 (N_18744,N_18545,N_18540);
nand U18745 (N_18745,N_18555,N_18516);
nand U18746 (N_18746,N_18553,N_18598);
nand U18747 (N_18747,N_18488,N_18544);
nor U18748 (N_18748,N_18596,N_18568);
xor U18749 (N_18749,N_18509,N_18546);
xnor U18750 (N_18750,N_18584,N_18492);
nor U18751 (N_18751,N_18472,N_18465);
nand U18752 (N_18752,N_18543,N_18433);
xnor U18753 (N_18753,N_18427,N_18477);
and U18754 (N_18754,N_18474,N_18584);
nor U18755 (N_18755,N_18543,N_18546);
nor U18756 (N_18756,N_18427,N_18508);
xor U18757 (N_18757,N_18472,N_18458);
nor U18758 (N_18758,N_18434,N_18495);
nand U18759 (N_18759,N_18430,N_18554);
nand U18760 (N_18760,N_18572,N_18491);
nand U18761 (N_18761,N_18521,N_18591);
nor U18762 (N_18762,N_18414,N_18468);
or U18763 (N_18763,N_18582,N_18419);
or U18764 (N_18764,N_18446,N_18408);
nand U18765 (N_18765,N_18500,N_18455);
xor U18766 (N_18766,N_18463,N_18510);
nor U18767 (N_18767,N_18489,N_18586);
nor U18768 (N_18768,N_18449,N_18461);
xnor U18769 (N_18769,N_18509,N_18587);
nand U18770 (N_18770,N_18522,N_18503);
nand U18771 (N_18771,N_18426,N_18453);
nand U18772 (N_18772,N_18511,N_18534);
or U18773 (N_18773,N_18499,N_18437);
nor U18774 (N_18774,N_18425,N_18510);
nand U18775 (N_18775,N_18553,N_18454);
xnor U18776 (N_18776,N_18487,N_18411);
xor U18777 (N_18777,N_18519,N_18529);
or U18778 (N_18778,N_18477,N_18507);
nor U18779 (N_18779,N_18494,N_18582);
or U18780 (N_18780,N_18532,N_18417);
or U18781 (N_18781,N_18544,N_18424);
xnor U18782 (N_18782,N_18420,N_18571);
or U18783 (N_18783,N_18403,N_18408);
nor U18784 (N_18784,N_18562,N_18542);
or U18785 (N_18785,N_18520,N_18425);
and U18786 (N_18786,N_18596,N_18484);
nand U18787 (N_18787,N_18494,N_18554);
nand U18788 (N_18788,N_18510,N_18451);
nor U18789 (N_18789,N_18561,N_18532);
xor U18790 (N_18790,N_18406,N_18530);
nand U18791 (N_18791,N_18598,N_18437);
nand U18792 (N_18792,N_18444,N_18473);
nand U18793 (N_18793,N_18459,N_18419);
or U18794 (N_18794,N_18499,N_18576);
nor U18795 (N_18795,N_18541,N_18424);
nor U18796 (N_18796,N_18496,N_18548);
xnor U18797 (N_18797,N_18507,N_18520);
and U18798 (N_18798,N_18460,N_18542);
xor U18799 (N_18799,N_18476,N_18401);
or U18800 (N_18800,N_18683,N_18769);
xor U18801 (N_18801,N_18775,N_18681);
nor U18802 (N_18802,N_18640,N_18666);
nand U18803 (N_18803,N_18672,N_18607);
xor U18804 (N_18804,N_18773,N_18653);
and U18805 (N_18805,N_18747,N_18776);
nor U18806 (N_18806,N_18600,N_18734);
nand U18807 (N_18807,N_18788,N_18667);
xnor U18808 (N_18808,N_18620,N_18657);
xor U18809 (N_18809,N_18625,N_18652);
and U18810 (N_18810,N_18619,N_18665);
xnor U18811 (N_18811,N_18694,N_18750);
or U18812 (N_18812,N_18799,N_18705);
or U18813 (N_18813,N_18612,N_18648);
nand U18814 (N_18814,N_18678,N_18797);
nand U18815 (N_18815,N_18616,N_18757);
and U18816 (N_18816,N_18661,N_18738);
xor U18817 (N_18817,N_18703,N_18767);
and U18818 (N_18818,N_18635,N_18763);
and U18819 (N_18819,N_18634,N_18723);
xor U18820 (N_18820,N_18755,N_18772);
nor U18821 (N_18821,N_18742,N_18671);
or U18822 (N_18822,N_18670,N_18736);
nor U18823 (N_18823,N_18646,N_18631);
xnor U18824 (N_18824,N_18602,N_18785);
nand U18825 (N_18825,N_18614,N_18752);
nor U18826 (N_18826,N_18641,N_18761);
nor U18827 (N_18827,N_18690,N_18730);
nand U18828 (N_18828,N_18603,N_18676);
and U18829 (N_18829,N_18731,N_18695);
and U18830 (N_18830,N_18726,N_18724);
nand U18831 (N_18831,N_18748,N_18664);
nor U18832 (N_18832,N_18781,N_18786);
or U18833 (N_18833,N_18768,N_18706);
nor U18834 (N_18834,N_18624,N_18792);
nor U18835 (N_18835,N_18649,N_18718);
nor U18836 (N_18836,N_18692,N_18639);
nor U18837 (N_18837,N_18746,N_18774);
xor U18838 (N_18838,N_18674,N_18693);
or U18839 (N_18839,N_18709,N_18663);
xnor U18840 (N_18840,N_18778,N_18754);
or U18841 (N_18841,N_18659,N_18737);
nor U18842 (N_18842,N_18739,N_18711);
or U18843 (N_18843,N_18637,N_18662);
xor U18844 (N_18844,N_18629,N_18656);
and U18845 (N_18845,N_18712,N_18698);
or U18846 (N_18846,N_18708,N_18735);
xnor U18847 (N_18847,N_18762,N_18604);
nand U18848 (N_18848,N_18759,N_18744);
nor U18849 (N_18849,N_18725,N_18645);
nand U18850 (N_18850,N_18721,N_18771);
nand U18851 (N_18851,N_18655,N_18633);
nand U18852 (N_18852,N_18675,N_18700);
nor U18853 (N_18853,N_18621,N_18686);
nor U18854 (N_18854,N_18701,N_18796);
or U18855 (N_18855,N_18784,N_18627);
or U18856 (N_18856,N_18651,N_18765);
nand U18857 (N_18857,N_18642,N_18687);
xnor U18858 (N_18858,N_18688,N_18668);
and U18859 (N_18859,N_18715,N_18791);
nand U18860 (N_18860,N_18628,N_18780);
nand U18861 (N_18861,N_18719,N_18632);
xnor U18862 (N_18862,N_18766,N_18793);
nor U18863 (N_18863,N_18689,N_18606);
or U18864 (N_18864,N_18758,N_18751);
or U18865 (N_18865,N_18722,N_18704);
or U18866 (N_18866,N_18608,N_18720);
xor U18867 (N_18867,N_18605,N_18729);
nand U18868 (N_18868,N_18611,N_18623);
and U18869 (N_18869,N_18601,N_18647);
nor U18870 (N_18870,N_18696,N_18743);
or U18871 (N_18871,N_18669,N_18626);
and U18872 (N_18872,N_18702,N_18679);
nor U18873 (N_18873,N_18677,N_18764);
xor U18874 (N_18874,N_18787,N_18717);
nor U18875 (N_18875,N_18610,N_18691);
nand U18876 (N_18876,N_18697,N_18795);
and U18877 (N_18877,N_18617,N_18749);
xnor U18878 (N_18878,N_18733,N_18745);
and U18879 (N_18879,N_18714,N_18622);
and U18880 (N_18880,N_18789,N_18732);
or U18881 (N_18881,N_18760,N_18613);
nor U18882 (N_18882,N_18756,N_18636);
nand U18883 (N_18883,N_18658,N_18770);
nor U18884 (N_18884,N_18777,N_18716);
nor U18885 (N_18885,N_18680,N_18713);
nand U18886 (N_18886,N_18782,N_18740);
and U18887 (N_18887,N_18710,N_18790);
xor U18888 (N_18888,N_18618,N_18654);
or U18889 (N_18889,N_18609,N_18699);
or U18890 (N_18890,N_18673,N_18727);
nand U18891 (N_18891,N_18630,N_18644);
or U18892 (N_18892,N_18753,N_18783);
xor U18893 (N_18893,N_18650,N_18615);
xor U18894 (N_18894,N_18638,N_18779);
or U18895 (N_18895,N_18794,N_18707);
xor U18896 (N_18896,N_18660,N_18741);
xor U18897 (N_18897,N_18643,N_18728);
and U18898 (N_18898,N_18682,N_18798);
nand U18899 (N_18899,N_18685,N_18684);
or U18900 (N_18900,N_18677,N_18656);
xnor U18901 (N_18901,N_18683,N_18626);
and U18902 (N_18902,N_18749,N_18629);
xnor U18903 (N_18903,N_18664,N_18747);
xor U18904 (N_18904,N_18652,N_18716);
nand U18905 (N_18905,N_18780,N_18736);
or U18906 (N_18906,N_18760,N_18631);
or U18907 (N_18907,N_18728,N_18744);
nor U18908 (N_18908,N_18714,N_18628);
xnor U18909 (N_18909,N_18632,N_18646);
nand U18910 (N_18910,N_18740,N_18628);
nand U18911 (N_18911,N_18785,N_18711);
and U18912 (N_18912,N_18658,N_18796);
and U18913 (N_18913,N_18758,N_18791);
nand U18914 (N_18914,N_18616,N_18791);
and U18915 (N_18915,N_18759,N_18798);
xnor U18916 (N_18916,N_18776,N_18761);
nor U18917 (N_18917,N_18772,N_18624);
nand U18918 (N_18918,N_18774,N_18625);
xnor U18919 (N_18919,N_18792,N_18604);
nor U18920 (N_18920,N_18779,N_18709);
and U18921 (N_18921,N_18684,N_18648);
nand U18922 (N_18922,N_18634,N_18734);
or U18923 (N_18923,N_18794,N_18698);
or U18924 (N_18924,N_18773,N_18667);
or U18925 (N_18925,N_18697,N_18682);
xor U18926 (N_18926,N_18637,N_18782);
nand U18927 (N_18927,N_18731,N_18691);
and U18928 (N_18928,N_18629,N_18611);
xor U18929 (N_18929,N_18694,N_18669);
and U18930 (N_18930,N_18709,N_18696);
nor U18931 (N_18931,N_18794,N_18795);
nand U18932 (N_18932,N_18653,N_18695);
or U18933 (N_18933,N_18749,N_18667);
xnor U18934 (N_18934,N_18682,N_18720);
and U18935 (N_18935,N_18648,N_18652);
and U18936 (N_18936,N_18662,N_18743);
and U18937 (N_18937,N_18797,N_18649);
xnor U18938 (N_18938,N_18669,N_18649);
xor U18939 (N_18939,N_18611,N_18716);
nor U18940 (N_18940,N_18731,N_18767);
and U18941 (N_18941,N_18679,N_18633);
nor U18942 (N_18942,N_18793,N_18674);
xor U18943 (N_18943,N_18645,N_18651);
or U18944 (N_18944,N_18759,N_18739);
nor U18945 (N_18945,N_18722,N_18789);
and U18946 (N_18946,N_18697,N_18662);
nand U18947 (N_18947,N_18730,N_18793);
xor U18948 (N_18948,N_18782,N_18607);
xor U18949 (N_18949,N_18772,N_18717);
or U18950 (N_18950,N_18748,N_18708);
and U18951 (N_18951,N_18676,N_18695);
and U18952 (N_18952,N_18713,N_18668);
nand U18953 (N_18953,N_18643,N_18724);
or U18954 (N_18954,N_18693,N_18787);
nor U18955 (N_18955,N_18694,N_18778);
xnor U18956 (N_18956,N_18756,N_18740);
and U18957 (N_18957,N_18689,N_18679);
or U18958 (N_18958,N_18771,N_18675);
or U18959 (N_18959,N_18706,N_18617);
or U18960 (N_18960,N_18675,N_18627);
or U18961 (N_18961,N_18748,N_18732);
or U18962 (N_18962,N_18789,N_18758);
or U18963 (N_18963,N_18748,N_18730);
xor U18964 (N_18964,N_18772,N_18656);
nand U18965 (N_18965,N_18697,N_18750);
nor U18966 (N_18966,N_18660,N_18665);
or U18967 (N_18967,N_18677,N_18711);
xor U18968 (N_18968,N_18685,N_18619);
nor U18969 (N_18969,N_18792,N_18633);
xor U18970 (N_18970,N_18603,N_18766);
nor U18971 (N_18971,N_18751,N_18745);
nor U18972 (N_18972,N_18674,N_18682);
xnor U18973 (N_18973,N_18781,N_18792);
nand U18974 (N_18974,N_18603,N_18688);
or U18975 (N_18975,N_18735,N_18722);
and U18976 (N_18976,N_18783,N_18796);
xnor U18977 (N_18977,N_18635,N_18621);
xnor U18978 (N_18978,N_18682,N_18698);
nand U18979 (N_18979,N_18727,N_18623);
xor U18980 (N_18980,N_18698,N_18755);
xor U18981 (N_18981,N_18776,N_18764);
nand U18982 (N_18982,N_18693,N_18728);
xnor U18983 (N_18983,N_18665,N_18760);
nand U18984 (N_18984,N_18754,N_18798);
nor U18985 (N_18985,N_18617,N_18707);
and U18986 (N_18986,N_18621,N_18752);
or U18987 (N_18987,N_18646,N_18660);
and U18988 (N_18988,N_18684,N_18755);
nor U18989 (N_18989,N_18768,N_18623);
or U18990 (N_18990,N_18604,N_18799);
nor U18991 (N_18991,N_18698,N_18766);
or U18992 (N_18992,N_18773,N_18675);
and U18993 (N_18993,N_18722,N_18733);
or U18994 (N_18994,N_18652,N_18671);
xor U18995 (N_18995,N_18636,N_18650);
and U18996 (N_18996,N_18649,N_18602);
nor U18997 (N_18997,N_18646,N_18712);
and U18998 (N_18998,N_18788,N_18698);
nor U18999 (N_18999,N_18659,N_18600);
or U19000 (N_19000,N_18983,N_18859);
nor U19001 (N_19001,N_18911,N_18829);
nand U19002 (N_19002,N_18955,N_18995);
nand U19003 (N_19003,N_18979,N_18866);
nor U19004 (N_19004,N_18969,N_18971);
or U19005 (N_19005,N_18894,N_18906);
and U19006 (N_19006,N_18813,N_18949);
nand U19007 (N_19007,N_18895,N_18918);
or U19008 (N_19008,N_18831,N_18824);
nor U19009 (N_19009,N_18963,N_18939);
xor U19010 (N_19010,N_18820,N_18899);
nor U19011 (N_19011,N_18986,N_18893);
xor U19012 (N_19012,N_18881,N_18830);
nor U19013 (N_19013,N_18970,N_18960);
or U19014 (N_19014,N_18966,N_18817);
nand U19015 (N_19015,N_18946,N_18961);
nor U19016 (N_19016,N_18887,N_18844);
nand U19017 (N_19017,N_18974,N_18815);
and U19018 (N_19018,N_18801,N_18802);
and U19019 (N_19019,N_18822,N_18948);
nor U19020 (N_19020,N_18843,N_18807);
nand U19021 (N_19021,N_18838,N_18953);
nor U19022 (N_19022,N_18922,N_18929);
or U19023 (N_19023,N_18886,N_18851);
nand U19024 (N_19024,N_18996,N_18848);
xnor U19025 (N_19025,N_18908,N_18913);
and U19026 (N_19026,N_18898,N_18823);
nor U19027 (N_19027,N_18873,N_18855);
nor U19028 (N_19028,N_18883,N_18840);
nor U19029 (N_19029,N_18858,N_18988);
and U19030 (N_19030,N_18880,N_18919);
and U19031 (N_19031,N_18806,N_18834);
nor U19032 (N_19032,N_18984,N_18944);
or U19033 (N_19033,N_18885,N_18910);
nand U19034 (N_19034,N_18932,N_18805);
and U19035 (N_19035,N_18941,N_18933);
nand U19036 (N_19036,N_18942,N_18863);
and U19037 (N_19037,N_18846,N_18987);
or U19038 (N_19038,N_18874,N_18990);
xnor U19039 (N_19039,N_18818,N_18812);
and U19040 (N_19040,N_18965,N_18950);
and U19041 (N_19041,N_18957,N_18958);
nand U19042 (N_19042,N_18900,N_18839);
or U19043 (N_19043,N_18860,N_18867);
or U19044 (N_19044,N_18803,N_18884);
or U19045 (N_19045,N_18879,N_18833);
nand U19046 (N_19046,N_18915,N_18973);
or U19047 (N_19047,N_18861,N_18976);
and U19048 (N_19048,N_18964,N_18914);
or U19049 (N_19049,N_18977,N_18877);
xor U19050 (N_19050,N_18980,N_18865);
or U19051 (N_19051,N_18892,N_18821);
nand U19052 (N_19052,N_18917,N_18875);
nand U19053 (N_19053,N_18921,N_18954);
xnor U19054 (N_19054,N_18937,N_18841);
or U19055 (N_19055,N_18835,N_18854);
xnor U19056 (N_19056,N_18907,N_18901);
and U19057 (N_19057,N_18868,N_18999);
nand U19058 (N_19058,N_18940,N_18943);
and U19059 (N_19059,N_18897,N_18952);
and U19060 (N_19060,N_18998,N_18808);
xnor U19061 (N_19061,N_18928,N_18945);
and U19062 (N_19062,N_18850,N_18967);
nor U19063 (N_19063,N_18981,N_18853);
or U19064 (N_19064,N_18878,N_18920);
nor U19065 (N_19065,N_18982,N_18814);
nand U19066 (N_19066,N_18852,N_18916);
xor U19067 (N_19067,N_18889,N_18876);
xnor U19068 (N_19068,N_18902,N_18827);
and U19069 (N_19069,N_18997,N_18882);
xnor U19070 (N_19070,N_18819,N_18804);
and U19071 (N_19071,N_18968,N_18930);
xor U19072 (N_19072,N_18828,N_18993);
or U19073 (N_19073,N_18869,N_18951);
or U19074 (N_19074,N_18978,N_18959);
nand U19075 (N_19075,N_18912,N_18836);
xnor U19076 (N_19076,N_18924,N_18862);
xor U19077 (N_19077,N_18856,N_18809);
and U19078 (N_19078,N_18832,N_18934);
xnor U19079 (N_19079,N_18925,N_18904);
xnor U19080 (N_19080,N_18888,N_18896);
nand U19081 (N_19081,N_18936,N_18926);
and U19082 (N_19082,N_18962,N_18956);
xor U19083 (N_19083,N_18857,N_18972);
or U19084 (N_19084,N_18864,N_18903);
nor U19085 (N_19085,N_18931,N_18870);
and U19086 (N_19086,N_18810,N_18842);
nor U19087 (N_19087,N_18816,N_18800);
nand U19088 (N_19088,N_18891,N_18905);
or U19089 (N_19089,N_18872,N_18923);
nand U19090 (N_19090,N_18890,N_18927);
nor U19091 (N_19091,N_18837,N_18985);
nor U19092 (N_19092,N_18811,N_18849);
nor U19093 (N_19093,N_18847,N_18909);
or U19094 (N_19094,N_18938,N_18935);
nand U19095 (N_19095,N_18947,N_18994);
or U19096 (N_19096,N_18871,N_18991);
xor U19097 (N_19097,N_18826,N_18845);
nor U19098 (N_19098,N_18975,N_18992);
and U19099 (N_19099,N_18989,N_18825);
nand U19100 (N_19100,N_18818,N_18822);
nor U19101 (N_19101,N_18815,N_18868);
nor U19102 (N_19102,N_18880,N_18865);
or U19103 (N_19103,N_18808,N_18996);
nand U19104 (N_19104,N_18972,N_18936);
or U19105 (N_19105,N_18824,N_18901);
or U19106 (N_19106,N_18903,N_18894);
xnor U19107 (N_19107,N_18879,N_18849);
or U19108 (N_19108,N_18900,N_18996);
nor U19109 (N_19109,N_18897,N_18930);
nor U19110 (N_19110,N_18816,N_18890);
and U19111 (N_19111,N_18808,N_18827);
nand U19112 (N_19112,N_18910,N_18956);
or U19113 (N_19113,N_18971,N_18937);
or U19114 (N_19114,N_18963,N_18816);
and U19115 (N_19115,N_18963,N_18837);
and U19116 (N_19116,N_18972,N_18959);
nand U19117 (N_19117,N_18843,N_18887);
or U19118 (N_19118,N_18931,N_18926);
or U19119 (N_19119,N_18808,N_18982);
xor U19120 (N_19120,N_18982,N_18962);
and U19121 (N_19121,N_18991,N_18962);
nor U19122 (N_19122,N_18907,N_18816);
nor U19123 (N_19123,N_18862,N_18994);
or U19124 (N_19124,N_18887,N_18868);
or U19125 (N_19125,N_18945,N_18989);
or U19126 (N_19126,N_18940,N_18993);
nor U19127 (N_19127,N_18955,N_18829);
nand U19128 (N_19128,N_18823,N_18828);
xor U19129 (N_19129,N_18828,N_18892);
or U19130 (N_19130,N_18969,N_18807);
and U19131 (N_19131,N_18985,N_18845);
xor U19132 (N_19132,N_18959,N_18970);
and U19133 (N_19133,N_18844,N_18903);
nand U19134 (N_19134,N_18848,N_18902);
nand U19135 (N_19135,N_18878,N_18950);
and U19136 (N_19136,N_18908,N_18866);
xor U19137 (N_19137,N_18971,N_18987);
or U19138 (N_19138,N_18998,N_18894);
and U19139 (N_19139,N_18950,N_18900);
nor U19140 (N_19140,N_18820,N_18888);
and U19141 (N_19141,N_18823,N_18839);
nand U19142 (N_19142,N_18970,N_18806);
nor U19143 (N_19143,N_18941,N_18919);
nor U19144 (N_19144,N_18853,N_18813);
nand U19145 (N_19145,N_18929,N_18940);
xor U19146 (N_19146,N_18943,N_18893);
or U19147 (N_19147,N_18835,N_18978);
nor U19148 (N_19148,N_18898,N_18860);
xnor U19149 (N_19149,N_18976,N_18906);
nand U19150 (N_19150,N_18940,N_18904);
nand U19151 (N_19151,N_18976,N_18886);
nand U19152 (N_19152,N_18916,N_18837);
or U19153 (N_19153,N_18872,N_18880);
and U19154 (N_19154,N_18857,N_18934);
xor U19155 (N_19155,N_18819,N_18852);
nor U19156 (N_19156,N_18906,N_18940);
and U19157 (N_19157,N_18999,N_18972);
nor U19158 (N_19158,N_18974,N_18825);
or U19159 (N_19159,N_18948,N_18960);
or U19160 (N_19160,N_18975,N_18859);
and U19161 (N_19161,N_18871,N_18839);
nand U19162 (N_19162,N_18948,N_18923);
nand U19163 (N_19163,N_18937,N_18864);
xor U19164 (N_19164,N_18906,N_18802);
and U19165 (N_19165,N_18993,N_18994);
xnor U19166 (N_19166,N_18830,N_18895);
nand U19167 (N_19167,N_18809,N_18904);
nand U19168 (N_19168,N_18946,N_18993);
nor U19169 (N_19169,N_18986,N_18938);
xor U19170 (N_19170,N_18930,N_18801);
and U19171 (N_19171,N_18837,N_18842);
and U19172 (N_19172,N_18936,N_18881);
or U19173 (N_19173,N_18848,N_18917);
xor U19174 (N_19174,N_18854,N_18999);
nor U19175 (N_19175,N_18983,N_18889);
xnor U19176 (N_19176,N_18983,N_18982);
nand U19177 (N_19177,N_18833,N_18958);
xor U19178 (N_19178,N_18834,N_18879);
nor U19179 (N_19179,N_18950,N_18936);
and U19180 (N_19180,N_18971,N_18963);
xor U19181 (N_19181,N_18987,N_18801);
xor U19182 (N_19182,N_18893,N_18886);
and U19183 (N_19183,N_18869,N_18931);
and U19184 (N_19184,N_18873,N_18879);
and U19185 (N_19185,N_18869,N_18989);
xor U19186 (N_19186,N_18913,N_18836);
and U19187 (N_19187,N_18822,N_18913);
and U19188 (N_19188,N_18914,N_18871);
nor U19189 (N_19189,N_18823,N_18879);
and U19190 (N_19190,N_18943,N_18970);
nand U19191 (N_19191,N_18950,N_18824);
or U19192 (N_19192,N_18980,N_18949);
and U19193 (N_19193,N_18989,N_18835);
xnor U19194 (N_19194,N_18916,N_18848);
nand U19195 (N_19195,N_18818,N_18842);
nand U19196 (N_19196,N_18885,N_18867);
nor U19197 (N_19197,N_18973,N_18841);
xnor U19198 (N_19198,N_18825,N_18884);
nor U19199 (N_19199,N_18888,N_18983);
xnor U19200 (N_19200,N_19070,N_19185);
nand U19201 (N_19201,N_19167,N_19138);
or U19202 (N_19202,N_19121,N_19170);
xnor U19203 (N_19203,N_19193,N_19106);
nand U19204 (N_19204,N_19110,N_19089);
nand U19205 (N_19205,N_19096,N_19151);
nor U19206 (N_19206,N_19149,N_19018);
or U19207 (N_19207,N_19086,N_19124);
nor U19208 (N_19208,N_19159,N_19144);
nand U19209 (N_19209,N_19067,N_19126);
nand U19210 (N_19210,N_19156,N_19006);
or U19211 (N_19211,N_19190,N_19194);
or U19212 (N_19212,N_19094,N_19078);
nor U19213 (N_19213,N_19036,N_19040);
nor U19214 (N_19214,N_19035,N_19174);
and U19215 (N_19215,N_19184,N_19157);
and U19216 (N_19216,N_19058,N_19047);
nor U19217 (N_19217,N_19196,N_19063);
or U19218 (N_19218,N_19111,N_19177);
nand U19219 (N_19219,N_19007,N_19175);
or U19220 (N_19220,N_19188,N_19142);
xnor U19221 (N_19221,N_19033,N_19164);
xnor U19222 (N_19222,N_19137,N_19066);
and U19223 (N_19223,N_19139,N_19163);
or U19224 (N_19224,N_19060,N_19014);
xnor U19225 (N_19225,N_19002,N_19027);
nor U19226 (N_19226,N_19038,N_19088);
nor U19227 (N_19227,N_19198,N_19084);
and U19228 (N_19228,N_19025,N_19054);
or U19229 (N_19229,N_19081,N_19039);
xor U19230 (N_19230,N_19132,N_19012);
xnor U19231 (N_19231,N_19104,N_19001);
nor U19232 (N_19232,N_19133,N_19152);
nor U19233 (N_19233,N_19055,N_19011);
and U19234 (N_19234,N_19093,N_19010);
or U19235 (N_19235,N_19071,N_19135);
and U19236 (N_19236,N_19119,N_19082);
or U19237 (N_19237,N_19136,N_19087);
and U19238 (N_19238,N_19048,N_19125);
nor U19239 (N_19239,N_19034,N_19160);
nand U19240 (N_19240,N_19107,N_19015);
nor U19241 (N_19241,N_19155,N_19130);
and U19242 (N_19242,N_19145,N_19100);
nor U19243 (N_19243,N_19113,N_19148);
and U19244 (N_19244,N_19032,N_19189);
nor U19245 (N_19245,N_19024,N_19114);
nand U19246 (N_19246,N_19052,N_19168);
or U19247 (N_19247,N_19091,N_19154);
nand U19248 (N_19248,N_19069,N_19150);
xor U19249 (N_19249,N_19080,N_19097);
nand U19250 (N_19250,N_19109,N_19068);
and U19251 (N_19251,N_19076,N_19192);
nand U19252 (N_19252,N_19199,N_19090);
xor U19253 (N_19253,N_19073,N_19045);
xor U19254 (N_19254,N_19146,N_19179);
and U19255 (N_19255,N_19083,N_19044);
and U19256 (N_19256,N_19131,N_19072);
or U19257 (N_19257,N_19161,N_19061);
and U19258 (N_19258,N_19005,N_19178);
nor U19259 (N_19259,N_19122,N_19141);
or U19260 (N_19260,N_19103,N_19013);
or U19261 (N_19261,N_19117,N_19108);
and U19262 (N_19262,N_19105,N_19147);
or U19263 (N_19263,N_19056,N_19112);
and U19264 (N_19264,N_19099,N_19102);
xor U19265 (N_19265,N_19059,N_19028);
and U19266 (N_19266,N_19127,N_19030);
nor U19267 (N_19267,N_19016,N_19075);
nand U19268 (N_19268,N_19004,N_19043);
or U19269 (N_19269,N_19162,N_19128);
and U19270 (N_19270,N_19116,N_19165);
xnor U19271 (N_19271,N_19023,N_19051);
xnor U19272 (N_19272,N_19031,N_19022);
and U19273 (N_19273,N_19003,N_19197);
nand U19274 (N_19274,N_19008,N_19079);
and U19275 (N_19275,N_19158,N_19118);
and U19276 (N_19276,N_19021,N_19101);
nor U19277 (N_19277,N_19049,N_19098);
xnor U19278 (N_19278,N_19172,N_19092);
nand U19279 (N_19279,N_19077,N_19134);
nor U19280 (N_19280,N_19000,N_19053);
nand U19281 (N_19281,N_19062,N_19176);
xnor U19282 (N_19282,N_19166,N_19095);
nor U19283 (N_19283,N_19129,N_19041);
nor U19284 (N_19284,N_19064,N_19115);
xnor U19285 (N_19285,N_19173,N_19120);
and U19286 (N_19286,N_19046,N_19181);
or U19287 (N_19287,N_19187,N_19019);
xnor U19288 (N_19288,N_19182,N_19074);
nand U19289 (N_19289,N_19029,N_19171);
nand U19290 (N_19290,N_19042,N_19026);
or U19291 (N_19291,N_19085,N_19037);
xor U19292 (N_19292,N_19195,N_19153);
or U19293 (N_19293,N_19020,N_19169);
nor U19294 (N_19294,N_19180,N_19191);
xor U19295 (N_19295,N_19143,N_19050);
and U19296 (N_19296,N_19009,N_19140);
and U19297 (N_19297,N_19017,N_19183);
nand U19298 (N_19298,N_19057,N_19065);
and U19299 (N_19299,N_19186,N_19123);
and U19300 (N_19300,N_19139,N_19061);
and U19301 (N_19301,N_19018,N_19091);
or U19302 (N_19302,N_19075,N_19098);
and U19303 (N_19303,N_19184,N_19051);
xnor U19304 (N_19304,N_19160,N_19142);
nand U19305 (N_19305,N_19144,N_19026);
nor U19306 (N_19306,N_19007,N_19041);
or U19307 (N_19307,N_19013,N_19021);
or U19308 (N_19308,N_19180,N_19129);
and U19309 (N_19309,N_19149,N_19113);
nor U19310 (N_19310,N_19184,N_19193);
and U19311 (N_19311,N_19059,N_19112);
or U19312 (N_19312,N_19160,N_19052);
and U19313 (N_19313,N_19013,N_19037);
and U19314 (N_19314,N_19099,N_19071);
nor U19315 (N_19315,N_19116,N_19125);
xor U19316 (N_19316,N_19047,N_19082);
or U19317 (N_19317,N_19129,N_19007);
or U19318 (N_19318,N_19135,N_19060);
and U19319 (N_19319,N_19033,N_19143);
or U19320 (N_19320,N_19139,N_19160);
or U19321 (N_19321,N_19025,N_19153);
and U19322 (N_19322,N_19059,N_19173);
nor U19323 (N_19323,N_19194,N_19047);
or U19324 (N_19324,N_19083,N_19127);
and U19325 (N_19325,N_19017,N_19106);
and U19326 (N_19326,N_19169,N_19131);
nand U19327 (N_19327,N_19186,N_19116);
and U19328 (N_19328,N_19125,N_19153);
or U19329 (N_19329,N_19034,N_19056);
and U19330 (N_19330,N_19088,N_19025);
and U19331 (N_19331,N_19046,N_19062);
nand U19332 (N_19332,N_19041,N_19019);
and U19333 (N_19333,N_19108,N_19170);
nand U19334 (N_19334,N_19116,N_19023);
xor U19335 (N_19335,N_19059,N_19131);
nor U19336 (N_19336,N_19069,N_19196);
xor U19337 (N_19337,N_19175,N_19034);
nand U19338 (N_19338,N_19111,N_19191);
xor U19339 (N_19339,N_19111,N_19145);
nand U19340 (N_19340,N_19095,N_19106);
nand U19341 (N_19341,N_19194,N_19022);
or U19342 (N_19342,N_19170,N_19017);
and U19343 (N_19343,N_19094,N_19020);
nor U19344 (N_19344,N_19131,N_19181);
xnor U19345 (N_19345,N_19073,N_19168);
nor U19346 (N_19346,N_19180,N_19025);
nor U19347 (N_19347,N_19040,N_19129);
nor U19348 (N_19348,N_19081,N_19122);
and U19349 (N_19349,N_19143,N_19025);
or U19350 (N_19350,N_19058,N_19084);
xor U19351 (N_19351,N_19009,N_19016);
nand U19352 (N_19352,N_19102,N_19087);
nand U19353 (N_19353,N_19169,N_19128);
xor U19354 (N_19354,N_19107,N_19192);
or U19355 (N_19355,N_19167,N_19050);
nor U19356 (N_19356,N_19122,N_19132);
xnor U19357 (N_19357,N_19149,N_19163);
and U19358 (N_19358,N_19097,N_19075);
xnor U19359 (N_19359,N_19093,N_19001);
or U19360 (N_19360,N_19040,N_19126);
xnor U19361 (N_19361,N_19152,N_19190);
xor U19362 (N_19362,N_19179,N_19093);
nor U19363 (N_19363,N_19023,N_19126);
nor U19364 (N_19364,N_19108,N_19023);
nor U19365 (N_19365,N_19080,N_19167);
nor U19366 (N_19366,N_19111,N_19192);
nand U19367 (N_19367,N_19169,N_19177);
nand U19368 (N_19368,N_19195,N_19185);
or U19369 (N_19369,N_19125,N_19122);
nand U19370 (N_19370,N_19058,N_19017);
xnor U19371 (N_19371,N_19092,N_19197);
or U19372 (N_19372,N_19041,N_19073);
and U19373 (N_19373,N_19163,N_19193);
nor U19374 (N_19374,N_19168,N_19104);
and U19375 (N_19375,N_19060,N_19183);
or U19376 (N_19376,N_19023,N_19190);
xnor U19377 (N_19377,N_19088,N_19137);
nor U19378 (N_19378,N_19024,N_19160);
nor U19379 (N_19379,N_19198,N_19097);
and U19380 (N_19380,N_19183,N_19098);
and U19381 (N_19381,N_19144,N_19132);
nand U19382 (N_19382,N_19043,N_19093);
and U19383 (N_19383,N_19168,N_19183);
nor U19384 (N_19384,N_19100,N_19047);
nand U19385 (N_19385,N_19145,N_19093);
nor U19386 (N_19386,N_19166,N_19010);
nand U19387 (N_19387,N_19160,N_19121);
nand U19388 (N_19388,N_19179,N_19149);
or U19389 (N_19389,N_19005,N_19184);
nor U19390 (N_19390,N_19159,N_19139);
and U19391 (N_19391,N_19028,N_19115);
or U19392 (N_19392,N_19192,N_19172);
or U19393 (N_19393,N_19058,N_19041);
nor U19394 (N_19394,N_19096,N_19191);
or U19395 (N_19395,N_19123,N_19163);
xnor U19396 (N_19396,N_19068,N_19175);
nand U19397 (N_19397,N_19074,N_19051);
and U19398 (N_19398,N_19131,N_19040);
and U19399 (N_19399,N_19101,N_19110);
and U19400 (N_19400,N_19238,N_19274);
and U19401 (N_19401,N_19252,N_19282);
xor U19402 (N_19402,N_19255,N_19295);
nand U19403 (N_19403,N_19325,N_19305);
xor U19404 (N_19404,N_19259,N_19234);
nor U19405 (N_19405,N_19390,N_19283);
and U19406 (N_19406,N_19268,N_19276);
and U19407 (N_19407,N_19351,N_19289);
nand U19408 (N_19408,N_19243,N_19270);
xor U19409 (N_19409,N_19303,N_19288);
nand U19410 (N_19410,N_19329,N_19235);
xnor U19411 (N_19411,N_19229,N_19355);
nand U19412 (N_19412,N_19218,N_19375);
nor U19413 (N_19413,N_19396,N_19300);
and U19414 (N_19414,N_19308,N_19392);
nor U19415 (N_19415,N_19393,N_19226);
nand U19416 (N_19416,N_19333,N_19233);
nor U19417 (N_19417,N_19379,N_19328);
nand U19418 (N_19418,N_19382,N_19315);
nand U19419 (N_19419,N_19262,N_19241);
or U19420 (N_19420,N_19245,N_19373);
and U19421 (N_19421,N_19266,N_19299);
nor U19422 (N_19422,N_19251,N_19365);
and U19423 (N_19423,N_19261,N_19369);
and U19424 (N_19424,N_19247,N_19356);
and U19425 (N_19425,N_19391,N_19237);
nand U19426 (N_19426,N_19254,N_19310);
or U19427 (N_19427,N_19334,N_19381);
nor U19428 (N_19428,N_19219,N_19336);
and U19429 (N_19429,N_19368,N_19264);
nand U19430 (N_19430,N_19222,N_19389);
or U19431 (N_19431,N_19388,N_19347);
nor U19432 (N_19432,N_19385,N_19367);
xnor U19433 (N_19433,N_19284,N_19285);
nor U19434 (N_19434,N_19205,N_19338);
and U19435 (N_19435,N_19204,N_19397);
nor U19436 (N_19436,N_19395,N_19387);
nand U19437 (N_19437,N_19307,N_19217);
nand U19438 (N_19438,N_19230,N_19281);
or U19439 (N_19439,N_19380,N_19249);
nor U19440 (N_19440,N_19220,N_19386);
and U19441 (N_19441,N_19311,N_19231);
nand U19442 (N_19442,N_19265,N_19340);
xor U19443 (N_19443,N_19312,N_19203);
and U19444 (N_19444,N_19363,N_19248);
nor U19445 (N_19445,N_19236,N_19301);
or U19446 (N_19446,N_19313,N_19354);
and U19447 (N_19447,N_19263,N_19292);
nor U19448 (N_19448,N_19349,N_19215);
and U19449 (N_19449,N_19346,N_19319);
nand U19450 (N_19450,N_19257,N_19240);
and U19451 (N_19451,N_19366,N_19232);
nor U19452 (N_19452,N_19309,N_19250);
and U19453 (N_19453,N_19253,N_19214);
and U19454 (N_19454,N_19374,N_19370);
nand U19455 (N_19455,N_19362,N_19302);
nor U19456 (N_19456,N_19296,N_19353);
nor U19457 (N_19457,N_19225,N_19271);
nand U19458 (N_19458,N_19260,N_19398);
xor U19459 (N_19459,N_19364,N_19201);
and U19460 (N_19460,N_19213,N_19286);
nor U19461 (N_19461,N_19272,N_19343);
nand U19462 (N_19462,N_19297,N_19287);
nand U19463 (N_19463,N_19377,N_19208);
xor U19464 (N_19464,N_19280,N_19357);
nor U19465 (N_19465,N_19290,N_19337);
nor U19466 (N_19466,N_19332,N_19202);
nand U19467 (N_19467,N_19314,N_19335);
nand U19468 (N_19468,N_19242,N_19275);
xnor U19469 (N_19469,N_19216,N_19360);
or U19470 (N_19470,N_19206,N_19352);
xnor U19471 (N_19471,N_19378,N_19239);
nand U19472 (N_19472,N_19223,N_19298);
nor U19473 (N_19473,N_19359,N_19269);
nor U19474 (N_19474,N_19372,N_19318);
xor U19475 (N_19475,N_19256,N_19345);
nand U19476 (N_19476,N_19321,N_19350);
and U19477 (N_19477,N_19330,N_19294);
or U19478 (N_19478,N_19291,N_19323);
nor U19479 (N_19479,N_19324,N_19399);
nor U19480 (N_19480,N_19279,N_19246);
xnor U19481 (N_19481,N_19227,N_19224);
nand U19482 (N_19482,N_19212,N_19383);
nor U19483 (N_19483,N_19339,N_19244);
and U19484 (N_19484,N_19293,N_19273);
nand U19485 (N_19485,N_19207,N_19384);
or U19486 (N_19486,N_19394,N_19278);
nand U19487 (N_19487,N_19200,N_19371);
and U19488 (N_19488,N_19306,N_19376);
or U19489 (N_19489,N_19228,N_19331);
or U19490 (N_19490,N_19304,N_19327);
nand U19491 (N_19491,N_19342,N_19317);
or U19492 (N_19492,N_19322,N_19209);
nand U19493 (N_19493,N_19210,N_19341);
nor U19494 (N_19494,N_19258,N_19361);
and U19495 (N_19495,N_19221,N_19277);
nor U19496 (N_19496,N_19316,N_19320);
and U19497 (N_19497,N_19358,N_19326);
xor U19498 (N_19498,N_19348,N_19344);
xnor U19499 (N_19499,N_19211,N_19267);
and U19500 (N_19500,N_19295,N_19341);
and U19501 (N_19501,N_19265,N_19234);
and U19502 (N_19502,N_19256,N_19297);
and U19503 (N_19503,N_19268,N_19267);
and U19504 (N_19504,N_19343,N_19296);
xnor U19505 (N_19505,N_19278,N_19352);
nor U19506 (N_19506,N_19232,N_19221);
and U19507 (N_19507,N_19352,N_19395);
nor U19508 (N_19508,N_19349,N_19234);
nor U19509 (N_19509,N_19219,N_19243);
nand U19510 (N_19510,N_19302,N_19330);
or U19511 (N_19511,N_19201,N_19207);
or U19512 (N_19512,N_19347,N_19326);
or U19513 (N_19513,N_19225,N_19252);
and U19514 (N_19514,N_19312,N_19398);
or U19515 (N_19515,N_19379,N_19384);
and U19516 (N_19516,N_19318,N_19361);
xor U19517 (N_19517,N_19251,N_19382);
xnor U19518 (N_19518,N_19358,N_19204);
and U19519 (N_19519,N_19284,N_19273);
nor U19520 (N_19520,N_19215,N_19354);
nand U19521 (N_19521,N_19246,N_19294);
or U19522 (N_19522,N_19394,N_19395);
xnor U19523 (N_19523,N_19392,N_19379);
xnor U19524 (N_19524,N_19346,N_19314);
xnor U19525 (N_19525,N_19258,N_19327);
xor U19526 (N_19526,N_19317,N_19216);
nor U19527 (N_19527,N_19207,N_19217);
nor U19528 (N_19528,N_19334,N_19321);
xnor U19529 (N_19529,N_19218,N_19308);
nand U19530 (N_19530,N_19208,N_19354);
or U19531 (N_19531,N_19316,N_19236);
nand U19532 (N_19532,N_19343,N_19380);
nand U19533 (N_19533,N_19200,N_19318);
nand U19534 (N_19534,N_19332,N_19388);
nor U19535 (N_19535,N_19207,N_19321);
xor U19536 (N_19536,N_19362,N_19369);
nand U19537 (N_19537,N_19333,N_19293);
and U19538 (N_19538,N_19270,N_19288);
xor U19539 (N_19539,N_19232,N_19395);
or U19540 (N_19540,N_19308,N_19278);
or U19541 (N_19541,N_19354,N_19271);
xor U19542 (N_19542,N_19208,N_19322);
or U19543 (N_19543,N_19214,N_19297);
and U19544 (N_19544,N_19318,N_19294);
or U19545 (N_19545,N_19336,N_19368);
xnor U19546 (N_19546,N_19342,N_19257);
nand U19547 (N_19547,N_19395,N_19205);
or U19548 (N_19548,N_19351,N_19332);
or U19549 (N_19549,N_19330,N_19251);
nor U19550 (N_19550,N_19228,N_19259);
xnor U19551 (N_19551,N_19314,N_19316);
and U19552 (N_19552,N_19237,N_19212);
xnor U19553 (N_19553,N_19377,N_19202);
nor U19554 (N_19554,N_19260,N_19345);
and U19555 (N_19555,N_19315,N_19326);
xor U19556 (N_19556,N_19292,N_19348);
nand U19557 (N_19557,N_19368,N_19265);
xor U19558 (N_19558,N_19205,N_19321);
xnor U19559 (N_19559,N_19326,N_19255);
nand U19560 (N_19560,N_19346,N_19304);
or U19561 (N_19561,N_19392,N_19233);
nor U19562 (N_19562,N_19287,N_19385);
and U19563 (N_19563,N_19339,N_19393);
xor U19564 (N_19564,N_19253,N_19231);
xnor U19565 (N_19565,N_19344,N_19354);
and U19566 (N_19566,N_19277,N_19256);
and U19567 (N_19567,N_19301,N_19231);
or U19568 (N_19568,N_19354,N_19259);
or U19569 (N_19569,N_19358,N_19214);
nand U19570 (N_19570,N_19314,N_19365);
or U19571 (N_19571,N_19380,N_19251);
nor U19572 (N_19572,N_19358,N_19391);
nand U19573 (N_19573,N_19357,N_19382);
nor U19574 (N_19574,N_19214,N_19327);
nand U19575 (N_19575,N_19216,N_19331);
xor U19576 (N_19576,N_19201,N_19297);
and U19577 (N_19577,N_19216,N_19320);
nor U19578 (N_19578,N_19220,N_19227);
nand U19579 (N_19579,N_19285,N_19392);
nand U19580 (N_19580,N_19266,N_19281);
xor U19581 (N_19581,N_19379,N_19353);
nor U19582 (N_19582,N_19392,N_19335);
or U19583 (N_19583,N_19278,N_19232);
nor U19584 (N_19584,N_19205,N_19203);
and U19585 (N_19585,N_19397,N_19335);
or U19586 (N_19586,N_19238,N_19398);
xor U19587 (N_19587,N_19339,N_19341);
or U19588 (N_19588,N_19293,N_19255);
xnor U19589 (N_19589,N_19354,N_19296);
or U19590 (N_19590,N_19379,N_19372);
nand U19591 (N_19591,N_19258,N_19394);
xor U19592 (N_19592,N_19300,N_19376);
and U19593 (N_19593,N_19384,N_19263);
nand U19594 (N_19594,N_19392,N_19223);
and U19595 (N_19595,N_19351,N_19207);
nand U19596 (N_19596,N_19283,N_19205);
nand U19597 (N_19597,N_19303,N_19247);
nor U19598 (N_19598,N_19365,N_19239);
nand U19599 (N_19599,N_19370,N_19229);
nand U19600 (N_19600,N_19560,N_19430);
or U19601 (N_19601,N_19444,N_19594);
or U19602 (N_19602,N_19402,N_19565);
or U19603 (N_19603,N_19581,N_19432);
or U19604 (N_19604,N_19544,N_19591);
nand U19605 (N_19605,N_19470,N_19448);
or U19606 (N_19606,N_19519,N_19436);
nand U19607 (N_19607,N_19445,N_19529);
nand U19608 (N_19608,N_19408,N_19439);
nor U19609 (N_19609,N_19466,N_19468);
nor U19610 (N_19610,N_19597,N_19458);
and U19611 (N_19611,N_19593,N_19542);
and U19612 (N_19612,N_19473,N_19481);
or U19613 (N_19613,N_19434,N_19440);
nand U19614 (N_19614,N_19454,N_19487);
nor U19615 (N_19615,N_19475,N_19412);
or U19616 (N_19616,N_19512,N_19419);
xor U19617 (N_19617,N_19451,N_19404);
xor U19618 (N_19618,N_19462,N_19520);
and U19619 (N_19619,N_19596,N_19514);
nor U19620 (N_19620,N_19447,N_19450);
nand U19621 (N_19621,N_19546,N_19584);
nand U19622 (N_19622,N_19522,N_19428);
or U19623 (N_19623,N_19575,N_19425);
nor U19624 (N_19624,N_19401,N_19421);
and U19625 (N_19625,N_19513,N_19505);
or U19626 (N_19626,N_19536,N_19477);
nand U19627 (N_19627,N_19453,N_19469);
nor U19628 (N_19628,N_19442,N_19443);
and U19629 (N_19629,N_19526,N_19449);
nor U19630 (N_19630,N_19418,N_19543);
and U19631 (N_19631,N_19472,N_19535);
or U19632 (N_19632,N_19501,N_19496);
nand U19633 (N_19633,N_19456,N_19463);
xnor U19634 (N_19634,N_19485,N_19518);
or U19635 (N_19635,N_19564,N_19574);
nand U19636 (N_19636,N_19455,N_19476);
xor U19637 (N_19637,N_19504,N_19493);
and U19638 (N_19638,N_19499,N_19530);
nor U19639 (N_19639,N_19561,N_19480);
or U19640 (N_19640,N_19557,N_19461);
nor U19641 (N_19641,N_19527,N_19427);
or U19642 (N_19642,N_19559,N_19503);
nand U19643 (N_19643,N_19416,N_19435);
xnor U19644 (N_19644,N_19558,N_19488);
and U19645 (N_19645,N_19516,N_19467);
nand U19646 (N_19646,N_19531,N_19506);
or U19647 (N_19647,N_19414,N_19491);
xor U19648 (N_19648,N_19452,N_19573);
and U19649 (N_19649,N_19465,N_19484);
and U19650 (N_19650,N_19563,N_19511);
and U19651 (N_19651,N_19579,N_19406);
and U19652 (N_19652,N_19423,N_19552);
xor U19653 (N_19653,N_19409,N_19599);
and U19654 (N_19654,N_19583,N_19495);
or U19655 (N_19655,N_19545,N_19494);
or U19656 (N_19656,N_19403,N_19437);
xnor U19657 (N_19657,N_19515,N_19420);
and U19658 (N_19658,N_19464,N_19407);
nand U19659 (N_19659,N_19582,N_19478);
xor U19660 (N_19660,N_19566,N_19446);
and U19661 (N_19661,N_19497,N_19482);
or U19662 (N_19662,N_19433,N_19441);
and U19663 (N_19663,N_19571,N_19498);
nor U19664 (N_19664,N_19509,N_19576);
or U19665 (N_19665,N_19417,N_19474);
and U19666 (N_19666,N_19580,N_19490);
nor U19667 (N_19667,N_19424,N_19537);
xnor U19668 (N_19668,N_19556,N_19521);
xnor U19669 (N_19669,N_19567,N_19569);
xor U19670 (N_19670,N_19460,N_19562);
or U19671 (N_19671,N_19479,N_19534);
or U19672 (N_19672,N_19525,N_19570);
or U19673 (N_19673,N_19429,N_19410);
nor U19674 (N_19674,N_19538,N_19587);
nor U19675 (N_19675,N_19411,N_19532);
nor U19676 (N_19676,N_19551,N_19595);
nand U19677 (N_19677,N_19426,N_19589);
or U19678 (N_19678,N_19549,N_19510);
xnor U19679 (N_19679,N_19586,N_19486);
nand U19680 (N_19680,N_19598,N_19492);
nand U19681 (N_19681,N_19502,N_19524);
or U19682 (N_19682,N_19568,N_19539);
nand U19683 (N_19683,N_19541,N_19459);
nor U19684 (N_19684,N_19523,N_19500);
nor U19685 (N_19685,N_19471,N_19431);
or U19686 (N_19686,N_19438,N_19577);
and U19687 (N_19687,N_19548,N_19588);
nand U19688 (N_19688,N_19508,N_19540);
and U19689 (N_19689,N_19554,N_19550);
and U19690 (N_19690,N_19400,N_19413);
xor U19691 (N_19691,N_19457,N_19405);
or U19692 (N_19692,N_19415,N_19555);
or U19693 (N_19693,N_19507,N_19590);
nor U19694 (N_19694,N_19572,N_19533);
xor U19695 (N_19695,N_19422,N_19553);
xor U19696 (N_19696,N_19547,N_19517);
nand U19697 (N_19697,N_19489,N_19585);
xnor U19698 (N_19698,N_19528,N_19483);
xnor U19699 (N_19699,N_19578,N_19592);
nand U19700 (N_19700,N_19565,N_19430);
nand U19701 (N_19701,N_19430,N_19499);
nor U19702 (N_19702,N_19440,N_19597);
nor U19703 (N_19703,N_19597,N_19420);
nand U19704 (N_19704,N_19553,N_19424);
xor U19705 (N_19705,N_19568,N_19407);
and U19706 (N_19706,N_19575,N_19592);
xnor U19707 (N_19707,N_19581,N_19475);
nor U19708 (N_19708,N_19489,N_19567);
and U19709 (N_19709,N_19469,N_19555);
nor U19710 (N_19710,N_19559,N_19556);
xor U19711 (N_19711,N_19489,N_19441);
and U19712 (N_19712,N_19530,N_19529);
xor U19713 (N_19713,N_19461,N_19492);
and U19714 (N_19714,N_19457,N_19477);
nor U19715 (N_19715,N_19561,N_19588);
or U19716 (N_19716,N_19475,N_19454);
nor U19717 (N_19717,N_19406,N_19423);
nor U19718 (N_19718,N_19515,N_19517);
nor U19719 (N_19719,N_19413,N_19586);
or U19720 (N_19720,N_19573,N_19506);
xor U19721 (N_19721,N_19461,N_19489);
and U19722 (N_19722,N_19559,N_19406);
nor U19723 (N_19723,N_19465,N_19492);
and U19724 (N_19724,N_19501,N_19441);
xor U19725 (N_19725,N_19409,N_19548);
nand U19726 (N_19726,N_19559,N_19588);
xnor U19727 (N_19727,N_19447,N_19410);
xor U19728 (N_19728,N_19447,N_19412);
nand U19729 (N_19729,N_19409,N_19567);
nor U19730 (N_19730,N_19439,N_19537);
or U19731 (N_19731,N_19488,N_19506);
nor U19732 (N_19732,N_19569,N_19556);
nand U19733 (N_19733,N_19470,N_19550);
nor U19734 (N_19734,N_19548,N_19401);
nor U19735 (N_19735,N_19500,N_19517);
and U19736 (N_19736,N_19462,N_19565);
nor U19737 (N_19737,N_19466,N_19583);
nor U19738 (N_19738,N_19590,N_19504);
nand U19739 (N_19739,N_19518,N_19476);
or U19740 (N_19740,N_19475,N_19408);
nor U19741 (N_19741,N_19457,N_19508);
xnor U19742 (N_19742,N_19567,N_19552);
xor U19743 (N_19743,N_19576,N_19408);
or U19744 (N_19744,N_19582,N_19458);
or U19745 (N_19745,N_19497,N_19500);
nor U19746 (N_19746,N_19568,N_19472);
xor U19747 (N_19747,N_19459,N_19561);
nor U19748 (N_19748,N_19457,N_19441);
and U19749 (N_19749,N_19562,N_19479);
nor U19750 (N_19750,N_19534,N_19408);
nor U19751 (N_19751,N_19478,N_19481);
or U19752 (N_19752,N_19469,N_19458);
xor U19753 (N_19753,N_19464,N_19460);
nor U19754 (N_19754,N_19580,N_19543);
xnor U19755 (N_19755,N_19438,N_19523);
or U19756 (N_19756,N_19405,N_19567);
nor U19757 (N_19757,N_19441,N_19537);
and U19758 (N_19758,N_19451,N_19579);
and U19759 (N_19759,N_19448,N_19450);
nand U19760 (N_19760,N_19539,N_19476);
and U19761 (N_19761,N_19548,N_19421);
xor U19762 (N_19762,N_19477,N_19581);
xnor U19763 (N_19763,N_19454,N_19575);
xor U19764 (N_19764,N_19427,N_19583);
or U19765 (N_19765,N_19422,N_19532);
or U19766 (N_19766,N_19414,N_19400);
or U19767 (N_19767,N_19556,N_19405);
nor U19768 (N_19768,N_19438,N_19582);
and U19769 (N_19769,N_19526,N_19542);
nor U19770 (N_19770,N_19419,N_19475);
xnor U19771 (N_19771,N_19510,N_19420);
and U19772 (N_19772,N_19552,N_19527);
or U19773 (N_19773,N_19522,N_19469);
xnor U19774 (N_19774,N_19451,N_19547);
and U19775 (N_19775,N_19507,N_19479);
xor U19776 (N_19776,N_19497,N_19452);
nor U19777 (N_19777,N_19400,N_19436);
nand U19778 (N_19778,N_19496,N_19483);
nor U19779 (N_19779,N_19459,N_19434);
nor U19780 (N_19780,N_19504,N_19453);
or U19781 (N_19781,N_19448,N_19512);
xnor U19782 (N_19782,N_19519,N_19477);
nor U19783 (N_19783,N_19512,N_19478);
xnor U19784 (N_19784,N_19541,N_19439);
nor U19785 (N_19785,N_19580,N_19450);
nand U19786 (N_19786,N_19515,N_19573);
and U19787 (N_19787,N_19456,N_19430);
and U19788 (N_19788,N_19530,N_19491);
xnor U19789 (N_19789,N_19469,N_19405);
nor U19790 (N_19790,N_19479,N_19520);
xor U19791 (N_19791,N_19447,N_19561);
nor U19792 (N_19792,N_19513,N_19490);
or U19793 (N_19793,N_19527,N_19438);
nand U19794 (N_19794,N_19557,N_19442);
or U19795 (N_19795,N_19540,N_19403);
nor U19796 (N_19796,N_19560,N_19557);
nand U19797 (N_19797,N_19408,N_19536);
or U19798 (N_19798,N_19455,N_19448);
or U19799 (N_19799,N_19519,N_19473);
nand U19800 (N_19800,N_19768,N_19668);
nor U19801 (N_19801,N_19744,N_19633);
nand U19802 (N_19802,N_19740,N_19636);
nor U19803 (N_19803,N_19784,N_19698);
or U19804 (N_19804,N_19734,N_19611);
or U19805 (N_19805,N_19653,N_19649);
and U19806 (N_19806,N_19767,N_19751);
nand U19807 (N_19807,N_19625,N_19618);
nor U19808 (N_19808,N_19728,N_19614);
or U19809 (N_19809,N_19689,N_19745);
nand U19810 (N_19810,N_19790,N_19778);
and U19811 (N_19811,N_19638,N_19796);
nand U19812 (N_19812,N_19712,N_19688);
or U19813 (N_19813,N_19798,N_19774);
and U19814 (N_19814,N_19770,N_19710);
xor U19815 (N_19815,N_19785,N_19732);
nor U19816 (N_19816,N_19755,N_19615);
and U19817 (N_19817,N_19766,N_19604);
nand U19818 (N_19818,N_19640,N_19754);
nand U19819 (N_19819,N_19686,N_19637);
and U19820 (N_19820,N_19717,N_19797);
nand U19821 (N_19821,N_19782,N_19634);
xnor U19822 (N_19822,N_19704,N_19619);
nand U19823 (N_19823,N_19721,N_19746);
nand U19824 (N_19824,N_19616,N_19613);
or U19825 (N_19825,N_19713,N_19656);
nor U19826 (N_19826,N_19666,N_19697);
nor U19827 (N_19827,N_19764,N_19641);
or U19828 (N_19828,N_19632,N_19772);
or U19829 (N_19829,N_19758,N_19642);
xnor U19830 (N_19830,N_19635,N_19724);
or U19831 (N_19831,N_19644,N_19693);
and U19832 (N_19832,N_19628,N_19718);
nand U19833 (N_19833,N_19765,N_19729);
xnor U19834 (N_19834,N_19756,N_19776);
nor U19835 (N_19835,N_19741,N_19675);
or U19836 (N_19836,N_19783,N_19752);
and U19837 (N_19837,N_19645,N_19696);
nor U19838 (N_19838,N_19786,N_19699);
and U19839 (N_19839,N_19791,N_19739);
or U19840 (N_19840,N_19660,N_19648);
nor U19841 (N_19841,N_19714,N_19690);
nor U19842 (N_19842,N_19674,N_19763);
xnor U19843 (N_19843,N_19682,N_19733);
or U19844 (N_19844,N_19759,N_19665);
xnor U19845 (N_19845,N_19792,N_19610);
nand U19846 (N_19846,N_19775,N_19622);
and U19847 (N_19847,N_19657,N_19671);
xnor U19848 (N_19848,N_19787,N_19694);
xnor U19849 (N_19849,N_19612,N_19700);
nor U19850 (N_19850,N_19701,N_19715);
nand U19851 (N_19851,N_19702,N_19651);
or U19852 (N_19852,N_19606,N_19670);
xor U19853 (N_19853,N_19624,N_19769);
nor U19854 (N_19854,N_19779,N_19788);
nor U19855 (N_19855,N_19655,N_19737);
nor U19856 (N_19856,N_19748,N_19692);
xnor U19857 (N_19857,N_19646,N_19603);
nor U19858 (N_19858,N_19771,N_19654);
nand U19859 (N_19859,N_19679,N_19757);
xor U19860 (N_19860,N_19673,N_19722);
and U19861 (N_19861,N_19685,N_19600);
and U19862 (N_19862,N_19680,N_19664);
nor U19863 (N_19863,N_19667,N_19760);
and U19864 (N_19864,N_19607,N_19709);
and U19865 (N_19865,N_19736,N_19761);
or U19866 (N_19866,N_19799,N_19683);
xor U19867 (N_19867,N_19726,N_19631);
nor U19868 (N_19868,N_19773,N_19708);
and U19869 (N_19869,N_19711,N_19602);
nand U19870 (N_19870,N_19691,N_19723);
nor U19871 (N_19871,N_19780,N_19695);
xnor U19872 (N_19872,N_19703,N_19630);
nand U19873 (N_19873,N_19661,N_19738);
xnor U19874 (N_19874,N_19753,N_19781);
and U19875 (N_19875,N_19663,N_19720);
and U19876 (N_19876,N_19747,N_19705);
xnor U19877 (N_19877,N_19681,N_19706);
or U19878 (N_19878,N_19731,N_19730);
xnor U19879 (N_19879,N_19662,N_19735);
nor U19880 (N_19880,N_19727,N_19777);
or U19881 (N_19881,N_19743,N_19750);
nor U19882 (N_19882,N_19620,N_19676);
or U19883 (N_19883,N_19601,N_19659);
and U19884 (N_19884,N_19742,N_19794);
nand U19885 (N_19885,N_19623,N_19789);
and U19886 (N_19886,N_19672,N_19678);
and U19887 (N_19887,N_19650,N_19647);
xor U19888 (N_19888,N_19687,N_19684);
or U19889 (N_19889,N_19793,N_19749);
or U19890 (N_19890,N_19719,N_19639);
nor U19891 (N_19891,N_19669,N_19627);
nand U19892 (N_19892,N_19652,N_19658);
xnor U19893 (N_19893,N_19629,N_19617);
nor U19894 (N_19894,N_19605,N_19725);
xor U19895 (N_19895,N_19626,N_19608);
nor U19896 (N_19896,N_19707,N_19621);
and U19897 (N_19897,N_19677,N_19609);
xor U19898 (N_19898,N_19762,N_19716);
or U19899 (N_19899,N_19643,N_19795);
xor U19900 (N_19900,N_19770,N_19607);
xnor U19901 (N_19901,N_19764,N_19686);
or U19902 (N_19902,N_19658,N_19671);
xor U19903 (N_19903,N_19737,N_19786);
or U19904 (N_19904,N_19790,N_19794);
nor U19905 (N_19905,N_19695,N_19616);
nor U19906 (N_19906,N_19779,N_19671);
nor U19907 (N_19907,N_19654,N_19660);
xor U19908 (N_19908,N_19774,N_19702);
or U19909 (N_19909,N_19668,N_19604);
nand U19910 (N_19910,N_19688,N_19663);
xor U19911 (N_19911,N_19677,N_19603);
xor U19912 (N_19912,N_19702,N_19659);
nor U19913 (N_19913,N_19692,N_19705);
nor U19914 (N_19914,N_19655,N_19635);
nand U19915 (N_19915,N_19617,N_19688);
nor U19916 (N_19916,N_19628,N_19779);
and U19917 (N_19917,N_19636,N_19625);
or U19918 (N_19918,N_19745,N_19799);
nor U19919 (N_19919,N_19663,N_19668);
xnor U19920 (N_19920,N_19627,N_19764);
xnor U19921 (N_19921,N_19745,N_19680);
or U19922 (N_19922,N_19638,N_19746);
xnor U19923 (N_19923,N_19729,N_19664);
or U19924 (N_19924,N_19761,N_19664);
and U19925 (N_19925,N_19651,N_19730);
and U19926 (N_19926,N_19739,N_19744);
xnor U19927 (N_19927,N_19684,N_19621);
and U19928 (N_19928,N_19653,N_19745);
nor U19929 (N_19929,N_19788,N_19607);
or U19930 (N_19930,N_19669,N_19696);
and U19931 (N_19931,N_19602,N_19613);
nand U19932 (N_19932,N_19603,N_19662);
nor U19933 (N_19933,N_19728,N_19764);
or U19934 (N_19934,N_19785,N_19751);
xor U19935 (N_19935,N_19733,N_19619);
nand U19936 (N_19936,N_19780,N_19659);
nand U19937 (N_19937,N_19600,N_19619);
nand U19938 (N_19938,N_19737,N_19612);
nor U19939 (N_19939,N_19701,N_19694);
and U19940 (N_19940,N_19732,N_19778);
xnor U19941 (N_19941,N_19760,N_19797);
nor U19942 (N_19942,N_19778,N_19667);
nand U19943 (N_19943,N_19625,N_19619);
nand U19944 (N_19944,N_19614,N_19696);
and U19945 (N_19945,N_19663,N_19687);
xor U19946 (N_19946,N_19630,N_19794);
or U19947 (N_19947,N_19752,N_19700);
or U19948 (N_19948,N_19750,N_19637);
and U19949 (N_19949,N_19781,N_19608);
or U19950 (N_19950,N_19726,N_19673);
or U19951 (N_19951,N_19607,N_19773);
nand U19952 (N_19952,N_19691,N_19693);
and U19953 (N_19953,N_19740,N_19601);
and U19954 (N_19954,N_19683,N_19723);
nor U19955 (N_19955,N_19741,N_19623);
xor U19956 (N_19956,N_19725,N_19637);
and U19957 (N_19957,N_19627,N_19656);
or U19958 (N_19958,N_19777,N_19607);
or U19959 (N_19959,N_19715,N_19748);
nand U19960 (N_19960,N_19618,N_19620);
nor U19961 (N_19961,N_19641,N_19607);
xor U19962 (N_19962,N_19701,N_19743);
or U19963 (N_19963,N_19674,N_19739);
or U19964 (N_19964,N_19684,N_19637);
xnor U19965 (N_19965,N_19657,N_19745);
nand U19966 (N_19966,N_19773,N_19711);
and U19967 (N_19967,N_19790,N_19672);
and U19968 (N_19968,N_19730,N_19718);
nor U19969 (N_19969,N_19723,N_19782);
nor U19970 (N_19970,N_19683,N_19769);
or U19971 (N_19971,N_19611,N_19633);
xor U19972 (N_19972,N_19665,N_19736);
or U19973 (N_19973,N_19658,N_19741);
nand U19974 (N_19974,N_19699,N_19650);
nand U19975 (N_19975,N_19622,N_19647);
and U19976 (N_19976,N_19672,N_19737);
nor U19977 (N_19977,N_19722,N_19769);
nor U19978 (N_19978,N_19749,N_19652);
xor U19979 (N_19979,N_19714,N_19795);
nand U19980 (N_19980,N_19777,N_19614);
nor U19981 (N_19981,N_19759,N_19604);
nor U19982 (N_19982,N_19783,N_19661);
nand U19983 (N_19983,N_19675,N_19605);
nand U19984 (N_19984,N_19676,N_19688);
nor U19985 (N_19985,N_19628,N_19661);
xor U19986 (N_19986,N_19632,N_19657);
xor U19987 (N_19987,N_19688,N_19742);
xor U19988 (N_19988,N_19784,N_19609);
nand U19989 (N_19989,N_19603,N_19609);
nand U19990 (N_19990,N_19618,N_19601);
xor U19991 (N_19991,N_19709,N_19698);
and U19992 (N_19992,N_19687,N_19675);
or U19993 (N_19993,N_19792,N_19611);
or U19994 (N_19994,N_19683,N_19636);
nand U19995 (N_19995,N_19743,N_19659);
and U19996 (N_19996,N_19693,N_19648);
nand U19997 (N_19997,N_19747,N_19713);
nor U19998 (N_19998,N_19602,N_19658);
nor U19999 (N_19999,N_19679,N_19657);
nand U20000 (N_20000,N_19967,N_19970);
nor U20001 (N_20001,N_19874,N_19871);
or U20002 (N_20002,N_19986,N_19857);
and U20003 (N_20003,N_19889,N_19906);
or U20004 (N_20004,N_19885,N_19966);
nor U20005 (N_20005,N_19983,N_19928);
nor U20006 (N_20006,N_19990,N_19861);
and U20007 (N_20007,N_19802,N_19817);
xnor U20008 (N_20008,N_19933,N_19914);
xnor U20009 (N_20009,N_19979,N_19932);
or U20010 (N_20010,N_19823,N_19921);
nor U20011 (N_20011,N_19930,N_19881);
or U20012 (N_20012,N_19877,N_19996);
nand U20013 (N_20013,N_19995,N_19856);
xor U20014 (N_20014,N_19926,N_19803);
or U20015 (N_20015,N_19903,N_19860);
nor U20016 (N_20016,N_19916,N_19841);
and U20017 (N_20017,N_19893,N_19950);
and U20018 (N_20018,N_19884,N_19956);
xor U20019 (N_20019,N_19837,N_19868);
nor U20020 (N_20020,N_19829,N_19890);
nor U20021 (N_20021,N_19887,N_19876);
nand U20022 (N_20022,N_19820,N_19867);
nor U20023 (N_20023,N_19934,N_19973);
and U20024 (N_20024,N_19961,N_19835);
and U20025 (N_20025,N_19862,N_19911);
and U20026 (N_20026,N_19988,N_19941);
xor U20027 (N_20027,N_19927,N_19946);
or U20028 (N_20028,N_19909,N_19818);
and U20029 (N_20029,N_19839,N_19917);
nor U20030 (N_20030,N_19883,N_19897);
nand U20031 (N_20031,N_19937,N_19858);
nor U20032 (N_20032,N_19985,N_19804);
xor U20033 (N_20033,N_19822,N_19910);
nand U20034 (N_20034,N_19845,N_19880);
and U20035 (N_20035,N_19851,N_19908);
or U20036 (N_20036,N_19975,N_19923);
and U20037 (N_20037,N_19824,N_19844);
or U20038 (N_20038,N_19846,N_19905);
nand U20039 (N_20039,N_19827,N_19832);
and U20040 (N_20040,N_19976,N_19936);
xor U20041 (N_20041,N_19865,N_19968);
nor U20042 (N_20042,N_19918,N_19848);
nand U20043 (N_20043,N_19819,N_19982);
xnor U20044 (N_20044,N_19952,N_19993);
xor U20045 (N_20045,N_19900,N_19863);
and U20046 (N_20046,N_19816,N_19987);
nand U20047 (N_20047,N_19869,N_19974);
nor U20048 (N_20048,N_19977,N_19945);
xor U20049 (N_20049,N_19999,N_19984);
or U20050 (N_20050,N_19944,N_19969);
and U20051 (N_20051,N_19895,N_19929);
xnor U20052 (N_20052,N_19931,N_19808);
xor U20053 (N_20053,N_19864,N_19899);
or U20054 (N_20054,N_19831,N_19947);
nand U20055 (N_20055,N_19898,N_19811);
and U20056 (N_20056,N_19812,N_19913);
xnor U20057 (N_20057,N_19994,N_19922);
or U20058 (N_20058,N_19924,N_19901);
or U20059 (N_20059,N_19888,N_19957);
nand U20060 (N_20060,N_19960,N_19904);
xor U20061 (N_20061,N_19830,N_19886);
and U20062 (N_20062,N_19849,N_19907);
xnor U20063 (N_20063,N_19853,N_19955);
and U20064 (N_20064,N_19843,N_19809);
and U20065 (N_20065,N_19891,N_19838);
and U20066 (N_20066,N_19954,N_19940);
or U20067 (N_20067,N_19821,N_19873);
or U20068 (N_20068,N_19972,N_19981);
and U20069 (N_20069,N_19892,N_19958);
nor U20070 (N_20070,N_19992,N_19836);
or U20071 (N_20071,N_19965,N_19855);
and U20072 (N_20072,N_19872,N_19813);
and U20073 (N_20073,N_19935,N_19964);
nand U20074 (N_20074,N_19805,N_19980);
nand U20075 (N_20075,N_19942,N_19879);
nand U20076 (N_20076,N_19943,N_19870);
nor U20077 (N_20077,N_19847,N_19854);
nor U20078 (N_20078,N_19810,N_19896);
nor U20079 (N_20079,N_19815,N_19806);
xor U20080 (N_20080,N_19894,N_19875);
nand U20081 (N_20081,N_19852,N_19801);
or U20082 (N_20082,N_19866,N_19962);
or U20083 (N_20083,N_19939,N_19807);
nor U20084 (N_20084,N_19951,N_19859);
nand U20085 (N_20085,N_19948,N_19991);
nand U20086 (N_20086,N_19919,N_19971);
xnor U20087 (N_20087,N_19938,N_19826);
nand U20088 (N_20088,N_19878,N_19800);
or U20089 (N_20089,N_19920,N_19997);
nand U20090 (N_20090,N_19912,N_19825);
nor U20091 (N_20091,N_19989,N_19953);
or U20092 (N_20092,N_19842,N_19850);
nand U20093 (N_20093,N_19834,N_19828);
or U20094 (N_20094,N_19814,N_19949);
nand U20095 (N_20095,N_19998,N_19840);
or U20096 (N_20096,N_19978,N_19925);
or U20097 (N_20097,N_19833,N_19959);
or U20098 (N_20098,N_19882,N_19902);
xnor U20099 (N_20099,N_19963,N_19915);
nor U20100 (N_20100,N_19935,N_19829);
nor U20101 (N_20101,N_19865,N_19814);
xnor U20102 (N_20102,N_19935,N_19996);
nor U20103 (N_20103,N_19938,N_19892);
xnor U20104 (N_20104,N_19944,N_19910);
xor U20105 (N_20105,N_19994,N_19921);
or U20106 (N_20106,N_19905,N_19918);
and U20107 (N_20107,N_19827,N_19966);
nand U20108 (N_20108,N_19984,N_19892);
or U20109 (N_20109,N_19915,N_19831);
xnor U20110 (N_20110,N_19858,N_19807);
nand U20111 (N_20111,N_19988,N_19882);
and U20112 (N_20112,N_19938,N_19970);
or U20113 (N_20113,N_19970,N_19820);
nor U20114 (N_20114,N_19973,N_19837);
nor U20115 (N_20115,N_19951,N_19984);
nor U20116 (N_20116,N_19842,N_19906);
and U20117 (N_20117,N_19857,N_19820);
or U20118 (N_20118,N_19800,N_19944);
xnor U20119 (N_20119,N_19862,N_19982);
nand U20120 (N_20120,N_19943,N_19937);
or U20121 (N_20121,N_19974,N_19841);
xor U20122 (N_20122,N_19951,N_19981);
or U20123 (N_20123,N_19936,N_19986);
xor U20124 (N_20124,N_19904,N_19881);
or U20125 (N_20125,N_19987,N_19989);
xor U20126 (N_20126,N_19949,N_19887);
xor U20127 (N_20127,N_19900,N_19857);
nor U20128 (N_20128,N_19927,N_19846);
or U20129 (N_20129,N_19980,N_19885);
xnor U20130 (N_20130,N_19838,N_19816);
or U20131 (N_20131,N_19881,N_19897);
nand U20132 (N_20132,N_19982,N_19826);
nor U20133 (N_20133,N_19800,N_19902);
nand U20134 (N_20134,N_19934,N_19930);
and U20135 (N_20135,N_19837,N_19967);
xnor U20136 (N_20136,N_19993,N_19942);
nor U20137 (N_20137,N_19867,N_19992);
nand U20138 (N_20138,N_19904,N_19914);
and U20139 (N_20139,N_19956,N_19833);
nor U20140 (N_20140,N_19903,N_19978);
nor U20141 (N_20141,N_19866,N_19935);
xor U20142 (N_20142,N_19854,N_19810);
or U20143 (N_20143,N_19845,N_19962);
xnor U20144 (N_20144,N_19978,N_19908);
and U20145 (N_20145,N_19845,N_19852);
xnor U20146 (N_20146,N_19980,N_19996);
and U20147 (N_20147,N_19988,N_19804);
or U20148 (N_20148,N_19958,N_19809);
and U20149 (N_20149,N_19910,N_19805);
nand U20150 (N_20150,N_19966,N_19854);
xnor U20151 (N_20151,N_19857,N_19800);
xor U20152 (N_20152,N_19953,N_19889);
nand U20153 (N_20153,N_19962,N_19814);
xnor U20154 (N_20154,N_19972,N_19893);
or U20155 (N_20155,N_19993,N_19978);
xnor U20156 (N_20156,N_19890,N_19911);
xnor U20157 (N_20157,N_19979,N_19824);
xnor U20158 (N_20158,N_19820,N_19841);
and U20159 (N_20159,N_19834,N_19872);
nor U20160 (N_20160,N_19923,N_19900);
nor U20161 (N_20161,N_19842,N_19836);
and U20162 (N_20162,N_19845,N_19803);
nand U20163 (N_20163,N_19904,N_19810);
nand U20164 (N_20164,N_19856,N_19879);
or U20165 (N_20165,N_19862,N_19904);
xor U20166 (N_20166,N_19951,N_19999);
nor U20167 (N_20167,N_19830,N_19834);
xnor U20168 (N_20168,N_19923,N_19862);
nor U20169 (N_20169,N_19815,N_19859);
nand U20170 (N_20170,N_19936,N_19863);
or U20171 (N_20171,N_19911,N_19934);
nor U20172 (N_20172,N_19883,N_19979);
and U20173 (N_20173,N_19887,N_19850);
nand U20174 (N_20174,N_19923,N_19818);
and U20175 (N_20175,N_19951,N_19901);
nand U20176 (N_20176,N_19942,N_19846);
and U20177 (N_20177,N_19962,N_19957);
and U20178 (N_20178,N_19820,N_19885);
and U20179 (N_20179,N_19966,N_19866);
xor U20180 (N_20180,N_19871,N_19830);
nand U20181 (N_20181,N_19969,N_19977);
and U20182 (N_20182,N_19996,N_19817);
and U20183 (N_20183,N_19993,N_19909);
nand U20184 (N_20184,N_19892,N_19821);
or U20185 (N_20185,N_19867,N_19819);
and U20186 (N_20186,N_19931,N_19800);
nand U20187 (N_20187,N_19932,N_19988);
and U20188 (N_20188,N_19890,N_19852);
xnor U20189 (N_20189,N_19804,N_19877);
and U20190 (N_20190,N_19939,N_19805);
or U20191 (N_20191,N_19961,N_19971);
or U20192 (N_20192,N_19831,N_19941);
xnor U20193 (N_20193,N_19981,N_19853);
nand U20194 (N_20194,N_19940,N_19822);
and U20195 (N_20195,N_19918,N_19887);
or U20196 (N_20196,N_19947,N_19811);
and U20197 (N_20197,N_19947,N_19866);
nand U20198 (N_20198,N_19819,N_19876);
xor U20199 (N_20199,N_19936,N_19922);
nand U20200 (N_20200,N_20117,N_20033);
nor U20201 (N_20201,N_20078,N_20017);
nor U20202 (N_20202,N_20138,N_20190);
and U20203 (N_20203,N_20199,N_20052);
xor U20204 (N_20204,N_20110,N_20161);
xnor U20205 (N_20205,N_20085,N_20049);
nand U20206 (N_20206,N_20015,N_20066);
nor U20207 (N_20207,N_20145,N_20135);
nand U20208 (N_20208,N_20077,N_20067);
xnor U20209 (N_20209,N_20086,N_20063);
nand U20210 (N_20210,N_20149,N_20099);
and U20211 (N_20211,N_20012,N_20150);
and U20212 (N_20212,N_20102,N_20089);
nand U20213 (N_20213,N_20171,N_20043);
or U20214 (N_20214,N_20178,N_20119);
xor U20215 (N_20215,N_20132,N_20127);
or U20216 (N_20216,N_20107,N_20108);
or U20217 (N_20217,N_20064,N_20196);
and U20218 (N_20218,N_20002,N_20047);
or U20219 (N_20219,N_20170,N_20098);
xor U20220 (N_20220,N_20073,N_20131);
xnor U20221 (N_20221,N_20082,N_20023);
nor U20222 (N_20222,N_20160,N_20187);
nand U20223 (N_20223,N_20021,N_20075);
or U20224 (N_20224,N_20134,N_20092);
or U20225 (N_20225,N_20139,N_20068);
nand U20226 (N_20226,N_20151,N_20143);
and U20227 (N_20227,N_20106,N_20120);
or U20228 (N_20228,N_20095,N_20070);
or U20229 (N_20229,N_20115,N_20079);
or U20230 (N_20230,N_20008,N_20177);
nand U20231 (N_20231,N_20100,N_20022);
xor U20232 (N_20232,N_20088,N_20137);
xor U20233 (N_20233,N_20175,N_20061);
and U20234 (N_20234,N_20028,N_20133);
and U20235 (N_20235,N_20162,N_20152);
nand U20236 (N_20236,N_20056,N_20093);
or U20237 (N_20237,N_20153,N_20129);
nor U20238 (N_20238,N_20105,N_20128);
or U20239 (N_20239,N_20164,N_20126);
nand U20240 (N_20240,N_20025,N_20122);
or U20241 (N_20241,N_20193,N_20116);
or U20242 (N_20242,N_20188,N_20158);
xor U20243 (N_20243,N_20024,N_20121);
nor U20244 (N_20244,N_20154,N_20059);
xnor U20245 (N_20245,N_20146,N_20189);
or U20246 (N_20246,N_20007,N_20032);
or U20247 (N_20247,N_20176,N_20148);
nand U20248 (N_20248,N_20060,N_20080);
or U20249 (N_20249,N_20091,N_20103);
and U20250 (N_20250,N_20186,N_20042);
nand U20251 (N_20251,N_20136,N_20019);
or U20252 (N_20252,N_20005,N_20010);
nor U20253 (N_20253,N_20183,N_20179);
and U20254 (N_20254,N_20046,N_20053);
xor U20255 (N_20255,N_20048,N_20014);
and U20256 (N_20256,N_20030,N_20011);
xor U20257 (N_20257,N_20191,N_20113);
nand U20258 (N_20258,N_20156,N_20141);
and U20259 (N_20259,N_20087,N_20071);
or U20260 (N_20260,N_20006,N_20026);
nor U20261 (N_20261,N_20197,N_20094);
xor U20262 (N_20262,N_20034,N_20055);
or U20263 (N_20263,N_20027,N_20018);
xnor U20264 (N_20264,N_20009,N_20147);
and U20265 (N_20265,N_20038,N_20084);
nor U20266 (N_20266,N_20112,N_20192);
xor U20267 (N_20267,N_20083,N_20004);
and U20268 (N_20268,N_20054,N_20173);
nor U20269 (N_20269,N_20044,N_20029);
and U20270 (N_20270,N_20140,N_20051);
and U20271 (N_20271,N_20035,N_20090);
nand U20272 (N_20272,N_20142,N_20155);
and U20273 (N_20273,N_20058,N_20167);
xnor U20274 (N_20274,N_20166,N_20076);
and U20275 (N_20275,N_20036,N_20081);
xnor U20276 (N_20276,N_20045,N_20037);
xor U20277 (N_20277,N_20169,N_20096);
xor U20278 (N_20278,N_20101,N_20041);
xor U20279 (N_20279,N_20111,N_20198);
or U20280 (N_20280,N_20185,N_20118);
nand U20281 (N_20281,N_20001,N_20031);
nor U20282 (N_20282,N_20016,N_20062);
nor U20283 (N_20283,N_20039,N_20065);
and U20284 (N_20284,N_20124,N_20174);
nand U20285 (N_20285,N_20050,N_20163);
nand U20286 (N_20286,N_20109,N_20069);
and U20287 (N_20287,N_20000,N_20165);
nand U20288 (N_20288,N_20040,N_20097);
nand U20289 (N_20289,N_20114,N_20057);
nand U20290 (N_20290,N_20003,N_20104);
nor U20291 (N_20291,N_20123,N_20144);
nor U20292 (N_20292,N_20194,N_20074);
and U20293 (N_20293,N_20180,N_20181);
nand U20294 (N_20294,N_20184,N_20072);
and U20295 (N_20295,N_20157,N_20195);
xor U20296 (N_20296,N_20159,N_20172);
and U20297 (N_20297,N_20130,N_20182);
nor U20298 (N_20298,N_20020,N_20168);
nor U20299 (N_20299,N_20013,N_20125);
or U20300 (N_20300,N_20176,N_20038);
and U20301 (N_20301,N_20118,N_20139);
or U20302 (N_20302,N_20134,N_20124);
nand U20303 (N_20303,N_20169,N_20056);
nor U20304 (N_20304,N_20092,N_20110);
and U20305 (N_20305,N_20046,N_20105);
xnor U20306 (N_20306,N_20093,N_20162);
or U20307 (N_20307,N_20059,N_20088);
and U20308 (N_20308,N_20054,N_20155);
xnor U20309 (N_20309,N_20074,N_20188);
and U20310 (N_20310,N_20115,N_20187);
xnor U20311 (N_20311,N_20029,N_20158);
or U20312 (N_20312,N_20089,N_20087);
nor U20313 (N_20313,N_20103,N_20082);
nand U20314 (N_20314,N_20087,N_20042);
and U20315 (N_20315,N_20160,N_20115);
or U20316 (N_20316,N_20123,N_20080);
or U20317 (N_20317,N_20162,N_20189);
or U20318 (N_20318,N_20046,N_20060);
and U20319 (N_20319,N_20190,N_20088);
nor U20320 (N_20320,N_20155,N_20075);
and U20321 (N_20321,N_20057,N_20005);
and U20322 (N_20322,N_20025,N_20064);
or U20323 (N_20323,N_20072,N_20010);
nor U20324 (N_20324,N_20170,N_20020);
nor U20325 (N_20325,N_20173,N_20021);
xnor U20326 (N_20326,N_20112,N_20070);
nor U20327 (N_20327,N_20077,N_20176);
xnor U20328 (N_20328,N_20050,N_20061);
and U20329 (N_20329,N_20195,N_20081);
or U20330 (N_20330,N_20113,N_20179);
xnor U20331 (N_20331,N_20124,N_20189);
nor U20332 (N_20332,N_20110,N_20033);
nor U20333 (N_20333,N_20064,N_20190);
xor U20334 (N_20334,N_20052,N_20030);
nor U20335 (N_20335,N_20088,N_20018);
xnor U20336 (N_20336,N_20156,N_20090);
nand U20337 (N_20337,N_20184,N_20071);
nand U20338 (N_20338,N_20133,N_20194);
nand U20339 (N_20339,N_20178,N_20125);
xnor U20340 (N_20340,N_20170,N_20147);
and U20341 (N_20341,N_20101,N_20046);
or U20342 (N_20342,N_20147,N_20044);
nor U20343 (N_20343,N_20146,N_20047);
nand U20344 (N_20344,N_20091,N_20014);
xnor U20345 (N_20345,N_20108,N_20192);
xor U20346 (N_20346,N_20124,N_20155);
and U20347 (N_20347,N_20135,N_20041);
or U20348 (N_20348,N_20186,N_20080);
nand U20349 (N_20349,N_20097,N_20195);
nor U20350 (N_20350,N_20076,N_20142);
or U20351 (N_20351,N_20005,N_20088);
or U20352 (N_20352,N_20155,N_20101);
nand U20353 (N_20353,N_20017,N_20034);
and U20354 (N_20354,N_20132,N_20152);
nand U20355 (N_20355,N_20117,N_20061);
or U20356 (N_20356,N_20044,N_20165);
nand U20357 (N_20357,N_20006,N_20065);
nor U20358 (N_20358,N_20191,N_20180);
xor U20359 (N_20359,N_20164,N_20124);
nor U20360 (N_20360,N_20037,N_20069);
nand U20361 (N_20361,N_20124,N_20040);
nor U20362 (N_20362,N_20159,N_20021);
or U20363 (N_20363,N_20149,N_20112);
and U20364 (N_20364,N_20187,N_20128);
nor U20365 (N_20365,N_20166,N_20177);
nor U20366 (N_20366,N_20039,N_20190);
nand U20367 (N_20367,N_20012,N_20162);
nor U20368 (N_20368,N_20078,N_20180);
nor U20369 (N_20369,N_20132,N_20088);
and U20370 (N_20370,N_20100,N_20012);
or U20371 (N_20371,N_20021,N_20041);
or U20372 (N_20372,N_20041,N_20141);
or U20373 (N_20373,N_20043,N_20150);
and U20374 (N_20374,N_20073,N_20194);
or U20375 (N_20375,N_20134,N_20032);
or U20376 (N_20376,N_20062,N_20046);
and U20377 (N_20377,N_20059,N_20052);
and U20378 (N_20378,N_20114,N_20141);
and U20379 (N_20379,N_20161,N_20030);
xnor U20380 (N_20380,N_20072,N_20032);
and U20381 (N_20381,N_20089,N_20145);
nor U20382 (N_20382,N_20058,N_20005);
nand U20383 (N_20383,N_20131,N_20046);
nand U20384 (N_20384,N_20121,N_20035);
and U20385 (N_20385,N_20072,N_20176);
and U20386 (N_20386,N_20017,N_20177);
or U20387 (N_20387,N_20198,N_20178);
xor U20388 (N_20388,N_20079,N_20055);
or U20389 (N_20389,N_20105,N_20194);
nor U20390 (N_20390,N_20095,N_20136);
nor U20391 (N_20391,N_20164,N_20063);
nor U20392 (N_20392,N_20159,N_20057);
nor U20393 (N_20393,N_20031,N_20040);
nor U20394 (N_20394,N_20171,N_20005);
or U20395 (N_20395,N_20148,N_20108);
or U20396 (N_20396,N_20044,N_20166);
nand U20397 (N_20397,N_20149,N_20053);
xor U20398 (N_20398,N_20133,N_20187);
or U20399 (N_20399,N_20001,N_20131);
nand U20400 (N_20400,N_20296,N_20341);
xnor U20401 (N_20401,N_20201,N_20247);
nand U20402 (N_20402,N_20287,N_20305);
or U20403 (N_20403,N_20350,N_20318);
or U20404 (N_20404,N_20313,N_20230);
xnor U20405 (N_20405,N_20309,N_20399);
xor U20406 (N_20406,N_20250,N_20256);
nand U20407 (N_20407,N_20385,N_20277);
or U20408 (N_20408,N_20294,N_20348);
or U20409 (N_20409,N_20332,N_20288);
or U20410 (N_20410,N_20244,N_20359);
nor U20411 (N_20411,N_20370,N_20384);
nand U20412 (N_20412,N_20395,N_20272);
or U20413 (N_20413,N_20209,N_20293);
nand U20414 (N_20414,N_20393,N_20324);
xor U20415 (N_20415,N_20358,N_20369);
nand U20416 (N_20416,N_20265,N_20327);
nand U20417 (N_20417,N_20255,N_20205);
nand U20418 (N_20418,N_20319,N_20392);
nand U20419 (N_20419,N_20295,N_20337);
nor U20420 (N_20420,N_20286,N_20284);
and U20421 (N_20421,N_20223,N_20326);
nor U20422 (N_20422,N_20300,N_20335);
or U20423 (N_20423,N_20377,N_20215);
xnor U20424 (N_20424,N_20371,N_20290);
nor U20425 (N_20425,N_20374,N_20356);
xnor U20426 (N_20426,N_20301,N_20264);
or U20427 (N_20427,N_20308,N_20389);
nor U20428 (N_20428,N_20396,N_20259);
nand U20429 (N_20429,N_20239,N_20345);
nand U20430 (N_20430,N_20200,N_20211);
or U20431 (N_20431,N_20343,N_20273);
or U20432 (N_20432,N_20258,N_20231);
nand U20433 (N_20433,N_20283,N_20360);
or U20434 (N_20434,N_20257,N_20373);
or U20435 (N_20435,N_20372,N_20333);
xnor U20436 (N_20436,N_20316,N_20275);
xor U20437 (N_20437,N_20346,N_20315);
nand U20438 (N_20438,N_20364,N_20251);
or U20439 (N_20439,N_20362,N_20241);
xnor U20440 (N_20440,N_20271,N_20357);
or U20441 (N_20441,N_20376,N_20234);
or U20442 (N_20442,N_20363,N_20276);
nand U20443 (N_20443,N_20367,N_20342);
nor U20444 (N_20444,N_20322,N_20391);
nor U20445 (N_20445,N_20352,N_20302);
nor U20446 (N_20446,N_20260,N_20334);
xor U20447 (N_20447,N_20289,N_20388);
xnor U20448 (N_20448,N_20262,N_20349);
nor U20449 (N_20449,N_20361,N_20387);
or U20450 (N_20450,N_20204,N_20394);
xor U20451 (N_20451,N_20226,N_20390);
and U20452 (N_20452,N_20268,N_20245);
nand U20453 (N_20453,N_20397,N_20236);
and U20454 (N_20454,N_20219,N_20323);
or U20455 (N_20455,N_20375,N_20366);
nor U20456 (N_20456,N_20202,N_20248);
nand U20457 (N_20457,N_20213,N_20380);
nand U20458 (N_20458,N_20218,N_20254);
and U20459 (N_20459,N_20381,N_20382);
or U20460 (N_20460,N_20225,N_20263);
and U20461 (N_20461,N_20207,N_20398);
nor U20462 (N_20462,N_20383,N_20206);
nor U20463 (N_20463,N_20238,N_20270);
xor U20464 (N_20464,N_20320,N_20365);
and U20465 (N_20465,N_20351,N_20214);
and U20466 (N_20466,N_20329,N_20306);
xnor U20467 (N_20467,N_20338,N_20210);
xnor U20468 (N_20468,N_20292,N_20355);
or U20469 (N_20469,N_20267,N_20208);
or U20470 (N_20470,N_20344,N_20321);
xnor U20471 (N_20471,N_20297,N_20330);
xnor U20472 (N_20472,N_20221,N_20378);
nand U20473 (N_20473,N_20229,N_20222);
or U20474 (N_20474,N_20278,N_20242);
and U20475 (N_20475,N_20228,N_20212);
nand U20476 (N_20476,N_20285,N_20331);
or U20477 (N_20477,N_20336,N_20253);
and U20478 (N_20478,N_20261,N_20340);
and U20479 (N_20479,N_20237,N_20291);
or U20480 (N_20480,N_20303,N_20246);
xnor U20481 (N_20481,N_20314,N_20347);
and U20482 (N_20482,N_20282,N_20307);
or U20483 (N_20483,N_20217,N_20353);
nand U20484 (N_20484,N_20224,N_20386);
or U20485 (N_20485,N_20339,N_20216);
or U20486 (N_20486,N_20249,N_20281);
or U20487 (N_20487,N_20227,N_20280);
xnor U20488 (N_20488,N_20240,N_20310);
nand U20489 (N_20489,N_20311,N_20235);
xnor U20490 (N_20490,N_20203,N_20266);
or U20491 (N_20491,N_20379,N_20312);
or U20492 (N_20492,N_20354,N_20298);
nor U20493 (N_20493,N_20274,N_20317);
nor U20494 (N_20494,N_20328,N_20368);
nand U20495 (N_20495,N_20299,N_20252);
or U20496 (N_20496,N_20220,N_20232);
and U20497 (N_20497,N_20243,N_20304);
and U20498 (N_20498,N_20269,N_20325);
or U20499 (N_20499,N_20233,N_20279);
xnor U20500 (N_20500,N_20320,N_20264);
nand U20501 (N_20501,N_20254,N_20223);
xor U20502 (N_20502,N_20342,N_20351);
or U20503 (N_20503,N_20297,N_20302);
xnor U20504 (N_20504,N_20239,N_20217);
nor U20505 (N_20505,N_20311,N_20223);
xor U20506 (N_20506,N_20260,N_20370);
nand U20507 (N_20507,N_20260,N_20235);
nor U20508 (N_20508,N_20376,N_20228);
and U20509 (N_20509,N_20276,N_20307);
and U20510 (N_20510,N_20393,N_20299);
nand U20511 (N_20511,N_20340,N_20370);
nor U20512 (N_20512,N_20359,N_20220);
or U20513 (N_20513,N_20206,N_20366);
or U20514 (N_20514,N_20328,N_20370);
xnor U20515 (N_20515,N_20386,N_20351);
nor U20516 (N_20516,N_20224,N_20332);
nor U20517 (N_20517,N_20356,N_20336);
nand U20518 (N_20518,N_20204,N_20315);
nand U20519 (N_20519,N_20366,N_20255);
nand U20520 (N_20520,N_20368,N_20279);
or U20521 (N_20521,N_20267,N_20379);
and U20522 (N_20522,N_20322,N_20287);
xnor U20523 (N_20523,N_20388,N_20347);
nand U20524 (N_20524,N_20335,N_20209);
or U20525 (N_20525,N_20294,N_20381);
or U20526 (N_20526,N_20249,N_20257);
nand U20527 (N_20527,N_20321,N_20389);
or U20528 (N_20528,N_20249,N_20284);
xor U20529 (N_20529,N_20248,N_20299);
nand U20530 (N_20530,N_20308,N_20276);
or U20531 (N_20531,N_20205,N_20332);
nand U20532 (N_20532,N_20221,N_20203);
or U20533 (N_20533,N_20298,N_20393);
nor U20534 (N_20534,N_20282,N_20398);
xor U20535 (N_20535,N_20201,N_20368);
xor U20536 (N_20536,N_20282,N_20350);
and U20537 (N_20537,N_20309,N_20231);
or U20538 (N_20538,N_20228,N_20324);
nand U20539 (N_20539,N_20284,N_20365);
and U20540 (N_20540,N_20249,N_20218);
nand U20541 (N_20541,N_20202,N_20395);
or U20542 (N_20542,N_20253,N_20370);
nand U20543 (N_20543,N_20253,N_20259);
nand U20544 (N_20544,N_20267,N_20342);
and U20545 (N_20545,N_20374,N_20324);
xnor U20546 (N_20546,N_20230,N_20317);
and U20547 (N_20547,N_20367,N_20394);
or U20548 (N_20548,N_20366,N_20289);
and U20549 (N_20549,N_20338,N_20357);
and U20550 (N_20550,N_20327,N_20378);
or U20551 (N_20551,N_20357,N_20266);
nor U20552 (N_20552,N_20342,N_20253);
nor U20553 (N_20553,N_20229,N_20294);
and U20554 (N_20554,N_20302,N_20306);
and U20555 (N_20555,N_20383,N_20225);
or U20556 (N_20556,N_20324,N_20249);
nor U20557 (N_20557,N_20211,N_20325);
or U20558 (N_20558,N_20291,N_20350);
nor U20559 (N_20559,N_20245,N_20375);
xor U20560 (N_20560,N_20386,N_20348);
nand U20561 (N_20561,N_20247,N_20354);
xnor U20562 (N_20562,N_20331,N_20219);
xnor U20563 (N_20563,N_20220,N_20208);
or U20564 (N_20564,N_20367,N_20387);
and U20565 (N_20565,N_20269,N_20290);
and U20566 (N_20566,N_20278,N_20360);
nor U20567 (N_20567,N_20333,N_20302);
nor U20568 (N_20568,N_20397,N_20297);
or U20569 (N_20569,N_20220,N_20308);
xnor U20570 (N_20570,N_20320,N_20226);
nor U20571 (N_20571,N_20236,N_20386);
xor U20572 (N_20572,N_20205,N_20309);
xnor U20573 (N_20573,N_20281,N_20205);
nand U20574 (N_20574,N_20352,N_20375);
nor U20575 (N_20575,N_20239,N_20245);
and U20576 (N_20576,N_20383,N_20221);
and U20577 (N_20577,N_20365,N_20342);
nor U20578 (N_20578,N_20208,N_20274);
nor U20579 (N_20579,N_20323,N_20230);
or U20580 (N_20580,N_20207,N_20231);
xnor U20581 (N_20581,N_20336,N_20285);
or U20582 (N_20582,N_20256,N_20384);
nor U20583 (N_20583,N_20221,N_20298);
or U20584 (N_20584,N_20318,N_20329);
nor U20585 (N_20585,N_20259,N_20313);
xor U20586 (N_20586,N_20394,N_20322);
or U20587 (N_20587,N_20213,N_20378);
nand U20588 (N_20588,N_20240,N_20320);
and U20589 (N_20589,N_20216,N_20287);
xnor U20590 (N_20590,N_20292,N_20242);
xnor U20591 (N_20591,N_20317,N_20240);
nand U20592 (N_20592,N_20209,N_20230);
xor U20593 (N_20593,N_20380,N_20381);
or U20594 (N_20594,N_20356,N_20217);
nand U20595 (N_20595,N_20307,N_20384);
and U20596 (N_20596,N_20391,N_20337);
nand U20597 (N_20597,N_20208,N_20251);
nor U20598 (N_20598,N_20385,N_20264);
nor U20599 (N_20599,N_20299,N_20267);
nor U20600 (N_20600,N_20453,N_20421);
xnor U20601 (N_20601,N_20450,N_20515);
or U20602 (N_20602,N_20591,N_20442);
nand U20603 (N_20603,N_20571,N_20495);
nand U20604 (N_20604,N_20523,N_20522);
and U20605 (N_20605,N_20463,N_20437);
and U20606 (N_20606,N_20461,N_20483);
xnor U20607 (N_20607,N_20576,N_20468);
and U20608 (N_20608,N_20537,N_20543);
and U20609 (N_20609,N_20562,N_20504);
or U20610 (N_20610,N_20434,N_20592);
nor U20611 (N_20611,N_20449,N_20406);
nand U20612 (N_20612,N_20502,N_20569);
or U20613 (N_20613,N_20503,N_20597);
and U20614 (N_20614,N_20519,N_20563);
nor U20615 (N_20615,N_20587,N_20538);
xor U20616 (N_20616,N_20459,N_20520);
or U20617 (N_20617,N_20521,N_20555);
nand U20618 (N_20618,N_20542,N_20478);
xnor U20619 (N_20619,N_20544,N_20477);
nor U20620 (N_20620,N_20526,N_20558);
and U20621 (N_20621,N_20496,N_20480);
and U20622 (N_20622,N_20428,N_20490);
xnor U20623 (N_20623,N_20551,N_20529);
or U20624 (N_20624,N_20401,N_20443);
or U20625 (N_20625,N_20582,N_20589);
xnor U20626 (N_20626,N_20455,N_20416);
and U20627 (N_20627,N_20420,N_20457);
nand U20628 (N_20628,N_20510,N_20512);
or U20629 (N_20629,N_20426,N_20586);
xor U20630 (N_20630,N_20432,N_20422);
and U20631 (N_20631,N_20511,N_20473);
or U20632 (N_20632,N_20417,N_20583);
nor U20633 (N_20633,N_20580,N_20404);
nand U20634 (N_20634,N_20516,N_20427);
nor U20635 (N_20635,N_20418,N_20472);
and U20636 (N_20636,N_20545,N_20524);
and U20637 (N_20637,N_20488,N_20445);
xnor U20638 (N_20638,N_20527,N_20460);
and U20639 (N_20639,N_20435,N_20448);
nand U20640 (N_20640,N_20541,N_20499);
and U20641 (N_20641,N_20439,N_20409);
and U20642 (N_20642,N_20474,N_20419);
nand U20643 (N_20643,N_20564,N_20424);
or U20644 (N_20644,N_20531,N_20475);
nor U20645 (N_20645,N_20407,N_20585);
and U20646 (N_20646,N_20400,N_20550);
nand U20647 (N_20647,N_20458,N_20476);
nor U20648 (N_20648,N_20412,N_20590);
nand U20649 (N_20649,N_20556,N_20567);
nor U20650 (N_20650,N_20436,N_20492);
xor U20651 (N_20651,N_20561,N_20467);
xor U20652 (N_20652,N_20414,N_20494);
nand U20653 (N_20653,N_20595,N_20506);
or U20654 (N_20654,N_20447,N_20441);
nand U20655 (N_20655,N_20493,N_20593);
nand U20656 (N_20656,N_20501,N_20572);
and U20657 (N_20657,N_20575,N_20464);
or U20658 (N_20658,N_20479,N_20540);
xnor U20659 (N_20659,N_20518,N_20484);
nand U20660 (N_20660,N_20568,N_20402);
xor U20661 (N_20661,N_20588,N_20456);
or U20662 (N_20662,N_20560,N_20599);
xnor U20663 (N_20663,N_20444,N_20451);
or U20664 (N_20664,N_20554,N_20430);
nor U20665 (N_20665,N_20565,N_20546);
xnor U20666 (N_20666,N_20471,N_20552);
or U20667 (N_20667,N_20415,N_20513);
or U20668 (N_20668,N_20462,N_20581);
xnor U20669 (N_20669,N_20548,N_20440);
xor U20670 (N_20670,N_20486,N_20525);
xor U20671 (N_20671,N_20465,N_20577);
nand U20672 (N_20672,N_20491,N_20466);
nor U20673 (N_20673,N_20429,N_20536);
and U20674 (N_20674,N_20509,N_20489);
or U20675 (N_20675,N_20514,N_20425);
xnor U20676 (N_20676,N_20532,N_20570);
xnor U20677 (N_20677,N_20549,N_20487);
or U20678 (N_20678,N_20553,N_20470);
and U20679 (N_20679,N_20584,N_20469);
xnor U20680 (N_20680,N_20578,N_20594);
and U20681 (N_20681,N_20534,N_20559);
or U20682 (N_20682,N_20533,N_20574);
nor U20683 (N_20683,N_20433,N_20598);
nand U20684 (N_20684,N_20517,N_20547);
xnor U20685 (N_20685,N_20403,N_20505);
xnor U20686 (N_20686,N_20454,N_20482);
and U20687 (N_20687,N_20530,N_20423);
nand U20688 (N_20688,N_20452,N_20438);
nor U20689 (N_20689,N_20413,N_20535);
or U20690 (N_20690,N_20596,N_20539);
nor U20691 (N_20691,N_20405,N_20500);
and U20692 (N_20692,N_20528,N_20411);
nand U20693 (N_20693,N_20557,N_20573);
xnor U20694 (N_20694,N_20507,N_20497);
and U20695 (N_20695,N_20579,N_20498);
and U20696 (N_20696,N_20508,N_20431);
xor U20697 (N_20697,N_20410,N_20481);
or U20698 (N_20698,N_20485,N_20446);
or U20699 (N_20699,N_20566,N_20408);
and U20700 (N_20700,N_20463,N_20527);
xnor U20701 (N_20701,N_20552,N_20544);
or U20702 (N_20702,N_20503,N_20469);
or U20703 (N_20703,N_20486,N_20497);
and U20704 (N_20704,N_20533,N_20514);
xnor U20705 (N_20705,N_20495,N_20507);
nand U20706 (N_20706,N_20437,N_20428);
or U20707 (N_20707,N_20551,N_20591);
or U20708 (N_20708,N_20486,N_20482);
nand U20709 (N_20709,N_20495,N_20425);
nor U20710 (N_20710,N_20486,N_20566);
nand U20711 (N_20711,N_20459,N_20563);
and U20712 (N_20712,N_20548,N_20473);
nand U20713 (N_20713,N_20403,N_20485);
or U20714 (N_20714,N_20494,N_20546);
xor U20715 (N_20715,N_20596,N_20433);
xnor U20716 (N_20716,N_20517,N_20476);
and U20717 (N_20717,N_20412,N_20494);
nor U20718 (N_20718,N_20435,N_20486);
or U20719 (N_20719,N_20498,N_20595);
xnor U20720 (N_20720,N_20579,N_20481);
xnor U20721 (N_20721,N_20523,N_20423);
nand U20722 (N_20722,N_20444,N_20593);
and U20723 (N_20723,N_20416,N_20427);
nand U20724 (N_20724,N_20581,N_20420);
nand U20725 (N_20725,N_20473,N_20515);
nor U20726 (N_20726,N_20522,N_20506);
nand U20727 (N_20727,N_20470,N_20442);
xnor U20728 (N_20728,N_20405,N_20404);
nand U20729 (N_20729,N_20484,N_20566);
nor U20730 (N_20730,N_20456,N_20586);
xor U20731 (N_20731,N_20515,N_20469);
or U20732 (N_20732,N_20443,N_20555);
nand U20733 (N_20733,N_20533,N_20543);
and U20734 (N_20734,N_20480,N_20483);
or U20735 (N_20735,N_20458,N_20452);
nor U20736 (N_20736,N_20400,N_20469);
and U20737 (N_20737,N_20479,N_20454);
or U20738 (N_20738,N_20419,N_20567);
xnor U20739 (N_20739,N_20569,N_20472);
nor U20740 (N_20740,N_20573,N_20536);
or U20741 (N_20741,N_20450,N_20475);
nor U20742 (N_20742,N_20451,N_20481);
nand U20743 (N_20743,N_20527,N_20474);
nor U20744 (N_20744,N_20434,N_20538);
and U20745 (N_20745,N_20513,N_20582);
and U20746 (N_20746,N_20466,N_20485);
nand U20747 (N_20747,N_20537,N_20554);
nand U20748 (N_20748,N_20500,N_20445);
and U20749 (N_20749,N_20456,N_20439);
nand U20750 (N_20750,N_20445,N_20438);
nor U20751 (N_20751,N_20528,N_20406);
xnor U20752 (N_20752,N_20498,N_20497);
nand U20753 (N_20753,N_20492,N_20475);
nor U20754 (N_20754,N_20580,N_20501);
xor U20755 (N_20755,N_20446,N_20555);
xor U20756 (N_20756,N_20589,N_20456);
and U20757 (N_20757,N_20502,N_20468);
nand U20758 (N_20758,N_20572,N_20549);
and U20759 (N_20759,N_20480,N_20577);
nor U20760 (N_20760,N_20556,N_20505);
nand U20761 (N_20761,N_20402,N_20459);
nand U20762 (N_20762,N_20400,N_20556);
nand U20763 (N_20763,N_20441,N_20513);
xor U20764 (N_20764,N_20453,N_20588);
nor U20765 (N_20765,N_20499,N_20468);
and U20766 (N_20766,N_20527,N_20472);
xor U20767 (N_20767,N_20468,N_20439);
xnor U20768 (N_20768,N_20456,N_20551);
and U20769 (N_20769,N_20493,N_20573);
xnor U20770 (N_20770,N_20563,N_20410);
xor U20771 (N_20771,N_20536,N_20587);
and U20772 (N_20772,N_20529,N_20530);
nand U20773 (N_20773,N_20507,N_20427);
nor U20774 (N_20774,N_20569,N_20411);
nor U20775 (N_20775,N_20516,N_20539);
or U20776 (N_20776,N_20450,N_20442);
and U20777 (N_20777,N_20502,N_20466);
nor U20778 (N_20778,N_20504,N_20599);
xor U20779 (N_20779,N_20571,N_20426);
nor U20780 (N_20780,N_20543,N_20498);
nand U20781 (N_20781,N_20463,N_20596);
nand U20782 (N_20782,N_20507,N_20540);
or U20783 (N_20783,N_20521,N_20441);
nor U20784 (N_20784,N_20500,N_20568);
nor U20785 (N_20785,N_20515,N_20488);
xor U20786 (N_20786,N_20509,N_20504);
and U20787 (N_20787,N_20455,N_20476);
nor U20788 (N_20788,N_20493,N_20539);
xnor U20789 (N_20789,N_20481,N_20510);
nor U20790 (N_20790,N_20465,N_20544);
and U20791 (N_20791,N_20571,N_20550);
nor U20792 (N_20792,N_20412,N_20520);
nand U20793 (N_20793,N_20506,N_20513);
and U20794 (N_20794,N_20430,N_20461);
nor U20795 (N_20795,N_20497,N_20463);
nand U20796 (N_20796,N_20529,N_20479);
or U20797 (N_20797,N_20419,N_20431);
nor U20798 (N_20798,N_20549,N_20428);
nand U20799 (N_20799,N_20486,N_20471);
xnor U20800 (N_20800,N_20737,N_20746);
xor U20801 (N_20801,N_20745,N_20715);
xnor U20802 (N_20802,N_20735,N_20644);
nor U20803 (N_20803,N_20654,N_20690);
xor U20804 (N_20804,N_20607,N_20664);
nand U20805 (N_20805,N_20641,N_20759);
nand U20806 (N_20806,N_20619,N_20733);
nand U20807 (N_20807,N_20718,N_20787);
and U20808 (N_20808,N_20772,N_20628);
xor U20809 (N_20809,N_20739,N_20642);
xor U20810 (N_20810,N_20716,N_20754);
xor U20811 (N_20811,N_20790,N_20647);
nor U20812 (N_20812,N_20680,N_20768);
nor U20813 (N_20813,N_20695,N_20722);
nor U20814 (N_20814,N_20663,N_20609);
nand U20815 (N_20815,N_20719,N_20688);
and U20816 (N_20816,N_20764,N_20639);
or U20817 (N_20817,N_20651,N_20789);
or U20818 (N_20818,N_20659,N_20625);
xnor U20819 (N_20819,N_20756,N_20649);
xor U20820 (N_20820,N_20721,N_20788);
nor U20821 (N_20821,N_20684,N_20742);
and U20822 (N_20822,N_20708,N_20705);
nor U20823 (N_20823,N_20623,N_20776);
or U20824 (N_20824,N_20694,N_20782);
nor U20825 (N_20825,N_20757,N_20668);
nor U20826 (N_20826,N_20773,N_20653);
nor U20827 (N_20827,N_20677,N_20687);
nor U20828 (N_20828,N_20741,N_20794);
nand U20829 (N_20829,N_20662,N_20701);
xor U20830 (N_20830,N_20646,N_20755);
xnor U20831 (N_20831,N_20784,N_20686);
xnor U20832 (N_20832,N_20732,N_20611);
nand U20833 (N_20833,N_20792,N_20614);
and U20834 (N_20834,N_20671,N_20748);
or U20835 (N_20835,N_20779,N_20658);
nand U20836 (N_20836,N_20743,N_20632);
nand U20837 (N_20837,N_20786,N_20697);
xnor U20838 (N_20838,N_20640,N_20744);
and U20839 (N_20839,N_20793,N_20622);
nand U20840 (N_20840,N_20774,N_20672);
nand U20841 (N_20841,N_20652,N_20669);
nand U20842 (N_20842,N_20600,N_20621);
xnor U20843 (N_20843,N_20712,N_20692);
xor U20844 (N_20844,N_20781,N_20747);
or U20845 (N_20845,N_20750,N_20796);
and U20846 (N_20846,N_20717,N_20758);
and U20847 (N_20847,N_20727,N_20630);
or U20848 (N_20848,N_20603,N_20724);
xnor U20849 (N_20849,N_20730,N_20615);
xnor U20850 (N_20850,N_20638,N_20656);
nor U20851 (N_20851,N_20637,N_20602);
xnor U20852 (N_20852,N_20673,N_20799);
or U20853 (N_20853,N_20728,N_20725);
xnor U20854 (N_20854,N_20685,N_20783);
and U20855 (N_20855,N_20766,N_20631);
xor U20856 (N_20856,N_20626,N_20665);
xor U20857 (N_20857,N_20765,N_20752);
xor U20858 (N_20858,N_20601,N_20740);
or U20859 (N_20859,N_20711,N_20679);
xnor U20860 (N_20860,N_20785,N_20612);
and U20861 (N_20861,N_20618,N_20797);
nor U20862 (N_20862,N_20780,N_20606);
or U20863 (N_20863,N_20667,N_20762);
and U20864 (N_20864,N_20770,N_20771);
nand U20865 (N_20865,N_20761,N_20749);
nand U20866 (N_20866,N_20734,N_20635);
xor U20867 (N_20867,N_20650,N_20643);
nor U20868 (N_20868,N_20702,N_20703);
nand U20869 (N_20869,N_20723,N_20699);
or U20870 (N_20870,N_20657,N_20798);
and U20871 (N_20871,N_20753,N_20666);
xnor U20872 (N_20872,N_20660,N_20674);
xnor U20873 (N_20873,N_20624,N_20605);
xnor U20874 (N_20874,N_20636,N_20736);
nand U20875 (N_20875,N_20707,N_20655);
or U20876 (N_20876,N_20729,N_20709);
or U20877 (N_20877,N_20629,N_20675);
or U20878 (N_20878,N_20769,N_20633);
xor U20879 (N_20879,N_20731,N_20610);
nor U20880 (N_20880,N_20682,N_20751);
xnor U20881 (N_20881,N_20700,N_20720);
xor U20882 (N_20882,N_20704,N_20706);
nor U20883 (N_20883,N_20613,N_20713);
or U20884 (N_20884,N_20645,N_20616);
nand U20885 (N_20885,N_20763,N_20693);
xor U20886 (N_20886,N_20777,N_20689);
xnor U20887 (N_20887,N_20791,N_20683);
xor U20888 (N_20888,N_20726,N_20676);
nor U20889 (N_20889,N_20767,N_20678);
nor U20890 (N_20890,N_20775,N_20604);
or U20891 (N_20891,N_20670,N_20648);
and U20892 (N_20892,N_20710,N_20620);
nor U20893 (N_20893,N_20634,N_20696);
xor U20894 (N_20894,N_20627,N_20714);
and U20895 (N_20895,N_20698,N_20617);
xnor U20896 (N_20896,N_20608,N_20681);
xnor U20897 (N_20897,N_20661,N_20760);
nand U20898 (N_20898,N_20778,N_20691);
xnor U20899 (N_20899,N_20738,N_20795);
or U20900 (N_20900,N_20622,N_20627);
nor U20901 (N_20901,N_20650,N_20680);
and U20902 (N_20902,N_20603,N_20702);
nor U20903 (N_20903,N_20654,N_20622);
nor U20904 (N_20904,N_20793,N_20768);
and U20905 (N_20905,N_20662,N_20609);
nor U20906 (N_20906,N_20666,N_20749);
and U20907 (N_20907,N_20607,N_20776);
xnor U20908 (N_20908,N_20716,N_20623);
and U20909 (N_20909,N_20612,N_20758);
xnor U20910 (N_20910,N_20748,N_20628);
nand U20911 (N_20911,N_20624,N_20601);
nand U20912 (N_20912,N_20784,N_20758);
xor U20913 (N_20913,N_20630,N_20698);
xor U20914 (N_20914,N_20604,N_20723);
nor U20915 (N_20915,N_20774,N_20754);
nand U20916 (N_20916,N_20794,N_20702);
nor U20917 (N_20917,N_20615,N_20797);
xor U20918 (N_20918,N_20667,N_20698);
and U20919 (N_20919,N_20685,N_20627);
and U20920 (N_20920,N_20604,N_20730);
or U20921 (N_20921,N_20610,N_20751);
nor U20922 (N_20922,N_20651,N_20630);
or U20923 (N_20923,N_20642,N_20737);
nand U20924 (N_20924,N_20607,N_20673);
nand U20925 (N_20925,N_20778,N_20768);
nand U20926 (N_20926,N_20666,N_20781);
and U20927 (N_20927,N_20659,N_20711);
xor U20928 (N_20928,N_20607,N_20723);
and U20929 (N_20929,N_20772,N_20723);
and U20930 (N_20930,N_20706,N_20761);
or U20931 (N_20931,N_20737,N_20761);
nand U20932 (N_20932,N_20753,N_20687);
and U20933 (N_20933,N_20609,N_20686);
and U20934 (N_20934,N_20733,N_20632);
nand U20935 (N_20935,N_20656,N_20610);
nand U20936 (N_20936,N_20624,N_20675);
nand U20937 (N_20937,N_20747,N_20610);
nor U20938 (N_20938,N_20766,N_20717);
nor U20939 (N_20939,N_20724,N_20738);
or U20940 (N_20940,N_20688,N_20627);
xor U20941 (N_20941,N_20607,N_20611);
xnor U20942 (N_20942,N_20774,N_20736);
nand U20943 (N_20943,N_20712,N_20720);
nor U20944 (N_20944,N_20607,N_20763);
and U20945 (N_20945,N_20752,N_20681);
or U20946 (N_20946,N_20747,N_20613);
and U20947 (N_20947,N_20771,N_20696);
nor U20948 (N_20948,N_20618,N_20733);
nor U20949 (N_20949,N_20609,N_20705);
xnor U20950 (N_20950,N_20783,N_20627);
nand U20951 (N_20951,N_20644,N_20645);
nor U20952 (N_20952,N_20753,N_20751);
nor U20953 (N_20953,N_20726,N_20718);
or U20954 (N_20954,N_20669,N_20776);
or U20955 (N_20955,N_20657,N_20727);
nor U20956 (N_20956,N_20695,N_20677);
or U20957 (N_20957,N_20684,N_20612);
nand U20958 (N_20958,N_20672,N_20775);
or U20959 (N_20959,N_20731,N_20765);
and U20960 (N_20960,N_20789,N_20736);
xnor U20961 (N_20961,N_20654,N_20776);
or U20962 (N_20962,N_20688,N_20635);
and U20963 (N_20963,N_20675,N_20663);
nor U20964 (N_20964,N_20663,N_20723);
nand U20965 (N_20965,N_20761,N_20798);
nor U20966 (N_20966,N_20608,N_20601);
or U20967 (N_20967,N_20641,N_20659);
or U20968 (N_20968,N_20683,N_20797);
nand U20969 (N_20969,N_20736,N_20623);
nor U20970 (N_20970,N_20654,N_20636);
nor U20971 (N_20971,N_20633,N_20626);
nand U20972 (N_20972,N_20645,N_20708);
and U20973 (N_20973,N_20686,N_20634);
or U20974 (N_20974,N_20699,N_20730);
or U20975 (N_20975,N_20615,N_20703);
and U20976 (N_20976,N_20637,N_20794);
and U20977 (N_20977,N_20703,N_20707);
xnor U20978 (N_20978,N_20755,N_20636);
or U20979 (N_20979,N_20612,N_20616);
nand U20980 (N_20980,N_20788,N_20736);
and U20981 (N_20981,N_20669,N_20730);
or U20982 (N_20982,N_20613,N_20690);
nand U20983 (N_20983,N_20657,N_20623);
nand U20984 (N_20984,N_20776,N_20752);
xnor U20985 (N_20985,N_20717,N_20645);
and U20986 (N_20986,N_20642,N_20674);
or U20987 (N_20987,N_20674,N_20639);
or U20988 (N_20988,N_20621,N_20651);
and U20989 (N_20989,N_20795,N_20799);
nor U20990 (N_20990,N_20730,N_20762);
nand U20991 (N_20991,N_20705,N_20744);
and U20992 (N_20992,N_20775,N_20654);
or U20993 (N_20993,N_20697,N_20699);
nor U20994 (N_20994,N_20678,N_20621);
nand U20995 (N_20995,N_20608,N_20783);
nand U20996 (N_20996,N_20638,N_20661);
nor U20997 (N_20997,N_20715,N_20613);
xnor U20998 (N_20998,N_20724,N_20670);
nor U20999 (N_20999,N_20702,N_20778);
nand U21000 (N_21000,N_20825,N_20991);
xor U21001 (N_21001,N_20901,N_20842);
or U21002 (N_21002,N_20909,N_20806);
nor U21003 (N_21003,N_20926,N_20998);
nor U21004 (N_21004,N_20813,N_20921);
or U21005 (N_21005,N_20963,N_20924);
nor U21006 (N_21006,N_20849,N_20876);
nand U21007 (N_21007,N_20829,N_20830);
and U21008 (N_21008,N_20939,N_20845);
nor U21009 (N_21009,N_20995,N_20967);
or U21010 (N_21010,N_20855,N_20992);
and U21011 (N_21011,N_20871,N_20920);
or U21012 (N_21012,N_20978,N_20917);
nor U21013 (N_21013,N_20893,N_20940);
xnor U21014 (N_21014,N_20905,N_20915);
xor U21015 (N_21015,N_20863,N_20900);
or U21016 (N_21016,N_20951,N_20859);
or U21017 (N_21017,N_20965,N_20867);
xor U21018 (N_21018,N_20885,N_20927);
xor U21019 (N_21019,N_20878,N_20950);
or U21020 (N_21020,N_20890,N_20922);
nor U21021 (N_21021,N_20898,N_20833);
or U21022 (N_21022,N_20862,N_20957);
or U21023 (N_21023,N_20902,N_20961);
xor U21024 (N_21024,N_20932,N_20837);
and U21025 (N_21025,N_20836,N_20895);
or U21026 (N_21026,N_20888,N_20925);
nor U21027 (N_21027,N_20903,N_20912);
nand U21028 (N_21028,N_20834,N_20857);
or U21029 (N_21029,N_20944,N_20962);
and U21030 (N_21030,N_20819,N_20843);
nor U21031 (N_21031,N_20960,N_20820);
nand U21032 (N_21032,N_20931,N_20919);
and U21033 (N_21033,N_20897,N_20838);
nand U21034 (N_21034,N_20841,N_20954);
nand U21035 (N_21035,N_20974,N_20907);
nor U21036 (N_21036,N_20881,N_20937);
xnor U21037 (N_21037,N_20981,N_20993);
xor U21038 (N_21038,N_20948,N_20800);
nor U21039 (N_21039,N_20983,N_20873);
nand U21040 (N_21040,N_20870,N_20977);
xor U21041 (N_21041,N_20914,N_20810);
or U21042 (N_21042,N_20848,N_20953);
nor U21043 (N_21043,N_20935,N_20846);
nor U21044 (N_21044,N_20987,N_20942);
and U21045 (N_21045,N_20990,N_20889);
or U21046 (N_21046,N_20852,N_20858);
nand U21047 (N_21047,N_20984,N_20887);
nand U21048 (N_21048,N_20817,N_20865);
xor U21049 (N_21049,N_20861,N_20807);
xnor U21050 (N_21050,N_20899,N_20997);
nand U21051 (N_21051,N_20853,N_20801);
xnor U21052 (N_21052,N_20938,N_20824);
xnor U21053 (N_21053,N_20856,N_20864);
nor U21054 (N_21054,N_20976,N_20815);
and U21055 (N_21055,N_20959,N_20949);
xnor U21056 (N_21056,N_20989,N_20911);
nand U21057 (N_21057,N_20869,N_20975);
nand U21058 (N_21058,N_20933,N_20928);
or U21059 (N_21059,N_20936,N_20854);
and U21060 (N_21060,N_20886,N_20946);
nor U21061 (N_21061,N_20910,N_20941);
nor U21062 (N_21062,N_20970,N_20958);
or U21063 (N_21063,N_20847,N_20908);
or U21064 (N_21064,N_20956,N_20877);
and U21065 (N_21065,N_20947,N_20929);
xor U21066 (N_21066,N_20966,N_20896);
nor U21067 (N_21067,N_20874,N_20811);
and U21068 (N_21068,N_20916,N_20808);
nand U21069 (N_21069,N_20973,N_20822);
or U21070 (N_21070,N_20969,N_20812);
nand U21071 (N_21071,N_20952,N_20844);
xnor U21072 (N_21072,N_20823,N_20994);
and U21073 (N_21073,N_20883,N_20809);
or U21074 (N_21074,N_20996,N_20804);
xnor U21075 (N_21075,N_20840,N_20979);
or U21076 (N_21076,N_20802,N_20866);
xnor U21077 (N_21077,N_20972,N_20999);
xnor U21078 (N_21078,N_20816,N_20803);
or U21079 (N_21079,N_20832,N_20955);
nand U21080 (N_21080,N_20880,N_20835);
xnor U21081 (N_21081,N_20985,N_20964);
xor U21082 (N_21082,N_20904,N_20988);
xnor U21083 (N_21083,N_20826,N_20872);
nor U21084 (N_21084,N_20818,N_20894);
or U21085 (N_21085,N_20971,N_20930);
nand U21086 (N_21086,N_20906,N_20827);
or U21087 (N_21087,N_20828,N_20879);
nand U21088 (N_21088,N_20891,N_20882);
xnor U21089 (N_21089,N_20884,N_20913);
xor U21090 (N_21090,N_20831,N_20821);
nand U21091 (N_21091,N_20860,N_20980);
and U21092 (N_21092,N_20982,N_20968);
or U21093 (N_21093,N_20918,N_20839);
and U21094 (N_21094,N_20805,N_20868);
nor U21095 (N_21095,N_20943,N_20892);
and U21096 (N_21096,N_20814,N_20851);
or U21097 (N_21097,N_20875,N_20850);
xnor U21098 (N_21098,N_20934,N_20923);
xnor U21099 (N_21099,N_20945,N_20986);
and U21100 (N_21100,N_20894,N_20866);
xnor U21101 (N_21101,N_20979,N_20953);
or U21102 (N_21102,N_20931,N_20966);
nand U21103 (N_21103,N_20878,N_20870);
nand U21104 (N_21104,N_20887,N_20810);
nor U21105 (N_21105,N_20967,N_20944);
nor U21106 (N_21106,N_20906,N_20813);
and U21107 (N_21107,N_20902,N_20854);
or U21108 (N_21108,N_20998,N_20854);
nor U21109 (N_21109,N_20804,N_20897);
nor U21110 (N_21110,N_20803,N_20907);
or U21111 (N_21111,N_20990,N_20839);
or U21112 (N_21112,N_20974,N_20961);
nor U21113 (N_21113,N_20947,N_20979);
nand U21114 (N_21114,N_20900,N_20993);
and U21115 (N_21115,N_20914,N_20833);
nand U21116 (N_21116,N_20810,N_20953);
or U21117 (N_21117,N_20809,N_20844);
and U21118 (N_21118,N_20921,N_20950);
nor U21119 (N_21119,N_20822,N_20803);
nand U21120 (N_21120,N_20919,N_20870);
or U21121 (N_21121,N_20821,N_20850);
and U21122 (N_21122,N_20918,N_20868);
nand U21123 (N_21123,N_20907,N_20918);
or U21124 (N_21124,N_20860,N_20933);
nor U21125 (N_21125,N_20906,N_20924);
nand U21126 (N_21126,N_20805,N_20814);
or U21127 (N_21127,N_20969,N_20874);
xnor U21128 (N_21128,N_20868,N_20940);
and U21129 (N_21129,N_20868,N_20952);
nand U21130 (N_21130,N_20962,N_20900);
nor U21131 (N_21131,N_20974,N_20815);
xor U21132 (N_21132,N_20961,N_20878);
xor U21133 (N_21133,N_20823,N_20989);
nand U21134 (N_21134,N_20914,N_20826);
or U21135 (N_21135,N_20997,N_20954);
nand U21136 (N_21136,N_20971,N_20857);
nand U21137 (N_21137,N_20824,N_20806);
xnor U21138 (N_21138,N_20898,N_20911);
or U21139 (N_21139,N_20957,N_20811);
and U21140 (N_21140,N_20999,N_20947);
nand U21141 (N_21141,N_20937,N_20812);
nand U21142 (N_21142,N_20809,N_20955);
xnor U21143 (N_21143,N_20831,N_20904);
or U21144 (N_21144,N_20803,N_20858);
xor U21145 (N_21145,N_20884,N_20886);
nand U21146 (N_21146,N_20952,N_20916);
or U21147 (N_21147,N_20837,N_20852);
or U21148 (N_21148,N_20970,N_20847);
and U21149 (N_21149,N_20813,N_20890);
nor U21150 (N_21150,N_20948,N_20923);
and U21151 (N_21151,N_20975,N_20903);
xor U21152 (N_21152,N_20925,N_20937);
and U21153 (N_21153,N_20881,N_20802);
nor U21154 (N_21154,N_20884,N_20964);
and U21155 (N_21155,N_20804,N_20845);
xor U21156 (N_21156,N_20919,N_20915);
and U21157 (N_21157,N_20855,N_20957);
and U21158 (N_21158,N_20979,N_20814);
xor U21159 (N_21159,N_20944,N_20984);
or U21160 (N_21160,N_20802,N_20855);
nand U21161 (N_21161,N_20966,N_20978);
or U21162 (N_21162,N_20812,N_20875);
and U21163 (N_21163,N_20821,N_20811);
nand U21164 (N_21164,N_20910,N_20885);
or U21165 (N_21165,N_20973,N_20916);
or U21166 (N_21166,N_20804,N_20910);
nand U21167 (N_21167,N_20990,N_20826);
or U21168 (N_21168,N_20902,N_20878);
or U21169 (N_21169,N_20808,N_20805);
nor U21170 (N_21170,N_20875,N_20963);
nand U21171 (N_21171,N_20825,N_20865);
and U21172 (N_21172,N_20804,N_20883);
nand U21173 (N_21173,N_20903,N_20823);
nor U21174 (N_21174,N_20853,N_20834);
or U21175 (N_21175,N_20891,N_20974);
nand U21176 (N_21176,N_20915,N_20872);
and U21177 (N_21177,N_20982,N_20887);
and U21178 (N_21178,N_20933,N_20876);
xnor U21179 (N_21179,N_20800,N_20884);
nand U21180 (N_21180,N_20918,N_20944);
or U21181 (N_21181,N_20843,N_20820);
nand U21182 (N_21182,N_20834,N_20885);
nor U21183 (N_21183,N_20952,N_20962);
nand U21184 (N_21184,N_20833,N_20972);
or U21185 (N_21185,N_20949,N_20982);
nand U21186 (N_21186,N_20914,N_20938);
nor U21187 (N_21187,N_20859,N_20928);
xnor U21188 (N_21188,N_20820,N_20850);
and U21189 (N_21189,N_20847,N_20879);
xor U21190 (N_21190,N_20988,N_20875);
or U21191 (N_21191,N_20871,N_20998);
or U21192 (N_21192,N_20896,N_20988);
nand U21193 (N_21193,N_20838,N_20987);
or U21194 (N_21194,N_20996,N_20813);
or U21195 (N_21195,N_20986,N_20880);
nand U21196 (N_21196,N_20990,N_20976);
xnor U21197 (N_21197,N_20822,N_20842);
xor U21198 (N_21198,N_20947,N_20828);
nor U21199 (N_21199,N_20984,N_20825);
or U21200 (N_21200,N_21139,N_21127);
and U21201 (N_21201,N_21074,N_21172);
and U21202 (N_21202,N_21148,N_21024);
or U21203 (N_21203,N_21002,N_21063);
xor U21204 (N_21204,N_21113,N_21088);
or U21205 (N_21205,N_21184,N_21035);
nand U21206 (N_21206,N_21106,N_21188);
or U21207 (N_21207,N_21053,N_21175);
nor U21208 (N_21208,N_21160,N_21046);
or U21209 (N_21209,N_21001,N_21022);
or U21210 (N_21210,N_21051,N_21173);
nor U21211 (N_21211,N_21038,N_21043);
xor U21212 (N_21212,N_21055,N_21159);
xnor U21213 (N_21213,N_21198,N_21126);
and U21214 (N_21214,N_21073,N_21199);
nor U21215 (N_21215,N_21177,N_21015);
and U21216 (N_21216,N_21170,N_21109);
and U21217 (N_21217,N_21012,N_21025);
nor U21218 (N_21218,N_21138,N_21026);
nor U21219 (N_21219,N_21179,N_21171);
and U21220 (N_21220,N_21111,N_21009);
nor U21221 (N_21221,N_21101,N_21047);
nor U21222 (N_21222,N_21118,N_21168);
and U21223 (N_21223,N_21189,N_21115);
xnor U21224 (N_21224,N_21069,N_21056);
and U21225 (N_21225,N_21132,N_21041);
xnor U21226 (N_21226,N_21163,N_21122);
nand U21227 (N_21227,N_21124,N_21186);
xnor U21228 (N_21228,N_21049,N_21146);
nor U21229 (N_21229,N_21057,N_21187);
nand U21230 (N_21230,N_21119,N_21104);
xnor U21231 (N_21231,N_21180,N_21037);
and U21232 (N_21232,N_21003,N_21135);
xnor U21233 (N_21233,N_21060,N_21040);
or U21234 (N_21234,N_21013,N_21176);
or U21235 (N_21235,N_21125,N_21108);
and U21236 (N_21236,N_21094,N_21105);
and U21237 (N_21237,N_21102,N_21085);
nor U21238 (N_21238,N_21143,N_21112);
xnor U21239 (N_21239,N_21150,N_21061);
and U21240 (N_21240,N_21082,N_21095);
and U21241 (N_21241,N_21091,N_21190);
and U21242 (N_21242,N_21165,N_21054);
xor U21243 (N_21243,N_21178,N_21029);
xnor U21244 (N_21244,N_21182,N_21000);
and U21245 (N_21245,N_21072,N_21020);
nor U21246 (N_21246,N_21005,N_21117);
nand U21247 (N_21247,N_21092,N_21174);
nand U21248 (N_21248,N_21155,N_21064);
or U21249 (N_21249,N_21083,N_21068);
nand U21250 (N_21250,N_21114,N_21081);
nor U21251 (N_21251,N_21030,N_21097);
xor U21252 (N_21252,N_21169,N_21193);
xor U21253 (N_21253,N_21133,N_21028);
xnor U21254 (N_21254,N_21129,N_21099);
xor U21255 (N_21255,N_21087,N_21027);
nand U21256 (N_21256,N_21075,N_21116);
nor U21257 (N_21257,N_21050,N_21007);
and U21258 (N_21258,N_21077,N_21137);
nand U21259 (N_21259,N_21098,N_21121);
xor U21260 (N_21260,N_21004,N_21036);
nor U21261 (N_21261,N_21164,N_21154);
or U21262 (N_21262,N_21136,N_21142);
and U21263 (N_21263,N_21016,N_21162);
and U21264 (N_21264,N_21079,N_21014);
xor U21265 (N_21265,N_21033,N_21145);
xor U21266 (N_21266,N_21089,N_21058);
xnor U21267 (N_21267,N_21152,N_21048);
and U21268 (N_21268,N_21034,N_21149);
and U21269 (N_21269,N_21044,N_21141);
nor U21270 (N_21270,N_21042,N_21134);
nand U21271 (N_21271,N_21019,N_21130);
nand U21272 (N_21272,N_21144,N_21008);
and U21273 (N_21273,N_21183,N_21181);
nor U21274 (N_21274,N_21062,N_21017);
xor U21275 (N_21275,N_21011,N_21120);
nor U21276 (N_21276,N_21191,N_21157);
and U21277 (N_21277,N_21018,N_21153);
nor U21278 (N_21278,N_21192,N_21093);
xor U21279 (N_21279,N_21021,N_21096);
nand U21280 (N_21280,N_21161,N_21032);
or U21281 (N_21281,N_21103,N_21185);
or U21282 (N_21282,N_21131,N_21123);
and U21283 (N_21283,N_21052,N_21107);
and U21284 (N_21284,N_21065,N_21045);
or U21285 (N_21285,N_21167,N_21156);
xor U21286 (N_21286,N_21194,N_21076);
nand U21287 (N_21287,N_21023,N_21166);
and U21288 (N_21288,N_21070,N_21140);
nor U21289 (N_21289,N_21084,N_21078);
or U21290 (N_21290,N_21080,N_21151);
nand U21291 (N_21291,N_21100,N_21195);
or U21292 (N_21292,N_21006,N_21010);
nor U21293 (N_21293,N_21067,N_21128);
nor U21294 (N_21294,N_21090,N_21158);
and U21295 (N_21295,N_21110,N_21197);
and U21296 (N_21296,N_21086,N_21071);
and U21297 (N_21297,N_21059,N_21031);
and U21298 (N_21298,N_21147,N_21039);
xor U21299 (N_21299,N_21066,N_21196);
nand U21300 (N_21300,N_21027,N_21175);
nor U21301 (N_21301,N_21023,N_21028);
nor U21302 (N_21302,N_21103,N_21089);
xor U21303 (N_21303,N_21086,N_21131);
nand U21304 (N_21304,N_21199,N_21084);
nor U21305 (N_21305,N_21122,N_21195);
nor U21306 (N_21306,N_21173,N_21188);
and U21307 (N_21307,N_21143,N_21091);
and U21308 (N_21308,N_21148,N_21057);
nor U21309 (N_21309,N_21069,N_21010);
xnor U21310 (N_21310,N_21176,N_21030);
nand U21311 (N_21311,N_21121,N_21002);
nand U21312 (N_21312,N_21181,N_21086);
nor U21313 (N_21313,N_21138,N_21137);
or U21314 (N_21314,N_21119,N_21047);
nand U21315 (N_21315,N_21167,N_21100);
xor U21316 (N_21316,N_21081,N_21055);
and U21317 (N_21317,N_21049,N_21160);
nand U21318 (N_21318,N_21005,N_21021);
nand U21319 (N_21319,N_21099,N_21073);
nor U21320 (N_21320,N_21149,N_21005);
nand U21321 (N_21321,N_21070,N_21064);
or U21322 (N_21322,N_21045,N_21173);
and U21323 (N_21323,N_21066,N_21011);
nor U21324 (N_21324,N_21129,N_21170);
or U21325 (N_21325,N_21178,N_21071);
nor U21326 (N_21326,N_21199,N_21165);
or U21327 (N_21327,N_21104,N_21152);
and U21328 (N_21328,N_21033,N_21067);
nor U21329 (N_21329,N_21196,N_21004);
nor U21330 (N_21330,N_21100,N_21196);
xor U21331 (N_21331,N_21030,N_21107);
xnor U21332 (N_21332,N_21086,N_21100);
nor U21333 (N_21333,N_21154,N_21015);
nand U21334 (N_21334,N_21136,N_21002);
nand U21335 (N_21335,N_21071,N_21157);
xor U21336 (N_21336,N_21176,N_21031);
and U21337 (N_21337,N_21057,N_21124);
and U21338 (N_21338,N_21193,N_21125);
xor U21339 (N_21339,N_21114,N_21162);
xor U21340 (N_21340,N_21030,N_21155);
xnor U21341 (N_21341,N_21047,N_21178);
nor U21342 (N_21342,N_21072,N_21028);
or U21343 (N_21343,N_21183,N_21012);
nor U21344 (N_21344,N_21110,N_21019);
nand U21345 (N_21345,N_21183,N_21112);
nand U21346 (N_21346,N_21146,N_21153);
xnor U21347 (N_21347,N_21112,N_21036);
and U21348 (N_21348,N_21094,N_21129);
nor U21349 (N_21349,N_21057,N_21083);
and U21350 (N_21350,N_21009,N_21008);
xor U21351 (N_21351,N_21070,N_21139);
or U21352 (N_21352,N_21053,N_21101);
or U21353 (N_21353,N_21053,N_21115);
xor U21354 (N_21354,N_21094,N_21045);
xor U21355 (N_21355,N_21009,N_21106);
xor U21356 (N_21356,N_21070,N_21010);
and U21357 (N_21357,N_21002,N_21071);
and U21358 (N_21358,N_21022,N_21071);
and U21359 (N_21359,N_21178,N_21028);
nor U21360 (N_21360,N_21059,N_21116);
or U21361 (N_21361,N_21133,N_21199);
nor U21362 (N_21362,N_21098,N_21119);
xor U21363 (N_21363,N_21100,N_21154);
xnor U21364 (N_21364,N_21043,N_21094);
xnor U21365 (N_21365,N_21075,N_21126);
nor U21366 (N_21366,N_21073,N_21102);
and U21367 (N_21367,N_21156,N_21022);
xnor U21368 (N_21368,N_21172,N_21023);
and U21369 (N_21369,N_21036,N_21171);
nand U21370 (N_21370,N_21103,N_21174);
or U21371 (N_21371,N_21118,N_21085);
xor U21372 (N_21372,N_21192,N_21017);
nand U21373 (N_21373,N_21198,N_21024);
nand U21374 (N_21374,N_21089,N_21167);
and U21375 (N_21375,N_21074,N_21029);
nor U21376 (N_21376,N_21091,N_21069);
xnor U21377 (N_21377,N_21011,N_21071);
nand U21378 (N_21378,N_21061,N_21090);
and U21379 (N_21379,N_21072,N_21012);
nand U21380 (N_21380,N_21061,N_21042);
xor U21381 (N_21381,N_21063,N_21004);
or U21382 (N_21382,N_21181,N_21124);
and U21383 (N_21383,N_21086,N_21098);
nor U21384 (N_21384,N_21190,N_21117);
xor U21385 (N_21385,N_21059,N_21173);
nand U21386 (N_21386,N_21114,N_21045);
nor U21387 (N_21387,N_21184,N_21143);
and U21388 (N_21388,N_21152,N_21149);
nor U21389 (N_21389,N_21094,N_21075);
or U21390 (N_21390,N_21098,N_21165);
nand U21391 (N_21391,N_21012,N_21123);
or U21392 (N_21392,N_21034,N_21093);
nor U21393 (N_21393,N_21150,N_21024);
nor U21394 (N_21394,N_21112,N_21100);
and U21395 (N_21395,N_21145,N_21152);
or U21396 (N_21396,N_21085,N_21101);
xnor U21397 (N_21397,N_21155,N_21016);
nand U21398 (N_21398,N_21034,N_21056);
nand U21399 (N_21399,N_21072,N_21133);
or U21400 (N_21400,N_21237,N_21304);
nand U21401 (N_21401,N_21272,N_21323);
nand U21402 (N_21402,N_21388,N_21344);
nand U21403 (N_21403,N_21274,N_21303);
or U21404 (N_21404,N_21213,N_21391);
xnor U21405 (N_21405,N_21340,N_21269);
xor U21406 (N_21406,N_21236,N_21318);
and U21407 (N_21407,N_21392,N_21308);
nand U21408 (N_21408,N_21216,N_21345);
nand U21409 (N_21409,N_21266,N_21399);
and U21410 (N_21410,N_21380,N_21370);
and U21411 (N_21411,N_21238,N_21267);
and U21412 (N_21412,N_21214,N_21288);
nor U21413 (N_21413,N_21351,N_21220);
nand U21414 (N_21414,N_21273,N_21261);
or U21415 (N_21415,N_21242,N_21217);
nor U21416 (N_21416,N_21275,N_21229);
and U21417 (N_21417,N_21330,N_21282);
xnor U21418 (N_21418,N_21290,N_21353);
and U21419 (N_21419,N_21324,N_21224);
nor U21420 (N_21420,N_21383,N_21257);
xnor U21421 (N_21421,N_21221,N_21270);
xor U21422 (N_21422,N_21325,N_21228);
nand U21423 (N_21423,N_21332,N_21377);
xor U21424 (N_21424,N_21295,N_21320);
xnor U21425 (N_21425,N_21335,N_21255);
or U21426 (N_21426,N_21243,N_21227);
and U21427 (N_21427,N_21240,N_21309);
or U21428 (N_21428,N_21210,N_21253);
xor U21429 (N_21429,N_21287,N_21393);
nand U21430 (N_21430,N_21381,N_21299);
nand U21431 (N_21431,N_21311,N_21336);
and U21432 (N_21432,N_21327,N_21293);
and U21433 (N_21433,N_21375,N_21204);
nand U21434 (N_21434,N_21235,N_21362);
xnor U21435 (N_21435,N_21306,N_21231);
or U21436 (N_21436,N_21321,N_21250);
and U21437 (N_21437,N_21346,N_21301);
or U21438 (N_21438,N_21387,N_21305);
or U21439 (N_21439,N_21200,N_21222);
or U21440 (N_21440,N_21209,N_21294);
and U21441 (N_21441,N_21234,N_21285);
nand U21442 (N_21442,N_21208,N_21349);
and U21443 (N_21443,N_21202,N_21252);
and U21444 (N_21444,N_21249,N_21331);
or U21445 (N_21445,N_21279,N_21302);
xor U21446 (N_21446,N_21355,N_21394);
xor U21447 (N_21447,N_21211,N_21310);
or U21448 (N_21448,N_21296,N_21322);
or U21449 (N_21449,N_21260,N_21339);
or U21450 (N_21450,N_21312,N_21374);
xnor U21451 (N_21451,N_21280,N_21360);
and U21452 (N_21452,N_21368,N_21307);
or U21453 (N_21453,N_21218,N_21247);
nand U21454 (N_21454,N_21365,N_21367);
and U21455 (N_21455,N_21315,N_21244);
nor U21456 (N_21456,N_21265,N_21230);
or U21457 (N_21457,N_21215,N_21263);
and U21458 (N_21458,N_21276,N_21254);
nand U21459 (N_21459,N_21379,N_21319);
or U21460 (N_21460,N_21378,N_21386);
nand U21461 (N_21461,N_21334,N_21212);
or U21462 (N_21462,N_21358,N_21205);
or U21463 (N_21463,N_21291,N_21326);
xor U21464 (N_21464,N_21384,N_21248);
nand U21465 (N_21465,N_21366,N_21354);
and U21466 (N_21466,N_21264,N_21256);
nand U21467 (N_21467,N_21298,N_21382);
and U21468 (N_21468,N_21259,N_21233);
nor U21469 (N_21469,N_21328,N_21300);
and U21470 (N_21470,N_21348,N_21363);
xnor U21471 (N_21471,N_21373,N_21350);
and U21472 (N_21472,N_21385,N_21232);
or U21473 (N_21473,N_21245,N_21284);
xor U21474 (N_21474,N_21219,N_21239);
xnor U21475 (N_21475,N_21333,N_21277);
xor U21476 (N_21476,N_21289,N_21342);
or U21477 (N_21477,N_21357,N_21223);
xor U21478 (N_21478,N_21395,N_21203);
or U21479 (N_21479,N_21397,N_21396);
xor U21480 (N_21480,N_21268,N_21206);
xnor U21481 (N_21481,N_21369,N_21372);
nand U21482 (N_21482,N_21292,N_21359);
xor U21483 (N_21483,N_21241,N_21390);
or U21484 (N_21484,N_21297,N_21389);
nand U21485 (N_21485,N_21317,N_21341);
nand U21486 (N_21486,N_21371,N_21226);
nand U21487 (N_21487,N_21225,N_21246);
and U21488 (N_21488,N_21316,N_21364);
nor U21489 (N_21489,N_21361,N_21258);
nand U21490 (N_21490,N_21201,N_21352);
and U21491 (N_21491,N_21278,N_21356);
nand U21492 (N_21492,N_21329,N_21313);
and U21493 (N_21493,N_21207,N_21338);
nand U21494 (N_21494,N_21314,N_21271);
nand U21495 (N_21495,N_21343,N_21262);
nand U21496 (N_21496,N_21376,N_21283);
or U21497 (N_21497,N_21347,N_21251);
and U21498 (N_21498,N_21286,N_21337);
or U21499 (N_21499,N_21398,N_21281);
nand U21500 (N_21500,N_21255,N_21243);
nor U21501 (N_21501,N_21242,N_21222);
nand U21502 (N_21502,N_21234,N_21316);
nand U21503 (N_21503,N_21265,N_21280);
xor U21504 (N_21504,N_21375,N_21360);
nor U21505 (N_21505,N_21353,N_21206);
xnor U21506 (N_21506,N_21266,N_21386);
nand U21507 (N_21507,N_21278,N_21315);
xnor U21508 (N_21508,N_21231,N_21327);
nand U21509 (N_21509,N_21379,N_21306);
or U21510 (N_21510,N_21331,N_21397);
xnor U21511 (N_21511,N_21310,N_21212);
and U21512 (N_21512,N_21215,N_21271);
and U21513 (N_21513,N_21242,N_21325);
xor U21514 (N_21514,N_21367,N_21265);
xor U21515 (N_21515,N_21331,N_21389);
and U21516 (N_21516,N_21355,N_21318);
or U21517 (N_21517,N_21204,N_21232);
or U21518 (N_21518,N_21320,N_21258);
nand U21519 (N_21519,N_21344,N_21253);
or U21520 (N_21520,N_21319,N_21310);
nand U21521 (N_21521,N_21219,N_21264);
and U21522 (N_21522,N_21291,N_21252);
nor U21523 (N_21523,N_21352,N_21296);
or U21524 (N_21524,N_21242,N_21264);
nor U21525 (N_21525,N_21367,N_21202);
nor U21526 (N_21526,N_21234,N_21280);
nor U21527 (N_21527,N_21367,N_21230);
nand U21528 (N_21528,N_21273,N_21251);
xnor U21529 (N_21529,N_21338,N_21358);
nand U21530 (N_21530,N_21248,N_21230);
nor U21531 (N_21531,N_21352,N_21357);
xnor U21532 (N_21532,N_21259,N_21295);
nor U21533 (N_21533,N_21218,N_21351);
or U21534 (N_21534,N_21241,N_21311);
xor U21535 (N_21535,N_21327,N_21215);
nand U21536 (N_21536,N_21247,N_21274);
nand U21537 (N_21537,N_21389,N_21356);
and U21538 (N_21538,N_21375,N_21379);
nor U21539 (N_21539,N_21375,N_21382);
xnor U21540 (N_21540,N_21369,N_21204);
xor U21541 (N_21541,N_21329,N_21320);
nor U21542 (N_21542,N_21277,N_21201);
or U21543 (N_21543,N_21267,N_21372);
nand U21544 (N_21544,N_21394,N_21348);
or U21545 (N_21545,N_21374,N_21324);
nand U21546 (N_21546,N_21243,N_21331);
nor U21547 (N_21547,N_21326,N_21394);
or U21548 (N_21548,N_21237,N_21290);
nand U21549 (N_21549,N_21351,N_21371);
or U21550 (N_21550,N_21283,N_21254);
xnor U21551 (N_21551,N_21323,N_21394);
nor U21552 (N_21552,N_21369,N_21358);
nor U21553 (N_21553,N_21206,N_21263);
nand U21554 (N_21554,N_21338,N_21284);
nor U21555 (N_21555,N_21287,N_21205);
or U21556 (N_21556,N_21307,N_21369);
nand U21557 (N_21557,N_21238,N_21231);
or U21558 (N_21558,N_21221,N_21304);
nor U21559 (N_21559,N_21205,N_21362);
and U21560 (N_21560,N_21353,N_21292);
nand U21561 (N_21561,N_21257,N_21202);
and U21562 (N_21562,N_21201,N_21288);
nor U21563 (N_21563,N_21207,N_21373);
nand U21564 (N_21564,N_21248,N_21240);
xor U21565 (N_21565,N_21246,N_21278);
nand U21566 (N_21566,N_21270,N_21355);
and U21567 (N_21567,N_21326,N_21318);
nor U21568 (N_21568,N_21203,N_21331);
xor U21569 (N_21569,N_21379,N_21329);
or U21570 (N_21570,N_21346,N_21294);
nor U21571 (N_21571,N_21256,N_21346);
nand U21572 (N_21572,N_21247,N_21294);
and U21573 (N_21573,N_21345,N_21340);
nand U21574 (N_21574,N_21268,N_21336);
and U21575 (N_21575,N_21232,N_21337);
and U21576 (N_21576,N_21281,N_21248);
nand U21577 (N_21577,N_21350,N_21252);
or U21578 (N_21578,N_21226,N_21382);
nand U21579 (N_21579,N_21267,N_21384);
nor U21580 (N_21580,N_21399,N_21228);
or U21581 (N_21581,N_21270,N_21362);
xnor U21582 (N_21582,N_21367,N_21386);
and U21583 (N_21583,N_21266,N_21213);
nand U21584 (N_21584,N_21345,N_21351);
and U21585 (N_21585,N_21229,N_21243);
and U21586 (N_21586,N_21268,N_21338);
xnor U21587 (N_21587,N_21352,N_21271);
and U21588 (N_21588,N_21325,N_21379);
nor U21589 (N_21589,N_21338,N_21345);
xnor U21590 (N_21590,N_21348,N_21259);
xnor U21591 (N_21591,N_21246,N_21217);
or U21592 (N_21592,N_21210,N_21391);
or U21593 (N_21593,N_21316,N_21366);
nand U21594 (N_21594,N_21392,N_21210);
and U21595 (N_21595,N_21280,N_21283);
or U21596 (N_21596,N_21364,N_21243);
nand U21597 (N_21597,N_21398,N_21375);
nor U21598 (N_21598,N_21211,N_21351);
xor U21599 (N_21599,N_21262,N_21297);
or U21600 (N_21600,N_21500,N_21440);
or U21601 (N_21601,N_21400,N_21401);
or U21602 (N_21602,N_21544,N_21411);
nor U21603 (N_21603,N_21415,N_21470);
and U21604 (N_21604,N_21468,N_21593);
or U21605 (N_21605,N_21536,N_21465);
and U21606 (N_21606,N_21487,N_21574);
or U21607 (N_21607,N_21432,N_21493);
xor U21608 (N_21608,N_21555,N_21525);
nor U21609 (N_21609,N_21418,N_21598);
and U21610 (N_21610,N_21515,N_21537);
nor U21611 (N_21611,N_21433,N_21522);
nand U21612 (N_21612,N_21452,N_21494);
nor U21613 (N_21613,N_21457,N_21510);
or U21614 (N_21614,N_21471,N_21558);
and U21615 (N_21615,N_21516,N_21480);
or U21616 (N_21616,N_21430,N_21526);
xor U21617 (N_21617,N_21429,N_21581);
nor U21618 (N_21618,N_21413,N_21441);
nor U21619 (N_21619,N_21595,N_21521);
nand U21620 (N_21620,N_21504,N_21548);
and U21621 (N_21621,N_21560,N_21421);
xor U21622 (N_21622,N_21546,N_21532);
nand U21623 (N_21623,N_21518,N_21442);
nor U21624 (N_21624,N_21476,N_21507);
or U21625 (N_21625,N_21424,N_21583);
or U21626 (N_21626,N_21431,N_21478);
nand U21627 (N_21627,N_21520,N_21408);
xor U21628 (N_21628,N_21576,N_21423);
or U21629 (N_21629,N_21445,N_21416);
or U21630 (N_21630,N_21466,N_21570);
xnor U21631 (N_21631,N_21483,N_21577);
nand U21632 (N_21632,N_21508,N_21488);
or U21633 (N_21633,N_21556,N_21502);
nand U21634 (N_21634,N_21410,N_21417);
xor U21635 (N_21635,N_21531,N_21551);
and U21636 (N_21636,N_21450,N_21509);
or U21637 (N_21637,N_21517,N_21484);
or U21638 (N_21638,N_21590,N_21464);
xor U21639 (N_21639,N_21584,N_21588);
nor U21640 (N_21640,N_21427,N_21420);
or U21641 (N_21641,N_21428,N_21477);
and U21642 (N_21642,N_21406,N_21527);
xor U21643 (N_21643,N_21565,N_21578);
or U21644 (N_21644,N_21535,N_21412);
nor U21645 (N_21645,N_21414,N_21472);
xor U21646 (N_21646,N_21454,N_21564);
or U21647 (N_21647,N_21482,N_21563);
nand U21648 (N_21648,N_21550,N_21485);
nand U21649 (N_21649,N_21512,N_21486);
or U21650 (N_21650,N_21443,N_21462);
or U21651 (N_21651,N_21497,N_21403);
nand U21652 (N_21652,N_21538,N_21467);
and U21653 (N_21653,N_21491,N_21597);
nand U21654 (N_21654,N_21419,N_21456);
nand U21655 (N_21655,N_21503,N_21501);
or U21656 (N_21656,N_21547,N_21489);
xor U21657 (N_21657,N_21409,N_21498);
and U21658 (N_21658,N_21586,N_21449);
nor U21659 (N_21659,N_21552,N_21529);
or U21660 (N_21660,N_21446,N_21549);
nand U21661 (N_21661,N_21425,N_21458);
and U21662 (N_21662,N_21539,N_21553);
nor U21663 (N_21663,N_21533,N_21463);
nand U21664 (N_21664,N_21479,N_21474);
xnor U21665 (N_21665,N_21437,N_21455);
nand U21666 (N_21666,N_21505,N_21451);
or U21667 (N_21667,N_21545,N_21575);
xnor U21668 (N_21668,N_21591,N_21438);
nor U21669 (N_21669,N_21436,N_21435);
or U21670 (N_21670,N_21530,N_21542);
nand U21671 (N_21671,N_21422,N_21534);
and U21672 (N_21672,N_21519,N_21434);
nor U21673 (N_21673,N_21571,N_21475);
xnor U21674 (N_21674,N_21543,N_21554);
nand U21675 (N_21675,N_21426,N_21459);
or U21676 (N_21676,N_21562,N_21573);
and U21677 (N_21677,N_21447,N_21481);
or U21678 (N_21678,N_21405,N_21566);
nor U21679 (N_21679,N_21524,N_21499);
xnor U21680 (N_21680,N_21492,N_21585);
nor U21681 (N_21681,N_21568,N_21592);
xor U21682 (N_21682,N_21580,N_21582);
nand U21683 (N_21683,N_21523,N_21513);
xnor U21684 (N_21684,N_21453,N_21448);
nand U21685 (N_21685,N_21596,N_21579);
or U21686 (N_21686,N_21557,N_21589);
nor U21687 (N_21687,N_21473,N_21439);
nand U21688 (N_21688,N_21402,N_21444);
and U21689 (N_21689,N_21490,N_21599);
nand U21690 (N_21690,N_21460,N_21404);
and U21691 (N_21691,N_21469,N_21506);
and U21692 (N_21692,N_21461,N_21561);
or U21693 (N_21693,N_21495,N_21511);
and U21694 (N_21694,N_21514,N_21496);
nand U21695 (N_21695,N_21572,N_21594);
xnor U21696 (N_21696,N_21567,N_21528);
nor U21697 (N_21697,N_21587,N_21559);
xnor U21698 (N_21698,N_21541,N_21540);
nor U21699 (N_21699,N_21407,N_21569);
nor U21700 (N_21700,N_21596,N_21423);
xor U21701 (N_21701,N_21445,N_21412);
or U21702 (N_21702,N_21489,N_21550);
xor U21703 (N_21703,N_21520,N_21490);
nand U21704 (N_21704,N_21434,N_21540);
or U21705 (N_21705,N_21429,N_21465);
xnor U21706 (N_21706,N_21419,N_21487);
or U21707 (N_21707,N_21517,N_21503);
nor U21708 (N_21708,N_21427,N_21505);
nor U21709 (N_21709,N_21554,N_21469);
nor U21710 (N_21710,N_21462,N_21494);
or U21711 (N_21711,N_21425,N_21492);
or U21712 (N_21712,N_21570,N_21510);
or U21713 (N_21713,N_21434,N_21493);
nand U21714 (N_21714,N_21524,N_21459);
and U21715 (N_21715,N_21558,N_21544);
nand U21716 (N_21716,N_21515,N_21544);
or U21717 (N_21717,N_21513,N_21499);
or U21718 (N_21718,N_21599,N_21427);
and U21719 (N_21719,N_21597,N_21439);
nor U21720 (N_21720,N_21426,N_21564);
nor U21721 (N_21721,N_21530,N_21457);
xnor U21722 (N_21722,N_21522,N_21475);
or U21723 (N_21723,N_21524,N_21419);
xor U21724 (N_21724,N_21538,N_21459);
and U21725 (N_21725,N_21560,N_21428);
nand U21726 (N_21726,N_21558,N_21556);
or U21727 (N_21727,N_21584,N_21435);
or U21728 (N_21728,N_21488,N_21449);
nor U21729 (N_21729,N_21457,N_21475);
nand U21730 (N_21730,N_21423,N_21478);
or U21731 (N_21731,N_21445,N_21518);
and U21732 (N_21732,N_21418,N_21539);
nor U21733 (N_21733,N_21565,N_21518);
or U21734 (N_21734,N_21595,N_21553);
and U21735 (N_21735,N_21420,N_21459);
or U21736 (N_21736,N_21453,N_21532);
nand U21737 (N_21737,N_21479,N_21561);
or U21738 (N_21738,N_21528,N_21470);
or U21739 (N_21739,N_21543,N_21438);
or U21740 (N_21740,N_21545,N_21506);
xor U21741 (N_21741,N_21551,N_21529);
nor U21742 (N_21742,N_21438,N_21497);
xnor U21743 (N_21743,N_21447,N_21494);
nand U21744 (N_21744,N_21577,N_21546);
or U21745 (N_21745,N_21436,N_21525);
or U21746 (N_21746,N_21598,N_21538);
or U21747 (N_21747,N_21489,N_21498);
and U21748 (N_21748,N_21555,N_21580);
nand U21749 (N_21749,N_21428,N_21546);
or U21750 (N_21750,N_21516,N_21423);
and U21751 (N_21751,N_21539,N_21422);
xnor U21752 (N_21752,N_21528,N_21415);
nand U21753 (N_21753,N_21593,N_21450);
nand U21754 (N_21754,N_21472,N_21424);
nand U21755 (N_21755,N_21575,N_21556);
nor U21756 (N_21756,N_21481,N_21475);
nand U21757 (N_21757,N_21594,N_21414);
nand U21758 (N_21758,N_21510,N_21437);
xnor U21759 (N_21759,N_21402,N_21545);
xor U21760 (N_21760,N_21598,N_21475);
and U21761 (N_21761,N_21470,N_21406);
or U21762 (N_21762,N_21461,N_21490);
and U21763 (N_21763,N_21564,N_21442);
or U21764 (N_21764,N_21597,N_21565);
nand U21765 (N_21765,N_21426,N_21420);
nand U21766 (N_21766,N_21557,N_21499);
xor U21767 (N_21767,N_21449,N_21509);
nor U21768 (N_21768,N_21525,N_21469);
nor U21769 (N_21769,N_21596,N_21555);
and U21770 (N_21770,N_21573,N_21553);
xor U21771 (N_21771,N_21521,N_21564);
nor U21772 (N_21772,N_21492,N_21404);
or U21773 (N_21773,N_21469,N_21550);
nand U21774 (N_21774,N_21463,N_21579);
or U21775 (N_21775,N_21539,N_21554);
xnor U21776 (N_21776,N_21558,N_21408);
and U21777 (N_21777,N_21535,N_21488);
or U21778 (N_21778,N_21586,N_21453);
and U21779 (N_21779,N_21598,N_21592);
xor U21780 (N_21780,N_21437,N_21436);
nor U21781 (N_21781,N_21453,N_21479);
xnor U21782 (N_21782,N_21493,N_21522);
and U21783 (N_21783,N_21429,N_21485);
xnor U21784 (N_21784,N_21494,N_21433);
nand U21785 (N_21785,N_21482,N_21500);
or U21786 (N_21786,N_21459,N_21441);
nor U21787 (N_21787,N_21599,N_21560);
or U21788 (N_21788,N_21447,N_21523);
and U21789 (N_21789,N_21540,N_21565);
nor U21790 (N_21790,N_21419,N_21448);
or U21791 (N_21791,N_21421,N_21509);
nor U21792 (N_21792,N_21509,N_21516);
xnor U21793 (N_21793,N_21575,N_21483);
nand U21794 (N_21794,N_21461,N_21426);
xor U21795 (N_21795,N_21557,N_21516);
and U21796 (N_21796,N_21527,N_21507);
nand U21797 (N_21797,N_21443,N_21486);
nor U21798 (N_21798,N_21404,N_21456);
or U21799 (N_21799,N_21574,N_21523);
and U21800 (N_21800,N_21656,N_21765);
xor U21801 (N_21801,N_21710,N_21706);
or U21802 (N_21802,N_21636,N_21603);
nand U21803 (N_21803,N_21642,N_21608);
and U21804 (N_21804,N_21663,N_21659);
and U21805 (N_21805,N_21627,N_21761);
nand U21806 (N_21806,N_21776,N_21707);
nand U21807 (N_21807,N_21641,N_21673);
or U21808 (N_21808,N_21749,N_21647);
nor U21809 (N_21809,N_21687,N_21668);
nand U21810 (N_21810,N_21727,N_21719);
nor U21811 (N_21811,N_21624,N_21681);
nor U21812 (N_21812,N_21733,N_21728);
nor U21813 (N_21813,N_21746,N_21742);
or U21814 (N_21814,N_21760,N_21700);
or U21815 (N_21815,N_21726,N_21714);
nand U21816 (N_21816,N_21633,N_21698);
and U21817 (N_21817,N_21721,N_21613);
or U21818 (N_21818,N_21783,N_21737);
xnor U21819 (N_21819,N_21601,N_21614);
nand U21820 (N_21820,N_21799,N_21638);
xor U21821 (N_21821,N_21735,N_21669);
nor U21822 (N_21822,N_21688,N_21650);
nor U21823 (N_21823,N_21731,N_21748);
and U21824 (N_21824,N_21685,N_21712);
or U21825 (N_21825,N_21632,N_21678);
and U21826 (N_21826,N_21730,N_21747);
xor U21827 (N_21827,N_21606,N_21766);
or U21828 (N_21828,N_21743,N_21779);
nand U21829 (N_21829,N_21769,N_21630);
nand U21830 (N_21830,N_21716,N_21757);
and U21831 (N_21831,N_21695,N_21657);
nor U21832 (N_21832,N_21792,N_21684);
xnor U21833 (N_21833,N_21751,N_21738);
and U21834 (N_21834,N_21639,N_21618);
xnor U21835 (N_21835,N_21628,N_21672);
or U21836 (N_21836,N_21750,N_21600);
and U21837 (N_21837,N_21649,N_21788);
nor U21838 (N_21838,N_21785,N_21696);
xnor U21839 (N_21839,N_21640,N_21789);
nor U21840 (N_21840,N_21667,N_21625);
xor U21841 (N_21841,N_21755,N_21637);
and U21842 (N_21842,N_21604,N_21736);
nor U21843 (N_21843,N_21619,N_21741);
xor U21844 (N_21844,N_21623,N_21715);
nand U21845 (N_21845,N_21734,N_21605);
nand U21846 (N_21846,N_21772,N_21708);
nor U21847 (N_21847,N_21732,N_21771);
and U21848 (N_21848,N_21790,N_21677);
and U21849 (N_21849,N_21683,N_21654);
or U21850 (N_21850,N_21781,N_21724);
xor U21851 (N_21851,N_21671,N_21674);
nor U21852 (N_21852,N_21795,N_21713);
nand U21853 (N_21853,N_21758,N_21768);
nand U21854 (N_21854,N_21645,N_21648);
or U21855 (N_21855,N_21665,N_21689);
xor U21856 (N_21856,N_21611,N_21609);
and U21857 (N_21857,N_21626,N_21753);
nand U21858 (N_21858,N_21703,N_21690);
nand U21859 (N_21859,N_21660,N_21679);
nand U21860 (N_21860,N_21631,N_21786);
or U21861 (N_21861,N_21740,N_21759);
nor U21862 (N_21862,N_21697,N_21782);
or U21863 (N_21863,N_21744,N_21644);
nand U21864 (N_21864,N_21770,N_21774);
or U21865 (N_21865,N_21691,N_21717);
nand U21866 (N_21866,N_21701,N_21686);
xor U21867 (N_21867,N_21777,N_21763);
or U21868 (N_21868,N_21620,N_21797);
nand U21869 (N_21869,N_21796,N_21780);
nor U21870 (N_21870,N_21702,N_21615);
or U21871 (N_21871,N_21670,N_21752);
nor U21872 (N_21872,N_21711,N_21622);
and U21873 (N_21873,N_21791,N_21699);
or U21874 (N_21874,N_21617,N_21662);
or U21875 (N_21875,N_21661,N_21655);
nand U21876 (N_21876,N_21798,N_21704);
nand U21877 (N_21877,N_21794,N_21718);
or U21878 (N_21878,N_21653,N_21725);
xnor U21879 (N_21879,N_21666,N_21705);
and U21880 (N_21880,N_21682,N_21767);
nand U21881 (N_21881,N_21646,N_21739);
nor U21882 (N_21882,N_21651,N_21692);
or U21883 (N_21883,N_21754,N_21756);
nand U21884 (N_21884,N_21778,N_21773);
nor U21885 (N_21885,N_21745,N_21762);
nand U21886 (N_21886,N_21729,N_21629);
nor U21887 (N_21887,N_21680,N_21787);
nand U21888 (N_21888,N_21722,N_21602);
or U21889 (N_21889,N_21607,N_21610);
nor U21890 (N_21890,N_21720,N_21643);
nor U21891 (N_21891,N_21621,N_21652);
nand U21892 (N_21892,N_21612,N_21764);
and U21893 (N_21893,N_21723,N_21784);
or U21894 (N_21894,N_21793,N_21664);
nand U21895 (N_21895,N_21775,N_21658);
nor U21896 (N_21896,N_21634,N_21675);
nand U21897 (N_21897,N_21616,N_21676);
nand U21898 (N_21898,N_21694,N_21709);
and U21899 (N_21899,N_21635,N_21693);
xnor U21900 (N_21900,N_21610,N_21622);
nand U21901 (N_21901,N_21617,N_21677);
and U21902 (N_21902,N_21649,N_21732);
or U21903 (N_21903,N_21654,N_21647);
nand U21904 (N_21904,N_21792,N_21726);
or U21905 (N_21905,N_21619,N_21706);
or U21906 (N_21906,N_21673,N_21768);
nand U21907 (N_21907,N_21677,N_21650);
nand U21908 (N_21908,N_21765,N_21761);
nand U21909 (N_21909,N_21726,N_21795);
xnor U21910 (N_21910,N_21782,N_21738);
xnor U21911 (N_21911,N_21713,N_21631);
nor U21912 (N_21912,N_21769,N_21738);
nor U21913 (N_21913,N_21794,N_21703);
xor U21914 (N_21914,N_21675,N_21790);
and U21915 (N_21915,N_21640,N_21657);
nand U21916 (N_21916,N_21757,N_21660);
nand U21917 (N_21917,N_21699,N_21626);
nand U21918 (N_21918,N_21729,N_21665);
and U21919 (N_21919,N_21694,N_21624);
and U21920 (N_21920,N_21658,N_21752);
xor U21921 (N_21921,N_21784,N_21675);
or U21922 (N_21922,N_21723,N_21696);
or U21923 (N_21923,N_21671,N_21709);
nand U21924 (N_21924,N_21707,N_21640);
nand U21925 (N_21925,N_21711,N_21754);
and U21926 (N_21926,N_21608,N_21610);
and U21927 (N_21927,N_21662,N_21657);
nor U21928 (N_21928,N_21765,N_21740);
nor U21929 (N_21929,N_21736,N_21693);
or U21930 (N_21930,N_21707,N_21756);
and U21931 (N_21931,N_21783,N_21653);
xnor U21932 (N_21932,N_21768,N_21747);
nand U21933 (N_21933,N_21707,N_21701);
and U21934 (N_21934,N_21665,N_21701);
and U21935 (N_21935,N_21663,N_21746);
nand U21936 (N_21936,N_21709,N_21668);
xor U21937 (N_21937,N_21757,N_21752);
nor U21938 (N_21938,N_21703,N_21726);
xnor U21939 (N_21939,N_21646,N_21632);
or U21940 (N_21940,N_21798,N_21674);
and U21941 (N_21941,N_21783,N_21654);
or U21942 (N_21942,N_21661,N_21639);
or U21943 (N_21943,N_21612,N_21691);
or U21944 (N_21944,N_21758,N_21684);
nand U21945 (N_21945,N_21772,N_21794);
or U21946 (N_21946,N_21769,N_21656);
nand U21947 (N_21947,N_21798,N_21743);
nand U21948 (N_21948,N_21683,N_21656);
or U21949 (N_21949,N_21670,N_21794);
or U21950 (N_21950,N_21711,N_21764);
and U21951 (N_21951,N_21708,N_21640);
nor U21952 (N_21952,N_21667,N_21607);
xor U21953 (N_21953,N_21724,N_21767);
nor U21954 (N_21954,N_21678,N_21714);
and U21955 (N_21955,N_21723,N_21778);
nor U21956 (N_21956,N_21701,N_21625);
or U21957 (N_21957,N_21739,N_21668);
and U21958 (N_21958,N_21785,N_21766);
nor U21959 (N_21959,N_21721,N_21730);
xnor U21960 (N_21960,N_21660,N_21756);
or U21961 (N_21961,N_21644,N_21663);
nand U21962 (N_21962,N_21667,N_21741);
and U21963 (N_21963,N_21667,N_21747);
nand U21964 (N_21964,N_21690,N_21664);
nand U21965 (N_21965,N_21789,N_21696);
and U21966 (N_21966,N_21620,N_21705);
nand U21967 (N_21967,N_21657,N_21795);
xnor U21968 (N_21968,N_21763,N_21771);
and U21969 (N_21969,N_21735,N_21668);
or U21970 (N_21970,N_21691,N_21790);
nand U21971 (N_21971,N_21652,N_21641);
nand U21972 (N_21972,N_21686,N_21747);
or U21973 (N_21973,N_21692,N_21799);
or U21974 (N_21974,N_21618,N_21695);
nand U21975 (N_21975,N_21601,N_21622);
or U21976 (N_21976,N_21719,N_21700);
and U21977 (N_21977,N_21608,N_21736);
xnor U21978 (N_21978,N_21784,N_21752);
xnor U21979 (N_21979,N_21710,N_21707);
xnor U21980 (N_21980,N_21723,N_21781);
xor U21981 (N_21981,N_21612,N_21617);
nor U21982 (N_21982,N_21733,N_21720);
and U21983 (N_21983,N_21651,N_21756);
or U21984 (N_21984,N_21798,N_21651);
xnor U21985 (N_21985,N_21630,N_21736);
nand U21986 (N_21986,N_21694,N_21783);
xor U21987 (N_21987,N_21773,N_21621);
xor U21988 (N_21988,N_21790,N_21725);
or U21989 (N_21989,N_21627,N_21738);
nor U21990 (N_21990,N_21669,N_21707);
nor U21991 (N_21991,N_21650,N_21682);
nor U21992 (N_21992,N_21731,N_21698);
nor U21993 (N_21993,N_21775,N_21788);
xor U21994 (N_21994,N_21767,N_21749);
nor U21995 (N_21995,N_21683,N_21700);
xor U21996 (N_21996,N_21753,N_21715);
xnor U21997 (N_21997,N_21733,N_21777);
and U21998 (N_21998,N_21752,N_21620);
nor U21999 (N_21999,N_21719,N_21699);
xnor U22000 (N_22000,N_21819,N_21916);
nor U22001 (N_22001,N_21977,N_21913);
nand U22002 (N_22002,N_21866,N_21828);
or U22003 (N_22003,N_21893,N_21870);
nand U22004 (N_22004,N_21938,N_21958);
and U22005 (N_22005,N_21848,N_21822);
or U22006 (N_22006,N_21820,N_21917);
nand U22007 (N_22007,N_21937,N_21817);
and U22008 (N_22008,N_21858,N_21874);
and U22009 (N_22009,N_21998,N_21800);
nand U22010 (N_22010,N_21924,N_21933);
xor U22011 (N_22011,N_21824,N_21871);
nor U22012 (N_22012,N_21829,N_21997);
xnor U22013 (N_22013,N_21966,N_21941);
and U22014 (N_22014,N_21812,N_21903);
nand U22015 (N_22015,N_21880,N_21897);
nand U22016 (N_22016,N_21877,N_21885);
and U22017 (N_22017,N_21801,N_21914);
and U22018 (N_22018,N_21811,N_21864);
nor U22019 (N_22019,N_21978,N_21845);
nand U22020 (N_22020,N_21849,N_21869);
or U22021 (N_22021,N_21971,N_21813);
or U22022 (N_22022,N_21951,N_21891);
and U22023 (N_22023,N_21974,N_21983);
xor U22024 (N_22024,N_21918,N_21825);
or U22025 (N_22025,N_21816,N_21876);
nor U22026 (N_22026,N_21863,N_21985);
xnor U22027 (N_22027,N_21953,N_21949);
or U22028 (N_22028,N_21855,N_21847);
or U22029 (N_22029,N_21803,N_21989);
xor U22030 (N_22030,N_21987,N_21909);
nand U22031 (N_22031,N_21954,N_21854);
and U22032 (N_22032,N_21972,N_21882);
or U22033 (N_22033,N_21818,N_21879);
and U22034 (N_22034,N_21968,N_21975);
or U22035 (N_22035,N_21996,N_21965);
xor U22036 (N_22036,N_21889,N_21920);
nand U22037 (N_22037,N_21842,N_21821);
xnor U22038 (N_22038,N_21804,N_21981);
or U22039 (N_22039,N_21900,N_21999);
nand U22040 (N_22040,N_21814,N_21927);
nor U22041 (N_22041,N_21905,N_21886);
or U22042 (N_22042,N_21901,N_21837);
nand U22043 (N_22043,N_21919,N_21826);
nand U22044 (N_22044,N_21894,N_21843);
and U22045 (N_22045,N_21890,N_21823);
nor U22046 (N_22046,N_21850,N_21973);
or U22047 (N_22047,N_21896,N_21995);
nor U22048 (N_22048,N_21898,N_21802);
xnor U22049 (N_22049,N_21827,N_21988);
nor U22050 (N_22050,N_21935,N_21810);
nor U22051 (N_22051,N_21959,N_21867);
xor U22052 (N_22052,N_21815,N_21970);
and U22053 (N_22053,N_21846,N_21943);
and U22054 (N_22054,N_21881,N_21915);
nor U22055 (N_22055,N_21952,N_21932);
xnor U22056 (N_22056,N_21836,N_21807);
xnor U22057 (N_22057,N_21895,N_21902);
nand U22058 (N_22058,N_21878,N_21872);
nor U22059 (N_22059,N_21934,N_21840);
nand U22060 (N_22060,N_21830,N_21851);
xor U22061 (N_22061,N_21831,N_21892);
xnor U22062 (N_22062,N_21936,N_21928);
or U22063 (N_22063,N_21904,N_21921);
nor U22064 (N_22064,N_21868,N_21926);
or U22065 (N_22065,N_21853,N_21962);
xnor U22066 (N_22066,N_21841,N_21925);
and U22067 (N_22067,N_21833,N_21946);
and U22068 (N_22068,N_21993,N_21839);
nand U22069 (N_22069,N_21859,N_21834);
nand U22070 (N_22070,N_21844,N_21888);
or U22071 (N_22071,N_21873,N_21950);
or U22072 (N_22072,N_21967,N_21994);
xnor U22073 (N_22073,N_21862,N_21808);
xnor U22074 (N_22074,N_21838,N_21990);
or U22075 (N_22075,N_21805,N_21912);
nor U22076 (N_22076,N_21806,N_21986);
xnor U22077 (N_22077,N_21884,N_21991);
or U22078 (N_22078,N_21942,N_21832);
or U22079 (N_22079,N_21857,N_21923);
or U22080 (N_22080,N_21908,N_21948);
xor U22081 (N_22081,N_21856,N_21931);
nand U22082 (N_22082,N_21906,N_21865);
nor U22083 (N_22083,N_21957,N_21907);
xnor U22084 (N_22084,N_21956,N_21969);
and U22085 (N_22085,N_21852,N_21960);
and U22086 (N_22086,N_21940,N_21944);
xnor U22087 (N_22087,N_21887,N_21910);
and U22088 (N_22088,N_21875,N_21982);
and U22089 (N_22089,N_21930,N_21979);
xor U22090 (N_22090,N_21963,N_21861);
and U22091 (N_22091,N_21947,N_21835);
and U22092 (N_22092,N_21980,N_21809);
xnor U22093 (N_22093,N_21939,N_21899);
xor U22094 (N_22094,N_21961,N_21911);
or U22095 (N_22095,N_21922,N_21929);
nand U22096 (N_22096,N_21945,N_21992);
or U22097 (N_22097,N_21984,N_21860);
and U22098 (N_22098,N_21964,N_21976);
or U22099 (N_22099,N_21955,N_21883);
xnor U22100 (N_22100,N_21820,N_21912);
nand U22101 (N_22101,N_21892,N_21918);
xor U22102 (N_22102,N_21925,N_21825);
or U22103 (N_22103,N_21864,N_21854);
nand U22104 (N_22104,N_21832,N_21982);
and U22105 (N_22105,N_21827,N_21932);
nor U22106 (N_22106,N_21854,N_21873);
or U22107 (N_22107,N_21948,N_21953);
nor U22108 (N_22108,N_21895,N_21865);
nand U22109 (N_22109,N_21986,N_21858);
and U22110 (N_22110,N_21892,N_21881);
xor U22111 (N_22111,N_21953,N_21988);
nor U22112 (N_22112,N_21823,N_21901);
nor U22113 (N_22113,N_21864,N_21814);
xnor U22114 (N_22114,N_21991,N_21942);
nor U22115 (N_22115,N_21904,N_21960);
and U22116 (N_22116,N_21937,N_21989);
xnor U22117 (N_22117,N_21956,N_21971);
nand U22118 (N_22118,N_21923,N_21969);
or U22119 (N_22119,N_21922,N_21906);
and U22120 (N_22120,N_21964,N_21877);
and U22121 (N_22121,N_21905,N_21865);
and U22122 (N_22122,N_21929,N_21837);
nor U22123 (N_22123,N_21915,N_21802);
nor U22124 (N_22124,N_21972,N_21937);
or U22125 (N_22125,N_21889,N_21840);
nand U22126 (N_22126,N_21840,N_21850);
xor U22127 (N_22127,N_21915,N_21960);
xor U22128 (N_22128,N_21802,N_21998);
and U22129 (N_22129,N_21840,N_21919);
xnor U22130 (N_22130,N_21878,N_21882);
nand U22131 (N_22131,N_21885,N_21956);
nor U22132 (N_22132,N_21946,N_21811);
nor U22133 (N_22133,N_21855,N_21938);
xor U22134 (N_22134,N_21928,N_21943);
or U22135 (N_22135,N_21975,N_21872);
nand U22136 (N_22136,N_21943,N_21948);
nor U22137 (N_22137,N_21927,N_21874);
xnor U22138 (N_22138,N_21843,N_21974);
xor U22139 (N_22139,N_21965,N_21878);
nand U22140 (N_22140,N_21993,N_21887);
nand U22141 (N_22141,N_21827,N_21976);
xnor U22142 (N_22142,N_21842,N_21982);
xor U22143 (N_22143,N_21968,N_21948);
or U22144 (N_22144,N_21804,N_21932);
and U22145 (N_22145,N_21910,N_21903);
nor U22146 (N_22146,N_21833,N_21878);
nand U22147 (N_22147,N_21911,N_21992);
or U22148 (N_22148,N_21947,N_21920);
and U22149 (N_22149,N_21828,N_21875);
and U22150 (N_22150,N_21805,N_21911);
nor U22151 (N_22151,N_21869,N_21902);
nand U22152 (N_22152,N_21974,N_21894);
and U22153 (N_22153,N_21933,N_21932);
and U22154 (N_22154,N_21964,N_21899);
and U22155 (N_22155,N_21924,N_21905);
nand U22156 (N_22156,N_21931,N_21863);
xnor U22157 (N_22157,N_21954,N_21911);
xor U22158 (N_22158,N_21851,N_21825);
xor U22159 (N_22159,N_21822,N_21911);
and U22160 (N_22160,N_21857,N_21882);
and U22161 (N_22161,N_21930,N_21894);
nor U22162 (N_22162,N_21845,N_21980);
and U22163 (N_22163,N_21994,N_21983);
xor U22164 (N_22164,N_21966,N_21927);
or U22165 (N_22165,N_21901,N_21922);
nand U22166 (N_22166,N_21982,N_21928);
nor U22167 (N_22167,N_21998,N_21931);
or U22168 (N_22168,N_21883,N_21961);
nand U22169 (N_22169,N_21931,N_21968);
nor U22170 (N_22170,N_21833,N_21970);
and U22171 (N_22171,N_21886,N_21953);
and U22172 (N_22172,N_21966,N_21916);
nor U22173 (N_22173,N_21862,N_21968);
nor U22174 (N_22174,N_21941,N_21813);
and U22175 (N_22175,N_21827,N_21805);
nand U22176 (N_22176,N_21970,N_21879);
xor U22177 (N_22177,N_21848,N_21841);
xor U22178 (N_22178,N_21894,N_21925);
nand U22179 (N_22179,N_21847,N_21858);
nand U22180 (N_22180,N_21820,N_21839);
or U22181 (N_22181,N_21871,N_21909);
or U22182 (N_22182,N_21938,N_21871);
or U22183 (N_22183,N_21806,N_21840);
nor U22184 (N_22184,N_21858,N_21963);
nand U22185 (N_22185,N_21827,N_21815);
or U22186 (N_22186,N_21904,N_21835);
and U22187 (N_22187,N_21851,N_21972);
or U22188 (N_22188,N_21890,N_21990);
or U22189 (N_22189,N_21899,N_21929);
nor U22190 (N_22190,N_21975,N_21842);
nor U22191 (N_22191,N_21930,N_21884);
nor U22192 (N_22192,N_21920,N_21956);
nor U22193 (N_22193,N_21941,N_21895);
nand U22194 (N_22194,N_21995,N_21898);
xor U22195 (N_22195,N_21977,N_21928);
xor U22196 (N_22196,N_21957,N_21926);
or U22197 (N_22197,N_21904,N_21913);
xor U22198 (N_22198,N_21891,N_21968);
xnor U22199 (N_22199,N_21867,N_21891);
xnor U22200 (N_22200,N_22022,N_22026);
xor U22201 (N_22201,N_22085,N_22060);
xnor U22202 (N_22202,N_22043,N_22028);
xor U22203 (N_22203,N_22053,N_22164);
or U22204 (N_22204,N_22143,N_22184);
xnor U22205 (N_22205,N_22191,N_22127);
nand U22206 (N_22206,N_22044,N_22054);
xnor U22207 (N_22207,N_22001,N_22166);
nand U22208 (N_22208,N_22175,N_22118);
xnor U22209 (N_22209,N_22177,N_22180);
nand U22210 (N_22210,N_22093,N_22038);
nor U22211 (N_22211,N_22120,N_22129);
and U22212 (N_22212,N_22097,N_22159);
and U22213 (N_22213,N_22122,N_22140);
and U22214 (N_22214,N_22141,N_22040);
nor U22215 (N_22215,N_22010,N_22183);
nand U22216 (N_22216,N_22113,N_22006);
or U22217 (N_22217,N_22000,N_22107);
nand U22218 (N_22218,N_22059,N_22124);
nand U22219 (N_22219,N_22103,N_22119);
xor U22220 (N_22220,N_22158,N_22055);
xnor U22221 (N_22221,N_22019,N_22156);
nor U22222 (N_22222,N_22037,N_22098);
nand U22223 (N_22223,N_22002,N_22075);
nand U22224 (N_22224,N_22015,N_22092);
nor U22225 (N_22225,N_22137,N_22090);
nand U22226 (N_22226,N_22178,N_22012);
nand U22227 (N_22227,N_22193,N_22115);
nand U22228 (N_22228,N_22069,N_22186);
nor U22229 (N_22229,N_22146,N_22018);
xnor U22230 (N_22230,N_22007,N_22050);
xnor U22231 (N_22231,N_22168,N_22039);
and U22232 (N_22232,N_22065,N_22128);
or U22233 (N_22233,N_22162,N_22154);
nor U22234 (N_22234,N_22041,N_22181);
xnor U22235 (N_22235,N_22135,N_22017);
nand U22236 (N_22236,N_22105,N_22032);
and U22237 (N_22237,N_22187,N_22068);
nand U22238 (N_22238,N_22117,N_22024);
xor U22239 (N_22239,N_22096,N_22099);
or U22240 (N_22240,N_22149,N_22023);
and U22241 (N_22241,N_22042,N_22004);
and U22242 (N_22242,N_22131,N_22188);
xor U22243 (N_22243,N_22031,N_22080);
nor U22244 (N_22244,N_22161,N_22163);
or U22245 (N_22245,N_22153,N_22104);
or U22246 (N_22246,N_22192,N_22013);
or U22247 (N_22247,N_22155,N_22025);
or U22248 (N_22248,N_22081,N_22114);
xor U22249 (N_22249,N_22151,N_22130);
and U22250 (N_22250,N_22198,N_22126);
or U22251 (N_22251,N_22150,N_22056);
xnor U22252 (N_22252,N_22199,N_22035);
or U22253 (N_22253,N_22109,N_22094);
nand U22254 (N_22254,N_22182,N_22144);
and U22255 (N_22255,N_22195,N_22136);
xor U22256 (N_22256,N_22070,N_22157);
xnor U22257 (N_22257,N_22049,N_22116);
xnor U22258 (N_22258,N_22170,N_22171);
or U22259 (N_22259,N_22167,N_22045);
nand U22260 (N_22260,N_22106,N_22078);
and U22261 (N_22261,N_22048,N_22008);
nor U22262 (N_22262,N_22088,N_22142);
or U22263 (N_22263,N_22021,N_22033);
or U22264 (N_22264,N_22016,N_22179);
or U22265 (N_22265,N_22086,N_22034);
nand U22266 (N_22266,N_22084,N_22087);
nor U22267 (N_22267,N_22100,N_22046);
or U22268 (N_22268,N_22169,N_22112);
nand U22269 (N_22269,N_22064,N_22132);
nand U22270 (N_22270,N_22091,N_22139);
nand U22271 (N_22271,N_22147,N_22196);
or U22272 (N_22272,N_22089,N_22145);
xnor U22273 (N_22273,N_22047,N_22102);
nand U22274 (N_22274,N_22072,N_22011);
nand U22275 (N_22275,N_22071,N_22082);
xor U22276 (N_22276,N_22036,N_22101);
or U22277 (N_22277,N_22062,N_22189);
nor U22278 (N_22278,N_22076,N_22051);
or U22279 (N_22279,N_22067,N_22174);
or U22280 (N_22280,N_22014,N_22003);
nand U22281 (N_22281,N_22125,N_22027);
or U22282 (N_22282,N_22197,N_22172);
nor U22283 (N_22283,N_22185,N_22160);
nor U22284 (N_22284,N_22110,N_22121);
nand U22285 (N_22285,N_22074,N_22029);
nor U22286 (N_22286,N_22057,N_22176);
nor U22287 (N_22287,N_22194,N_22061);
nand U22288 (N_22288,N_22066,N_22030);
and U22289 (N_22289,N_22173,N_22152);
or U22290 (N_22290,N_22058,N_22095);
and U22291 (N_22291,N_22083,N_22165);
and U22292 (N_22292,N_22077,N_22133);
or U22293 (N_22293,N_22190,N_22123);
nand U22294 (N_22294,N_22148,N_22108);
and U22295 (N_22295,N_22138,N_22020);
nor U22296 (N_22296,N_22005,N_22063);
and U22297 (N_22297,N_22009,N_22079);
nor U22298 (N_22298,N_22111,N_22073);
and U22299 (N_22299,N_22052,N_22134);
xor U22300 (N_22300,N_22073,N_22148);
nand U22301 (N_22301,N_22078,N_22065);
nand U22302 (N_22302,N_22094,N_22104);
nand U22303 (N_22303,N_22163,N_22053);
and U22304 (N_22304,N_22057,N_22195);
and U22305 (N_22305,N_22188,N_22003);
nand U22306 (N_22306,N_22091,N_22145);
nor U22307 (N_22307,N_22157,N_22074);
xnor U22308 (N_22308,N_22138,N_22121);
and U22309 (N_22309,N_22112,N_22158);
xnor U22310 (N_22310,N_22036,N_22144);
or U22311 (N_22311,N_22199,N_22043);
or U22312 (N_22312,N_22064,N_22092);
and U22313 (N_22313,N_22166,N_22109);
and U22314 (N_22314,N_22127,N_22051);
nand U22315 (N_22315,N_22132,N_22176);
nor U22316 (N_22316,N_22185,N_22001);
or U22317 (N_22317,N_22097,N_22028);
nand U22318 (N_22318,N_22127,N_22118);
and U22319 (N_22319,N_22123,N_22058);
nor U22320 (N_22320,N_22165,N_22131);
or U22321 (N_22321,N_22009,N_22163);
nand U22322 (N_22322,N_22027,N_22189);
xor U22323 (N_22323,N_22130,N_22067);
xnor U22324 (N_22324,N_22043,N_22101);
nand U22325 (N_22325,N_22097,N_22105);
xor U22326 (N_22326,N_22044,N_22007);
nand U22327 (N_22327,N_22163,N_22007);
and U22328 (N_22328,N_22118,N_22149);
nand U22329 (N_22329,N_22134,N_22054);
nand U22330 (N_22330,N_22046,N_22112);
and U22331 (N_22331,N_22033,N_22196);
nand U22332 (N_22332,N_22118,N_22110);
or U22333 (N_22333,N_22054,N_22052);
and U22334 (N_22334,N_22007,N_22000);
nand U22335 (N_22335,N_22121,N_22008);
nor U22336 (N_22336,N_22117,N_22059);
nand U22337 (N_22337,N_22097,N_22158);
nor U22338 (N_22338,N_22162,N_22034);
or U22339 (N_22339,N_22135,N_22167);
or U22340 (N_22340,N_22101,N_22114);
nand U22341 (N_22341,N_22111,N_22159);
nor U22342 (N_22342,N_22091,N_22198);
nand U22343 (N_22343,N_22097,N_22162);
nor U22344 (N_22344,N_22001,N_22188);
nor U22345 (N_22345,N_22026,N_22068);
or U22346 (N_22346,N_22015,N_22137);
nor U22347 (N_22347,N_22109,N_22131);
or U22348 (N_22348,N_22024,N_22190);
or U22349 (N_22349,N_22018,N_22038);
xor U22350 (N_22350,N_22119,N_22034);
or U22351 (N_22351,N_22052,N_22132);
and U22352 (N_22352,N_22012,N_22163);
nor U22353 (N_22353,N_22162,N_22174);
and U22354 (N_22354,N_22187,N_22067);
xnor U22355 (N_22355,N_22173,N_22066);
xnor U22356 (N_22356,N_22161,N_22009);
xnor U22357 (N_22357,N_22010,N_22171);
nor U22358 (N_22358,N_22136,N_22014);
and U22359 (N_22359,N_22124,N_22136);
and U22360 (N_22360,N_22196,N_22093);
and U22361 (N_22361,N_22177,N_22035);
nor U22362 (N_22362,N_22146,N_22166);
or U22363 (N_22363,N_22034,N_22025);
nor U22364 (N_22364,N_22089,N_22136);
nor U22365 (N_22365,N_22045,N_22180);
or U22366 (N_22366,N_22073,N_22048);
nand U22367 (N_22367,N_22022,N_22100);
or U22368 (N_22368,N_22007,N_22061);
xnor U22369 (N_22369,N_22171,N_22179);
nor U22370 (N_22370,N_22156,N_22186);
nor U22371 (N_22371,N_22002,N_22069);
or U22372 (N_22372,N_22089,N_22014);
nor U22373 (N_22373,N_22077,N_22177);
xnor U22374 (N_22374,N_22167,N_22095);
xnor U22375 (N_22375,N_22163,N_22041);
or U22376 (N_22376,N_22130,N_22072);
and U22377 (N_22377,N_22100,N_22089);
and U22378 (N_22378,N_22109,N_22198);
nand U22379 (N_22379,N_22084,N_22082);
nor U22380 (N_22380,N_22024,N_22139);
or U22381 (N_22381,N_22153,N_22036);
nor U22382 (N_22382,N_22110,N_22101);
xnor U22383 (N_22383,N_22099,N_22086);
nand U22384 (N_22384,N_22013,N_22196);
xnor U22385 (N_22385,N_22087,N_22099);
nor U22386 (N_22386,N_22199,N_22026);
or U22387 (N_22387,N_22092,N_22160);
or U22388 (N_22388,N_22178,N_22170);
and U22389 (N_22389,N_22031,N_22022);
xnor U22390 (N_22390,N_22016,N_22121);
nand U22391 (N_22391,N_22031,N_22021);
and U22392 (N_22392,N_22117,N_22152);
xor U22393 (N_22393,N_22146,N_22028);
nand U22394 (N_22394,N_22026,N_22081);
nand U22395 (N_22395,N_22039,N_22182);
or U22396 (N_22396,N_22133,N_22116);
nand U22397 (N_22397,N_22039,N_22161);
and U22398 (N_22398,N_22009,N_22015);
nor U22399 (N_22399,N_22057,N_22032);
or U22400 (N_22400,N_22254,N_22245);
nor U22401 (N_22401,N_22299,N_22339);
and U22402 (N_22402,N_22267,N_22382);
nor U22403 (N_22403,N_22266,N_22209);
nor U22404 (N_22404,N_22268,N_22309);
or U22405 (N_22405,N_22256,N_22274);
and U22406 (N_22406,N_22287,N_22272);
and U22407 (N_22407,N_22248,N_22333);
or U22408 (N_22408,N_22255,N_22228);
or U22409 (N_22409,N_22352,N_22354);
nand U22410 (N_22410,N_22356,N_22235);
or U22411 (N_22411,N_22211,N_22342);
or U22412 (N_22412,N_22362,N_22317);
or U22413 (N_22413,N_22384,N_22286);
xnor U22414 (N_22414,N_22224,N_22264);
nor U22415 (N_22415,N_22258,N_22281);
xor U22416 (N_22416,N_22217,N_22334);
nor U22417 (N_22417,N_22238,N_22388);
xnor U22418 (N_22418,N_22251,N_22395);
and U22419 (N_22419,N_22216,N_22207);
xnor U22420 (N_22420,N_22364,N_22358);
nor U22421 (N_22421,N_22225,N_22372);
and U22422 (N_22422,N_22381,N_22365);
nor U22423 (N_22423,N_22316,N_22212);
xnor U22424 (N_22424,N_22366,N_22293);
xor U22425 (N_22425,N_22392,N_22232);
xor U22426 (N_22426,N_22233,N_22234);
nand U22427 (N_22427,N_22368,N_22208);
and U22428 (N_22428,N_22304,N_22307);
and U22429 (N_22429,N_22306,N_22222);
xor U22430 (N_22430,N_22283,N_22303);
and U22431 (N_22431,N_22341,N_22376);
nand U22432 (N_22432,N_22231,N_22244);
or U22433 (N_22433,N_22318,N_22284);
nand U22434 (N_22434,N_22340,N_22262);
or U22435 (N_22435,N_22300,N_22326);
nor U22436 (N_22436,N_22355,N_22247);
nor U22437 (N_22437,N_22383,N_22369);
and U22438 (N_22438,N_22329,N_22302);
and U22439 (N_22439,N_22374,N_22230);
nand U22440 (N_22440,N_22218,N_22292);
xnor U22441 (N_22441,N_22312,N_22350);
nand U22442 (N_22442,N_22393,N_22335);
and U22443 (N_22443,N_22296,N_22347);
xor U22444 (N_22444,N_22398,N_22305);
xor U22445 (N_22445,N_22219,N_22246);
and U22446 (N_22446,N_22371,N_22270);
and U22447 (N_22447,N_22315,N_22394);
nand U22448 (N_22448,N_22322,N_22277);
nor U22449 (N_22449,N_22203,N_22377);
or U22450 (N_22450,N_22269,N_22205);
or U22451 (N_22451,N_22204,N_22390);
and U22452 (N_22452,N_22370,N_22263);
nand U22453 (N_22453,N_22385,N_22226);
nand U22454 (N_22454,N_22288,N_22221);
nand U22455 (N_22455,N_22261,N_22353);
xnor U22456 (N_22456,N_22386,N_22397);
and U22457 (N_22457,N_22301,N_22249);
xor U22458 (N_22458,N_22239,N_22375);
nor U22459 (N_22459,N_22319,N_22260);
or U22460 (N_22460,N_22242,N_22379);
xor U22461 (N_22461,N_22321,N_22399);
and U22462 (N_22462,N_22273,N_22215);
xor U22463 (N_22463,N_22210,N_22298);
or U22464 (N_22464,N_22285,N_22373);
nor U22465 (N_22465,N_22324,N_22250);
or U22466 (N_22466,N_22240,N_22332);
xor U22467 (N_22467,N_22200,N_22265);
nor U22468 (N_22468,N_22378,N_22201);
xor U22469 (N_22469,N_22311,N_22336);
or U22470 (N_22470,N_22280,N_22348);
and U22471 (N_22471,N_22325,N_22361);
and U22472 (N_22472,N_22236,N_22331);
nand U22473 (N_22473,N_22396,N_22271);
nor U22474 (N_22474,N_22295,N_22360);
xor U22475 (N_22475,N_22227,N_22253);
or U22476 (N_22476,N_22351,N_22343);
xor U22477 (N_22477,N_22387,N_22367);
or U22478 (N_22478,N_22357,N_22363);
nor U22479 (N_22479,N_22206,N_22289);
nand U22480 (N_22480,N_22297,N_22391);
or U22481 (N_22481,N_22323,N_22241);
xor U22482 (N_22482,N_22337,N_22243);
nand U22483 (N_22483,N_22327,N_22346);
nor U22484 (N_22484,N_22294,N_22237);
xor U22485 (N_22485,N_22223,N_22338);
or U22486 (N_22486,N_22314,N_22252);
and U22487 (N_22487,N_22313,N_22220);
and U22488 (N_22488,N_22330,N_22275);
nor U22489 (N_22489,N_22282,N_22290);
nand U22490 (N_22490,N_22380,N_22279);
or U22491 (N_22491,N_22349,N_22276);
and U22492 (N_22492,N_22257,N_22359);
nor U22493 (N_22493,N_22310,N_22259);
xor U22494 (N_22494,N_22229,N_22213);
nor U22495 (N_22495,N_22308,N_22345);
or U22496 (N_22496,N_22328,N_22320);
nor U22497 (N_22497,N_22214,N_22291);
xnor U22498 (N_22498,N_22202,N_22278);
or U22499 (N_22499,N_22389,N_22344);
and U22500 (N_22500,N_22389,N_22223);
and U22501 (N_22501,N_22216,N_22236);
xor U22502 (N_22502,N_22282,N_22353);
and U22503 (N_22503,N_22349,N_22298);
nand U22504 (N_22504,N_22341,N_22312);
nor U22505 (N_22505,N_22392,N_22279);
and U22506 (N_22506,N_22349,N_22346);
or U22507 (N_22507,N_22301,N_22368);
nor U22508 (N_22508,N_22333,N_22323);
and U22509 (N_22509,N_22290,N_22316);
nand U22510 (N_22510,N_22214,N_22206);
or U22511 (N_22511,N_22256,N_22292);
and U22512 (N_22512,N_22377,N_22222);
nor U22513 (N_22513,N_22231,N_22364);
and U22514 (N_22514,N_22369,N_22203);
nor U22515 (N_22515,N_22269,N_22211);
nor U22516 (N_22516,N_22325,N_22370);
xor U22517 (N_22517,N_22219,N_22334);
or U22518 (N_22518,N_22213,N_22396);
nor U22519 (N_22519,N_22255,N_22220);
nor U22520 (N_22520,N_22315,N_22200);
or U22521 (N_22521,N_22213,N_22375);
or U22522 (N_22522,N_22343,N_22303);
or U22523 (N_22523,N_22368,N_22337);
or U22524 (N_22524,N_22213,N_22272);
and U22525 (N_22525,N_22330,N_22367);
nand U22526 (N_22526,N_22314,N_22328);
or U22527 (N_22527,N_22347,N_22336);
nand U22528 (N_22528,N_22325,N_22288);
or U22529 (N_22529,N_22293,N_22308);
or U22530 (N_22530,N_22332,N_22294);
nand U22531 (N_22531,N_22211,N_22227);
nor U22532 (N_22532,N_22234,N_22297);
nor U22533 (N_22533,N_22323,N_22399);
xor U22534 (N_22534,N_22208,N_22274);
and U22535 (N_22535,N_22340,N_22213);
nor U22536 (N_22536,N_22245,N_22318);
and U22537 (N_22537,N_22344,N_22353);
or U22538 (N_22538,N_22313,N_22238);
nand U22539 (N_22539,N_22301,N_22330);
xnor U22540 (N_22540,N_22360,N_22272);
or U22541 (N_22541,N_22310,N_22336);
nand U22542 (N_22542,N_22376,N_22329);
nand U22543 (N_22543,N_22264,N_22371);
or U22544 (N_22544,N_22376,N_22215);
nand U22545 (N_22545,N_22345,N_22306);
and U22546 (N_22546,N_22260,N_22357);
nor U22547 (N_22547,N_22319,N_22217);
nor U22548 (N_22548,N_22386,N_22395);
or U22549 (N_22549,N_22347,N_22235);
xor U22550 (N_22550,N_22229,N_22309);
nor U22551 (N_22551,N_22236,N_22374);
or U22552 (N_22552,N_22316,N_22381);
nand U22553 (N_22553,N_22323,N_22226);
and U22554 (N_22554,N_22265,N_22266);
nand U22555 (N_22555,N_22268,N_22277);
nor U22556 (N_22556,N_22387,N_22283);
nor U22557 (N_22557,N_22313,N_22273);
or U22558 (N_22558,N_22243,N_22253);
and U22559 (N_22559,N_22397,N_22318);
or U22560 (N_22560,N_22390,N_22354);
and U22561 (N_22561,N_22249,N_22201);
nand U22562 (N_22562,N_22254,N_22359);
nor U22563 (N_22563,N_22393,N_22392);
and U22564 (N_22564,N_22284,N_22221);
xor U22565 (N_22565,N_22219,N_22240);
nor U22566 (N_22566,N_22335,N_22214);
or U22567 (N_22567,N_22244,N_22294);
nor U22568 (N_22568,N_22333,N_22344);
nor U22569 (N_22569,N_22229,N_22204);
xor U22570 (N_22570,N_22304,N_22343);
nor U22571 (N_22571,N_22374,N_22210);
xor U22572 (N_22572,N_22308,N_22281);
xor U22573 (N_22573,N_22306,N_22280);
xnor U22574 (N_22574,N_22330,N_22226);
and U22575 (N_22575,N_22334,N_22303);
nor U22576 (N_22576,N_22238,N_22354);
nand U22577 (N_22577,N_22391,N_22260);
nor U22578 (N_22578,N_22230,N_22255);
nand U22579 (N_22579,N_22327,N_22383);
xor U22580 (N_22580,N_22228,N_22302);
or U22581 (N_22581,N_22382,N_22209);
nand U22582 (N_22582,N_22386,N_22273);
or U22583 (N_22583,N_22275,N_22321);
or U22584 (N_22584,N_22383,N_22227);
and U22585 (N_22585,N_22357,N_22246);
nor U22586 (N_22586,N_22285,N_22250);
nand U22587 (N_22587,N_22283,N_22276);
or U22588 (N_22588,N_22387,N_22275);
and U22589 (N_22589,N_22219,N_22352);
nor U22590 (N_22590,N_22391,N_22386);
and U22591 (N_22591,N_22337,N_22205);
or U22592 (N_22592,N_22222,N_22389);
nand U22593 (N_22593,N_22233,N_22339);
or U22594 (N_22594,N_22220,N_22224);
xnor U22595 (N_22595,N_22239,N_22271);
nor U22596 (N_22596,N_22318,N_22206);
xor U22597 (N_22597,N_22265,N_22254);
nor U22598 (N_22598,N_22230,N_22205);
and U22599 (N_22599,N_22233,N_22348);
nor U22600 (N_22600,N_22469,N_22506);
xor U22601 (N_22601,N_22455,N_22486);
nand U22602 (N_22602,N_22449,N_22546);
and U22603 (N_22603,N_22560,N_22419);
nor U22604 (N_22604,N_22588,N_22575);
nand U22605 (N_22605,N_22597,N_22513);
xnor U22606 (N_22606,N_22539,N_22565);
nand U22607 (N_22607,N_22443,N_22529);
or U22608 (N_22608,N_22428,N_22500);
nand U22609 (N_22609,N_22467,N_22499);
and U22610 (N_22610,N_22498,N_22453);
and U22611 (N_22611,N_22519,N_22490);
nand U22612 (N_22612,N_22482,N_22562);
xnor U22613 (N_22613,N_22445,N_22439);
xor U22614 (N_22614,N_22440,N_22491);
or U22615 (N_22615,N_22466,N_22454);
or U22616 (N_22616,N_22582,N_22502);
nand U22617 (N_22617,N_22462,N_22592);
or U22618 (N_22618,N_22432,N_22464);
nand U22619 (N_22619,N_22510,N_22563);
nor U22620 (N_22620,N_22417,N_22504);
and U22621 (N_22621,N_22574,N_22535);
nor U22622 (N_22622,N_22508,N_22568);
nand U22623 (N_22623,N_22576,N_22438);
nor U22624 (N_22624,N_22450,N_22558);
xor U22625 (N_22625,N_22473,N_22525);
and U22626 (N_22626,N_22475,N_22401);
or U22627 (N_22627,N_22514,N_22404);
xnor U22628 (N_22628,N_22516,N_22520);
xor U22629 (N_22629,N_22433,N_22412);
xor U22630 (N_22630,N_22522,N_22460);
nand U22631 (N_22631,N_22489,N_22556);
or U22632 (N_22632,N_22583,N_22465);
nand U22633 (N_22633,N_22590,N_22481);
and U22634 (N_22634,N_22434,N_22418);
or U22635 (N_22635,N_22420,N_22495);
and U22636 (N_22636,N_22400,N_22569);
and U22637 (N_22637,N_22541,N_22451);
nand U22638 (N_22638,N_22446,N_22487);
nor U22639 (N_22639,N_22543,N_22414);
or U22640 (N_22640,N_22551,N_22552);
and U22641 (N_22641,N_22571,N_22470);
nand U22642 (N_22642,N_22554,N_22409);
and U22643 (N_22643,N_22485,N_22458);
and U22644 (N_22644,N_22483,N_22599);
xor U22645 (N_22645,N_22530,N_22488);
or U22646 (N_22646,N_22403,N_22457);
or U22647 (N_22647,N_22584,N_22477);
and U22648 (N_22648,N_22544,N_22447);
or U22649 (N_22649,N_22427,N_22593);
or U22650 (N_22650,N_22468,N_22456);
nor U22651 (N_22651,N_22523,N_22426);
nand U22652 (N_22652,N_22577,N_22415);
nand U22653 (N_22653,N_22542,N_22559);
or U22654 (N_22654,N_22596,N_22547);
nor U22655 (N_22655,N_22461,N_22586);
and U22656 (N_22656,N_22578,N_22431);
or U22657 (N_22657,N_22598,N_22573);
xor U22658 (N_22658,N_22503,N_22509);
xor U22659 (N_22659,N_22416,N_22570);
or U22660 (N_22660,N_22476,N_22517);
or U22661 (N_22661,N_22531,N_22555);
or U22662 (N_22662,N_22527,N_22534);
and U22663 (N_22663,N_22526,N_22407);
nand U22664 (N_22664,N_22423,N_22474);
xnor U22665 (N_22665,N_22553,N_22507);
or U22666 (N_22666,N_22484,N_22540);
or U22667 (N_22667,N_22436,N_22532);
and U22668 (N_22668,N_22478,N_22448);
or U22669 (N_22669,N_22594,N_22581);
or U22670 (N_22670,N_22413,N_22545);
nand U22671 (N_22671,N_22494,N_22561);
nor U22672 (N_22672,N_22463,N_22567);
and U22673 (N_22673,N_22548,N_22472);
nand U22674 (N_22674,N_22579,N_22496);
xnor U22675 (N_22675,N_22505,N_22549);
or U22676 (N_22676,N_22444,N_22512);
xnor U22677 (N_22677,N_22480,N_22492);
nand U22678 (N_22678,N_22422,N_22585);
nand U22679 (N_22679,N_22429,N_22493);
nor U22680 (N_22680,N_22425,N_22437);
nand U22681 (N_22681,N_22538,N_22471);
or U22682 (N_22682,N_22564,N_22536);
and U22683 (N_22683,N_22528,N_22497);
or U22684 (N_22684,N_22591,N_22572);
and U22685 (N_22685,N_22430,N_22587);
nand U22686 (N_22686,N_22406,N_22557);
or U22687 (N_22687,N_22566,N_22442);
and U22688 (N_22688,N_22589,N_22518);
and U22689 (N_22689,N_22595,N_22511);
or U22690 (N_22690,N_22515,N_22452);
nor U22691 (N_22691,N_22521,N_22402);
nor U22692 (N_22692,N_22421,N_22424);
and U22693 (N_22693,N_22459,N_22550);
nand U22694 (N_22694,N_22501,N_22441);
nor U22695 (N_22695,N_22580,N_22435);
nor U22696 (N_22696,N_22411,N_22524);
nand U22697 (N_22697,N_22537,N_22479);
and U22698 (N_22698,N_22405,N_22410);
or U22699 (N_22699,N_22408,N_22533);
nor U22700 (N_22700,N_22575,N_22407);
or U22701 (N_22701,N_22488,N_22479);
xor U22702 (N_22702,N_22503,N_22476);
xnor U22703 (N_22703,N_22453,N_22468);
or U22704 (N_22704,N_22465,N_22512);
and U22705 (N_22705,N_22550,N_22492);
nand U22706 (N_22706,N_22483,N_22412);
nand U22707 (N_22707,N_22402,N_22575);
nor U22708 (N_22708,N_22469,N_22454);
or U22709 (N_22709,N_22504,N_22437);
or U22710 (N_22710,N_22583,N_22575);
nand U22711 (N_22711,N_22586,N_22525);
and U22712 (N_22712,N_22521,N_22536);
nor U22713 (N_22713,N_22465,N_22426);
or U22714 (N_22714,N_22495,N_22519);
xor U22715 (N_22715,N_22445,N_22466);
nor U22716 (N_22716,N_22490,N_22503);
xnor U22717 (N_22717,N_22469,N_22586);
or U22718 (N_22718,N_22479,N_22531);
and U22719 (N_22719,N_22404,N_22466);
nor U22720 (N_22720,N_22586,N_22414);
or U22721 (N_22721,N_22542,N_22525);
xnor U22722 (N_22722,N_22584,N_22577);
nand U22723 (N_22723,N_22528,N_22593);
and U22724 (N_22724,N_22486,N_22558);
or U22725 (N_22725,N_22550,N_22521);
or U22726 (N_22726,N_22415,N_22536);
nor U22727 (N_22727,N_22426,N_22418);
or U22728 (N_22728,N_22572,N_22584);
and U22729 (N_22729,N_22479,N_22553);
nand U22730 (N_22730,N_22517,N_22523);
or U22731 (N_22731,N_22556,N_22541);
nor U22732 (N_22732,N_22442,N_22554);
and U22733 (N_22733,N_22427,N_22569);
xnor U22734 (N_22734,N_22540,N_22411);
xnor U22735 (N_22735,N_22453,N_22542);
nor U22736 (N_22736,N_22575,N_22509);
or U22737 (N_22737,N_22413,N_22530);
nor U22738 (N_22738,N_22597,N_22441);
or U22739 (N_22739,N_22424,N_22439);
nor U22740 (N_22740,N_22591,N_22489);
xor U22741 (N_22741,N_22527,N_22535);
and U22742 (N_22742,N_22552,N_22595);
or U22743 (N_22743,N_22526,N_22554);
or U22744 (N_22744,N_22454,N_22440);
nor U22745 (N_22745,N_22471,N_22510);
nor U22746 (N_22746,N_22568,N_22572);
or U22747 (N_22747,N_22516,N_22413);
or U22748 (N_22748,N_22549,N_22496);
xor U22749 (N_22749,N_22583,N_22565);
nor U22750 (N_22750,N_22502,N_22549);
or U22751 (N_22751,N_22590,N_22591);
and U22752 (N_22752,N_22563,N_22501);
nand U22753 (N_22753,N_22546,N_22528);
nand U22754 (N_22754,N_22433,N_22527);
and U22755 (N_22755,N_22471,N_22485);
nor U22756 (N_22756,N_22404,N_22475);
nor U22757 (N_22757,N_22470,N_22440);
or U22758 (N_22758,N_22578,N_22566);
nand U22759 (N_22759,N_22585,N_22546);
nor U22760 (N_22760,N_22514,N_22599);
and U22761 (N_22761,N_22416,N_22453);
nand U22762 (N_22762,N_22578,N_22447);
xor U22763 (N_22763,N_22412,N_22444);
xor U22764 (N_22764,N_22449,N_22551);
or U22765 (N_22765,N_22524,N_22446);
or U22766 (N_22766,N_22461,N_22405);
or U22767 (N_22767,N_22531,N_22548);
nor U22768 (N_22768,N_22451,N_22521);
and U22769 (N_22769,N_22552,N_22560);
or U22770 (N_22770,N_22488,N_22425);
nand U22771 (N_22771,N_22583,N_22476);
xor U22772 (N_22772,N_22496,N_22516);
and U22773 (N_22773,N_22404,N_22566);
nor U22774 (N_22774,N_22418,N_22501);
and U22775 (N_22775,N_22468,N_22583);
nand U22776 (N_22776,N_22539,N_22410);
or U22777 (N_22777,N_22427,N_22567);
xnor U22778 (N_22778,N_22532,N_22477);
xnor U22779 (N_22779,N_22490,N_22516);
or U22780 (N_22780,N_22565,N_22509);
nand U22781 (N_22781,N_22480,N_22448);
nor U22782 (N_22782,N_22543,N_22457);
and U22783 (N_22783,N_22479,N_22534);
nand U22784 (N_22784,N_22496,N_22403);
and U22785 (N_22785,N_22447,N_22598);
xor U22786 (N_22786,N_22486,N_22529);
nor U22787 (N_22787,N_22424,N_22571);
xnor U22788 (N_22788,N_22560,N_22595);
xor U22789 (N_22789,N_22499,N_22585);
nand U22790 (N_22790,N_22406,N_22444);
or U22791 (N_22791,N_22486,N_22565);
nor U22792 (N_22792,N_22564,N_22493);
and U22793 (N_22793,N_22413,N_22430);
and U22794 (N_22794,N_22483,N_22493);
or U22795 (N_22795,N_22468,N_22544);
nor U22796 (N_22796,N_22587,N_22573);
and U22797 (N_22797,N_22507,N_22467);
xnor U22798 (N_22798,N_22555,N_22547);
nor U22799 (N_22799,N_22476,N_22464);
nor U22800 (N_22800,N_22642,N_22686);
xor U22801 (N_22801,N_22794,N_22661);
nand U22802 (N_22802,N_22692,N_22679);
xnor U22803 (N_22803,N_22699,N_22775);
nor U22804 (N_22804,N_22729,N_22685);
and U22805 (N_22805,N_22782,N_22610);
and U22806 (N_22806,N_22749,N_22655);
or U22807 (N_22807,N_22615,N_22601);
nor U22808 (N_22808,N_22694,N_22622);
xor U22809 (N_22809,N_22653,N_22788);
and U22810 (N_22810,N_22616,N_22764);
and U22811 (N_22811,N_22735,N_22602);
xnor U22812 (N_22812,N_22753,N_22627);
or U22813 (N_22813,N_22693,N_22639);
or U22814 (N_22814,N_22776,N_22718);
or U22815 (N_22815,N_22633,N_22746);
and U22816 (N_22816,N_22760,N_22673);
nand U22817 (N_22817,N_22695,N_22668);
nand U22818 (N_22818,N_22757,N_22798);
nor U22819 (N_22819,N_22779,N_22637);
nand U22820 (N_22820,N_22607,N_22751);
xnor U22821 (N_22821,N_22644,N_22707);
xnor U22822 (N_22822,N_22783,N_22606);
and U22823 (N_22823,N_22657,N_22613);
nand U22824 (N_22824,N_22645,N_22726);
nor U22825 (N_22825,N_22747,N_22678);
nand U22826 (N_22826,N_22682,N_22715);
and U22827 (N_22827,N_22756,N_22629);
and U22828 (N_22828,N_22758,N_22600);
and U22829 (N_22829,N_22612,N_22636);
or U22830 (N_22830,N_22786,N_22667);
nand U22831 (N_22831,N_22730,N_22769);
nor U22832 (N_22832,N_22632,N_22618);
xor U22833 (N_22833,N_22706,N_22752);
nand U22834 (N_22834,N_22720,N_22641);
or U22835 (N_22835,N_22683,N_22670);
nand U22836 (N_22836,N_22654,N_22680);
nor U22837 (N_22837,N_22659,N_22689);
and U22838 (N_22838,N_22789,N_22743);
or U22839 (N_22839,N_22643,N_22732);
nor U22840 (N_22840,N_22701,N_22611);
xor U22841 (N_22841,N_22647,N_22792);
nor U22842 (N_22842,N_22620,N_22698);
xnor U22843 (N_22843,N_22778,N_22733);
nand U22844 (N_22844,N_22684,N_22703);
and U22845 (N_22845,N_22740,N_22625);
and U22846 (N_22846,N_22717,N_22750);
xor U22847 (N_22847,N_22772,N_22754);
or U22848 (N_22848,N_22777,N_22731);
nor U22849 (N_22849,N_22796,N_22608);
nor U22850 (N_22850,N_22635,N_22799);
nand U22851 (N_22851,N_22716,N_22650);
and U22852 (N_22852,N_22674,N_22797);
xor U22853 (N_22853,N_22711,N_22604);
nor U22854 (N_22854,N_22744,N_22704);
and U22855 (N_22855,N_22614,N_22666);
nand U22856 (N_22856,N_22742,N_22761);
and U22857 (N_22857,N_22675,N_22708);
nor U22858 (N_22858,N_22739,N_22765);
nor U22859 (N_22859,N_22759,N_22624);
nor U22860 (N_22860,N_22710,N_22738);
xnor U22861 (N_22861,N_22734,N_22790);
nor U22862 (N_22862,N_22631,N_22623);
and U22863 (N_22863,N_22619,N_22605);
or U22864 (N_22864,N_22669,N_22793);
nand U22865 (N_22865,N_22724,N_22691);
nor U22866 (N_22866,N_22660,N_22630);
nor U22867 (N_22867,N_22714,N_22648);
nor U22868 (N_22868,N_22727,N_22651);
xor U22869 (N_22869,N_22728,N_22787);
xor U22870 (N_22870,N_22664,N_22649);
nor U22871 (N_22871,N_22713,N_22736);
nand U22872 (N_22872,N_22662,N_22652);
or U22873 (N_22873,N_22656,N_22681);
or U22874 (N_22874,N_22671,N_22791);
xnor U22875 (N_22875,N_22721,N_22621);
or U22876 (N_22876,N_22634,N_22626);
and U22877 (N_22877,N_22745,N_22773);
xnor U22878 (N_22878,N_22663,N_22665);
and U22879 (N_22879,N_22774,N_22628);
nand U22880 (N_22880,N_22741,N_22690);
nor U22881 (N_22881,N_22617,N_22638);
nor U22882 (N_22882,N_22781,N_22609);
or U22883 (N_22883,N_22697,N_22737);
and U22884 (N_22884,N_22603,N_22709);
and U22885 (N_22885,N_22767,N_22702);
and U22886 (N_22886,N_22780,N_22725);
nand U22887 (N_22887,N_22700,N_22677);
nand U22888 (N_22888,N_22763,N_22722);
and U22889 (N_22889,N_22712,N_22755);
nand U22890 (N_22890,N_22795,N_22672);
xnor U22891 (N_22891,N_22785,N_22748);
xor U22892 (N_22892,N_22658,N_22766);
and U22893 (N_22893,N_22688,N_22719);
or U22894 (N_22894,N_22687,N_22705);
nor U22895 (N_22895,N_22784,N_22762);
or U22896 (N_22896,N_22723,N_22676);
nand U22897 (N_22897,N_22771,N_22646);
nor U22898 (N_22898,N_22770,N_22640);
nor U22899 (N_22899,N_22696,N_22768);
nor U22900 (N_22900,N_22778,N_22750);
xor U22901 (N_22901,N_22706,N_22718);
xnor U22902 (N_22902,N_22662,N_22720);
nor U22903 (N_22903,N_22673,N_22717);
xnor U22904 (N_22904,N_22670,N_22795);
and U22905 (N_22905,N_22736,N_22753);
and U22906 (N_22906,N_22707,N_22794);
or U22907 (N_22907,N_22715,N_22733);
or U22908 (N_22908,N_22785,N_22763);
xnor U22909 (N_22909,N_22701,N_22652);
or U22910 (N_22910,N_22734,N_22784);
nor U22911 (N_22911,N_22688,N_22777);
or U22912 (N_22912,N_22677,N_22680);
xor U22913 (N_22913,N_22783,N_22604);
xnor U22914 (N_22914,N_22649,N_22758);
nand U22915 (N_22915,N_22694,N_22761);
nor U22916 (N_22916,N_22754,N_22652);
nand U22917 (N_22917,N_22681,N_22799);
or U22918 (N_22918,N_22649,N_22612);
and U22919 (N_22919,N_22689,N_22787);
xnor U22920 (N_22920,N_22793,N_22765);
or U22921 (N_22921,N_22614,N_22785);
or U22922 (N_22922,N_22628,N_22757);
or U22923 (N_22923,N_22672,N_22761);
nor U22924 (N_22924,N_22707,N_22614);
or U22925 (N_22925,N_22789,N_22763);
xor U22926 (N_22926,N_22693,N_22771);
and U22927 (N_22927,N_22679,N_22684);
xnor U22928 (N_22928,N_22712,N_22798);
nor U22929 (N_22929,N_22606,N_22621);
nand U22930 (N_22930,N_22794,N_22780);
and U22931 (N_22931,N_22706,N_22745);
nand U22932 (N_22932,N_22637,N_22610);
nand U22933 (N_22933,N_22745,N_22701);
or U22934 (N_22934,N_22765,N_22641);
nor U22935 (N_22935,N_22658,N_22606);
or U22936 (N_22936,N_22722,N_22696);
or U22937 (N_22937,N_22674,N_22660);
and U22938 (N_22938,N_22628,N_22688);
or U22939 (N_22939,N_22730,N_22741);
or U22940 (N_22940,N_22700,N_22734);
or U22941 (N_22941,N_22690,N_22621);
xor U22942 (N_22942,N_22677,N_22725);
nand U22943 (N_22943,N_22763,N_22729);
or U22944 (N_22944,N_22724,N_22687);
nor U22945 (N_22945,N_22721,N_22666);
and U22946 (N_22946,N_22649,N_22786);
and U22947 (N_22947,N_22637,N_22770);
and U22948 (N_22948,N_22736,N_22648);
or U22949 (N_22949,N_22768,N_22783);
nor U22950 (N_22950,N_22633,N_22638);
xor U22951 (N_22951,N_22663,N_22762);
nand U22952 (N_22952,N_22679,N_22608);
and U22953 (N_22953,N_22700,N_22690);
nand U22954 (N_22954,N_22606,N_22767);
xnor U22955 (N_22955,N_22728,N_22620);
or U22956 (N_22956,N_22678,N_22603);
xor U22957 (N_22957,N_22720,N_22738);
xnor U22958 (N_22958,N_22781,N_22756);
xnor U22959 (N_22959,N_22714,N_22621);
nand U22960 (N_22960,N_22767,N_22616);
nor U22961 (N_22961,N_22744,N_22755);
or U22962 (N_22962,N_22682,N_22755);
xor U22963 (N_22963,N_22796,N_22630);
nor U22964 (N_22964,N_22676,N_22785);
nand U22965 (N_22965,N_22714,N_22764);
nor U22966 (N_22966,N_22678,N_22626);
nor U22967 (N_22967,N_22639,N_22629);
nor U22968 (N_22968,N_22723,N_22747);
and U22969 (N_22969,N_22645,N_22606);
and U22970 (N_22970,N_22612,N_22639);
or U22971 (N_22971,N_22601,N_22621);
or U22972 (N_22972,N_22667,N_22633);
nor U22973 (N_22973,N_22766,N_22742);
nand U22974 (N_22974,N_22670,N_22623);
and U22975 (N_22975,N_22655,N_22728);
and U22976 (N_22976,N_22729,N_22786);
or U22977 (N_22977,N_22757,N_22731);
xnor U22978 (N_22978,N_22638,N_22793);
nand U22979 (N_22979,N_22659,N_22610);
xnor U22980 (N_22980,N_22606,N_22676);
xor U22981 (N_22981,N_22602,N_22757);
or U22982 (N_22982,N_22780,N_22612);
xnor U22983 (N_22983,N_22710,N_22729);
nor U22984 (N_22984,N_22711,N_22660);
and U22985 (N_22985,N_22719,N_22655);
xnor U22986 (N_22986,N_22687,N_22697);
xnor U22987 (N_22987,N_22662,N_22648);
or U22988 (N_22988,N_22735,N_22678);
or U22989 (N_22989,N_22799,N_22735);
and U22990 (N_22990,N_22708,N_22748);
nor U22991 (N_22991,N_22643,N_22627);
xor U22992 (N_22992,N_22778,N_22685);
or U22993 (N_22993,N_22691,N_22740);
nand U22994 (N_22994,N_22619,N_22670);
xor U22995 (N_22995,N_22757,N_22799);
nor U22996 (N_22996,N_22665,N_22636);
nor U22997 (N_22997,N_22782,N_22690);
nand U22998 (N_22998,N_22656,N_22687);
xnor U22999 (N_22999,N_22731,N_22780);
xnor U23000 (N_23000,N_22911,N_22843);
nor U23001 (N_23001,N_22828,N_22856);
nor U23002 (N_23002,N_22853,N_22859);
or U23003 (N_23003,N_22937,N_22998);
and U23004 (N_23004,N_22972,N_22973);
or U23005 (N_23005,N_22835,N_22925);
nor U23006 (N_23006,N_22882,N_22826);
and U23007 (N_23007,N_22806,N_22905);
nor U23008 (N_23008,N_22906,N_22938);
xnor U23009 (N_23009,N_22935,N_22840);
xor U23010 (N_23010,N_22805,N_22804);
xnor U23011 (N_23011,N_22893,N_22866);
nor U23012 (N_23012,N_22999,N_22966);
nand U23013 (N_23013,N_22936,N_22967);
xor U23014 (N_23014,N_22931,N_22957);
nand U23015 (N_23015,N_22946,N_22948);
nor U23016 (N_23016,N_22894,N_22941);
xor U23017 (N_23017,N_22961,N_22824);
xnor U23018 (N_23018,N_22845,N_22953);
xnor U23019 (N_23019,N_22872,N_22993);
or U23020 (N_23020,N_22817,N_22958);
xnor U23021 (N_23021,N_22907,N_22871);
or U23022 (N_23022,N_22991,N_22877);
and U23023 (N_23023,N_22858,N_22811);
or U23024 (N_23024,N_22968,N_22976);
nor U23025 (N_23025,N_22926,N_22801);
or U23026 (N_23026,N_22880,N_22965);
or U23027 (N_23027,N_22832,N_22841);
xor U23028 (N_23028,N_22848,N_22921);
xnor U23029 (N_23029,N_22833,N_22932);
nor U23030 (N_23030,N_22974,N_22943);
or U23031 (N_23031,N_22971,N_22928);
nand U23032 (N_23032,N_22977,N_22881);
and U23033 (N_23033,N_22969,N_22949);
and U23034 (N_23034,N_22803,N_22890);
and U23035 (N_23035,N_22989,N_22984);
or U23036 (N_23036,N_22908,N_22836);
and U23037 (N_23037,N_22954,N_22887);
nand U23038 (N_23038,N_22838,N_22822);
nand U23039 (N_23039,N_22963,N_22896);
nor U23040 (N_23040,N_22997,N_22874);
nor U23041 (N_23041,N_22883,N_22952);
xnor U23042 (N_23042,N_22902,N_22915);
or U23043 (N_23043,N_22903,N_22947);
xor U23044 (N_23044,N_22844,N_22919);
nand U23045 (N_23045,N_22829,N_22873);
nor U23046 (N_23046,N_22852,N_22847);
nor U23047 (N_23047,N_22855,N_22885);
nor U23048 (N_23048,N_22809,N_22980);
nor U23049 (N_23049,N_22864,N_22945);
xor U23050 (N_23050,N_22970,N_22960);
nor U23051 (N_23051,N_22933,N_22955);
nor U23052 (N_23052,N_22854,N_22900);
nor U23053 (N_23053,N_22819,N_22850);
nand U23054 (N_23054,N_22994,N_22897);
xnor U23055 (N_23055,N_22918,N_22888);
or U23056 (N_23056,N_22862,N_22892);
nand U23057 (N_23057,N_22868,N_22870);
nor U23058 (N_23058,N_22879,N_22816);
nand U23059 (N_23059,N_22812,N_22814);
nor U23060 (N_23060,N_22962,N_22810);
nor U23061 (N_23061,N_22807,N_22867);
nand U23062 (N_23062,N_22861,N_22820);
nor U23063 (N_23063,N_22985,N_22982);
nor U23064 (N_23064,N_22916,N_22878);
nand U23065 (N_23065,N_22964,N_22979);
nand U23066 (N_23066,N_22899,N_22863);
or U23067 (N_23067,N_22975,N_22865);
xnor U23068 (N_23068,N_22914,N_22901);
nor U23069 (N_23069,N_22808,N_22818);
nand U23070 (N_23070,N_22889,N_22800);
nand U23071 (N_23071,N_22951,N_22912);
xnor U23072 (N_23072,N_22825,N_22891);
nor U23073 (N_23073,N_22988,N_22875);
or U23074 (N_23074,N_22851,N_22815);
nor U23075 (N_23075,N_22940,N_22830);
or U23076 (N_23076,N_22959,N_22986);
or U23077 (N_23077,N_22860,N_22922);
or U23078 (N_23078,N_22942,N_22929);
nand U23079 (N_23079,N_22813,N_22834);
and U23080 (N_23080,N_22857,N_22823);
nand U23081 (N_23081,N_22944,N_22884);
and U23082 (N_23082,N_22898,N_22924);
or U23083 (N_23083,N_22895,N_22930);
xnor U23084 (N_23084,N_22827,N_22842);
or U23085 (N_23085,N_22992,N_22869);
and U23086 (N_23086,N_22923,N_22996);
or U23087 (N_23087,N_22983,N_22990);
xor U23088 (N_23088,N_22846,N_22939);
nand U23089 (N_23089,N_22978,N_22904);
and U23090 (N_23090,N_22876,N_22920);
xnor U23091 (N_23091,N_22839,N_22802);
xnor U23092 (N_23092,N_22910,N_22913);
or U23093 (N_23093,N_22981,N_22950);
xor U23094 (N_23094,N_22934,N_22886);
xor U23095 (N_23095,N_22927,N_22995);
nor U23096 (N_23096,N_22909,N_22837);
xor U23097 (N_23097,N_22821,N_22987);
nand U23098 (N_23098,N_22917,N_22849);
or U23099 (N_23099,N_22956,N_22831);
and U23100 (N_23100,N_22899,N_22957);
nand U23101 (N_23101,N_22976,N_22906);
or U23102 (N_23102,N_22853,N_22851);
and U23103 (N_23103,N_22845,N_22874);
nand U23104 (N_23104,N_22986,N_22911);
nor U23105 (N_23105,N_22967,N_22953);
xor U23106 (N_23106,N_22922,N_22854);
nor U23107 (N_23107,N_22927,N_22924);
and U23108 (N_23108,N_22800,N_22856);
xnor U23109 (N_23109,N_22826,N_22986);
nand U23110 (N_23110,N_22945,N_22926);
or U23111 (N_23111,N_22846,N_22894);
and U23112 (N_23112,N_22901,N_22905);
nand U23113 (N_23113,N_22902,N_22944);
and U23114 (N_23114,N_22821,N_22889);
nor U23115 (N_23115,N_22945,N_22821);
nor U23116 (N_23116,N_22835,N_22927);
xnor U23117 (N_23117,N_22821,N_22817);
nand U23118 (N_23118,N_22800,N_22969);
nand U23119 (N_23119,N_22916,N_22800);
and U23120 (N_23120,N_22903,N_22869);
nor U23121 (N_23121,N_22844,N_22806);
xor U23122 (N_23122,N_22909,N_22962);
nor U23123 (N_23123,N_22956,N_22896);
nand U23124 (N_23124,N_22999,N_22959);
xor U23125 (N_23125,N_22941,N_22954);
nand U23126 (N_23126,N_22809,N_22916);
or U23127 (N_23127,N_22947,N_22841);
xor U23128 (N_23128,N_22834,N_22995);
xnor U23129 (N_23129,N_22968,N_22855);
and U23130 (N_23130,N_22972,N_22977);
xnor U23131 (N_23131,N_22959,N_22850);
nand U23132 (N_23132,N_22861,N_22813);
or U23133 (N_23133,N_22973,N_22949);
nand U23134 (N_23134,N_22878,N_22997);
nand U23135 (N_23135,N_22897,N_22900);
or U23136 (N_23136,N_22987,N_22803);
or U23137 (N_23137,N_22980,N_22953);
xor U23138 (N_23138,N_22955,N_22869);
nand U23139 (N_23139,N_22917,N_22837);
or U23140 (N_23140,N_22900,N_22940);
or U23141 (N_23141,N_22984,N_22897);
xnor U23142 (N_23142,N_22895,N_22938);
nand U23143 (N_23143,N_22877,N_22985);
nand U23144 (N_23144,N_22815,N_22807);
nand U23145 (N_23145,N_22803,N_22978);
xnor U23146 (N_23146,N_22982,N_22938);
nand U23147 (N_23147,N_22873,N_22869);
xor U23148 (N_23148,N_22823,N_22929);
nand U23149 (N_23149,N_22972,N_22889);
xor U23150 (N_23150,N_22821,N_22941);
or U23151 (N_23151,N_22903,N_22800);
and U23152 (N_23152,N_22883,N_22936);
xnor U23153 (N_23153,N_22949,N_22921);
or U23154 (N_23154,N_22988,N_22964);
nor U23155 (N_23155,N_22820,N_22944);
and U23156 (N_23156,N_22927,N_22905);
or U23157 (N_23157,N_22941,N_22825);
xnor U23158 (N_23158,N_22945,N_22810);
and U23159 (N_23159,N_22947,N_22956);
and U23160 (N_23160,N_22983,N_22818);
or U23161 (N_23161,N_22873,N_22934);
and U23162 (N_23162,N_22874,N_22903);
xor U23163 (N_23163,N_22999,N_22834);
nor U23164 (N_23164,N_22940,N_22943);
nand U23165 (N_23165,N_22838,N_22961);
xnor U23166 (N_23166,N_22927,N_22844);
or U23167 (N_23167,N_22918,N_22812);
and U23168 (N_23168,N_22872,N_22895);
and U23169 (N_23169,N_22881,N_22832);
nand U23170 (N_23170,N_22987,N_22929);
nand U23171 (N_23171,N_22969,N_22978);
and U23172 (N_23172,N_22846,N_22893);
or U23173 (N_23173,N_22829,N_22819);
xor U23174 (N_23174,N_22885,N_22918);
xor U23175 (N_23175,N_22944,N_22979);
nor U23176 (N_23176,N_22872,N_22847);
nand U23177 (N_23177,N_22906,N_22962);
or U23178 (N_23178,N_22893,N_22860);
nand U23179 (N_23179,N_22912,N_22952);
nor U23180 (N_23180,N_22946,N_22958);
xor U23181 (N_23181,N_22977,N_22847);
and U23182 (N_23182,N_22816,N_22847);
nand U23183 (N_23183,N_22976,N_22840);
and U23184 (N_23184,N_22919,N_22804);
nor U23185 (N_23185,N_22958,N_22803);
and U23186 (N_23186,N_22974,N_22877);
and U23187 (N_23187,N_22952,N_22925);
or U23188 (N_23188,N_22906,N_22972);
nand U23189 (N_23189,N_22874,N_22842);
nand U23190 (N_23190,N_22823,N_22849);
xnor U23191 (N_23191,N_22929,N_22818);
nor U23192 (N_23192,N_22867,N_22983);
nor U23193 (N_23193,N_22936,N_22870);
nand U23194 (N_23194,N_22953,N_22820);
or U23195 (N_23195,N_22943,N_22936);
and U23196 (N_23196,N_22954,N_22990);
xnor U23197 (N_23197,N_22859,N_22949);
nor U23198 (N_23198,N_22998,N_22995);
nand U23199 (N_23199,N_22882,N_22920);
or U23200 (N_23200,N_23192,N_23167);
nor U23201 (N_23201,N_23103,N_23182);
and U23202 (N_23202,N_23164,N_23187);
and U23203 (N_23203,N_23124,N_23175);
nand U23204 (N_23204,N_23156,N_23041);
and U23205 (N_23205,N_23189,N_23030);
xnor U23206 (N_23206,N_23151,N_23054);
or U23207 (N_23207,N_23093,N_23057);
xnor U23208 (N_23208,N_23018,N_23010);
or U23209 (N_23209,N_23078,N_23110);
xnor U23210 (N_23210,N_23123,N_23120);
nor U23211 (N_23211,N_23162,N_23101);
nor U23212 (N_23212,N_23085,N_23102);
nor U23213 (N_23213,N_23161,N_23111);
nor U23214 (N_23214,N_23193,N_23027);
xor U23215 (N_23215,N_23055,N_23038);
nor U23216 (N_23216,N_23056,N_23084);
nand U23217 (N_23217,N_23002,N_23012);
and U23218 (N_23218,N_23152,N_23019);
nor U23219 (N_23219,N_23034,N_23097);
nor U23220 (N_23220,N_23089,N_23092);
xnor U23221 (N_23221,N_23134,N_23170);
nor U23222 (N_23222,N_23113,N_23063);
and U23223 (N_23223,N_23122,N_23090);
and U23224 (N_23224,N_23119,N_23032);
and U23225 (N_23225,N_23100,N_23066);
nor U23226 (N_23226,N_23118,N_23068);
or U23227 (N_23227,N_23052,N_23138);
and U23228 (N_23228,N_23165,N_23195);
xnor U23229 (N_23229,N_23194,N_23053);
nand U23230 (N_23230,N_23001,N_23174);
and U23231 (N_23231,N_23070,N_23000);
nand U23232 (N_23232,N_23091,N_23033);
xnor U23233 (N_23233,N_23076,N_23062);
xnor U23234 (N_23234,N_23140,N_23139);
and U23235 (N_23235,N_23177,N_23096);
nor U23236 (N_23236,N_23005,N_23071);
and U23237 (N_23237,N_23011,N_23014);
or U23238 (N_23238,N_23108,N_23130);
xnor U23239 (N_23239,N_23025,N_23022);
and U23240 (N_23240,N_23143,N_23171);
nand U23241 (N_23241,N_23135,N_23048);
and U23242 (N_23242,N_23147,N_23026);
or U23243 (N_23243,N_23109,N_23107);
and U23244 (N_23244,N_23043,N_23039);
xnor U23245 (N_23245,N_23186,N_23080);
and U23246 (N_23246,N_23094,N_23082);
or U23247 (N_23247,N_23172,N_23028);
nor U23248 (N_23248,N_23035,N_23188);
xnor U23249 (N_23249,N_23146,N_23099);
or U23250 (N_23250,N_23142,N_23159);
and U23251 (N_23251,N_23088,N_23023);
nor U23252 (N_23252,N_23067,N_23045);
nand U23253 (N_23253,N_23169,N_23003);
nor U23254 (N_23254,N_23006,N_23086);
nand U23255 (N_23255,N_23069,N_23051);
nor U23256 (N_23256,N_23058,N_23180);
nand U23257 (N_23257,N_23029,N_23197);
nor U23258 (N_23258,N_23072,N_23061);
nand U23259 (N_23259,N_23105,N_23129);
nor U23260 (N_23260,N_23112,N_23144);
and U23261 (N_23261,N_23149,N_23168);
nand U23262 (N_23262,N_23148,N_23004);
nand U23263 (N_23263,N_23199,N_23037);
and U23264 (N_23264,N_23183,N_23074);
nand U23265 (N_23265,N_23166,N_23160);
nor U23266 (N_23266,N_23191,N_23184);
or U23267 (N_23267,N_23150,N_23190);
and U23268 (N_23268,N_23021,N_23024);
nor U23269 (N_23269,N_23128,N_23073);
or U23270 (N_23270,N_23137,N_23009);
nor U23271 (N_23271,N_23007,N_23181);
nand U23272 (N_23272,N_23013,N_23098);
or U23273 (N_23273,N_23046,N_23136);
nor U23274 (N_23274,N_23008,N_23075);
or U23275 (N_23275,N_23040,N_23017);
nand U23276 (N_23276,N_23042,N_23083);
or U23277 (N_23277,N_23047,N_23020);
nor U23278 (N_23278,N_23015,N_23115);
nand U23279 (N_23279,N_23117,N_23153);
and U23280 (N_23280,N_23060,N_23157);
nor U23281 (N_23281,N_23087,N_23064);
xor U23282 (N_23282,N_23125,N_23065);
nand U23283 (N_23283,N_23196,N_23121);
nand U23284 (N_23284,N_23114,N_23176);
nand U23285 (N_23285,N_23059,N_23106);
or U23286 (N_23286,N_23116,N_23127);
and U23287 (N_23287,N_23185,N_23154);
and U23288 (N_23288,N_23179,N_23016);
and U23289 (N_23289,N_23158,N_23081);
or U23290 (N_23290,N_23126,N_23095);
nor U23291 (N_23291,N_23131,N_23173);
or U23292 (N_23292,N_23031,N_23077);
or U23293 (N_23293,N_23198,N_23163);
xnor U23294 (N_23294,N_23050,N_23133);
xor U23295 (N_23295,N_23132,N_23141);
nand U23296 (N_23296,N_23104,N_23145);
xor U23297 (N_23297,N_23178,N_23079);
or U23298 (N_23298,N_23036,N_23049);
and U23299 (N_23299,N_23155,N_23044);
or U23300 (N_23300,N_23070,N_23109);
nand U23301 (N_23301,N_23029,N_23199);
nand U23302 (N_23302,N_23198,N_23083);
nand U23303 (N_23303,N_23001,N_23190);
nand U23304 (N_23304,N_23045,N_23080);
nor U23305 (N_23305,N_23133,N_23068);
nand U23306 (N_23306,N_23037,N_23017);
or U23307 (N_23307,N_23006,N_23134);
nand U23308 (N_23308,N_23048,N_23170);
and U23309 (N_23309,N_23152,N_23128);
or U23310 (N_23310,N_23196,N_23003);
or U23311 (N_23311,N_23063,N_23131);
and U23312 (N_23312,N_23112,N_23164);
nor U23313 (N_23313,N_23073,N_23011);
and U23314 (N_23314,N_23097,N_23088);
nand U23315 (N_23315,N_23032,N_23033);
and U23316 (N_23316,N_23095,N_23123);
nor U23317 (N_23317,N_23164,N_23166);
and U23318 (N_23318,N_23003,N_23173);
or U23319 (N_23319,N_23092,N_23054);
nand U23320 (N_23320,N_23042,N_23157);
and U23321 (N_23321,N_23164,N_23146);
nor U23322 (N_23322,N_23035,N_23141);
or U23323 (N_23323,N_23122,N_23139);
or U23324 (N_23324,N_23156,N_23024);
nand U23325 (N_23325,N_23004,N_23172);
or U23326 (N_23326,N_23041,N_23167);
or U23327 (N_23327,N_23082,N_23009);
and U23328 (N_23328,N_23159,N_23132);
nand U23329 (N_23329,N_23004,N_23040);
xnor U23330 (N_23330,N_23130,N_23128);
xor U23331 (N_23331,N_23105,N_23067);
and U23332 (N_23332,N_23188,N_23059);
nor U23333 (N_23333,N_23036,N_23128);
or U23334 (N_23334,N_23107,N_23058);
or U23335 (N_23335,N_23162,N_23125);
nand U23336 (N_23336,N_23109,N_23166);
xnor U23337 (N_23337,N_23157,N_23088);
or U23338 (N_23338,N_23058,N_23025);
or U23339 (N_23339,N_23073,N_23157);
nor U23340 (N_23340,N_23175,N_23119);
or U23341 (N_23341,N_23095,N_23146);
nand U23342 (N_23342,N_23187,N_23112);
and U23343 (N_23343,N_23142,N_23060);
and U23344 (N_23344,N_23184,N_23050);
or U23345 (N_23345,N_23045,N_23111);
nor U23346 (N_23346,N_23167,N_23026);
nand U23347 (N_23347,N_23112,N_23129);
nand U23348 (N_23348,N_23166,N_23184);
nor U23349 (N_23349,N_23170,N_23043);
nand U23350 (N_23350,N_23053,N_23001);
nand U23351 (N_23351,N_23178,N_23142);
or U23352 (N_23352,N_23022,N_23018);
and U23353 (N_23353,N_23083,N_23039);
nor U23354 (N_23354,N_23179,N_23156);
and U23355 (N_23355,N_23028,N_23058);
and U23356 (N_23356,N_23036,N_23180);
or U23357 (N_23357,N_23136,N_23188);
and U23358 (N_23358,N_23168,N_23188);
xor U23359 (N_23359,N_23083,N_23024);
nor U23360 (N_23360,N_23149,N_23117);
xnor U23361 (N_23361,N_23148,N_23101);
and U23362 (N_23362,N_23042,N_23170);
nor U23363 (N_23363,N_23111,N_23064);
nand U23364 (N_23364,N_23179,N_23069);
nor U23365 (N_23365,N_23075,N_23148);
or U23366 (N_23366,N_23060,N_23019);
nor U23367 (N_23367,N_23092,N_23062);
xor U23368 (N_23368,N_23154,N_23072);
nand U23369 (N_23369,N_23071,N_23155);
and U23370 (N_23370,N_23170,N_23117);
and U23371 (N_23371,N_23011,N_23182);
nand U23372 (N_23372,N_23035,N_23184);
nor U23373 (N_23373,N_23126,N_23010);
nand U23374 (N_23374,N_23054,N_23008);
xnor U23375 (N_23375,N_23180,N_23169);
and U23376 (N_23376,N_23186,N_23173);
or U23377 (N_23377,N_23027,N_23111);
nand U23378 (N_23378,N_23139,N_23034);
or U23379 (N_23379,N_23010,N_23033);
and U23380 (N_23380,N_23039,N_23172);
or U23381 (N_23381,N_23184,N_23117);
nor U23382 (N_23382,N_23141,N_23007);
xor U23383 (N_23383,N_23115,N_23095);
or U23384 (N_23384,N_23023,N_23060);
nand U23385 (N_23385,N_23123,N_23075);
and U23386 (N_23386,N_23056,N_23195);
xnor U23387 (N_23387,N_23180,N_23140);
nand U23388 (N_23388,N_23168,N_23139);
nand U23389 (N_23389,N_23171,N_23037);
or U23390 (N_23390,N_23062,N_23052);
xor U23391 (N_23391,N_23074,N_23098);
or U23392 (N_23392,N_23166,N_23097);
nor U23393 (N_23393,N_23165,N_23126);
nor U23394 (N_23394,N_23193,N_23178);
nor U23395 (N_23395,N_23152,N_23130);
xor U23396 (N_23396,N_23015,N_23155);
nand U23397 (N_23397,N_23166,N_23016);
and U23398 (N_23398,N_23195,N_23064);
nor U23399 (N_23399,N_23045,N_23125);
nand U23400 (N_23400,N_23261,N_23395);
xor U23401 (N_23401,N_23228,N_23327);
nor U23402 (N_23402,N_23341,N_23264);
nor U23403 (N_23403,N_23263,N_23353);
nor U23404 (N_23404,N_23206,N_23396);
and U23405 (N_23405,N_23233,N_23271);
nand U23406 (N_23406,N_23212,N_23289);
nand U23407 (N_23407,N_23336,N_23201);
and U23408 (N_23408,N_23399,N_23290);
and U23409 (N_23409,N_23256,N_23235);
nand U23410 (N_23410,N_23314,N_23357);
xnor U23411 (N_23411,N_23282,N_23268);
nor U23412 (N_23412,N_23223,N_23234);
nor U23413 (N_23413,N_23245,N_23346);
nor U23414 (N_23414,N_23302,N_23269);
nor U23415 (N_23415,N_23366,N_23277);
xor U23416 (N_23416,N_23211,N_23205);
or U23417 (N_23417,N_23296,N_23279);
nor U23418 (N_23418,N_23257,N_23318);
nand U23419 (N_23419,N_23379,N_23326);
nand U23420 (N_23420,N_23320,N_23335);
or U23421 (N_23421,N_23309,N_23312);
and U23422 (N_23422,N_23363,N_23342);
nand U23423 (N_23423,N_23299,N_23325);
and U23424 (N_23424,N_23242,N_23390);
nor U23425 (N_23425,N_23291,N_23221);
xor U23426 (N_23426,N_23367,N_23267);
and U23427 (N_23427,N_23361,N_23344);
and U23428 (N_23428,N_23255,N_23238);
nor U23429 (N_23429,N_23278,N_23338);
nand U23430 (N_23430,N_23392,N_23208);
nand U23431 (N_23431,N_23343,N_23377);
or U23432 (N_23432,N_23224,N_23324);
or U23433 (N_23433,N_23382,N_23337);
nand U23434 (N_23434,N_23253,N_23360);
and U23435 (N_23435,N_23378,N_23281);
xor U23436 (N_23436,N_23389,N_23213);
and U23437 (N_23437,N_23200,N_23293);
nor U23438 (N_23438,N_23297,N_23243);
nand U23439 (N_23439,N_23215,N_23207);
nand U23440 (N_23440,N_23246,N_23348);
and U23441 (N_23441,N_23364,N_23219);
and U23442 (N_23442,N_23316,N_23359);
or U23443 (N_23443,N_23301,N_23210);
nand U23444 (N_23444,N_23373,N_23332);
nand U23445 (N_23445,N_23352,N_23250);
xnor U23446 (N_23446,N_23249,N_23272);
or U23447 (N_23447,N_23376,N_23305);
xor U23448 (N_23448,N_23322,N_23231);
nand U23449 (N_23449,N_23329,N_23240);
nor U23450 (N_23450,N_23273,N_23350);
nor U23451 (N_23451,N_23230,N_23391);
xor U23452 (N_23452,N_23217,N_23384);
or U23453 (N_23453,N_23274,N_23260);
xor U23454 (N_23454,N_23351,N_23317);
or U23455 (N_23455,N_23345,N_23303);
nand U23456 (N_23456,N_23319,N_23298);
or U23457 (N_23457,N_23294,N_23209);
nor U23458 (N_23458,N_23270,N_23365);
or U23459 (N_23459,N_23368,N_23288);
nand U23460 (N_23460,N_23331,N_23333);
nand U23461 (N_23461,N_23374,N_23387);
nor U23462 (N_23462,N_23306,N_23244);
xnor U23463 (N_23463,N_23330,N_23258);
xor U23464 (N_23464,N_23315,N_23251);
nand U23465 (N_23465,N_23356,N_23310);
xor U23466 (N_23466,N_23248,N_23383);
xnor U23467 (N_23467,N_23328,N_23216);
or U23468 (N_23468,N_23292,N_23227);
or U23469 (N_23469,N_23241,N_23236);
nand U23470 (N_23470,N_23225,N_23304);
nand U23471 (N_23471,N_23375,N_23283);
xor U23472 (N_23472,N_23295,N_23347);
and U23473 (N_23473,N_23266,N_23308);
xnor U23474 (N_23474,N_23385,N_23321);
and U23475 (N_23475,N_23388,N_23218);
nand U23476 (N_23476,N_23203,N_23204);
nand U23477 (N_23477,N_23394,N_23226);
nor U23478 (N_23478,N_23202,N_23254);
or U23479 (N_23479,N_23354,N_23370);
or U23480 (N_23480,N_23280,N_23334);
nand U23481 (N_23481,N_23339,N_23232);
xnor U23482 (N_23482,N_23259,N_23276);
or U23483 (N_23483,N_23252,N_23313);
nor U23484 (N_23484,N_23284,N_23371);
nand U23485 (N_23485,N_23340,N_23393);
nor U23486 (N_23486,N_23237,N_23311);
nor U23487 (N_23487,N_23398,N_23369);
or U23488 (N_23488,N_23286,N_23381);
and U23489 (N_23489,N_23323,N_23372);
and U23490 (N_23490,N_23229,N_23214);
nor U23491 (N_23491,N_23355,N_23220);
and U23492 (N_23492,N_23285,N_23275);
and U23493 (N_23493,N_23307,N_23358);
nor U23494 (N_23494,N_23262,N_23265);
or U23495 (N_23495,N_23222,N_23349);
nand U23496 (N_23496,N_23362,N_23247);
nand U23497 (N_23497,N_23287,N_23397);
and U23498 (N_23498,N_23380,N_23300);
and U23499 (N_23499,N_23239,N_23386);
xor U23500 (N_23500,N_23216,N_23244);
nand U23501 (N_23501,N_23324,N_23357);
xnor U23502 (N_23502,N_23260,N_23212);
nor U23503 (N_23503,N_23244,N_23335);
xnor U23504 (N_23504,N_23222,N_23247);
nand U23505 (N_23505,N_23218,N_23398);
nand U23506 (N_23506,N_23375,N_23271);
or U23507 (N_23507,N_23311,N_23328);
and U23508 (N_23508,N_23356,N_23240);
nor U23509 (N_23509,N_23275,N_23339);
nand U23510 (N_23510,N_23311,N_23368);
nor U23511 (N_23511,N_23330,N_23260);
nand U23512 (N_23512,N_23383,N_23230);
nand U23513 (N_23513,N_23281,N_23290);
or U23514 (N_23514,N_23211,N_23361);
and U23515 (N_23515,N_23388,N_23282);
xor U23516 (N_23516,N_23215,N_23370);
nor U23517 (N_23517,N_23219,N_23288);
and U23518 (N_23518,N_23274,N_23319);
or U23519 (N_23519,N_23374,N_23298);
nand U23520 (N_23520,N_23383,N_23354);
xor U23521 (N_23521,N_23305,N_23313);
and U23522 (N_23522,N_23228,N_23316);
and U23523 (N_23523,N_23291,N_23354);
xnor U23524 (N_23524,N_23326,N_23213);
nand U23525 (N_23525,N_23351,N_23390);
nor U23526 (N_23526,N_23208,N_23366);
xor U23527 (N_23527,N_23238,N_23319);
xnor U23528 (N_23528,N_23311,N_23292);
nand U23529 (N_23529,N_23358,N_23250);
nor U23530 (N_23530,N_23231,N_23300);
and U23531 (N_23531,N_23303,N_23233);
nand U23532 (N_23532,N_23362,N_23376);
or U23533 (N_23533,N_23286,N_23240);
nor U23534 (N_23534,N_23393,N_23325);
xor U23535 (N_23535,N_23335,N_23358);
nand U23536 (N_23536,N_23350,N_23391);
xor U23537 (N_23537,N_23340,N_23241);
xor U23538 (N_23538,N_23282,N_23288);
and U23539 (N_23539,N_23295,N_23383);
xnor U23540 (N_23540,N_23353,N_23314);
nor U23541 (N_23541,N_23383,N_23214);
nand U23542 (N_23542,N_23310,N_23334);
xnor U23543 (N_23543,N_23343,N_23257);
xor U23544 (N_23544,N_23231,N_23360);
nor U23545 (N_23545,N_23360,N_23295);
nor U23546 (N_23546,N_23318,N_23384);
xnor U23547 (N_23547,N_23354,N_23379);
nor U23548 (N_23548,N_23365,N_23325);
nand U23549 (N_23549,N_23392,N_23382);
xnor U23550 (N_23550,N_23226,N_23359);
nand U23551 (N_23551,N_23373,N_23229);
nor U23552 (N_23552,N_23324,N_23300);
nand U23553 (N_23553,N_23272,N_23289);
nor U23554 (N_23554,N_23239,N_23231);
xnor U23555 (N_23555,N_23226,N_23279);
and U23556 (N_23556,N_23315,N_23388);
and U23557 (N_23557,N_23348,N_23280);
nand U23558 (N_23558,N_23225,N_23220);
or U23559 (N_23559,N_23336,N_23347);
nand U23560 (N_23560,N_23209,N_23253);
nand U23561 (N_23561,N_23226,N_23305);
xnor U23562 (N_23562,N_23367,N_23236);
and U23563 (N_23563,N_23216,N_23373);
nor U23564 (N_23564,N_23231,N_23293);
xnor U23565 (N_23565,N_23208,N_23239);
and U23566 (N_23566,N_23220,N_23375);
or U23567 (N_23567,N_23369,N_23272);
nor U23568 (N_23568,N_23202,N_23277);
xor U23569 (N_23569,N_23247,N_23316);
and U23570 (N_23570,N_23278,N_23391);
and U23571 (N_23571,N_23252,N_23217);
xor U23572 (N_23572,N_23287,N_23344);
and U23573 (N_23573,N_23380,N_23293);
or U23574 (N_23574,N_23394,N_23253);
or U23575 (N_23575,N_23395,N_23355);
nor U23576 (N_23576,N_23202,N_23228);
and U23577 (N_23577,N_23325,N_23354);
or U23578 (N_23578,N_23376,N_23246);
nor U23579 (N_23579,N_23291,N_23200);
xnor U23580 (N_23580,N_23302,N_23255);
nor U23581 (N_23581,N_23225,N_23354);
nor U23582 (N_23582,N_23371,N_23307);
nand U23583 (N_23583,N_23364,N_23323);
and U23584 (N_23584,N_23306,N_23259);
nor U23585 (N_23585,N_23288,N_23375);
and U23586 (N_23586,N_23352,N_23259);
xnor U23587 (N_23587,N_23387,N_23222);
nand U23588 (N_23588,N_23218,N_23248);
nand U23589 (N_23589,N_23233,N_23238);
nor U23590 (N_23590,N_23213,N_23385);
nor U23591 (N_23591,N_23295,N_23319);
xnor U23592 (N_23592,N_23255,N_23321);
nor U23593 (N_23593,N_23361,N_23308);
or U23594 (N_23594,N_23281,N_23372);
xnor U23595 (N_23595,N_23371,N_23247);
or U23596 (N_23596,N_23225,N_23387);
or U23597 (N_23597,N_23360,N_23269);
nand U23598 (N_23598,N_23317,N_23361);
nand U23599 (N_23599,N_23248,N_23315);
xnor U23600 (N_23600,N_23530,N_23436);
nand U23601 (N_23601,N_23489,N_23487);
and U23602 (N_23602,N_23539,N_23567);
nor U23603 (N_23603,N_23572,N_23494);
nor U23604 (N_23604,N_23553,N_23479);
nand U23605 (N_23605,N_23552,N_23455);
or U23606 (N_23606,N_23412,N_23585);
nand U23607 (N_23607,N_23467,N_23537);
nand U23608 (N_23608,N_23451,N_23501);
nand U23609 (N_23609,N_23546,N_23437);
nor U23610 (N_23610,N_23497,N_23584);
or U23611 (N_23611,N_23513,N_23470);
and U23612 (N_23612,N_23531,N_23444);
nand U23613 (N_23613,N_23575,N_23550);
nor U23614 (N_23614,N_23430,N_23402);
and U23615 (N_23615,N_23466,N_23411);
nor U23616 (N_23616,N_23505,N_23562);
and U23617 (N_23617,N_23508,N_23596);
nor U23618 (N_23618,N_23533,N_23483);
and U23619 (N_23619,N_23532,N_23558);
xor U23620 (N_23620,N_23565,N_23594);
or U23621 (N_23621,N_23439,N_23473);
and U23622 (N_23622,N_23538,N_23586);
or U23623 (N_23623,N_23477,N_23571);
xor U23624 (N_23624,N_23579,N_23568);
and U23625 (N_23625,N_23516,N_23410);
xnor U23626 (N_23626,N_23441,N_23589);
nand U23627 (N_23627,N_23576,N_23449);
and U23628 (N_23628,N_23559,N_23401);
or U23629 (N_23629,N_23514,N_23423);
xnor U23630 (N_23630,N_23545,N_23534);
and U23631 (N_23631,N_23518,N_23418);
xor U23632 (N_23632,N_23519,N_23464);
xor U23633 (N_23633,N_23438,N_23493);
nand U23634 (N_23634,N_23422,N_23569);
nor U23635 (N_23635,N_23597,N_23485);
nor U23636 (N_23636,N_23446,N_23599);
and U23637 (N_23637,N_23471,N_23529);
nand U23638 (N_23638,N_23406,N_23465);
nand U23639 (N_23639,N_23595,N_23443);
nand U23640 (N_23640,N_23475,N_23424);
nor U23641 (N_23641,N_23598,N_23445);
or U23642 (N_23642,N_23510,N_23442);
xor U23643 (N_23643,N_23582,N_23592);
or U23644 (N_23644,N_23491,N_23428);
nor U23645 (N_23645,N_23419,N_23570);
nand U23646 (N_23646,N_23499,N_23560);
and U23647 (N_23647,N_23506,N_23481);
or U23648 (N_23648,N_23407,N_23504);
and U23649 (N_23649,N_23425,N_23456);
nand U23650 (N_23650,N_23503,N_23429);
nand U23651 (N_23651,N_23408,N_23440);
or U23652 (N_23652,N_23566,N_23509);
nand U23653 (N_23653,N_23453,N_23486);
and U23654 (N_23654,N_23405,N_23452);
xnor U23655 (N_23655,N_23525,N_23414);
and U23656 (N_23656,N_23426,N_23415);
and U23657 (N_23657,N_23502,N_23498);
and U23658 (N_23658,N_23547,N_23581);
nand U23659 (N_23659,N_23578,N_23457);
nand U23660 (N_23660,N_23484,N_23458);
nand U23661 (N_23661,N_23573,N_23536);
nor U23662 (N_23662,N_23587,N_23472);
xnor U23663 (N_23663,N_23432,N_23561);
or U23664 (N_23664,N_23555,N_23522);
xnor U23665 (N_23665,N_23400,N_23460);
and U23666 (N_23666,N_23563,N_23450);
nand U23667 (N_23667,N_23541,N_23462);
nor U23668 (N_23668,N_23459,N_23490);
nand U23669 (N_23669,N_23526,N_23417);
nor U23670 (N_23670,N_23447,N_23461);
nor U23671 (N_23671,N_23556,N_23591);
nor U23672 (N_23672,N_23527,N_23433);
xnor U23673 (N_23673,N_23404,N_23590);
or U23674 (N_23674,N_23434,N_23492);
xnor U23675 (N_23675,N_23517,N_23478);
xnor U23676 (N_23676,N_23403,N_23574);
nand U23677 (N_23677,N_23524,N_23515);
nand U23678 (N_23678,N_23431,N_23463);
xor U23679 (N_23679,N_23495,N_23593);
or U23680 (N_23680,N_23577,N_23482);
xnor U23681 (N_23681,N_23416,N_23488);
nor U23682 (N_23682,N_23549,N_23521);
and U23683 (N_23683,N_23496,N_23557);
nor U23684 (N_23684,N_23548,N_23420);
and U23685 (N_23685,N_23421,N_23454);
nand U23686 (N_23686,N_23500,N_23512);
or U23687 (N_23687,N_23523,N_23551);
and U23688 (N_23688,N_23542,N_23535);
or U23689 (N_23689,N_23543,N_23448);
or U23690 (N_23690,N_23554,N_23480);
nor U23691 (N_23691,N_23427,N_23580);
or U23692 (N_23692,N_23409,N_23476);
nand U23693 (N_23693,N_23413,N_23507);
xnor U23694 (N_23694,N_23520,N_23544);
xnor U23695 (N_23695,N_23583,N_23540);
and U23696 (N_23696,N_23468,N_23588);
nand U23697 (N_23697,N_23474,N_23435);
or U23698 (N_23698,N_23564,N_23469);
or U23699 (N_23699,N_23511,N_23528);
nor U23700 (N_23700,N_23436,N_23572);
nand U23701 (N_23701,N_23413,N_23503);
and U23702 (N_23702,N_23594,N_23404);
and U23703 (N_23703,N_23476,N_23558);
nor U23704 (N_23704,N_23559,N_23490);
nand U23705 (N_23705,N_23469,N_23407);
nand U23706 (N_23706,N_23461,N_23465);
and U23707 (N_23707,N_23449,N_23436);
and U23708 (N_23708,N_23461,N_23443);
or U23709 (N_23709,N_23539,N_23505);
nand U23710 (N_23710,N_23422,N_23453);
and U23711 (N_23711,N_23567,N_23422);
nor U23712 (N_23712,N_23470,N_23590);
nor U23713 (N_23713,N_23466,N_23471);
xor U23714 (N_23714,N_23543,N_23408);
nor U23715 (N_23715,N_23423,N_23589);
and U23716 (N_23716,N_23551,N_23427);
or U23717 (N_23717,N_23518,N_23581);
nand U23718 (N_23718,N_23476,N_23442);
xor U23719 (N_23719,N_23597,N_23563);
and U23720 (N_23720,N_23427,N_23490);
nand U23721 (N_23721,N_23504,N_23468);
and U23722 (N_23722,N_23567,N_23463);
nor U23723 (N_23723,N_23592,N_23466);
nand U23724 (N_23724,N_23539,N_23433);
xor U23725 (N_23725,N_23551,N_23521);
or U23726 (N_23726,N_23572,N_23575);
or U23727 (N_23727,N_23559,N_23548);
and U23728 (N_23728,N_23409,N_23495);
nand U23729 (N_23729,N_23586,N_23590);
nor U23730 (N_23730,N_23571,N_23584);
or U23731 (N_23731,N_23492,N_23578);
nor U23732 (N_23732,N_23547,N_23482);
or U23733 (N_23733,N_23503,N_23443);
nand U23734 (N_23734,N_23453,N_23420);
and U23735 (N_23735,N_23439,N_23547);
nor U23736 (N_23736,N_23563,N_23575);
nor U23737 (N_23737,N_23458,N_23400);
or U23738 (N_23738,N_23590,N_23428);
or U23739 (N_23739,N_23458,N_23485);
xor U23740 (N_23740,N_23498,N_23400);
and U23741 (N_23741,N_23432,N_23518);
nor U23742 (N_23742,N_23446,N_23478);
or U23743 (N_23743,N_23542,N_23562);
and U23744 (N_23744,N_23581,N_23596);
nor U23745 (N_23745,N_23417,N_23523);
or U23746 (N_23746,N_23573,N_23540);
or U23747 (N_23747,N_23494,N_23528);
xor U23748 (N_23748,N_23456,N_23578);
nand U23749 (N_23749,N_23437,N_23478);
and U23750 (N_23750,N_23535,N_23421);
xnor U23751 (N_23751,N_23592,N_23577);
or U23752 (N_23752,N_23401,N_23415);
nand U23753 (N_23753,N_23492,N_23579);
and U23754 (N_23754,N_23543,N_23493);
and U23755 (N_23755,N_23456,N_23522);
xor U23756 (N_23756,N_23571,N_23476);
nor U23757 (N_23757,N_23430,N_23545);
xnor U23758 (N_23758,N_23411,N_23410);
or U23759 (N_23759,N_23552,N_23539);
xnor U23760 (N_23760,N_23573,N_23478);
nand U23761 (N_23761,N_23436,N_23554);
or U23762 (N_23762,N_23410,N_23478);
nor U23763 (N_23763,N_23539,N_23465);
or U23764 (N_23764,N_23463,N_23473);
and U23765 (N_23765,N_23467,N_23500);
nor U23766 (N_23766,N_23541,N_23586);
and U23767 (N_23767,N_23526,N_23597);
xor U23768 (N_23768,N_23421,N_23426);
and U23769 (N_23769,N_23531,N_23474);
and U23770 (N_23770,N_23500,N_23424);
or U23771 (N_23771,N_23448,N_23568);
and U23772 (N_23772,N_23543,N_23462);
nor U23773 (N_23773,N_23596,N_23436);
nand U23774 (N_23774,N_23556,N_23503);
or U23775 (N_23775,N_23448,N_23554);
or U23776 (N_23776,N_23540,N_23519);
nor U23777 (N_23777,N_23466,N_23585);
nand U23778 (N_23778,N_23587,N_23588);
and U23779 (N_23779,N_23522,N_23544);
and U23780 (N_23780,N_23404,N_23438);
nor U23781 (N_23781,N_23449,N_23521);
xor U23782 (N_23782,N_23569,N_23494);
nand U23783 (N_23783,N_23523,N_23565);
nor U23784 (N_23784,N_23431,N_23541);
and U23785 (N_23785,N_23466,N_23492);
and U23786 (N_23786,N_23504,N_23535);
nor U23787 (N_23787,N_23526,N_23461);
nand U23788 (N_23788,N_23552,N_23522);
or U23789 (N_23789,N_23454,N_23459);
nor U23790 (N_23790,N_23566,N_23588);
and U23791 (N_23791,N_23498,N_23518);
or U23792 (N_23792,N_23543,N_23595);
xor U23793 (N_23793,N_23482,N_23410);
or U23794 (N_23794,N_23536,N_23470);
nor U23795 (N_23795,N_23424,N_23427);
and U23796 (N_23796,N_23517,N_23582);
xnor U23797 (N_23797,N_23595,N_23415);
or U23798 (N_23798,N_23493,N_23554);
or U23799 (N_23799,N_23552,N_23566);
nor U23800 (N_23800,N_23718,N_23620);
xor U23801 (N_23801,N_23613,N_23780);
xnor U23802 (N_23802,N_23666,N_23767);
and U23803 (N_23803,N_23657,N_23698);
or U23804 (N_23804,N_23717,N_23719);
nor U23805 (N_23805,N_23757,N_23798);
or U23806 (N_23806,N_23762,N_23749);
and U23807 (N_23807,N_23612,N_23754);
xor U23808 (N_23808,N_23652,N_23658);
and U23809 (N_23809,N_23634,N_23627);
or U23810 (N_23810,N_23624,N_23655);
or U23811 (N_23811,N_23761,N_23637);
xor U23812 (N_23812,N_23726,N_23660);
nor U23813 (N_23813,N_23677,N_23701);
nand U23814 (N_23814,N_23741,N_23667);
nor U23815 (N_23815,N_23645,N_23714);
and U23816 (N_23816,N_23723,N_23687);
nor U23817 (N_23817,N_23695,N_23676);
xnor U23818 (N_23818,N_23689,N_23720);
xnor U23819 (N_23819,N_23721,N_23686);
and U23820 (N_23820,N_23673,N_23632);
nor U23821 (N_23821,N_23748,N_23656);
or U23822 (N_23822,N_23693,N_23685);
and U23823 (N_23823,N_23646,N_23758);
xnor U23824 (N_23824,N_23630,N_23766);
or U23825 (N_23825,N_23788,N_23750);
or U23826 (N_23826,N_23653,N_23638);
xnor U23827 (N_23827,N_23648,N_23680);
or U23828 (N_23828,N_23752,N_23775);
and U23829 (N_23829,N_23765,N_23699);
nand U23830 (N_23830,N_23618,N_23705);
nand U23831 (N_23831,N_23784,N_23697);
xnor U23832 (N_23832,N_23796,N_23737);
xor U23833 (N_23833,N_23715,N_23614);
nand U23834 (N_23834,N_23755,N_23734);
or U23835 (N_23835,N_23616,N_23644);
nor U23836 (N_23836,N_23702,N_23746);
nor U23837 (N_23837,N_23662,N_23626);
nand U23838 (N_23838,N_23739,N_23759);
or U23839 (N_23839,N_23793,N_23777);
or U23840 (N_23840,N_23785,N_23782);
or U23841 (N_23841,N_23799,N_23610);
xnor U23842 (N_23842,N_23773,N_23747);
or U23843 (N_23843,N_23679,N_23684);
or U23844 (N_23844,N_23708,N_23724);
nor U23845 (N_23845,N_23743,N_23635);
nand U23846 (N_23846,N_23651,N_23760);
and U23847 (N_23847,N_23706,N_23642);
nor U23848 (N_23848,N_23732,N_23674);
nor U23849 (N_23849,N_23670,N_23795);
and U23850 (N_23850,N_23625,N_23738);
and U23851 (N_23851,N_23659,N_23727);
nor U23852 (N_23852,N_23690,N_23753);
nand U23853 (N_23853,N_23751,N_23731);
nor U23854 (N_23854,N_23682,N_23707);
nor U23855 (N_23855,N_23792,N_23769);
xor U23856 (N_23856,N_23602,N_23619);
nand U23857 (N_23857,N_23608,N_23694);
or U23858 (N_23858,N_23607,N_23641);
xor U23859 (N_23859,N_23604,N_23744);
or U23860 (N_23860,N_23688,N_23633);
xnor U23861 (N_23861,N_23671,N_23609);
or U23862 (N_23862,N_23764,N_23742);
or U23863 (N_23863,N_23763,N_23643);
or U23864 (N_23864,N_23647,N_23768);
nor U23865 (N_23865,N_23740,N_23663);
and U23866 (N_23866,N_23664,N_23735);
nor U23867 (N_23867,N_23611,N_23756);
or U23868 (N_23868,N_23640,N_23745);
xnor U23869 (N_23869,N_23700,N_23733);
or U23870 (N_23870,N_23683,N_23661);
or U23871 (N_23871,N_23730,N_23786);
and U23872 (N_23872,N_23696,N_23711);
nor U23873 (N_23873,N_23691,N_23791);
xnor U23874 (N_23874,N_23709,N_23728);
and U23875 (N_23875,N_23654,N_23675);
xor U23876 (N_23876,N_23629,N_23781);
and U23877 (N_23877,N_23600,N_23669);
and U23878 (N_23878,N_23649,N_23692);
nor U23879 (N_23879,N_23716,N_23621);
nand U23880 (N_23880,N_23665,N_23623);
or U23881 (N_23881,N_23797,N_23712);
xnor U23882 (N_23882,N_23704,N_23710);
and U23883 (N_23883,N_23789,N_23603);
xnor U23884 (N_23884,N_23771,N_23722);
nand U23885 (N_23885,N_23672,N_23770);
xnor U23886 (N_23886,N_23650,N_23778);
nor U23887 (N_23887,N_23729,N_23668);
or U23888 (N_23888,N_23622,N_23601);
and U23889 (N_23889,N_23628,N_23725);
nor U23890 (N_23890,N_23615,N_23779);
nand U23891 (N_23891,N_23631,N_23617);
xor U23892 (N_23892,N_23703,N_23776);
nand U23893 (N_23893,N_23636,N_23772);
or U23894 (N_23894,N_23678,N_23606);
nor U23895 (N_23895,N_23639,N_23605);
or U23896 (N_23896,N_23794,N_23713);
xnor U23897 (N_23897,N_23783,N_23681);
or U23898 (N_23898,N_23787,N_23736);
nand U23899 (N_23899,N_23774,N_23790);
and U23900 (N_23900,N_23776,N_23663);
nand U23901 (N_23901,N_23627,N_23753);
or U23902 (N_23902,N_23715,N_23752);
and U23903 (N_23903,N_23644,N_23763);
or U23904 (N_23904,N_23625,N_23621);
xor U23905 (N_23905,N_23733,N_23743);
and U23906 (N_23906,N_23727,N_23632);
xor U23907 (N_23907,N_23674,N_23796);
or U23908 (N_23908,N_23695,N_23613);
nand U23909 (N_23909,N_23713,N_23639);
or U23910 (N_23910,N_23796,N_23604);
nor U23911 (N_23911,N_23694,N_23626);
or U23912 (N_23912,N_23680,N_23637);
nand U23913 (N_23913,N_23647,N_23747);
or U23914 (N_23914,N_23735,N_23712);
nor U23915 (N_23915,N_23725,N_23627);
or U23916 (N_23916,N_23770,N_23752);
xor U23917 (N_23917,N_23743,N_23603);
xor U23918 (N_23918,N_23777,N_23623);
xor U23919 (N_23919,N_23615,N_23645);
nor U23920 (N_23920,N_23635,N_23750);
xnor U23921 (N_23921,N_23713,N_23702);
nand U23922 (N_23922,N_23793,N_23646);
and U23923 (N_23923,N_23616,N_23690);
xor U23924 (N_23924,N_23643,N_23754);
nand U23925 (N_23925,N_23744,N_23794);
and U23926 (N_23926,N_23693,N_23612);
nor U23927 (N_23927,N_23648,N_23781);
xnor U23928 (N_23928,N_23793,N_23665);
nor U23929 (N_23929,N_23621,N_23623);
nand U23930 (N_23930,N_23608,N_23722);
nand U23931 (N_23931,N_23634,N_23677);
xnor U23932 (N_23932,N_23711,N_23697);
nor U23933 (N_23933,N_23719,N_23750);
xor U23934 (N_23934,N_23727,N_23777);
xnor U23935 (N_23935,N_23692,N_23735);
xnor U23936 (N_23936,N_23760,N_23750);
and U23937 (N_23937,N_23755,N_23737);
nor U23938 (N_23938,N_23663,N_23639);
nand U23939 (N_23939,N_23700,N_23781);
nand U23940 (N_23940,N_23798,N_23726);
or U23941 (N_23941,N_23675,N_23649);
nand U23942 (N_23942,N_23787,N_23671);
or U23943 (N_23943,N_23601,N_23779);
nor U23944 (N_23944,N_23742,N_23607);
xnor U23945 (N_23945,N_23737,N_23742);
nor U23946 (N_23946,N_23693,N_23695);
and U23947 (N_23947,N_23759,N_23794);
or U23948 (N_23948,N_23663,N_23767);
and U23949 (N_23949,N_23728,N_23608);
nand U23950 (N_23950,N_23755,N_23780);
nor U23951 (N_23951,N_23748,N_23612);
and U23952 (N_23952,N_23758,N_23697);
and U23953 (N_23953,N_23640,N_23798);
xor U23954 (N_23954,N_23610,N_23789);
nand U23955 (N_23955,N_23706,N_23760);
nor U23956 (N_23956,N_23736,N_23721);
and U23957 (N_23957,N_23707,N_23638);
and U23958 (N_23958,N_23666,N_23788);
xnor U23959 (N_23959,N_23788,N_23699);
and U23960 (N_23960,N_23714,N_23692);
and U23961 (N_23961,N_23677,N_23600);
nand U23962 (N_23962,N_23749,N_23799);
nand U23963 (N_23963,N_23659,N_23799);
nor U23964 (N_23964,N_23706,N_23615);
nor U23965 (N_23965,N_23643,N_23629);
or U23966 (N_23966,N_23621,N_23604);
or U23967 (N_23967,N_23605,N_23650);
nor U23968 (N_23968,N_23785,N_23724);
and U23969 (N_23969,N_23607,N_23650);
nand U23970 (N_23970,N_23785,N_23753);
or U23971 (N_23971,N_23760,N_23780);
or U23972 (N_23972,N_23759,N_23738);
nor U23973 (N_23973,N_23730,N_23780);
xor U23974 (N_23974,N_23693,N_23650);
or U23975 (N_23975,N_23671,N_23764);
and U23976 (N_23976,N_23612,N_23631);
nand U23977 (N_23977,N_23704,N_23618);
and U23978 (N_23978,N_23628,N_23660);
nand U23979 (N_23979,N_23648,N_23796);
or U23980 (N_23980,N_23798,N_23674);
and U23981 (N_23981,N_23689,N_23658);
nor U23982 (N_23982,N_23604,N_23720);
xnor U23983 (N_23983,N_23609,N_23785);
xor U23984 (N_23984,N_23737,N_23678);
and U23985 (N_23985,N_23725,N_23624);
nand U23986 (N_23986,N_23614,N_23664);
nor U23987 (N_23987,N_23640,N_23669);
nand U23988 (N_23988,N_23628,N_23749);
nand U23989 (N_23989,N_23729,N_23769);
and U23990 (N_23990,N_23628,N_23658);
nor U23991 (N_23991,N_23677,N_23653);
and U23992 (N_23992,N_23672,N_23753);
or U23993 (N_23993,N_23735,N_23724);
or U23994 (N_23994,N_23601,N_23684);
xnor U23995 (N_23995,N_23706,N_23625);
nor U23996 (N_23996,N_23729,N_23605);
and U23997 (N_23997,N_23716,N_23624);
and U23998 (N_23998,N_23664,N_23657);
nor U23999 (N_23999,N_23697,N_23707);
xor U24000 (N_24000,N_23966,N_23917);
and U24001 (N_24001,N_23940,N_23856);
or U24002 (N_24002,N_23929,N_23840);
nor U24003 (N_24003,N_23896,N_23818);
nand U24004 (N_24004,N_23826,N_23993);
nand U24005 (N_24005,N_23845,N_23920);
or U24006 (N_24006,N_23982,N_23942);
nor U24007 (N_24007,N_23975,N_23863);
nor U24008 (N_24008,N_23974,N_23997);
xnor U24009 (N_24009,N_23860,N_23956);
and U24010 (N_24010,N_23830,N_23957);
xnor U24011 (N_24011,N_23871,N_23914);
nand U24012 (N_24012,N_23816,N_23802);
xor U24013 (N_24013,N_23904,N_23971);
xor U24014 (N_24014,N_23815,N_23877);
nand U24015 (N_24015,N_23883,N_23927);
nor U24016 (N_24016,N_23989,N_23949);
and U24017 (N_24017,N_23944,N_23908);
and U24018 (N_24018,N_23804,N_23855);
nor U24019 (N_24019,N_23801,N_23879);
or U24020 (N_24020,N_23808,N_23979);
or U24021 (N_24021,N_23918,N_23889);
xor U24022 (N_24022,N_23945,N_23867);
or U24023 (N_24023,N_23913,N_23948);
nor U24024 (N_24024,N_23968,N_23864);
xor U24025 (N_24025,N_23836,N_23960);
nand U24026 (N_24026,N_23911,N_23903);
and U24027 (N_24027,N_23839,N_23905);
or U24028 (N_24028,N_23881,N_23963);
and U24029 (N_24029,N_23819,N_23946);
nand U24030 (N_24030,N_23870,N_23842);
and U24031 (N_24031,N_23869,N_23961);
nor U24032 (N_24032,N_23866,N_23925);
nor U24033 (N_24033,N_23959,N_23928);
nand U24034 (N_24034,N_23894,N_23827);
nor U24035 (N_24035,N_23983,N_23841);
nor U24036 (N_24036,N_23969,N_23906);
xor U24037 (N_24037,N_23874,N_23831);
nor U24038 (N_24038,N_23807,N_23857);
or U24039 (N_24039,N_23932,N_23978);
nor U24040 (N_24040,N_23813,N_23843);
nand U24041 (N_24041,N_23909,N_23833);
xor U24042 (N_24042,N_23829,N_23977);
xnor U24043 (N_24043,N_23990,N_23844);
nand U24044 (N_24044,N_23964,N_23995);
and U24045 (N_24045,N_23919,N_23850);
xor U24046 (N_24046,N_23972,N_23885);
or U24047 (N_24047,N_23937,N_23882);
nand U24048 (N_24048,N_23976,N_23891);
nor U24049 (N_24049,N_23922,N_23910);
nor U24050 (N_24050,N_23846,N_23953);
or U24051 (N_24051,N_23888,N_23973);
and U24052 (N_24052,N_23876,N_23924);
xor U24053 (N_24053,N_23800,N_23951);
xor U24054 (N_24054,N_23921,N_23851);
and U24055 (N_24055,N_23861,N_23967);
or U24056 (N_24056,N_23886,N_23854);
xor U24057 (N_24057,N_23941,N_23998);
nor U24058 (N_24058,N_23992,N_23811);
xnor U24059 (N_24059,N_23915,N_23986);
xor U24060 (N_24060,N_23900,N_23892);
nor U24061 (N_24061,N_23952,N_23930);
xor U24062 (N_24062,N_23803,N_23858);
and U24063 (N_24063,N_23822,N_23933);
or U24064 (N_24064,N_23847,N_23890);
and U24065 (N_24065,N_23947,N_23878);
xnor U24066 (N_24066,N_23887,N_23884);
or U24067 (N_24067,N_23901,N_23981);
xnor U24068 (N_24068,N_23936,N_23824);
and U24069 (N_24069,N_23838,N_23849);
nor U24070 (N_24070,N_23825,N_23865);
xor U24071 (N_24071,N_23987,N_23821);
and U24072 (N_24072,N_23938,N_23996);
xor U24073 (N_24073,N_23958,N_23812);
xor U24074 (N_24074,N_23923,N_23814);
or U24075 (N_24075,N_23991,N_23943);
nor U24076 (N_24076,N_23809,N_23962);
nand U24077 (N_24077,N_23898,N_23994);
nand U24078 (N_24078,N_23985,N_23970);
xnor U24079 (N_24079,N_23931,N_23902);
and U24080 (N_24080,N_23848,N_23862);
and U24081 (N_24081,N_23873,N_23935);
nand U24082 (N_24082,N_23835,N_23868);
xnor U24083 (N_24083,N_23875,N_23988);
and U24084 (N_24084,N_23999,N_23893);
or U24085 (N_24085,N_23872,N_23950);
xor U24086 (N_24086,N_23817,N_23852);
nand U24087 (N_24087,N_23926,N_23810);
xor U24088 (N_24088,N_23820,N_23828);
nand U24089 (N_24089,N_23859,N_23837);
nand U24090 (N_24090,N_23895,N_23897);
xnor U24091 (N_24091,N_23912,N_23853);
nor U24092 (N_24092,N_23939,N_23832);
xor U24093 (N_24093,N_23907,N_23984);
xor U24094 (N_24094,N_23806,N_23916);
and U24095 (N_24095,N_23980,N_23954);
and U24096 (N_24096,N_23899,N_23805);
or U24097 (N_24097,N_23834,N_23965);
xnor U24098 (N_24098,N_23880,N_23823);
and U24099 (N_24099,N_23955,N_23934);
nand U24100 (N_24100,N_23907,N_23827);
and U24101 (N_24101,N_23923,N_23873);
or U24102 (N_24102,N_23954,N_23916);
nor U24103 (N_24103,N_23828,N_23836);
nor U24104 (N_24104,N_23877,N_23826);
xnor U24105 (N_24105,N_23989,N_23981);
and U24106 (N_24106,N_23870,N_23847);
xnor U24107 (N_24107,N_23913,N_23839);
nor U24108 (N_24108,N_23800,N_23845);
or U24109 (N_24109,N_23843,N_23828);
and U24110 (N_24110,N_23891,N_23857);
and U24111 (N_24111,N_23941,N_23816);
xnor U24112 (N_24112,N_23890,N_23820);
and U24113 (N_24113,N_23941,N_23842);
nor U24114 (N_24114,N_23940,N_23959);
or U24115 (N_24115,N_23853,N_23866);
and U24116 (N_24116,N_23851,N_23857);
nor U24117 (N_24117,N_23915,N_23844);
nor U24118 (N_24118,N_23842,N_23833);
xor U24119 (N_24119,N_23909,N_23805);
xor U24120 (N_24120,N_23910,N_23962);
and U24121 (N_24121,N_23940,N_23862);
nor U24122 (N_24122,N_23882,N_23978);
nand U24123 (N_24123,N_23932,N_23814);
and U24124 (N_24124,N_23912,N_23879);
nand U24125 (N_24125,N_23892,N_23803);
xnor U24126 (N_24126,N_23970,N_23913);
nor U24127 (N_24127,N_23962,N_23830);
and U24128 (N_24128,N_23881,N_23996);
nand U24129 (N_24129,N_23928,N_23993);
xor U24130 (N_24130,N_23976,N_23981);
xor U24131 (N_24131,N_23850,N_23989);
or U24132 (N_24132,N_23853,N_23872);
nor U24133 (N_24133,N_23938,N_23840);
or U24134 (N_24134,N_23954,N_23851);
xor U24135 (N_24135,N_23985,N_23801);
or U24136 (N_24136,N_23875,N_23952);
xor U24137 (N_24137,N_23847,N_23831);
and U24138 (N_24138,N_23935,N_23851);
xor U24139 (N_24139,N_23985,N_23849);
and U24140 (N_24140,N_23906,N_23909);
or U24141 (N_24141,N_23993,N_23930);
nand U24142 (N_24142,N_23977,N_23863);
nor U24143 (N_24143,N_23973,N_23843);
and U24144 (N_24144,N_23989,N_23841);
or U24145 (N_24145,N_23845,N_23947);
or U24146 (N_24146,N_23854,N_23966);
nor U24147 (N_24147,N_23978,N_23881);
or U24148 (N_24148,N_23863,N_23828);
or U24149 (N_24149,N_23845,N_23999);
or U24150 (N_24150,N_23972,N_23945);
and U24151 (N_24151,N_23924,N_23882);
xor U24152 (N_24152,N_23991,N_23844);
nor U24153 (N_24153,N_23919,N_23807);
nand U24154 (N_24154,N_23918,N_23827);
nand U24155 (N_24155,N_23831,N_23887);
or U24156 (N_24156,N_23877,N_23930);
nor U24157 (N_24157,N_23954,N_23929);
nor U24158 (N_24158,N_23985,N_23845);
nand U24159 (N_24159,N_23913,N_23925);
or U24160 (N_24160,N_23914,N_23806);
or U24161 (N_24161,N_23827,N_23974);
nand U24162 (N_24162,N_23864,N_23920);
xor U24163 (N_24163,N_23898,N_23910);
nor U24164 (N_24164,N_23896,N_23948);
nand U24165 (N_24165,N_23968,N_23875);
and U24166 (N_24166,N_23965,N_23895);
xnor U24167 (N_24167,N_23879,N_23993);
xnor U24168 (N_24168,N_23942,N_23804);
nand U24169 (N_24169,N_23845,N_23847);
or U24170 (N_24170,N_23880,N_23825);
nand U24171 (N_24171,N_23873,N_23979);
or U24172 (N_24172,N_23975,N_23924);
and U24173 (N_24173,N_23899,N_23944);
or U24174 (N_24174,N_23833,N_23965);
nand U24175 (N_24175,N_23956,N_23835);
xor U24176 (N_24176,N_23822,N_23852);
and U24177 (N_24177,N_23934,N_23999);
or U24178 (N_24178,N_23888,N_23930);
and U24179 (N_24179,N_23972,N_23863);
and U24180 (N_24180,N_23823,N_23958);
nor U24181 (N_24181,N_23994,N_23966);
xnor U24182 (N_24182,N_23976,N_23998);
xnor U24183 (N_24183,N_23853,N_23902);
xnor U24184 (N_24184,N_23983,N_23807);
or U24185 (N_24185,N_23984,N_23832);
or U24186 (N_24186,N_23930,N_23890);
and U24187 (N_24187,N_23941,N_23955);
nand U24188 (N_24188,N_23942,N_23805);
nor U24189 (N_24189,N_23964,N_23969);
or U24190 (N_24190,N_23866,N_23833);
or U24191 (N_24191,N_23929,N_23876);
and U24192 (N_24192,N_23943,N_23982);
nor U24193 (N_24193,N_23975,N_23861);
or U24194 (N_24194,N_23952,N_23845);
or U24195 (N_24195,N_23953,N_23870);
xnor U24196 (N_24196,N_23892,N_23854);
and U24197 (N_24197,N_23848,N_23953);
and U24198 (N_24198,N_23897,N_23977);
and U24199 (N_24199,N_23935,N_23949);
nand U24200 (N_24200,N_24183,N_24086);
and U24201 (N_24201,N_24006,N_24131);
or U24202 (N_24202,N_24096,N_24057);
nor U24203 (N_24203,N_24017,N_24124);
nor U24204 (N_24204,N_24071,N_24178);
nor U24205 (N_24205,N_24186,N_24104);
xnor U24206 (N_24206,N_24145,N_24164);
and U24207 (N_24207,N_24182,N_24043);
nand U24208 (N_24208,N_24160,N_24168);
xnor U24209 (N_24209,N_24013,N_24171);
xnor U24210 (N_24210,N_24002,N_24047);
or U24211 (N_24211,N_24022,N_24097);
or U24212 (N_24212,N_24115,N_24078);
nor U24213 (N_24213,N_24062,N_24197);
xor U24214 (N_24214,N_24005,N_24173);
xor U24215 (N_24215,N_24016,N_24158);
nand U24216 (N_24216,N_24014,N_24109);
xnor U24217 (N_24217,N_24166,N_24020);
nor U24218 (N_24218,N_24174,N_24147);
or U24219 (N_24219,N_24134,N_24095);
and U24220 (N_24220,N_24007,N_24105);
or U24221 (N_24221,N_24079,N_24117);
xnor U24222 (N_24222,N_24187,N_24179);
nor U24223 (N_24223,N_24037,N_24041);
or U24224 (N_24224,N_24159,N_24148);
nand U24225 (N_24225,N_24051,N_24100);
xor U24226 (N_24226,N_24108,N_24039);
nand U24227 (N_24227,N_24025,N_24198);
and U24228 (N_24228,N_24021,N_24075);
nor U24229 (N_24229,N_24107,N_24130);
xor U24230 (N_24230,N_24122,N_24093);
and U24231 (N_24231,N_24061,N_24012);
or U24232 (N_24232,N_24136,N_24082);
nand U24233 (N_24233,N_24127,N_24029);
nand U24234 (N_24234,N_24089,N_24137);
nand U24235 (N_24235,N_24118,N_24068);
and U24236 (N_24236,N_24045,N_24081);
xnor U24237 (N_24237,N_24150,N_24146);
and U24238 (N_24238,N_24060,N_24112);
xor U24239 (N_24239,N_24032,N_24190);
and U24240 (N_24240,N_24114,N_24170);
or U24241 (N_24241,N_24125,N_24181);
nand U24242 (N_24242,N_24073,N_24149);
nand U24243 (N_24243,N_24080,N_24035);
and U24244 (N_24244,N_24143,N_24034);
or U24245 (N_24245,N_24052,N_24087);
nand U24246 (N_24246,N_24092,N_24154);
nor U24247 (N_24247,N_24046,N_24055);
or U24248 (N_24248,N_24111,N_24050);
nand U24249 (N_24249,N_24138,N_24119);
and U24250 (N_24250,N_24157,N_24026);
and U24251 (N_24251,N_24053,N_24027);
xnor U24252 (N_24252,N_24008,N_24099);
xnor U24253 (N_24253,N_24036,N_24167);
or U24254 (N_24254,N_24191,N_24165);
or U24255 (N_24255,N_24001,N_24058);
nor U24256 (N_24256,N_24193,N_24188);
nand U24257 (N_24257,N_24175,N_24024);
nand U24258 (N_24258,N_24072,N_24196);
nand U24259 (N_24259,N_24121,N_24155);
xor U24260 (N_24260,N_24019,N_24110);
and U24261 (N_24261,N_24177,N_24044);
xor U24262 (N_24262,N_24015,N_24056);
and U24263 (N_24263,N_24169,N_24031);
nor U24264 (N_24264,N_24028,N_24059);
or U24265 (N_24265,N_24133,N_24054);
nor U24266 (N_24266,N_24033,N_24199);
nand U24267 (N_24267,N_24064,N_24069);
nand U24268 (N_24268,N_24066,N_24084);
or U24269 (N_24269,N_24085,N_24048);
xor U24270 (N_24270,N_24094,N_24113);
nor U24271 (N_24271,N_24194,N_24088);
and U24272 (N_24272,N_24153,N_24156);
nor U24273 (N_24273,N_24018,N_24101);
and U24274 (N_24274,N_24152,N_24009);
and U24275 (N_24275,N_24102,N_24038);
nor U24276 (N_24276,N_24184,N_24195);
nand U24277 (N_24277,N_24070,N_24049);
and U24278 (N_24278,N_24163,N_24139);
nand U24279 (N_24279,N_24128,N_24192);
xor U24280 (N_24280,N_24140,N_24011);
nor U24281 (N_24281,N_24116,N_24142);
and U24282 (N_24282,N_24074,N_24185);
or U24283 (N_24283,N_24000,N_24023);
or U24284 (N_24284,N_24103,N_24151);
xnor U24285 (N_24285,N_24063,N_24189);
or U24286 (N_24286,N_24132,N_24120);
nor U24287 (N_24287,N_24126,N_24040);
nor U24288 (N_24288,N_24091,N_24161);
xnor U24289 (N_24289,N_24004,N_24172);
nor U24290 (N_24290,N_24076,N_24010);
xnor U24291 (N_24291,N_24098,N_24090);
nor U24292 (N_24292,N_24129,N_24135);
and U24293 (N_24293,N_24030,N_24083);
and U24294 (N_24294,N_24176,N_24180);
or U24295 (N_24295,N_24106,N_24042);
nand U24296 (N_24296,N_24003,N_24067);
nor U24297 (N_24297,N_24077,N_24141);
or U24298 (N_24298,N_24144,N_24162);
or U24299 (N_24299,N_24123,N_24065);
and U24300 (N_24300,N_24116,N_24062);
xnor U24301 (N_24301,N_24177,N_24036);
and U24302 (N_24302,N_24183,N_24029);
nor U24303 (N_24303,N_24188,N_24089);
nor U24304 (N_24304,N_24123,N_24012);
nor U24305 (N_24305,N_24063,N_24066);
and U24306 (N_24306,N_24091,N_24187);
or U24307 (N_24307,N_24005,N_24010);
and U24308 (N_24308,N_24175,N_24063);
xor U24309 (N_24309,N_24145,N_24126);
nor U24310 (N_24310,N_24052,N_24083);
nor U24311 (N_24311,N_24194,N_24030);
xor U24312 (N_24312,N_24014,N_24153);
nor U24313 (N_24313,N_24044,N_24170);
and U24314 (N_24314,N_24102,N_24143);
or U24315 (N_24315,N_24014,N_24069);
nor U24316 (N_24316,N_24025,N_24004);
and U24317 (N_24317,N_24029,N_24194);
nor U24318 (N_24318,N_24071,N_24081);
xor U24319 (N_24319,N_24180,N_24068);
and U24320 (N_24320,N_24087,N_24155);
xnor U24321 (N_24321,N_24133,N_24089);
or U24322 (N_24322,N_24130,N_24175);
or U24323 (N_24323,N_24106,N_24181);
or U24324 (N_24324,N_24090,N_24119);
or U24325 (N_24325,N_24102,N_24105);
nor U24326 (N_24326,N_24087,N_24006);
and U24327 (N_24327,N_24157,N_24151);
nand U24328 (N_24328,N_24090,N_24113);
and U24329 (N_24329,N_24025,N_24117);
nor U24330 (N_24330,N_24073,N_24187);
and U24331 (N_24331,N_24054,N_24170);
xnor U24332 (N_24332,N_24100,N_24096);
and U24333 (N_24333,N_24112,N_24010);
or U24334 (N_24334,N_24196,N_24145);
xor U24335 (N_24335,N_24050,N_24009);
xor U24336 (N_24336,N_24147,N_24149);
or U24337 (N_24337,N_24169,N_24123);
nand U24338 (N_24338,N_24104,N_24029);
nor U24339 (N_24339,N_24113,N_24134);
xnor U24340 (N_24340,N_24031,N_24102);
and U24341 (N_24341,N_24121,N_24154);
nand U24342 (N_24342,N_24172,N_24129);
xnor U24343 (N_24343,N_24034,N_24106);
or U24344 (N_24344,N_24060,N_24169);
xnor U24345 (N_24345,N_24197,N_24156);
nand U24346 (N_24346,N_24103,N_24017);
or U24347 (N_24347,N_24195,N_24053);
nand U24348 (N_24348,N_24185,N_24154);
and U24349 (N_24349,N_24046,N_24038);
nor U24350 (N_24350,N_24045,N_24152);
or U24351 (N_24351,N_24122,N_24140);
nor U24352 (N_24352,N_24170,N_24187);
or U24353 (N_24353,N_24069,N_24053);
nand U24354 (N_24354,N_24072,N_24085);
xor U24355 (N_24355,N_24126,N_24070);
nor U24356 (N_24356,N_24020,N_24162);
xor U24357 (N_24357,N_24172,N_24006);
and U24358 (N_24358,N_24117,N_24099);
nand U24359 (N_24359,N_24107,N_24168);
xnor U24360 (N_24360,N_24084,N_24196);
nor U24361 (N_24361,N_24053,N_24160);
or U24362 (N_24362,N_24167,N_24021);
nand U24363 (N_24363,N_24163,N_24029);
nor U24364 (N_24364,N_24056,N_24158);
nor U24365 (N_24365,N_24106,N_24060);
xor U24366 (N_24366,N_24038,N_24024);
or U24367 (N_24367,N_24196,N_24108);
xor U24368 (N_24368,N_24179,N_24006);
nor U24369 (N_24369,N_24108,N_24193);
or U24370 (N_24370,N_24175,N_24102);
and U24371 (N_24371,N_24091,N_24090);
or U24372 (N_24372,N_24183,N_24199);
xnor U24373 (N_24373,N_24102,N_24101);
and U24374 (N_24374,N_24055,N_24156);
xor U24375 (N_24375,N_24078,N_24062);
and U24376 (N_24376,N_24052,N_24165);
nand U24377 (N_24377,N_24054,N_24106);
xor U24378 (N_24378,N_24054,N_24188);
or U24379 (N_24379,N_24008,N_24174);
xnor U24380 (N_24380,N_24084,N_24077);
and U24381 (N_24381,N_24145,N_24104);
or U24382 (N_24382,N_24053,N_24117);
nor U24383 (N_24383,N_24152,N_24148);
and U24384 (N_24384,N_24038,N_24151);
nand U24385 (N_24385,N_24160,N_24057);
nand U24386 (N_24386,N_24058,N_24164);
nor U24387 (N_24387,N_24159,N_24136);
xor U24388 (N_24388,N_24030,N_24036);
nand U24389 (N_24389,N_24169,N_24057);
xor U24390 (N_24390,N_24198,N_24006);
nand U24391 (N_24391,N_24140,N_24095);
nor U24392 (N_24392,N_24021,N_24120);
nand U24393 (N_24393,N_24057,N_24146);
or U24394 (N_24394,N_24005,N_24034);
nor U24395 (N_24395,N_24136,N_24030);
nand U24396 (N_24396,N_24039,N_24075);
nand U24397 (N_24397,N_24030,N_24162);
xor U24398 (N_24398,N_24166,N_24051);
xnor U24399 (N_24399,N_24124,N_24098);
nand U24400 (N_24400,N_24204,N_24384);
nor U24401 (N_24401,N_24219,N_24383);
nand U24402 (N_24402,N_24304,N_24207);
and U24403 (N_24403,N_24330,N_24392);
xor U24404 (N_24404,N_24296,N_24336);
nor U24405 (N_24405,N_24310,N_24297);
or U24406 (N_24406,N_24231,N_24335);
nand U24407 (N_24407,N_24294,N_24273);
nor U24408 (N_24408,N_24390,N_24205);
nor U24409 (N_24409,N_24361,N_24343);
or U24410 (N_24410,N_24292,N_24394);
nand U24411 (N_24411,N_24378,N_24222);
and U24412 (N_24412,N_24397,N_24291);
and U24413 (N_24413,N_24346,N_24278);
or U24414 (N_24414,N_24260,N_24389);
nor U24415 (N_24415,N_24360,N_24327);
nor U24416 (N_24416,N_24325,N_24253);
nand U24417 (N_24417,N_24313,N_24312);
or U24418 (N_24418,N_24283,N_24276);
nor U24419 (N_24419,N_24328,N_24270);
nand U24420 (N_24420,N_24373,N_24263);
xor U24421 (N_24421,N_24299,N_24208);
and U24422 (N_24422,N_24215,N_24357);
nand U24423 (N_24423,N_24301,N_24201);
nand U24424 (N_24424,N_24286,N_24329);
nor U24425 (N_24425,N_24355,N_24240);
and U24426 (N_24426,N_24254,N_24369);
and U24427 (N_24427,N_24305,N_24290);
or U24428 (N_24428,N_24332,N_24348);
nor U24429 (N_24429,N_24224,N_24344);
and U24430 (N_24430,N_24381,N_24251);
xor U24431 (N_24431,N_24236,N_24368);
nor U24432 (N_24432,N_24250,N_24352);
xor U24433 (N_24433,N_24298,N_24238);
nand U24434 (N_24434,N_24351,N_24206);
xnor U24435 (N_24435,N_24387,N_24303);
nor U24436 (N_24436,N_24309,N_24244);
xor U24437 (N_24437,N_24265,N_24264);
or U24438 (N_24438,N_24277,N_24233);
nor U24439 (N_24439,N_24248,N_24306);
nand U24440 (N_24440,N_24372,N_24293);
and U24441 (N_24441,N_24356,N_24225);
xnor U24442 (N_24442,N_24308,N_24223);
xnor U24443 (N_24443,N_24345,N_24243);
and U24444 (N_24444,N_24227,N_24320);
nand U24445 (N_24445,N_24342,N_24229);
and U24446 (N_24446,N_24377,N_24334);
nor U24447 (N_24447,N_24282,N_24235);
nand U24448 (N_24448,N_24341,N_24275);
nor U24449 (N_24449,N_24274,N_24375);
nor U24450 (N_24450,N_24364,N_24212);
nor U24451 (N_24451,N_24391,N_24242);
and U24452 (N_24452,N_24359,N_24380);
or U24453 (N_24453,N_24363,N_24272);
and U24454 (N_24454,N_24221,N_24281);
or U24455 (N_24455,N_24210,N_24367);
or U24456 (N_24456,N_24268,N_24202);
xor U24457 (N_24457,N_24370,N_24241);
or U24458 (N_24458,N_24262,N_24258);
or U24459 (N_24459,N_24230,N_24388);
nand U24460 (N_24460,N_24339,N_24333);
nand U24461 (N_24461,N_24379,N_24209);
nor U24462 (N_24462,N_24289,N_24358);
or U24463 (N_24463,N_24216,N_24256);
and U24464 (N_24464,N_24213,N_24228);
nor U24465 (N_24465,N_24217,N_24319);
nand U24466 (N_24466,N_24261,N_24393);
and U24467 (N_24467,N_24318,N_24316);
and U24468 (N_24468,N_24331,N_24324);
or U24469 (N_24469,N_24317,N_24396);
or U24470 (N_24470,N_24245,N_24323);
and U24471 (N_24471,N_24371,N_24218);
or U24472 (N_24472,N_24302,N_24314);
xor U24473 (N_24473,N_24259,N_24295);
nand U24474 (N_24474,N_24280,N_24326);
xor U24475 (N_24475,N_24214,N_24252);
nor U24476 (N_24476,N_24321,N_24288);
and U24477 (N_24477,N_24285,N_24255);
nand U24478 (N_24478,N_24382,N_24311);
nor U24479 (N_24479,N_24365,N_24200);
nand U24480 (N_24480,N_24232,N_24362);
nand U24481 (N_24481,N_24300,N_24239);
and U24482 (N_24482,N_24386,N_24220);
xnor U24483 (N_24483,N_24246,N_24385);
and U24484 (N_24484,N_24398,N_24211);
or U24485 (N_24485,N_24234,N_24249);
and U24486 (N_24486,N_24340,N_24353);
and U24487 (N_24487,N_24284,N_24337);
nor U24488 (N_24488,N_24399,N_24366);
or U24489 (N_24489,N_24203,N_24322);
nand U24490 (N_24490,N_24354,N_24395);
nor U24491 (N_24491,N_24226,N_24349);
xnor U24492 (N_24492,N_24237,N_24338);
or U24493 (N_24493,N_24269,N_24267);
xor U24494 (N_24494,N_24247,N_24350);
and U24495 (N_24495,N_24279,N_24315);
nand U24496 (N_24496,N_24257,N_24374);
nand U24497 (N_24497,N_24307,N_24347);
nand U24498 (N_24498,N_24376,N_24271);
xnor U24499 (N_24499,N_24266,N_24287);
and U24500 (N_24500,N_24268,N_24367);
and U24501 (N_24501,N_24300,N_24233);
or U24502 (N_24502,N_24293,N_24248);
nor U24503 (N_24503,N_24214,N_24289);
xnor U24504 (N_24504,N_24261,N_24251);
nand U24505 (N_24505,N_24252,N_24242);
or U24506 (N_24506,N_24374,N_24384);
nand U24507 (N_24507,N_24393,N_24270);
and U24508 (N_24508,N_24373,N_24253);
nor U24509 (N_24509,N_24280,N_24214);
and U24510 (N_24510,N_24358,N_24227);
and U24511 (N_24511,N_24324,N_24273);
or U24512 (N_24512,N_24307,N_24234);
or U24513 (N_24513,N_24307,N_24348);
nand U24514 (N_24514,N_24394,N_24399);
nand U24515 (N_24515,N_24380,N_24287);
nor U24516 (N_24516,N_24255,N_24262);
or U24517 (N_24517,N_24237,N_24319);
xor U24518 (N_24518,N_24203,N_24321);
or U24519 (N_24519,N_24238,N_24338);
or U24520 (N_24520,N_24383,N_24397);
xor U24521 (N_24521,N_24230,N_24221);
and U24522 (N_24522,N_24236,N_24252);
or U24523 (N_24523,N_24318,N_24278);
or U24524 (N_24524,N_24376,N_24296);
nor U24525 (N_24525,N_24225,N_24283);
nand U24526 (N_24526,N_24264,N_24289);
nand U24527 (N_24527,N_24336,N_24347);
or U24528 (N_24528,N_24223,N_24215);
nand U24529 (N_24529,N_24274,N_24325);
nand U24530 (N_24530,N_24398,N_24324);
xor U24531 (N_24531,N_24279,N_24291);
and U24532 (N_24532,N_24378,N_24391);
or U24533 (N_24533,N_24261,N_24284);
nand U24534 (N_24534,N_24225,N_24355);
nand U24535 (N_24535,N_24352,N_24328);
and U24536 (N_24536,N_24378,N_24232);
and U24537 (N_24537,N_24274,N_24286);
xnor U24538 (N_24538,N_24271,N_24205);
nor U24539 (N_24539,N_24308,N_24217);
xor U24540 (N_24540,N_24283,N_24311);
or U24541 (N_24541,N_24242,N_24208);
nand U24542 (N_24542,N_24291,N_24259);
and U24543 (N_24543,N_24320,N_24389);
nor U24544 (N_24544,N_24204,N_24244);
and U24545 (N_24545,N_24304,N_24289);
or U24546 (N_24546,N_24279,N_24203);
and U24547 (N_24547,N_24374,N_24327);
or U24548 (N_24548,N_24264,N_24247);
nand U24549 (N_24549,N_24329,N_24226);
xor U24550 (N_24550,N_24277,N_24322);
and U24551 (N_24551,N_24266,N_24261);
nand U24552 (N_24552,N_24393,N_24236);
xor U24553 (N_24553,N_24213,N_24298);
nor U24554 (N_24554,N_24221,N_24328);
nand U24555 (N_24555,N_24388,N_24337);
nor U24556 (N_24556,N_24244,N_24209);
and U24557 (N_24557,N_24281,N_24271);
xor U24558 (N_24558,N_24252,N_24306);
xnor U24559 (N_24559,N_24241,N_24201);
and U24560 (N_24560,N_24271,N_24307);
or U24561 (N_24561,N_24221,N_24241);
xor U24562 (N_24562,N_24295,N_24398);
nand U24563 (N_24563,N_24243,N_24247);
nor U24564 (N_24564,N_24348,N_24317);
or U24565 (N_24565,N_24205,N_24399);
and U24566 (N_24566,N_24345,N_24254);
xnor U24567 (N_24567,N_24334,N_24326);
or U24568 (N_24568,N_24321,N_24280);
and U24569 (N_24569,N_24229,N_24367);
or U24570 (N_24570,N_24282,N_24353);
or U24571 (N_24571,N_24323,N_24266);
nand U24572 (N_24572,N_24296,N_24317);
and U24573 (N_24573,N_24245,N_24276);
nand U24574 (N_24574,N_24304,N_24233);
nor U24575 (N_24575,N_24295,N_24355);
nor U24576 (N_24576,N_24343,N_24209);
nor U24577 (N_24577,N_24301,N_24296);
xnor U24578 (N_24578,N_24394,N_24216);
xor U24579 (N_24579,N_24208,N_24336);
nor U24580 (N_24580,N_24246,N_24268);
or U24581 (N_24581,N_24231,N_24360);
and U24582 (N_24582,N_24381,N_24274);
nand U24583 (N_24583,N_24291,N_24245);
nor U24584 (N_24584,N_24346,N_24301);
nor U24585 (N_24585,N_24278,N_24380);
nand U24586 (N_24586,N_24397,N_24307);
and U24587 (N_24587,N_24372,N_24307);
xor U24588 (N_24588,N_24359,N_24321);
xnor U24589 (N_24589,N_24278,N_24273);
nand U24590 (N_24590,N_24255,N_24235);
nor U24591 (N_24591,N_24384,N_24289);
nor U24592 (N_24592,N_24234,N_24295);
xnor U24593 (N_24593,N_24250,N_24327);
nor U24594 (N_24594,N_24322,N_24215);
and U24595 (N_24595,N_24331,N_24257);
and U24596 (N_24596,N_24312,N_24297);
nand U24597 (N_24597,N_24374,N_24376);
nor U24598 (N_24598,N_24368,N_24246);
xnor U24599 (N_24599,N_24299,N_24325);
and U24600 (N_24600,N_24475,N_24466);
or U24601 (N_24601,N_24402,N_24497);
nor U24602 (N_24602,N_24429,N_24517);
xor U24603 (N_24603,N_24558,N_24538);
nor U24604 (N_24604,N_24505,N_24559);
and U24605 (N_24605,N_24582,N_24536);
or U24606 (N_24606,N_24504,N_24455);
or U24607 (N_24607,N_24498,N_24562);
or U24608 (N_24608,N_24526,N_24436);
nor U24609 (N_24609,N_24550,N_24572);
nor U24610 (N_24610,N_24537,N_24420);
xnor U24611 (N_24611,N_24564,N_24452);
xor U24612 (N_24612,N_24431,N_24584);
and U24613 (N_24613,N_24464,N_24408);
nand U24614 (N_24614,N_24440,N_24503);
nor U24615 (N_24615,N_24579,N_24568);
xor U24616 (N_24616,N_24400,N_24456);
or U24617 (N_24617,N_24424,N_24423);
nand U24618 (N_24618,N_24404,N_24591);
xor U24619 (N_24619,N_24439,N_24478);
nand U24620 (N_24620,N_24560,N_24535);
and U24621 (N_24621,N_24586,N_24547);
nor U24622 (N_24622,N_24576,N_24570);
nor U24623 (N_24623,N_24453,N_24565);
nand U24624 (N_24624,N_24414,N_24409);
nor U24625 (N_24625,N_24418,N_24575);
and U24626 (N_24626,N_24479,N_24494);
or U24627 (N_24627,N_24460,N_24415);
and U24628 (N_24628,N_24461,N_24527);
and U24629 (N_24629,N_24519,N_24444);
and U24630 (N_24630,N_24510,N_24549);
and U24631 (N_24631,N_24502,N_24412);
nor U24632 (N_24632,N_24506,N_24462);
xnor U24633 (N_24633,N_24546,N_24442);
xor U24634 (N_24634,N_24445,N_24581);
or U24635 (N_24635,N_24594,N_24512);
or U24636 (N_24636,N_24515,N_24544);
nor U24637 (N_24637,N_24525,N_24446);
or U24638 (N_24638,N_24499,N_24493);
nor U24639 (N_24639,N_24441,N_24428);
nor U24640 (N_24640,N_24553,N_24542);
xor U24641 (N_24641,N_24573,N_24589);
xor U24642 (N_24642,N_24548,N_24580);
nand U24643 (N_24643,N_24435,N_24477);
and U24644 (N_24644,N_24492,N_24458);
nand U24645 (N_24645,N_24486,N_24578);
nand U24646 (N_24646,N_24407,N_24567);
and U24647 (N_24647,N_24593,N_24432);
and U24648 (N_24648,N_24511,N_24545);
nor U24649 (N_24649,N_24513,N_24596);
and U24650 (N_24650,N_24474,N_24532);
nor U24651 (N_24651,N_24543,N_24590);
nand U24652 (N_24652,N_24557,N_24422);
or U24653 (N_24653,N_24469,N_24595);
nand U24654 (N_24654,N_24433,N_24416);
and U24655 (N_24655,N_24410,N_24419);
and U24656 (N_24656,N_24574,N_24483);
or U24657 (N_24657,N_24533,N_24495);
nor U24658 (N_24658,N_24468,N_24588);
xnor U24659 (N_24659,N_24489,N_24447);
nand U24660 (N_24660,N_24470,N_24585);
or U24661 (N_24661,N_24500,N_24430);
xnor U24662 (N_24662,N_24531,N_24514);
nor U24663 (N_24663,N_24485,N_24472);
nand U24664 (N_24664,N_24426,N_24599);
or U24665 (N_24665,N_24443,N_24507);
nor U24666 (N_24666,N_24484,N_24411);
nand U24667 (N_24667,N_24501,N_24561);
xor U24668 (N_24668,N_24521,N_24571);
and U24669 (N_24669,N_24516,N_24437);
xnor U24670 (N_24670,N_24450,N_24598);
and U24671 (N_24671,N_24438,N_24480);
and U24672 (N_24672,N_24551,N_24496);
nor U24673 (N_24673,N_24597,N_24459);
nand U24674 (N_24674,N_24569,N_24471);
nor U24675 (N_24675,N_24530,N_24522);
and U24676 (N_24676,N_24434,N_24481);
and U24677 (N_24677,N_24413,N_24583);
xor U24678 (N_24678,N_24491,N_24528);
or U24679 (N_24679,N_24509,N_24563);
nor U24680 (N_24680,N_24427,N_24473);
xnor U24681 (N_24681,N_24555,N_24592);
xor U24682 (N_24682,N_24482,N_24540);
nand U24683 (N_24683,N_24508,N_24539);
xnor U24684 (N_24684,N_24587,N_24577);
xor U24685 (N_24685,N_24523,N_24401);
xor U24686 (N_24686,N_24465,N_24554);
xnor U24687 (N_24687,N_24524,N_24534);
and U24688 (N_24688,N_24425,N_24490);
xnor U24689 (N_24689,N_24488,N_24457);
xnor U24690 (N_24690,N_24518,N_24406);
and U24691 (N_24691,N_24556,N_24529);
or U24692 (N_24692,N_24566,N_24541);
nor U24693 (N_24693,N_24405,N_24487);
nand U24694 (N_24694,N_24467,N_24449);
xnor U24695 (N_24695,N_24520,N_24421);
and U24696 (N_24696,N_24552,N_24454);
xor U24697 (N_24697,N_24476,N_24403);
nor U24698 (N_24698,N_24417,N_24451);
and U24699 (N_24699,N_24463,N_24448);
nand U24700 (N_24700,N_24490,N_24555);
or U24701 (N_24701,N_24508,N_24543);
nand U24702 (N_24702,N_24535,N_24596);
nor U24703 (N_24703,N_24562,N_24420);
or U24704 (N_24704,N_24422,N_24451);
or U24705 (N_24705,N_24511,N_24430);
or U24706 (N_24706,N_24567,N_24476);
or U24707 (N_24707,N_24429,N_24528);
nor U24708 (N_24708,N_24486,N_24461);
nor U24709 (N_24709,N_24406,N_24497);
or U24710 (N_24710,N_24534,N_24547);
nor U24711 (N_24711,N_24583,N_24415);
nand U24712 (N_24712,N_24474,N_24454);
xnor U24713 (N_24713,N_24584,N_24550);
nand U24714 (N_24714,N_24541,N_24463);
or U24715 (N_24715,N_24511,N_24548);
nor U24716 (N_24716,N_24503,N_24579);
or U24717 (N_24717,N_24449,N_24411);
nor U24718 (N_24718,N_24472,N_24400);
and U24719 (N_24719,N_24564,N_24595);
nor U24720 (N_24720,N_24579,N_24432);
xor U24721 (N_24721,N_24543,N_24452);
nand U24722 (N_24722,N_24563,N_24590);
nor U24723 (N_24723,N_24550,N_24412);
and U24724 (N_24724,N_24432,N_24522);
xor U24725 (N_24725,N_24438,N_24553);
xor U24726 (N_24726,N_24543,N_24572);
xor U24727 (N_24727,N_24444,N_24427);
nand U24728 (N_24728,N_24483,N_24589);
nand U24729 (N_24729,N_24527,N_24424);
nor U24730 (N_24730,N_24523,N_24562);
or U24731 (N_24731,N_24405,N_24435);
or U24732 (N_24732,N_24458,N_24585);
and U24733 (N_24733,N_24578,N_24547);
or U24734 (N_24734,N_24565,N_24521);
and U24735 (N_24735,N_24438,N_24520);
and U24736 (N_24736,N_24557,N_24525);
nand U24737 (N_24737,N_24465,N_24415);
and U24738 (N_24738,N_24599,N_24457);
nand U24739 (N_24739,N_24581,N_24572);
and U24740 (N_24740,N_24485,N_24502);
nor U24741 (N_24741,N_24458,N_24531);
xor U24742 (N_24742,N_24447,N_24532);
and U24743 (N_24743,N_24543,N_24489);
and U24744 (N_24744,N_24414,N_24469);
or U24745 (N_24745,N_24502,N_24562);
or U24746 (N_24746,N_24530,N_24427);
nand U24747 (N_24747,N_24512,N_24502);
xnor U24748 (N_24748,N_24409,N_24504);
or U24749 (N_24749,N_24428,N_24518);
and U24750 (N_24750,N_24574,N_24556);
or U24751 (N_24751,N_24468,N_24444);
nor U24752 (N_24752,N_24581,N_24405);
xor U24753 (N_24753,N_24508,N_24567);
nor U24754 (N_24754,N_24439,N_24420);
xor U24755 (N_24755,N_24565,N_24463);
xnor U24756 (N_24756,N_24419,N_24529);
and U24757 (N_24757,N_24512,N_24415);
nor U24758 (N_24758,N_24420,N_24584);
and U24759 (N_24759,N_24531,N_24579);
or U24760 (N_24760,N_24518,N_24407);
nor U24761 (N_24761,N_24465,N_24461);
nor U24762 (N_24762,N_24533,N_24584);
xnor U24763 (N_24763,N_24541,N_24591);
nand U24764 (N_24764,N_24590,N_24514);
nand U24765 (N_24765,N_24453,N_24468);
or U24766 (N_24766,N_24594,N_24518);
nand U24767 (N_24767,N_24407,N_24419);
and U24768 (N_24768,N_24453,N_24452);
nand U24769 (N_24769,N_24499,N_24490);
nand U24770 (N_24770,N_24544,N_24537);
or U24771 (N_24771,N_24401,N_24511);
nand U24772 (N_24772,N_24520,N_24521);
nor U24773 (N_24773,N_24502,N_24407);
or U24774 (N_24774,N_24582,N_24515);
and U24775 (N_24775,N_24469,N_24486);
nor U24776 (N_24776,N_24580,N_24414);
xnor U24777 (N_24777,N_24486,N_24431);
nand U24778 (N_24778,N_24527,N_24449);
and U24779 (N_24779,N_24541,N_24430);
xnor U24780 (N_24780,N_24454,N_24456);
xor U24781 (N_24781,N_24436,N_24568);
nor U24782 (N_24782,N_24565,N_24408);
nor U24783 (N_24783,N_24545,N_24460);
or U24784 (N_24784,N_24450,N_24578);
or U24785 (N_24785,N_24450,N_24465);
xnor U24786 (N_24786,N_24589,N_24598);
and U24787 (N_24787,N_24577,N_24409);
nand U24788 (N_24788,N_24505,N_24549);
xor U24789 (N_24789,N_24592,N_24581);
xnor U24790 (N_24790,N_24444,N_24584);
and U24791 (N_24791,N_24516,N_24582);
nor U24792 (N_24792,N_24574,N_24462);
or U24793 (N_24793,N_24462,N_24566);
or U24794 (N_24794,N_24598,N_24543);
nor U24795 (N_24795,N_24537,N_24448);
or U24796 (N_24796,N_24465,N_24400);
xor U24797 (N_24797,N_24486,N_24562);
or U24798 (N_24798,N_24585,N_24426);
nor U24799 (N_24799,N_24485,N_24597);
nor U24800 (N_24800,N_24788,N_24752);
or U24801 (N_24801,N_24651,N_24789);
and U24802 (N_24802,N_24775,N_24658);
xor U24803 (N_24803,N_24680,N_24707);
nand U24804 (N_24804,N_24674,N_24758);
or U24805 (N_24805,N_24636,N_24696);
xor U24806 (N_24806,N_24777,N_24664);
xor U24807 (N_24807,N_24672,N_24670);
xor U24808 (N_24808,N_24647,N_24695);
and U24809 (N_24809,N_24710,N_24717);
xnor U24810 (N_24810,N_24702,N_24605);
nand U24811 (N_24811,N_24759,N_24669);
xnor U24812 (N_24812,N_24730,N_24621);
nor U24813 (N_24813,N_24635,N_24741);
nor U24814 (N_24814,N_24629,N_24649);
xor U24815 (N_24815,N_24754,N_24798);
nand U24816 (N_24816,N_24682,N_24746);
and U24817 (N_24817,N_24609,N_24760);
xor U24818 (N_24818,N_24701,N_24653);
or U24819 (N_24819,N_24604,N_24665);
and U24820 (N_24820,N_24633,N_24632);
and U24821 (N_24821,N_24634,N_24638);
nand U24822 (N_24822,N_24761,N_24771);
nand U24823 (N_24823,N_24666,N_24763);
nand U24824 (N_24824,N_24697,N_24673);
xor U24825 (N_24825,N_24641,N_24768);
and U24826 (N_24826,N_24753,N_24713);
xor U24827 (N_24827,N_24755,N_24659);
or U24828 (N_24828,N_24620,N_24765);
or U24829 (N_24829,N_24679,N_24602);
and U24830 (N_24830,N_24721,N_24607);
nand U24831 (N_24831,N_24734,N_24684);
and U24832 (N_24832,N_24625,N_24631);
nand U24833 (N_24833,N_24729,N_24790);
and U24834 (N_24834,N_24643,N_24736);
nand U24835 (N_24835,N_24750,N_24694);
nor U24836 (N_24836,N_24691,N_24622);
xnor U24837 (N_24837,N_24725,N_24692);
xor U24838 (N_24838,N_24712,N_24606);
nand U24839 (N_24839,N_24688,N_24764);
and U24840 (N_24840,N_24732,N_24785);
or U24841 (N_24841,N_24709,N_24690);
nand U24842 (N_24842,N_24787,N_24667);
and U24843 (N_24843,N_24738,N_24623);
xnor U24844 (N_24844,N_24745,N_24781);
xnor U24845 (N_24845,N_24731,N_24716);
nand U24846 (N_24846,N_24627,N_24793);
xor U24847 (N_24847,N_24723,N_24624);
xor U24848 (N_24848,N_24608,N_24699);
and U24849 (N_24849,N_24693,N_24644);
and U24850 (N_24850,N_24720,N_24698);
or U24851 (N_24851,N_24685,N_24614);
or U24852 (N_24852,N_24747,N_24645);
and U24853 (N_24853,N_24778,N_24796);
or U24854 (N_24854,N_24650,N_24612);
nor U24855 (N_24855,N_24705,N_24774);
and U24856 (N_24856,N_24792,N_24782);
nor U24857 (N_24857,N_24773,N_24617);
or U24858 (N_24858,N_24637,N_24655);
and U24859 (N_24859,N_24600,N_24769);
and U24860 (N_24860,N_24776,N_24786);
xnor U24861 (N_24861,N_24708,N_24648);
and U24862 (N_24862,N_24718,N_24611);
nor U24863 (N_24863,N_24681,N_24715);
nor U24864 (N_24864,N_24751,N_24727);
nand U24865 (N_24865,N_24652,N_24704);
nand U24866 (N_24866,N_24714,N_24628);
nand U24867 (N_24867,N_24756,N_24668);
and U24868 (N_24868,N_24615,N_24728);
nor U24869 (N_24869,N_24626,N_24757);
nand U24870 (N_24870,N_24657,N_24743);
xnor U24871 (N_24871,N_24639,N_24726);
nand U24872 (N_24872,N_24646,N_24724);
nand U24873 (N_24873,N_24766,N_24687);
nand U24874 (N_24874,N_24661,N_24749);
nor U24875 (N_24875,N_24737,N_24794);
nand U24876 (N_24876,N_24663,N_24795);
nor U24877 (N_24877,N_24706,N_24739);
nor U24878 (N_24878,N_24671,N_24618);
or U24879 (N_24879,N_24784,N_24744);
nand U24880 (N_24880,N_24719,N_24767);
and U24881 (N_24881,N_24770,N_24662);
nand U24882 (N_24882,N_24748,N_24703);
xor U24883 (N_24883,N_24733,N_24613);
nor U24884 (N_24884,N_24762,N_24779);
or U24885 (N_24885,N_24683,N_24601);
nand U24886 (N_24886,N_24654,N_24740);
and U24887 (N_24887,N_24678,N_24610);
xor U24888 (N_24888,N_24722,N_24603);
nand U24889 (N_24889,N_24619,N_24675);
xnor U24890 (N_24890,N_24656,N_24700);
xor U24891 (N_24891,N_24735,N_24660);
nor U24892 (N_24892,N_24791,N_24640);
and U24893 (N_24893,N_24742,N_24677);
xnor U24894 (N_24894,N_24630,N_24616);
nand U24895 (N_24895,N_24686,N_24783);
nor U24896 (N_24896,N_24797,N_24676);
nor U24897 (N_24897,N_24642,N_24772);
nand U24898 (N_24898,N_24799,N_24711);
nand U24899 (N_24899,N_24689,N_24780);
and U24900 (N_24900,N_24682,N_24678);
xnor U24901 (N_24901,N_24669,N_24779);
and U24902 (N_24902,N_24724,N_24718);
nor U24903 (N_24903,N_24699,N_24633);
and U24904 (N_24904,N_24721,N_24661);
and U24905 (N_24905,N_24749,N_24675);
nand U24906 (N_24906,N_24779,N_24780);
and U24907 (N_24907,N_24609,N_24771);
xnor U24908 (N_24908,N_24743,N_24764);
nor U24909 (N_24909,N_24720,N_24656);
and U24910 (N_24910,N_24600,N_24755);
nand U24911 (N_24911,N_24778,N_24690);
xnor U24912 (N_24912,N_24677,N_24664);
or U24913 (N_24913,N_24751,N_24705);
or U24914 (N_24914,N_24687,N_24725);
and U24915 (N_24915,N_24745,N_24682);
or U24916 (N_24916,N_24690,N_24647);
nand U24917 (N_24917,N_24668,N_24799);
nor U24918 (N_24918,N_24790,N_24713);
nand U24919 (N_24919,N_24749,N_24648);
nand U24920 (N_24920,N_24728,N_24633);
or U24921 (N_24921,N_24621,N_24681);
nor U24922 (N_24922,N_24671,N_24698);
or U24923 (N_24923,N_24685,N_24759);
and U24924 (N_24924,N_24609,N_24660);
nor U24925 (N_24925,N_24664,N_24789);
xor U24926 (N_24926,N_24743,N_24705);
xnor U24927 (N_24927,N_24619,N_24682);
nand U24928 (N_24928,N_24752,N_24793);
or U24929 (N_24929,N_24684,N_24794);
or U24930 (N_24930,N_24732,N_24724);
or U24931 (N_24931,N_24765,N_24662);
and U24932 (N_24932,N_24762,N_24645);
or U24933 (N_24933,N_24757,N_24782);
nand U24934 (N_24934,N_24666,N_24757);
nor U24935 (N_24935,N_24602,N_24658);
and U24936 (N_24936,N_24745,N_24629);
xor U24937 (N_24937,N_24657,N_24777);
nand U24938 (N_24938,N_24614,N_24630);
nand U24939 (N_24939,N_24633,N_24735);
and U24940 (N_24940,N_24693,N_24711);
and U24941 (N_24941,N_24752,N_24659);
or U24942 (N_24942,N_24654,N_24721);
nor U24943 (N_24943,N_24743,N_24765);
or U24944 (N_24944,N_24779,N_24709);
nor U24945 (N_24945,N_24673,N_24691);
or U24946 (N_24946,N_24744,N_24780);
nor U24947 (N_24947,N_24788,N_24753);
nor U24948 (N_24948,N_24626,N_24762);
xnor U24949 (N_24949,N_24709,N_24739);
xor U24950 (N_24950,N_24785,N_24673);
nor U24951 (N_24951,N_24793,N_24749);
or U24952 (N_24952,N_24742,N_24672);
nor U24953 (N_24953,N_24615,N_24754);
and U24954 (N_24954,N_24774,N_24762);
nand U24955 (N_24955,N_24798,N_24746);
xor U24956 (N_24956,N_24631,N_24771);
and U24957 (N_24957,N_24629,N_24763);
xor U24958 (N_24958,N_24656,N_24636);
nor U24959 (N_24959,N_24720,N_24785);
or U24960 (N_24960,N_24634,N_24681);
xor U24961 (N_24961,N_24616,N_24641);
and U24962 (N_24962,N_24688,N_24697);
or U24963 (N_24963,N_24621,N_24795);
nand U24964 (N_24964,N_24636,N_24776);
nor U24965 (N_24965,N_24796,N_24671);
xnor U24966 (N_24966,N_24764,N_24637);
nor U24967 (N_24967,N_24617,N_24772);
nor U24968 (N_24968,N_24624,N_24687);
nor U24969 (N_24969,N_24637,N_24709);
or U24970 (N_24970,N_24789,N_24686);
nor U24971 (N_24971,N_24668,N_24692);
nand U24972 (N_24972,N_24697,N_24609);
xor U24973 (N_24973,N_24776,N_24639);
or U24974 (N_24974,N_24636,N_24611);
nor U24975 (N_24975,N_24688,N_24663);
or U24976 (N_24976,N_24779,N_24705);
xor U24977 (N_24977,N_24737,N_24696);
and U24978 (N_24978,N_24724,N_24722);
and U24979 (N_24979,N_24728,N_24624);
xnor U24980 (N_24980,N_24608,N_24745);
nand U24981 (N_24981,N_24668,N_24767);
xnor U24982 (N_24982,N_24610,N_24728);
xor U24983 (N_24983,N_24612,N_24665);
or U24984 (N_24984,N_24684,N_24635);
or U24985 (N_24985,N_24762,N_24751);
nand U24986 (N_24986,N_24739,N_24648);
nand U24987 (N_24987,N_24704,N_24749);
and U24988 (N_24988,N_24744,N_24618);
xor U24989 (N_24989,N_24673,N_24705);
xnor U24990 (N_24990,N_24771,N_24718);
and U24991 (N_24991,N_24639,N_24763);
xor U24992 (N_24992,N_24607,N_24773);
xor U24993 (N_24993,N_24739,N_24623);
or U24994 (N_24994,N_24733,N_24624);
or U24995 (N_24995,N_24690,N_24649);
nand U24996 (N_24996,N_24733,N_24617);
nand U24997 (N_24997,N_24641,N_24610);
and U24998 (N_24998,N_24707,N_24734);
nand U24999 (N_24999,N_24729,N_24693);
xnor UO_0 (O_0,N_24930,N_24858);
nor UO_1 (O_1,N_24842,N_24873);
or UO_2 (O_2,N_24823,N_24992);
xnor UO_3 (O_3,N_24815,N_24839);
nand UO_4 (O_4,N_24817,N_24949);
and UO_5 (O_5,N_24890,N_24897);
nor UO_6 (O_6,N_24855,N_24923);
nor UO_7 (O_7,N_24971,N_24834);
or UO_8 (O_8,N_24970,N_24850);
or UO_9 (O_9,N_24937,N_24803);
xor UO_10 (O_10,N_24812,N_24991);
nand UO_11 (O_11,N_24905,N_24904);
xor UO_12 (O_12,N_24857,N_24848);
and UO_13 (O_13,N_24888,N_24926);
nor UO_14 (O_14,N_24969,N_24861);
nor UO_15 (O_15,N_24977,N_24898);
xnor UO_16 (O_16,N_24827,N_24875);
or UO_17 (O_17,N_24979,N_24957);
xnor UO_18 (O_18,N_24835,N_24990);
and UO_19 (O_19,N_24993,N_24843);
and UO_20 (O_20,N_24882,N_24879);
nand UO_21 (O_21,N_24880,N_24961);
xnor UO_22 (O_22,N_24872,N_24996);
nor UO_23 (O_23,N_24844,N_24901);
or UO_24 (O_24,N_24954,N_24945);
xor UO_25 (O_25,N_24852,N_24947);
nand UO_26 (O_26,N_24938,N_24856);
and UO_27 (O_27,N_24909,N_24907);
nand UO_28 (O_28,N_24874,N_24900);
xnor UO_29 (O_29,N_24838,N_24982);
xnor UO_30 (O_30,N_24942,N_24801);
nand UO_31 (O_31,N_24948,N_24944);
and UO_32 (O_32,N_24840,N_24972);
nand UO_33 (O_33,N_24809,N_24849);
nor UO_34 (O_34,N_24864,N_24928);
or UO_35 (O_35,N_24925,N_24881);
and UO_36 (O_36,N_24955,N_24895);
and UO_37 (O_37,N_24959,N_24952);
or UO_38 (O_38,N_24927,N_24813);
nor UO_39 (O_39,N_24988,N_24821);
nand UO_40 (O_40,N_24941,N_24885);
and UO_41 (O_41,N_24963,N_24946);
or UO_42 (O_42,N_24884,N_24894);
nor UO_43 (O_43,N_24912,N_24981);
nand UO_44 (O_44,N_24870,N_24968);
nor UO_45 (O_45,N_24903,N_24865);
xnor UO_46 (O_46,N_24965,N_24915);
xor UO_47 (O_47,N_24820,N_24899);
and UO_48 (O_48,N_24859,N_24845);
and UO_49 (O_49,N_24924,N_24953);
nand UO_50 (O_50,N_24985,N_24931);
xor UO_51 (O_51,N_24964,N_24829);
and UO_52 (O_52,N_24854,N_24832);
and UO_53 (O_53,N_24935,N_24878);
nand UO_54 (O_54,N_24847,N_24974);
or UO_55 (O_55,N_24920,N_24833);
and UO_56 (O_56,N_24814,N_24987);
nor UO_57 (O_57,N_24999,N_24860);
xor UO_58 (O_58,N_24911,N_24913);
and UO_59 (O_59,N_24916,N_24922);
xnor UO_60 (O_60,N_24932,N_24933);
nor UO_61 (O_61,N_24891,N_24863);
nor UO_62 (O_62,N_24984,N_24994);
xor UO_63 (O_63,N_24997,N_24950);
xor UO_64 (O_64,N_24975,N_24818);
nand UO_65 (O_65,N_24816,N_24846);
or UO_66 (O_66,N_24921,N_24837);
nand UO_67 (O_67,N_24826,N_24883);
or UO_68 (O_68,N_24986,N_24804);
and UO_69 (O_69,N_24828,N_24914);
nand UO_70 (O_70,N_24973,N_24887);
and UO_71 (O_71,N_24934,N_24917);
nor UO_72 (O_72,N_24951,N_24902);
and UO_73 (O_73,N_24807,N_24966);
nor UO_74 (O_74,N_24800,N_24805);
and UO_75 (O_75,N_24893,N_24998);
and UO_76 (O_76,N_24976,N_24978);
and UO_77 (O_77,N_24886,N_24811);
xnor UO_78 (O_78,N_24868,N_24802);
xor UO_79 (O_79,N_24906,N_24841);
and UO_80 (O_80,N_24836,N_24995);
or UO_81 (O_81,N_24851,N_24867);
and UO_82 (O_82,N_24824,N_24983);
xor UO_83 (O_83,N_24960,N_24876);
and UO_84 (O_84,N_24853,N_24936);
or UO_85 (O_85,N_24958,N_24980);
and UO_86 (O_86,N_24889,N_24810);
xor UO_87 (O_87,N_24939,N_24943);
or UO_88 (O_88,N_24896,N_24967);
and UO_89 (O_89,N_24910,N_24877);
nand UO_90 (O_90,N_24869,N_24866);
xnor UO_91 (O_91,N_24825,N_24822);
or UO_92 (O_92,N_24989,N_24862);
xor UO_93 (O_93,N_24808,N_24908);
nor UO_94 (O_94,N_24919,N_24892);
xor UO_95 (O_95,N_24830,N_24806);
nor UO_96 (O_96,N_24962,N_24956);
or UO_97 (O_97,N_24940,N_24929);
and UO_98 (O_98,N_24871,N_24819);
nand UO_99 (O_99,N_24831,N_24918);
or UO_100 (O_100,N_24936,N_24906);
or UO_101 (O_101,N_24983,N_24931);
or UO_102 (O_102,N_24992,N_24947);
xnor UO_103 (O_103,N_24817,N_24869);
xnor UO_104 (O_104,N_24974,N_24940);
xor UO_105 (O_105,N_24899,N_24948);
and UO_106 (O_106,N_24917,N_24944);
and UO_107 (O_107,N_24987,N_24938);
xor UO_108 (O_108,N_24809,N_24873);
nor UO_109 (O_109,N_24949,N_24825);
or UO_110 (O_110,N_24843,N_24877);
and UO_111 (O_111,N_24940,N_24973);
xor UO_112 (O_112,N_24880,N_24933);
xnor UO_113 (O_113,N_24986,N_24829);
xnor UO_114 (O_114,N_24808,N_24860);
nand UO_115 (O_115,N_24803,N_24876);
xnor UO_116 (O_116,N_24944,N_24836);
xor UO_117 (O_117,N_24864,N_24811);
xnor UO_118 (O_118,N_24954,N_24832);
nor UO_119 (O_119,N_24807,N_24844);
and UO_120 (O_120,N_24889,N_24812);
and UO_121 (O_121,N_24931,N_24844);
and UO_122 (O_122,N_24908,N_24925);
nand UO_123 (O_123,N_24936,N_24807);
or UO_124 (O_124,N_24846,N_24937);
nand UO_125 (O_125,N_24879,N_24904);
nor UO_126 (O_126,N_24937,N_24978);
nor UO_127 (O_127,N_24884,N_24877);
xor UO_128 (O_128,N_24969,N_24808);
nand UO_129 (O_129,N_24909,N_24813);
nand UO_130 (O_130,N_24810,N_24937);
xnor UO_131 (O_131,N_24918,N_24868);
nor UO_132 (O_132,N_24842,N_24958);
and UO_133 (O_133,N_24840,N_24883);
xor UO_134 (O_134,N_24878,N_24951);
or UO_135 (O_135,N_24997,N_24917);
xor UO_136 (O_136,N_24865,N_24945);
nand UO_137 (O_137,N_24881,N_24819);
nor UO_138 (O_138,N_24928,N_24849);
and UO_139 (O_139,N_24921,N_24952);
nor UO_140 (O_140,N_24992,N_24899);
and UO_141 (O_141,N_24809,N_24938);
nor UO_142 (O_142,N_24961,N_24945);
nand UO_143 (O_143,N_24842,N_24950);
nand UO_144 (O_144,N_24911,N_24894);
xnor UO_145 (O_145,N_24851,N_24882);
and UO_146 (O_146,N_24812,N_24819);
nand UO_147 (O_147,N_24958,N_24916);
nor UO_148 (O_148,N_24915,N_24936);
xnor UO_149 (O_149,N_24928,N_24917);
nor UO_150 (O_150,N_24977,N_24957);
or UO_151 (O_151,N_24924,N_24880);
and UO_152 (O_152,N_24856,N_24926);
or UO_153 (O_153,N_24992,N_24973);
and UO_154 (O_154,N_24866,N_24910);
nor UO_155 (O_155,N_24831,N_24857);
nand UO_156 (O_156,N_24882,N_24956);
xor UO_157 (O_157,N_24976,N_24827);
xnor UO_158 (O_158,N_24800,N_24924);
nor UO_159 (O_159,N_24960,N_24949);
nand UO_160 (O_160,N_24858,N_24875);
and UO_161 (O_161,N_24821,N_24805);
nand UO_162 (O_162,N_24893,N_24921);
nor UO_163 (O_163,N_24953,N_24939);
and UO_164 (O_164,N_24925,N_24857);
and UO_165 (O_165,N_24863,N_24934);
nand UO_166 (O_166,N_24846,N_24912);
xnor UO_167 (O_167,N_24918,N_24882);
xnor UO_168 (O_168,N_24868,N_24979);
xor UO_169 (O_169,N_24968,N_24929);
nor UO_170 (O_170,N_24845,N_24858);
xor UO_171 (O_171,N_24874,N_24833);
and UO_172 (O_172,N_24851,N_24824);
nor UO_173 (O_173,N_24977,N_24961);
or UO_174 (O_174,N_24872,N_24807);
and UO_175 (O_175,N_24846,N_24809);
nand UO_176 (O_176,N_24830,N_24964);
xor UO_177 (O_177,N_24812,N_24913);
nor UO_178 (O_178,N_24864,N_24872);
or UO_179 (O_179,N_24990,N_24890);
and UO_180 (O_180,N_24800,N_24957);
and UO_181 (O_181,N_24805,N_24919);
nor UO_182 (O_182,N_24809,N_24902);
nor UO_183 (O_183,N_24907,N_24883);
or UO_184 (O_184,N_24964,N_24957);
nand UO_185 (O_185,N_24911,N_24989);
nor UO_186 (O_186,N_24902,N_24981);
or UO_187 (O_187,N_24980,N_24868);
nand UO_188 (O_188,N_24957,N_24891);
or UO_189 (O_189,N_24833,N_24891);
and UO_190 (O_190,N_24939,N_24981);
or UO_191 (O_191,N_24853,N_24873);
and UO_192 (O_192,N_24800,N_24992);
nor UO_193 (O_193,N_24963,N_24978);
nand UO_194 (O_194,N_24839,N_24820);
nor UO_195 (O_195,N_24863,N_24920);
or UO_196 (O_196,N_24933,N_24808);
nand UO_197 (O_197,N_24936,N_24892);
nand UO_198 (O_198,N_24929,N_24880);
or UO_199 (O_199,N_24990,N_24930);
nor UO_200 (O_200,N_24952,N_24878);
nor UO_201 (O_201,N_24954,N_24975);
nor UO_202 (O_202,N_24939,N_24924);
and UO_203 (O_203,N_24958,N_24996);
and UO_204 (O_204,N_24881,N_24998);
and UO_205 (O_205,N_24875,N_24895);
and UO_206 (O_206,N_24995,N_24894);
and UO_207 (O_207,N_24820,N_24904);
nor UO_208 (O_208,N_24864,N_24802);
nor UO_209 (O_209,N_24844,N_24867);
or UO_210 (O_210,N_24877,N_24841);
xor UO_211 (O_211,N_24812,N_24873);
and UO_212 (O_212,N_24865,N_24972);
or UO_213 (O_213,N_24832,N_24893);
nand UO_214 (O_214,N_24818,N_24947);
and UO_215 (O_215,N_24969,N_24869);
or UO_216 (O_216,N_24943,N_24935);
nand UO_217 (O_217,N_24881,N_24849);
xor UO_218 (O_218,N_24858,N_24850);
and UO_219 (O_219,N_24824,N_24898);
and UO_220 (O_220,N_24855,N_24924);
or UO_221 (O_221,N_24810,N_24878);
nand UO_222 (O_222,N_24889,N_24974);
and UO_223 (O_223,N_24879,N_24811);
and UO_224 (O_224,N_24991,N_24910);
and UO_225 (O_225,N_24982,N_24935);
nand UO_226 (O_226,N_24947,N_24843);
or UO_227 (O_227,N_24931,N_24998);
or UO_228 (O_228,N_24871,N_24904);
nor UO_229 (O_229,N_24914,N_24885);
nand UO_230 (O_230,N_24946,N_24972);
xnor UO_231 (O_231,N_24937,N_24957);
and UO_232 (O_232,N_24832,N_24818);
nor UO_233 (O_233,N_24814,N_24835);
or UO_234 (O_234,N_24883,N_24830);
xor UO_235 (O_235,N_24879,N_24852);
nand UO_236 (O_236,N_24928,N_24867);
or UO_237 (O_237,N_24950,N_24898);
or UO_238 (O_238,N_24994,N_24860);
nor UO_239 (O_239,N_24970,N_24818);
or UO_240 (O_240,N_24936,N_24884);
nor UO_241 (O_241,N_24910,N_24916);
nor UO_242 (O_242,N_24866,N_24830);
and UO_243 (O_243,N_24895,N_24872);
xnor UO_244 (O_244,N_24816,N_24917);
nand UO_245 (O_245,N_24957,N_24973);
and UO_246 (O_246,N_24805,N_24892);
or UO_247 (O_247,N_24849,N_24922);
xor UO_248 (O_248,N_24987,N_24831);
nand UO_249 (O_249,N_24833,N_24946);
nor UO_250 (O_250,N_24850,N_24839);
or UO_251 (O_251,N_24813,N_24922);
and UO_252 (O_252,N_24835,N_24970);
or UO_253 (O_253,N_24856,N_24873);
or UO_254 (O_254,N_24921,N_24812);
and UO_255 (O_255,N_24836,N_24915);
nor UO_256 (O_256,N_24906,N_24813);
and UO_257 (O_257,N_24837,N_24816);
nand UO_258 (O_258,N_24878,N_24815);
nand UO_259 (O_259,N_24893,N_24985);
or UO_260 (O_260,N_24832,N_24998);
xor UO_261 (O_261,N_24901,N_24984);
nor UO_262 (O_262,N_24929,N_24973);
nor UO_263 (O_263,N_24936,N_24976);
xor UO_264 (O_264,N_24840,N_24954);
and UO_265 (O_265,N_24939,N_24960);
and UO_266 (O_266,N_24855,N_24828);
and UO_267 (O_267,N_24885,N_24833);
or UO_268 (O_268,N_24878,N_24859);
xor UO_269 (O_269,N_24841,N_24892);
and UO_270 (O_270,N_24917,N_24832);
nor UO_271 (O_271,N_24889,N_24891);
nand UO_272 (O_272,N_24882,N_24917);
or UO_273 (O_273,N_24854,N_24955);
and UO_274 (O_274,N_24978,N_24901);
nand UO_275 (O_275,N_24883,N_24964);
xnor UO_276 (O_276,N_24986,N_24926);
nand UO_277 (O_277,N_24922,N_24893);
nor UO_278 (O_278,N_24802,N_24956);
nand UO_279 (O_279,N_24913,N_24885);
xnor UO_280 (O_280,N_24895,N_24820);
nor UO_281 (O_281,N_24949,N_24923);
nand UO_282 (O_282,N_24860,N_24854);
or UO_283 (O_283,N_24802,N_24884);
xor UO_284 (O_284,N_24841,N_24858);
nor UO_285 (O_285,N_24911,N_24810);
nor UO_286 (O_286,N_24972,N_24829);
or UO_287 (O_287,N_24994,N_24995);
xnor UO_288 (O_288,N_24934,N_24923);
and UO_289 (O_289,N_24927,N_24845);
nand UO_290 (O_290,N_24875,N_24889);
xor UO_291 (O_291,N_24845,N_24926);
xor UO_292 (O_292,N_24975,N_24908);
or UO_293 (O_293,N_24936,N_24898);
xnor UO_294 (O_294,N_24911,N_24869);
or UO_295 (O_295,N_24982,N_24939);
xor UO_296 (O_296,N_24808,N_24843);
and UO_297 (O_297,N_24962,N_24909);
xnor UO_298 (O_298,N_24914,N_24982);
nor UO_299 (O_299,N_24925,N_24905);
nand UO_300 (O_300,N_24845,N_24936);
nor UO_301 (O_301,N_24977,N_24929);
nand UO_302 (O_302,N_24978,N_24864);
and UO_303 (O_303,N_24984,N_24924);
xor UO_304 (O_304,N_24835,N_24898);
xor UO_305 (O_305,N_24805,N_24984);
xor UO_306 (O_306,N_24805,N_24977);
or UO_307 (O_307,N_24843,N_24977);
nor UO_308 (O_308,N_24958,N_24837);
xor UO_309 (O_309,N_24897,N_24802);
nand UO_310 (O_310,N_24824,N_24936);
and UO_311 (O_311,N_24983,N_24831);
nor UO_312 (O_312,N_24901,N_24972);
or UO_313 (O_313,N_24864,N_24859);
and UO_314 (O_314,N_24906,N_24991);
xnor UO_315 (O_315,N_24909,N_24803);
nor UO_316 (O_316,N_24966,N_24853);
and UO_317 (O_317,N_24837,N_24898);
xor UO_318 (O_318,N_24875,N_24924);
nand UO_319 (O_319,N_24828,N_24867);
and UO_320 (O_320,N_24992,N_24898);
nor UO_321 (O_321,N_24995,N_24823);
nand UO_322 (O_322,N_24896,N_24812);
nor UO_323 (O_323,N_24914,N_24964);
nor UO_324 (O_324,N_24993,N_24962);
xor UO_325 (O_325,N_24945,N_24829);
nand UO_326 (O_326,N_24901,N_24862);
or UO_327 (O_327,N_24994,N_24924);
or UO_328 (O_328,N_24967,N_24803);
xor UO_329 (O_329,N_24838,N_24882);
xor UO_330 (O_330,N_24919,N_24876);
or UO_331 (O_331,N_24884,N_24983);
xor UO_332 (O_332,N_24986,N_24896);
xor UO_333 (O_333,N_24886,N_24830);
nand UO_334 (O_334,N_24896,N_24945);
or UO_335 (O_335,N_24890,N_24971);
and UO_336 (O_336,N_24958,N_24850);
and UO_337 (O_337,N_24961,N_24993);
xnor UO_338 (O_338,N_24964,N_24986);
or UO_339 (O_339,N_24956,N_24860);
nand UO_340 (O_340,N_24871,N_24903);
xnor UO_341 (O_341,N_24922,N_24866);
or UO_342 (O_342,N_24905,N_24990);
nor UO_343 (O_343,N_24898,N_24906);
nand UO_344 (O_344,N_24941,N_24863);
or UO_345 (O_345,N_24986,N_24925);
nand UO_346 (O_346,N_24882,N_24912);
nor UO_347 (O_347,N_24954,N_24952);
nand UO_348 (O_348,N_24941,N_24956);
and UO_349 (O_349,N_24945,N_24803);
nor UO_350 (O_350,N_24914,N_24847);
nand UO_351 (O_351,N_24945,N_24956);
and UO_352 (O_352,N_24877,N_24952);
and UO_353 (O_353,N_24912,N_24990);
or UO_354 (O_354,N_24931,N_24915);
and UO_355 (O_355,N_24859,N_24986);
nand UO_356 (O_356,N_24964,N_24996);
or UO_357 (O_357,N_24858,N_24919);
nor UO_358 (O_358,N_24949,N_24835);
nor UO_359 (O_359,N_24977,N_24963);
or UO_360 (O_360,N_24803,N_24820);
xor UO_361 (O_361,N_24952,N_24876);
and UO_362 (O_362,N_24833,N_24890);
and UO_363 (O_363,N_24869,N_24899);
nor UO_364 (O_364,N_24978,N_24853);
nor UO_365 (O_365,N_24933,N_24841);
nor UO_366 (O_366,N_24829,N_24912);
nand UO_367 (O_367,N_24852,N_24992);
nand UO_368 (O_368,N_24943,N_24927);
and UO_369 (O_369,N_24861,N_24899);
or UO_370 (O_370,N_24826,N_24936);
nand UO_371 (O_371,N_24894,N_24918);
and UO_372 (O_372,N_24964,N_24905);
nor UO_373 (O_373,N_24962,N_24860);
and UO_374 (O_374,N_24834,N_24955);
xnor UO_375 (O_375,N_24986,N_24850);
xnor UO_376 (O_376,N_24976,N_24910);
or UO_377 (O_377,N_24895,N_24949);
nor UO_378 (O_378,N_24912,N_24815);
xnor UO_379 (O_379,N_24896,N_24992);
nor UO_380 (O_380,N_24837,N_24871);
nand UO_381 (O_381,N_24832,N_24834);
nand UO_382 (O_382,N_24947,N_24900);
or UO_383 (O_383,N_24992,N_24881);
or UO_384 (O_384,N_24991,N_24995);
nor UO_385 (O_385,N_24923,N_24823);
and UO_386 (O_386,N_24813,N_24822);
nand UO_387 (O_387,N_24800,N_24958);
or UO_388 (O_388,N_24872,N_24938);
xor UO_389 (O_389,N_24870,N_24987);
or UO_390 (O_390,N_24986,N_24807);
and UO_391 (O_391,N_24967,N_24913);
and UO_392 (O_392,N_24884,N_24821);
xor UO_393 (O_393,N_24946,N_24805);
xor UO_394 (O_394,N_24865,N_24983);
xor UO_395 (O_395,N_24933,N_24824);
and UO_396 (O_396,N_24867,N_24982);
and UO_397 (O_397,N_24803,N_24801);
xnor UO_398 (O_398,N_24855,N_24938);
and UO_399 (O_399,N_24801,N_24877);
nor UO_400 (O_400,N_24899,N_24847);
nand UO_401 (O_401,N_24919,N_24934);
nand UO_402 (O_402,N_24848,N_24832);
xor UO_403 (O_403,N_24809,N_24898);
or UO_404 (O_404,N_24959,N_24936);
xor UO_405 (O_405,N_24970,N_24962);
and UO_406 (O_406,N_24909,N_24993);
nand UO_407 (O_407,N_24944,N_24835);
xor UO_408 (O_408,N_24850,N_24991);
nor UO_409 (O_409,N_24966,N_24816);
nand UO_410 (O_410,N_24969,N_24858);
xnor UO_411 (O_411,N_24987,N_24955);
or UO_412 (O_412,N_24984,N_24946);
xnor UO_413 (O_413,N_24910,N_24967);
nand UO_414 (O_414,N_24803,N_24954);
nor UO_415 (O_415,N_24926,N_24925);
and UO_416 (O_416,N_24992,N_24959);
or UO_417 (O_417,N_24800,N_24861);
nand UO_418 (O_418,N_24812,N_24966);
xnor UO_419 (O_419,N_24911,N_24909);
xnor UO_420 (O_420,N_24931,N_24847);
nand UO_421 (O_421,N_24962,N_24804);
and UO_422 (O_422,N_24839,N_24830);
and UO_423 (O_423,N_24907,N_24807);
nor UO_424 (O_424,N_24878,N_24985);
xnor UO_425 (O_425,N_24901,N_24973);
nor UO_426 (O_426,N_24903,N_24820);
xor UO_427 (O_427,N_24856,N_24850);
and UO_428 (O_428,N_24831,N_24937);
or UO_429 (O_429,N_24936,N_24841);
and UO_430 (O_430,N_24841,N_24871);
nor UO_431 (O_431,N_24929,N_24990);
xor UO_432 (O_432,N_24807,N_24836);
xnor UO_433 (O_433,N_24824,N_24967);
or UO_434 (O_434,N_24884,N_24883);
and UO_435 (O_435,N_24894,N_24933);
or UO_436 (O_436,N_24826,N_24991);
nor UO_437 (O_437,N_24934,N_24911);
nand UO_438 (O_438,N_24805,N_24807);
nand UO_439 (O_439,N_24950,N_24879);
nand UO_440 (O_440,N_24840,N_24865);
and UO_441 (O_441,N_24866,N_24907);
or UO_442 (O_442,N_24833,N_24978);
nor UO_443 (O_443,N_24800,N_24834);
nand UO_444 (O_444,N_24983,N_24985);
and UO_445 (O_445,N_24936,N_24856);
nand UO_446 (O_446,N_24940,N_24831);
or UO_447 (O_447,N_24919,N_24976);
nor UO_448 (O_448,N_24834,N_24953);
nand UO_449 (O_449,N_24802,N_24887);
and UO_450 (O_450,N_24920,N_24816);
nor UO_451 (O_451,N_24831,N_24966);
or UO_452 (O_452,N_24972,N_24897);
nor UO_453 (O_453,N_24940,N_24923);
nor UO_454 (O_454,N_24925,N_24836);
or UO_455 (O_455,N_24919,N_24814);
xor UO_456 (O_456,N_24806,N_24974);
nand UO_457 (O_457,N_24863,N_24987);
xnor UO_458 (O_458,N_24940,N_24801);
or UO_459 (O_459,N_24896,N_24803);
or UO_460 (O_460,N_24930,N_24991);
nand UO_461 (O_461,N_24907,N_24863);
nand UO_462 (O_462,N_24915,N_24917);
xor UO_463 (O_463,N_24867,N_24808);
or UO_464 (O_464,N_24850,N_24995);
nand UO_465 (O_465,N_24977,N_24923);
and UO_466 (O_466,N_24854,N_24834);
or UO_467 (O_467,N_24979,N_24920);
xor UO_468 (O_468,N_24963,N_24839);
and UO_469 (O_469,N_24863,N_24972);
and UO_470 (O_470,N_24991,N_24863);
or UO_471 (O_471,N_24870,N_24931);
or UO_472 (O_472,N_24865,N_24907);
and UO_473 (O_473,N_24814,N_24881);
nand UO_474 (O_474,N_24805,N_24847);
nor UO_475 (O_475,N_24866,N_24801);
xnor UO_476 (O_476,N_24852,N_24873);
nand UO_477 (O_477,N_24910,N_24961);
and UO_478 (O_478,N_24935,N_24839);
and UO_479 (O_479,N_24931,N_24900);
xnor UO_480 (O_480,N_24908,N_24819);
and UO_481 (O_481,N_24955,N_24892);
nor UO_482 (O_482,N_24817,N_24800);
nor UO_483 (O_483,N_24878,N_24814);
nor UO_484 (O_484,N_24907,N_24995);
nand UO_485 (O_485,N_24816,N_24869);
xor UO_486 (O_486,N_24890,N_24950);
nor UO_487 (O_487,N_24829,N_24856);
nor UO_488 (O_488,N_24890,N_24884);
xnor UO_489 (O_489,N_24834,N_24992);
nand UO_490 (O_490,N_24922,N_24886);
or UO_491 (O_491,N_24890,N_24824);
nor UO_492 (O_492,N_24847,N_24904);
nand UO_493 (O_493,N_24817,N_24933);
xor UO_494 (O_494,N_24997,N_24860);
xnor UO_495 (O_495,N_24839,N_24939);
xnor UO_496 (O_496,N_24966,N_24844);
xnor UO_497 (O_497,N_24849,N_24956);
and UO_498 (O_498,N_24969,N_24919);
or UO_499 (O_499,N_24930,N_24935);
nor UO_500 (O_500,N_24981,N_24958);
and UO_501 (O_501,N_24949,N_24831);
nand UO_502 (O_502,N_24927,N_24850);
nor UO_503 (O_503,N_24853,N_24959);
and UO_504 (O_504,N_24834,N_24803);
xor UO_505 (O_505,N_24802,N_24819);
xor UO_506 (O_506,N_24869,N_24910);
or UO_507 (O_507,N_24909,N_24942);
nor UO_508 (O_508,N_24897,N_24904);
or UO_509 (O_509,N_24990,N_24972);
nor UO_510 (O_510,N_24950,N_24886);
and UO_511 (O_511,N_24859,N_24821);
or UO_512 (O_512,N_24813,N_24864);
and UO_513 (O_513,N_24849,N_24905);
or UO_514 (O_514,N_24939,N_24954);
and UO_515 (O_515,N_24808,N_24934);
nor UO_516 (O_516,N_24981,N_24995);
or UO_517 (O_517,N_24864,N_24901);
nor UO_518 (O_518,N_24865,N_24812);
or UO_519 (O_519,N_24973,N_24871);
xor UO_520 (O_520,N_24907,N_24918);
xor UO_521 (O_521,N_24887,N_24942);
or UO_522 (O_522,N_24985,N_24949);
nand UO_523 (O_523,N_24842,N_24844);
nand UO_524 (O_524,N_24872,N_24979);
or UO_525 (O_525,N_24821,N_24803);
nand UO_526 (O_526,N_24800,N_24967);
nor UO_527 (O_527,N_24908,N_24992);
nor UO_528 (O_528,N_24937,N_24842);
and UO_529 (O_529,N_24920,N_24902);
nand UO_530 (O_530,N_24873,N_24867);
xor UO_531 (O_531,N_24975,N_24872);
or UO_532 (O_532,N_24935,N_24888);
or UO_533 (O_533,N_24835,N_24865);
xor UO_534 (O_534,N_24843,N_24944);
or UO_535 (O_535,N_24975,N_24944);
or UO_536 (O_536,N_24838,N_24862);
xnor UO_537 (O_537,N_24914,N_24978);
xor UO_538 (O_538,N_24989,N_24889);
xor UO_539 (O_539,N_24917,N_24950);
nand UO_540 (O_540,N_24928,N_24853);
xnor UO_541 (O_541,N_24922,N_24984);
or UO_542 (O_542,N_24914,N_24809);
nor UO_543 (O_543,N_24903,N_24821);
nand UO_544 (O_544,N_24949,N_24860);
or UO_545 (O_545,N_24868,N_24961);
or UO_546 (O_546,N_24830,N_24800);
nand UO_547 (O_547,N_24977,N_24816);
nand UO_548 (O_548,N_24888,N_24969);
nand UO_549 (O_549,N_24841,N_24986);
nand UO_550 (O_550,N_24976,N_24917);
xnor UO_551 (O_551,N_24914,N_24803);
nand UO_552 (O_552,N_24899,N_24986);
and UO_553 (O_553,N_24864,N_24969);
xnor UO_554 (O_554,N_24866,N_24841);
nor UO_555 (O_555,N_24933,N_24988);
or UO_556 (O_556,N_24844,N_24968);
nor UO_557 (O_557,N_24953,N_24946);
nand UO_558 (O_558,N_24978,N_24928);
nand UO_559 (O_559,N_24917,N_24901);
or UO_560 (O_560,N_24834,N_24959);
and UO_561 (O_561,N_24943,N_24825);
or UO_562 (O_562,N_24810,N_24952);
and UO_563 (O_563,N_24817,N_24904);
nor UO_564 (O_564,N_24915,N_24971);
xor UO_565 (O_565,N_24883,N_24932);
or UO_566 (O_566,N_24882,N_24930);
nor UO_567 (O_567,N_24932,N_24973);
or UO_568 (O_568,N_24940,N_24891);
or UO_569 (O_569,N_24910,N_24805);
nand UO_570 (O_570,N_24913,N_24896);
nor UO_571 (O_571,N_24971,N_24814);
or UO_572 (O_572,N_24994,N_24820);
and UO_573 (O_573,N_24995,N_24977);
nand UO_574 (O_574,N_24871,N_24836);
and UO_575 (O_575,N_24933,N_24898);
or UO_576 (O_576,N_24897,N_24948);
and UO_577 (O_577,N_24896,N_24820);
nand UO_578 (O_578,N_24966,N_24841);
xnor UO_579 (O_579,N_24905,N_24881);
nand UO_580 (O_580,N_24808,N_24983);
or UO_581 (O_581,N_24888,N_24992);
nand UO_582 (O_582,N_24852,N_24886);
nand UO_583 (O_583,N_24997,N_24853);
and UO_584 (O_584,N_24864,N_24883);
nor UO_585 (O_585,N_24841,N_24836);
nor UO_586 (O_586,N_24809,N_24847);
xor UO_587 (O_587,N_24821,N_24807);
nor UO_588 (O_588,N_24809,N_24947);
and UO_589 (O_589,N_24972,N_24845);
and UO_590 (O_590,N_24810,N_24805);
xnor UO_591 (O_591,N_24821,N_24802);
or UO_592 (O_592,N_24912,N_24888);
or UO_593 (O_593,N_24901,N_24995);
nand UO_594 (O_594,N_24871,N_24925);
or UO_595 (O_595,N_24953,N_24889);
xor UO_596 (O_596,N_24807,N_24984);
nor UO_597 (O_597,N_24890,N_24804);
xor UO_598 (O_598,N_24817,N_24897);
nand UO_599 (O_599,N_24866,N_24938);
xnor UO_600 (O_600,N_24986,N_24895);
and UO_601 (O_601,N_24948,N_24882);
nor UO_602 (O_602,N_24878,N_24837);
nand UO_603 (O_603,N_24824,N_24818);
nand UO_604 (O_604,N_24807,N_24949);
and UO_605 (O_605,N_24858,N_24839);
nor UO_606 (O_606,N_24924,N_24842);
nand UO_607 (O_607,N_24852,N_24939);
or UO_608 (O_608,N_24983,N_24804);
and UO_609 (O_609,N_24956,N_24954);
or UO_610 (O_610,N_24823,N_24884);
nand UO_611 (O_611,N_24887,N_24974);
nor UO_612 (O_612,N_24943,N_24964);
and UO_613 (O_613,N_24863,N_24917);
and UO_614 (O_614,N_24920,N_24887);
and UO_615 (O_615,N_24866,N_24918);
nand UO_616 (O_616,N_24812,N_24911);
nand UO_617 (O_617,N_24939,N_24800);
nor UO_618 (O_618,N_24823,N_24967);
and UO_619 (O_619,N_24962,N_24884);
or UO_620 (O_620,N_24950,N_24887);
and UO_621 (O_621,N_24854,N_24911);
nor UO_622 (O_622,N_24931,N_24947);
nor UO_623 (O_623,N_24982,N_24997);
and UO_624 (O_624,N_24976,N_24802);
nor UO_625 (O_625,N_24870,N_24949);
and UO_626 (O_626,N_24923,N_24879);
xnor UO_627 (O_627,N_24885,N_24858);
and UO_628 (O_628,N_24836,N_24860);
xor UO_629 (O_629,N_24981,N_24921);
and UO_630 (O_630,N_24930,N_24865);
or UO_631 (O_631,N_24919,N_24886);
nor UO_632 (O_632,N_24897,N_24842);
and UO_633 (O_633,N_24965,N_24933);
nand UO_634 (O_634,N_24910,N_24941);
nor UO_635 (O_635,N_24906,N_24918);
xnor UO_636 (O_636,N_24887,N_24985);
nor UO_637 (O_637,N_24800,N_24835);
or UO_638 (O_638,N_24842,N_24917);
or UO_639 (O_639,N_24960,N_24984);
and UO_640 (O_640,N_24838,N_24993);
or UO_641 (O_641,N_24896,N_24844);
or UO_642 (O_642,N_24915,N_24808);
nand UO_643 (O_643,N_24988,N_24889);
nor UO_644 (O_644,N_24969,N_24815);
or UO_645 (O_645,N_24877,N_24993);
or UO_646 (O_646,N_24916,N_24906);
nor UO_647 (O_647,N_24926,N_24832);
xnor UO_648 (O_648,N_24820,N_24972);
xnor UO_649 (O_649,N_24986,N_24892);
xnor UO_650 (O_650,N_24927,N_24887);
nor UO_651 (O_651,N_24903,N_24901);
nor UO_652 (O_652,N_24814,N_24950);
nand UO_653 (O_653,N_24935,N_24957);
nor UO_654 (O_654,N_24883,N_24920);
or UO_655 (O_655,N_24944,N_24925);
nand UO_656 (O_656,N_24853,N_24987);
or UO_657 (O_657,N_24917,N_24806);
and UO_658 (O_658,N_24980,N_24818);
nor UO_659 (O_659,N_24846,N_24928);
xnor UO_660 (O_660,N_24918,N_24801);
xnor UO_661 (O_661,N_24875,N_24902);
nor UO_662 (O_662,N_24837,N_24939);
and UO_663 (O_663,N_24979,N_24910);
and UO_664 (O_664,N_24808,N_24941);
nor UO_665 (O_665,N_24879,N_24877);
nand UO_666 (O_666,N_24923,N_24865);
nand UO_667 (O_667,N_24961,N_24994);
nand UO_668 (O_668,N_24959,N_24846);
xor UO_669 (O_669,N_24947,N_24973);
or UO_670 (O_670,N_24928,N_24991);
and UO_671 (O_671,N_24977,N_24857);
nor UO_672 (O_672,N_24837,N_24857);
and UO_673 (O_673,N_24899,N_24917);
or UO_674 (O_674,N_24871,N_24975);
or UO_675 (O_675,N_24981,N_24852);
nor UO_676 (O_676,N_24809,N_24901);
nor UO_677 (O_677,N_24923,N_24805);
nand UO_678 (O_678,N_24969,N_24837);
xnor UO_679 (O_679,N_24803,N_24811);
and UO_680 (O_680,N_24802,N_24930);
or UO_681 (O_681,N_24885,N_24918);
nand UO_682 (O_682,N_24832,N_24835);
or UO_683 (O_683,N_24873,N_24976);
or UO_684 (O_684,N_24820,N_24931);
or UO_685 (O_685,N_24978,N_24803);
or UO_686 (O_686,N_24887,N_24939);
nor UO_687 (O_687,N_24957,N_24898);
and UO_688 (O_688,N_24947,N_24923);
xor UO_689 (O_689,N_24915,N_24831);
and UO_690 (O_690,N_24925,N_24878);
and UO_691 (O_691,N_24972,N_24970);
or UO_692 (O_692,N_24860,N_24835);
or UO_693 (O_693,N_24888,N_24886);
nor UO_694 (O_694,N_24881,N_24847);
or UO_695 (O_695,N_24814,N_24986);
or UO_696 (O_696,N_24806,N_24937);
xor UO_697 (O_697,N_24941,N_24882);
nor UO_698 (O_698,N_24950,N_24965);
or UO_699 (O_699,N_24935,N_24836);
nand UO_700 (O_700,N_24907,N_24964);
nor UO_701 (O_701,N_24991,N_24907);
xor UO_702 (O_702,N_24803,N_24985);
nor UO_703 (O_703,N_24806,N_24906);
or UO_704 (O_704,N_24965,N_24856);
or UO_705 (O_705,N_24911,N_24944);
nand UO_706 (O_706,N_24916,N_24913);
and UO_707 (O_707,N_24991,N_24921);
xor UO_708 (O_708,N_24907,N_24838);
and UO_709 (O_709,N_24924,N_24922);
xor UO_710 (O_710,N_24875,N_24956);
and UO_711 (O_711,N_24960,N_24914);
nor UO_712 (O_712,N_24997,N_24992);
nand UO_713 (O_713,N_24958,N_24987);
nor UO_714 (O_714,N_24808,N_24937);
nor UO_715 (O_715,N_24969,N_24882);
and UO_716 (O_716,N_24825,N_24826);
or UO_717 (O_717,N_24901,N_24982);
nor UO_718 (O_718,N_24893,N_24914);
or UO_719 (O_719,N_24995,N_24820);
nand UO_720 (O_720,N_24807,N_24843);
nor UO_721 (O_721,N_24967,N_24898);
nand UO_722 (O_722,N_24986,N_24952);
xnor UO_723 (O_723,N_24956,N_24932);
nor UO_724 (O_724,N_24989,N_24915);
nand UO_725 (O_725,N_24968,N_24839);
and UO_726 (O_726,N_24923,N_24824);
xnor UO_727 (O_727,N_24843,N_24903);
and UO_728 (O_728,N_24937,N_24848);
nor UO_729 (O_729,N_24913,N_24803);
or UO_730 (O_730,N_24874,N_24854);
nand UO_731 (O_731,N_24957,N_24949);
and UO_732 (O_732,N_24987,N_24959);
and UO_733 (O_733,N_24812,N_24993);
and UO_734 (O_734,N_24826,N_24917);
or UO_735 (O_735,N_24883,N_24990);
nor UO_736 (O_736,N_24857,N_24951);
or UO_737 (O_737,N_24894,N_24829);
and UO_738 (O_738,N_24898,N_24902);
xor UO_739 (O_739,N_24896,N_24952);
nor UO_740 (O_740,N_24915,N_24805);
nand UO_741 (O_741,N_24890,N_24923);
nor UO_742 (O_742,N_24951,N_24881);
and UO_743 (O_743,N_24938,N_24858);
xnor UO_744 (O_744,N_24992,N_24941);
and UO_745 (O_745,N_24982,N_24815);
nand UO_746 (O_746,N_24850,N_24996);
or UO_747 (O_747,N_24856,N_24888);
nand UO_748 (O_748,N_24823,N_24899);
xnor UO_749 (O_749,N_24938,N_24917);
xnor UO_750 (O_750,N_24962,N_24953);
nand UO_751 (O_751,N_24902,N_24832);
or UO_752 (O_752,N_24956,N_24841);
nor UO_753 (O_753,N_24943,N_24881);
or UO_754 (O_754,N_24813,N_24992);
or UO_755 (O_755,N_24960,N_24882);
nor UO_756 (O_756,N_24975,N_24866);
nor UO_757 (O_757,N_24957,N_24877);
xnor UO_758 (O_758,N_24987,N_24951);
xnor UO_759 (O_759,N_24965,N_24989);
and UO_760 (O_760,N_24873,N_24997);
or UO_761 (O_761,N_24878,N_24874);
and UO_762 (O_762,N_24909,N_24898);
xnor UO_763 (O_763,N_24944,N_24805);
nand UO_764 (O_764,N_24934,N_24847);
nand UO_765 (O_765,N_24802,N_24804);
xnor UO_766 (O_766,N_24829,N_24841);
nor UO_767 (O_767,N_24904,N_24806);
and UO_768 (O_768,N_24841,N_24917);
nor UO_769 (O_769,N_24961,N_24818);
nor UO_770 (O_770,N_24863,N_24819);
xor UO_771 (O_771,N_24866,N_24899);
nor UO_772 (O_772,N_24857,N_24872);
nand UO_773 (O_773,N_24999,N_24882);
xor UO_774 (O_774,N_24878,N_24932);
nor UO_775 (O_775,N_24827,N_24883);
nand UO_776 (O_776,N_24938,N_24942);
or UO_777 (O_777,N_24981,N_24918);
nand UO_778 (O_778,N_24815,N_24989);
nor UO_779 (O_779,N_24968,N_24987);
and UO_780 (O_780,N_24813,N_24984);
nor UO_781 (O_781,N_24872,N_24977);
or UO_782 (O_782,N_24853,N_24975);
nand UO_783 (O_783,N_24804,N_24885);
nor UO_784 (O_784,N_24884,N_24832);
nor UO_785 (O_785,N_24854,N_24869);
xor UO_786 (O_786,N_24936,N_24903);
or UO_787 (O_787,N_24832,N_24935);
or UO_788 (O_788,N_24841,N_24955);
xnor UO_789 (O_789,N_24935,N_24857);
nand UO_790 (O_790,N_24894,N_24983);
xor UO_791 (O_791,N_24964,N_24864);
nor UO_792 (O_792,N_24926,N_24968);
nand UO_793 (O_793,N_24960,N_24811);
or UO_794 (O_794,N_24942,N_24899);
nand UO_795 (O_795,N_24868,N_24924);
nand UO_796 (O_796,N_24848,N_24881);
or UO_797 (O_797,N_24936,N_24944);
nor UO_798 (O_798,N_24824,N_24836);
xor UO_799 (O_799,N_24801,N_24897);
nor UO_800 (O_800,N_24888,N_24947);
nand UO_801 (O_801,N_24963,N_24858);
and UO_802 (O_802,N_24924,N_24848);
xor UO_803 (O_803,N_24938,N_24807);
nor UO_804 (O_804,N_24950,N_24858);
or UO_805 (O_805,N_24860,N_24867);
nor UO_806 (O_806,N_24912,N_24956);
and UO_807 (O_807,N_24983,N_24863);
and UO_808 (O_808,N_24848,N_24884);
or UO_809 (O_809,N_24821,N_24816);
nand UO_810 (O_810,N_24839,N_24967);
nor UO_811 (O_811,N_24998,N_24899);
or UO_812 (O_812,N_24980,N_24927);
nand UO_813 (O_813,N_24980,N_24801);
nor UO_814 (O_814,N_24820,N_24864);
xor UO_815 (O_815,N_24836,N_24949);
nor UO_816 (O_816,N_24883,N_24908);
or UO_817 (O_817,N_24819,N_24858);
nor UO_818 (O_818,N_24925,N_24936);
and UO_819 (O_819,N_24814,N_24893);
and UO_820 (O_820,N_24803,N_24884);
nand UO_821 (O_821,N_24819,N_24920);
and UO_822 (O_822,N_24868,N_24884);
or UO_823 (O_823,N_24895,N_24987);
nand UO_824 (O_824,N_24901,N_24910);
nor UO_825 (O_825,N_24815,N_24809);
and UO_826 (O_826,N_24891,N_24913);
and UO_827 (O_827,N_24818,N_24946);
nand UO_828 (O_828,N_24848,N_24887);
nor UO_829 (O_829,N_24931,N_24802);
nor UO_830 (O_830,N_24835,N_24907);
and UO_831 (O_831,N_24941,N_24981);
nand UO_832 (O_832,N_24857,N_24971);
xor UO_833 (O_833,N_24924,N_24817);
and UO_834 (O_834,N_24931,N_24849);
nand UO_835 (O_835,N_24868,N_24881);
xnor UO_836 (O_836,N_24946,N_24879);
xnor UO_837 (O_837,N_24899,N_24803);
xor UO_838 (O_838,N_24974,N_24893);
and UO_839 (O_839,N_24975,N_24935);
nand UO_840 (O_840,N_24864,N_24982);
nor UO_841 (O_841,N_24855,N_24988);
and UO_842 (O_842,N_24878,N_24937);
and UO_843 (O_843,N_24941,N_24898);
xor UO_844 (O_844,N_24925,N_24861);
xnor UO_845 (O_845,N_24854,N_24805);
and UO_846 (O_846,N_24817,N_24981);
nand UO_847 (O_847,N_24919,N_24808);
nand UO_848 (O_848,N_24815,N_24817);
xnor UO_849 (O_849,N_24857,N_24838);
nand UO_850 (O_850,N_24821,N_24991);
nor UO_851 (O_851,N_24803,N_24822);
and UO_852 (O_852,N_24834,N_24898);
xor UO_853 (O_853,N_24839,N_24928);
and UO_854 (O_854,N_24852,N_24988);
xor UO_855 (O_855,N_24980,N_24943);
xor UO_856 (O_856,N_24807,N_24890);
nand UO_857 (O_857,N_24926,N_24928);
nand UO_858 (O_858,N_24929,N_24885);
and UO_859 (O_859,N_24857,N_24936);
xnor UO_860 (O_860,N_24992,N_24810);
xnor UO_861 (O_861,N_24833,N_24912);
xnor UO_862 (O_862,N_24866,N_24969);
or UO_863 (O_863,N_24927,N_24849);
xor UO_864 (O_864,N_24965,N_24837);
nor UO_865 (O_865,N_24955,N_24829);
nand UO_866 (O_866,N_24827,N_24952);
xnor UO_867 (O_867,N_24895,N_24844);
nor UO_868 (O_868,N_24898,N_24953);
nand UO_869 (O_869,N_24930,N_24866);
or UO_870 (O_870,N_24907,N_24928);
and UO_871 (O_871,N_24871,N_24811);
and UO_872 (O_872,N_24965,N_24831);
or UO_873 (O_873,N_24988,N_24854);
or UO_874 (O_874,N_24987,N_24825);
nand UO_875 (O_875,N_24803,N_24824);
xnor UO_876 (O_876,N_24808,N_24862);
xnor UO_877 (O_877,N_24886,N_24906);
xor UO_878 (O_878,N_24988,N_24857);
nor UO_879 (O_879,N_24901,N_24935);
nor UO_880 (O_880,N_24845,N_24821);
nor UO_881 (O_881,N_24929,N_24895);
and UO_882 (O_882,N_24870,N_24815);
or UO_883 (O_883,N_24903,N_24814);
nor UO_884 (O_884,N_24873,N_24915);
or UO_885 (O_885,N_24908,N_24845);
xor UO_886 (O_886,N_24904,N_24858);
or UO_887 (O_887,N_24806,N_24878);
nor UO_888 (O_888,N_24884,N_24857);
nor UO_889 (O_889,N_24862,N_24885);
nor UO_890 (O_890,N_24834,N_24848);
xnor UO_891 (O_891,N_24801,N_24901);
nor UO_892 (O_892,N_24978,N_24835);
xnor UO_893 (O_893,N_24981,N_24934);
nand UO_894 (O_894,N_24814,N_24972);
and UO_895 (O_895,N_24904,N_24957);
nand UO_896 (O_896,N_24868,N_24954);
and UO_897 (O_897,N_24902,N_24819);
nand UO_898 (O_898,N_24901,N_24897);
or UO_899 (O_899,N_24947,N_24871);
nand UO_900 (O_900,N_24910,N_24867);
nand UO_901 (O_901,N_24842,N_24800);
xor UO_902 (O_902,N_24922,N_24869);
nor UO_903 (O_903,N_24839,N_24956);
nor UO_904 (O_904,N_24997,N_24839);
xor UO_905 (O_905,N_24919,N_24848);
and UO_906 (O_906,N_24939,N_24870);
nand UO_907 (O_907,N_24824,N_24956);
xnor UO_908 (O_908,N_24915,N_24863);
nand UO_909 (O_909,N_24828,N_24845);
xor UO_910 (O_910,N_24885,N_24897);
or UO_911 (O_911,N_24920,N_24965);
and UO_912 (O_912,N_24902,N_24838);
nor UO_913 (O_913,N_24816,N_24943);
or UO_914 (O_914,N_24909,N_24899);
and UO_915 (O_915,N_24814,N_24982);
or UO_916 (O_916,N_24926,N_24829);
xor UO_917 (O_917,N_24923,N_24876);
xnor UO_918 (O_918,N_24838,N_24908);
xor UO_919 (O_919,N_24947,N_24889);
and UO_920 (O_920,N_24892,N_24933);
xor UO_921 (O_921,N_24814,N_24870);
xnor UO_922 (O_922,N_24843,N_24885);
and UO_923 (O_923,N_24978,N_24818);
or UO_924 (O_924,N_24868,N_24816);
xor UO_925 (O_925,N_24978,N_24945);
and UO_926 (O_926,N_24942,N_24873);
and UO_927 (O_927,N_24997,N_24935);
or UO_928 (O_928,N_24996,N_24997);
or UO_929 (O_929,N_24932,N_24881);
xnor UO_930 (O_930,N_24880,N_24897);
and UO_931 (O_931,N_24970,N_24853);
nor UO_932 (O_932,N_24822,N_24926);
xnor UO_933 (O_933,N_24871,N_24881);
nand UO_934 (O_934,N_24813,N_24926);
or UO_935 (O_935,N_24869,N_24956);
or UO_936 (O_936,N_24899,N_24848);
or UO_937 (O_937,N_24898,N_24907);
or UO_938 (O_938,N_24896,N_24826);
or UO_939 (O_939,N_24887,N_24830);
and UO_940 (O_940,N_24888,N_24838);
and UO_941 (O_941,N_24860,N_24901);
xor UO_942 (O_942,N_24843,N_24887);
and UO_943 (O_943,N_24859,N_24967);
and UO_944 (O_944,N_24830,N_24975);
nor UO_945 (O_945,N_24917,N_24921);
nor UO_946 (O_946,N_24816,N_24885);
or UO_947 (O_947,N_24892,N_24844);
nor UO_948 (O_948,N_24861,N_24830);
or UO_949 (O_949,N_24999,N_24840);
nand UO_950 (O_950,N_24833,N_24870);
or UO_951 (O_951,N_24967,N_24903);
or UO_952 (O_952,N_24972,N_24975);
nand UO_953 (O_953,N_24874,N_24951);
or UO_954 (O_954,N_24930,N_24846);
or UO_955 (O_955,N_24967,N_24883);
xor UO_956 (O_956,N_24907,N_24980);
xor UO_957 (O_957,N_24854,N_24995);
xor UO_958 (O_958,N_24950,N_24999);
xor UO_959 (O_959,N_24927,N_24868);
or UO_960 (O_960,N_24864,N_24996);
nor UO_961 (O_961,N_24825,N_24818);
xor UO_962 (O_962,N_24826,N_24970);
or UO_963 (O_963,N_24955,N_24960);
nand UO_964 (O_964,N_24964,N_24852);
or UO_965 (O_965,N_24924,N_24949);
and UO_966 (O_966,N_24926,N_24909);
nor UO_967 (O_967,N_24983,N_24893);
and UO_968 (O_968,N_24887,N_24870);
and UO_969 (O_969,N_24902,N_24839);
nor UO_970 (O_970,N_24948,N_24832);
and UO_971 (O_971,N_24903,N_24961);
or UO_972 (O_972,N_24972,N_24993);
or UO_973 (O_973,N_24997,N_24872);
nor UO_974 (O_974,N_24902,N_24893);
and UO_975 (O_975,N_24839,N_24854);
nand UO_976 (O_976,N_24820,N_24813);
xor UO_977 (O_977,N_24991,N_24871);
nor UO_978 (O_978,N_24944,N_24803);
nand UO_979 (O_979,N_24867,N_24875);
nor UO_980 (O_980,N_24826,N_24985);
and UO_981 (O_981,N_24911,N_24969);
and UO_982 (O_982,N_24845,N_24824);
nand UO_983 (O_983,N_24904,N_24821);
or UO_984 (O_984,N_24851,N_24970);
or UO_985 (O_985,N_24837,N_24832);
and UO_986 (O_986,N_24977,N_24925);
or UO_987 (O_987,N_24972,N_24857);
xnor UO_988 (O_988,N_24902,N_24932);
xnor UO_989 (O_989,N_24865,N_24844);
or UO_990 (O_990,N_24950,N_24870);
and UO_991 (O_991,N_24885,N_24800);
xnor UO_992 (O_992,N_24850,N_24870);
nor UO_993 (O_993,N_24869,N_24984);
nor UO_994 (O_994,N_24844,N_24987);
nor UO_995 (O_995,N_24891,N_24906);
or UO_996 (O_996,N_24805,N_24964);
and UO_997 (O_997,N_24826,N_24943);
and UO_998 (O_998,N_24831,N_24833);
xor UO_999 (O_999,N_24925,N_24960);
nand UO_1000 (O_1000,N_24823,N_24830);
xor UO_1001 (O_1001,N_24933,N_24978);
or UO_1002 (O_1002,N_24895,N_24930);
xor UO_1003 (O_1003,N_24868,N_24866);
xnor UO_1004 (O_1004,N_24990,N_24956);
xnor UO_1005 (O_1005,N_24966,N_24847);
nor UO_1006 (O_1006,N_24848,N_24991);
and UO_1007 (O_1007,N_24868,N_24987);
nand UO_1008 (O_1008,N_24890,N_24898);
nor UO_1009 (O_1009,N_24810,N_24936);
nor UO_1010 (O_1010,N_24825,N_24924);
nor UO_1011 (O_1011,N_24939,N_24845);
or UO_1012 (O_1012,N_24984,N_24938);
nand UO_1013 (O_1013,N_24961,N_24962);
or UO_1014 (O_1014,N_24958,N_24995);
nor UO_1015 (O_1015,N_24973,N_24909);
and UO_1016 (O_1016,N_24964,N_24935);
nor UO_1017 (O_1017,N_24845,N_24835);
or UO_1018 (O_1018,N_24990,N_24804);
nor UO_1019 (O_1019,N_24801,N_24948);
and UO_1020 (O_1020,N_24947,N_24913);
and UO_1021 (O_1021,N_24945,N_24915);
nor UO_1022 (O_1022,N_24947,N_24842);
xnor UO_1023 (O_1023,N_24810,N_24881);
nor UO_1024 (O_1024,N_24890,N_24811);
nand UO_1025 (O_1025,N_24963,N_24916);
and UO_1026 (O_1026,N_24879,N_24836);
xor UO_1027 (O_1027,N_24988,N_24864);
and UO_1028 (O_1028,N_24925,N_24824);
nand UO_1029 (O_1029,N_24855,N_24929);
xor UO_1030 (O_1030,N_24959,N_24879);
or UO_1031 (O_1031,N_24804,N_24801);
and UO_1032 (O_1032,N_24961,N_24824);
or UO_1033 (O_1033,N_24856,N_24997);
nand UO_1034 (O_1034,N_24939,N_24844);
nand UO_1035 (O_1035,N_24975,N_24849);
and UO_1036 (O_1036,N_24982,N_24873);
and UO_1037 (O_1037,N_24952,N_24880);
or UO_1038 (O_1038,N_24992,N_24804);
and UO_1039 (O_1039,N_24980,N_24863);
xnor UO_1040 (O_1040,N_24811,N_24831);
nand UO_1041 (O_1041,N_24855,N_24849);
and UO_1042 (O_1042,N_24925,N_24879);
or UO_1043 (O_1043,N_24930,N_24806);
or UO_1044 (O_1044,N_24951,N_24814);
nand UO_1045 (O_1045,N_24950,N_24969);
nor UO_1046 (O_1046,N_24965,N_24961);
or UO_1047 (O_1047,N_24968,N_24889);
and UO_1048 (O_1048,N_24958,N_24992);
nand UO_1049 (O_1049,N_24858,N_24890);
xnor UO_1050 (O_1050,N_24895,N_24973);
nand UO_1051 (O_1051,N_24996,N_24930);
xor UO_1052 (O_1052,N_24935,N_24819);
nor UO_1053 (O_1053,N_24966,N_24889);
nand UO_1054 (O_1054,N_24886,N_24990);
nand UO_1055 (O_1055,N_24941,N_24960);
nor UO_1056 (O_1056,N_24896,N_24968);
xnor UO_1057 (O_1057,N_24822,N_24927);
xor UO_1058 (O_1058,N_24940,N_24825);
nand UO_1059 (O_1059,N_24956,N_24946);
and UO_1060 (O_1060,N_24808,N_24855);
and UO_1061 (O_1061,N_24963,N_24832);
nand UO_1062 (O_1062,N_24926,N_24993);
nor UO_1063 (O_1063,N_24876,N_24886);
xor UO_1064 (O_1064,N_24964,N_24838);
and UO_1065 (O_1065,N_24962,N_24878);
and UO_1066 (O_1066,N_24901,N_24840);
xor UO_1067 (O_1067,N_24817,N_24824);
nor UO_1068 (O_1068,N_24939,N_24964);
nand UO_1069 (O_1069,N_24987,N_24851);
nand UO_1070 (O_1070,N_24910,N_24945);
nand UO_1071 (O_1071,N_24999,N_24939);
nand UO_1072 (O_1072,N_24961,N_24800);
nor UO_1073 (O_1073,N_24856,N_24855);
or UO_1074 (O_1074,N_24869,N_24848);
or UO_1075 (O_1075,N_24871,N_24986);
nor UO_1076 (O_1076,N_24838,N_24891);
nor UO_1077 (O_1077,N_24869,N_24831);
nor UO_1078 (O_1078,N_24806,N_24884);
nand UO_1079 (O_1079,N_24925,N_24974);
and UO_1080 (O_1080,N_24911,N_24895);
nand UO_1081 (O_1081,N_24800,N_24857);
or UO_1082 (O_1082,N_24999,N_24803);
xor UO_1083 (O_1083,N_24934,N_24803);
nand UO_1084 (O_1084,N_24983,N_24895);
nor UO_1085 (O_1085,N_24982,N_24863);
nand UO_1086 (O_1086,N_24932,N_24952);
or UO_1087 (O_1087,N_24928,N_24804);
nor UO_1088 (O_1088,N_24986,N_24962);
xnor UO_1089 (O_1089,N_24900,N_24985);
or UO_1090 (O_1090,N_24989,N_24951);
or UO_1091 (O_1091,N_24988,N_24817);
or UO_1092 (O_1092,N_24860,N_24976);
xnor UO_1093 (O_1093,N_24812,N_24922);
and UO_1094 (O_1094,N_24996,N_24820);
or UO_1095 (O_1095,N_24893,N_24930);
and UO_1096 (O_1096,N_24952,N_24860);
xnor UO_1097 (O_1097,N_24831,N_24920);
nor UO_1098 (O_1098,N_24882,N_24872);
nor UO_1099 (O_1099,N_24897,N_24920);
or UO_1100 (O_1100,N_24994,N_24938);
or UO_1101 (O_1101,N_24884,N_24804);
xor UO_1102 (O_1102,N_24908,N_24871);
xnor UO_1103 (O_1103,N_24844,N_24920);
xnor UO_1104 (O_1104,N_24809,N_24876);
or UO_1105 (O_1105,N_24870,N_24892);
nand UO_1106 (O_1106,N_24996,N_24986);
or UO_1107 (O_1107,N_24992,N_24801);
and UO_1108 (O_1108,N_24916,N_24819);
nor UO_1109 (O_1109,N_24854,N_24993);
xor UO_1110 (O_1110,N_24954,N_24974);
nand UO_1111 (O_1111,N_24832,N_24868);
xnor UO_1112 (O_1112,N_24820,N_24938);
xnor UO_1113 (O_1113,N_24863,N_24858);
and UO_1114 (O_1114,N_24808,N_24841);
nor UO_1115 (O_1115,N_24923,N_24922);
and UO_1116 (O_1116,N_24816,N_24901);
or UO_1117 (O_1117,N_24952,N_24924);
and UO_1118 (O_1118,N_24998,N_24957);
nor UO_1119 (O_1119,N_24801,N_24856);
or UO_1120 (O_1120,N_24847,N_24997);
and UO_1121 (O_1121,N_24907,N_24832);
and UO_1122 (O_1122,N_24877,N_24964);
nor UO_1123 (O_1123,N_24838,N_24939);
and UO_1124 (O_1124,N_24838,N_24959);
and UO_1125 (O_1125,N_24968,N_24964);
nand UO_1126 (O_1126,N_24985,N_24870);
and UO_1127 (O_1127,N_24830,N_24878);
nor UO_1128 (O_1128,N_24906,N_24828);
and UO_1129 (O_1129,N_24824,N_24927);
xnor UO_1130 (O_1130,N_24901,N_24889);
or UO_1131 (O_1131,N_24929,N_24850);
nor UO_1132 (O_1132,N_24807,N_24985);
and UO_1133 (O_1133,N_24987,N_24854);
nor UO_1134 (O_1134,N_24923,N_24861);
and UO_1135 (O_1135,N_24985,N_24945);
nor UO_1136 (O_1136,N_24885,N_24878);
nor UO_1137 (O_1137,N_24949,N_24874);
nand UO_1138 (O_1138,N_24968,N_24973);
and UO_1139 (O_1139,N_24886,N_24977);
nand UO_1140 (O_1140,N_24838,N_24936);
xnor UO_1141 (O_1141,N_24836,N_24826);
or UO_1142 (O_1142,N_24873,N_24893);
or UO_1143 (O_1143,N_24914,N_24834);
xnor UO_1144 (O_1144,N_24902,N_24948);
nand UO_1145 (O_1145,N_24941,N_24912);
and UO_1146 (O_1146,N_24836,N_24886);
nand UO_1147 (O_1147,N_24831,N_24828);
nand UO_1148 (O_1148,N_24932,N_24866);
or UO_1149 (O_1149,N_24873,N_24813);
nand UO_1150 (O_1150,N_24978,N_24929);
nand UO_1151 (O_1151,N_24906,N_24846);
nand UO_1152 (O_1152,N_24853,N_24960);
xnor UO_1153 (O_1153,N_24955,N_24821);
or UO_1154 (O_1154,N_24981,N_24888);
or UO_1155 (O_1155,N_24879,N_24804);
nand UO_1156 (O_1156,N_24820,N_24966);
nor UO_1157 (O_1157,N_24920,N_24896);
xor UO_1158 (O_1158,N_24800,N_24827);
and UO_1159 (O_1159,N_24932,N_24968);
nand UO_1160 (O_1160,N_24951,N_24892);
xnor UO_1161 (O_1161,N_24870,N_24893);
or UO_1162 (O_1162,N_24926,N_24985);
or UO_1163 (O_1163,N_24919,N_24991);
or UO_1164 (O_1164,N_24838,N_24880);
xnor UO_1165 (O_1165,N_24916,N_24892);
xnor UO_1166 (O_1166,N_24801,N_24815);
xnor UO_1167 (O_1167,N_24916,N_24865);
and UO_1168 (O_1168,N_24871,N_24970);
nor UO_1169 (O_1169,N_24881,N_24941);
xor UO_1170 (O_1170,N_24837,N_24847);
nand UO_1171 (O_1171,N_24913,N_24852);
nand UO_1172 (O_1172,N_24911,N_24821);
or UO_1173 (O_1173,N_24826,N_24919);
and UO_1174 (O_1174,N_24810,N_24932);
nor UO_1175 (O_1175,N_24856,N_24950);
nor UO_1176 (O_1176,N_24952,N_24950);
xnor UO_1177 (O_1177,N_24846,N_24998);
nand UO_1178 (O_1178,N_24824,N_24991);
or UO_1179 (O_1179,N_24818,N_24812);
nor UO_1180 (O_1180,N_24863,N_24903);
or UO_1181 (O_1181,N_24867,N_24811);
nor UO_1182 (O_1182,N_24966,N_24860);
nor UO_1183 (O_1183,N_24992,N_24875);
and UO_1184 (O_1184,N_24932,N_24911);
nand UO_1185 (O_1185,N_24826,N_24846);
nor UO_1186 (O_1186,N_24864,N_24983);
nor UO_1187 (O_1187,N_24956,N_24866);
xor UO_1188 (O_1188,N_24857,N_24839);
xor UO_1189 (O_1189,N_24809,N_24896);
xor UO_1190 (O_1190,N_24935,N_24931);
nand UO_1191 (O_1191,N_24990,N_24831);
nand UO_1192 (O_1192,N_24899,N_24926);
xor UO_1193 (O_1193,N_24979,N_24982);
or UO_1194 (O_1194,N_24900,N_24831);
and UO_1195 (O_1195,N_24860,N_24832);
xnor UO_1196 (O_1196,N_24947,N_24997);
nand UO_1197 (O_1197,N_24928,N_24810);
and UO_1198 (O_1198,N_24817,N_24999);
xor UO_1199 (O_1199,N_24954,N_24957);
or UO_1200 (O_1200,N_24879,N_24921);
nor UO_1201 (O_1201,N_24920,N_24867);
nand UO_1202 (O_1202,N_24839,N_24832);
or UO_1203 (O_1203,N_24859,N_24953);
and UO_1204 (O_1204,N_24992,N_24925);
xnor UO_1205 (O_1205,N_24802,N_24896);
or UO_1206 (O_1206,N_24907,N_24998);
or UO_1207 (O_1207,N_24962,N_24996);
and UO_1208 (O_1208,N_24838,N_24865);
xor UO_1209 (O_1209,N_24982,N_24879);
nor UO_1210 (O_1210,N_24806,N_24892);
or UO_1211 (O_1211,N_24953,N_24931);
or UO_1212 (O_1212,N_24899,N_24911);
nand UO_1213 (O_1213,N_24855,N_24913);
and UO_1214 (O_1214,N_24930,N_24857);
and UO_1215 (O_1215,N_24867,N_24930);
or UO_1216 (O_1216,N_24808,N_24852);
or UO_1217 (O_1217,N_24976,N_24871);
nor UO_1218 (O_1218,N_24807,N_24970);
and UO_1219 (O_1219,N_24889,N_24864);
xnor UO_1220 (O_1220,N_24815,N_24958);
xnor UO_1221 (O_1221,N_24922,N_24856);
nand UO_1222 (O_1222,N_24902,N_24922);
or UO_1223 (O_1223,N_24810,N_24896);
xor UO_1224 (O_1224,N_24997,N_24877);
or UO_1225 (O_1225,N_24970,N_24930);
nand UO_1226 (O_1226,N_24876,N_24971);
or UO_1227 (O_1227,N_24868,N_24949);
and UO_1228 (O_1228,N_24813,N_24988);
nor UO_1229 (O_1229,N_24928,N_24952);
nor UO_1230 (O_1230,N_24934,N_24867);
nand UO_1231 (O_1231,N_24943,N_24945);
and UO_1232 (O_1232,N_24853,N_24845);
and UO_1233 (O_1233,N_24984,N_24958);
xnor UO_1234 (O_1234,N_24841,N_24896);
xnor UO_1235 (O_1235,N_24863,N_24899);
nand UO_1236 (O_1236,N_24973,N_24923);
nor UO_1237 (O_1237,N_24985,N_24879);
xor UO_1238 (O_1238,N_24969,N_24982);
or UO_1239 (O_1239,N_24826,N_24802);
or UO_1240 (O_1240,N_24846,N_24821);
xor UO_1241 (O_1241,N_24970,N_24922);
or UO_1242 (O_1242,N_24890,N_24815);
or UO_1243 (O_1243,N_24856,N_24925);
or UO_1244 (O_1244,N_24825,N_24967);
xnor UO_1245 (O_1245,N_24830,N_24948);
xnor UO_1246 (O_1246,N_24982,N_24816);
or UO_1247 (O_1247,N_24919,N_24818);
and UO_1248 (O_1248,N_24983,N_24926);
nor UO_1249 (O_1249,N_24991,N_24986);
or UO_1250 (O_1250,N_24915,N_24819);
nor UO_1251 (O_1251,N_24977,N_24825);
nor UO_1252 (O_1252,N_24888,N_24847);
xnor UO_1253 (O_1253,N_24945,N_24839);
nand UO_1254 (O_1254,N_24918,N_24971);
nand UO_1255 (O_1255,N_24861,N_24857);
or UO_1256 (O_1256,N_24986,N_24933);
and UO_1257 (O_1257,N_24841,N_24951);
xor UO_1258 (O_1258,N_24904,N_24969);
or UO_1259 (O_1259,N_24868,N_24858);
and UO_1260 (O_1260,N_24964,N_24818);
nor UO_1261 (O_1261,N_24845,N_24868);
xnor UO_1262 (O_1262,N_24884,N_24898);
nor UO_1263 (O_1263,N_24814,N_24839);
and UO_1264 (O_1264,N_24954,N_24873);
and UO_1265 (O_1265,N_24866,N_24963);
xor UO_1266 (O_1266,N_24909,N_24821);
nor UO_1267 (O_1267,N_24861,N_24995);
nor UO_1268 (O_1268,N_24910,N_24891);
nor UO_1269 (O_1269,N_24830,N_24801);
xnor UO_1270 (O_1270,N_24811,N_24878);
nand UO_1271 (O_1271,N_24803,N_24886);
or UO_1272 (O_1272,N_24969,N_24845);
or UO_1273 (O_1273,N_24831,N_24893);
and UO_1274 (O_1274,N_24863,N_24804);
or UO_1275 (O_1275,N_24883,N_24944);
and UO_1276 (O_1276,N_24881,N_24939);
xor UO_1277 (O_1277,N_24966,N_24900);
and UO_1278 (O_1278,N_24996,N_24892);
xnor UO_1279 (O_1279,N_24817,N_24855);
and UO_1280 (O_1280,N_24942,N_24841);
and UO_1281 (O_1281,N_24827,N_24974);
and UO_1282 (O_1282,N_24827,N_24865);
or UO_1283 (O_1283,N_24976,N_24986);
nand UO_1284 (O_1284,N_24875,N_24832);
nand UO_1285 (O_1285,N_24960,N_24877);
nor UO_1286 (O_1286,N_24854,N_24904);
and UO_1287 (O_1287,N_24822,N_24952);
and UO_1288 (O_1288,N_24801,N_24812);
nand UO_1289 (O_1289,N_24940,N_24902);
or UO_1290 (O_1290,N_24812,N_24824);
nand UO_1291 (O_1291,N_24964,N_24881);
xor UO_1292 (O_1292,N_24963,N_24945);
nor UO_1293 (O_1293,N_24897,N_24809);
and UO_1294 (O_1294,N_24881,N_24965);
nand UO_1295 (O_1295,N_24850,N_24965);
nor UO_1296 (O_1296,N_24898,N_24956);
nand UO_1297 (O_1297,N_24853,N_24999);
nand UO_1298 (O_1298,N_24813,N_24882);
xnor UO_1299 (O_1299,N_24814,N_24965);
nand UO_1300 (O_1300,N_24964,N_24861);
nand UO_1301 (O_1301,N_24828,N_24873);
nor UO_1302 (O_1302,N_24822,N_24957);
xor UO_1303 (O_1303,N_24944,N_24907);
xnor UO_1304 (O_1304,N_24951,N_24870);
xnor UO_1305 (O_1305,N_24969,N_24966);
and UO_1306 (O_1306,N_24980,N_24987);
or UO_1307 (O_1307,N_24806,N_24818);
nor UO_1308 (O_1308,N_24824,N_24905);
xor UO_1309 (O_1309,N_24814,N_24897);
and UO_1310 (O_1310,N_24852,N_24849);
nand UO_1311 (O_1311,N_24989,N_24929);
and UO_1312 (O_1312,N_24930,N_24922);
or UO_1313 (O_1313,N_24910,N_24982);
nand UO_1314 (O_1314,N_24841,N_24935);
and UO_1315 (O_1315,N_24916,N_24982);
nand UO_1316 (O_1316,N_24980,N_24860);
nor UO_1317 (O_1317,N_24801,N_24883);
xor UO_1318 (O_1318,N_24801,N_24952);
xor UO_1319 (O_1319,N_24846,N_24945);
xor UO_1320 (O_1320,N_24906,N_24892);
nand UO_1321 (O_1321,N_24844,N_24902);
or UO_1322 (O_1322,N_24874,N_24858);
nor UO_1323 (O_1323,N_24886,N_24825);
xor UO_1324 (O_1324,N_24994,N_24987);
or UO_1325 (O_1325,N_24806,N_24942);
or UO_1326 (O_1326,N_24806,N_24845);
nor UO_1327 (O_1327,N_24940,N_24863);
or UO_1328 (O_1328,N_24950,N_24998);
xor UO_1329 (O_1329,N_24818,N_24908);
and UO_1330 (O_1330,N_24806,N_24946);
or UO_1331 (O_1331,N_24903,N_24988);
xor UO_1332 (O_1332,N_24834,N_24875);
or UO_1333 (O_1333,N_24916,N_24852);
and UO_1334 (O_1334,N_24995,N_24999);
nor UO_1335 (O_1335,N_24854,N_24974);
nand UO_1336 (O_1336,N_24953,N_24849);
nor UO_1337 (O_1337,N_24851,N_24809);
and UO_1338 (O_1338,N_24990,N_24857);
nand UO_1339 (O_1339,N_24853,N_24804);
xnor UO_1340 (O_1340,N_24899,N_24806);
nor UO_1341 (O_1341,N_24910,N_24856);
nand UO_1342 (O_1342,N_24840,N_24929);
or UO_1343 (O_1343,N_24830,N_24918);
nand UO_1344 (O_1344,N_24814,N_24990);
nand UO_1345 (O_1345,N_24884,N_24935);
nor UO_1346 (O_1346,N_24999,N_24922);
and UO_1347 (O_1347,N_24952,N_24851);
and UO_1348 (O_1348,N_24975,N_24991);
xor UO_1349 (O_1349,N_24898,N_24984);
nand UO_1350 (O_1350,N_24902,N_24960);
and UO_1351 (O_1351,N_24870,N_24848);
and UO_1352 (O_1352,N_24946,N_24864);
or UO_1353 (O_1353,N_24915,N_24826);
and UO_1354 (O_1354,N_24836,N_24984);
or UO_1355 (O_1355,N_24863,N_24822);
and UO_1356 (O_1356,N_24824,N_24984);
or UO_1357 (O_1357,N_24891,N_24812);
nand UO_1358 (O_1358,N_24967,N_24925);
xor UO_1359 (O_1359,N_24912,N_24802);
or UO_1360 (O_1360,N_24876,N_24814);
nor UO_1361 (O_1361,N_24887,N_24941);
nand UO_1362 (O_1362,N_24950,N_24915);
nor UO_1363 (O_1363,N_24938,N_24923);
and UO_1364 (O_1364,N_24816,N_24941);
nand UO_1365 (O_1365,N_24889,N_24931);
xor UO_1366 (O_1366,N_24951,N_24855);
or UO_1367 (O_1367,N_24936,N_24872);
and UO_1368 (O_1368,N_24902,N_24870);
nand UO_1369 (O_1369,N_24804,N_24984);
nand UO_1370 (O_1370,N_24813,N_24914);
nand UO_1371 (O_1371,N_24842,N_24803);
and UO_1372 (O_1372,N_24810,N_24968);
or UO_1373 (O_1373,N_24852,N_24822);
xor UO_1374 (O_1374,N_24882,N_24801);
nor UO_1375 (O_1375,N_24944,N_24880);
or UO_1376 (O_1376,N_24933,N_24962);
or UO_1377 (O_1377,N_24956,N_24868);
nand UO_1378 (O_1378,N_24895,N_24976);
nand UO_1379 (O_1379,N_24912,N_24997);
and UO_1380 (O_1380,N_24834,N_24923);
nor UO_1381 (O_1381,N_24960,N_24824);
and UO_1382 (O_1382,N_24957,N_24958);
and UO_1383 (O_1383,N_24862,N_24968);
or UO_1384 (O_1384,N_24916,N_24811);
nor UO_1385 (O_1385,N_24863,N_24913);
and UO_1386 (O_1386,N_24861,N_24858);
nor UO_1387 (O_1387,N_24800,N_24810);
nor UO_1388 (O_1388,N_24818,N_24859);
and UO_1389 (O_1389,N_24841,N_24822);
and UO_1390 (O_1390,N_24927,N_24917);
nor UO_1391 (O_1391,N_24939,N_24866);
and UO_1392 (O_1392,N_24956,N_24982);
and UO_1393 (O_1393,N_24895,N_24974);
nand UO_1394 (O_1394,N_24860,N_24885);
xnor UO_1395 (O_1395,N_24807,N_24855);
and UO_1396 (O_1396,N_24875,N_24962);
xnor UO_1397 (O_1397,N_24888,N_24916);
or UO_1398 (O_1398,N_24985,N_24855);
or UO_1399 (O_1399,N_24959,N_24934);
and UO_1400 (O_1400,N_24898,N_24937);
xnor UO_1401 (O_1401,N_24835,N_24935);
nor UO_1402 (O_1402,N_24953,N_24956);
nor UO_1403 (O_1403,N_24977,N_24948);
nor UO_1404 (O_1404,N_24888,N_24942);
and UO_1405 (O_1405,N_24888,N_24878);
and UO_1406 (O_1406,N_24886,N_24848);
and UO_1407 (O_1407,N_24960,N_24970);
xor UO_1408 (O_1408,N_24802,N_24880);
or UO_1409 (O_1409,N_24902,N_24887);
nand UO_1410 (O_1410,N_24909,N_24890);
nor UO_1411 (O_1411,N_24941,N_24809);
xnor UO_1412 (O_1412,N_24843,N_24845);
nor UO_1413 (O_1413,N_24874,N_24879);
or UO_1414 (O_1414,N_24907,N_24869);
nor UO_1415 (O_1415,N_24904,N_24827);
and UO_1416 (O_1416,N_24870,N_24969);
xnor UO_1417 (O_1417,N_24914,N_24806);
xnor UO_1418 (O_1418,N_24832,N_24881);
and UO_1419 (O_1419,N_24954,N_24980);
xor UO_1420 (O_1420,N_24849,N_24867);
or UO_1421 (O_1421,N_24921,N_24886);
nor UO_1422 (O_1422,N_24877,N_24870);
nand UO_1423 (O_1423,N_24977,N_24845);
or UO_1424 (O_1424,N_24930,N_24981);
nand UO_1425 (O_1425,N_24903,N_24829);
nor UO_1426 (O_1426,N_24826,N_24949);
nor UO_1427 (O_1427,N_24827,N_24908);
nor UO_1428 (O_1428,N_24941,N_24891);
nand UO_1429 (O_1429,N_24822,N_24832);
or UO_1430 (O_1430,N_24812,N_24949);
and UO_1431 (O_1431,N_24940,N_24896);
xnor UO_1432 (O_1432,N_24829,N_24947);
nand UO_1433 (O_1433,N_24956,N_24928);
or UO_1434 (O_1434,N_24832,N_24823);
or UO_1435 (O_1435,N_24813,N_24933);
or UO_1436 (O_1436,N_24944,N_24821);
and UO_1437 (O_1437,N_24875,N_24801);
nor UO_1438 (O_1438,N_24964,N_24965);
nor UO_1439 (O_1439,N_24919,N_24800);
or UO_1440 (O_1440,N_24945,N_24968);
or UO_1441 (O_1441,N_24930,N_24954);
and UO_1442 (O_1442,N_24879,N_24940);
nor UO_1443 (O_1443,N_24911,N_24832);
or UO_1444 (O_1444,N_24891,N_24840);
nand UO_1445 (O_1445,N_24927,N_24924);
xor UO_1446 (O_1446,N_24934,N_24879);
nor UO_1447 (O_1447,N_24907,N_24818);
xor UO_1448 (O_1448,N_24998,N_24919);
or UO_1449 (O_1449,N_24938,N_24989);
and UO_1450 (O_1450,N_24852,N_24812);
and UO_1451 (O_1451,N_24979,N_24913);
nand UO_1452 (O_1452,N_24802,N_24809);
xor UO_1453 (O_1453,N_24830,N_24847);
and UO_1454 (O_1454,N_24850,N_24800);
or UO_1455 (O_1455,N_24840,N_24950);
and UO_1456 (O_1456,N_24824,N_24938);
xnor UO_1457 (O_1457,N_24949,N_24927);
nand UO_1458 (O_1458,N_24851,N_24960);
nor UO_1459 (O_1459,N_24917,N_24924);
xnor UO_1460 (O_1460,N_24836,N_24800);
nor UO_1461 (O_1461,N_24868,N_24926);
or UO_1462 (O_1462,N_24966,N_24879);
nand UO_1463 (O_1463,N_24966,N_24814);
nor UO_1464 (O_1464,N_24920,N_24873);
nor UO_1465 (O_1465,N_24962,N_24949);
or UO_1466 (O_1466,N_24991,N_24926);
nor UO_1467 (O_1467,N_24978,N_24870);
xnor UO_1468 (O_1468,N_24817,N_24900);
nand UO_1469 (O_1469,N_24852,N_24898);
nor UO_1470 (O_1470,N_24844,N_24904);
and UO_1471 (O_1471,N_24897,N_24856);
xor UO_1472 (O_1472,N_24990,N_24977);
or UO_1473 (O_1473,N_24982,N_24973);
and UO_1474 (O_1474,N_24898,N_24893);
nor UO_1475 (O_1475,N_24905,N_24870);
and UO_1476 (O_1476,N_24888,N_24959);
nand UO_1477 (O_1477,N_24812,N_24831);
xnor UO_1478 (O_1478,N_24943,N_24896);
and UO_1479 (O_1479,N_24826,N_24903);
xor UO_1480 (O_1480,N_24819,N_24865);
nor UO_1481 (O_1481,N_24806,N_24813);
xnor UO_1482 (O_1482,N_24986,N_24805);
and UO_1483 (O_1483,N_24954,N_24858);
or UO_1484 (O_1484,N_24924,N_24857);
nor UO_1485 (O_1485,N_24876,N_24973);
or UO_1486 (O_1486,N_24880,N_24850);
or UO_1487 (O_1487,N_24995,N_24872);
nand UO_1488 (O_1488,N_24831,N_24819);
xnor UO_1489 (O_1489,N_24818,N_24820);
or UO_1490 (O_1490,N_24886,N_24885);
nand UO_1491 (O_1491,N_24872,N_24920);
nand UO_1492 (O_1492,N_24941,N_24827);
nor UO_1493 (O_1493,N_24959,N_24890);
nor UO_1494 (O_1494,N_24954,N_24857);
and UO_1495 (O_1495,N_24859,N_24958);
and UO_1496 (O_1496,N_24829,N_24983);
nand UO_1497 (O_1497,N_24988,N_24875);
nor UO_1498 (O_1498,N_24933,N_24918);
xnor UO_1499 (O_1499,N_24852,N_24874);
xnor UO_1500 (O_1500,N_24813,N_24875);
nand UO_1501 (O_1501,N_24811,N_24857);
or UO_1502 (O_1502,N_24901,N_24872);
nand UO_1503 (O_1503,N_24817,N_24998);
or UO_1504 (O_1504,N_24933,N_24989);
xnor UO_1505 (O_1505,N_24931,N_24833);
or UO_1506 (O_1506,N_24833,N_24945);
or UO_1507 (O_1507,N_24800,N_24846);
nand UO_1508 (O_1508,N_24968,N_24979);
or UO_1509 (O_1509,N_24979,N_24861);
nand UO_1510 (O_1510,N_24894,N_24837);
or UO_1511 (O_1511,N_24988,N_24837);
and UO_1512 (O_1512,N_24914,N_24886);
nand UO_1513 (O_1513,N_24895,N_24945);
nor UO_1514 (O_1514,N_24963,N_24967);
xnor UO_1515 (O_1515,N_24852,N_24807);
nand UO_1516 (O_1516,N_24913,N_24829);
xnor UO_1517 (O_1517,N_24959,N_24964);
nand UO_1518 (O_1518,N_24903,N_24873);
nor UO_1519 (O_1519,N_24903,N_24803);
nand UO_1520 (O_1520,N_24921,N_24872);
xnor UO_1521 (O_1521,N_24922,N_24808);
or UO_1522 (O_1522,N_24848,N_24916);
or UO_1523 (O_1523,N_24835,N_24985);
nand UO_1524 (O_1524,N_24848,N_24873);
nor UO_1525 (O_1525,N_24869,N_24859);
and UO_1526 (O_1526,N_24919,N_24891);
xor UO_1527 (O_1527,N_24886,N_24915);
or UO_1528 (O_1528,N_24948,N_24995);
nand UO_1529 (O_1529,N_24963,N_24830);
and UO_1530 (O_1530,N_24981,N_24989);
nor UO_1531 (O_1531,N_24940,N_24967);
or UO_1532 (O_1532,N_24992,N_24946);
nor UO_1533 (O_1533,N_24948,N_24846);
nor UO_1534 (O_1534,N_24990,N_24941);
xor UO_1535 (O_1535,N_24899,N_24960);
nor UO_1536 (O_1536,N_24913,N_24982);
and UO_1537 (O_1537,N_24880,N_24876);
nand UO_1538 (O_1538,N_24821,N_24936);
nand UO_1539 (O_1539,N_24911,N_24977);
or UO_1540 (O_1540,N_24902,N_24871);
nand UO_1541 (O_1541,N_24913,N_24822);
xor UO_1542 (O_1542,N_24873,N_24871);
xnor UO_1543 (O_1543,N_24827,N_24937);
nand UO_1544 (O_1544,N_24962,N_24959);
nor UO_1545 (O_1545,N_24900,N_24871);
nor UO_1546 (O_1546,N_24843,N_24940);
or UO_1547 (O_1547,N_24816,N_24946);
xnor UO_1548 (O_1548,N_24922,N_24851);
and UO_1549 (O_1549,N_24985,N_24954);
nand UO_1550 (O_1550,N_24834,N_24978);
nand UO_1551 (O_1551,N_24816,N_24953);
nand UO_1552 (O_1552,N_24929,N_24881);
nand UO_1553 (O_1553,N_24928,N_24831);
or UO_1554 (O_1554,N_24900,N_24976);
xor UO_1555 (O_1555,N_24952,N_24939);
and UO_1556 (O_1556,N_24953,N_24982);
nor UO_1557 (O_1557,N_24912,N_24873);
and UO_1558 (O_1558,N_24867,N_24950);
and UO_1559 (O_1559,N_24936,N_24919);
and UO_1560 (O_1560,N_24930,N_24887);
nor UO_1561 (O_1561,N_24932,N_24844);
nand UO_1562 (O_1562,N_24932,N_24985);
nand UO_1563 (O_1563,N_24995,N_24904);
xnor UO_1564 (O_1564,N_24989,N_24816);
xor UO_1565 (O_1565,N_24926,N_24816);
nand UO_1566 (O_1566,N_24986,N_24821);
nand UO_1567 (O_1567,N_24949,N_24910);
or UO_1568 (O_1568,N_24821,N_24806);
or UO_1569 (O_1569,N_24951,N_24879);
nor UO_1570 (O_1570,N_24807,N_24934);
nand UO_1571 (O_1571,N_24843,N_24979);
or UO_1572 (O_1572,N_24909,N_24943);
nor UO_1573 (O_1573,N_24843,N_24911);
xnor UO_1574 (O_1574,N_24838,N_24943);
nor UO_1575 (O_1575,N_24898,N_24983);
nand UO_1576 (O_1576,N_24946,N_24853);
nand UO_1577 (O_1577,N_24907,N_24917);
nand UO_1578 (O_1578,N_24827,N_24903);
and UO_1579 (O_1579,N_24930,N_24915);
or UO_1580 (O_1580,N_24949,N_24875);
and UO_1581 (O_1581,N_24974,N_24826);
xor UO_1582 (O_1582,N_24975,N_24973);
or UO_1583 (O_1583,N_24874,N_24871);
nor UO_1584 (O_1584,N_24901,N_24861);
nor UO_1585 (O_1585,N_24950,N_24993);
or UO_1586 (O_1586,N_24896,N_24969);
or UO_1587 (O_1587,N_24903,N_24861);
nand UO_1588 (O_1588,N_24942,N_24839);
nand UO_1589 (O_1589,N_24817,N_24854);
xor UO_1590 (O_1590,N_24907,N_24810);
nand UO_1591 (O_1591,N_24838,N_24819);
and UO_1592 (O_1592,N_24935,N_24979);
nand UO_1593 (O_1593,N_24875,N_24936);
nand UO_1594 (O_1594,N_24889,N_24927);
nand UO_1595 (O_1595,N_24814,N_24911);
nor UO_1596 (O_1596,N_24911,N_24976);
or UO_1597 (O_1597,N_24820,N_24907);
and UO_1598 (O_1598,N_24829,N_24871);
and UO_1599 (O_1599,N_24850,N_24852);
nand UO_1600 (O_1600,N_24822,N_24839);
nand UO_1601 (O_1601,N_24860,N_24981);
nand UO_1602 (O_1602,N_24904,N_24896);
nand UO_1603 (O_1603,N_24913,N_24844);
xnor UO_1604 (O_1604,N_24973,N_24856);
or UO_1605 (O_1605,N_24833,N_24908);
nand UO_1606 (O_1606,N_24879,N_24832);
nor UO_1607 (O_1607,N_24851,N_24816);
nor UO_1608 (O_1608,N_24961,N_24909);
and UO_1609 (O_1609,N_24927,N_24829);
xnor UO_1610 (O_1610,N_24967,N_24923);
xnor UO_1611 (O_1611,N_24843,N_24958);
nor UO_1612 (O_1612,N_24981,N_24956);
or UO_1613 (O_1613,N_24871,N_24890);
nor UO_1614 (O_1614,N_24915,N_24860);
or UO_1615 (O_1615,N_24808,N_24976);
and UO_1616 (O_1616,N_24979,N_24909);
and UO_1617 (O_1617,N_24820,N_24869);
or UO_1618 (O_1618,N_24824,N_24823);
or UO_1619 (O_1619,N_24958,N_24864);
and UO_1620 (O_1620,N_24834,N_24861);
xor UO_1621 (O_1621,N_24942,N_24937);
and UO_1622 (O_1622,N_24855,N_24896);
and UO_1623 (O_1623,N_24971,N_24970);
xor UO_1624 (O_1624,N_24857,N_24814);
xnor UO_1625 (O_1625,N_24922,N_24824);
and UO_1626 (O_1626,N_24800,N_24914);
nand UO_1627 (O_1627,N_24992,N_24990);
nand UO_1628 (O_1628,N_24995,N_24911);
and UO_1629 (O_1629,N_24904,N_24967);
and UO_1630 (O_1630,N_24979,N_24898);
nor UO_1631 (O_1631,N_24852,N_24840);
or UO_1632 (O_1632,N_24975,N_24827);
xnor UO_1633 (O_1633,N_24880,N_24853);
and UO_1634 (O_1634,N_24922,N_24834);
or UO_1635 (O_1635,N_24925,N_24832);
nand UO_1636 (O_1636,N_24851,N_24912);
nand UO_1637 (O_1637,N_24852,N_24885);
or UO_1638 (O_1638,N_24998,N_24909);
nor UO_1639 (O_1639,N_24943,N_24934);
nor UO_1640 (O_1640,N_24987,N_24926);
xnor UO_1641 (O_1641,N_24811,N_24978);
nand UO_1642 (O_1642,N_24980,N_24874);
or UO_1643 (O_1643,N_24950,N_24912);
or UO_1644 (O_1644,N_24800,N_24932);
or UO_1645 (O_1645,N_24883,N_24859);
nor UO_1646 (O_1646,N_24918,N_24991);
and UO_1647 (O_1647,N_24977,N_24812);
nand UO_1648 (O_1648,N_24871,N_24843);
nor UO_1649 (O_1649,N_24810,N_24825);
xnor UO_1650 (O_1650,N_24890,N_24865);
xor UO_1651 (O_1651,N_24899,N_24925);
and UO_1652 (O_1652,N_24882,N_24916);
or UO_1653 (O_1653,N_24956,N_24812);
xnor UO_1654 (O_1654,N_24925,N_24930);
xor UO_1655 (O_1655,N_24849,N_24924);
xnor UO_1656 (O_1656,N_24860,N_24928);
xnor UO_1657 (O_1657,N_24956,N_24960);
and UO_1658 (O_1658,N_24892,N_24907);
or UO_1659 (O_1659,N_24895,N_24985);
xnor UO_1660 (O_1660,N_24853,N_24961);
and UO_1661 (O_1661,N_24901,N_24963);
and UO_1662 (O_1662,N_24800,N_24980);
nor UO_1663 (O_1663,N_24923,N_24908);
and UO_1664 (O_1664,N_24905,N_24971);
xor UO_1665 (O_1665,N_24960,N_24905);
nand UO_1666 (O_1666,N_24836,N_24821);
or UO_1667 (O_1667,N_24943,N_24910);
or UO_1668 (O_1668,N_24819,N_24964);
nand UO_1669 (O_1669,N_24947,N_24845);
nor UO_1670 (O_1670,N_24899,N_24828);
and UO_1671 (O_1671,N_24817,N_24868);
nand UO_1672 (O_1672,N_24894,N_24989);
or UO_1673 (O_1673,N_24883,N_24962);
nor UO_1674 (O_1674,N_24968,N_24842);
nor UO_1675 (O_1675,N_24801,N_24991);
xnor UO_1676 (O_1676,N_24945,N_24960);
nand UO_1677 (O_1677,N_24949,N_24971);
xnor UO_1678 (O_1678,N_24996,N_24842);
or UO_1679 (O_1679,N_24858,N_24882);
nor UO_1680 (O_1680,N_24996,N_24941);
nor UO_1681 (O_1681,N_24992,N_24984);
or UO_1682 (O_1682,N_24889,N_24807);
or UO_1683 (O_1683,N_24878,N_24902);
xor UO_1684 (O_1684,N_24869,N_24937);
nand UO_1685 (O_1685,N_24893,N_24860);
nor UO_1686 (O_1686,N_24961,N_24969);
and UO_1687 (O_1687,N_24965,N_24845);
nor UO_1688 (O_1688,N_24893,N_24823);
nor UO_1689 (O_1689,N_24958,N_24954);
nor UO_1690 (O_1690,N_24949,N_24959);
and UO_1691 (O_1691,N_24933,N_24926);
or UO_1692 (O_1692,N_24846,N_24870);
and UO_1693 (O_1693,N_24998,N_24966);
nand UO_1694 (O_1694,N_24930,N_24919);
xor UO_1695 (O_1695,N_24869,N_24864);
or UO_1696 (O_1696,N_24907,N_24831);
or UO_1697 (O_1697,N_24823,N_24828);
nor UO_1698 (O_1698,N_24869,N_24915);
nor UO_1699 (O_1699,N_24905,N_24846);
nor UO_1700 (O_1700,N_24865,N_24978);
or UO_1701 (O_1701,N_24853,N_24998);
xor UO_1702 (O_1702,N_24807,N_24837);
or UO_1703 (O_1703,N_24839,N_24962);
nor UO_1704 (O_1704,N_24852,N_24977);
or UO_1705 (O_1705,N_24803,N_24936);
nor UO_1706 (O_1706,N_24810,N_24833);
and UO_1707 (O_1707,N_24992,N_24931);
xnor UO_1708 (O_1708,N_24817,N_24821);
nor UO_1709 (O_1709,N_24990,N_24999);
or UO_1710 (O_1710,N_24993,N_24907);
xnor UO_1711 (O_1711,N_24902,N_24971);
nand UO_1712 (O_1712,N_24859,N_24941);
xnor UO_1713 (O_1713,N_24819,N_24827);
or UO_1714 (O_1714,N_24818,N_24956);
nand UO_1715 (O_1715,N_24884,N_24895);
nor UO_1716 (O_1716,N_24812,N_24998);
xnor UO_1717 (O_1717,N_24908,N_24936);
nand UO_1718 (O_1718,N_24994,N_24818);
or UO_1719 (O_1719,N_24989,N_24802);
and UO_1720 (O_1720,N_24972,N_24856);
xnor UO_1721 (O_1721,N_24960,N_24958);
nand UO_1722 (O_1722,N_24811,N_24852);
nor UO_1723 (O_1723,N_24834,N_24919);
or UO_1724 (O_1724,N_24961,N_24888);
xnor UO_1725 (O_1725,N_24802,N_24993);
or UO_1726 (O_1726,N_24870,N_24849);
xnor UO_1727 (O_1727,N_24800,N_24901);
xor UO_1728 (O_1728,N_24975,N_24810);
nand UO_1729 (O_1729,N_24915,N_24908);
or UO_1730 (O_1730,N_24982,N_24853);
or UO_1731 (O_1731,N_24903,N_24947);
or UO_1732 (O_1732,N_24847,N_24896);
nor UO_1733 (O_1733,N_24971,N_24977);
nor UO_1734 (O_1734,N_24984,N_24810);
nand UO_1735 (O_1735,N_24971,N_24853);
and UO_1736 (O_1736,N_24808,N_24833);
nor UO_1737 (O_1737,N_24899,N_24997);
xor UO_1738 (O_1738,N_24908,N_24968);
nand UO_1739 (O_1739,N_24870,N_24938);
nand UO_1740 (O_1740,N_24995,N_24932);
nor UO_1741 (O_1741,N_24809,N_24860);
xnor UO_1742 (O_1742,N_24804,N_24910);
xor UO_1743 (O_1743,N_24817,N_24818);
nor UO_1744 (O_1744,N_24877,N_24824);
nand UO_1745 (O_1745,N_24908,N_24802);
nor UO_1746 (O_1746,N_24841,N_24804);
or UO_1747 (O_1747,N_24846,N_24806);
and UO_1748 (O_1748,N_24913,N_24876);
nand UO_1749 (O_1749,N_24845,N_24963);
nor UO_1750 (O_1750,N_24904,N_24988);
and UO_1751 (O_1751,N_24882,N_24817);
nor UO_1752 (O_1752,N_24828,N_24969);
and UO_1753 (O_1753,N_24898,N_24851);
nand UO_1754 (O_1754,N_24945,N_24966);
xor UO_1755 (O_1755,N_24986,N_24978);
or UO_1756 (O_1756,N_24814,N_24945);
or UO_1757 (O_1757,N_24888,N_24927);
or UO_1758 (O_1758,N_24987,N_24852);
and UO_1759 (O_1759,N_24913,N_24805);
nand UO_1760 (O_1760,N_24989,N_24809);
xor UO_1761 (O_1761,N_24863,N_24986);
and UO_1762 (O_1762,N_24838,N_24924);
nand UO_1763 (O_1763,N_24853,N_24954);
or UO_1764 (O_1764,N_24900,N_24897);
xor UO_1765 (O_1765,N_24800,N_24907);
and UO_1766 (O_1766,N_24839,N_24930);
or UO_1767 (O_1767,N_24828,N_24803);
nor UO_1768 (O_1768,N_24859,N_24881);
and UO_1769 (O_1769,N_24812,N_24901);
nor UO_1770 (O_1770,N_24858,N_24978);
and UO_1771 (O_1771,N_24878,N_24808);
or UO_1772 (O_1772,N_24814,N_24953);
nor UO_1773 (O_1773,N_24804,N_24887);
nor UO_1774 (O_1774,N_24960,N_24847);
xnor UO_1775 (O_1775,N_24893,N_24993);
or UO_1776 (O_1776,N_24987,N_24930);
and UO_1777 (O_1777,N_24989,N_24860);
xnor UO_1778 (O_1778,N_24957,N_24821);
nor UO_1779 (O_1779,N_24808,N_24952);
nand UO_1780 (O_1780,N_24896,N_24956);
nor UO_1781 (O_1781,N_24949,N_24884);
nand UO_1782 (O_1782,N_24815,N_24810);
or UO_1783 (O_1783,N_24984,N_24950);
nor UO_1784 (O_1784,N_24972,N_24954);
or UO_1785 (O_1785,N_24860,N_24826);
and UO_1786 (O_1786,N_24910,N_24969);
xnor UO_1787 (O_1787,N_24970,N_24832);
nand UO_1788 (O_1788,N_24887,N_24818);
nand UO_1789 (O_1789,N_24999,N_24941);
and UO_1790 (O_1790,N_24941,N_24954);
and UO_1791 (O_1791,N_24872,N_24878);
nand UO_1792 (O_1792,N_24834,N_24829);
nor UO_1793 (O_1793,N_24887,N_24826);
xor UO_1794 (O_1794,N_24814,N_24864);
nand UO_1795 (O_1795,N_24915,N_24902);
or UO_1796 (O_1796,N_24955,N_24954);
or UO_1797 (O_1797,N_24966,N_24976);
nor UO_1798 (O_1798,N_24822,N_24909);
nand UO_1799 (O_1799,N_24986,N_24870);
or UO_1800 (O_1800,N_24972,N_24862);
xor UO_1801 (O_1801,N_24960,N_24885);
xnor UO_1802 (O_1802,N_24940,N_24888);
nand UO_1803 (O_1803,N_24905,N_24852);
nand UO_1804 (O_1804,N_24967,N_24884);
nand UO_1805 (O_1805,N_24924,N_24883);
or UO_1806 (O_1806,N_24844,N_24905);
or UO_1807 (O_1807,N_24895,N_24916);
nand UO_1808 (O_1808,N_24824,N_24918);
and UO_1809 (O_1809,N_24822,N_24829);
nand UO_1810 (O_1810,N_24967,N_24936);
or UO_1811 (O_1811,N_24969,N_24946);
and UO_1812 (O_1812,N_24963,N_24898);
xnor UO_1813 (O_1813,N_24885,N_24943);
nor UO_1814 (O_1814,N_24888,N_24877);
nand UO_1815 (O_1815,N_24819,N_24911);
or UO_1816 (O_1816,N_24854,N_24940);
nor UO_1817 (O_1817,N_24830,N_24957);
nor UO_1818 (O_1818,N_24849,N_24960);
or UO_1819 (O_1819,N_24861,N_24992);
nor UO_1820 (O_1820,N_24967,N_24976);
nor UO_1821 (O_1821,N_24973,N_24840);
xnor UO_1822 (O_1822,N_24903,N_24868);
xor UO_1823 (O_1823,N_24879,N_24807);
nand UO_1824 (O_1824,N_24837,N_24811);
xor UO_1825 (O_1825,N_24851,N_24925);
xor UO_1826 (O_1826,N_24818,N_24842);
or UO_1827 (O_1827,N_24813,N_24911);
nor UO_1828 (O_1828,N_24807,N_24976);
nor UO_1829 (O_1829,N_24802,N_24999);
nand UO_1830 (O_1830,N_24991,N_24892);
xnor UO_1831 (O_1831,N_24942,N_24878);
xnor UO_1832 (O_1832,N_24899,N_24946);
nor UO_1833 (O_1833,N_24883,N_24960);
or UO_1834 (O_1834,N_24959,N_24849);
and UO_1835 (O_1835,N_24870,N_24991);
and UO_1836 (O_1836,N_24838,N_24963);
nand UO_1837 (O_1837,N_24921,N_24910);
nand UO_1838 (O_1838,N_24819,N_24810);
or UO_1839 (O_1839,N_24982,N_24996);
and UO_1840 (O_1840,N_24889,N_24932);
nor UO_1841 (O_1841,N_24832,N_24815);
nand UO_1842 (O_1842,N_24862,N_24987);
nor UO_1843 (O_1843,N_24905,N_24968);
xnor UO_1844 (O_1844,N_24981,N_24886);
or UO_1845 (O_1845,N_24897,N_24834);
nor UO_1846 (O_1846,N_24976,N_24992);
and UO_1847 (O_1847,N_24859,N_24816);
xor UO_1848 (O_1848,N_24848,N_24952);
xor UO_1849 (O_1849,N_24810,N_24946);
xor UO_1850 (O_1850,N_24934,N_24946);
or UO_1851 (O_1851,N_24923,N_24926);
nor UO_1852 (O_1852,N_24910,N_24852);
nor UO_1853 (O_1853,N_24902,N_24882);
xor UO_1854 (O_1854,N_24968,N_24917);
nand UO_1855 (O_1855,N_24999,N_24910);
nor UO_1856 (O_1856,N_24892,N_24860);
nand UO_1857 (O_1857,N_24923,N_24885);
xor UO_1858 (O_1858,N_24968,N_24851);
or UO_1859 (O_1859,N_24812,N_24962);
nand UO_1860 (O_1860,N_24847,N_24920);
xor UO_1861 (O_1861,N_24908,N_24944);
and UO_1862 (O_1862,N_24949,N_24966);
nand UO_1863 (O_1863,N_24876,N_24804);
and UO_1864 (O_1864,N_24968,N_24832);
nor UO_1865 (O_1865,N_24891,N_24975);
and UO_1866 (O_1866,N_24898,N_24999);
and UO_1867 (O_1867,N_24978,N_24944);
nand UO_1868 (O_1868,N_24983,N_24830);
nand UO_1869 (O_1869,N_24962,N_24983);
nand UO_1870 (O_1870,N_24972,N_24803);
and UO_1871 (O_1871,N_24803,N_24925);
nand UO_1872 (O_1872,N_24925,N_24943);
nand UO_1873 (O_1873,N_24806,N_24824);
nand UO_1874 (O_1874,N_24991,N_24858);
nand UO_1875 (O_1875,N_24908,N_24815);
and UO_1876 (O_1876,N_24994,N_24934);
or UO_1877 (O_1877,N_24965,N_24884);
nand UO_1878 (O_1878,N_24979,N_24879);
nor UO_1879 (O_1879,N_24871,N_24974);
xnor UO_1880 (O_1880,N_24984,N_24969);
nand UO_1881 (O_1881,N_24987,N_24819);
or UO_1882 (O_1882,N_24857,N_24817);
xor UO_1883 (O_1883,N_24854,N_24979);
xor UO_1884 (O_1884,N_24893,N_24812);
or UO_1885 (O_1885,N_24953,N_24930);
nor UO_1886 (O_1886,N_24995,N_24965);
nand UO_1887 (O_1887,N_24874,N_24926);
nand UO_1888 (O_1888,N_24883,N_24844);
xnor UO_1889 (O_1889,N_24986,N_24921);
nor UO_1890 (O_1890,N_24874,N_24962);
and UO_1891 (O_1891,N_24916,N_24893);
nor UO_1892 (O_1892,N_24873,N_24835);
nand UO_1893 (O_1893,N_24953,N_24985);
nand UO_1894 (O_1894,N_24808,N_24921);
xor UO_1895 (O_1895,N_24916,N_24943);
nand UO_1896 (O_1896,N_24817,N_24948);
or UO_1897 (O_1897,N_24832,N_24901);
nand UO_1898 (O_1898,N_24996,N_24957);
nor UO_1899 (O_1899,N_24886,N_24832);
and UO_1900 (O_1900,N_24819,N_24872);
nand UO_1901 (O_1901,N_24956,N_24920);
and UO_1902 (O_1902,N_24828,N_24961);
and UO_1903 (O_1903,N_24962,N_24882);
nor UO_1904 (O_1904,N_24880,N_24989);
xnor UO_1905 (O_1905,N_24917,N_24859);
xnor UO_1906 (O_1906,N_24972,N_24979);
nand UO_1907 (O_1907,N_24924,N_24909);
xor UO_1908 (O_1908,N_24827,N_24972);
and UO_1909 (O_1909,N_24840,N_24815);
nor UO_1910 (O_1910,N_24854,N_24877);
and UO_1911 (O_1911,N_24975,N_24811);
xnor UO_1912 (O_1912,N_24800,N_24870);
and UO_1913 (O_1913,N_24962,N_24806);
xor UO_1914 (O_1914,N_24834,N_24860);
or UO_1915 (O_1915,N_24858,N_24933);
nor UO_1916 (O_1916,N_24944,N_24817);
or UO_1917 (O_1917,N_24830,N_24991);
nand UO_1918 (O_1918,N_24926,N_24811);
nand UO_1919 (O_1919,N_24849,N_24943);
xnor UO_1920 (O_1920,N_24959,N_24974);
xnor UO_1921 (O_1921,N_24867,N_24909);
or UO_1922 (O_1922,N_24992,N_24860);
xor UO_1923 (O_1923,N_24925,N_24889);
nand UO_1924 (O_1924,N_24966,N_24981);
xnor UO_1925 (O_1925,N_24999,N_24997);
nor UO_1926 (O_1926,N_24846,N_24902);
xor UO_1927 (O_1927,N_24984,N_24932);
xnor UO_1928 (O_1928,N_24914,N_24818);
or UO_1929 (O_1929,N_24837,N_24823);
nand UO_1930 (O_1930,N_24917,N_24954);
or UO_1931 (O_1931,N_24956,N_24984);
or UO_1932 (O_1932,N_24876,N_24859);
nand UO_1933 (O_1933,N_24963,N_24841);
and UO_1934 (O_1934,N_24866,N_24835);
nor UO_1935 (O_1935,N_24806,N_24820);
nor UO_1936 (O_1936,N_24968,N_24829);
nand UO_1937 (O_1937,N_24975,N_24873);
xor UO_1938 (O_1938,N_24803,N_24882);
nor UO_1939 (O_1939,N_24886,N_24896);
and UO_1940 (O_1940,N_24859,N_24962);
xor UO_1941 (O_1941,N_24899,N_24877);
xnor UO_1942 (O_1942,N_24840,N_24977);
and UO_1943 (O_1943,N_24818,N_24918);
nor UO_1944 (O_1944,N_24804,N_24856);
nand UO_1945 (O_1945,N_24973,N_24835);
or UO_1946 (O_1946,N_24963,N_24868);
nor UO_1947 (O_1947,N_24979,N_24801);
nand UO_1948 (O_1948,N_24889,N_24973);
nand UO_1949 (O_1949,N_24891,N_24960);
nand UO_1950 (O_1950,N_24970,N_24843);
or UO_1951 (O_1951,N_24893,N_24887);
and UO_1952 (O_1952,N_24863,N_24854);
xor UO_1953 (O_1953,N_24814,N_24920);
nor UO_1954 (O_1954,N_24822,N_24824);
and UO_1955 (O_1955,N_24947,N_24815);
nand UO_1956 (O_1956,N_24849,N_24951);
nor UO_1957 (O_1957,N_24815,N_24881);
and UO_1958 (O_1958,N_24903,N_24939);
or UO_1959 (O_1959,N_24968,N_24921);
xor UO_1960 (O_1960,N_24882,N_24909);
nor UO_1961 (O_1961,N_24860,N_24960);
nand UO_1962 (O_1962,N_24806,N_24836);
nor UO_1963 (O_1963,N_24887,N_24991);
nor UO_1964 (O_1964,N_24938,N_24964);
nor UO_1965 (O_1965,N_24905,N_24923);
and UO_1966 (O_1966,N_24914,N_24949);
nor UO_1967 (O_1967,N_24823,N_24808);
and UO_1968 (O_1968,N_24841,N_24941);
nand UO_1969 (O_1969,N_24945,N_24947);
and UO_1970 (O_1970,N_24912,N_24946);
nand UO_1971 (O_1971,N_24939,N_24879);
and UO_1972 (O_1972,N_24965,N_24946);
nor UO_1973 (O_1973,N_24965,N_24821);
or UO_1974 (O_1974,N_24936,N_24934);
xor UO_1975 (O_1975,N_24840,N_24992);
nor UO_1976 (O_1976,N_24914,N_24826);
nor UO_1977 (O_1977,N_24937,N_24961);
or UO_1978 (O_1978,N_24863,N_24951);
xor UO_1979 (O_1979,N_24828,N_24838);
nor UO_1980 (O_1980,N_24896,N_24876);
or UO_1981 (O_1981,N_24858,N_24814);
nand UO_1982 (O_1982,N_24947,N_24851);
nor UO_1983 (O_1983,N_24812,N_24841);
and UO_1984 (O_1984,N_24947,N_24814);
and UO_1985 (O_1985,N_24996,N_24943);
and UO_1986 (O_1986,N_24931,N_24852);
nor UO_1987 (O_1987,N_24932,N_24864);
nor UO_1988 (O_1988,N_24900,N_24812);
nor UO_1989 (O_1989,N_24904,N_24978);
xor UO_1990 (O_1990,N_24913,N_24846);
xor UO_1991 (O_1991,N_24828,N_24861);
and UO_1992 (O_1992,N_24842,N_24923);
and UO_1993 (O_1993,N_24898,N_24943);
xnor UO_1994 (O_1994,N_24867,N_24918);
xnor UO_1995 (O_1995,N_24825,N_24864);
xor UO_1996 (O_1996,N_24885,N_24845);
xor UO_1997 (O_1997,N_24989,N_24985);
nand UO_1998 (O_1998,N_24890,N_24861);
nor UO_1999 (O_1999,N_24942,N_24815);
and UO_2000 (O_2000,N_24952,N_24809);
or UO_2001 (O_2001,N_24903,N_24933);
xor UO_2002 (O_2002,N_24943,N_24815);
xor UO_2003 (O_2003,N_24897,N_24999);
or UO_2004 (O_2004,N_24920,N_24921);
nor UO_2005 (O_2005,N_24817,N_24848);
or UO_2006 (O_2006,N_24903,N_24910);
or UO_2007 (O_2007,N_24804,N_24923);
xor UO_2008 (O_2008,N_24915,N_24960);
or UO_2009 (O_2009,N_24823,N_24857);
and UO_2010 (O_2010,N_24989,N_24993);
nor UO_2011 (O_2011,N_24851,N_24820);
and UO_2012 (O_2012,N_24856,N_24824);
or UO_2013 (O_2013,N_24927,N_24925);
or UO_2014 (O_2014,N_24975,N_24940);
or UO_2015 (O_2015,N_24834,N_24891);
nand UO_2016 (O_2016,N_24907,N_24940);
xor UO_2017 (O_2017,N_24940,N_24884);
and UO_2018 (O_2018,N_24850,N_24826);
xor UO_2019 (O_2019,N_24882,N_24980);
xor UO_2020 (O_2020,N_24847,N_24895);
and UO_2021 (O_2021,N_24989,N_24888);
or UO_2022 (O_2022,N_24810,N_24951);
and UO_2023 (O_2023,N_24955,N_24925);
nor UO_2024 (O_2024,N_24898,N_24853);
nand UO_2025 (O_2025,N_24883,N_24836);
xnor UO_2026 (O_2026,N_24873,N_24844);
or UO_2027 (O_2027,N_24961,N_24954);
nand UO_2028 (O_2028,N_24984,N_24847);
xor UO_2029 (O_2029,N_24941,N_24944);
or UO_2030 (O_2030,N_24992,N_24850);
nand UO_2031 (O_2031,N_24941,N_24835);
and UO_2032 (O_2032,N_24819,N_24808);
and UO_2033 (O_2033,N_24935,N_24870);
nand UO_2034 (O_2034,N_24850,N_24872);
nor UO_2035 (O_2035,N_24985,N_24964);
or UO_2036 (O_2036,N_24826,N_24962);
nand UO_2037 (O_2037,N_24925,N_24863);
or UO_2038 (O_2038,N_24930,N_24914);
or UO_2039 (O_2039,N_24990,N_24966);
nor UO_2040 (O_2040,N_24975,N_24994);
nor UO_2041 (O_2041,N_24942,N_24905);
or UO_2042 (O_2042,N_24920,N_24948);
nand UO_2043 (O_2043,N_24837,N_24877);
or UO_2044 (O_2044,N_24886,N_24892);
xor UO_2045 (O_2045,N_24861,N_24905);
and UO_2046 (O_2046,N_24825,N_24814);
and UO_2047 (O_2047,N_24929,N_24871);
nand UO_2048 (O_2048,N_24857,N_24941);
or UO_2049 (O_2049,N_24967,N_24922);
or UO_2050 (O_2050,N_24832,N_24802);
nor UO_2051 (O_2051,N_24957,N_24970);
nor UO_2052 (O_2052,N_24853,N_24872);
xnor UO_2053 (O_2053,N_24860,N_24945);
nand UO_2054 (O_2054,N_24915,N_24893);
and UO_2055 (O_2055,N_24968,N_24952);
and UO_2056 (O_2056,N_24970,N_24973);
nand UO_2057 (O_2057,N_24985,N_24832);
nand UO_2058 (O_2058,N_24917,N_24904);
nor UO_2059 (O_2059,N_24802,N_24863);
nand UO_2060 (O_2060,N_24842,N_24922);
xor UO_2061 (O_2061,N_24980,N_24901);
or UO_2062 (O_2062,N_24871,N_24983);
or UO_2063 (O_2063,N_24840,N_24860);
xor UO_2064 (O_2064,N_24843,N_24828);
nand UO_2065 (O_2065,N_24890,N_24998);
nor UO_2066 (O_2066,N_24908,N_24822);
nand UO_2067 (O_2067,N_24979,N_24830);
and UO_2068 (O_2068,N_24886,N_24980);
or UO_2069 (O_2069,N_24945,N_24820);
nand UO_2070 (O_2070,N_24810,N_24887);
and UO_2071 (O_2071,N_24915,N_24953);
xnor UO_2072 (O_2072,N_24994,N_24846);
xnor UO_2073 (O_2073,N_24882,N_24936);
or UO_2074 (O_2074,N_24996,N_24918);
xor UO_2075 (O_2075,N_24864,N_24900);
nand UO_2076 (O_2076,N_24935,N_24872);
nand UO_2077 (O_2077,N_24836,N_24896);
or UO_2078 (O_2078,N_24874,N_24803);
nand UO_2079 (O_2079,N_24964,N_24930);
nand UO_2080 (O_2080,N_24817,N_24953);
xnor UO_2081 (O_2081,N_24921,N_24936);
nor UO_2082 (O_2082,N_24804,N_24827);
and UO_2083 (O_2083,N_24832,N_24889);
xnor UO_2084 (O_2084,N_24951,N_24907);
and UO_2085 (O_2085,N_24954,N_24892);
nand UO_2086 (O_2086,N_24914,N_24932);
and UO_2087 (O_2087,N_24858,N_24949);
xor UO_2088 (O_2088,N_24888,N_24826);
or UO_2089 (O_2089,N_24896,N_24988);
or UO_2090 (O_2090,N_24842,N_24954);
or UO_2091 (O_2091,N_24946,N_24804);
or UO_2092 (O_2092,N_24975,N_24943);
xor UO_2093 (O_2093,N_24937,N_24868);
xor UO_2094 (O_2094,N_24824,N_24874);
and UO_2095 (O_2095,N_24850,N_24892);
nor UO_2096 (O_2096,N_24864,N_24949);
or UO_2097 (O_2097,N_24867,N_24850);
nand UO_2098 (O_2098,N_24895,N_24862);
nand UO_2099 (O_2099,N_24982,N_24946);
xor UO_2100 (O_2100,N_24858,N_24906);
or UO_2101 (O_2101,N_24924,N_24834);
nor UO_2102 (O_2102,N_24960,N_24947);
nor UO_2103 (O_2103,N_24943,N_24921);
xnor UO_2104 (O_2104,N_24948,N_24888);
nand UO_2105 (O_2105,N_24918,N_24929);
nand UO_2106 (O_2106,N_24946,N_24851);
nor UO_2107 (O_2107,N_24883,N_24820);
nor UO_2108 (O_2108,N_24971,N_24849);
xnor UO_2109 (O_2109,N_24812,N_24925);
nand UO_2110 (O_2110,N_24953,N_24902);
nand UO_2111 (O_2111,N_24861,N_24820);
and UO_2112 (O_2112,N_24946,N_24886);
or UO_2113 (O_2113,N_24851,N_24939);
and UO_2114 (O_2114,N_24973,N_24824);
and UO_2115 (O_2115,N_24961,N_24955);
xnor UO_2116 (O_2116,N_24902,N_24831);
nor UO_2117 (O_2117,N_24922,N_24876);
or UO_2118 (O_2118,N_24939,N_24861);
xnor UO_2119 (O_2119,N_24802,N_24806);
or UO_2120 (O_2120,N_24876,N_24883);
nand UO_2121 (O_2121,N_24810,N_24964);
and UO_2122 (O_2122,N_24893,N_24910);
nor UO_2123 (O_2123,N_24934,N_24967);
or UO_2124 (O_2124,N_24970,N_24982);
nor UO_2125 (O_2125,N_24835,N_24999);
nand UO_2126 (O_2126,N_24968,N_24834);
and UO_2127 (O_2127,N_24924,N_24899);
nand UO_2128 (O_2128,N_24919,N_24951);
or UO_2129 (O_2129,N_24923,N_24906);
nor UO_2130 (O_2130,N_24999,N_24899);
or UO_2131 (O_2131,N_24909,N_24988);
and UO_2132 (O_2132,N_24906,N_24879);
xor UO_2133 (O_2133,N_24898,N_24822);
xor UO_2134 (O_2134,N_24870,N_24965);
nand UO_2135 (O_2135,N_24936,N_24990);
or UO_2136 (O_2136,N_24817,N_24951);
nand UO_2137 (O_2137,N_24818,N_24991);
xnor UO_2138 (O_2138,N_24898,N_24931);
xor UO_2139 (O_2139,N_24993,N_24939);
xnor UO_2140 (O_2140,N_24959,N_24976);
or UO_2141 (O_2141,N_24843,N_24868);
nor UO_2142 (O_2142,N_24964,N_24815);
nand UO_2143 (O_2143,N_24931,N_24995);
nand UO_2144 (O_2144,N_24985,N_24881);
xnor UO_2145 (O_2145,N_24868,N_24925);
nor UO_2146 (O_2146,N_24845,N_24857);
or UO_2147 (O_2147,N_24889,N_24842);
and UO_2148 (O_2148,N_24969,N_24800);
and UO_2149 (O_2149,N_24877,N_24847);
and UO_2150 (O_2150,N_24841,N_24815);
nand UO_2151 (O_2151,N_24943,N_24993);
nor UO_2152 (O_2152,N_24893,N_24857);
or UO_2153 (O_2153,N_24875,N_24860);
xor UO_2154 (O_2154,N_24847,N_24933);
xnor UO_2155 (O_2155,N_24936,N_24816);
xnor UO_2156 (O_2156,N_24969,N_24991);
or UO_2157 (O_2157,N_24913,N_24868);
nor UO_2158 (O_2158,N_24875,N_24843);
and UO_2159 (O_2159,N_24802,N_24853);
nor UO_2160 (O_2160,N_24914,N_24872);
nand UO_2161 (O_2161,N_24803,N_24847);
xnor UO_2162 (O_2162,N_24889,N_24803);
or UO_2163 (O_2163,N_24990,N_24988);
nand UO_2164 (O_2164,N_24848,N_24837);
xnor UO_2165 (O_2165,N_24914,N_24820);
nor UO_2166 (O_2166,N_24894,N_24951);
nand UO_2167 (O_2167,N_24856,N_24834);
xnor UO_2168 (O_2168,N_24832,N_24863);
or UO_2169 (O_2169,N_24962,N_24913);
xor UO_2170 (O_2170,N_24846,N_24933);
or UO_2171 (O_2171,N_24924,N_24846);
nand UO_2172 (O_2172,N_24815,N_24930);
xnor UO_2173 (O_2173,N_24954,N_24879);
xor UO_2174 (O_2174,N_24927,N_24960);
nand UO_2175 (O_2175,N_24814,N_24831);
nand UO_2176 (O_2176,N_24940,N_24810);
nor UO_2177 (O_2177,N_24903,N_24960);
nor UO_2178 (O_2178,N_24808,N_24985);
nand UO_2179 (O_2179,N_24826,N_24988);
and UO_2180 (O_2180,N_24842,N_24850);
nor UO_2181 (O_2181,N_24873,N_24870);
nand UO_2182 (O_2182,N_24883,N_24850);
and UO_2183 (O_2183,N_24850,N_24969);
nand UO_2184 (O_2184,N_24947,N_24963);
xor UO_2185 (O_2185,N_24885,N_24959);
nor UO_2186 (O_2186,N_24958,N_24948);
and UO_2187 (O_2187,N_24816,N_24914);
nand UO_2188 (O_2188,N_24951,N_24950);
xnor UO_2189 (O_2189,N_24973,N_24916);
xor UO_2190 (O_2190,N_24931,N_24879);
nor UO_2191 (O_2191,N_24824,N_24969);
and UO_2192 (O_2192,N_24896,N_24832);
nand UO_2193 (O_2193,N_24982,N_24907);
and UO_2194 (O_2194,N_24972,N_24818);
xor UO_2195 (O_2195,N_24805,N_24902);
nand UO_2196 (O_2196,N_24978,N_24848);
or UO_2197 (O_2197,N_24916,N_24991);
nand UO_2198 (O_2198,N_24899,N_24908);
xor UO_2199 (O_2199,N_24896,N_24806);
or UO_2200 (O_2200,N_24885,N_24925);
nor UO_2201 (O_2201,N_24824,N_24931);
nand UO_2202 (O_2202,N_24907,N_24962);
nor UO_2203 (O_2203,N_24827,N_24884);
nor UO_2204 (O_2204,N_24894,N_24974);
nor UO_2205 (O_2205,N_24893,N_24901);
and UO_2206 (O_2206,N_24826,N_24945);
or UO_2207 (O_2207,N_24879,N_24926);
and UO_2208 (O_2208,N_24942,N_24805);
nand UO_2209 (O_2209,N_24842,N_24846);
nor UO_2210 (O_2210,N_24885,N_24818);
nor UO_2211 (O_2211,N_24903,N_24804);
xor UO_2212 (O_2212,N_24962,N_24999);
xor UO_2213 (O_2213,N_24986,N_24876);
nand UO_2214 (O_2214,N_24825,N_24875);
or UO_2215 (O_2215,N_24925,N_24811);
nor UO_2216 (O_2216,N_24822,N_24989);
xor UO_2217 (O_2217,N_24899,N_24827);
nor UO_2218 (O_2218,N_24888,N_24891);
xor UO_2219 (O_2219,N_24954,N_24971);
xnor UO_2220 (O_2220,N_24934,N_24820);
nand UO_2221 (O_2221,N_24865,N_24848);
nand UO_2222 (O_2222,N_24947,N_24839);
nor UO_2223 (O_2223,N_24802,N_24875);
xor UO_2224 (O_2224,N_24998,N_24938);
nand UO_2225 (O_2225,N_24974,N_24891);
nand UO_2226 (O_2226,N_24825,N_24956);
and UO_2227 (O_2227,N_24826,N_24806);
xnor UO_2228 (O_2228,N_24952,N_24843);
and UO_2229 (O_2229,N_24935,N_24828);
or UO_2230 (O_2230,N_24945,N_24875);
nor UO_2231 (O_2231,N_24932,N_24841);
nor UO_2232 (O_2232,N_24906,N_24843);
nor UO_2233 (O_2233,N_24841,N_24862);
xor UO_2234 (O_2234,N_24892,N_24808);
and UO_2235 (O_2235,N_24804,N_24866);
and UO_2236 (O_2236,N_24956,N_24985);
xnor UO_2237 (O_2237,N_24810,N_24924);
and UO_2238 (O_2238,N_24856,N_24908);
nor UO_2239 (O_2239,N_24880,N_24988);
and UO_2240 (O_2240,N_24817,N_24905);
nor UO_2241 (O_2241,N_24912,N_24945);
xnor UO_2242 (O_2242,N_24942,N_24833);
xnor UO_2243 (O_2243,N_24852,N_24962);
or UO_2244 (O_2244,N_24871,N_24901);
nand UO_2245 (O_2245,N_24887,N_24907);
nor UO_2246 (O_2246,N_24991,N_24861);
or UO_2247 (O_2247,N_24905,N_24821);
nand UO_2248 (O_2248,N_24939,N_24934);
and UO_2249 (O_2249,N_24986,N_24979);
or UO_2250 (O_2250,N_24883,N_24997);
xnor UO_2251 (O_2251,N_24835,N_24914);
nand UO_2252 (O_2252,N_24950,N_24909);
xnor UO_2253 (O_2253,N_24851,N_24931);
nor UO_2254 (O_2254,N_24943,N_24835);
and UO_2255 (O_2255,N_24868,N_24833);
or UO_2256 (O_2256,N_24858,N_24804);
nand UO_2257 (O_2257,N_24844,N_24884);
nor UO_2258 (O_2258,N_24872,N_24887);
xnor UO_2259 (O_2259,N_24905,N_24931);
or UO_2260 (O_2260,N_24843,N_24882);
xnor UO_2261 (O_2261,N_24800,N_24956);
and UO_2262 (O_2262,N_24892,N_24837);
xor UO_2263 (O_2263,N_24886,N_24867);
or UO_2264 (O_2264,N_24992,N_24835);
nand UO_2265 (O_2265,N_24942,N_24982);
nand UO_2266 (O_2266,N_24898,N_24955);
xor UO_2267 (O_2267,N_24887,N_24871);
xnor UO_2268 (O_2268,N_24921,N_24866);
xor UO_2269 (O_2269,N_24808,N_24910);
nor UO_2270 (O_2270,N_24862,N_24951);
and UO_2271 (O_2271,N_24854,N_24808);
and UO_2272 (O_2272,N_24872,N_24825);
and UO_2273 (O_2273,N_24839,N_24931);
or UO_2274 (O_2274,N_24963,N_24856);
nor UO_2275 (O_2275,N_24969,N_24868);
or UO_2276 (O_2276,N_24964,N_24911);
and UO_2277 (O_2277,N_24971,N_24986);
or UO_2278 (O_2278,N_24812,N_24892);
or UO_2279 (O_2279,N_24994,N_24853);
nor UO_2280 (O_2280,N_24881,N_24893);
and UO_2281 (O_2281,N_24965,N_24863);
or UO_2282 (O_2282,N_24902,N_24927);
and UO_2283 (O_2283,N_24955,N_24936);
nand UO_2284 (O_2284,N_24936,N_24952);
xnor UO_2285 (O_2285,N_24822,N_24883);
xnor UO_2286 (O_2286,N_24863,N_24942);
nor UO_2287 (O_2287,N_24953,N_24856);
nand UO_2288 (O_2288,N_24904,N_24814);
xnor UO_2289 (O_2289,N_24831,N_24804);
and UO_2290 (O_2290,N_24818,N_24901);
or UO_2291 (O_2291,N_24849,N_24923);
xor UO_2292 (O_2292,N_24993,N_24930);
and UO_2293 (O_2293,N_24946,N_24867);
nand UO_2294 (O_2294,N_24925,N_24933);
xnor UO_2295 (O_2295,N_24960,N_24913);
xnor UO_2296 (O_2296,N_24832,N_24958);
or UO_2297 (O_2297,N_24914,N_24931);
nor UO_2298 (O_2298,N_24807,N_24878);
nand UO_2299 (O_2299,N_24823,N_24925);
and UO_2300 (O_2300,N_24930,N_24924);
xor UO_2301 (O_2301,N_24823,N_24991);
or UO_2302 (O_2302,N_24977,N_24966);
or UO_2303 (O_2303,N_24843,N_24909);
xor UO_2304 (O_2304,N_24813,N_24809);
xnor UO_2305 (O_2305,N_24857,N_24828);
nor UO_2306 (O_2306,N_24874,N_24941);
xor UO_2307 (O_2307,N_24826,N_24971);
nand UO_2308 (O_2308,N_24932,N_24938);
xnor UO_2309 (O_2309,N_24837,N_24874);
and UO_2310 (O_2310,N_24951,N_24847);
or UO_2311 (O_2311,N_24928,N_24834);
nor UO_2312 (O_2312,N_24976,N_24956);
or UO_2313 (O_2313,N_24962,N_24922);
xnor UO_2314 (O_2314,N_24900,N_24937);
nor UO_2315 (O_2315,N_24981,N_24942);
and UO_2316 (O_2316,N_24973,N_24969);
or UO_2317 (O_2317,N_24978,N_24876);
and UO_2318 (O_2318,N_24835,N_24876);
nor UO_2319 (O_2319,N_24933,N_24901);
nand UO_2320 (O_2320,N_24960,N_24999);
xnor UO_2321 (O_2321,N_24887,N_24841);
xnor UO_2322 (O_2322,N_24991,N_24922);
and UO_2323 (O_2323,N_24807,N_24893);
or UO_2324 (O_2324,N_24979,N_24829);
and UO_2325 (O_2325,N_24905,N_24918);
nand UO_2326 (O_2326,N_24905,N_24810);
or UO_2327 (O_2327,N_24859,N_24815);
nand UO_2328 (O_2328,N_24907,N_24955);
nand UO_2329 (O_2329,N_24842,N_24906);
nor UO_2330 (O_2330,N_24802,N_24971);
nand UO_2331 (O_2331,N_24830,N_24844);
nor UO_2332 (O_2332,N_24919,N_24966);
nor UO_2333 (O_2333,N_24941,N_24930);
nor UO_2334 (O_2334,N_24939,N_24821);
nor UO_2335 (O_2335,N_24992,N_24955);
or UO_2336 (O_2336,N_24864,N_24938);
or UO_2337 (O_2337,N_24887,N_24881);
nand UO_2338 (O_2338,N_24817,N_24959);
xor UO_2339 (O_2339,N_24944,N_24807);
or UO_2340 (O_2340,N_24843,N_24841);
nand UO_2341 (O_2341,N_24817,N_24802);
nand UO_2342 (O_2342,N_24934,N_24927);
and UO_2343 (O_2343,N_24842,N_24966);
xnor UO_2344 (O_2344,N_24939,N_24933);
nand UO_2345 (O_2345,N_24835,N_24972);
nor UO_2346 (O_2346,N_24939,N_24890);
and UO_2347 (O_2347,N_24834,N_24852);
nor UO_2348 (O_2348,N_24859,N_24838);
nand UO_2349 (O_2349,N_24809,N_24923);
or UO_2350 (O_2350,N_24810,N_24803);
or UO_2351 (O_2351,N_24976,N_24874);
or UO_2352 (O_2352,N_24901,N_24989);
or UO_2353 (O_2353,N_24839,N_24844);
nor UO_2354 (O_2354,N_24836,N_24902);
or UO_2355 (O_2355,N_24891,N_24958);
nand UO_2356 (O_2356,N_24953,N_24871);
nand UO_2357 (O_2357,N_24931,N_24994);
nor UO_2358 (O_2358,N_24833,N_24979);
nor UO_2359 (O_2359,N_24808,N_24903);
xnor UO_2360 (O_2360,N_24819,N_24841);
and UO_2361 (O_2361,N_24880,N_24845);
nor UO_2362 (O_2362,N_24850,N_24879);
or UO_2363 (O_2363,N_24803,N_24940);
xnor UO_2364 (O_2364,N_24936,N_24912);
or UO_2365 (O_2365,N_24994,N_24854);
xor UO_2366 (O_2366,N_24885,N_24987);
and UO_2367 (O_2367,N_24924,N_24886);
nand UO_2368 (O_2368,N_24891,N_24831);
and UO_2369 (O_2369,N_24852,N_24942);
or UO_2370 (O_2370,N_24901,N_24880);
and UO_2371 (O_2371,N_24985,N_24856);
and UO_2372 (O_2372,N_24814,N_24978);
nor UO_2373 (O_2373,N_24861,N_24922);
and UO_2374 (O_2374,N_24956,N_24829);
and UO_2375 (O_2375,N_24835,N_24827);
or UO_2376 (O_2376,N_24845,N_24950);
or UO_2377 (O_2377,N_24937,N_24901);
nor UO_2378 (O_2378,N_24881,N_24987);
xnor UO_2379 (O_2379,N_24855,N_24857);
or UO_2380 (O_2380,N_24904,N_24804);
xnor UO_2381 (O_2381,N_24946,N_24812);
or UO_2382 (O_2382,N_24998,N_24895);
nand UO_2383 (O_2383,N_24872,N_24967);
xnor UO_2384 (O_2384,N_24952,N_24813);
nand UO_2385 (O_2385,N_24836,N_24916);
nor UO_2386 (O_2386,N_24857,N_24832);
xor UO_2387 (O_2387,N_24900,N_24841);
nor UO_2388 (O_2388,N_24970,N_24893);
nor UO_2389 (O_2389,N_24995,N_24925);
or UO_2390 (O_2390,N_24855,N_24928);
and UO_2391 (O_2391,N_24835,N_24921);
nor UO_2392 (O_2392,N_24908,N_24965);
nor UO_2393 (O_2393,N_24931,N_24807);
xor UO_2394 (O_2394,N_24904,N_24882);
nor UO_2395 (O_2395,N_24947,N_24803);
nand UO_2396 (O_2396,N_24878,N_24927);
and UO_2397 (O_2397,N_24829,N_24863);
nand UO_2398 (O_2398,N_24874,N_24923);
xor UO_2399 (O_2399,N_24959,N_24989);
nand UO_2400 (O_2400,N_24830,N_24923);
nor UO_2401 (O_2401,N_24996,N_24822);
nand UO_2402 (O_2402,N_24962,N_24829);
and UO_2403 (O_2403,N_24815,N_24921);
or UO_2404 (O_2404,N_24910,N_24951);
nor UO_2405 (O_2405,N_24902,N_24918);
xor UO_2406 (O_2406,N_24934,N_24813);
xor UO_2407 (O_2407,N_24830,N_24929);
xor UO_2408 (O_2408,N_24882,N_24850);
nand UO_2409 (O_2409,N_24906,N_24902);
nor UO_2410 (O_2410,N_24810,N_24944);
nor UO_2411 (O_2411,N_24953,N_24819);
xnor UO_2412 (O_2412,N_24805,N_24929);
and UO_2413 (O_2413,N_24921,N_24933);
or UO_2414 (O_2414,N_24946,N_24979);
nor UO_2415 (O_2415,N_24980,N_24881);
nor UO_2416 (O_2416,N_24955,N_24938);
and UO_2417 (O_2417,N_24888,N_24964);
or UO_2418 (O_2418,N_24964,N_24995);
or UO_2419 (O_2419,N_24974,N_24836);
xor UO_2420 (O_2420,N_24896,N_24807);
and UO_2421 (O_2421,N_24952,N_24882);
nor UO_2422 (O_2422,N_24808,N_24905);
xnor UO_2423 (O_2423,N_24823,N_24993);
xnor UO_2424 (O_2424,N_24812,N_24809);
xor UO_2425 (O_2425,N_24932,N_24855);
nand UO_2426 (O_2426,N_24825,N_24876);
or UO_2427 (O_2427,N_24853,N_24858);
and UO_2428 (O_2428,N_24908,N_24938);
xor UO_2429 (O_2429,N_24850,N_24957);
xnor UO_2430 (O_2430,N_24973,N_24827);
nor UO_2431 (O_2431,N_24842,N_24951);
and UO_2432 (O_2432,N_24962,N_24872);
xor UO_2433 (O_2433,N_24804,N_24943);
xor UO_2434 (O_2434,N_24882,N_24800);
nand UO_2435 (O_2435,N_24932,N_24940);
xor UO_2436 (O_2436,N_24949,N_24933);
and UO_2437 (O_2437,N_24828,N_24983);
nor UO_2438 (O_2438,N_24834,N_24944);
nand UO_2439 (O_2439,N_24820,N_24808);
or UO_2440 (O_2440,N_24902,N_24895);
and UO_2441 (O_2441,N_24942,N_24947);
nor UO_2442 (O_2442,N_24868,N_24915);
nand UO_2443 (O_2443,N_24986,N_24878);
xor UO_2444 (O_2444,N_24845,N_24933);
nand UO_2445 (O_2445,N_24898,N_24878);
xor UO_2446 (O_2446,N_24839,N_24879);
or UO_2447 (O_2447,N_24897,N_24945);
or UO_2448 (O_2448,N_24917,N_24922);
xnor UO_2449 (O_2449,N_24894,N_24820);
nor UO_2450 (O_2450,N_24909,N_24868);
nand UO_2451 (O_2451,N_24993,N_24835);
nand UO_2452 (O_2452,N_24846,N_24825);
nand UO_2453 (O_2453,N_24991,N_24911);
nor UO_2454 (O_2454,N_24856,N_24840);
or UO_2455 (O_2455,N_24974,N_24960);
xor UO_2456 (O_2456,N_24860,N_24982);
nor UO_2457 (O_2457,N_24916,N_24927);
and UO_2458 (O_2458,N_24985,N_24909);
xnor UO_2459 (O_2459,N_24890,N_24828);
xnor UO_2460 (O_2460,N_24954,N_24987);
xor UO_2461 (O_2461,N_24838,N_24961);
nor UO_2462 (O_2462,N_24853,N_24835);
nand UO_2463 (O_2463,N_24919,N_24851);
nor UO_2464 (O_2464,N_24863,N_24842);
or UO_2465 (O_2465,N_24879,N_24996);
or UO_2466 (O_2466,N_24911,N_24804);
and UO_2467 (O_2467,N_24816,N_24959);
nand UO_2468 (O_2468,N_24943,N_24843);
nor UO_2469 (O_2469,N_24889,N_24823);
nor UO_2470 (O_2470,N_24936,N_24847);
and UO_2471 (O_2471,N_24800,N_24831);
nand UO_2472 (O_2472,N_24951,N_24900);
or UO_2473 (O_2473,N_24958,N_24961);
xnor UO_2474 (O_2474,N_24879,N_24898);
xnor UO_2475 (O_2475,N_24923,N_24894);
or UO_2476 (O_2476,N_24815,N_24957);
or UO_2477 (O_2477,N_24997,N_24870);
xnor UO_2478 (O_2478,N_24974,N_24862);
nor UO_2479 (O_2479,N_24931,N_24978);
or UO_2480 (O_2480,N_24848,N_24878);
or UO_2481 (O_2481,N_24896,N_24951);
and UO_2482 (O_2482,N_24910,N_24885);
xnor UO_2483 (O_2483,N_24899,N_24989);
nand UO_2484 (O_2484,N_24838,N_24999);
or UO_2485 (O_2485,N_24915,N_24850);
xor UO_2486 (O_2486,N_24900,N_24903);
nor UO_2487 (O_2487,N_24920,N_24870);
or UO_2488 (O_2488,N_24945,N_24878);
nand UO_2489 (O_2489,N_24998,N_24975);
and UO_2490 (O_2490,N_24847,N_24831);
and UO_2491 (O_2491,N_24814,N_24801);
nor UO_2492 (O_2492,N_24967,N_24842);
nor UO_2493 (O_2493,N_24938,N_24914);
xor UO_2494 (O_2494,N_24944,N_24984);
nor UO_2495 (O_2495,N_24880,N_24966);
or UO_2496 (O_2496,N_24949,N_24977);
or UO_2497 (O_2497,N_24897,N_24927);
nand UO_2498 (O_2498,N_24961,N_24836);
and UO_2499 (O_2499,N_24979,N_24941);
nand UO_2500 (O_2500,N_24953,N_24884);
or UO_2501 (O_2501,N_24948,N_24956);
or UO_2502 (O_2502,N_24828,N_24904);
and UO_2503 (O_2503,N_24998,N_24815);
xnor UO_2504 (O_2504,N_24894,N_24869);
nor UO_2505 (O_2505,N_24975,N_24982);
and UO_2506 (O_2506,N_24839,N_24843);
and UO_2507 (O_2507,N_24857,N_24818);
or UO_2508 (O_2508,N_24977,N_24806);
nor UO_2509 (O_2509,N_24905,N_24834);
and UO_2510 (O_2510,N_24876,N_24870);
nand UO_2511 (O_2511,N_24918,N_24975);
nand UO_2512 (O_2512,N_24869,N_24941);
nand UO_2513 (O_2513,N_24807,N_24977);
or UO_2514 (O_2514,N_24932,N_24918);
nand UO_2515 (O_2515,N_24812,N_24827);
nor UO_2516 (O_2516,N_24970,N_24856);
or UO_2517 (O_2517,N_24981,N_24901);
or UO_2518 (O_2518,N_24853,N_24866);
and UO_2519 (O_2519,N_24937,N_24826);
xor UO_2520 (O_2520,N_24851,N_24806);
nor UO_2521 (O_2521,N_24935,N_24970);
xnor UO_2522 (O_2522,N_24877,N_24917);
and UO_2523 (O_2523,N_24990,N_24867);
or UO_2524 (O_2524,N_24881,N_24828);
nor UO_2525 (O_2525,N_24965,N_24893);
nand UO_2526 (O_2526,N_24889,N_24918);
nand UO_2527 (O_2527,N_24877,N_24972);
nor UO_2528 (O_2528,N_24901,N_24969);
xor UO_2529 (O_2529,N_24958,N_24888);
nand UO_2530 (O_2530,N_24855,N_24902);
or UO_2531 (O_2531,N_24975,N_24832);
or UO_2532 (O_2532,N_24908,N_24895);
xor UO_2533 (O_2533,N_24840,N_24853);
nor UO_2534 (O_2534,N_24928,N_24895);
and UO_2535 (O_2535,N_24873,N_24894);
xnor UO_2536 (O_2536,N_24895,N_24980);
and UO_2537 (O_2537,N_24833,N_24968);
and UO_2538 (O_2538,N_24846,N_24901);
or UO_2539 (O_2539,N_24863,N_24932);
nor UO_2540 (O_2540,N_24831,N_24842);
or UO_2541 (O_2541,N_24926,N_24836);
nor UO_2542 (O_2542,N_24904,N_24973);
nor UO_2543 (O_2543,N_24916,N_24881);
nand UO_2544 (O_2544,N_24931,N_24951);
nand UO_2545 (O_2545,N_24856,N_24900);
and UO_2546 (O_2546,N_24979,N_24908);
and UO_2547 (O_2547,N_24953,N_24971);
nor UO_2548 (O_2548,N_24802,N_24954);
and UO_2549 (O_2549,N_24909,N_24895);
nand UO_2550 (O_2550,N_24864,N_24887);
nor UO_2551 (O_2551,N_24835,N_24962);
xor UO_2552 (O_2552,N_24971,N_24851);
or UO_2553 (O_2553,N_24855,N_24907);
and UO_2554 (O_2554,N_24873,N_24910);
and UO_2555 (O_2555,N_24835,N_24854);
nor UO_2556 (O_2556,N_24888,N_24976);
and UO_2557 (O_2557,N_24930,N_24917);
or UO_2558 (O_2558,N_24947,N_24940);
or UO_2559 (O_2559,N_24812,N_24838);
nor UO_2560 (O_2560,N_24852,N_24914);
and UO_2561 (O_2561,N_24859,N_24903);
and UO_2562 (O_2562,N_24979,N_24847);
xnor UO_2563 (O_2563,N_24913,N_24937);
xor UO_2564 (O_2564,N_24876,N_24829);
or UO_2565 (O_2565,N_24891,N_24984);
nand UO_2566 (O_2566,N_24894,N_24862);
nand UO_2567 (O_2567,N_24942,N_24987);
or UO_2568 (O_2568,N_24910,N_24813);
or UO_2569 (O_2569,N_24854,N_24917);
nor UO_2570 (O_2570,N_24993,N_24928);
xnor UO_2571 (O_2571,N_24999,N_24883);
and UO_2572 (O_2572,N_24805,N_24951);
nor UO_2573 (O_2573,N_24929,N_24867);
and UO_2574 (O_2574,N_24850,N_24871);
nand UO_2575 (O_2575,N_24901,N_24887);
or UO_2576 (O_2576,N_24874,N_24811);
nor UO_2577 (O_2577,N_24904,N_24955);
xor UO_2578 (O_2578,N_24985,N_24819);
nand UO_2579 (O_2579,N_24917,N_24831);
xor UO_2580 (O_2580,N_24826,N_24884);
nor UO_2581 (O_2581,N_24878,N_24842);
or UO_2582 (O_2582,N_24813,N_24940);
and UO_2583 (O_2583,N_24886,N_24838);
and UO_2584 (O_2584,N_24851,N_24951);
and UO_2585 (O_2585,N_24828,N_24907);
and UO_2586 (O_2586,N_24988,N_24955);
and UO_2587 (O_2587,N_24915,N_24999);
nor UO_2588 (O_2588,N_24873,N_24822);
xor UO_2589 (O_2589,N_24868,N_24916);
or UO_2590 (O_2590,N_24884,N_24972);
xor UO_2591 (O_2591,N_24984,N_24948);
nor UO_2592 (O_2592,N_24822,N_24821);
xnor UO_2593 (O_2593,N_24872,N_24980);
and UO_2594 (O_2594,N_24934,N_24855);
nand UO_2595 (O_2595,N_24953,N_24886);
nor UO_2596 (O_2596,N_24888,N_24839);
or UO_2597 (O_2597,N_24826,N_24981);
nor UO_2598 (O_2598,N_24888,N_24928);
nand UO_2599 (O_2599,N_24882,N_24911);
nor UO_2600 (O_2600,N_24998,N_24819);
xor UO_2601 (O_2601,N_24957,N_24890);
and UO_2602 (O_2602,N_24829,N_24963);
xor UO_2603 (O_2603,N_24985,N_24977);
nand UO_2604 (O_2604,N_24836,N_24978);
or UO_2605 (O_2605,N_24822,N_24966);
and UO_2606 (O_2606,N_24995,N_24864);
nand UO_2607 (O_2607,N_24996,N_24915);
nor UO_2608 (O_2608,N_24944,N_24840);
or UO_2609 (O_2609,N_24982,N_24926);
nor UO_2610 (O_2610,N_24818,N_24895);
nand UO_2611 (O_2611,N_24839,N_24853);
and UO_2612 (O_2612,N_24801,N_24941);
or UO_2613 (O_2613,N_24846,N_24980);
nor UO_2614 (O_2614,N_24840,N_24962);
nor UO_2615 (O_2615,N_24966,N_24922);
and UO_2616 (O_2616,N_24814,N_24850);
nor UO_2617 (O_2617,N_24954,N_24907);
nor UO_2618 (O_2618,N_24864,N_24925);
nand UO_2619 (O_2619,N_24942,N_24826);
and UO_2620 (O_2620,N_24820,N_24805);
xor UO_2621 (O_2621,N_24891,N_24851);
nand UO_2622 (O_2622,N_24878,N_24820);
or UO_2623 (O_2623,N_24872,N_24884);
nor UO_2624 (O_2624,N_24856,N_24820);
xor UO_2625 (O_2625,N_24991,N_24962);
xor UO_2626 (O_2626,N_24895,N_24866);
or UO_2627 (O_2627,N_24987,N_24829);
nor UO_2628 (O_2628,N_24846,N_24975);
nor UO_2629 (O_2629,N_24908,N_24995);
xnor UO_2630 (O_2630,N_24966,N_24952);
xnor UO_2631 (O_2631,N_24928,N_24891);
nor UO_2632 (O_2632,N_24997,N_24904);
and UO_2633 (O_2633,N_24803,N_24992);
or UO_2634 (O_2634,N_24854,N_24948);
and UO_2635 (O_2635,N_24931,N_24846);
or UO_2636 (O_2636,N_24826,N_24891);
xnor UO_2637 (O_2637,N_24927,N_24959);
nor UO_2638 (O_2638,N_24860,N_24807);
and UO_2639 (O_2639,N_24879,N_24869);
or UO_2640 (O_2640,N_24868,N_24869);
nor UO_2641 (O_2641,N_24855,N_24886);
or UO_2642 (O_2642,N_24916,N_24979);
nand UO_2643 (O_2643,N_24952,N_24823);
and UO_2644 (O_2644,N_24846,N_24843);
or UO_2645 (O_2645,N_24892,N_24923);
xor UO_2646 (O_2646,N_24950,N_24974);
xnor UO_2647 (O_2647,N_24957,N_24818);
or UO_2648 (O_2648,N_24862,N_24983);
xor UO_2649 (O_2649,N_24908,N_24870);
nor UO_2650 (O_2650,N_24980,N_24889);
nor UO_2651 (O_2651,N_24919,N_24943);
nor UO_2652 (O_2652,N_24909,N_24952);
nand UO_2653 (O_2653,N_24942,N_24846);
or UO_2654 (O_2654,N_24980,N_24964);
nor UO_2655 (O_2655,N_24920,N_24949);
and UO_2656 (O_2656,N_24870,N_24859);
xnor UO_2657 (O_2657,N_24835,N_24874);
and UO_2658 (O_2658,N_24982,N_24931);
and UO_2659 (O_2659,N_24896,N_24944);
nand UO_2660 (O_2660,N_24813,N_24900);
nor UO_2661 (O_2661,N_24808,N_24863);
or UO_2662 (O_2662,N_24962,N_24873);
nor UO_2663 (O_2663,N_24920,N_24987);
nand UO_2664 (O_2664,N_24906,N_24946);
nor UO_2665 (O_2665,N_24946,N_24844);
or UO_2666 (O_2666,N_24936,N_24830);
or UO_2667 (O_2667,N_24879,N_24933);
nand UO_2668 (O_2668,N_24805,N_24992);
xor UO_2669 (O_2669,N_24993,N_24902);
nand UO_2670 (O_2670,N_24924,N_24898);
and UO_2671 (O_2671,N_24844,N_24841);
or UO_2672 (O_2672,N_24987,N_24996);
xnor UO_2673 (O_2673,N_24856,N_24848);
nor UO_2674 (O_2674,N_24924,N_24928);
nand UO_2675 (O_2675,N_24846,N_24932);
or UO_2676 (O_2676,N_24909,N_24893);
or UO_2677 (O_2677,N_24994,N_24944);
nor UO_2678 (O_2678,N_24995,N_24910);
nor UO_2679 (O_2679,N_24814,N_24918);
or UO_2680 (O_2680,N_24802,N_24881);
or UO_2681 (O_2681,N_24824,N_24996);
xor UO_2682 (O_2682,N_24848,N_24830);
xor UO_2683 (O_2683,N_24853,N_24890);
nand UO_2684 (O_2684,N_24989,N_24927);
and UO_2685 (O_2685,N_24880,N_24805);
or UO_2686 (O_2686,N_24849,N_24891);
xor UO_2687 (O_2687,N_24958,N_24893);
xor UO_2688 (O_2688,N_24944,N_24841);
nand UO_2689 (O_2689,N_24852,N_24979);
or UO_2690 (O_2690,N_24834,N_24866);
nand UO_2691 (O_2691,N_24954,N_24910);
nor UO_2692 (O_2692,N_24999,N_24810);
xor UO_2693 (O_2693,N_24974,N_24910);
or UO_2694 (O_2694,N_24885,N_24901);
nand UO_2695 (O_2695,N_24938,N_24902);
nor UO_2696 (O_2696,N_24975,N_24890);
xor UO_2697 (O_2697,N_24849,N_24866);
and UO_2698 (O_2698,N_24936,N_24848);
and UO_2699 (O_2699,N_24951,N_24975);
and UO_2700 (O_2700,N_24913,N_24930);
or UO_2701 (O_2701,N_24825,N_24821);
nor UO_2702 (O_2702,N_24954,N_24861);
nor UO_2703 (O_2703,N_24943,N_24966);
nand UO_2704 (O_2704,N_24912,N_24920);
nand UO_2705 (O_2705,N_24980,N_24861);
nand UO_2706 (O_2706,N_24919,N_24830);
and UO_2707 (O_2707,N_24999,N_24935);
or UO_2708 (O_2708,N_24895,N_24966);
and UO_2709 (O_2709,N_24933,N_24943);
nor UO_2710 (O_2710,N_24972,N_24855);
nor UO_2711 (O_2711,N_24899,N_24868);
and UO_2712 (O_2712,N_24979,N_24849);
xnor UO_2713 (O_2713,N_24872,N_24939);
or UO_2714 (O_2714,N_24976,N_24844);
or UO_2715 (O_2715,N_24895,N_24800);
and UO_2716 (O_2716,N_24966,N_24850);
nor UO_2717 (O_2717,N_24996,N_24808);
or UO_2718 (O_2718,N_24961,N_24859);
and UO_2719 (O_2719,N_24979,N_24993);
xor UO_2720 (O_2720,N_24828,N_24849);
or UO_2721 (O_2721,N_24890,N_24896);
or UO_2722 (O_2722,N_24997,N_24820);
xor UO_2723 (O_2723,N_24926,N_24970);
or UO_2724 (O_2724,N_24858,N_24956);
nand UO_2725 (O_2725,N_24877,N_24892);
nand UO_2726 (O_2726,N_24967,N_24944);
or UO_2727 (O_2727,N_24971,N_24889);
nor UO_2728 (O_2728,N_24805,N_24862);
nor UO_2729 (O_2729,N_24806,N_24902);
nand UO_2730 (O_2730,N_24851,N_24972);
or UO_2731 (O_2731,N_24925,N_24821);
or UO_2732 (O_2732,N_24933,N_24954);
xor UO_2733 (O_2733,N_24855,N_24976);
nand UO_2734 (O_2734,N_24813,N_24903);
and UO_2735 (O_2735,N_24865,N_24910);
nor UO_2736 (O_2736,N_24887,N_24849);
and UO_2737 (O_2737,N_24820,N_24898);
nor UO_2738 (O_2738,N_24939,N_24811);
nand UO_2739 (O_2739,N_24893,N_24878);
nor UO_2740 (O_2740,N_24830,N_24860);
or UO_2741 (O_2741,N_24940,N_24953);
or UO_2742 (O_2742,N_24842,N_24847);
and UO_2743 (O_2743,N_24969,N_24906);
nor UO_2744 (O_2744,N_24840,N_24930);
and UO_2745 (O_2745,N_24989,N_24812);
nand UO_2746 (O_2746,N_24822,N_24912);
nor UO_2747 (O_2747,N_24960,N_24907);
and UO_2748 (O_2748,N_24909,N_24928);
xnor UO_2749 (O_2749,N_24846,N_24973);
xnor UO_2750 (O_2750,N_24923,N_24857);
nand UO_2751 (O_2751,N_24954,N_24822);
nor UO_2752 (O_2752,N_24822,N_24923);
nor UO_2753 (O_2753,N_24999,N_24906);
or UO_2754 (O_2754,N_24801,N_24813);
nor UO_2755 (O_2755,N_24801,N_24947);
nand UO_2756 (O_2756,N_24957,N_24934);
nor UO_2757 (O_2757,N_24846,N_24849);
or UO_2758 (O_2758,N_24819,N_24942);
nor UO_2759 (O_2759,N_24891,N_24971);
nor UO_2760 (O_2760,N_24925,N_24816);
or UO_2761 (O_2761,N_24972,N_24996);
and UO_2762 (O_2762,N_24871,N_24889);
nor UO_2763 (O_2763,N_24951,N_24808);
xnor UO_2764 (O_2764,N_24898,N_24998);
or UO_2765 (O_2765,N_24835,N_24896);
or UO_2766 (O_2766,N_24904,N_24936);
nand UO_2767 (O_2767,N_24989,N_24891);
and UO_2768 (O_2768,N_24849,N_24838);
nand UO_2769 (O_2769,N_24894,N_24917);
nor UO_2770 (O_2770,N_24877,N_24985);
xnor UO_2771 (O_2771,N_24856,N_24960);
and UO_2772 (O_2772,N_24928,N_24908);
xnor UO_2773 (O_2773,N_24805,N_24914);
xor UO_2774 (O_2774,N_24817,N_24838);
or UO_2775 (O_2775,N_24829,N_24879);
nor UO_2776 (O_2776,N_24876,N_24822);
nand UO_2777 (O_2777,N_24995,N_24986);
or UO_2778 (O_2778,N_24978,N_24959);
xnor UO_2779 (O_2779,N_24893,N_24905);
nand UO_2780 (O_2780,N_24945,N_24993);
or UO_2781 (O_2781,N_24822,N_24994);
or UO_2782 (O_2782,N_24895,N_24870);
and UO_2783 (O_2783,N_24992,N_24831);
nand UO_2784 (O_2784,N_24938,N_24939);
or UO_2785 (O_2785,N_24998,N_24999);
nor UO_2786 (O_2786,N_24941,N_24987);
nor UO_2787 (O_2787,N_24865,N_24867);
xnor UO_2788 (O_2788,N_24907,N_24900);
nor UO_2789 (O_2789,N_24932,N_24906);
and UO_2790 (O_2790,N_24890,N_24987);
nor UO_2791 (O_2791,N_24956,N_24854);
and UO_2792 (O_2792,N_24841,N_24948);
and UO_2793 (O_2793,N_24896,N_24899);
and UO_2794 (O_2794,N_24965,N_24980);
nand UO_2795 (O_2795,N_24843,N_24804);
nand UO_2796 (O_2796,N_24913,N_24977);
or UO_2797 (O_2797,N_24973,N_24874);
and UO_2798 (O_2798,N_24838,N_24800);
and UO_2799 (O_2799,N_24991,N_24827);
nand UO_2800 (O_2800,N_24953,N_24906);
nor UO_2801 (O_2801,N_24899,N_24962);
xor UO_2802 (O_2802,N_24930,N_24819);
or UO_2803 (O_2803,N_24947,N_24863);
xor UO_2804 (O_2804,N_24953,N_24848);
or UO_2805 (O_2805,N_24839,N_24801);
nor UO_2806 (O_2806,N_24990,N_24878);
nand UO_2807 (O_2807,N_24852,N_24863);
nand UO_2808 (O_2808,N_24899,N_24947);
or UO_2809 (O_2809,N_24920,N_24874);
nand UO_2810 (O_2810,N_24896,N_24866);
or UO_2811 (O_2811,N_24902,N_24967);
or UO_2812 (O_2812,N_24940,N_24937);
nor UO_2813 (O_2813,N_24977,N_24896);
or UO_2814 (O_2814,N_24921,N_24930);
or UO_2815 (O_2815,N_24828,N_24945);
nor UO_2816 (O_2816,N_24932,N_24942);
or UO_2817 (O_2817,N_24965,N_24909);
nand UO_2818 (O_2818,N_24986,N_24819);
or UO_2819 (O_2819,N_24970,N_24949);
or UO_2820 (O_2820,N_24974,N_24877);
or UO_2821 (O_2821,N_24993,N_24847);
nor UO_2822 (O_2822,N_24896,N_24900);
nand UO_2823 (O_2823,N_24931,N_24909);
and UO_2824 (O_2824,N_24969,N_24947);
nand UO_2825 (O_2825,N_24962,N_24891);
or UO_2826 (O_2826,N_24869,N_24875);
nor UO_2827 (O_2827,N_24994,N_24925);
nand UO_2828 (O_2828,N_24977,N_24846);
nor UO_2829 (O_2829,N_24997,N_24942);
or UO_2830 (O_2830,N_24888,N_24819);
xnor UO_2831 (O_2831,N_24803,N_24835);
nand UO_2832 (O_2832,N_24837,N_24870);
nand UO_2833 (O_2833,N_24930,N_24985);
or UO_2834 (O_2834,N_24903,N_24999);
and UO_2835 (O_2835,N_24873,N_24936);
xor UO_2836 (O_2836,N_24851,N_24957);
and UO_2837 (O_2837,N_24819,N_24984);
or UO_2838 (O_2838,N_24932,N_24912);
xnor UO_2839 (O_2839,N_24993,N_24857);
xnor UO_2840 (O_2840,N_24992,N_24977);
nand UO_2841 (O_2841,N_24913,N_24845);
nand UO_2842 (O_2842,N_24915,N_24839);
or UO_2843 (O_2843,N_24860,N_24984);
and UO_2844 (O_2844,N_24974,N_24958);
xnor UO_2845 (O_2845,N_24930,N_24834);
xnor UO_2846 (O_2846,N_24903,N_24828);
nor UO_2847 (O_2847,N_24903,N_24800);
xnor UO_2848 (O_2848,N_24833,N_24815);
and UO_2849 (O_2849,N_24878,N_24976);
and UO_2850 (O_2850,N_24836,N_24801);
xnor UO_2851 (O_2851,N_24966,N_24897);
nor UO_2852 (O_2852,N_24928,N_24820);
xor UO_2853 (O_2853,N_24977,N_24969);
and UO_2854 (O_2854,N_24922,N_24840);
and UO_2855 (O_2855,N_24895,N_24997);
nand UO_2856 (O_2856,N_24950,N_24978);
xnor UO_2857 (O_2857,N_24852,N_24821);
nand UO_2858 (O_2858,N_24916,N_24899);
and UO_2859 (O_2859,N_24858,N_24959);
nor UO_2860 (O_2860,N_24972,N_24874);
xor UO_2861 (O_2861,N_24839,N_24899);
and UO_2862 (O_2862,N_24904,N_24818);
nor UO_2863 (O_2863,N_24871,N_24964);
nor UO_2864 (O_2864,N_24924,N_24866);
nor UO_2865 (O_2865,N_24920,N_24934);
nand UO_2866 (O_2866,N_24817,N_24839);
nand UO_2867 (O_2867,N_24829,N_24989);
nor UO_2868 (O_2868,N_24812,N_24945);
xor UO_2869 (O_2869,N_24862,N_24916);
nand UO_2870 (O_2870,N_24920,N_24963);
and UO_2871 (O_2871,N_24941,N_24915);
nand UO_2872 (O_2872,N_24874,N_24946);
xor UO_2873 (O_2873,N_24872,N_24972);
nand UO_2874 (O_2874,N_24845,N_24808);
or UO_2875 (O_2875,N_24892,N_24961);
nand UO_2876 (O_2876,N_24978,N_24806);
nand UO_2877 (O_2877,N_24975,N_24950);
xor UO_2878 (O_2878,N_24801,N_24962);
or UO_2879 (O_2879,N_24982,N_24845);
nand UO_2880 (O_2880,N_24870,N_24979);
nand UO_2881 (O_2881,N_24882,N_24846);
xor UO_2882 (O_2882,N_24946,N_24891);
nand UO_2883 (O_2883,N_24953,N_24827);
xnor UO_2884 (O_2884,N_24821,N_24924);
and UO_2885 (O_2885,N_24993,N_24927);
xor UO_2886 (O_2886,N_24901,N_24821);
and UO_2887 (O_2887,N_24972,N_24947);
nor UO_2888 (O_2888,N_24965,N_24903);
xor UO_2889 (O_2889,N_24803,N_24923);
or UO_2890 (O_2890,N_24882,N_24964);
and UO_2891 (O_2891,N_24934,N_24817);
or UO_2892 (O_2892,N_24978,N_24804);
or UO_2893 (O_2893,N_24918,N_24893);
or UO_2894 (O_2894,N_24977,N_24927);
and UO_2895 (O_2895,N_24959,N_24829);
and UO_2896 (O_2896,N_24930,N_24801);
nor UO_2897 (O_2897,N_24925,N_24963);
nand UO_2898 (O_2898,N_24871,N_24864);
or UO_2899 (O_2899,N_24946,N_24908);
or UO_2900 (O_2900,N_24914,N_24804);
nand UO_2901 (O_2901,N_24859,N_24802);
or UO_2902 (O_2902,N_24939,N_24996);
nand UO_2903 (O_2903,N_24834,N_24954);
nand UO_2904 (O_2904,N_24890,N_24916);
xnor UO_2905 (O_2905,N_24873,N_24914);
and UO_2906 (O_2906,N_24844,N_24802);
and UO_2907 (O_2907,N_24849,N_24915);
or UO_2908 (O_2908,N_24876,N_24902);
nand UO_2909 (O_2909,N_24893,N_24919);
nand UO_2910 (O_2910,N_24958,N_24823);
and UO_2911 (O_2911,N_24805,N_24980);
nand UO_2912 (O_2912,N_24829,N_24973);
or UO_2913 (O_2913,N_24890,N_24906);
nor UO_2914 (O_2914,N_24972,N_24892);
xor UO_2915 (O_2915,N_24802,N_24834);
xor UO_2916 (O_2916,N_24816,N_24815);
xor UO_2917 (O_2917,N_24989,N_24863);
or UO_2918 (O_2918,N_24948,N_24999);
nor UO_2919 (O_2919,N_24813,N_24833);
nor UO_2920 (O_2920,N_24920,N_24893);
xnor UO_2921 (O_2921,N_24973,N_24919);
or UO_2922 (O_2922,N_24923,N_24883);
or UO_2923 (O_2923,N_24907,N_24950);
nor UO_2924 (O_2924,N_24853,N_24956);
nor UO_2925 (O_2925,N_24975,N_24962);
or UO_2926 (O_2926,N_24988,N_24975);
nand UO_2927 (O_2927,N_24840,N_24875);
or UO_2928 (O_2928,N_24834,N_24988);
xnor UO_2929 (O_2929,N_24966,N_24972);
nor UO_2930 (O_2930,N_24986,N_24843);
or UO_2931 (O_2931,N_24843,N_24945);
or UO_2932 (O_2932,N_24905,N_24982);
xor UO_2933 (O_2933,N_24946,N_24885);
xor UO_2934 (O_2934,N_24800,N_24944);
and UO_2935 (O_2935,N_24962,N_24931);
nand UO_2936 (O_2936,N_24882,N_24978);
nand UO_2937 (O_2937,N_24961,N_24907);
or UO_2938 (O_2938,N_24896,N_24860);
nor UO_2939 (O_2939,N_24821,N_24934);
nor UO_2940 (O_2940,N_24932,N_24869);
or UO_2941 (O_2941,N_24854,N_24931);
and UO_2942 (O_2942,N_24832,N_24918);
nand UO_2943 (O_2943,N_24888,N_24840);
or UO_2944 (O_2944,N_24828,N_24889);
or UO_2945 (O_2945,N_24993,N_24869);
nor UO_2946 (O_2946,N_24881,N_24927);
or UO_2947 (O_2947,N_24989,N_24821);
or UO_2948 (O_2948,N_24844,N_24943);
nor UO_2949 (O_2949,N_24820,N_24970);
xor UO_2950 (O_2950,N_24984,N_24829);
nor UO_2951 (O_2951,N_24997,N_24940);
and UO_2952 (O_2952,N_24888,N_24868);
xor UO_2953 (O_2953,N_24940,N_24821);
or UO_2954 (O_2954,N_24992,N_24928);
and UO_2955 (O_2955,N_24926,N_24946);
nand UO_2956 (O_2956,N_24853,N_24822);
xor UO_2957 (O_2957,N_24979,N_24921);
nand UO_2958 (O_2958,N_24971,N_24869);
nor UO_2959 (O_2959,N_24954,N_24876);
nand UO_2960 (O_2960,N_24980,N_24844);
nor UO_2961 (O_2961,N_24915,N_24974);
xor UO_2962 (O_2962,N_24849,N_24901);
or UO_2963 (O_2963,N_24870,N_24903);
or UO_2964 (O_2964,N_24846,N_24957);
nand UO_2965 (O_2965,N_24801,N_24846);
and UO_2966 (O_2966,N_24801,N_24809);
and UO_2967 (O_2967,N_24820,N_24887);
or UO_2968 (O_2968,N_24886,N_24984);
xnor UO_2969 (O_2969,N_24867,N_24870);
and UO_2970 (O_2970,N_24953,N_24891);
and UO_2971 (O_2971,N_24868,N_24877);
or UO_2972 (O_2972,N_24864,N_24816);
or UO_2973 (O_2973,N_24829,N_24975);
nor UO_2974 (O_2974,N_24809,N_24829);
nor UO_2975 (O_2975,N_24830,N_24967);
xor UO_2976 (O_2976,N_24857,N_24862);
or UO_2977 (O_2977,N_24924,N_24916);
nand UO_2978 (O_2978,N_24860,N_24811);
nand UO_2979 (O_2979,N_24805,N_24822);
and UO_2980 (O_2980,N_24839,N_24877);
nor UO_2981 (O_2981,N_24829,N_24891);
or UO_2982 (O_2982,N_24813,N_24930);
nor UO_2983 (O_2983,N_24955,N_24894);
nand UO_2984 (O_2984,N_24901,N_24956);
and UO_2985 (O_2985,N_24808,N_24947);
xnor UO_2986 (O_2986,N_24830,N_24813);
or UO_2987 (O_2987,N_24886,N_24859);
nor UO_2988 (O_2988,N_24824,N_24831);
and UO_2989 (O_2989,N_24826,N_24847);
xor UO_2990 (O_2990,N_24882,N_24991);
nor UO_2991 (O_2991,N_24888,N_24900);
xnor UO_2992 (O_2992,N_24883,N_24925);
nor UO_2993 (O_2993,N_24935,N_24939);
xnor UO_2994 (O_2994,N_24871,N_24984);
and UO_2995 (O_2995,N_24987,N_24857);
nor UO_2996 (O_2996,N_24833,N_24809);
nand UO_2997 (O_2997,N_24930,N_24939);
and UO_2998 (O_2998,N_24892,N_24943);
nor UO_2999 (O_2999,N_24873,N_24921);
endmodule