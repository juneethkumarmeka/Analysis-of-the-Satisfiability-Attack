module basic_750_5000_1000_5_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_477,In_736);
nand U1 (N_1,In_270,In_565);
xnor U2 (N_2,In_646,In_570);
or U3 (N_3,In_398,In_380);
nor U4 (N_4,In_702,In_617);
nor U5 (N_5,In_231,In_444);
and U6 (N_6,In_379,In_159);
and U7 (N_7,In_253,In_674);
nor U8 (N_8,In_619,In_557);
xor U9 (N_9,In_337,In_55);
nor U10 (N_10,In_338,In_500);
nor U11 (N_11,In_208,In_3);
nor U12 (N_12,In_598,In_693);
nand U13 (N_13,In_239,In_120);
nand U14 (N_14,In_371,In_490);
nor U15 (N_15,In_236,In_436);
nor U16 (N_16,In_660,In_108);
and U17 (N_17,In_414,In_20);
nor U18 (N_18,In_672,In_165);
and U19 (N_19,In_421,In_321);
and U20 (N_20,In_652,In_378);
or U21 (N_21,In_508,In_536);
nand U22 (N_22,In_48,In_302);
nor U23 (N_23,In_242,In_217);
and U24 (N_24,In_320,In_26);
or U25 (N_25,In_675,In_558);
or U26 (N_26,In_692,In_654);
or U27 (N_27,In_475,In_293);
nand U28 (N_28,In_252,In_211);
nor U29 (N_29,In_527,In_233);
nand U30 (N_30,In_173,In_637);
and U31 (N_31,In_458,In_716);
nor U32 (N_32,In_463,In_435);
nand U33 (N_33,In_132,In_548);
nand U34 (N_34,In_445,In_370);
or U35 (N_35,In_519,In_152);
nand U36 (N_36,In_341,In_709);
xor U37 (N_37,In_656,In_501);
xnor U38 (N_38,In_104,In_461);
nor U39 (N_39,In_474,In_95);
nand U40 (N_40,In_438,In_171);
nor U41 (N_41,In_151,In_535);
nor U42 (N_42,In_417,In_294);
nand U43 (N_43,In_305,In_650);
xor U44 (N_44,In_331,In_110);
and U45 (N_45,In_561,In_45);
and U46 (N_46,In_392,In_624);
and U47 (N_47,In_385,In_591);
and U48 (N_48,In_189,In_142);
nor U49 (N_49,In_114,In_473);
xor U50 (N_50,In_663,In_39);
nor U51 (N_51,In_581,In_54);
nor U52 (N_52,In_595,In_21);
or U53 (N_53,In_453,In_86);
nand U54 (N_54,In_641,In_254);
and U55 (N_55,In_205,In_512);
xnor U56 (N_56,In_323,In_101);
xnor U57 (N_57,In_92,In_122);
xor U58 (N_58,In_734,In_116);
nor U59 (N_59,In_694,In_216);
and U60 (N_60,In_450,In_291);
nor U61 (N_61,In_32,In_618);
nor U62 (N_62,In_166,In_707);
xnor U63 (N_63,In_545,In_249);
nor U64 (N_64,In_287,In_639);
nor U65 (N_65,In_144,In_374);
xor U66 (N_66,In_63,In_9);
and U67 (N_67,In_107,In_203);
or U68 (N_68,In_353,In_313);
or U69 (N_69,In_636,In_213);
and U70 (N_70,In_464,In_14);
nand U71 (N_71,In_13,In_356);
or U72 (N_72,In_629,In_456);
xnor U73 (N_73,In_488,In_739);
and U74 (N_74,In_603,In_185);
xor U75 (N_75,In_533,In_89);
xnor U76 (N_76,In_505,In_257);
nor U77 (N_77,In_585,In_145);
and U78 (N_78,In_19,In_590);
or U79 (N_79,In_292,In_223);
xor U80 (N_80,In_691,In_608);
nand U81 (N_81,In_573,In_564);
or U82 (N_82,In_669,In_429);
nor U83 (N_83,In_404,In_743);
and U84 (N_84,In_224,In_83);
or U85 (N_85,In_43,In_16);
nor U86 (N_86,In_383,In_186);
and U87 (N_87,In_180,In_687);
nor U88 (N_88,In_362,In_727);
or U89 (N_89,In_187,In_470);
nand U90 (N_90,In_497,In_411);
or U91 (N_91,In_266,In_677);
nor U92 (N_92,In_409,In_679);
xnor U93 (N_93,In_218,In_179);
or U94 (N_94,In_296,In_673);
nand U95 (N_95,In_682,In_161);
nor U96 (N_96,In_419,In_626);
nand U97 (N_97,In_431,In_748);
nor U98 (N_98,In_572,In_82);
xor U99 (N_99,In_269,In_345);
xnor U100 (N_100,In_277,In_622);
or U101 (N_101,In_552,In_153);
and U102 (N_102,In_592,In_11);
or U103 (N_103,In_350,In_664);
or U104 (N_104,In_246,In_317);
or U105 (N_105,In_157,In_407);
nand U106 (N_106,In_88,In_480);
nand U107 (N_107,In_715,In_551);
or U108 (N_108,In_125,In_632);
nor U109 (N_109,In_18,In_70);
xor U110 (N_110,In_123,In_128);
and U111 (N_111,In_600,In_538);
and U112 (N_112,In_103,In_507);
nand U113 (N_113,In_457,In_586);
or U114 (N_114,In_683,In_206);
or U115 (N_115,In_469,In_606);
and U116 (N_116,In_587,In_274);
and U117 (N_117,In_271,In_332);
xnor U118 (N_118,In_244,In_631);
and U119 (N_119,In_680,In_405);
xnor U120 (N_120,In_701,In_181);
or U121 (N_121,In_658,In_455);
nor U122 (N_122,In_522,In_136);
xnor U123 (N_123,In_209,In_342);
nand U124 (N_124,In_330,In_708);
nand U125 (N_125,In_403,In_28);
nor U126 (N_126,In_61,In_51);
nor U127 (N_127,In_158,In_476);
nor U128 (N_128,In_521,In_238);
nor U129 (N_129,In_726,In_721);
and U130 (N_130,In_695,In_644);
xnor U131 (N_131,In_413,In_183);
and U132 (N_132,In_35,In_174);
or U133 (N_133,In_381,In_594);
and U134 (N_134,In_465,In_578);
and U135 (N_135,In_229,In_584);
nand U136 (N_136,In_588,In_361);
or U137 (N_137,In_645,In_418);
nand U138 (N_138,In_248,In_127);
or U139 (N_139,In_325,In_719);
nor U140 (N_140,In_495,In_259);
or U141 (N_141,In_279,In_700);
nand U142 (N_142,In_310,In_526);
xnor U143 (N_143,In_577,In_78);
xnor U144 (N_144,In_503,In_201);
xor U145 (N_145,In_191,In_449);
nand U146 (N_146,In_454,In_426);
xnor U147 (N_147,In_138,In_443);
nor U148 (N_148,In_344,In_176);
nor U149 (N_149,In_729,In_569);
nor U150 (N_150,In_499,In_234);
nor U151 (N_151,In_303,In_44);
nand U152 (N_152,In_704,In_684);
or U153 (N_153,In_77,In_485);
or U154 (N_154,In_681,In_738);
xnor U155 (N_155,In_363,In_542);
xnor U156 (N_156,In_697,In_155);
and U157 (N_157,In_64,In_232);
and U158 (N_158,In_498,In_496);
nor U159 (N_159,In_528,In_447);
and U160 (N_160,In_247,In_288);
nand U161 (N_161,In_427,In_327);
xor U162 (N_162,In_264,In_550);
xnor U163 (N_163,In_184,In_525);
nor U164 (N_164,In_459,In_139);
nor U165 (N_165,In_312,In_642);
nand U166 (N_166,In_689,In_52);
or U167 (N_167,In_258,In_75);
or U168 (N_168,In_129,In_532);
and U169 (N_169,In_393,In_7);
xor U170 (N_170,In_59,In_676);
xnor U171 (N_171,In_286,In_448);
or U172 (N_172,In_597,In_517);
nand U173 (N_173,In_0,In_182);
or U174 (N_174,In_657,In_486);
nor U175 (N_175,In_8,In_731);
or U176 (N_176,In_530,In_640);
or U177 (N_177,In_580,In_442);
and U178 (N_178,In_237,In_29);
xor U179 (N_179,In_610,In_214);
or U180 (N_180,In_467,In_333);
nor U181 (N_181,In_339,In_481);
and U182 (N_182,In_699,In_628);
nand U183 (N_183,In_487,In_712);
and U184 (N_184,In_219,In_204);
or U185 (N_185,In_566,In_416);
or U186 (N_186,In_102,In_308);
nor U187 (N_187,In_539,In_424);
or U188 (N_188,In_290,In_670);
xnor U189 (N_189,In_74,In_560);
nand U190 (N_190,In_156,In_100);
xor U191 (N_191,In_627,In_41);
nor U192 (N_192,In_390,In_343);
and U193 (N_193,In_10,In_415);
xor U194 (N_194,In_314,In_135);
nor U195 (N_195,In_170,In_164);
nor U196 (N_196,In_275,In_479);
nor U197 (N_197,In_661,In_131);
nand U198 (N_198,In_620,In_93);
nand U199 (N_199,In_309,In_420);
or U200 (N_200,In_38,In_12);
and U201 (N_201,In_2,In_717);
xnor U202 (N_202,In_80,In_53);
nor U203 (N_203,In_441,In_567);
and U204 (N_204,In_267,In_1);
or U205 (N_205,In_740,In_358);
or U206 (N_206,In_553,In_98);
nor U207 (N_207,In_388,In_169);
or U208 (N_208,In_196,In_79);
xnor U209 (N_209,In_547,In_718);
nand U210 (N_210,In_601,In_384);
and U211 (N_211,In_703,In_730);
xor U212 (N_212,In_732,In_372);
and U213 (N_213,In_579,In_397);
nor U214 (N_214,In_596,In_194);
and U215 (N_215,In_87,In_276);
nor U216 (N_216,In_531,In_112);
or U217 (N_217,In_177,In_66);
and U218 (N_218,In_386,In_630);
nor U219 (N_219,In_199,In_315);
nor U220 (N_220,In_671,In_105);
xor U221 (N_221,In_741,In_147);
xnor U222 (N_222,In_746,In_349);
and U223 (N_223,In_148,In_141);
or U224 (N_224,In_281,In_735);
nand U225 (N_225,In_84,In_555);
xor U226 (N_226,In_364,In_367);
and U227 (N_227,In_278,In_130);
nand U228 (N_228,In_635,In_382);
nor U229 (N_229,In_306,In_160);
nand U230 (N_230,In_50,In_262);
xor U231 (N_231,In_17,In_4);
or U232 (N_232,In_440,In_227);
or U233 (N_233,In_430,In_516);
and U234 (N_234,In_42,In_33);
nor U235 (N_235,In_260,In_376);
or U236 (N_236,In_58,In_605);
nand U237 (N_237,In_690,In_324);
or U238 (N_238,In_94,In_667);
xnor U239 (N_239,In_285,In_520);
nand U240 (N_240,In_513,In_698);
and U241 (N_241,In_614,In_126);
nand U242 (N_242,In_647,In_273);
nand U243 (N_243,In_225,In_328);
nand U244 (N_244,In_462,In_556);
nand U245 (N_245,In_23,In_146);
xnor U246 (N_246,In_576,In_506);
nor U247 (N_247,In_119,In_625);
and U248 (N_248,In_408,In_289);
or U249 (N_249,In_336,In_615);
or U250 (N_250,In_283,In_493);
or U251 (N_251,In_149,In_190);
nand U252 (N_252,In_616,In_210);
nor U253 (N_253,In_478,In_412);
or U254 (N_254,In_651,In_117);
xor U255 (N_255,In_633,In_22);
and U256 (N_256,In_549,In_713);
xnor U257 (N_257,In_401,In_562);
or U258 (N_258,In_534,In_154);
nor U259 (N_259,In_623,In_659);
nor U260 (N_260,In_452,In_282);
and U261 (N_261,In_221,In_192);
nor U262 (N_262,In_583,In_728);
nor U263 (N_263,In_688,In_433);
nor U264 (N_264,In_662,In_256);
or U265 (N_265,In_391,In_347);
xnor U266 (N_266,In_649,In_744);
and U267 (N_267,In_668,In_563);
or U268 (N_268,In_168,In_40);
xnor U269 (N_269,In_255,In_137);
or U270 (N_270,In_696,In_612);
and U271 (N_271,In_428,In_432);
nand U272 (N_272,In_607,In_124);
xor U273 (N_273,In_593,In_472);
nand U274 (N_274,In_73,In_373);
and U275 (N_275,In_178,In_354);
nor U276 (N_276,In_706,In_37);
and U277 (N_277,In_720,In_446);
nand U278 (N_278,In_280,In_742);
and U279 (N_279,In_140,In_106);
nand U280 (N_280,In_471,In_634);
nand U281 (N_281,In_509,In_121);
and U282 (N_282,In_326,In_34);
nor U283 (N_283,In_434,In_396);
nand U284 (N_284,In_163,In_298);
or U285 (N_285,In_143,In_554);
xor U286 (N_286,In_489,In_394);
nand U287 (N_287,In_638,In_60);
nor U288 (N_288,In_46,In_665);
or U289 (N_289,In_423,In_198);
xnor U290 (N_290,In_460,In_263);
or U291 (N_291,In_540,In_439);
and U292 (N_292,In_582,In_91);
or U293 (N_293,In_195,In_523);
and U294 (N_294,In_352,In_643);
nand U295 (N_295,In_511,In_482);
nor U296 (N_296,In_56,In_118);
or U297 (N_297,In_604,In_311);
nand U298 (N_298,In_559,In_133);
or U299 (N_299,In_510,In_574);
nor U300 (N_300,In_24,In_115);
nand U301 (N_301,In_724,In_369);
or U302 (N_302,In_25,In_351);
nor U303 (N_303,In_268,In_395);
or U304 (N_304,In_747,In_514);
or U305 (N_305,In_99,In_334);
or U306 (N_306,In_705,In_723);
or U307 (N_307,In_483,In_749);
nand U308 (N_308,In_722,In_544);
nand U309 (N_309,In_57,In_150);
nand U310 (N_310,In_360,In_389);
nor U311 (N_311,In_272,In_36);
or U312 (N_312,In_737,In_67);
xor U313 (N_313,In_466,In_284);
or U314 (N_314,In_340,In_265);
nor U315 (N_315,In_599,In_492);
or U316 (N_316,In_329,In_611);
or U317 (N_317,In_215,In_243);
xor U318 (N_318,In_322,In_491);
and U319 (N_319,In_15,In_301);
and U320 (N_320,In_241,In_111);
and U321 (N_321,In_113,In_653);
and U322 (N_322,In_134,In_524);
or U323 (N_323,In_76,In_589);
nand U324 (N_324,In_537,In_200);
and U325 (N_325,In_745,In_235);
or U326 (N_326,In_613,In_175);
xor U327 (N_327,In_31,In_68);
nand U328 (N_328,In_47,In_109);
nand U329 (N_329,In_541,In_245);
and U330 (N_330,In_297,In_655);
or U331 (N_331,In_346,In_193);
or U332 (N_332,In_172,In_316);
or U333 (N_333,In_365,In_502);
nor U334 (N_334,In_410,In_299);
or U335 (N_335,In_359,In_733);
xnor U336 (N_336,In_85,In_648);
nand U337 (N_337,In_250,In_240);
nand U338 (N_338,In_81,In_197);
xnor U339 (N_339,In_402,In_504);
nor U340 (N_340,In_678,In_300);
nor U341 (N_341,In_307,In_377);
nand U342 (N_342,In_202,In_725);
xnor U343 (N_343,In_666,In_400);
nor U344 (N_344,In_97,In_71);
nor U345 (N_345,In_621,In_228);
or U346 (N_346,In_30,In_188);
xor U347 (N_347,In_222,In_406);
and U348 (N_348,In_212,In_27);
or U349 (N_349,In_518,In_69);
xnor U350 (N_350,In_251,In_468);
or U351 (N_351,In_529,In_543);
nor U352 (N_352,In_304,In_207);
or U353 (N_353,In_546,In_714);
or U354 (N_354,In_90,In_357);
xor U355 (N_355,In_368,In_6);
and U356 (N_356,In_602,In_261);
nor U357 (N_357,In_568,In_96);
and U358 (N_358,In_226,In_686);
and U359 (N_359,In_437,In_571);
or U360 (N_360,In_494,In_399);
and U361 (N_361,In_710,In_375);
and U362 (N_362,In_609,In_319);
and U363 (N_363,In_49,In_515);
and U364 (N_364,In_65,In_387);
and U365 (N_365,In_162,In_335);
nand U366 (N_366,In_366,In_451);
xnor U367 (N_367,In_355,In_295);
nand U368 (N_368,In_425,In_230);
and U369 (N_369,In_72,In_484);
nand U370 (N_370,In_348,In_167);
or U371 (N_371,In_575,In_711);
nor U372 (N_372,In_62,In_422);
xor U373 (N_373,In_220,In_318);
nand U374 (N_374,In_685,In_5);
nor U375 (N_375,In_514,In_699);
xnor U376 (N_376,In_507,In_582);
nand U377 (N_377,In_206,In_669);
xnor U378 (N_378,In_474,In_47);
or U379 (N_379,In_556,In_332);
nand U380 (N_380,In_530,In_511);
and U381 (N_381,In_425,In_237);
xor U382 (N_382,In_449,In_353);
xor U383 (N_383,In_293,In_154);
or U384 (N_384,In_271,In_653);
and U385 (N_385,In_737,In_484);
xnor U386 (N_386,In_119,In_460);
or U387 (N_387,In_394,In_83);
and U388 (N_388,In_340,In_155);
nor U389 (N_389,In_194,In_51);
and U390 (N_390,In_88,In_692);
or U391 (N_391,In_101,In_467);
nand U392 (N_392,In_415,In_595);
nor U393 (N_393,In_289,In_718);
xor U394 (N_394,In_708,In_729);
nand U395 (N_395,In_141,In_72);
or U396 (N_396,In_548,In_662);
nand U397 (N_397,In_32,In_128);
or U398 (N_398,In_476,In_482);
xnor U399 (N_399,In_310,In_297);
or U400 (N_400,In_650,In_502);
or U401 (N_401,In_372,In_504);
xor U402 (N_402,In_505,In_55);
or U403 (N_403,In_577,In_498);
xnor U404 (N_404,In_55,In_418);
nand U405 (N_405,In_626,In_457);
or U406 (N_406,In_66,In_669);
nor U407 (N_407,In_172,In_226);
nand U408 (N_408,In_403,In_541);
nand U409 (N_409,In_63,In_572);
nor U410 (N_410,In_83,In_529);
and U411 (N_411,In_61,In_734);
nor U412 (N_412,In_732,In_54);
nor U413 (N_413,In_722,In_553);
xnor U414 (N_414,In_256,In_69);
xnor U415 (N_415,In_722,In_217);
xor U416 (N_416,In_500,In_448);
xor U417 (N_417,In_573,In_458);
or U418 (N_418,In_450,In_76);
xor U419 (N_419,In_606,In_236);
and U420 (N_420,In_672,In_267);
nand U421 (N_421,In_58,In_424);
and U422 (N_422,In_92,In_469);
and U423 (N_423,In_26,In_641);
nand U424 (N_424,In_124,In_320);
nor U425 (N_425,In_297,In_270);
and U426 (N_426,In_53,In_38);
nor U427 (N_427,In_50,In_585);
nand U428 (N_428,In_159,In_515);
xor U429 (N_429,In_68,In_674);
xnor U430 (N_430,In_599,In_520);
and U431 (N_431,In_728,In_523);
nor U432 (N_432,In_481,In_489);
and U433 (N_433,In_8,In_117);
nand U434 (N_434,In_155,In_231);
and U435 (N_435,In_433,In_489);
and U436 (N_436,In_611,In_537);
nand U437 (N_437,In_486,In_225);
and U438 (N_438,In_664,In_680);
or U439 (N_439,In_252,In_745);
xor U440 (N_440,In_447,In_636);
xnor U441 (N_441,In_442,In_124);
nand U442 (N_442,In_56,In_631);
nor U443 (N_443,In_694,In_329);
or U444 (N_444,In_739,In_419);
or U445 (N_445,In_269,In_434);
and U446 (N_446,In_386,In_402);
and U447 (N_447,In_147,In_3);
and U448 (N_448,In_257,In_566);
xnor U449 (N_449,In_177,In_14);
or U450 (N_450,In_279,In_126);
nand U451 (N_451,In_296,In_537);
and U452 (N_452,In_127,In_206);
and U453 (N_453,In_50,In_484);
nor U454 (N_454,In_292,In_169);
or U455 (N_455,In_193,In_217);
xnor U456 (N_456,In_563,In_389);
nor U457 (N_457,In_196,In_693);
and U458 (N_458,In_409,In_467);
or U459 (N_459,In_735,In_82);
nor U460 (N_460,In_5,In_198);
and U461 (N_461,In_415,In_679);
xor U462 (N_462,In_621,In_236);
nor U463 (N_463,In_169,In_182);
xnor U464 (N_464,In_290,In_181);
nand U465 (N_465,In_354,In_202);
or U466 (N_466,In_684,In_581);
nor U467 (N_467,In_638,In_239);
or U468 (N_468,In_540,In_696);
and U469 (N_469,In_361,In_342);
or U470 (N_470,In_680,In_249);
and U471 (N_471,In_123,In_125);
and U472 (N_472,In_221,In_742);
or U473 (N_473,In_611,In_334);
or U474 (N_474,In_20,In_16);
or U475 (N_475,In_251,In_664);
and U476 (N_476,In_394,In_481);
xnor U477 (N_477,In_80,In_182);
nor U478 (N_478,In_655,In_378);
nand U479 (N_479,In_496,In_421);
nand U480 (N_480,In_89,In_510);
xnor U481 (N_481,In_705,In_179);
and U482 (N_482,In_749,In_168);
nand U483 (N_483,In_439,In_398);
and U484 (N_484,In_405,In_406);
or U485 (N_485,In_106,In_628);
and U486 (N_486,In_52,In_196);
nand U487 (N_487,In_698,In_13);
or U488 (N_488,In_291,In_377);
nor U489 (N_489,In_534,In_193);
xor U490 (N_490,In_445,In_424);
nor U491 (N_491,In_194,In_524);
or U492 (N_492,In_471,In_155);
xnor U493 (N_493,In_133,In_413);
or U494 (N_494,In_376,In_461);
nor U495 (N_495,In_439,In_443);
nor U496 (N_496,In_736,In_392);
or U497 (N_497,In_33,In_377);
or U498 (N_498,In_154,In_361);
and U499 (N_499,In_269,In_241);
nand U500 (N_500,In_611,In_374);
and U501 (N_501,In_652,In_192);
nor U502 (N_502,In_242,In_168);
nor U503 (N_503,In_430,In_136);
or U504 (N_504,In_260,In_25);
and U505 (N_505,In_222,In_16);
nor U506 (N_506,In_431,In_645);
and U507 (N_507,In_572,In_347);
nor U508 (N_508,In_36,In_658);
or U509 (N_509,In_649,In_564);
nand U510 (N_510,In_285,In_434);
and U511 (N_511,In_737,In_37);
nand U512 (N_512,In_484,In_570);
and U513 (N_513,In_247,In_63);
and U514 (N_514,In_602,In_452);
and U515 (N_515,In_117,In_39);
or U516 (N_516,In_588,In_515);
nor U517 (N_517,In_482,In_343);
nor U518 (N_518,In_586,In_184);
nor U519 (N_519,In_187,In_338);
or U520 (N_520,In_97,In_698);
nand U521 (N_521,In_406,In_360);
nor U522 (N_522,In_643,In_447);
xor U523 (N_523,In_688,In_289);
or U524 (N_524,In_280,In_568);
nand U525 (N_525,In_586,In_666);
nor U526 (N_526,In_651,In_273);
nand U527 (N_527,In_153,In_475);
or U528 (N_528,In_338,In_122);
or U529 (N_529,In_503,In_497);
and U530 (N_530,In_164,In_619);
and U531 (N_531,In_318,In_268);
or U532 (N_532,In_36,In_293);
xor U533 (N_533,In_195,In_681);
nand U534 (N_534,In_553,In_469);
or U535 (N_535,In_407,In_408);
nand U536 (N_536,In_5,In_659);
nor U537 (N_537,In_113,In_735);
and U538 (N_538,In_709,In_299);
nand U539 (N_539,In_95,In_617);
or U540 (N_540,In_93,In_10);
or U541 (N_541,In_121,In_156);
xor U542 (N_542,In_732,In_185);
nand U543 (N_543,In_243,In_587);
or U544 (N_544,In_585,In_413);
or U545 (N_545,In_293,In_357);
and U546 (N_546,In_426,In_78);
or U547 (N_547,In_310,In_498);
nor U548 (N_548,In_490,In_382);
or U549 (N_549,In_448,In_89);
and U550 (N_550,In_599,In_457);
xor U551 (N_551,In_224,In_743);
xnor U552 (N_552,In_5,In_102);
and U553 (N_553,In_69,In_403);
and U554 (N_554,In_281,In_459);
or U555 (N_555,In_630,In_253);
or U556 (N_556,In_482,In_576);
nand U557 (N_557,In_403,In_219);
nor U558 (N_558,In_407,In_253);
nand U559 (N_559,In_438,In_105);
nor U560 (N_560,In_438,In_370);
xnor U561 (N_561,In_259,In_160);
nand U562 (N_562,In_276,In_84);
and U563 (N_563,In_680,In_398);
or U564 (N_564,In_539,In_264);
xnor U565 (N_565,In_186,In_267);
or U566 (N_566,In_232,In_335);
nor U567 (N_567,In_308,In_95);
nor U568 (N_568,In_204,In_207);
or U569 (N_569,In_274,In_428);
nand U570 (N_570,In_391,In_213);
nand U571 (N_571,In_263,In_487);
or U572 (N_572,In_669,In_351);
nand U573 (N_573,In_312,In_23);
or U574 (N_574,In_91,In_51);
xnor U575 (N_575,In_103,In_308);
nor U576 (N_576,In_484,In_178);
nand U577 (N_577,In_135,In_590);
nor U578 (N_578,In_456,In_378);
and U579 (N_579,In_122,In_25);
nor U580 (N_580,In_372,In_536);
nor U581 (N_581,In_464,In_596);
xor U582 (N_582,In_94,In_596);
or U583 (N_583,In_582,In_82);
nand U584 (N_584,In_342,In_118);
nor U585 (N_585,In_593,In_142);
xnor U586 (N_586,In_380,In_745);
nor U587 (N_587,In_498,In_204);
and U588 (N_588,In_74,In_493);
and U589 (N_589,In_683,In_335);
nand U590 (N_590,In_719,In_617);
or U591 (N_591,In_436,In_359);
or U592 (N_592,In_654,In_639);
or U593 (N_593,In_151,In_457);
nand U594 (N_594,In_317,In_39);
nand U595 (N_595,In_368,In_270);
xor U596 (N_596,In_478,In_460);
nor U597 (N_597,In_258,In_206);
nand U598 (N_598,In_472,In_139);
or U599 (N_599,In_593,In_202);
or U600 (N_600,In_729,In_544);
nor U601 (N_601,In_348,In_202);
xor U602 (N_602,In_270,In_382);
nor U603 (N_603,In_681,In_109);
nor U604 (N_604,In_10,In_683);
and U605 (N_605,In_250,In_168);
nor U606 (N_606,In_493,In_120);
xnor U607 (N_607,In_395,In_481);
xnor U608 (N_608,In_736,In_109);
and U609 (N_609,In_408,In_585);
xor U610 (N_610,In_152,In_515);
and U611 (N_611,In_644,In_475);
xor U612 (N_612,In_421,In_153);
nor U613 (N_613,In_514,In_613);
or U614 (N_614,In_220,In_331);
or U615 (N_615,In_133,In_499);
xor U616 (N_616,In_285,In_447);
xnor U617 (N_617,In_160,In_125);
nor U618 (N_618,In_508,In_411);
nand U619 (N_619,In_33,In_191);
nor U620 (N_620,In_587,In_442);
or U621 (N_621,In_200,In_225);
or U622 (N_622,In_563,In_495);
nand U623 (N_623,In_216,In_529);
xor U624 (N_624,In_236,In_656);
or U625 (N_625,In_251,In_390);
nand U626 (N_626,In_587,In_78);
and U627 (N_627,In_413,In_607);
nor U628 (N_628,In_362,In_333);
nor U629 (N_629,In_691,In_114);
nor U630 (N_630,In_728,In_571);
xnor U631 (N_631,In_215,In_618);
xor U632 (N_632,In_142,In_447);
nand U633 (N_633,In_680,In_287);
and U634 (N_634,In_686,In_294);
nand U635 (N_635,In_234,In_52);
xor U636 (N_636,In_693,In_141);
xnor U637 (N_637,In_43,In_702);
nor U638 (N_638,In_285,In_377);
and U639 (N_639,In_472,In_132);
or U640 (N_640,In_13,In_377);
or U641 (N_641,In_529,In_287);
nand U642 (N_642,In_637,In_350);
nor U643 (N_643,In_271,In_198);
nand U644 (N_644,In_107,In_144);
nand U645 (N_645,In_309,In_462);
nor U646 (N_646,In_292,In_653);
xor U647 (N_647,In_116,In_541);
nor U648 (N_648,In_460,In_240);
nor U649 (N_649,In_161,In_102);
xnor U650 (N_650,In_409,In_694);
nand U651 (N_651,In_67,In_34);
and U652 (N_652,In_500,In_182);
nor U653 (N_653,In_249,In_655);
and U654 (N_654,In_420,In_267);
nand U655 (N_655,In_302,In_244);
or U656 (N_656,In_123,In_700);
or U657 (N_657,In_714,In_560);
xnor U658 (N_658,In_10,In_16);
nand U659 (N_659,In_1,In_19);
or U660 (N_660,In_631,In_722);
xor U661 (N_661,In_490,In_620);
nand U662 (N_662,In_387,In_440);
xor U663 (N_663,In_614,In_177);
and U664 (N_664,In_330,In_191);
xor U665 (N_665,In_215,In_638);
xnor U666 (N_666,In_712,In_336);
nor U667 (N_667,In_539,In_114);
nor U668 (N_668,In_111,In_623);
xnor U669 (N_669,In_64,In_94);
xnor U670 (N_670,In_462,In_135);
nor U671 (N_671,In_726,In_181);
nor U672 (N_672,In_624,In_1);
nand U673 (N_673,In_180,In_483);
nand U674 (N_674,In_713,In_347);
nor U675 (N_675,In_619,In_676);
nor U676 (N_676,In_291,In_139);
or U677 (N_677,In_741,In_744);
xnor U678 (N_678,In_139,In_263);
nand U679 (N_679,In_701,In_421);
and U680 (N_680,In_735,In_736);
and U681 (N_681,In_2,In_287);
or U682 (N_682,In_281,In_257);
or U683 (N_683,In_163,In_398);
or U684 (N_684,In_355,In_216);
and U685 (N_685,In_396,In_347);
nand U686 (N_686,In_185,In_139);
nor U687 (N_687,In_644,In_367);
and U688 (N_688,In_635,In_747);
nand U689 (N_689,In_6,In_536);
nand U690 (N_690,In_726,In_349);
xor U691 (N_691,In_18,In_240);
xor U692 (N_692,In_371,In_501);
nand U693 (N_693,In_369,In_361);
or U694 (N_694,In_57,In_99);
and U695 (N_695,In_222,In_418);
or U696 (N_696,In_31,In_649);
nor U697 (N_697,In_463,In_323);
nand U698 (N_698,In_49,In_324);
nand U699 (N_699,In_660,In_715);
and U700 (N_700,In_555,In_201);
or U701 (N_701,In_655,In_243);
and U702 (N_702,In_170,In_196);
and U703 (N_703,In_472,In_292);
or U704 (N_704,In_377,In_49);
nor U705 (N_705,In_240,In_663);
nand U706 (N_706,In_15,In_709);
and U707 (N_707,In_599,In_589);
and U708 (N_708,In_87,In_267);
and U709 (N_709,In_231,In_69);
or U710 (N_710,In_110,In_106);
nor U711 (N_711,In_224,In_745);
nand U712 (N_712,In_94,In_84);
nand U713 (N_713,In_704,In_730);
xnor U714 (N_714,In_617,In_589);
xor U715 (N_715,In_716,In_526);
xor U716 (N_716,In_448,In_562);
or U717 (N_717,In_688,In_455);
and U718 (N_718,In_636,In_105);
nor U719 (N_719,In_270,In_223);
nor U720 (N_720,In_380,In_564);
nor U721 (N_721,In_520,In_642);
xnor U722 (N_722,In_336,In_319);
and U723 (N_723,In_730,In_645);
nand U724 (N_724,In_360,In_201);
xor U725 (N_725,In_195,In_273);
xor U726 (N_726,In_632,In_401);
and U727 (N_727,In_714,In_31);
xor U728 (N_728,In_359,In_497);
and U729 (N_729,In_695,In_407);
or U730 (N_730,In_652,In_713);
nand U731 (N_731,In_641,In_730);
xnor U732 (N_732,In_412,In_638);
and U733 (N_733,In_601,In_630);
xor U734 (N_734,In_407,In_538);
nor U735 (N_735,In_139,In_546);
nand U736 (N_736,In_668,In_81);
or U737 (N_737,In_551,In_528);
nand U738 (N_738,In_621,In_449);
nand U739 (N_739,In_635,In_699);
xor U740 (N_740,In_212,In_666);
nor U741 (N_741,In_655,In_397);
xnor U742 (N_742,In_743,In_562);
nor U743 (N_743,In_443,In_251);
or U744 (N_744,In_3,In_68);
or U745 (N_745,In_119,In_226);
or U746 (N_746,In_383,In_117);
or U747 (N_747,In_271,In_131);
nand U748 (N_748,In_92,In_12);
nor U749 (N_749,In_409,In_236);
nor U750 (N_750,In_42,In_145);
or U751 (N_751,In_33,In_66);
xor U752 (N_752,In_173,In_237);
or U753 (N_753,In_66,In_610);
or U754 (N_754,In_330,In_215);
and U755 (N_755,In_363,In_19);
and U756 (N_756,In_118,In_557);
nand U757 (N_757,In_481,In_732);
and U758 (N_758,In_381,In_648);
and U759 (N_759,In_564,In_395);
or U760 (N_760,In_381,In_260);
or U761 (N_761,In_310,In_587);
nand U762 (N_762,In_585,In_459);
and U763 (N_763,In_623,In_388);
xnor U764 (N_764,In_731,In_553);
and U765 (N_765,In_490,In_572);
or U766 (N_766,In_499,In_167);
nand U767 (N_767,In_352,In_337);
or U768 (N_768,In_268,In_316);
and U769 (N_769,In_152,In_472);
xor U770 (N_770,In_734,In_323);
xnor U771 (N_771,In_378,In_388);
nand U772 (N_772,In_579,In_417);
nand U773 (N_773,In_173,In_313);
or U774 (N_774,In_251,In_430);
xor U775 (N_775,In_568,In_149);
nand U776 (N_776,In_611,In_182);
and U777 (N_777,In_289,In_618);
nand U778 (N_778,In_112,In_246);
and U779 (N_779,In_79,In_59);
nor U780 (N_780,In_312,In_84);
or U781 (N_781,In_119,In_221);
or U782 (N_782,In_120,In_655);
xor U783 (N_783,In_669,In_440);
xor U784 (N_784,In_31,In_49);
or U785 (N_785,In_156,In_475);
xor U786 (N_786,In_347,In_35);
and U787 (N_787,In_535,In_422);
and U788 (N_788,In_725,In_268);
or U789 (N_789,In_466,In_271);
xnor U790 (N_790,In_294,In_252);
or U791 (N_791,In_746,In_638);
and U792 (N_792,In_705,In_238);
or U793 (N_793,In_547,In_331);
or U794 (N_794,In_627,In_638);
xnor U795 (N_795,In_34,In_724);
nor U796 (N_796,In_618,In_111);
and U797 (N_797,In_469,In_60);
xnor U798 (N_798,In_69,In_730);
and U799 (N_799,In_595,In_702);
and U800 (N_800,In_455,In_431);
nor U801 (N_801,In_403,In_661);
and U802 (N_802,In_706,In_171);
nand U803 (N_803,In_582,In_558);
xnor U804 (N_804,In_15,In_729);
xnor U805 (N_805,In_361,In_385);
xnor U806 (N_806,In_696,In_721);
and U807 (N_807,In_652,In_549);
and U808 (N_808,In_19,In_729);
nor U809 (N_809,In_301,In_583);
or U810 (N_810,In_215,In_453);
nor U811 (N_811,In_567,In_477);
xnor U812 (N_812,In_438,In_146);
or U813 (N_813,In_125,In_18);
nand U814 (N_814,In_354,In_639);
and U815 (N_815,In_301,In_302);
nor U816 (N_816,In_528,In_165);
or U817 (N_817,In_688,In_709);
xor U818 (N_818,In_502,In_736);
and U819 (N_819,In_667,In_660);
or U820 (N_820,In_454,In_408);
xor U821 (N_821,In_584,In_441);
and U822 (N_822,In_466,In_157);
xor U823 (N_823,In_142,In_124);
or U824 (N_824,In_574,In_443);
xnor U825 (N_825,In_192,In_305);
nor U826 (N_826,In_391,In_582);
nand U827 (N_827,In_214,In_675);
nand U828 (N_828,In_133,In_317);
and U829 (N_829,In_105,In_661);
and U830 (N_830,In_108,In_575);
or U831 (N_831,In_187,In_471);
xnor U832 (N_832,In_315,In_519);
or U833 (N_833,In_55,In_241);
nor U834 (N_834,In_607,In_85);
nand U835 (N_835,In_525,In_557);
or U836 (N_836,In_610,In_474);
and U837 (N_837,In_14,In_611);
and U838 (N_838,In_11,In_336);
and U839 (N_839,In_446,In_627);
or U840 (N_840,In_256,In_60);
nand U841 (N_841,In_60,In_682);
or U842 (N_842,In_71,In_706);
or U843 (N_843,In_704,In_379);
nor U844 (N_844,In_380,In_583);
nor U845 (N_845,In_32,In_476);
nand U846 (N_846,In_329,In_402);
xor U847 (N_847,In_1,In_106);
and U848 (N_848,In_237,In_589);
or U849 (N_849,In_407,In_136);
nor U850 (N_850,In_473,In_402);
nor U851 (N_851,In_273,In_394);
nand U852 (N_852,In_712,In_728);
xor U853 (N_853,In_44,In_591);
and U854 (N_854,In_301,In_731);
xor U855 (N_855,In_48,In_543);
or U856 (N_856,In_658,In_456);
and U857 (N_857,In_12,In_242);
nor U858 (N_858,In_393,In_71);
nand U859 (N_859,In_412,In_471);
nor U860 (N_860,In_484,In_181);
and U861 (N_861,In_137,In_290);
nand U862 (N_862,In_538,In_616);
and U863 (N_863,In_471,In_271);
xor U864 (N_864,In_100,In_115);
or U865 (N_865,In_54,In_145);
nand U866 (N_866,In_720,In_385);
and U867 (N_867,In_195,In_705);
or U868 (N_868,In_14,In_433);
xnor U869 (N_869,In_418,In_462);
and U870 (N_870,In_606,In_51);
or U871 (N_871,In_740,In_730);
nor U872 (N_872,In_307,In_352);
nor U873 (N_873,In_719,In_207);
or U874 (N_874,In_216,In_693);
nor U875 (N_875,In_555,In_390);
nand U876 (N_876,In_418,In_16);
or U877 (N_877,In_739,In_666);
nor U878 (N_878,In_21,In_264);
xor U879 (N_879,In_42,In_740);
or U880 (N_880,In_52,In_743);
nor U881 (N_881,In_609,In_300);
nand U882 (N_882,In_372,In_327);
nand U883 (N_883,In_75,In_113);
nand U884 (N_884,In_567,In_374);
nand U885 (N_885,In_595,In_308);
nor U886 (N_886,In_349,In_661);
or U887 (N_887,In_575,In_168);
or U888 (N_888,In_42,In_672);
or U889 (N_889,In_526,In_334);
nand U890 (N_890,In_567,In_687);
nand U891 (N_891,In_327,In_318);
xor U892 (N_892,In_108,In_554);
xor U893 (N_893,In_560,In_317);
nor U894 (N_894,In_636,In_343);
xor U895 (N_895,In_745,In_663);
xor U896 (N_896,In_182,In_584);
and U897 (N_897,In_307,In_410);
or U898 (N_898,In_673,In_424);
nor U899 (N_899,In_657,In_165);
and U900 (N_900,In_667,In_592);
nor U901 (N_901,In_541,In_558);
xor U902 (N_902,In_211,In_656);
or U903 (N_903,In_320,In_591);
and U904 (N_904,In_38,In_425);
nor U905 (N_905,In_140,In_568);
nand U906 (N_906,In_155,In_75);
xor U907 (N_907,In_443,In_268);
or U908 (N_908,In_484,In_693);
nand U909 (N_909,In_233,In_640);
xor U910 (N_910,In_375,In_689);
nor U911 (N_911,In_14,In_401);
or U912 (N_912,In_438,In_361);
nor U913 (N_913,In_228,In_574);
or U914 (N_914,In_678,In_358);
nand U915 (N_915,In_323,In_582);
nor U916 (N_916,In_306,In_639);
and U917 (N_917,In_667,In_170);
xnor U918 (N_918,In_182,In_748);
and U919 (N_919,In_70,In_577);
nand U920 (N_920,In_662,In_595);
xor U921 (N_921,In_699,In_311);
nand U922 (N_922,In_726,In_96);
nor U923 (N_923,In_402,In_622);
nand U924 (N_924,In_539,In_58);
nor U925 (N_925,In_273,In_217);
nor U926 (N_926,In_688,In_548);
or U927 (N_927,In_556,In_284);
or U928 (N_928,In_180,In_312);
nor U929 (N_929,In_422,In_380);
nor U930 (N_930,In_150,In_476);
and U931 (N_931,In_274,In_401);
and U932 (N_932,In_285,In_61);
xnor U933 (N_933,In_643,In_41);
or U934 (N_934,In_6,In_741);
or U935 (N_935,In_410,In_733);
nand U936 (N_936,In_433,In_402);
nor U937 (N_937,In_399,In_115);
xor U938 (N_938,In_590,In_448);
or U939 (N_939,In_62,In_73);
nand U940 (N_940,In_60,In_548);
nor U941 (N_941,In_143,In_175);
and U942 (N_942,In_77,In_349);
xnor U943 (N_943,In_50,In_296);
nor U944 (N_944,In_495,In_231);
nand U945 (N_945,In_549,In_366);
nor U946 (N_946,In_272,In_678);
and U947 (N_947,In_579,In_396);
nand U948 (N_948,In_7,In_529);
or U949 (N_949,In_434,In_440);
nor U950 (N_950,In_724,In_360);
and U951 (N_951,In_436,In_251);
nand U952 (N_952,In_674,In_10);
nand U953 (N_953,In_560,In_157);
xor U954 (N_954,In_368,In_145);
and U955 (N_955,In_591,In_481);
and U956 (N_956,In_578,In_289);
nor U957 (N_957,In_655,In_288);
nor U958 (N_958,In_185,In_74);
or U959 (N_959,In_281,In_39);
xnor U960 (N_960,In_200,In_383);
and U961 (N_961,In_190,In_597);
nor U962 (N_962,In_357,In_290);
nand U963 (N_963,In_139,In_677);
and U964 (N_964,In_692,In_296);
xnor U965 (N_965,In_469,In_150);
nand U966 (N_966,In_553,In_264);
or U967 (N_967,In_641,In_718);
nand U968 (N_968,In_494,In_719);
or U969 (N_969,In_655,In_498);
nor U970 (N_970,In_88,In_562);
or U971 (N_971,In_696,In_69);
nand U972 (N_972,In_76,In_103);
or U973 (N_973,In_231,In_242);
nor U974 (N_974,In_440,In_620);
xnor U975 (N_975,In_215,In_591);
nor U976 (N_976,In_322,In_735);
xor U977 (N_977,In_86,In_680);
xor U978 (N_978,In_586,In_165);
and U979 (N_979,In_553,In_209);
and U980 (N_980,In_643,In_624);
nor U981 (N_981,In_172,In_324);
nand U982 (N_982,In_450,In_444);
and U983 (N_983,In_273,In_462);
xnor U984 (N_984,In_682,In_581);
nor U985 (N_985,In_206,In_662);
nand U986 (N_986,In_565,In_654);
nand U987 (N_987,In_398,In_543);
nand U988 (N_988,In_112,In_43);
nor U989 (N_989,In_641,In_529);
xnor U990 (N_990,In_644,In_614);
nor U991 (N_991,In_231,In_16);
or U992 (N_992,In_144,In_288);
nor U993 (N_993,In_256,In_332);
or U994 (N_994,In_710,In_298);
or U995 (N_995,In_96,In_316);
nand U996 (N_996,In_8,In_97);
and U997 (N_997,In_165,In_356);
or U998 (N_998,In_140,In_4);
nand U999 (N_999,In_148,In_481);
nand U1000 (N_1000,N_938,N_82);
nor U1001 (N_1001,N_507,N_640);
and U1002 (N_1002,N_733,N_496);
nor U1003 (N_1003,N_371,N_296);
xnor U1004 (N_1004,N_59,N_861);
xor U1005 (N_1005,N_977,N_990);
and U1006 (N_1006,N_577,N_474);
xor U1007 (N_1007,N_94,N_58);
nor U1008 (N_1008,N_659,N_319);
and U1009 (N_1009,N_83,N_948);
xor U1010 (N_1010,N_501,N_802);
xnor U1011 (N_1011,N_596,N_553);
nand U1012 (N_1012,N_744,N_632);
nand U1013 (N_1013,N_687,N_548);
nand U1014 (N_1014,N_105,N_634);
nor U1015 (N_1015,N_79,N_0);
nand U1016 (N_1016,N_797,N_865);
nor U1017 (N_1017,N_897,N_809);
and U1018 (N_1018,N_901,N_737);
and U1019 (N_1019,N_48,N_668);
nor U1020 (N_1020,N_346,N_651);
xor U1021 (N_1021,N_525,N_671);
or U1022 (N_1022,N_870,N_568);
and U1023 (N_1023,N_199,N_884);
or U1024 (N_1024,N_88,N_110);
nand U1025 (N_1025,N_402,N_449);
and U1026 (N_1026,N_421,N_223);
xor U1027 (N_1027,N_149,N_180);
and U1028 (N_1028,N_476,N_799);
and U1029 (N_1029,N_647,N_258);
xnor U1030 (N_1030,N_335,N_812);
xnor U1031 (N_1031,N_282,N_782);
or U1032 (N_1032,N_114,N_805);
xor U1033 (N_1033,N_593,N_838);
nor U1034 (N_1034,N_516,N_313);
or U1035 (N_1035,N_871,N_993);
xor U1036 (N_1036,N_530,N_646);
nor U1037 (N_1037,N_173,N_312);
and U1038 (N_1038,N_228,N_832);
and U1039 (N_1039,N_610,N_849);
nand U1040 (N_1040,N_1,N_906);
xnor U1041 (N_1041,N_450,N_243);
xnor U1042 (N_1042,N_112,N_852);
or U1043 (N_1043,N_144,N_187);
nand U1044 (N_1044,N_4,N_947);
and U1045 (N_1045,N_473,N_834);
nand U1046 (N_1046,N_379,N_193);
or U1047 (N_1047,N_281,N_480);
and U1048 (N_1048,N_196,N_249);
and U1049 (N_1049,N_381,N_669);
nand U1050 (N_1050,N_815,N_287);
and U1051 (N_1051,N_700,N_750);
nor U1052 (N_1052,N_975,N_418);
xnor U1053 (N_1053,N_814,N_683);
and U1054 (N_1054,N_686,N_195);
nand U1055 (N_1055,N_494,N_134);
nor U1056 (N_1056,N_210,N_68);
xnor U1057 (N_1057,N_888,N_298);
xnor U1058 (N_1058,N_625,N_984);
nand U1059 (N_1059,N_150,N_587);
nand U1060 (N_1060,N_672,N_181);
nor U1061 (N_1061,N_177,N_122);
or U1062 (N_1062,N_344,N_622);
or U1063 (N_1063,N_562,N_30);
xor U1064 (N_1064,N_775,N_257);
xor U1065 (N_1065,N_445,N_332);
nor U1066 (N_1066,N_305,N_950);
nand U1067 (N_1067,N_845,N_104);
or U1068 (N_1068,N_855,N_23);
nand U1069 (N_1069,N_154,N_486);
or U1070 (N_1070,N_125,N_503);
nor U1071 (N_1071,N_167,N_835);
xor U1072 (N_1072,N_179,N_760);
and U1073 (N_1073,N_369,N_616);
or U1074 (N_1074,N_570,N_469);
nor U1075 (N_1075,N_263,N_495);
nand U1076 (N_1076,N_464,N_168);
and U1077 (N_1077,N_475,N_617);
and U1078 (N_1078,N_505,N_752);
nand U1079 (N_1079,N_270,N_423);
xor U1080 (N_1080,N_726,N_292);
nor U1081 (N_1081,N_841,N_138);
or U1082 (N_1082,N_771,N_801);
and U1083 (N_1083,N_631,N_293);
or U1084 (N_1084,N_766,N_793);
xor U1085 (N_1085,N_624,N_183);
and U1086 (N_1086,N_370,N_716);
nand U1087 (N_1087,N_970,N_818);
or U1088 (N_1088,N_595,N_27);
nor U1089 (N_1089,N_946,N_719);
or U1090 (N_1090,N_119,N_356);
xor U1091 (N_1091,N_635,N_512);
xnor U1092 (N_1092,N_283,N_951);
nor U1093 (N_1093,N_848,N_483);
xor U1094 (N_1094,N_885,N_958);
or U1095 (N_1095,N_869,N_19);
and U1096 (N_1096,N_803,N_35);
nand U1097 (N_1097,N_859,N_277);
nor U1098 (N_1098,N_485,N_117);
xnor U1099 (N_1099,N_666,N_656);
and U1100 (N_1100,N_755,N_32);
or U1101 (N_1101,N_482,N_31);
nor U1102 (N_1102,N_236,N_256);
nand U1103 (N_1103,N_215,N_408);
and U1104 (N_1104,N_499,N_101);
and U1105 (N_1105,N_202,N_996);
nand U1106 (N_1106,N_93,N_365);
or U1107 (N_1107,N_247,N_235);
nor U1108 (N_1108,N_537,N_890);
nand U1109 (N_1109,N_761,N_601);
or U1110 (N_1110,N_91,N_80);
nand U1111 (N_1111,N_866,N_633);
nand U1112 (N_1112,N_376,N_390);
nand U1113 (N_1113,N_739,N_234);
nor U1114 (N_1114,N_410,N_52);
nand U1115 (N_1115,N_265,N_787);
or U1116 (N_1116,N_62,N_437);
nand U1117 (N_1117,N_969,N_364);
xor U1118 (N_1118,N_693,N_362);
xor U1119 (N_1119,N_38,N_205);
nor U1120 (N_1120,N_338,N_20);
nand U1121 (N_1121,N_627,N_268);
and U1122 (N_1122,N_417,N_567);
xnor U1123 (N_1123,N_456,N_533);
nor U1124 (N_1124,N_978,N_422);
and U1125 (N_1125,N_269,N_128);
xor U1126 (N_1126,N_862,N_842);
and U1127 (N_1127,N_974,N_189);
and U1128 (N_1128,N_73,N_334);
or U1129 (N_1129,N_17,N_148);
nor U1130 (N_1130,N_614,N_513);
nor U1131 (N_1131,N_560,N_384);
xor U1132 (N_1132,N_307,N_341);
xor U1133 (N_1133,N_166,N_743);
xor U1134 (N_1134,N_571,N_825);
xor U1135 (N_1135,N_13,N_591);
nand U1136 (N_1136,N_481,N_358);
or U1137 (N_1137,N_574,N_826);
nand U1138 (N_1138,N_100,N_979);
nor U1139 (N_1139,N_392,N_213);
and U1140 (N_1140,N_345,N_688);
xnor U1141 (N_1141,N_251,N_140);
xor U1142 (N_1142,N_352,N_290);
or U1143 (N_1143,N_426,N_230);
xnor U1144 (N_1144,N_65,N_881);
nor U1145 (N_1145,N_526,N_924);
nand U1146 (N_1146,N_2,N_331);
nor U1147 (N_1147,N_113,N_465);
or U1148 (N_1148,N_323,N_718);
or U1149 (N_1149,N_203,N_244);
xnor U1150 (N_1150,N_300,N_78);
nor U1151 (N_1151,N_51,N_639);
or U1152 (N_1152,N_880,N_252);
and U1153 (N_1153,N_34,N_543);
xor U1154 (N_1154,N_831,N_657);
and U1155 (N_1155,N_648,N_808);
nand U1156 (N_1156,N_549,N_92);
xnor U1157 (N_1157,N_925,N_147);
and U1158 (N_1158,N_676,N_642);
and U1159 (N_1159,N_403,N_877);
xnor U1160 (N_1160,N_583,N_337);
nand U1161 (N_1161,N_348,N_145);
or U1162 (N_1162,N_891,N_679);
nand U1163 (N_1163,N_488,N_57);
nand U1164 (N_1164,N_777,N_790);
or U1165 (N_1165,N_538,N_299);
or U1166 (N_1166,N_40,N_798);
and U1167 (N_1167,N_608,N_724);
xor U1168 (N_1168,N_414,N_689);
and U1169 (N_1169,N_791,N_372);
nor U1170 (N_1170,N_347,N_532);
nor U1171 (N_1171,N_830,N_33);
xnor U1172 (N_1172,N_603,N_261);
or U1173 (N_1173,N_912,N_455);
or U1174 (N_1174,N_53,N_661);
nand U1175 (N_1175,N_222,N_111);
nor U1176 (N_1176,N_515,N_673);
nor U1177 (N_1177,N_441,N_204);
xnor U1178 (N_1178,N_190,N_836);
nor U1179 (N_1179,N_121,N_50);
xor U1180 (N_1180,N_262,N_663);
or U1181 (N_1181,N_206,N_468);
or U1182 (N_1182,N_594,N_157);
nand U1183 (N_1183,N_734,N_741);
xor U1184 (N_1184,N_641,N_588);
or U1185 (N_1185,N_905,N_774);
nand U1186 (N_1186,N_662,N_697);
xor U1187 (N_1187,N_927,N_493);
nand U1188 (N_1188,N_813,N_564);
or U1189 (N_1189,N_238,N_514);
nor U1190 (N_1190,N_442,N_887);
and U1191 (N_1191,N_250,N_382);
nor U1192 (N_1192,N_922,N_288);
xor U1193 (N_1193,N_178,N_188);
or U1194 (N_1194,N_18,N_174);
nor U1195 (N_1195,N_615,N_619);
nand U1196 (N_1196,N_872,N_172);
and U1197 (N_1197,N_366,N_573);
or U1198 (N_1198,N_611,N_637);
or U1199 (N_1199,N_318,N_458);
and U1200 (N_1200,N_966,N_321);
xor U1201 (N_1201,N_999,N_440);
nand U1202 (N_1202,N_191,N_267);
and U1203 (N_1203,N_769,N_674);
xnor U1204 (N_1204,N_67,N_508);
xnor U1205 (N_1205,N_721,N_109);
xor U1206 (N_1206,N_155,N_224);
or U1207 (N_1207,N_699,N_326);
and U1208 (N_1208,N_463,N_899);
nand U1209 (N_1209,N_943,N_14);
nand U1210 (N_1210,N_329,N_702);
nor U1211 (N_1211,N_916,N_584);
and U1212 (N_1212,N_165,N_729);
xnor U1213 (N_1213,N_433,N_945);
nand U1214 (N_1214,N_375,N_524);
and U1215 (N_1215,N_606,N_649);
nand U1216 (N_1216,N_6,N_569);
and U1217 (N_1217,N_850,N_416);
xnor U1218 (N_1218,N_3,N_156);
or U1219 (N_1219,N_708,N_36);
and U1220 (N_1220,N_81,N_989);
nor U1221 (N_1221,N_137,N_275);
or U1222 (N_1222,N_259,N_280);
xor U1223 (N_1223,N_504,N_86);
nor U1224 (N_1224,N_860,N_731);
nor U1225 (N_1225,N_833,N_717);
and U1226 (N_1226,N_868,N_69);
nor U1227 (N_1227,N_896,N_415);
or U1228 (N_1228,N_139,N_698);
nor U1229 (N_1229,N_971,N_509);
nand U1230 (N_1230,N_598,N_506);
nor U1231 (N_1231,N_160,N_580);
xor U1232 (N_1232,N_998,N_457);
and U1233 (N_1233,N_972,N_161);
xnor U1234 (N_1234,N_395,N_658);
nor U1235 (N_1235,N_237,N_443);
nand U1236 (N_1236,N_960,N_563);
and U1237 (N_1237,N_411,N_904);
nand U1238 (N_1238,N_11,N_522);
or U1239 (N_1239,N_311,N_982);
xor U1240 (N_1240,N_22,N_518);
xnor U1241 (N_1241,N_492,N_759);
and U1242 (N_1242,N_857,N_767);
nor U1243 (N_1243,N_201,N_550);
and U1244 (N_1244,N_24,N_936);
nor U1245 (N_1245,N_720,N_397);
nand U1246 (N_1246,N_858,N_824);
nand U1247 (N_1247,N_90,N_712);
or U1248 (N_1248,N_60,N_353);
nor U1249 (N_1249,N_478,N_531);
and U1250 (N_1250,N_409,N_843);
nand U1251 (N_1251,N_911,N_367);
xor U1252 (N_1252,N_609,N_272);
and U1253 (N_1253,N_645,N_597);
or U1254 (N_1254,N_714,N_194);
and U1255 (N_1255,N_253,N_219);
nor U1256 (N_1256,N_665,N_920);
nand U1257 (N_1257,N_730,N_54);
and U1258 (N_1258,N_847,N_439);
xnor U1259 (N_1259,N_419,N_921);
nand U1260 (N_1260,N_400,N_879);
and U1261 (N_1261,N_607,N_363);
nand U1262 (N_1262,N_264,N_451);
and U1263 (N_1263,N_745,N_991);
nand U1264 (N_1264,N_162,N_361);
nor U1265 (N_1265,N_484,N_581);
nand U1266 (N_1266,N_490,N_602);
and U1267 (N_1267,N_394,N_722);
nor U1268 (N_1268,N_876,N_931);
nand U1269 (N_1269,N_854,N_102);
nand U1270 (N_1270,N_127,N_208);
and U1271 (N_1271,N_785,N_350);
nand U1272 (N_1272,N_255,N_378);
nand U1273 (N_1273,N_952,N_227);
and U1274 (N_1274,N_917,N_875);
and U1275 (N_1275,N_650,N_377);
nor U1276 (N_1276,N_297,N_245);
nor U1277 (N_1277,N_959,N_976);
and U1278 (N_1278,N_690,N_837);
xor U1279 (N_1279,N_64,N_233);
xnor U1280 (N_1280,N_856,N_432);
or U1281 (N_1281,N_556,N_176);
nand U1282 (N_1282,N_198,N_436);
or U1283 (N_1283,N_407,N_962);
nor U1284 (N_1284,N_146,N_466);
or U1285 (N_1285,N_953,N_910);
and U1286 (N_1286,N_209,N_973);
nor U1287 (N_1287,N_274,N_796);
xor U1288 (N_1288,N_820,N_9);
nor U1289 (N_1289,N_749,N_98);
or U1290 (N_1290,N_851,N_7);
xnor U1291 (N_1291,N_339,N_96);
and U1292 (N_1292,N_29,N_85);
and U1293 (N_1293,N_398,N_314);
and U1294 (N_1294,N_453,N_343);
nand U1295 (N_1295,N_70,N_351);
or U1296 (N_1296,N_618,N_342);
and U1297 (N_1297,N_430,N_542);
xor U1298 (N_1298,N_497,N_304);
nand U1299 (N_1299,N_828,N_8);
and U1300 (N_1300,N_72,N_401);
nor U1301 (N_1301,N_354,N_599);
or U1302 (N_1302,N_184,N_42);
nand U1303 (N_1303,N_185,N_106);
nor U1304 (N_1304,N_949,N_907);
xnor U1305 (N_1305,N_628,N_751);
nand U1306 (N_1306,N_118,N_963);
or U1307 (N_1307,N_16,N_368);
or U1308 (N_1308,N_291,N_710);
and U1309 (N_1309,N_428,N_170);
nand U1310 (N_1310,N_742,N_360);
xnor U1311 (N_1311,N_489,N_586);
nor U1312 (N_1312,N_932,N_612);
nand U1313 (N_1313,N_295,N_819);
and U1314 (N_1314,N_152,N_472);
nand U1315 (N_1315,N_477,N_630);
and U1316 (N_1316,N_792,N_240);
xnor U1317 (N_1317,N_218,N_557);
nor U1318 (N_1318,N_142,N_279);
nor U1319 (N_1319,N_930,N_653);
or U1320 (N_1320,N_286,N_968);
nor U1321 (N_1321,N_260,N_399);
and U1322 (N_1322,N_883,N_386);
xnor U1323 (N_1323,N_10,N_600);
or U1324 (N_1324,N_768,N_840);
or U1325 (N_1325,N_431,N_983);
nand U1326 (N_1326,N_212,N_207);
and U1327 (N_1327,N_55,N_997);
xnor U1328 (N_1328,N_87,N_954);
nor U1329 (N_1329,N_315,N_76);
or U1330 (N_1330,N_623,N_446);
xnor U1331 (N_1331,N_328,N_789);
or U1332 (N_1332,N_680,N_678);
xnor U1333 (N_1333,N_412,N_124);
nor U1334 (N_1334,N_909,N_636);
or U1335 (N_1335,N_214,N_670);
and U1336 (N_1336,N_221,N_903);
and U1337 (N_1337,N_874,N_479);
xor U1338 (N_1338,N_302,N_765);
and U1339 (N_1339,N_45,N_780);
nor U1340 (N_1340,N_510,N_655);
nor U1341 (N_1341,N_452,N_448);
nand U1342 (N_1342,N_933,N_694);
xor U1343 (N_1343,N_133,N_462);
or U1344 (N_1344,N_758,N_115);
xnor U1345 (N_1345,N_706,N_540);
nor U1346 (N_1346,N_898,N_511);
or U1347 (N_1347,N_278,N_727);
xnor U1348 (N_1348,N_301,N_310);
nand U1349 (N_1349,N_229,N_327);
and U1350 (N_1350,N_44,N_781);
or U1351 (N_1351,N_39,N_273);
or U1352 (N_1352,N_613,N_585);
nand U1353 (N_1353,N_783,N_406);
xnor U1354 (N_1354,N_349,N_728);
and U1355 (N_1355,N_985,N_703);
xor U1356 (N_1356,N_795,N_49);
xor U1357 (N_1357,N_956,N_527);
and U1358 (N_1358,N_566,N_192);
or U1359 (N_1359,N_547,N_380);
and U1360 (N_1360,N_807,N_271);
nor U1361 (N_1361,N_391,N_487);
and U1362 (N_1362,N_317,N_644);
nor U1363 (N_1363,N_89,N_660);
nand U1364 (N_1364,N_225,N_558);
xnor U1365 (N_1365,N_817,N_873);
nor U1366 (N_1366,N_823,N_308);
or U1367 (N_1367,N_715,N_685);
xnor U1368 (N_1368,N_772,N_43);
nand U1369 (N_1369,N_151,N_732);
and U1370 (N_1370,N_359,N_705);
and U1371 (N_1371,N_454,N_158);
nand U1372 (N_1372,N_846,N_248);
nor U1373 (N_1373,N_12,N_541);
and U1374 (N_1374,N_56,N_589);
nand U1375 (N_1375,N_544,N_746);
nand U1376 (N_1376,N_141,N_535);
and U1377 (N_1377,N_736,N_794);
xnor U1378 (N_1378,N_957,N_919);
nor U1379 (N_1379,N_340,N_882);
xnor U1380 (N_1380,N_434,N_216);
or U1381 (N_1381,N_886,N_713);
or U1382 (N_1382,N_981,N_276);
xor U1383 (N_1383,N_889,N_373);
xor U1384 (N_1384,N_915,N_582);
and U1385 (N_1385,N_779,N_220);
xor U1386 (N_1386,N_429,N_107);
and U1387 (N_1387,N_704,N_839);
nor U1388 (N_1388,N_941,N_413);
and U1389 (N_1389,N_467,N_763);
nor U1390 (N_1390,N_895,N_652);
and U1391 (N_1391,N_682,N_773);
nand U1392 (N_1392,N_306,N_561);
and U1393 (N_1393,N_695,N_75);
and U1394 (N_1394,N_491,N_116);
nor U1395 (N_1395,N_605,N_800);
or U1396 (N_1396,N_424,N_461);
and U1397 (N_1397,N_565,N_664);
nor U1398 (N_1398,N_175,N_675);
or U1399 (N_1399,N_143,N_576);
and U1400 (N_1400,N_575,N_757);
and U1401 (N_1401,N_806,N_97);
nor U1402 (N_1402,N_226,N_554);
or U1403 (N_1403,N_523,N_994);
xnor U1404 (N_1404,N_427,N_438);
nor U1405 (N_1405,N_389,N_322);
or U1406 (N_1406,N_829,N_816);
nor U1407 (N_1407,N_123,N_444);
or U1408 (N_1408,N_935,N_169);
nand U1409 (N_1409,N_84,N_944);
or U1410 (N_1410,N_231,N_536);
or U1411 (N_1411,N_555,N_691);
nor U1412 (N_1412,N_374,N_995);
xnor U1413 (N_1413,N_63,N_324);
or U1414 (N_1414,N_735,N_129);
nand U1415 (N_1415,N_788,N_878);
nor U1416 (N_1416,N_393,N_626);
nand U1417 (N_1417,N_711,N_71);
nor U1418 (N_1418,N_420,N_551);
or U1419 (N_1419,N_894,N_844);
nor U1420 (N_1420,N_926,N_590);
and U1421 (N_1421,N_471,N_764);
or U1422 (N_1422,N_131,N_171);
nand U1423 (N_1423,N_756,N_534);
nor U1424 (N_1424,N_762,N_748);
xor U1425 (N_1425,N_638,N_709);
and U1426 (N_1426,N_753,N_908);
and U1427 (N_1427,N_942,N_629);
and U1428 (N_1428,N_132,N_182);
nand U1429 (N_1429,N_961,N_108);
or U1430 (N_1430,N_232,N_460);
nor U1431 (N_1431,N_241,N_578);
nor U1432 (N_1432,N_545,N_821);
and U1433 (N_1433,N_289,N_325);
xor U1434 (N_1434,N_738,N_388);
and U1435 (N_1435,N_120,N_747);
xor U1436 (N_1436,N_822,N_681);
xor U1437 (N_1437,N_164,N_929);
xor U1438 (N_1438,N_254,N_784);
nor U1439 (N_1439,N_539,N_552);
or U1440 (N_1440,N_425,N_965);
xnor U1441 (N_1441,N_707,N_103);
nor U1442 (N_1442,N_643,N_186);
or U1443 (N_1443,N_520,N_25);
nor U1444 (N_1444,N_980,N_572);
or U1445 (N_1445,N_285,N_159);
xnor U1446 (N_1446,N_330,N_383);
nor U1447 (N_1447,N_579,N_900);
nor U1448 (N_1448,N_913,N_163);
or U1449 (N_1449,N_988,N_99);
nand U1450 (N_1450,N_867,N_521);
and U1451 (N_1451,N_677,N_940);
nand U1452 (N_1452,N_502,N_811);
or U1453 (N_1453,N_239,N_266);
xor U1454 (N_1454,N_294,N_667);
and U1455 (N_1455,N_385,N_654);
and U1456 (N_1456,N_136,N_853);
and U1457 (N_1457,N_778,N_316);
xnor U1458 (N_1458,N_21,N_333);
nand U1459 (N_1459,N_5,N_470);
nand U1460 (N_1460,N_211,N_309);
xnor U1461 (N_1461,N_498,N_46);
nand U1462 (N_1462,N_740,N_77);
xor U1463 (N_1463,N_939,N_986);
xor U1464 (N_1464,N_546,N_320);
nor U1465 (N_1465,N_621,N_864);
nand U1466 (N_1466,N_902,N_41);
or U1467 (N_1467,N_15,N_519);
and U1468 (N_1468,N_47,N_918);
nor U1469 (N_1469,N_559,N_246);
xor U1470 (N_1470,N_684,N_28);
or U1471 (N_1471,N_303,N_336);
or U1472 (N_1472,N_37,N_725);
and U1473 (N_1473,N_200,N_447);
nand U1474 (N_1474,N_604,N_74);
xnor U1475 (N_1475,N_284,N_197);
or U1476 (N_1476,N_357,N_804);
or U1477 (N_1477,N_964,N_459);
nor U1478 (N_1478,N_61,N_923);
nor U1479 (N_1479,N_517,N_934);
nor U1480 (N_1480,N_26,N_135);
xnor U1481 (N_1481,N_754,N_692);
nor U1482 (N_1482,N_928,N_967);
xnor U1483 (N_1483,N_528,N_776);
xnor U1484 (N_1484,N_992,N_987);
nor U1485 (N_1485,N_217,N_500);
nand U1486 (N_1486,N_405,N_355);
and U1487 (N_1487,N_701,N_955);
or U1488 (N_1488,N_892,N_387);
or U1489 (N_1489,N_620,N_893);
or U1490 (N_1490,N_770,N_723);
xnor U1491 (N_1491,N_435,N_529);
nand U1492 (N_1492,N_786,N_937);
and U1493 (N_1493,N_126,N_696);
nor U1494 (N_1494,N_66,N_130);
xor U1495 (N_1495,N_242,N_592);
nand U1496 (N_1496,N_404,N_153);
xnor U1497 (N_1497,N_827,N_914);
nand U1498 (N_1498,N_396,N_810);
or U1499 (N_1499,N_863,N_95);
and U1500 (N_1500,N_689,N_757);
xnor U1501 (N_1501,N_659,N_221);
and U1502 (N_1502,N_475,N_947);
nand U1503 (N_1503,N_574,N_646);
nand U1504 (N_1504,N_981,N_374);
or U1505 (N_1505,N_167,N_953);
nor U1506 (N_1506,N_357,N_931);
and U1507 (N_1507,N_462,N_397);
xor U1508 (N_1508,N_622,N_866);
xor U1509 (N_1509,N_778,N_732);
nor U1510 (N_1510,N_188,N_783);
nor U1511 (N_1511,N_488,N_890);
xnor U1512 (N_1512,N_688,N_393);
and U1513 (N_1513,N_730,N_319);
nand U1514 (N_1514,N_780,N_578);
or U1515 (N_1515,N_397,N_349);
nand U1516 (N_1516,N_595,N_475);
or U1517 (N_1517,N_24,N_526);
nor U1518 (N_1518,N_666,N_10);
nand U1519 (N_1519,N_724,N_952);
or U1520 (N_1520,N_804,N_4);
or U1521 (N_1521,N_747,N_532);
nand U1522 (N_1522,N_689,N_669);
xor U1523 (N_1523,N_305,N_413);
and U1524 (N_1524,N_954,N_442);
nor U1525 (N_1525,N_16,N_985);
nand U1526 (N_1526,N_828,N_68);
nand U1527 (N_1527,N_276,N_624);
nor U1528 (N_1528,N_275,N_447);
xor U1529 (N_1529,N_929,N_329);
nand U1530 (N_1530,N_253,N_913);
nand U1531 (N_1531,N_139,N_457);
nor U1532 (N_1532,N_426,N_387);
and U1533 (N_1533,N_104,N_144);
xor U1534 (N_1534,N_176,N_715);
nor U1535 (N_1535,N_150,N_818);
xor U1536 (N_1536,N_275,N_251);
xnor U1537 (N_1537,N_153,N_449);
or U1538 (N_1538,N_334,N_847);
or U1539 (N_1539,N_97,N_252);
or U1540 (N_1540,N_662,N_480);
or U1541 (N_1541,N_329,N_909);
nor U1542 (N_1542,N_147,N_799);
and U1543 (N_1543,N_564,N_217);
or U1544 (N_1544,N_244,N_342);
or U1545 (N_1545,N_592,N_948);
xnor U1546 (N_1546,N_586,N_564);
xnor U1547 (N_1547,N_481,N_693);
nor U1548 (N_1548,N_121,N_805);
and U1549 (N_1549,N_22,N_528);
nor U1550 (N_1550,N_236,N_125);
or U1551 (N_1551,N_948,N_98);
xnor U1552 (N_1552,N_776,N_780);
nor U1553 (N_1553,N_215,N_908);
nor U1554 (N_1554,N_347,N_552);
xnor U1555 (N_1555,N_974,N_682);
or U1556 (N_1556,N_845,N_43);
xor U1557 (N_1557,N_514,N_556);
and U1558 (N_1558,N_442,N_259);
nor U1559 (N_1559,N_422,N_239);
nor U1560 (N_1560,N_848,N_777);
or U1561 (N_1561,N_204,N_981);
nand U1562 (N_1562,N_210,N_425);
and U1563 (N_1563,N_599,N_441);
and U1564 (N_1564,N_558,N_540);
xnor U1565 (N_1565,N_607,N_98);
xnor U1566 (N_1566,N_302,N_348);
nor U1567 (N_1567,N_769,N_836);
and U1568 (N_1568,N_955,N_866);
nand U1569 (N_1569,N_578,N_877);
nand U1570 (N_1570,N_475,N_31);
and U1571 (N_1571,N_51,N_292);
nor U1572 (N_1572,N_537,N_448);
nand U1573 (N_1573,N_828,N_608);
nand U1574 (N_1574,N_517,N_106);
xor U1575 (N_1575,N_309,N_894);
nand U1576 (N_1576,N_38,N_46);
nor U1577 (N_1577,N_465,N_621);
nor U1578 (N_1578,N_494,N_907);
or U1579 (N_1579,N_521,N_389);
and U1580 (N_1580,N_254,N_10);
and U1581 (N_1581,N_573,N_167);
xnor U1582 (N_1582,N_491,N_931);
and U1583 (N_1583,N_925,N_381);
and U1584 (N_1584,N_618,N_819);
and U1585 (N_1585,N_917,N_751);
xor U1586 (N_1586,N_787,N_673);
or U1587 (N_1587,N_32,N_708);
nand U1588 (N_1588,N_478,N_881);
nor U1589 (N_1589,N_801,N_278);
nand U1590 (N_1590,N_478,N_331);
nand U1591 (N_1591,N_187,N_152);
or U1592 (N_1592,N_935,N_747);
xnor U1593 (N_1593,N_257,N_227);
xnor U1594 (N_1594,N_939,N_106);
nor U1595 (N_1595,N_42,N_440);
nor U1596 (N_1596,N_553,N_395);
or U1597 (N_1597,N_311,N_679);
nor U1598 (N_1598,N_663,N_598);
and U1599 (N_1599,N_316,N_2);
or U1600 (N_1600,N_893,N_796);
and U1601 (N_1601,N_653,N_633);
or U1602 (N_1602,N_865,N_956);
or U1603 (N_1603,N_212,N_468);
xnor U1604 (N_1604,N_442,N_385);
xor U1605 (N_1605,N_95,N_729);
nor U1606 (N_1606,N_346,N_117);
nor U1607 (N_1607,N_989,N_640);
and U1608 (N_1608,N_448,N_739);
nor U1609 (N_1609,N_488,N_32);
nor U1610 (N_1610,N_448,N_125);
xnor U1611 (N_1611,N_535,N_823);
nand U1612 (N_1612,N_634,N_335);
nor U1613 (N_1613,N_879,N_622);
nand U1614 (N_1614,N_97,N_469);
xor U1615 (N_1615,N_16,N_166);
and U1616 (N_1616,N_875,N_426);
or U1617 (N_1617,N_212,N_195);
xnor U1618 (N_1618,N_824,N_848);
nor U1619 (N_1619,N_401,N_893);
or U1620 (N_1620,N_122,N_114);
or U1621 (N_1621,N_801,N_574);
or U1622 (N_1622,N_543,N_77);
nor U1623 (N_1623,N_845,N_101);
nand U1624 (N_1624,N_47,N_600);
nand U1625 (N_1625,N_258,N_526);
or U1626 (N_1626,N_261,N_27);
or U1627 (N_1627,N_488,N_981);
or U1628 (N_1628,N_288,N_597);
nand U1629 (N_1629,N_631,N_352);
and U1630 (N_1630,N_125,N_946);
or U1631 (N_1631,N_983,N_839);
xor U1632 (N_1632,N_6,N_275);
nor U1633 (N_1633,N_137,N_650);
nand U1634 (N_1634,N_553,N_679);
or U1635 (N_1635,N_912,N_711);
nand U1636 (N_1636,N_187,N_876);
xnor U1637 (N_1637,N_782,N_984);
xnor U1638 (N_1638,N_166,N_39);
nand U1639 (N_1639,N_113,N_859);
nand U1640 (N_1640,N_516,N_950);
nor U1641 (N_1641,N_9,N_907);
nor U1642 (N_1642,N_997,N_577);
or U1643 (N_1643,N_867,N_114);
and U1644 (N_1644,N_467,N_802);
nand U1645 (N_1645,N_274,N_226);
xor U1646 (N_1646,N_550,N_316);
or U1647 (N_1647,N_831,N_775);
nor U1648 (N_1648,N_452,N_141);
and U1649 (N_1649,N_194,N_454);
or U1650 (N_1650,N_205,N_918);
nor U1651 (N_1651,N_591,N_781);
nand U1652 (N_1652,N_268,N_199);
nand U1653 (N_1653,N_932,N_462);
nand U1654 (N_1654,N_207,N_669);
nor U1655 (N_1655,N_920,N_50);
xor U1656 (N_1656,N_780,N_657);
nand U1657 (N_1657,N_242,N_946);
nor U1658 (N_1658,N_775,N_852);
nor U1659 (N_1659,N_237,N_22);
nand U1660 (N_1660,N_298,N_29);
nor U1661 (N_1661,N_510,N_274);
or U1662 (N_1662,N_262,N_609);
xnor U1663 (N_1663,N_458,N_221);
and U1664 (N_1664,N_698,N_556);
or U1665 (N_1665,N_634,N_887);
or U1666 (N_1666,N_202,N_284);
xor U1667 (N_1667,N_552,N_344);
xnor U1668 (N_1668,N_960,N_925);
or U1669 (N_1669,N_282,N_9);
xor U1670 (N_1670,N_260,N_749);
or U1671 (N_1671,N_806,N_313);
nor U1672 (N_1672,N_340,N_127);
and U1673 (N_1673,N_857,N_450);
xor U1674 (N_1674,N_899,N_424);
and U1675 (N_1675,N_241,N_711);
xnor U1676 (N_1676,N_563,N_928);
xor U1677 (N_1677,N_501,N_480);
nand U1678 (N_1678,N_535,N_467);
and U1679 (N_1679,N_598,N_375);
and U1680 (N_1680,N_811,N_429);
and U1681 (N_1681,N_715,N_513);
nand U1682 (N_1682,N_970,N_538);
and U1683 (N_1683,N_115,N_733);
xor U1684 (N_1684,N_897,N_778);
or U1685 (N_1685,N_943,N_838);
or U1686 (N_1686,N_19,N_651);
xor U1687 (N_1687,N_855,N_808);
nor U1688 (N_1688,N_110,N_709);
nand U1689 (N_1689,N_694,N_396);
or U1690 (N_1690,N_765,N_32);
and U1691 (N_1691,N_813,N_484);
and U1692 (N_1692,N_586,N_792);
nor U1693 (N_1693,N_764,N_787);
nor U1694 (N_1694,N_905,N_475);
or U1695 (N_1695,N_111,N_942);
nand U1696 (N_1696,N_767,N_473);
or U1697 (N_1697,N_842,N_728);
xnor U1698 (N_1698,N_821,N_687);
or U1699 (N_1699,N_667,N_689);
nor U1700 (N_1700,N_220,N_130);
nand U1701 (N_1701,N_826,N_390);
or U1702 (N_1702,N_383,N_970);
or U1703 (N_1703,N_446,N_178);
or U1704 (N_1704,N_946,N_426);
and U1705 (N_1705,N_162,N_580);
xor U1706 (N_1706,N_430,N_596);
or U1707 (N_1707,N_221,N_128);
or U1708 (N_1708,N_351,N_139);
nor U1709 (N_1709,N_19,N_254);
and U1710 (N_1710,N_359,N_739);
and U1711 (N_1711,N_780,N_174);
nand U1712 (N_1712,N_24,N_996);
and U1713 (N_1713,N_232,N_93);
xnor U1714 (N_1714,N_506,N_794);
and U1715 (N_1715,N_515,N_790);
nand U1716 (N_1716,N_893,N_288);
or U1717 (N_1717,N_941,N_184);
nor U1718 (N_1718,N_239,N_182);
nand U1719 (N_1719,N_776,N_872);
nor U1720 (N_1720,N_694,N_492);
or U1721 (N_1721,N_703,N_113);
nor U1722 (N_1722,N_33,N_728);
and U1723 (N_1723,N_985,N_952);
xor U1724 (N_1724,N_941,N_970);
xnor U1725 (N_1725,N_941,N_479);
or U1726 (N_1726,N_990,N_775);
xor U1727 (N_1727,N_303,N_323);
or U1728 (N_1728,N_466,N_906);
xnor U1729 (N_1729,N_312,N_61);
or U1730 (N_1730,N_351,N_769);
and U1731 (N_1731,N_851,N_656);
and U1732 (N_1732,N_43,N_347);
xnor U1733 (N_1733,N_360,N_496);
and U1734 (N_1734,N_884,N_325);
or U1735 (N_1735,N_953,N_303);
xor U1736 (N_1736,N_624,N_554);
nor U1737 (N_1737,N_942,N_927);
nand U1738 (N_1738,N_808,N_899);
and U1739 (N_1739,N_606,N_741);
nand U1740 (N_1740,N_35,N_22);
or U1741 (N_1741,N_407,N_235);
and U1742 (N_1742,N_337,N_854);
nor U1743 (N_1743,N_762,N_192);
or U1744 (N_1744,N_799,N_904);
nand U1745 (N_1745,N_10,N_672);
nand U1746 (N_1746,N_628,N_41);
nand U1747 (N_1747,N_414,N_643);
and U1748 (N_1748,N_155,N_368);
or U1749 (N_1749,N_692,N_531);
or U1750 (N_1750,N_812,N_258);
and U1751 (N_1751,N_576,N_584);
nor U1752 (N_1752,N_803,N_127);
or U1753 (N_1753,N_970,N_593);
xnor U1754 (N_1754,N_371,N_193);
nor U1755 (N_1755,N_334,N_48);
xnor U1756 (N_1756,N_700,N_353);
and U1757 (N_1757,N_722,N_497);
nor U1758 (N_1758,N_189,N_725);
or U1759 (N_1759,N_406,N_16);
xor U1760 (N_1760,N_878,N_123);
xnor U1761 (N_1761,N_448,N_259);
nor U1762 (N_1762,N_565,N_769);
and U1763 (N_1763,N_416,N_70);
xnor U1764 (N_1764,N_505,N_29);
or U1765 (N_1765,N_819,N_717);
nand U1766 (N_1766,N_482,N_710);
or U1767 (N_1767,N_702,N_974);
or U1768 (N_1768,N_493,N_247);
or U1769 (N_1769,N_577,N_67);
and U1770 (N_1770,N_899,N_446);
or U1771 (N_1771,N_787,N_535);
nor U1772 (N_1772,N_145,N_170);
nand U1773 (N_1773,N_822,N_31);
and U1774 (N_1774,N_524,N_822);
or U1775 (N_1775,N_733,N_965);
and U1776 (N_1776,N_774,N_961);
nor U1777 (N_1777,N_315,N_222);
and U1778 (N_1778,N_88,N_312);
nor U1779 (N_1779,N_875,N_71);
xnor U1780 (N_1780,N_256,N_527);
xnor U1781 (N_1781,N_424,N_612);
nor U1782 (N_1782,N_460,N_450);
nand U1783 (N_1783,N_890,N_359);
and U1784 (N_1784,N_135,N_117);
nand U1785 (N_1785,N_238,N_897);
nand U1786 (N_1786,N_574,N_473);
and U1787 (N_1787,N_824,N_234);
and U1788 (N_1788,N_896,N_22);
or U1789 (N_1789,N_598,N_923);
and U1790 (N_1790,N_236,N_228);
nor U1791 (N_1791,N_170,N_451);
nor U1792 (N_1792,N_306,N_486);
nor U1793 (N_1793,N_652,N_368);
xor U1794 (N_1794,N_302,N_968);
nor U1795 (N_1795,N_158,N_260);
or U1796 (N_1796,N_747,N_616);
xor U1797 (N_1797,N_801,N_516);
nand U1798 (N_1798,N_533,N_557);
and U1799 (N_1799,N_934,N_632);
xnor U1800 (N_1800,N_1,N_833);
and U1801 (N_1801,N_81,N_672);
or U1802 (N_1802,N_549,N_321);
xnor U1803 (N_1803,N_344,N_486);
or U1804 (N_1804,N_692,N_567);
or U1805 (N_1805,N_834,N_420);
nor U1806 (N_1806,N_327,N_239);
nand U1807 (N_1807,N_411,N_979);
and U1808 (N_1808,N_32,N_615);
xnor U1809 (N_1809,N_589,N_837);
or U1810 (N_1810,N_384,N_57);
nand U1811 (N_1811,N_451,N_513);
nand U1812 (N_1812,N_491,N_608);
nand U1813 (N_1813,N_255,N_771);
nand U1814 (N_1814,N_985,N_198);
nand U1815 (N_1815,N_876,N_367);
and U1816 (N_1816,N_328,N_259);
or U1817 (N_1817,N_586,N_196);
xor U1818 (N_1818,N_982,N_592);
or U1819 (N_1819,N_169,N_580);
or U1820 (N_1820,N_670,N_105);
and U1821 (N_1821,N_167,N_930);
xnor U1822 (N_1822,N_927,N_299);
xnor U1823 (N_1823,N_432,N_765);
nor U1824 (N_1824,N_530,N_101);
nand U1825 (N_1825,N_401,N_435);
nand U1826 (N_1826,N_797,N_725);
and U1827 (N_1827,N_941,N_820);
xnor U1828 (N_1828,N_109,N_235);
and U1829 (N_1829,N_790,N_222);
and U1830 (N_1830,N_956,N_283);
nor U1831 (N_1831,N_860,N_170);
and U1832 (N_1832,N_332,N_212);
or U1833 (N_1833,N_859,N_472);
or U1834 (N_1834,N_415,N_411);
or U1835 (N_1835,N_265,N_71);
or U1836 (N_1836,N_932,N_747);
xnor U1837 (N_1837,N_611,N_466);
xnor U1838 (N_1838,N_90,N_666);
nand U1839 (N_1839,N_818,N_754);
and U1840 (N_1840,N_266,N_245);
or U1841 (N_1841,N_858,N_44);
nand U1842 (N_1842,N_620,N_488);
xor U1843 (N_1843,N_669,N_893);
nand U1844 (N_1844,N_654,N_991);
or U1845 (N_1845,N_523,N_800);
nor U1846 (N_1846,N_76,N_980);
nor U1847 (N_1847,N_47,N_679);
xnor U1848 (N_1848,N_644,N_508);
and U1849 (N_1849,N_961,N_606);
xnor U1850 (N_1850,N_432,N_866);
nand U1851 (N_1851,N_642,N_542);
nor U1852 (N_1852,N_516,N_114);
nor U1853 (N_1853,N_798,N_768);
or U1854 (N_1854,N_875,N_206);
and U1855 (N_1855,N_806,N_983);
nor U1856 (N_1856,N_637,N_948);
and U1857 (N_1857,N_565,N_577);
nand U1858 (N_1858,N_598,N_878);
and U1859 (N_1859,N_416,N_526);
xor U1860 (N_1860,N_267,N_258);
nor U1861 (N_1861,N_288,N_414);
nand U1862 (N_1862,N_235,N_795);
nor U1863 (N_1863,N_907,N_415);
and U1864 (N_1864,N_636,N_264);
or U1865 (N_1865,N_747,N_530);
or U1866 (N_1866,N_216,N_211);
xnor U1867 (N_1867,N_798,N_981);
and U1868 (N_1868,N_561,N_360);
xnor U1869 (N_1869,N_123,N_322);
nor U1870 (N_1870,N_500,N_870);
or U1871 (N_1871,N_58,N_374);
nor U1872 (N_1872,N_463,N_556);
xnor U1873 (N_1873,N_840,N_989);
nor U1874 (N_1874,N_106,N_854);
or U1875 (N_1875,N_773,N_496);
nor U1876 (N_1876,N_669,N_453);
xor U1877 (N_1877,N_957,N_709);
nand U1878 (N_1878,N_294,N_715);
nor U1879 (N_1879,N_610,N_62);
and U1880 (N_1880,N_99,N_459);
and U1881 (N_1881,N_434,N_320);
nor U1882 (N_1882,N_733,N_659);
xor U1883 (N_1883,N_857,N_415);
nand U1884 (N_1884,N_321,N_401);
xor U1885 (N_1885,N_948,N_104);
nand U1886 (N_1886,N_925,N_256);
nor U1887 (N_1887,N_223,N_388);
nor U1888 (N_1888,N_773,N_520);
xnor U1889 (N_1889,N_603,N_203);
or U1890 (N_1890,N_186,N_843);
or U1891 (N_1891,N_334,N_198);
or U1892 (N_1892,N_849,N_232);
or U1893 (N_1893,N_511,N_123);
nor U1894 (N_1894,N_509,N_871);
nor U1895 (N_1895,N_113,N_748);
or U1896 (N_1896,N_616,N_30);
or U1897 (N_1897,N_41,N_277);
nor U1898 (N_1898,N_36,N_389);
nor U1899 (N_1899,N_907,N_549);
and U1900 (N_1900,N_828,N_805);
nor U1901 (N_1901,N_110,N_460);
and U1902 (N_1902,N_666,N_441);
xnor U1903 (N_1903,N_910,N_975);
nand U1904 (N_1904,N_64,N_138);
xor U1905 (N_1905,N_974,N_40);
xnor U1906 (N_1906,N_456,N_592);
nand U1907 (N_1907,N_547,N_65);
nand U1908 (N_1908,N_295,N_650);
nand U1909 (N_1909,N_394,N_547);
or U1910 (N_1910,N_808,N_712);
or U1911 (N_1911,N_535,N_958);
nor U1912 (N_1912,N_248,N_450);
xnor U1913 (N_1913,N_803,N_197);
or U1914 (N_1914,N_820,N_899);
or U1915 (N_1915,N_64,N_136);
nor U1916 (N_1916,N_982,N_261);
and U1917 (N_1917,N_145,N_380);
nand U1918 (N_1918,N_390,N_560);
or U1919 (N_1919,N_857,N_852);
nor U1920 (N_1920,N_100,N_171);
xor U1921 (N_1921,N_755,N_545);
and U1922 (N_1922,N_849,N_393);
and U1923 (N_1923,N_532,N_158);
nor U1924 (N_1924,N_297,N_630);
nor U1925 (N_1925,N_422,N_187);
or U1926 (N_1926,N_35,N_412);
or U1927 (N_1927,N_573,N_447);
or U1928 (N_1928,N_556,N_7);
nand U1929 (N_1929,N_537,N_129);
or U1930 (N_1930,N_859,N_360);
nand U1931 (N_1931,N_765,N_453);
xnor U1932 (N_1932,N_622,N_163);
nor U1933 (N_1933,N_770,N_992);
or U1934 (N_1934,N_670,N_855);
xor U1935 (N_1935,N_404,N_179);
nand U1936 (N_1936,N_254,N_351);
or U1937 (N_1937,N_65,N_334);
xor U1938 (N_1938,N_284,N_211);
or U1939 (N_1939,N_693,N_301);
or U1940 (N_1940,N_462,N_32);
or U1941 (N_1941,N_786,N_454);
nor U1942 (N_1942,N_455,N_859);
xor U1943 (N_1943,N_453,N_220);
and U1944 (N_1944,N_859,N_391);
or U1945 (N_1945,N_261,N_16);
nand U1946 (N_1946,N_45,N_472);
nand U1947 (N_1947,N_124,N_816);
xor U1948 (N_1948,N_874,N_965);
xnor U1949 (N_1949,N_40,N_111);
nand U1950 (N_1950,N_901,N_584);
or U1951 (N_1951,N_422,N_913);
nand U1952 (N_1952,N_983,N_234);
or U1953 (N_1953,N_782,N_284);
nand U1954 (N_1954,N_168,N_54);
xor U1955 (N_1955,N_172,N_895);
xnor U1956 (N_1956,N_636,N_942);
xnor U1957 (N_1957,N_508,N_871);
or U1958 (N_1958,N_356,N_226);
and U1959 (N_1959,N_233,N_749);
nor U1960 (N_1960,N_956,N_505);
or U1961 (N_1961,N_20,N_526);
xor U1962 (N_1962,N_88,N_469);
nand U1963 (N_1963,N_943,N_276);
xnor U1964 (N_1964,N_427,N_75);
xnor U1965 (N_1965,N_212,N_632);
nand U1966 (N_1966,N_578,N_333);
nand U1967 (N_1967,N_210,N_417);
and U1968 (N_1968,N_521,N_453);
and U1969 (N_1969,N_326,N_367);
or U1970 (N_1970,N_788,N_45);
and U1971 (N_1971,N_436,N_143);
xnor U1972 (N_1972,N_263,N_572);
or U1973 (N_1973,N_699,N_761);
xnor U1974 (N_1974,N_353,N_238);
and U1975 (N_1975,N_621,N_44);
and U1976 (N_1976,N_164,N_810);
xnor U1977 (N_1977,N_3,N_48);
or U1978 (N_1978,N_961,N_306);
xnor U1979 (N_1979,N_703,N_368);
nor U1980 (N_1980,N_552,N_784);
nor U1981 (N_1981,N_114,N_829);
nand U1982 (N_1982,N_317,N_68);
nor U1983 (N_1983,N_818,N_586);
nand U1984 (N_1984,N_61,N_209);
or U1985 (N_1985,N_69,N_276);
nand U1986 (N_1986,N_666,N_39);
or U1987 (N_1987,N_908,N_54);
or U1988 (N_1988,N_380,N_529);
nor U1989 (N_1989,N_457,N_546);
nand U1990 (N_1990,N_148,N_456);
or U1991 (N_1991,N_311,N_230);
xor U1992 (N_1992,N_732,N_499);
nand U1993 (N_1993,N_277,N_469);
or U1994 (N_1994,N_550,N_481);
nand U1995 (N_1995,N_367,N_25);
nand U1996 (N_1996,N_66,N_309);
and U1997 (N_1997,N_865,N_731);
nor U1998 (N_1998,N_563,N_250);
and U1999 (N_1999,N_218,N_38);
nor U2000 (N_2000,N_1634,N_1477);
nand U2001 (N_2001,N_1445,N_1573);
and U2002 (N_2002,N_1959,N_1216);
and U2003 (N_2003,N_1533,N_1977);
and U2004 (N_2004,N_1479,N_1384);
xnor U2005 (N_2005,N_1065,N_1379);
nor U2006 (N_2006,N_1036,N_1425);
nor U2007 (N_2007,N_1488,N_1772);
or U2008 (N_2008,N_1773,N_1450);
and U2009 (N_2009,N_1745,N_1486);
nor U2010 (N_2010,N_1810,N_1242);
nor U2011 (N_2011,N_1124,N_1496);
nor U2012 (N_2012,N_1386,N_1354);
or U2013 (N_2013,N_1514,N_1034);
nand U2014 (N_2014,N_1805,N_1195);
or U2015 (N_2015,N_1865,N_1649);
xor U2016 (N_2016,N_1301,N_1013);
xor U2017 (N_2017,N_1393,N_1665);
xor U2018 (N_2018,N_1908,N_1516);
or U2019 (N_2019,N_1997,N_1989);
or U2020 (N_2020,N_1343,N_1397);
xnor U2021 (N_2021,N_1349,N_1846);
and U2022 (N_2022,N_1706,N_1220);
and U2023 (N_2023,N_1956,N_1342);
xor U2024 (N_2024,N_1261,N_1139);
or U2025 (N_2025,N_1537,N_1376);
nor U2026 (N_2026,N_1099,N_1899);
and U2027 (N_2027,N_1125,N_1587);
nand U2028 (N_2028,N_1686,N_1842);
or U2029 (N_2029,N_1315,N_1276);
xnor U2030 (N_2030,N_1272,N_1655);
and U2031 (N_2031,N_1159,N_1560);
nand U2032 (N_2032,N_1757,N_1682);
nand U2033 (N_2033,N_1027,N_1401);
or U2034 (N_2034,N_1302,N_1359);
and U2035 (N_2035,N_1375,N_1677);
nand U2036 (N_2036,N_1118,N_1346);
or U2037 (N_2037,N_1121,N_1919);
or U2038 (N_2038,N_1999,N_1565);
xnor U2039 (N_2039,N_1184,N_1699);
nor U2040 (N_2040,N_1607,N_1681);
and U2041 (N_2041,N_1453,N_1187);
and U2042 (N_2042,N_1843,N_1804);
nor U2043 (N_2043,N_1168,N_1991);
xnor U2044 (N_2044,N_1513,N_1471);
nor U2045 (N_2045,N_1597,N_1490);
or U2046 (N_2046,N_1392,N_1851);
or U2047 (N_2047,N_1247,N_1737);
and U2048 (N_2048,N_1645,N_1660);
and U2049 (N_2049,N_1658,N_1172);
xnor U2050 (N_2050,N_1844,N_1581);
nand U2051 (N_2051,N_1311,N_1023);
and U2052 (N_2052,N_1288,N_1189);
or U2053 (N_2053,N_1265,N_1830);
and U2054 (N_2054,N_1057,N_1404);
nor U2055 (N_2055,N_1632,N_1300);
and U2056 (N_2056,N_1669,N_1715);
nor U2057 (N_2057,N_1416,N_1148);
nand U2058 (N_2058,N_1402,N_1833);
and U2059 (N_2059,N_1019,N_1567);
xnor U2060 (N_2060,N_1792,N_1671);
or U2061 (N_2061,N_1492,N_1904);
nor U2062 (N_2062,N_1628,N_1569);
or U2063 (N_2063,N_1538,N_1047);
and U2064 (N_2064,N_1434,N_1941);
or U2065 (N_2065,N_1031,N_1781);
or U2066 (N_2066,N_1334,N_1519);
xor U2067 (N_2067,N_1618,N_1962);
nor U2068 (N_2068,N_1405,N_1633);
or U2069 (N_2069,N_1924,N_1720);
nor U2070 (N_2070,N_1561,N_1190);
or U2071 (N_2071,N_1612,N_1421);
or U2072 (N_2072,N_1077,N_1791);
and U2073 (N_2073,N_1394,N_1193);
nor U2074 (N_2074,N_1930,N_1713);
xor U2075 (N_2075,N_1039,N_1091);
xnor U2076 (N_2076,N_1884,N_1203);
nand U2077 (N_2077,N_1433,N_1818);
nor U2078 (N_2078,N_1233,N_1796);
nor U2079 (N_2079,N_1601,N_1724);
and U2080 (N_2080,N_1408,N_1528);
nand U2081 (N_2081,N_1028,N_1259);
and U2082 (N_2082,N_1022,N_1606);
nand U2083 (N_2083,N_1372,N_1071);
nor U2084 (N_2084,N_1964,N_1178);
nor U2085 (N_2085,N_1205,N_1897);
xor U2086 (N_2086,N_1279,N_1312);
nand U2087 (N_2087,N_1491,N_1695);
and U2088 (N_2088,N_1155,N_1223);
nor U2089 (N_2089,N_1106,N_1867);
xor U2090 (N_2090,N_1010,N_1616);
or U2091 (N_2091,N_1115,N_1679);
xnor U2092 (N_2092,N_1710,N_1024);
or U2093 (N_2093,N_1199,N_1317);
and U2094 (N_2094,N_1268,N_1389);
xor U2095 (N_2095,N_1794,N_1219);
and U2096 (N_2096,N_1950,N_1138);
or U2097 (N_2097,N_1263,N_1310);
or U2098 (N_2098,N_1497,N_1666);
nand U2099 (N_2099,N_1562,N_1870);
and U2100 (N_2100,N_1641,N_1369);
nor U2101 (N_2101,N_1826,N_1151);
xor U2102 (N_2102,N_1546,N_1202);
xor U2103 (N_2103,N_1274,N_1848);
xor U2104 (N_2104,N_1446,N_1002);
or U2105 (N_2105,N_1503,N_1008);
and U2106 (N_2106,N_1850,N_1938);
or U2107 (N_2107,N_1438,N_1994);
or U2108 (N_2108,N_1149,N_1755);
or U2109 (N_2109,N_1275,N_1378);
and U2110 (N_2110,N_1961,N_1456);
nand U2111 (N_2111,N_1322,N_1108);
and U2112 (N_2112,N_1722,N_1473);
or U2113 (N_2113,N_1933,N_1819);
nor U2114 (N_2114,N_1365,N_1893);
xor U2115 (N_2115,N_1165,N_1308);
xnor U2116 (N_2116,N_1700,N_1101);
nor U2117 (N_2117,N_1017,N_1449);
and U2118 (N_2118,N_1198,N_1014);
or U2119 (N_2119,N_1692,N_1776);
or U2120 (N_2120,N_1240,N_1140);
and U2121 (N_2121,N_1171,N_1335);
or U2122 (N_2122,N_1784,N_1079);
and U2123 (N_2123,N_1509,N_1415);
nor U2124 (N_2124,N_1257,N_1185);
nor U2125 (N_2125,N_1500,N_1923);
and U2126 (N_2126,N_1583,N_1617);
nor U2127 (N_2127,N_1370,N_1760);
and U2128 (N_2128,N_1179,N_1610);
nor U2129 (N_2129,N_1998,N_1926);
nand U2130 (N_2130,N_1042,N_1856);
and U2131 (N_2131,N_1901,N_1986);
or U2132 (N_2132,N_1245,N_1662);
xnor U2133 (N_2133,N_1622,N_1283);
xnor U2134 (N_2134,N_1642,N_1750);
or U2135 (N_2135,N_1968,N_1451);
xnor U2136 (N_2136,N_1454,N_1107);
or U2137 (N_2137,N_1802,N_1771);
or U2138 (N_2138,N_1277,N_1762);
or U2139 (N_2139,N_1066,N_1838);
nor U2140 (N_2140,N_1549,N_1466);
and U2141 (N_2141,N_1174,N_1798);
and U2142 (N_2142,N_1258,N_1507);
nor U2143 (N_2143,N_1452,N_1545);
xor U2144 (N_2144,N_1126,N_1196);
nand U2145 (N_2145,N_1134,N_1464);
xnor U2146 (N_2146,N_1508,N_1747);
xnor U2147 (N_2147,N_1297,N_1663);
or U2148 (N_2148,N_1738,N_1906);
and U2149 (N_2149,N_1939,N_1358);
xnor U2150 (N_2150,N_1996,N_1424);
or U2151 (N_2151,N_1889,N_1038);
nor U2152 (N_2152,N_1707,N_1879);
nand U2153 (N_2153,N_1221,N_1535);
or U2154 (N_2154,N_1868,N_1748);
or U2155 (N_2155,N_1542,N_1230);
and U2156 (N_2156,N_1602,N_1915);
or U2157 (N_2157,N_1820,N_1352);
xor U2158 (N_2158,N_1417,N_1578);
nand U2159 (N_2159,N_1011,N_1048);
nor U2160 (N_2160,N_1858,N_1058);
or U2161 (N_2161,N_1878,N_1419);
and U2162 (N_2162,N_1368,N_1319);
or U2163 (N_2163,N_1291,N_1307);
nor U2164 (N_2164,N_1357,N_1777);
and U2165 (N_2165,N_1068,N_1152);
nand U2166 (N_2166,N_1098,N_1815);
and U2167 (N_2167,N_1696,N_1429);
and U2168 (N_2168,N_1215,N_1303);
and U2169 (N_2169,N_1212,N_1990);
or U2170 (N_2170,N_1504,N_1056);
xor U2171 (N_2171,N_1391,N_1156);
and U2172 (N_2172,N_1269,N_1207);
xor U2173 (N_2173,N_1461,N_1954);
nor U2174 (N_2174,N_1166,N_1350);
nand U2175 (N_2175,N_1880,N_1410);
xor U2176 (N_2176,N_1521,N_1898);
nand U2177 (N_2177,N_1552,N_1059);
nand U2178 (N_2178,N_1611,N_1030);
and U2179 (N_2179,N_1494,N_1458);
nand U2180 (N_2180,N_1704,N_1966);
and U2181 (N_2181,N_1648,N_1361);
nand U2182 (N_2182,N_1520,N_1817);
or U2183 (N_2183,N_1387,N_1383);
nor U2184 (N_2184,N_1063,N_1570);
or U2185 (N_2185,N_1162,N_1110);
and U2186 (N_2186,N_1734,N_1592);
nand U2187 (N_2187,N_1217,N_1875);
or U2188 (N_2188,N_1931,N_1824);
or U2189 (N_2189,N_1102,N_1459);
nor U2190 (N_2190,N_1957,N_1921);
and U2191 (N_2191,N_1348,N_1321);
xor U2192 (N_2192,N_1061,N_1227);
nand U2193 (N_2193,N_1427,N_1123);
and U2194 (N_2194,N_1111,N_1351);
and U2195 (N_2195,N_1554,N_1866);
or U2196 (N_2196,N_1644,N_1736);
and U2197 (N_2197,N_1708,N_1169);
or U2198 (N_2198,N_1270,N_1176);
nor U2199 (N_2199,N_1328,N_1287);
nor U2200 (N_2200,N_1339,N_1412);
nand U2201 (N_2201,N_1631,N_1800);
and U2202 (N_2202,N_1114,N_1158);
nor U2203 (N_2203,N_1595,N_1982);
and U2204 (N_2204,N_1705,N_1891);
nor U2205 (N_2205,N_1385,N_1603);
nand U2206 (N_2206,N_1987,N_1442);
and U2207 (N_2207,N_1661,N_1907);
and U2208 (N_2208,N_1852,N_1356);
nand U2209 (N_2209,N_1313,N_1487);
or U2210 (N_2210,N_1070,N_1579);
nand U2211 (N_2211,N_1764,N_1399);
xor U2212 (N_2212,N_1044,N_1046);
xor U2213 (N_2213,N_1636,N_1180);
xor U2214 (N_2214,N_1330,N_1090);
nor U2215 (N_2215,N_1192,N_1337);
or U2216 (N_2216,N_1462,N_1130);
and U2217 (N_2217,N_1656,N_1652);
or U2218 (N_2218,N_1484,N_1555);
nor U2219 (N_2219,N_1382,N_1837);
and U2220 (N_2220,N_1709,N_1676);
xnor U2221 (N_2221,N_1741,N_1472);
xnor U2222 (N_2222,N_1120,N_1857);
or U2223 (N_2223,N_1053,N_1078);
nand U2224 (N_2224,N_1292,N_1512);
nor U2225 (N_2225,N_1096,N_1822);
nor U2226 (N_2226,N_1135,N_1971);
nand U2227 (N_2227,N_1702,N_1083);
nor U2228 (N_2228,N_1447,N_1087);
xor U2229 (N_2229,N_1763,N_1116);
nand U2230 (N_2230,N_1483,N_1113);
or U2231 (N_2231,N_1344,N_1129);
xor U2232 (N_2232,N_1910,N_1353);
nand U2233 (N_2233,N_1574,N_1886);
nor U2234 (N_2234,N_1638,N_1532);
nor U2235 (N_2235,N_1340,N_1949);
or U2236 (N_2236,N_1441,N_1685);
xnor U2237 (N_2237,N_1625,N_1626);
and U2238 (N_2238,N_1007,N_1530);
nor U2239 (N_2239,N_1244,N_1122);
nand U2240 (N_2240,N_1236,N_1790);
nand U2241 (N_2241,N_1905,N_1281);
nand U2242 (N_2242,N_1834,N_1770);
nor U2243 (N_2243,N_1539,N_1718);
xnor U2244 (N_2244,N_1237,N_1463);
nand U2245 (N_2245,N_1373,N_1694);
and U2246 (N_2246,N_1000,N_1803);
nor U2247 (N_2247,N_1672,N_1947);
or U2248 (N_2248,N_1067,N_1992);
or U2249 (N_2249,N_1320,N_1150);
and U2250 (N_2250,N_1041,N_1586);
or U2251 (N_2251,N_1828,N_1559);
xnor U2252 (N_2252,N_1160,N_1759);
nand U2253 (N_2253,N_1970,N_1728);
xor U2254 (N_2254,N_1614,N_1501);
nor U2255 (N_2255,N_1547,N_1224);
nand U2256 (N_2256,N_1254,N_1659);
or U2257 (N_2257,N_1100,N_1323);
xor U2258 (N_2258,N_1588,N_1188);
nor U2259 (N_2259,N_1204,N_1985);
xnor U2260 (N_2260,N_1782,N_1860);
nand U2261 (N_2261,N_1716,N_1495);
xnor U2262 (N_2262,N_1448,N_1756);
or U2263 (N_2263,N_1690,N_1765);
or U2264 (N_2264,N_1827,N_1945);
nor U2265 (N_2265,N_1871,N_1197);
or U2266 (N_2266,N_1609,N_1754);
xnor U2267 (N_2267,N_1831,N_1654);
nand U2268 (N_2268,N_1331,N_1437);
xor U2269 (N_2269,N_1476,N_1955);
nand U2270 (N_2270,N_1511,N_1670);
nor U2271 (N_2271,N_1325,N_1440);
and U2272 (N_2272,N_1299,N_1793);
xor U2273 (N_2273,N_1009,N_1208);
xnor U2274 (N_2274,N_1829,N_1814);
xnor U2275 (N_2275,N_1289,N_1714);
or U2276 (N_2276,N_1929,N_1304);
and U2277 (N_2277,N_1423,N_1841);
nor U2278 (N_2278,N_1914,N_1251);
xor U2279 (N_2279,N_1481,N_1235);
nor U2280 (N_2280,N_1089,N_1266);
nor U2281 (N_2281,N_1329,N_1572);
nor U2282 (N_2282,N_1246,N_1637);
xor U2283 (N_2283,N_1717,N_1175);
nand U2284 (N_2284,N_1684,N_1095);
and U2285 (N_2285,N_1548,N_1436);
or U2286 (N_2286,N_1482,N_1983);
nor U2287 (N_2287,N_1136,N_1876);
and U2288 (N_2288,N_1229,N_1069);
and U2289 (N_2289,N_1881,N_1214);
nand U2290 (N_2290,N_1531,N_1598);
nor U2291 (N_2291,N_1164,N_1580);
nand U2292 (N_2292,N_1502,N_1557);
nor U2293 (N_2293,N_1726,N_1267);
xor U2294 (N_2294,N_1604,N_1012);
or U2295 (N_2295,N_1953,N_1286);
and U2296 (N_2296,N_1167,N_1248);
nand U2297 (N_2297,N_1049,N_1576);
xor U2298 (N_2298,N_1062,N_1518);
xnor U2299 (N_2299,N_1799,N_1026);
nand U2300 (N_2300,N_1273,N_1021);
xnor U2301 (N_2301,N_1935,N_1558);
nand U2302 (N_2302,N_1485,N_1418);
or U2303 (N_2303,N_1522,N_1206);
nand U2304 (N_2304,N_1916,N_1944);
or U2305 (N_2305,N_1563,N_1786);
and U2306 (N_2306,N_1324,N_1527);
xnor U2307 (N_2307,N_1468,N_1157);
xnor U2308 (N_2308,N_1544,N_1743);
and U2309 (N_2309,N_1590,N_1211);
and U2310 (N_2310,N_1769,N_1627);
nand U2311 (N_2311,N_1499,N_1173);
nand U2312 (N_2312,N_1161,N_1298);
and U2313 (N_2313,N_1589,N_1816);
or U2314 (N_2314,N_1887,N_1144);
xnor U2315 (N_2315,N_1571,N_1925);
or U2316 (N_2316,N_1238,N_1836);
xor U2317 (N_2317,N_1988,N_1080);
nand U2318 (N_2318,N_1146,N_1367);
and U2319 (N_2319,N_1541,N_1639);
nand U2320 (N_2320,N_1568,N_1969);
nand U2321 (N_2321,N_1226,N_1624);
xnor U2322 (N_2322,N_1647,N_1920);
xor U2323 (N_2323,N_1885,N_1825);
nand U2324 (N_2324,N_1296,N_1594);
nand U2325 (N_2325,N_1054,N_1543);
nor U2326 (N_2326,N_1869,N_1154);
nor U2327 (N_2327,N_1742,N_1145);
nor U2328 (N_2328,N_1775,N_1979);
or U2329 (N_2329,N_1855,N_1043);
nand U2330 (N_2330,N_1788,N_1976);
xor U2331 (N_2331,N_1131,N_1643);
nor U2332 (N_2332,N_1882,N_1396);
nand U2333 (N_2333,N_1678,N_1225);
nor U2334 (N_2334,N_1582,N_1029);
or U2335 (N_2335,N_1282,N_1444);
nand U2336 (N_2336,N_1839,N_1474);
nor U2337 (N_2337,N_1951,N_1751);
xor U2338 (N_2338,N_1599,N_1094);
and U2339 (N_2339,N_1422,N_1657);
nor U2340 (N_2340,N_1064,N_1132);
and U2341 (N_2341,N_1536,N_1355);
xnor U2342 (N_2342,N_1697,N_1621);
or U2343 (N_2343,N_1290,N_1840);
and U2344 (N_2344,N_1097,N_1613);
xor U2345 (N_2345,N_1912,N_1293);
and U2346 (N_2346,N_1210,N_1761);
or U2347 (N_2347,N_1128,N_1877);
xnor U2348 (N_2348,N_1060,N_1721);
xnor U2349 (N_2349,N_1664,N_1963);
or U2350 (N_2350,N_1918,N_1050);
or U2351 (N_2351,N_1902,N_1200);
nand U2352 (N_2352,N_1163,N_1779);
and U2353 (N_2353,N_1687,N_1927);
nand U2354 (N_2354,N_1584,N_1711);
xnor U2355 (N_2355,N_1911,N_1316);
nor U2356 (N_2356,N_1086,N_1406);
nor U2357 (N_2357,N_1585,N_1255);
nand U2358 (N_2358,N_1515,N_1455);
nor U2359 (N_2359,N_1278,N_1993);
and U2360 (N_2360,N_1318,N_1109);
xor U2361 (N_2361,N_1018,N_1377);
and U2362 (N_2362,N_1363,N_1081);
nor U2363 (N_2363,N_1228,N_1457);
nand U2364 (N_2364,N_1730,N_1698);
or U2365 (N_2365,N_1766,N_1435);
nor U2366 (N_2366,N_1250,N_1942);
and U2367 (N_2367,N_1032,N_1693);
xor U2368 (N_2368,N_1306,N_1774);
and U2369 (N_2369,N_1127,N_1593);
and U2370 (N_2370,N_1142,N_1407);
or U2371 (N_2371,N_1896,N_1088);
or U2372 (N_2372,N_1467,N_1073);
xnor U2373 (N_2373,N_1524,N_1629);
nand U2374 (N_2374,N_1783,N_1845);
and U2375 (N_2375,N_1525,N_1605);
and U2376 (N_2376,N_1103,N_1523);
nor U2377 (N_2377,N_1443,N_1691);
nand U2378 (N_2378,N_1006,N_1366);
and U2379 (N_2379,N_1498,N_1295);
nor U2380 (N_2380,N_1428,N_1020);
or U2381 (N_2381,N_1689,N_1640);
nand U2382 (N_2382,N_1821,N_1170);
nand U2383 (N_2383,N_1808,N_1092);
nor U2384 (N_2384,N_1338,N_1853);
or U2385 (N_2385,N_1739,N_1209);
xnor U2386 (N_2386,N_1811,N_1758);
nand U2387 (N_2387,N_1493,N_1909);
or U2388 (N_2388,N_1575,N_1940);
xnor U2389 (N_2389,N_1465,N_1016);
and U2390 (N_2390,N_1510,N_1650);
nand U2391 (N_2391,N_1892,N_1615);
or U2392 (N_2392,N_1795,N_1787);
and U2393 (N_2393,N_1608,N_1936);
nand U2394 (N_2394,N_1812,N_1972);
or U2395 (N_2395,N_1731,N_1668);
and U2396 (N_2396,N_1540,N_1327);
xor U2397 (N_2397,N_1137,N_1015);
and U2398 (N_2398,N_1967,N_1778);
or U2399 (N_2399,N_1823,N_1439);
and U2400 (N_2400,N_1785,N_1117);
and U2401 (N_2401,N_1556,N_1347);
nor U2402 (N_2402,N_1403,N_1566);
xnor U2403 (N_2403,N_1958,N_1517);
nor U2404 (N_2404,N_1431,N_1703);
nand U2405 (N_2405,N_1390,N_1591);
nor U2406 (N_2406,N_1832,N_1271);
or U2407 (N_2407,N_1232,N_1733);
nand U2408 (N_2408,N_1943,N_1314);
xor U2409 (N_2409,N_1143,N_1928);
or U2410 (N_2410,N_1995,N_1577);
nor U2411 (N_2411,N_1280,N_1674);
nand U2412 (N_2412,N_1045,N_1600);
xor U2413 (N_2413,N_1284,N_1854);
nor U2414 (N_2414,N_1505,N_1980);
xor U2415 (N_2415,N_1051,N_1432);
nor U2416 (N_2416,N_1529,N_1890);
and U2417 (N_2417,N_1932,N_1680);
nor U2418 (N_2418,N_1234,N_1336);
or U2419 (N_2419,N_1182,N_1974);
and U2420 (N_2420,N_1035,N_1388);
xnor U2421 (N_2421,N_1201,N_1667);
nor U2422 (N_2422,N_1740,N_1241);
nand U2423 (N_2423,N_1469,N_1813);
or U2424 (N_2424,N_1735,N_1861);
or U2425 (N_2425,N_1478,N_1470);
nor U2426 (N_2426,N_1768,N_1859);
and U2427 (N_2427,N_1005,N_1332);
xnor U2428 (N_2428,N_1719,N_1104);
nand U2429 (N_2429,N_1364,N_1243);
nand U2430 (N_2430,N_1239,N_1948);
xor U2431 (N_2431,N_1285,N_1978);
xor U2432 (N_2432,N_1973,N_1112);
nand U2433 (N_2433,N_1147,N_1849);
xor U2434 (N_2434,N_1630,N_1635);
xor U2435 (N_2435,N_1746,N_1862);
xor U2436 (N_2436,N_1653,N_1398);
and U2437 (N_2437,N_1218,N_1025);
and U2438 (N_2438,N_1534,N_1732);
or U2439 (N_2439,N_1801,N_1186);
nor U2440 (N_2440,N_1305,N_1231);
and U2441 (N_2441,N_1550,N_1683);
nor U2442 (N_2442,N_1075,N_1260);
nor U2443 (N_2443,N_1752,N_1371);
and U2444 (N_2444,N_1133,N_1252);
nand U2445 (N_2445,N_1253,N_1727);
nand U2446 (N_2446,N_1333,N_1430);
or U2447 (N_2447,N_1725,N_1141);
nor U2448 (N_2448,N_1620,N_1913);
or U2449 (N_2449,N_1809,N_1222);
xor U2450 (N_2450,N_1003,N_1093);
or U2451 (N_2451,N_1183,N_1119);
and U2452 (N_2452,N_1551,N_1895);
nand U2453 (N_2453,N_1675,N_1863);
nand U2454 (N_2454,N_1723,N_1326);
and U2455 (N_2455,N_1374,N_1177);
xor U2456 (N_2456,N_1806,N_1213);
xnor U2457 (N_2457,N_1181,N_1341);
and U2458 (N_2458,N_1489,N_1360);
and U2459 (N_2459,N_1780,N_1981);
and U2460 (N_2460,N_1744,N_1040);
xor U2461 (N_2461,N_1380,N_1729);
or U2462 (N_2462,N_1872,N_1767);
and U2463 (N_2463,N_1409,N_1249);
or U2464 (N_2464,N_1847,N_1712);
nand U2465 (N_2465,N_1984,N_1673);
xor U2466 (N_2466,N_1960,N_1413);
xor U2467 (N_2467,N_1052,N_1835);
nand U2468 (N_2468,N_1153,N_1864);
nand U2469 (N_2469,N_1426,N_1701);
nand U2470 (N_2470,N_1874,N_1414);
nand U2471 (N_2471,N_1037,N_1894);
and U2472 (N_2472,N_1475,N_1688);
and U2473 (N_2473,N_1420,N_1965);
nand U2474 (N_2474,N_1460,N_1309);
nor U2475 (N_2475,N_1345,N_1553);
xnor U2476 (N_2476,N_1072,N_1082);
nor U2477 (N_2477,N_1749,N_1362);
xor U2478 (N_2478,N_1807,N_1395);
or U2479 (N_2479,N_1264,N_1411);
and U2480 (N_2480,N_1975,N_1033);
or U2481 (N_2481,N_1623,N_1055);
xor U2482 (N_2482,N_1085,N_1526);
or U2483 (N_2483,N_1917,N_1262);
xnor U2484 (N_2484,N_1789,N_1564);
and U2485 (N_2485,N_1903,N_1646);
nor U2486 (N_2486,N_1952,N_1105);
xor U2487 (N_2487,N_1194,N_1004);
nor U2488 (N_2488,N_1922,N_1596);
nand U2489 (N_2489,N_1753,N_1797);
xor U2490 (N_2490,N_1294,N_1900);
nand U2491 (N_2491,N_1480,N_1883);
xor U2492 (N_2492,N_1506,N_1651);
and U2493 (N_2493,N_1946,N_1934);
nand U2494 (N_2494,N_1619,N_1256);
and U2495 (N_2495,N_1400,N_1888);
or U2496 (N_2496,N_1001,N_1074);
nand U2497 (N_2497,N_1381,N_1076);
xnor U2498 (N_2498,N_1937,N_1873);
nor U2499 (N_2499,N_1084,N_1191);
or U2500 (N_2500,N_1416,N_1672);
nor U2501 (N_2501,N_1573,N_1811);
nor U2502 (N_2502,N_1515,N_1256);
xor U2503 (N_2503,N_1790,N_1648);
nor U2504 (N_2504,N_1614,N_1480);
and U2505 (N_2505,N_1296,N_1649);
xnor U2506 (N_2506,N_1925,N_1262);
nor U2507 (N_2507,N_1483,N_1086);
or U2508 (N_2508,N_1997,N_1583);
nor U2509 (N_2509,N_1312,N_1338);
nand U2510 (N_2510,N_1054,N_1260);
nand U2511 (N_2511,N_1603,N_1241);
xor U2512 (N_2512,N_1598,N_1914);
xnor U2513 (N_2513,N_1434,N_1665);
xor U2514 (N_2514,N_1506,N_1110);
or U2515 (N_2515,N_1514,N_1168);
xnor U2516 (N_2516,N_1502,N_1909);
xnor U2517 (N_2517,N_1123,N_1709);
or U2518 (N_2518,N_1812,N_1527);
xnor U2519 (N_2519,N_1414,N_1385);
nand U2520 (N_2520,N_1702,N_1180);
and U2521 (N_2521,N_1423,N_1188);
nand U2522 (N_2522,N_1401,N_1687);
nand U2523 (N_2523,N_1723,N_1775);
and U2524 (N_2524,N_1828,N_1291);
nor U2525 (N_2525,N_1669,N_1685);
and U2526 (N_2526,N_1854,N_1852);
nor U2527 (N_2527,N_1686,N_1733);
and U2528 (N_2528,N_1595,N_1917);
xnor U2529 (N_2529,N_1068,N_1505);
nand U2530 (N_2530,N_1845,N_1846);
or U2531 (N_2531,N_1490,N_1752);
and U2532 (N_2532,N_1507,N_1756);
or U2533 (N_2533,N_1816,N_1292);
nor U2534 (N_2534,N_1306,N_1113);
and U2535 (N_2535,N_1316,N_1817);
or U2536 (N_2536,N_1644,N_1947);
xnor U2537 (N_2537,N_1996,N_1312);
or U2538 (N_2538,N_1644,N_1322);
nor U2539 (N_2539,N_1725,N_1594);
nor U2540 (N_2540,N_1527,N_1909);
nor U2541 (N_2541,N_1875,N_1323);
nand U2542 (N_2542,N_1478,N_1491);
or U2543 (N_2543,N_1493,N_1268);
nor U2544 (N_2544,N_1995,N_1956);
nand U2545 (N_2545,N_1948,N_1072);
xnor U2546 (N_2546,N_1943,N_1970);
nand U2547 (N_2547,N_1364,N_1680);
nor U2548 (N_2548,N_1198,N_1312);
nor U2549 (N_2549,N_1160,N_1903);
and U2550 (N_2550,N_1500,N_1562);
nand U2551 (N_2551,N_1490,N_1126);
and U2552 (N_2552,N_1658,N_1750);
or U2553 (N_2553,N_1765,N_1860);
or U2554 (N_2554,N_1013,N_1587);
nand U2555 (N_2555,N_1338,N_1078);
nor U2556 (N_2556,N_1820,N_1060);
nor U2557 (N_2557,N_1190,N_1423);
xor U2558 (N_2558,N_1022,N_1216);
xnor U2559 (N_2559,N_1538,N_1629);
or U2560 (N_2560,N_1506,N_1105);
nand U2561 (N_2561,N_1176,N_1674);
or U2562 (N_2562,N_1247,N_1119);
xor U2563 (N_2563,N_1668,N_1326);
and U2564 (N_2564,N_1850,N_1776);
and U2565 (N_2565,N_1359,N_1923);
and U2566 (N_2566,N_1104,N_1695);
nand U2567 (N_2567,N_1016,N_1848);
nand U2568 (N_2568,N_1175,N_1906);
nand U2569 (N_2569,N_1247,N_1812);
nand U2570 (N_2570,N_1705,N_1959);
xnor U2571 (N_2571,N_1016,N_1811);
and U2572 (N_2572,N_1735,N_1387);
nor U2573 (N_2573,N_1026,N_1704);
xor U2574 (N_2574,N_1432,N_1977);
or U2575 (N_2575,N_1757,N_1457);
nor U2576 (N_2576,N_1630,N_1912);
xor U2577 (N_2577,N_1160,N_1956);
or U2578 (N_2578,N_1963,N_1856);
xnor U2579 (N_2579,N_1117,N_1822);
or U2580 (N_2580,N_1656,N_1907);
or U2581 (N_2581,N_1252,N_1625);
xor U2582 (N_2582,N_1607,N_1062);
xnor U2583 (N_2583,N_1616,N_1189);
or U2584 (N_2584,N_1875,N_1559);
and U2585 (N_2585,N_1517,N_1589);
nand U2586 (N_2586,N_1984,N_1817);
or U2587 (N_2587,N_1691,N_1224);
and U2588 (N_2588,N_1957,N_1809);
xor U2589 (N_2589,N_1407,N_1478);
and U2590 (N_2590,N_1424,N_1429);
xnor U2591 (N_2591,N_1501,N_1472);
nand U2592 (N_2592,N_1990,N_1647);
and U2593 (N_2593,N_1751,N_1796);
and U2594 (N_2594,N_1815,N_1729);
nand U2595 (N_2595,N_1513,N_1855);
nor U2596 (N_2596,N_1805,N_1700);
or U2597 (N_2597,N_1907,N_1767);
and U2598 (N_2598,N_1922,N_1144);
and U2599 (N_2599,N_1315,N_1559);
nand U2600 (N_2600,N_1702,N_1402);
nand U2601 (N_2601,N_1187,N_1244);
or U2602 (N_2602,N_1040,N_1625);
nand U2603 (N_2603,N_1504,N_1902);
or U2604 (N_2604,N_1274,N_1033);
nand U2605 (N_2605,N_1912,N_1677);
nand U2606 (N_2606,N_1485,N_1667);
or U2607 (N_2607,N_1613,N_1383);
nor U2608 (N_2608,N_1811,N_1254);
and U2609 (N_2609,N_1692,N_1805);
or U2610 (N_2610,N_1630,N_1079);
xnor U2611 (N_2611,N_1098,N_1770);
xnor U2612 (N_2612,N_1715,N_1082);
or U2613 (N_2613,N_1828,N_1227);
nor U2614 (N_2614,N_1371,N_1360);
nor U2615 (N_2615,N_1813,N_1316);
or U2616 (N_2616,N_1037,N_1593);
nor U2617 (N_2617,N_1248,N_1490);
nand U2618 (N_2618,N_1216,N_1797);
nand U2619 (N_2619,N_1182,N_1125);
or U2620 (N_2620,N_1505,N_1327);
or U2621 (N_2621,N_1595,N_1518);
xor U2622 (N_2622,N_1512,N_1732);
xnor U2623 (N_2623,N_1013,N_1200);
or U2624 (N_2624,N_1207,N_1300);
and U2625 (N_2625,N_1935,N_1475);
nor U2626 (N_2626,N_1919,N_1140);
xnor U2627 (N_2627,N_1973,N_1482);
or U2628 (N_2628,N_1215,N_1262);
nand U2629 (N_2629,N_1369,N_1424);
and U2630 (N_2630,N_1817,N_1273);
and U2631 (N_2631,N_1476,N_1202);
nor U2632 (N_2632,N_1277,N_1419);
and U2633 (N_2633,N_1126,N_1224);
or U2634 (N_2634,N_1610,N_1396);
nand U2635 (N_2635,N_1400,N_1044);
nor U2636 (N_2636,N_1701,N_1289);
xor U2637 (N_2637,N_1831,N_1102);
or U2638 (N_2638,N_1823,N_1679);
xnor U2639 (N_2639,N_1118,N_1324);
and U2640 (N_2640,N_1136,N_1517);
nand U2641 (N_2641,N_1321,N_1248);
nor U2642 (N_2642,N_1052,N_1119);
nor U2643 (N_2643,N_1350,N_1670);
or U2644 (N_2644,N_1324,N_1883);
xor U2645 (N_2645,N_1676,N_1752);
and U2646 (N_2646,N_1738,N_1001);
nor U2647 (N_2647,N_1107,N_1542);
or U2648 (N_2648,N_1417,N_1608);
and U2649 (N_2649,N_1893,N_1654);
nor U2650 (N_2650,N_1859,N_1012);
nand U2651 (N_2651,N_1972,N_1311);
nand U2652 (N_2652,N_1713,N_1846);
or U2653 (N_2653,N_1072,N_1981);
xnor U2654 (N_2654,N_1363,N_1369);
nand U2655 (N_2655,N_1935,N_1567);
and U2656 (N_2656,N_1328,N_1197);
nor U2657 (N_2657,N_1510,N_1308);
nor U2658 (N_2658,N_1845,N_1579);
nor U2659 (N_2659,N_1733,N_1730);
xor U2660 (N_2660,N_1805,N_1000);
nand U2661 (N_2661,N_1980,N_1163);
nor U2662 (N_2662,N_1704,N_1947);
nor U2663 (N_2663,N_1797,N_1881);
nor U2664 (N_2664,N_1509,N_1744);
or U2665 (N_2665,N_1347,N_1580);
nor U2666 (N_2666,N_1230,N_1443);
and U2667 (N_2667,N_1656,N_1698);
nor U2668 (N_2668,N_1001,N_1000);
or U2669 (N_2669,N_1087,N_1914);
nor U2670 (N_2670,N_1546,N_1704);
and U2671 (N_2671,N_1989,N_1166);
xor U2672 (N_2672,N_1480,N_1967);
nor U2673 (N_2673,N_1877,N_1850);
xnor U2674 (N_2674,N_1680,N_1575);
nand U2675 (N_2675,N_1904,N_1972);
nand U2676 (N_2676,N_1659,N_1399);
xnor U2677 (N_2677,N_1397,N_1098);
nor U2678 (N_2678,N_1721,N_1615);
xor U2679 (N_2679,N_1095,N_1675);
xnor U2680 (N_2680,N_1207,N_1329);
xnor U2681 (N_2681,N_1001,N_1230);
nand U2682 (N_2682,N_1571,N_1974);
xnor U2683 (N_2683,N_1948,N_1167);
nand U2684 (N_2684,N_1720,N_1955);
nand U2685 (N_2685,N_1156,N_1324);
nor U2686 (N_2686,N_1627,N_1257);
or U2687 (N_2687,N_1682,N_1290);
xor U2688 (N_2688,N_1095,N_1740);
nor U2689 (N_2689,N_1699,N_1790);
and U2690 (N_2690,N_1898,N_1138);
nor U2691 (N_2691,N_1787,N_1604);
xor U2692 (N_2692,N_1750,N_1125);
nand U2693 (N_2693,N_1242,N_1990);
and U2694 (N_2694,N_1272,N_1232);
nor U2695 (N_2695,N_1746,N_1502);
nor U2696 (N_2696,N_1358,N_1027);
xor U2697 (N_2697,N_1039,N_1095);
xnor U2698 (N_2698,N_1627,N_1574);
nand U2699 (N_2699,N_1110,N_1167);
xnor U2700 (N_2700,N_1384,N_1306);
xnor U2701 (N_2701,N_1381,N_1723);
or U2702 (N_2702,N_1573,N_1851);
and U2703 (N_2703,N_1077,N_1218);
and U2704 (N_2704,N_1685,N_1010);
xnor U2705 (N_2705,N_1688,N_1023);
nor U2706 (N_2706,N_1350,N_1414);
xor U2707 (N_2707,N_1666,N_1185);
or U2708 (N_2708,N_1629,N_1392);
xnor U2709 (N_2709,N_1113,N_1819);
nand U2710 (N_2710,N_1277,N_1534);
nor U2711 (N_2711,N_1780,N_1673);
or U2712 (N_2712,N_1908,N_1901);
nand U2713 (N_2713,N_1875,N_1908);
or U2714 (N_2714,N_1403,N_1841);
and U2715 (N_2715,N_1349,N_1107);
and U2716 (N_2716,N_1425,N_1927);
or U2717 (N_2717,N_1285,N_1228);
nor U2718 (N_2718,N_1978,N_1043);
nor U2719 (N_2719,N_1299,N_1667);
nand U2720 (N_2720,N_1080,N_1894);
nand U2721 (N_2721,N_1661,N_1107);
or U2722 (N_2722,N_1423,N_1831);
xnor U2723 (N_2723,N_1527,N_1130);
and U2724 (N_2724,N_1528,N_1350);
nor U2725 (N_2725,N_1772,N_1133);
or U2726 (N_2726,N_1444,N_1866);
or U2727 (N_2727,N_1377,N_1759);
nand U2728 (N_2728,N_1193,N_1534);
nor U2729 (N_2729,N_1078,N_1253);
and U2730 (N_2730,N_1999,N_1968);
nand U2731 (N_2731,N_1870,N_1194);
nor U2732 (N_2732,N_1287,N_1251);
nor U2733 (N_2733,N_1713,N_1330);
nand U2734 (N_2734,N_1362,N_1854);
nand U2735 (N_2735,N_1542,N_1183);
nor U2736 (N_2736,N_1092,N_1629);
nor U2737 (N_2737,N_1947,N_1626);
xnor U2738 (N_2738,N_1333,N_1670);
xnor U2739 (N_2739,N_1411,N_1260);
or U2740 (N_2740,N_1904,N_1074);
xnor U2741 (N_2741,N_1141,N_1390);
or U2742 (N_2742,N_1053,N_1109);
nand U2743 (N_2743,N_1878,N_1443);
nand U2744 (N_2744,N_1973,N_1116);
nand U2745 (N_2745,N_1757,N_1873);
or U2746 (N_2746,N_1512,N_1063);
xnor U2747 (N_2747,N_1201,N_1643);
and U2748 (N_2748,N_1177,N_1230);
nand U2749 (N_2749,N_1815,N_1478);
nor U2750 (N_2750,N_1776,N_1538);
nor U2751 (N_2751,N_1440,N_1228);
xor U2752 (N_2752,N_1227,N_1160);
nor U2753 (N_2753,N_1376,N_1669);
and U2754 (N_2754,N_1141,N_1157);
and U2755 (N_2755,N_1611,N_1125);
or U2756 (N_2756,N_1936,N_1077);
or U2757 (N_2757,N_1426,N_1430);
nand U2758 (N_2758,N_1374,N_1557);
nand U2759 (N_2759,N_1001,N_1096);
nor U2760 (N_2760,N_1807,N_1738);
or U2761 (N_2761,N_1170,N_1894);
nand U2762 (N_2762,N_1881,N_1200);
nor U2763 (N_2763,N_1134,N_1884);
xnor U2764 (N_2764,N_1016,N_1266);
nor U2765 (N_2765,N_1109,N_1240);
nor U2766 (N_2766,N_1436,N_1901);
nand U2767 (N_2767,N_1241,N_1630);
and U2768 (N_2768,N_1905,N_1693);
xor U2769 (N_2769,N_1338,N_1329);
or U2770 (N_2770,N_1051,N_1726);
or U2771 (N_2771,N_1135,N_1572);
nor U2772 (N_2772,N_1562,N_1413);
nor U2773 (N_2773,N_1180,N_1820);
and U2774 (N_2774,N_1660,N_1701);
or U2775 (N_2775,N_1795,N_1894);
nand U2776 (N_2776,N_1208,N_1340);
or U2777 (N_2777,N_1672,N_1365);
and U2778 (N_2778,N_1681,N_1091);
nor U2779 (N_2779,N_1457,N_1659);
or U2780 (N_2780,N_1405,N_1419);
nand U2781 (N_2781,N_1733,N_1864);
nand U2782 (N_2782,N_1142,N_1806);
nor U2783 (N_2783,N_1707,N_1765);
nand U2784 (N_2784,N_1007,N_1843);
xnor U2785 (N_2785,N_1229,N_1253);
nand U2786 (N_2786,N_1914,N_1680);
nand U2787 (N_2787,N_1177,N_1294);
nor U2788 (N_2788,N_1919,N_1155);
nor U2789 (N_2789,N_1232,N_1438);
nand U2790 (N_2790,N_1084,N_1044);
xor U2791 (N_2791,N_1845,N_1036);
and U2792 (N_2792,N_1873,N_1616);
nand U2793 (N_2793,N_1057,N_1396);
and U2794 (N_2794,N_1963,N_1512);
and U2795 (N_2795,N_1709,N_1671);
nand U2796 (N_2796,N_1147,N_1153);
xor U2797 (N_2797,N_1292,N_1470);
xnor U2798 (N_2798,N_1486,N_1589);
nor U2799 (N_2799,N_1250,N_1533);
xor U2800 (N_2800,N_1330,N_1958);
nand U2801 (N_2801,N_1299,N_1783);
nor U2802 (N_2802,N_1271,N_1879);
or U2803 (N_2803,N_1698,N_1541);
and U2804 (N_2804,N_1098,N_1218);
or U2805 (N_2805,N_1819,N_1032);
nand U2806 (N_2806,N_1710,N_1953);
nand U2807 (N_2807,N_1365,N_1478);
nand U2808 (N_2808,N_1192,N_1466);
xor U2809 (N_2809,N_1034,N_1711);
or U2810 (N_2810,N_1009,N_1618);
nand U2811 (N_2811,N_1178,N_1198);
xnor U2812 (N_2812,N_1771,N_1058);
or U2813 (N_2813,N_1520,N_1674);
nand U2814 (N_2814,N_1883,N_1623);
nand U2815 (N_2815,N_1351,N_1871);
nand U2816 (N_2816,N_1955,N_1435);
xnor U2817 (N_2817,N_1008,N_1321);
nor U2818 (N_2818,N_1342,N_1491);
nor U2819 (N_2819,N_1524,N_1449);
and U2820 (N_2820,N_1024,N_1215);
nor U2821 (N_2821,N_1106,N_1894);
nor U2822 (N_2822,N_1152,N_1126);
xnor U2823 (N_2823,N_1973,N_1583);
xor U2824 (N_2824,N_1481,N_1931);
nor U2825 (N_2825,N_1546,N_1011);
nor U2826 (N_2826,N_1935,N_1924);
xor U2827 (N_2827,N_1317,N_1530);
xor U2828 (N_2828,N_1692,N_1341);
nand U2829 (N_2829,N_1488,N_1915);
nand U2830 (N_2830,N_1008,N_1945);
and U2831 (N_2831,N_1211,N_1299);
nand U2832 (N_2832,N_1098,N_1270);
nor U2833 (N_2833,N_1178,N_1221);
nand U2834 (N_2834,N_1156,N_1897);
nor U2835 (N_2835,N_1703,N_1386);
or U2836 (N_2836,N_1402,N_1813);
xor U2837 (N_2837,N_1168,N_1833);
nor U2838 (N_2838,N_1778,N_1649);
nand U2839 (N_2839,N_1899,N_1303);
nand U2840 (N_2840,N_1211,N_1635);
nor U2841 (N_2841,N_1404,N_1624);
xor U2842 (N_2842,N_1512,N_1366);
xnor U2843 (N_2843,N_1608,N_1140);
nand U2844 (N_2844,N_1135,N_1333);
xor U2845 (N_2845,N_1772,N_1632);
xor U2846 (N_2846,N_1260,N_1742);
or U2847 (N_2847,N_1212,N_1531);
nor U2848 (N_2848,N_1406,N_1065);
nor U2849 (N_2849,N_1079,N_1237);
and U2850 (N_2850,N_1179,N_1040);
and U2851 (N_2851,N_1496,N_1649);
nor U2852 (N_2852,N_1048,N_1112);
nand U2853 (N_2853,N_1721,N_1554);
nand U2854 (N_2854,N_1256,N_1005);
nor U2855 (N_2855,N_1075,N_1688);
and U2856 (N_2856,N_1947,N_1484);
nor U2857 (N_2857,N_1990,N_1208);
nand U2858 (N_2858,N_1989,N_1593);
nor U2859 (N_2859,N_1267,N_1846);
or U2860 (N_2860,N_1381,N_1065);
nor U2861 (N_2861,N_1604,N_1677);
and U2862 (N_2862,N_1603,N_1077);
xor U2863 (N_2863,N_1031,N_1575);
xor U2864 (N_2864,N_1037,N_1657);
xor U2865 (N_2865,N_1946,N_1112);
nand U2866 (N_2866,N_1580,N_1147);
and U2867 (N_2867,N_1382,N_1704);
or U2868 (N_2868,N_1577,N_1556);
and U2869 (N_2869,N_1247,N_1898);
nor U2870 (N_2870,N_1133,N_1701);
xnor U2871 (N_2871,N_1548,N_1837);
and U2872 (N_2872,N_1852,N_1869);
nand U2873 (N_2873,N_1733,N_1732);
nor U2874 (N_2874,N_1881,N_1167);
or U2875 (N_2875,N_1073,N_1504);
nand U2876 (N_2876,N_1591,N_1376);
nand U2877 (N_2877,N_1140,N_1043);
nor U2878 (N_2878,N_1538,N_1374);
nor U2879 (N_2879,N_1604,N_1262);
nand U2880 (N_2880,N_1679,N_1507);
nand U2881 (N_2881,N_1101,N_1117);
nand U2882 (N_2882,N_1124,N_1079);
or U2883 (N_2883,N_1779,N_1290);
nand U2884 (N_2884,N_1374,N_1466);
xnor U2885 (N_2885,N_1918,N_1371);
nand U2886 (N_2886,N_1768,N_1286);
nand U2887 (N_2887,N_1365,N_1604);
nand U2888 (N_2888,N_1581,N_1278);
and U2889 (N_2889,N_1924,N_1393);
nand U2890 (N_2890,N_1081,N_1982);
nor U2891 (N_2891,N_1181,N_1073);
nor U2892 (N_2892,N_1239,N_1048);
or U2893 (N_2893,N_1680,N_1524);
nand U2894 (N_2894,N_1215,N_1216);
or U2895 (N_2895,N_1746,N_1099);
or U2896 (N_2896,N_1450,N_1452);
nor U2897 (N_2897,N_1902,N_1059);
or U2898 (N_2898,N_1027,N_1049);
and U2899 (N_2899,N_1557,N_1281);
nand U2900 (N_2900,N_1963,N_1050);
xnor U2901 (N_2901,N_1027,N_1336);
nand U2902 (N_2902,N_1129,N_1353);
nand U2903 (N_2903,N_1270,N_1109);
or U2904 (N_2904,N_1300,N_1884);
and U2905 (N_2905,N_1378,N_1188);
nor U2906 (N_2906,N_1431,N_1140);
xor U2907 (N_2907,N_1964,N_1427);
and U2908 (N_2908,N_1454,N_1865);
xor U2909 (N_2909,N_1294,N_1702);
or U2910 (N_2910,N_1515,N_1187);
or U2911 (N_2911,N_1192,N_1095);
and U2912 (N_2912,N_1430,N_1037);
xnor U2913 (N_2913,N_1338,N_1336);
nor U2914 (N_2914,N_1749,N_1514);
or U2915 (N_2915,N_1193,N_1674);
and U2916 (N_2916,N_1935,N_1241);
nand U2917 (N_2917,N_1300,N_1438);
or U2918 (N_2918,N_1337,N_1812);
nor U2919 (N_2919,N_1543,N_1207);
and U2920 (N_2920,N_1390,N_1310);
xor U2921 (N_2921,N_1809,N_1870);
xor U2922 (N_2922,N_1419,N_1078);
xor U2923 (N_2923,N_1185,N_1777);
nor U2924 (N_2924,N_1443,N_1114);
nand U2925 (N_2925,N_1612,N_1320);
and U2926 (N_2926,N_1512,N_1916);
and U2927 (N_2927,N_1589,N_1470);
nand U2928 (N_2928,N_1764,N_1576);
or U2929 (N_2929,N_1664,N_1755);
nand U2930 (N_2930,N_1106,N_1474);
or U2931 (N_2931,N_1724,N_1258);
nand U2932 (N_2932,N_1324,N_1674);
xor U2933 (N_2933,N_1891,N_1476);
and U2934 (N_2934,N_1996,N_1348);
or U2935 (N_2935,N_1984,N_1469);
nand U2936 (N_2936,N_1814,N_1155);
xor U2937 (N_2937,N_1793,N_1124);
xor U2938 (N_2938,N_1544,N_1162);
xor U2939 (N_2939,N_1799,N_1681);
nor U2940 (N_2940,N_1161,N_1992);
and U2941 (N_2941,N_1686,N_1894);
nor U2942 (N_2942,N_1547,N_1111);
xnor U2943 (N_2943,N_1178,N_1849);
nor U2944 (N_2944,N_1423,N_1053);
nand U2945 (N_2945,N_1569,N_1260);
or U2946 (N_2946,N_1451,N_1706);
or U2947 (N_2947,N_1884,N_1181);
nand U2948 (N_2948,N_1366,N_1763);
nand U2949 (N_2949,N_1222,N_1916);
and U2950 (N_2950,N_1229,N_1084);
xnor U2951 (N_2951,N_1930,N_1044);
and U2952 (N_2952,N_1818,N_1249);
nor U2953 (N_2953,N_1088,N_1785);
xor U2954 (N_2954,N_1301,N_1300);
or U2955 (N_2955,N_1747,N_1938);
xor U2956 (N_2956,N_1627,N_1302);
nand U2957 (N_2957,N_1797,N_1652);
nand U2958 (N_2958,N_1347,N_1991);
xor U2959 (N_2959,N_1269,N_1372);
nand U2960 (N_2960,N_1183,N_1207);
or U2961 (N_2961,N_1447,N_1104);
and U2962 (N_2962,N_1495,N_1631);
and U2963 (N_2963,N_1083,N_1301);
or U2964 (N_2964,N_1249,N_1902);
nor U2965 (N_2965,N_1275,N_1012);
nor U2966 (N_2966,N_1110,N_1556);
and U2967 (N_2967,N_1206,N_1749);
nor U2968 (N_2968,N_1769,N_1023);
nand U2969 (N_2969,N_1070,N_1353);
nor U2970 (N_2970,N_1958,N_1830);
xnor U2971 (N_2971,N_1548,N_1563);
and U2972 (N_2972,N_1318,N_1644);
xnor U2973 (N_2973,N_1535,N_1264);
xor U2974 (N_2974,N_1956,N_1565);
or U2975 (N_2975,N_1312,N_1514);
or U2976 (N_2976,N_1637,N_1290);
xor U2977 (N_2977,N_1444,N_1637);
xor U2978 (N_2978,N_1438,N_1653);
and U2979 (N_2979,N_1822,N_1271);
nor U2980 (N_2980,N_1977,N_1646);
nor U2981 (N_2981,N_1524,N_1381);
and U2982 (N_2982,N_1658,N_1293);
nand U2983 (N_2983,N_1058,N_1422);
or U2984 (N_2984,N_1517,N_1761);
xnor U2985 (N_2985,N_1308,N_1160);
xor U2986 (N_2986,N_1437,N_1716);
or U2987 (N_2987,N_1154,N_1657);
nand U2988 (N_2988,N_1861,N_1451);
nor U2989 (N_2989,N_1874,N_1586);
nand U2990 (N_2990,N_1963,N_1041);
or U2991 (N_2991,N_1035,N_1532);
xor U2992 (N_2992,N_1469,N_1032);
nor U2993 (N_2993,N_1707,N_1635);
nand U2994 (N_2994,N_1796,N_1755);
and U2995 (N_2995,N_1091,N_1478);
nand U2996 (N_2996,N_1336,N_1620);
or U2997 (N_2997,N_1187,N_1348);
nor U2998 (N_2998,N_1882,N_1546);
nor U2999 (N_2999,N_1740,N_1059);
nand U3000 (N_3000,N_2206,N_2606);
xnor U3001 (N_3001,N_2719,N_2250);
and U3002 (N_3002,N_2420,N_2360);
xnor U3003 (N_3003,N_2462,N_2866);
nor U3004 (N_3004,N_2991,N_2044);
nor U3005 (N_3005,N_2026,N_2445);
nand U3006 (N_3006,N_2262,N_2550);
and U3007 (N_3007,N_2123,N_2717);
nand U3008 (N_3008,N_2261,N_2336);
and U3009 (N_3009,N_2624,N_2192);
nand U3010 (N_3010,N_2549,N_2100);
nand U3011 (N_3011,N_2040,N_2971);
nand U3012 (N_3012,N_2503,N_2332);
and U3013 (N_3013,N_2917,N_2881);
and U3014 (N_3014,N_2337,N_2467);
nand U3015 (N_3015,N_2022,N_2576);
or U3016 (N_3016,N_2778,N_2290);
and U3017 (N_3017,N_2889,N_2253);
xor U3018 (N_3018,N_2615,N_2754);
and U3019 (N_3019,N_2797,N_2543);
xnor U3020 (N_3020,N_2806,N_2659);
or U3021 (N_3021,N_2374,N_2820);
and U3022 (N_3022,N_2449,N_2484);
xor U3023 (N_3023,N_2024,N_2311);
xor U3024 (N_3024,N_2498,N_2059);
nor U3025 (N_3025,N_2201,N_2354);
or U3026 (N_3026,N_2494,N_2007);
and U3027 (N_3027,N_2070,N_2173);
xnor U3028 (N_3028,N_2531,N_2637);
and U3029 (N_3029,N_2214,N_2695);
nor U3030 (N_3030,N_2565,N_2838);
nand U3031 (N_3031,N_2929,N_2181);
nand U3032 (N_3032,N_2770,N_2443);
nand U3033 (N_3033,N_2135,N_2194);
and U3034 (N_3034,N_2987,N_2692);
nor U3035 (N_3035,N_2776,N_2456);
or U3036 (N_3036,N_2865,N_2678);
xor U3037 (N_3037,N_2712,N_2595);
and U3038 (N_3038,N_2108,N_2897);
or U3039 (N_3039,N_2249,N_2003);
or U3040 (N_3040,N_2620,N_2874);
and U3041 (N_3041,N_2020,N_2793);
or U3042 (N_3042,N_2068,N_2720);
nor U3043 (N_3043,N_2621,N_2184);
or U3044 (N_3044,N_2483,N_2682);
and U3045 (N_3045,N_2441,N_2221);
xor U3046 (N_3046,N_2023,N_2087);
nor U3047 (N_3047,N_2736,N_2145);
nand U3048 (N_3048,N_2422,N_2398);
xor U3049 (N_3049,N_2223,N_2168);
and U3050 (N_3050,N_2744,N_2596);
and U3051 (N_3051,N_2907,N_2120);
and U3052 (N_3052,N_2156,N_2506);
or U3053 (N_3053,N_2153,N_2718);
xnor U3054 (N_3054,N_2780,N_2801);
and U3055 (N_3055,N_2928,N_2590);
xor U3056 (N_3056,N_2243,N_2798);
nand U3057 (N_3057,N_2492,N_2419);
and U3058 (N_3058,N_2064,N_2157);
or U3059 (N_3059,N_2365,N_2603);
nor U3060 (N_3060,N_2564,N_2571);
nor U3061 (N_3061,N_2132,N_2459);
xnor U3062 (N_3062,N_2623,N_2700);
and U3063 (N_3063,N_2488,N_2705);
or U3064 (N_3064,N_2957,N_2774);
nor U3065 (N_3065,N_2371,N_2964);
xor U3066 (N_3066,N_2500,N_2724);
nor U3067 (N_3067,N_2322,N_2179);
and U3068 (N_3068,N_2267,N_2055);
nor U3069 (N_3069,N_2584,N_2217);
and U3070 (N_3070,N_2393,N_2187);
or U3071 (N_3071,N_2517,N_2539);
or U3072 (N_3072,N_2349,N_2034);
nor U3073 (N_3073,N_2491,N_2417);
nor U3074 (N_3074,N_2756,N_2962);
or U3075 (N_3075,N_2481,N_2742);
nor U3076 (N_3076,N_2256,N_2418);
xor U3077 (N_3077,N_2979,N_2379);
nand U3078 (N_3078,N_2010,N_2893);
nor U3079 (N_3079,N_2788,N_2434);
and U3080 (N_3080,N_2739,N_2279);
or U3081 (N_3081,N_2380,N_2828);
nor U3082 (N_3082,N_2972,N_2876);
or U3083 (N_3083,N_2499,N_2288);
or U3084 (N_3084,N_2661,N_2586);
nand U3085 (N_3085,N_2813,N_2092);
nand U3086 (N_3086,N_2077,N_2567);
xnor U3087 (N_3087,N_2170,N_2944);
and U3088 (N_3088,N_2570,N_2910);
nor U3089 (N_3089,N_2468,N_2836);
xnor U3090 (N_3090,N_2293,N_2004);
nand U3091 (N_3091,N_2954,N_2761);
and U3092 (N_3092,N_2591,N_2284);
xor U3093 (N_3093,N_2631,N_2103);
or U3094 (N_3094,N_2205,N_2746);
xor U3095 (N_3095,N_2189,N_2296);
xor U3096 (N_3096,N_2572,N_2435);
nor U3097 (N_3097,N_2509,N_2347);
nor U3098 (N_3098,N_2822,N_2653);
nor U3099 (N_3099,N_2546,N_2588);
nor U3100 (N_3100,N_2630,N_2628);
and U3101 (N_3101,N_2106,N_2837);
nor U3102 (N_3102,N_2751,N_2924);
nor U3103 (N_3103,N_2704,N_2901);
nor U3104 (N_3104,N_2834,N_2921);
and U3105 (N_3105,N_2966,N_2554);
nand U3106 (N_3106,N_2018,N_2952);
xnor U3107 (N_3107,N_2320,N_2016);
xor U3108 (N_3108,N_2597,N_2592);
xnor U3109 (N_3109,N_2264,N_2232);
nor U3110 (N_3110,N_2299,N_2846);
xor U3111 (N_3111,N_2263,N_2860);
xnor U3112 (N_3112,N_2461,N_2457);
and U3113 (N_3113,N_2297,N_2812);
nor U3114 (N_3114,N_2392,N_2873);
nand U3115 (N_3115,N_2903,N_2460);
nand U3116 (N_3116,N_2634,N_2415);
xnor U3117 (N_3117,N_2314,N_2555);
nor U3118 (N_3118,N_2547,N_2162);
nand U3119 (N_3119,N_2969,N_2672);
and U3120 (N_3120,N_2961,N_2790);
or U3121 (N_3121,N_2052,N_2946);
nand U3122 (N_3122,N_2765,N_2622);
nand U3123 (N_3123,N_2519,N_2078);
nor U3124 (N_3124,N_2625,N_2376);
nand U3125 (N_3125,N_2632,N_2088);
nor U3126 (N_3126,N_2920,N_2098);
or U3127 (N_3127,N_2548,N_2617);
xnor U3128 (N_3128,N_2673,N_2696);
xor U3129 (N_3129,N_2829,N_2502);
or U3130 (N_3130,N_2760,N_2694);
nand U3131 (N_3131,N_2286,N_2265);
or U3132 (N_3132,N_2693,N_2755);
nor U3133 (N_3133,N_2729,N_2891);
or U3134 (N_3134,N_2489,N_2627);
nor U3135 (N_3135,N_2394,N_2520);
and U3136 (N_3136,N_2438,N_2803);
and U3137 (N_3137,N_2741,N_2312);
nand U3138 (N_3138,N_2691,N_2183);
xnor U3139 (N_3139,N_2421,N_2568);
nand U3140 (N_3140,N_2633,N_2686);
or U3141 (N_3141,N_2166,N_2626);
nor U3142 (N_3142,N_2259,N_2497);
nor U3143 (N_3143,N_2642,N_2442);
and U3144 (N_3144,N_2252,N_2389);
and U3145 (N_3145,N_2171,N_2285);
and U3146 (N_3146,N_2953,N_2242);
nand U3147 (N_3147,N_2525,N_2681);
nor U3148 (N_3148,N_2839,N_2282);
xor U3149 (N_3149,N_2799,N_2992);
or U3150 (N_3150,N_2976,N_2999);
and U3151 (N_3151,N_2104,N_2875);
or U3152 (N_3152,N_2527,N_2802);
nand U3153 (N_3153,N_2240,N_2896);
and U3154 (N_3154,N_2919,N_2446);
nand U3155 (N_3155,N_2951,N_2725);
nand U3156 (N_3156,N_2099,N_2825);
nand U3157 (N_3157,N_2167,N_2819);
xnor U3158 (N_3158,N_2469,N_2308);
and U3159 (N_3159,N_2786,N_2902);
nor U3160 (N_3160,N_2111,N_2702);
or U3161 (N_3161,N_2072,N_2847);
or U3162 (N_3162,N_2811,N_2649);
xnor U3163 (N_3163,N_2967,N_2378);
xnor U3164 (N_3164,N_2607,N_2333);
xnor U3165 (N_3165,N_2769,N_2529);
xor U3166 (N_3166,N_2130,N_2067);
nand U3167 (N_3167,N_2413,N_2660);
nor U3168 (N_3168,N_2960,N_2747);
and U3169 (N_3169,N_2056,N_2410);
nor U3170 (N_3170,N_2644,N_2496);
or U3171 (N_3171,N_2504,N_2589);
or U3172 (N_3172,N_2204,N_2028);
nor U3173 (N_3173,N_2313,N_2149);
xnor U3174 (N_3174,N_2058,N_2368);
xor U3175 (N_3175,N_2523,N_2164);
and U3176 (N_3176,N_2083,N_2609);
and U3177 (N_3177,N_2391,N_2594);
nor U3178 (N_3178,N_2940,N_2464);
xnor U3179 (N_3179,N_2518,N_2352);
and U3180 (N_3180,N_2001,N_2050);
xor U3181 (N_3181,N_2863,N_2941);
xor U3182 (N_3182,N_2241,N_2683);
or U3183 (N_3183,N_2090,N_2619);
nand U3184 (N_3184,N_2711,N_2880);
nand U3185 (N_3185,N_2269,N_2689);
nand U3186 (N_3186,N_2832,N_2515);
nor U3187 (N_3187,N_2292,N_2791);
and U3188 (N_3188,N_2931,N_2089);
nand U3189 (N_3189,N_2722,N_2664);
nor U3190 (N_3190,N_2213,N_2381);
and U3191 (N_3191,N_2854,N_2914);
nand U3192 (N_3192,N_2476,N_2824);
and U3193 (N_3193,N_2408,N_2033);
and U3194 (N_3194,N_2465,N_2327);
xor U3195 (N_3195,N_2447,N_2879);
and U3196 (N_3196,N_2716,N_2015);
or U3197 (N_3197,N_2763,N_2043);
nor U3198 (N_3198,N_2403,N_2859);
nand U3199 (N_3199,N_2444,N_2122);
nor U3200 (N_3200,N_2886,N_2738);
nor U3201 (N_3201,N_2175,N_2566);
and U3202 (N_3202,N_2244,N_2735);
or U3203 (N_3203,N_2508,N_2767);
and U3204 (N_3204,N_2377,N_2562);
and U3205 (N_3205,N_2593,N_2757);
nor U3206 (N_3206,N_2815,N_2151);
nor U3207 (N_3207,N_2382,N_2493);
nor U3208 (N_3208,N_2762,N_2795);
nand U3209 (N_3209,N_2406,N_2871);
nand U3210 (N_3210,N_2121,N_2017);
nor U3211 (N_3211,N_2580,N_2582);
or U3212 (N_3212,N_2198,N_2236);
nor U3213 (N_3213,N_2323,N_2317);
and U3214 (N_3214,N_2578,N_2247);
nor U3215 (N_3215,N_2538,N_2697);
nand U3216 (N_3216,N_2909,N_2703);
nand U3217 (N_3217,N_2480,N_2366);
and U3218 (N_3218,N_2316,N_2350);
xnor U3219 (N_3219,N_2983,N_2390);
nor U3220 (N_3220,N_2611,N_2933);
or U3221 (N_3221,N_2107,N_2387);
nand U3222 (N_3222,N_2600,N_2309);
nand U3223 (N_3223,N_2161,N_2848);
or U3224 (N_3224,N_2598,N_2861);
nor U3225 (N_3225,N_2521,N_2061);
or U3226 (N_3226,N_2396,N_2537);
and U3227 (N_3227,N_2490,N_2911);
nand U3228 (N_3228,N_2726,N_2129);
nand U3229 (N_3229,N_2388,N_2342);
and U3230 (N_3230,N_2709,N_2195);
nand U3231 (N_3231,N_2690,N_2516);
xnor U3232 (N_3232,N_2974,N_2669);
xor U3233 (N_3233,N_2759,N_2344);
xnor U3234 (N_3234,N_2950,N_2160);
xor U3235 (N_3235,N_2916,N_2027);
xor U3236 (N_3236,N_2199,N_2021);
nor U3237 (N_3237,N_2101,N_2036);
or U3238 (N_3238,N_2049,N_2321);
nand U3239 (N_3239,N_2535,N_2601);
and U3240 (N_3240,N_2330,N_2677);
nor U3241 (N_3241,N_2948,N_2805);
nor U3242 (N_3242,N_2370,N_2000);
or U3243 (N_3243,N_2857,N_2215);
xnor U3244 (N_3244,N_2533,N_2125);
or U3245 (N_3245,N_2610,N_2714);
xor U3246 (N_3246,N_2781,N_2472);
and U3247 (N_3247,N_2348,N_2266);
and U3248 (N_3248,N_2012,N_2958);
or U3249 (N_3249,N_2715,N_2039);
xnor U3250 (N_3250,N_2466,N_2994);
or U3251 (N_3251,N_2947,N_2890);
and U3252 (N_3252,N_2985,N_2830);
or U3253 (N_3253,N_2512,N_2656);
nand U3254 (N_3254,N_2884,N_2645);
or U3255 (N_3255,N_2577,N_2478);
or U3256 (N_3256,N_2455,N_2667);
nor U3257 (N_3257,N_2114,N_2850);
and U3258 (N_3258,N_2110,N_2208);
nor U3259 (N_3259,N_2339,N_2237);
nand U3260 (N_3260,N_2505,N_2808);
nand U3261 (N_3261,N_2638,N_2325);
nor U3262 (N_3262,N_2084,N_2687);
and U3263 (N_3263,N_2305,N_2477);
or U3264 (N_3264,N_2530,N_2710);
and U3265 (N_3265,N_2202,N_2454);
or U3266 (N_3266,N_2427,N_2431);
and U3267 (N_3267,N_2923,N_2984);
xor U3268 (N_3268,N_2915,N_2654);
or U3269 (N_3269,N_2556,N_2423);
and U3270 (N_3270,N_2732,N_2275);
and U3271 (N_3271,N_2180,N_2340);
nor U3272 (N_3272,N_2045,N_2826);
and U3273 (N_3273,N_2258,N_2126);
and U3274 (N_3274,N_2482,N_2587);
xnor U3275 (N_3275,N_2112,N_2425);
nand U3276 (N_3276,N_2796,N_2599);
and U3277 (N_3277,N_2248,N_2817);
xnor U3278 (N_3278,N_2163,N_2009);
nor U3279 (N_3279,N_2605,N_2764);
nor U3280 (N_3280,N_2440,N_2988);
and U3281 (N_3281,N_2225,N_2536);
or U3282 (N_3282,N_2959,N_2351);
xnor U3283 (N_3283,N_2925,N_2663);
xnor U3284 (N_3284,N_2137,N_2032);
xor U3285 (N_3285,N_2066,N_2641);
or U3286 (N_3286,N_2142,N_2646);
and U3287 (N_3287,N_2116,N_2783);
nor U3288 (N_3288,N_2291,N_2804);
and U3289 (N_3289,N_2949,N_2479);
and U3290 (N_3290,N_2560,N_2772);
and U3291 (N_3291,N_2864,N_2355);
xor U3292 (N_3292,N_2583,N_2361);
nand U3293 (N_3293,N_2346,N_2768);
and U3294 (N_3294,N_2289,N_2684);
or U3295 (N_3295,N_2113,N_2436);
and U3296 (N_3296,N_2437,N_2143);
nor U3297 (N_3297,N_2154,N_2616);
or U3298 (N_3298,N_2750,N_2287);
xor U3299 (N_3299,N_2298,N_2172);
xnor U3300 (N_3300,N_2532,N_2074);
xnor U3301 (N_3301,N_2118,N_2397);
nand U3302 (N_3302,N_2414,N_2485);
nor U3303 (N_3303,N_2063,N_2251);
nor U3304 (N_3304,N_2670,N_2109);
nor U3305 (N_3305,N_2727,N_2816);
xor U3306 (N_3306,N_2981,N_2668);
and U3307 (N_3307,N_2307,N_2989);
xor U3308 (N_3308,N_2785,N_2561);
and U3309 (N_3309,N_2662,N_2939);
xor U3310 (N_3310,N_2883,N_2773);
or U3311 (N_3311,N_2405,N_2574);
nor U3312 (N_3312,N_2930,N_2014);
xor U3313 (N_3313,N_2060,N_2869);
nor U3314 (N_3314,N_2943,N_2159);
nand U3315 (N_3315,N_2006,N_2229);
xnor U3316 (N_3316,N_2048,N_2424);
and U3317 (N_3317,N_2216,N_2524);
nand U3318 (N_3318,N_2526,N_2495);
or U3319 (N_3319,N_2051,N_2094);
or U3320 (N_3320,N_2775,N_2190);
nand U3321 (N_3321,N_2986,N_2233);
nand U3322 (N_3322,N_2823,N_2272);
xnor U3323 (N_3323,N_2185,N_2463);
and U3324 (N_3324,N_2385,N_2450);
nor U3325 (N_3325,N_2618,N_2399);
xor U3326 (N_3326,N_2035,N_2581);
nand U3327 (N_3327,N_2220,N_2053);
nor U3328 (N_3328,N_2341,N_2230);
and U3329 (N_3329,N_2737,N_2679);
or U3330 (N_3330,N_2038,N_2219);
or U3331 (N_3331,N_2193,N_2302);
nor U3332 (N_3332,N_2698,N_2671);
nor U3333 (N_3333,N_2970,N_2510);
nor U3334 (N_3334,N_2150,N_2882);
and U3335 (N_3335,N_2085,N_2655);
and U3336 (N_3336,N_2973,N_2271);
nand U3337 (N_3337,N_2228,N_2528);
or U3338 (N_3338,N_2814,N_2752);
nand U3339 (N_3339,N_2575,N_2995);
nand U3340 (N_3340,N_2963,N_2658);
xnor U3341 (N_3341,N_2428,N_2501);
or U3342 (N_3342,N_2993,N_2073);
xnor U3343 (N_3343,N_2766,N_2842);
nand U3344 (N_3344,N_2551,N_2614);
nand U3345 (N_3345,N_2097,N_2648);
nand U3346 (N_3346,N_2643,N_2294);
and U3347 (N_3347,N_2281,N_2133);
xnor U3348 (N_3348,N_2522,N_2174);
nand U3349 (N_3349,N_2375,N_2942);
nor U3350 (N_3350,N_2276,N_2545);
or U3351 (N_3351,N_2395,N_2926);
and U3352 (N_3352,N_2856,N_2870);
xnor U3353 (N_3353,N_2277,N_2409);
and U3354 (N_3354,N_2412,N_2639);
nor U3355 (N_3355,N_2980,N_2810);
nor U3356 (N_3356,N_2912,N_2486);
xnor U3357 (N_3357,N_2753,N_2473);
and U3358 (N_3358,N_2862,N_2025);
nand U3359 (N_3359,N_2140,N_2065);
nand U3360 (N_3360,N_2845,N_2978);
nand U3361 (N_3361,N_2934,N_2707);
and U3362 (N_3362,N_2013,N_2807);
and U3363 (N_3363,N_2226,N_2868);
nor U3364 (N_3364,N_2784,N_2148);
nand U3365 (N_3365,N_2471,N_2260);
nor U3366 (N_3366,N_2833,N_2008);
nand U3367 (N_3367,N_2407,N_2867);
or U3368 (N_3368,N_2840,N_2573);
nor U3369 (N_3369,N_2657,N_2274);
and U3370 (N_3370,N_2900,N_2743);
nor U3371 (N_3371,N_2115,N_2326);
or U3372 (N_3372,N_2334,N_2134);
nor U3373 (N_3373,N_2429,N_2602);
nor U3374 (N_3374,N_2372,N_2404);
and U3375 (N_3375,N_2268,N_2373);
and U3376 (N_3376,N_2885,N_2283);
nand U3377 (N_3377,N_2069,N_2042);
xnor U3378 (N_3378,N_2936,N_2758);
and U3379 (N_3379,N_2888,N_2304);
nand U3380 (N_3380,N_2188,N_2075);
nand U3381 (N_3381,N_2922,N_2635);
nor U3382 (N_3382,N_2777,N_2779);
nand U3383 (N_3383,N_2734,N_2892);
xnor U3384 (N_3384,N_2386,N_2701);
or U3385 (N_3385,N_2029,N_2794);
and U3386 (N_3386,N_2451,N_2977);
or U3387 (N_3387,N_2629,N_2511);
nor U3388 (N_3388,N_2270,N_2945);
xor U3389 (N_3389,N_2353,N_2218);
nor U3390 (N_3390,N_2918,N_2932);
nor U3391 (N_3391,N_2362,N_2328);
or U3392 (N_3392,N_2367,N_2238);
xor U3393 (N_3393,N_2182,N_2563);
nor U3394 (N_3394,N_2165,N_2843);
nor U3395 (N_3395,N_2740,N_2534);
nand U3396 (N_3396,N_2086,N_2728);
nand U3397 (N_3397,N_2818,N_2851);
or U3398 (N_3398,N_2212,N_2146);
or U3399 (N_3399,N_2255,N_2310);
or U3400 (N_3400,N_2138,N_2031);
or U3401 (N_3401,N_2913,N_2513);
and U3402 (N_3402,N_2191,N_2558);
nand U3403 (N_3403,N_2895,N_2057);
nor U3404 (N_3404,N_2080,N_2877);
or U3405 (N_3405,N_2675,N_2329);
nand U3406 (N_3406,N_2540,N_2062);
or U3407 (N_3407,N_2047,N_2699);
or U3408 (N_3408,N_2169,N_2082);
nand U3409 (N_3409,N_2127,N_2612);
or U3410 (N_3410,N_2507,N_2005);
xor U3411 (N_3411,N_2652,N_2585);
xnor U3412 (N_3412,N_2608,N_2666);
and U3413 (N_3413,N_2343,N_2904);
nor U3414 (N_3414,N_2178,N_2899);
nand U3415 (N_3415,N_2894,N_2095);
or U3416 (N_3416,N_2731,N_2458);
nor U3417 (N_3417,N_2782,N_2831);
xnor U3418 (N_3418,N_2651,N_2079);
nor U3419 (N_3419,N_2384,N_2853);
or U3420 (N_3420,N_2105,N_2898);
xor U3421 (N_3421,N_2002,N_2997);
and U3422 (N_3422,N_2432,N_2359);
or U3423 (N_3423,N_2723,N_2800);
or U3424 (N_3424,N_2541,N_2426);
or U3425 (N_3425,N_2273,N_2306);
and U3426 (N_3426,N_2186,N_2557);
nor U3427 (N_3427,N_2955,N_2400);
nor U3428 (N_3428,N_2730,N_2071);
xor U3429 (N_3429,N_2054,N_2358);
or U3430 (N_3430,N_2745,N_2542);
nand U3431 (N_3431,N_2155,N_2210);
nand U3432 (N_3432,N_2552,N_2096);
or U3433 (N_3433,N_2433,N_2245);
or U3434 (N_3434,N_2878,N_2514);
nor U3435 (N_3435,N_2345,N_2324);
or U3436 (N_3436,N_2771,N_2835);
or U3437 (N_3437,N_2748,N_2301);
xnor U3438 (N_3438,N_2119,N_2319);
and U3439 (N_3439,N_2544,N_2102);
or U3440 (N_3440,N_2402,N_2235);
xnor U3441 (N_3441,N_2613,N_2401);
xor U3442 (N_3442,N_2474,N_2996);
and U3443 (N_3443,N_2676,N_2076);
and U3444 (N_3444,N_2211,N_2430);
nand U3445 (N_3445,N_2559,N_2280);
nand U3446 (N_3446,N_2196,N_2295);
and U3447 (N_3447,N_2685,N_2411);
nand U3448 (N_3448,N_2141,N_2224);
and U3449 (N_3449,N_2733,N_2300);
nand U3450 (N_3450,N_2453,N_2369);
nor U3451 (N_3451,N_2363,N_2650);
nor U3452 (N_3452,N_2030,N_2357);
and U3453 (N_3453,N_2278,N_2091);
nor U3454 (N_3454,N_2855,N_2246);
nor U3455 (N_3455,N_2139,N_2315);
nand U3456 (N_3456,N_2207,N_2688);
xnor U3457 (N_3457,N_2553,N_2203);
or U3458 (N_3458,N_2680,N_2257);
and U3459 (N_3459,N_2093,N_2222);
and U3460 (N_3460,N_2227,N_2338);
nor U3461 (N_3461,N_2965,N_2046);
xnor U3462 (N_3462,N_2197,N_2849);
or U3463 (N_3463,N_2708,N_2416);
xor U3464 (N_3464,N_2579,N_2858);
xor U3465 (N_3465,N_2124,N_2131);
xnor U3466 (N_3466,N_2905,N_2117);
xnor U3467 (N_3467,N_2908,N_2674);
or U3468 (N_3468,N_2844,N_2239);
nor U3469 (N_3469,N_2128,N_2990);
xnor U3470 (N_3470,N_2136,N_2927);
nand U3471 (N_3471,N_2439,N_2152);
xor U3472 (N_3472,N_2636,N_2147);
nand U3473 (N_3473,N_2231,N_2841);
nand U3474 (N_3474,N_2318,N_2640);
nor U3475 (N_3475,N_2647,N_2713);
nor U3476 (N_3476,N_2158,N_2037);
nor U3477 (N_3477,N_2081,N_2383);
nor U3478 (N_3478,N_2364,N_2749);
nand U3479 (N_3479,N_2144,N_2487);
nor U3480 (N_3480,N_2968,N_2176);
and U3481 (N_3481,N_2827,N_2569);
nor U3482 (N_3482,N_2019,N_2041);
or U3483 (N_3483,N_2975,N_2887);
or U3484 (N_3484,N_2792,N_2935);
nor U3485 (N_3485,N_2200,N_2254);
nand U3486 (N_3486,N_2706,N_2721);
or U3487 (N_3487,N_2303,N_2938);
nor U3488 (N_3488,N_2475,N_2177);
and U3489 (N_3489,N_2982,N_2787);
xnor U3490 (N_3490,N_2821,N_2452);
or U3491 (N_3491,N_2470,N_2872);
xnor U3492 (N_3492,N_2789,N_2335);
nor U3493 (N_3493,N_2956,N_2331);
or U3494 (N_3494,N_2209,N_2665);
xnor U3495 (N_3495,N_2998,N_2906);
nand U3496 (N_3496,N_2809,N_2604);
and U3497 (N_3497,N_2356,N_2011);
nand U3498 (N_3498,N_2448,N_2234);
xor U3499 (N_3499,N_2852,N_2937);
and U3500 (N_3500,N_2777,N_2353);
or U3501 (N_3501,N_2541,N_2146);
or U3502 (N_3502,N_2312,N_2638);
xnor U3503 (N_3503,N_2906,N_2990);
and U3504 (N_3504,N_2980,N_2180);
nand U3505 (N_3505,N_2700,N_2213);
or U3506 (N_3506,N_2808,N_2086);
or U3507 (N_3507,N_2819,N_2333);
xnor U3508 (N_3508,N_2242,N_2511);
xnor U3509 (N_3509,N_2637,N_2062);
nor U3510 (N_3510,N_2973,N_2355);
and U3511 (N_3511,N_2274,N_2467);
or U3512 (N_3512,N_2121,N_2840);
xnor U3513 (N_3513,N_2548,N_2316);
or U3514 (N_3514,N_2931,N_2262);
nand U3515 (N_3515,N_2966,N_2459);
or U3516 (N_3516,N_2068,N_2808);
nor U3517 (N_3517,N_2060,N_2537);
and U3518 (N_3518,N_2209,N_2657);
nand U3519 (N_3519,N_2371,N_2342);
and U3520 (N_3520,N_2997,N_2711);
or U3521 (N_3521,N_2704,N_2737);
xnor U3522 (N_3522,N_2555,N_2758);
or U3523 (N_3523,N_2092,N_2930);
nor U3524 (N_3524,N_2767,N_2905);
xnor U3525 (N_3525,N_2118,N_2161);
nand U3526 (N_3526,N_2455,N_2580);
nor U3527 (N_3527,N_2443,N_2789);
nand U3528 (N_3528,N_2538,N_2859);
and U3529 (N_3529,N_2466,N_2011);
and U3530 (N_3530,N_2428,N_2557);
xor U3531 (N_3531,N_2610,N_2009);
and U3532 (N_3532,N_2774,N_2256);
xnor U3533 (N_3533,N_2492,N_2152);
nor U3534 (N_3534,N_2615,N_2177);
xor U3535 (N_3535,N_2828,N_2867);
nand U3536 (N_3536,N_2247,N_2923);
nor U3537 (N_3537,N_2317,N_2735);
nor U3538 (N_3538,N_2199,N_2275);
nor U3539 (N_3539,N_2864,N_2487);
or U3540 (N_3540,N_2123,N_2711);
xnor U3541 (N_3541,N_2383,N_2000);
nand U3542 (N_3542,N_2122,N_2457);
xnor U3543 (N_3543,N_2544,N_2640);
nor U3544 (N_3544,N_2437,N_2450);
nor U3545 (N_3545,N_2734,N_2592);
nand U3546 (N_3546,N_2994,N_2672);
or U3547 (N_3547,N_2440,N_2332);
xnor U3548 (N_3548,N_2084,N_2211);
xor U3549 (N_3549,N_2892,N_2327);
nand U3550 (N_3550,N_2578,N_2640);
nand U3551 (N_3551,N_2860,N_2901);
nand U3552 (N_3552,N_2297,N_2326);
xor U3553 (N_3553,N_2768,N_2804);
nand U3554 (N_3554,N_2558,N_2262);
and U3555 (N_3555,N_2522,N_2460);
or U3556 (N_3556,N_2220,N_2239);
xor U3557 (N_3557,N_2066,N_2691);
nand U3558 (N_3558,N_2750,N_2282);
xor U3559 (N_3559,N_2942,N_2392);
xnor U3560 (N_3560,N_2696,N_2873);
nor U3561 (N_3561,N_2472,N_2382);
or U3562 (N_3562,N_2897,N_2095);
xor U3563 (N_3563,N_2145,N_2496);
nand U3564 (N_3564,N_2158,N_2231);
nor U3565 (N_3565,N_2886,N_2541);
or U3566 (N_3566,N_2312,N_2840);
nor U3567 (N_3567,N_2786,N_2156);
xnor U3568 (N_3568,N_2117,N_2423);
and U3569 (N_3569,N_2594,N_2670);
and U3570 (N_3570,N_2455,N_2105);
xnor U3571 (N_3571,N_2695,N_2045);
nand U3572 (N_3572,N_2925,N_2986);
nand U3573 (N_3573,N_2313,N_2765);
and U3574 (N_3574,N_2234,N_2380);
or U3575 (N_3575,N_2756,N_2134);
nor U3576 (N_3576,N_2707,N_2273);
or U3577 (N_3577,N_2410,N_2987);
nand U3578 (N_3578,N_2417,N_2096);
or U3579 (N_3579,N_2691,N_2957);
xor U3580 (N_3580,N_2884,N_2801);
nand U3581 (N_3581,N_2794,N_2709);
nor U3582 (N_3582,N_2756,N_2312);
and U3583 (N_3583,N_2915,N_2598);
or U3584 (N_3584,N_2456,N_2669);
xnor U3585 (N_3585,N_2736,N_2208);
or U3586 (N_3586,N_2113,N_2261);
xnor U3587 (N_3587,N_2388,N_2766);
or U3588 (N_3588,N_2125,N_2613);
nand U3589 (N_3589,N_2254,N_2421);
xnor U3590 (N_3590,N_2175,N_2616);
and U3591 (N_3591,N_2433,N_2740);
or U3592 (N_3592,N_2259,N_2407);
xnor U3593 (N_3593,N_2666,N_2263);
nor U3594 (N_3594,N_2549,N_2401);
or U3595 (N_3595,N_2541,N_2048);
and U3596 (N_3596,N_2291,N_2803);
nor U3597 (N_3597,N_2718,N_2215);
xnor U3598 (N_3598,N_2723,N_2882);
xor U3599 (N_3599,N_2213,N_2854);
xor U3600 (N_3600,N_2822,N_2389);
xnor U3601 (N_3601,N_2284,N_2126);
nand U3602 (N_3602,N_2808,N_2275);
xor U3603 (N_3603,N_2951,N_2718);
nor U3604 (N_3604,N_2709,N_2111);
nor U3605 (N_3605,N_2699,N_2154);
and U3606 (N_3606,N_2274,N_2301);
or U3607 (N_3607,N_2705,N_2660);
or U3608 (N_3608,N_2993,N_2463);
or U3609 (N_3609,N_2592,N_2460);
nand U3610 (N_3610,N_2474,N_2046);
and U3611 (N_3611,N_2920,N_2796);
nor U3612 (N_3612,N_2682,N_2674);
or U3613 (N_3613,N_2209,N_2010);
xor U3614 (N_3614,N_2931,N_2208);
xor U3615 (N_3615,N_2462,N_2441);
or U3616 (N_3616,N_2885,N_2574);
xor U3617 (N_3617,N_2906,N_2227);
and U3618 (N_3618,N_2541,N_2083);
xnor U3619 (N_3619,N_2321,N_2670);
or U3620 (N_3620,N_2022,N_2980);
nor U3621 (N_3621,N_2367,N_2749);
or U3622 (N_3622,N_2140,N_2842);
nor U3623 (N_3623,N_2569,N_2453);
or U3624 (N_3624,N_2402,N_2431);
and U3625 (N_3625,N_2698,N_2244);
nand U3626 (N_3626,N_2996,N_2504);
nor U3627 (N_3627,N_2320,N_2232);
xnor U3628 (N_3628,N_2630,N_2335);
nand U3629 (N_3629,N_2432,N_2250);
nand U3630 (N_3630,N_2920,N_2462);
or U3631 (N_3631,N_2612,N_2658);
nor U3632 (N_3632,N_2936,N_2927);
or U3633 (N_3633,N_2539,N_2141);
nor U3634 (N_3634,N_2910,N_2779);
nand U3635 (N_3635,N_2927,N_2629);
and U3636 (N_3636,N_2779,N_2106);
nand U3637 (N_3637,N_2385,N_2810);
or U3638 (N_3638,N_2347,N_2383);
or U3639 (N_3639,N_2573,N_2596);
xor U3640 (N_3640,N_2120,N_2623);
xnor U3641 (N_3641,N_2039,N_2721);
nand U3642 (N_3642,N_2110,N_2274);
xor U3643 (N_3643,N_2417,N_2984);
nor U3644 (N_3644,N_2980,N_2767);
and U3645 (N_3645,N_2625,N_2722);
and U3646 (N_3646,N_2106,N_2076);
nor U3647 (N_3647,N_2383,N_2197);
xor U3648 (N_3648,N_2781,N_2325);
nand U3649 (N_3649,N_2911,N_2965);
and U3650 (N_3650,N_2516,N_2268);
nand U3651 (N_3651,N_2414,N_2577);
nor U3652 (N_3652,N_2096,N_2254);
nor U3653 (N_3653,N_2334,N_2684);
or U3654 (N_3654,N_2757,N_2037);
and U3655 (N_3655,N_2329,N_2337);
nor U3656 (N_3656,N_2457,N_2642);
nor U3657 (N_3657,N_2105,N_2267);
or U3658 (N_3658,N_2629,N_2736);
xor U3659 (N_3659,N_2862,N_2143);
or U3660 (N_3660,N_2379,N_2146);
xnor U3661 (N_3661,N_2240,N_2860);
xor U3662 (N_3662,N_2939,N_2872);
and U3663 (N_3663,N_2220,N_2614);
or U3664 (N_3664,N_2759,N_2084);
xor U3665 (N_3665,N_2219,N_2241);
or U3666 (N_3666,N_2519,N_2628);
nor U3667 (N_3667,N_2713,N_2006);
nand U3668 (N_3668,N_2519,N_2128);
or U3669 (N_3669,N_2056,N_2827);
nand U3670 (N_3670,N_2762,N_2680);
and U3671 (N_3671,N_2524,N_2444);
nor U3672 (N_3672,N_2173,N_2249);
xnor U3673 (N_3673,N_2426,N_2886);
and U3674 (N_3674,N_2320,N_2180);
nand U3675 (N_3675,N_2971,N_2514);
nand U3676 (N_3676,N_2186,N_2264);
and U3677 (N_3677,N_2647,N_2182);
and U3678 (N_3678,N_2020,N_2699);
and U3679 (N_3679,N_2500,N_2530);
and U3680 (N_3680,N_2575,N_2818);
and U3681 (N_3681,N_2845,N_2170);
nor U3682 (N_3682,N_2540,N_2439);
xor U3683 (N_3683,N_2075,N_2093);
nand U3684 (N_3684,N_2604,N_2921);
xnor U3685 (N_3685,N_2592,N_2990);
nand U3686 (N_3686,N_2199,N_2601);
xor U3687 (N_3687,N_2652,N_2542);
xnor U3688 (N_3688,N_2808,N_2186);
xnor U3689 (N_3689,N_2084,N_2613);
nor U3690 (N_3690,N_2145,N_2517);
and U3691 (N_3691,N_2787,N_2725);
xor U3692 (N_3692,N_2777,N_2893);
and U3693 (N_3693,N_2962,N_2351);
and U3694 (N_3694,N_2612,N_2975);
xnor U3695 (N_3695,N_2933,N_2761);
nor U3696 (N_3696,N_2718,N_2106);
or U3697 (N_3697,N_2486,N_2533);
nand U3698 (N_3698,N_2777,N_2056);
xor U3699 (N_3699,N_2296,N_2704);
xor U3700 (N_3700,N_2605,N_2992);
nor U3701 (N_3701,N_2668,N_2408);
xnor U3702 (N_3702,N_2918,N_2542);
nand U3703 (N_3703,N_2117,N_2462);
nand U3704 (N_3704,N_2191,N_2163);
nor U3705 (N_3705,N_2968,N_2048);
and U3706 (N_3706,N_2794,N_2086);
nor U3707 (N_3707,N_2680,N_2534);
and U3708 (N_3708,N_2508,N_2805);
or U3709 (N_3709,N_2770,N_2084);
and U3710 (N_3710,N_2328,N_2511);
or U3711 (N_3711,N_2979,N_2905);
xor U3712 (N_3712,N_2646,N_2027);
xor U3713 (N_3713,N_2786,N_2618);
nand U3714 (N_3714,N_2516,N_2274);
and U3715 (N_3715,N_2140,N_2839);
nor U3716 (N_3716,N_2825,N_2285);
and U3717 (N_3717,N_2438,N_2641);
or U3718 (N_3718,N_2519,N_2943);
xor U3719 (N_3719,N_2037,N_2312);
and U3720 (N_3720,N_2622,N_2081);
nand U3721 (N_3721,N_2081,N_2744);
nand U3722 (N_3722,N_2336,N_2876);
xor U3723 (N_3723,N_2873,N_2786);
nor U3724 (N_3724,N_2256,N_2854);
or U3725 (N_3725,N_2024,N_2737);
xor U3726 (N_3726,N_2130,N_2313);
or U3727 (N_3727,N_2250,N_2005);
or U3728 (N_3728,N_2067,N_2401);
and U3729 (N_3729,N_2530,N_2368);
nand U3730 (N_3730,N_2744,N_2925);
and U3731 (N_3731,N_2289,N_2666);
nor U3732 (N_3732,N_2554,N_2415);
nor U3733 (N_3733,N_2409,N_2768);
xor U3734 (N_3734,N_2535,N_2636);
xnor U3735 (N_3735,N_2779,N_2014);
or U3736 (N_3736,N_2521,N_2177);
or U3737 (N_3737,N_2890,N_2839);
or U3738 (N_3738,N_2524,N_2146);
and U3739 (N_3739,N_2659,N_2599);
xnor U3740 (N_3740,N_2914,N_2412);
or U3741 (N_3741,N_2494,N_2785);
or U3742 (N_3742,N_2539,N_2041);
and U3743 (N_3743,N_2398,N_2439);
or U3744 (N_3744,N_2491,N_2603);
and U3745 (N_3745,N_2949,N_2686);
and U3746 (N_3746,N_2028,N_2667);
xnor U3747 (N_3747,N_2651,N_2954);
nor U3748 (N_3748,N_2758,N_2475);
nand U3749 (N_3749,N_2207,N_2767);
nand U3750 (N_3750,N_2339,N_2102);
and U3751 (N_3751,N_2946,N_2670);
nand U3752 (N_3752,N_2464,N_2545);
or U3753 (N_3753,N_2083,N_2361);
or U3754 (N_3754,N_2741,N_2549);
xnor U3755 (N_3755,N_2783,N_2234);
or U3756 (N_3756,N_2387,N_2348);
xnor U3757 (N_3757,N_2838,N_2757);
nor U3758 (N_3758,N_2290,N_2814);
or U3759 (N_3759,N_2382,N_2664);
nand U3760 (N_3760,N_2626,N_2981);
and U3761 (N_3761,N_2845,N_2142);
xor U3762 (N_3762,N_2393,N_2929);
xor U3763 (N_3763,N_2856,N_2414);
or U3764 (N_3764,N_2161,N_2832);
nor U3765 (N_3765,N_2592,N_2757);
nand U3766 (N_3766,N_2349,N_2351);
xor U3767 (N_3767,N_2795,N_2103);
nor U3768 (N_3768,N_2062,N_2848);
xnor U3769 (N_3769,N_2758,N_2823);
nor U3770 (N_3770,N_2562,N_2789);
or U3771 (N_3771,N_2064,N_2164);
and U3772 (N_3772,N_2923,N_2993);
and U3773 (N_3773,N_2178,N_2681);
nand U3774 (N_3774,N_2923,N_2462);
or U3775 (N_3775,N_2384,N_2763);
or U3776 (N_3776,N_2833,N_2014);
xor U3777 (N_3777,N_2086,N_2061);
and U3778 (N_3778,N_2838,N_2362);
xor U3779 (N_3779,N_2355,N_2422);
nand U3780 (N_3780,N_2433,N_2354);
nand U3781 (N_3781,N_2619,N_2730);
and U3782 (N_3782,N_2568,N_2649);
nor U3783 (N_3783,N_2677,N_2584);
nand U3784 (N_3784,N_2133,N_2435);
xor U3785 (N_3785,N_2469,N_2036);
or U3786 (N_3786,N_2110,N_2463);
nor U3787 (N_3787,N_2440,N_2718);
xnor U3788 (N_3788,N_2937,N_2896);
or U3789 (N_3789,N_2924,N_2351);
or U3790 (N_3790,N_2902,N_2781);
nand U3791 (N_3791,N_2750,N_2652);
or U3792 (N_3792,N_2889,N_2332);
xor U3793 (N_3793,N_2236,N_2733);
nand U3794 (N_3794,N_2411,N_2323);
nand U3795 (N_3795,N_2915,N_2818);
and U3796 (N_3796,N_2767,N_2112);
and U3797 (N_3797,N_2221,N_2334);
nand U3798 (N_3798,N_2117,N_2949);
xnor U3799 (N_3799,N_2353,N_2271);
or U3800 (N_3800,N_2164,N_2777);
nand U3801 (N_3801,N_2247,N_2099);
nor U3802 (N_3802,N_2989,N_2917);
xnor U3803 (N_3803,N_2072,N_2894);
nand U3804 (N_3804,N_2291,N_2900);
or U3805 (N_3805,N_2489,N_2142);
nand U3806 (N_3806,N_2553,N_2541);
nand U3807 (N_3807,N_2314,N_2711);
nor U3808 (N_3808,N_2601,N_2896);
nor U3809 (N_3809,N_2597,N_2339);
or U3810 (N_3810,N_2746,N_2436);
or U3811 (N_3811,N_2805,N_2609);
nand U3812 (N_3812,N_2614,N_2924);
and U3813 (N_3813,N_2757,N_2654);
nor U3814 (N_3814,N_2773,N_2830);
xor U3815 (N_3815,N_2551,N_2617);
and U3816 (N_3816,N_2430,N_2924);
nor U3817 (N_3817,N_2392,N_2766);
or U3818 (N_3818,N_2676,N_2858);
and U3819 (N_3819,N_2751,N_2667);
xnor U3820 (N_3820,N_2499,N_2413);
and U3821 (N_3821,N_2250,N_2955);
nor U3822 (N_3822,N_2843,N_2122);
nor U3823 (N_3823,N_2796,N_2465);
and U3824 (N_3824,N_2433,N_2111);
or U3825 (N_3825,N_2120,N_2456);
and U3826 (N_3826,N_2685,N_2393);
or U3827 (N_3827,N_2010,N_2721);
xnor U3828 (N_3828,N_2968,N_2549);
nand U3829 (N_3829,N_2676,N_2937);
and U3830 (N_3830,N_2106,N_2611);
and U3831 (N_3831,N_2158,N_2770);
or U3832 (N_3832,N_2143,N_2279);
xor U3833 (N_3833,N_2452,N_2129);
xor U3834 (N_3834,N_2784,N_2870);
nor U3835 (N_3835,N_2924,N_2112);
xnor U3836 (N_3836,N_2453,N_2902);
xor U3837 (N_3837,N_2419,N_2528);
and U3838 (N_3838,N_2530,N_2213);
nand U3839 (N_3839,N_2635,N_2419);
or U3840 (N_3840,N_2640,N_2582);
or U3841 (N_3841,N_2772,N_2974);
xnor U3842 (N_3842,N_2778,N_2869);
or U3843 (N_3843,N_2711,N_2464);
nand U3844 (N_3844,N_2378,N_2664);
nor U3845 (N_3845,N_2866,N_2120);
and U3846 (N_3846,N_2536,N_2293);
nand U3847 (N_3847,N_2988,N_2721);
and U3848 (N_3848,N_2012,N_2318);
nor U3849 (N_3849,N_2470,N_2897);
nand U3850 (N_3850,N_2235,N_2412);
nand U3851 (N_3851,N_2803,N_2425);
nand U3852 (N_3852,N_2545,N_2343);
xnor U3853 (N_3853,N_2293,N_2981);
or U3854 (N_3854,N_2946,N_2118);
and U3855 (N_3855,N_2165,N_2108);
xor U3856 (N_3856,N_2980,N_2424);
or U3857 (N_3857,N_2190,N_2339);
xnor U3858 (N_3858,N_2488,N_2339);
and U3859 (N_3859,N_2450,N_2359);
nor U3860 (N_3860,N_2982,N_2891);
nand U3861 (N_3861,N_2657,N_2442);
and U3862 (N_3862,N_2090,N_2486);
nor U3863 (N_3863,N_2349,N_2745);
and U3864 (N_3864,N_2326,N_2586);
or U3865 (N_3865,N_2980,N_2136);
xor U3866 (N_3866,N_2988,N_2524);
or U3867 (N_3867,N_2456,N_2782);
nand U3868 (N_3868,N_2175,N_2613);
xor U3869 (N_3869,N_2124,N_2485);
or U3870 (N_3870,N_2279,N_2385);
or U3871 (N_3871,N_2527,N_2812);
nand U3872 (N_3872,N_2888,N_2934);
nor U3873 (N_3873,N_2582,N_2759);
nor U3874 (N_3874,N_2993,N_2171);
xor U3875 (N_3875,N_2969,N_2994);
or U3876 (N_3876,N_2919,N_2169);
or U3877 (N_3877,N_2877,N_2327);
nor U3878 (N_3878,N_2084,N_2414);
nand U3879 (N_3879,N_2787,N_2585);
or U3880 (N_3880,N_2485,N_2438);
nand U3881 (N_3881,N_2920,N_2272);
or U3882 (N_3882,N_2323,N_2034);
and U3883 (N_3883,N_2720,N_2571);
and U3884 (N_3884,N_2587,N_2928);
or U3885 (N_3885,N_2578,N_2417);
and U3886 (N_3886,N_2823,N_2169);
xnor U3887 (N_3887,N_2669,N_2934);
xnor U3888 (N_3888,N_2764,N_2318);
nor U3889 (N_3889,N_2919,N_2297);
or U3890 (N_3890,N_2460,N_2726);
nand U3891 (N_3891,N_2462,N_2904);
nand U3892 (N_3892,N_2714,N_2080);
nor U3893 (N_3893,N_2189,N_2610);
nand U3894 (N_3894,N_2306,N_2007);
or U3895 (N_3895,N_2764,N_2547);
or U3896 (N_3896,N_2342,N_2023);
nand U3897 (N_3897,N_2522,N_2877);
nor U3898 (N_3898,N_2699,N_2949);
nor U3899 (N_3899,N_2144,N_2394);
nand U3900 (N_3900,N_2113,N_2857);
nor U3901 (N_3901,N_2148,N_2145);
nor U3902 (N_3902,N_2260,N_2334);
or U3903 (N_3903,N_2952,N_2004);
and U3904 (N_3904,N_2914,N_2923);
and U3905 (N_3905,N_2430,N_2110);
nor U3906 (N_3906,N_2809,N_2882);
and U3907 (N_3907,N_2917,N_2698);
or U3908 (N_3908,N_2284,N_2404);
xnor U3909 (N_3909,N_2486,N_2482);
nor U3910 (N_3910,N_2768,N_2460);
nand U3911 (N_3911,N_2626,N_2974);
or U3912 (N_3912,N_2723,N_2871);
xor U3913 (N_3913,N_2716,N_2412);
or U3914 (N_3914,N_2230,N_2688);
or U3915 (N_3915,N_2950,N_2143);
xor U3916 (N_3916,N_2077,N_2355);
and U3917 (N_3917,N_2133,N_2966);
xnor U3918 (N_3918,N_2221,N_2224);
xor U3919 (N_3919,N_2062,N_2614);
and U3920 (N_3920,N_2744,N_2236);
and U3921 (N_3921,N_2208,N_2225);
nand U3922 (N_3922,N_2784,N_2679);
and U3923 (N_3923,N_2189,N_2513);
xor U3924 (N_3924,N_2914,N_2017);
or U3925 (N_3925,N_2295,N_2521);
xor U3926 (N_3926,N_2048,N_2722);
and U3927 (N_3927,N_2796,N_2553);
nand U3928 (N_3928,N_2523,N_2454);
or U3929 (N_3929,N_2385,N_2522);
nand U3930 (N_3930,N_2374,N_2456);
and U3931 (N_3931,N_2468,N_2821);
or U3932 (N_3932,N_2823,N_2230);
nand U3933 (N_3933,N_2342,N_2159);
and U3934 (N_3934,N_2519,N_2169);
xor U3935 (N_3935,N_2183,N_2814);
or U3936 (N_3936,N_2270,N_2108);
xnor U3937 (N_3937,N_2971,N_2619);
nand U3938 (N_3938,N_2770,N_2582);
and U3939 (N_3939,N_2254,N_2045);
xor U3940 (N_3940,N_2771,N_2401);
xnor U3941 (N_3941,N_2451,N_2755);
nand U3942 (N_3942,N_2719,N_2022);
xnor U3943 (N_3943,N_2733,N_2511);
nand U3944 (N_3944,N_2607,N_2001);
and U3945 (N_3945,N_2052,N_2398);
nor U3946 (N_3946,N_2099,N_2233);
and U3947 (N_3947,N_2423,N_2105);
nand U3948 (N_3948,N_2119,N_2912);
nor U3949 (N_3949,N_2136,N_2701);
or U3950 (N_3950,N_2842,N_2916);
nand U3951 (N_3951,N_2960,N_2195);
and U3952 (N_3952,N_2822,N_2969);
nand U3953 (N_3953,N_2235,N_2943);
nor U3954 (N_3954,N_2447,N_2436);
nor U3955 (N_3955,N_2387,N_2325);
nor U3956 (N_3956,N_2256,N_2045);
xor U3957 (N_3957,N_2988,N_2248);
or U3958 (N_3958,N_2541,N_2884);
or U3959 (N_3959,N_2882,N_2685);
nor U3960 (N_3960,N_2816,N_2454);
nor U3961 (N_3961,N_2762,N_2027);
nand U3962 (N_3962,N_2668,N_2514);
nand U3963 (N_3963,N_2399,N_2712);
and U3964 (N_3964,N_2669,N_2518);
nand U3965 (N_3965,N_2950,N_2132);
or U3966 (N_3966,N_2674,N_2424);
and U3967 (N_3967,N_2419,N_2911);
and U3968 (N_3968,N_2804,N_2380);
or U3969 (N_3969,N_2305,N_2717);
and U3970 (N_3970,N_2289,N_2657);
nand U3971 (N_3971,N_2892,N_2608);
xor U3972 (N_3972,N_2718,N_2988);
or U3973 (N_3973,N_2235,N_2705);
and U3974 (N_3974,N_2395,N_2005);
or U3975 (N_3975,N_2552,N_2123);
and U3976 (N_3976,N_2525,N_2991);
or U3977 (N_3977,N_2784,N_2017);
nor U3978 (N_3978,N_2266,N_2905);
or U3979 (N_3979,N_2265,N_2165);
and U3980 (N_3980,N_2833,N_2938);
xor U3981 (N_3981,N_2727,N_2921);
nand U3982 (N_3982,N_2118,N_2319);
or U3983 (N_3983,N_2455,N_2749);
xor U3984 (N_3984,N_2419,N_2592);
nand U3985 (N_3985,N_2475,N_2550);
nor U3986 (N_3986,N_2273,N_2053);
xor U3987 (N_3987,N_2254,N_2606);
nand U3988 (N_3988,N_2919,N_2726);
xor U3989 (N_3989,N_2031,N_2007);
and U3990 (N_3990,N_2518,N_2787);
or U3991 (N_3991,N_2582,N_2409);
or U3992 (N_3992,N_2029,N_2006);
xor U3993 (N_3993,N_2982,N_2753);
or U3994 (N_3994,N_2120,N_2327);
nand U3995 (N_3995,N_2203,N_2606);
or U3996 (N_3996,N_2896,N_2638);
nand U3997 (N_3997,N_2789,N_2532);
nand U3998 (N_3998,N_2514,N_2577);
or U3999 (N_3999,N_2597,N_2111);
and U4000 (N_4000,N_3613,N_3276);
xnor U4001 (N_4001,N_3031,N_3505);
or U4002 (N_4002,N_3644,N_3479);
nor U4003 (N_4003,N_3730,N_3658);
nor U4004 (N_4004,N_3928,N_3709);
or U4005 (N_4005,N_3669,N_3428);
nand U4006 (N_4006,N_3225,N_3786);
or U4007 (N_4007,N_3553,N_3596);
or U4008 (N_4008,N_3676,N_3387);
nand U4009 (N_4009,N_3421,N_3643);
nand U4010 (N_4010,N_3010,N_3747);
xor U4011 (N_4011,N_3180,N_3196);
or U4012 (N_4012,N_3626,N_3967);
xor U4013 (N_4013,N_3798,N_3602);
and U4014 (N_4014,N_3329,N_3558);
nand U4015 (N_4015,N_3344,N_3272);
and U4016 (N_4016,N_3172,N_3406);
and U4017 (N_4017,N_3788,N_3131);
xor U4018 (N_4018,N_3695,N_3525);
nor U4019 (N_4019,N_3774,N_3229);
and U4020 (N_4020,N_3544,N_3909);
or U4021 (N_4021,N_3463,N_3023);
xor U4022 (N_4022,N_3865,N_3480);
xor U4023 (N_4023,N_3609,N_3371);
nor U4024 (N_4024,N_3866,N_3187);
nand U4025 (N_4025,N_3870,N_3726);
or U4026 (N_4026,N_3426,N_3762);
or U4027 (N_4027,N_3794,N_3259);
or U4028 (N_4028,N_3815,N_3791);
xnor U4029 (N_4029,N_3929,N_3179);
or U4030 (N_4030,N_3482,N_3130);
and U4031 (N_4031,N_3470,N_3099);
and U4032 (N_4032,N_3852,N_3649);
nand U4033 (N_4033,N_3170,N_3316);
nand U4034 (N_4034,N_3917,N_3535);
nand U4035 (N_4035,N_3156,N_3921);
nand U4036 (N_4036,N_3279,N_3230);
and U4037 (N_4037,N_3337,N_3955);
nand U4038 (N_4038,N_3696,N_3026);
nand U4039 (N_4039,N_3627,N_3390);
xor U4040 (N_4040,N_3030,N_3656);
nor U4041 (N_4041,N_3019,N_3171);
nor U4042 (N_4042,N_3894,N_3440);
nor U4043 (N_4043,N_3902,N_3206);
and U4044 (N_4044,N_3410,N_3261);
nor U4045 (N_4045,N_3855,N_3098);
and U4046 (N_4046,N_3391,N_3783);
or U4047 (N_4047,N_3085,N_3930);
and U4048 (N_4048,N_3255,N_3615);
nand U4049 (N_4049,N_3409,N_3300);
or U4050 (N_4050,N_3880,N_3045);
nand U4051 (N_4051,N_3516,N_3086);
and U4052 (N_4052,N_3503,N_3598);
nand U4053 (N_4053,N_3400,N_3079);
xor U4054 (N_4054,N_3799,N_3373);
or U4055 (N_4055,N_3041,N_3741);
xor U4056 (N_4056,N_3071,N_3446);
nand U4057 (N_4057,N_3096,N_3608);
nand U4058 (N_4058,N_3322,N_3563);
nor U4059 (N_4059,N_3236,N_3435);
nand U4060 (N_4060,N_3612,N_3139);
xnor U4061 (N_4061,N_3439,N_3000);
xor U4062 (N_4062,N_3106,N_3304);
and U4063 (N_4063,N_3281,N_3205);
nand U4064 (N_4064,N_3490,N_3862);
or U4065 (N_4065,N_3018,N_3780);
or U4066 (N_4066,N_3804,N_3665);
or U4067 (N_4067,N_3853,N_3933);
nor U4068 (N_4068,N_3244,N_3605);
nor U4069 (N_4069,N_3012,N_3222);
nor U4070 (N_4070,N_3534,N_3924);
nor U4071 (N_4071,N_3966,N_3506);
xnor U4072 (N_4072,N_3364,N_3825);
xor U4073 (N_4073,N_3444,N_3215);
nand U4074 (N_4074,N_3266,N_3290);
nor U4075 (N_4075,N_3867,N_3270);
xnor U4076 (N_4076,N_3303,N_3500);
xnor U4077 (N_4077,N_3177,N_3168);
and U4078 (N_4078,N_3744,N_3820);
or U4079 (N_4079,N_3745,N_3722);
nor U4080 (N_4080,N_3581,N_3697);
xor U4081 (N_4081,N_3403,N_3640);
xor U4082 (N_4082,N_3668,N_3580);
and U4083 (N_4083,N_3264,N_3631);
or U4084 (N_4084,N_3424,N_3953);
and U4085 (N_4085,N_3739,N_3672);
or U4086 (N_4086,N_3822,N_3884);
and U4087 (N_4087,N_3007,N_3311);
nand U4088 (N_4088,N_3477,N_3349);
xnor U4089 (N_4089,N_3105,N_3671);
nand U4090 (N_4090,N_3190,N_3746);
nand U4091 (N_4091,N_3552,N_3734);
nand U4092 (N_4092,N_3578,N_3389);
and U4093 (N_4093,N_3429,N_3195);
nand U4094 (N_4094,N_3214,N_3160);
and U4095 (N_4095,N_3358,N_3607);
xor U4096 (N_4096,N_3343,N_3081);
and U4097 (N_4097,N_3194,N_3978);
and U4098 (N_4098,N_3451,N_3020);
and U4099 (N_4099,N_3869,N_3724);
xnor U4100 (N_4100,N_3134,N_3785);
xnor U4101 (N_4101,N_3268,N_3413);
xnor U4102 (N_4102,N_3845,N_3473);
nor U4103 (N_4103,N_3981,N_3011);
nor U4104 (N_4104,N_3748,N_3811);
nand U4105 (N_4105,N_3795,N_3976);
or U4106 (N_4106,N_3650,N_3342);
xnor U4107 (N_4107,N_3245,N_3033);
and U4108 (N_4108,N_3842,N_3934);
and U4109 (N_4109,N_3393,N_3646);
xor U4110 (N_4110,N_3634,N_3637);
nor U4111 (N_4111,N_3806,N_3948);
nor U4112 (N_4112,N_3996,N_3285);
nor U4113 (N_4113,N_3919,N_3595);
or U4114 (N_4114,N_3882,N_3629);
nor U4115 (N_4115,N_3569,N_3227);
nor U4116 (N_4116,N_3495,N_3496);
and U4117 (N_4117,N_3143,N_3936);
or U4118 (N_4118,N_3474,N_3169);
nor U4119 (N_4119,N_3199,N_3904);
nand U4120 (N_4120,N_3843,N_3462);
xor U4121 (N_4121,N_3913,N_3947);
and U4122 (N_4122,N_3049,N_3557);
and U4123 (N_4123,N_3993,N_3887);
xnor U4124 (N_4124,N_3567,N_3088);
and U4125 (N_4125,N_3336,N_3540);
nor U4126 (N_4126,N_3465,N_3386);
nand U4127 (N_4127,N_3392,N_3009);
nor U4128 (N_4128,N_3528,N_3568);
and U4129 (N_4129,N_3127,N_3326);
and U4130 (N_4130,N_3959,N_3140);
nor U4131 (N_4131,N_3241,N_3193);
or U4132 (N_4132,N_3353,N_3767);
nand U4133 (N_4133,N_3221,N_3778);
and U4134 (N_4134,N_3454,N_3813);
nor U4135 (N_4135,N_3911,N_3588);
xor U4136 (N_4136,N_3514,N_3830);
or U4137 (N_4137,N_3164,N_3619);
nand U4138 (N_4138,N_3827,N_3548);
or U4139 (N_4139,N_3114,N_3128);
nor U4140 (N_4140,N_3135,N_3828);
nand U4141 (N_4141,N_3625,N_3498);
or U4142 (N_4142,N_3162,N_3069);
and U4143 (N_4143,N_3287,N_3059);
or U4144 (N_4144,N_3448,N_3362);
nor U4145 (N_4145,N_3513,N_3365);
and U4146 (N_4146,N_3814,N_3301);
or U4147 (N_4147,N_3916,N_3288);
xnor U4148 (N_4148,N_3152,N_3562);
and U4149 (N_4149,N_3754,N_3396);
or U4150 (N_4150,N_3111,N_3136);
and U4151 (N_4151,N_3103,N_3632);
xor U4152 (N_4152,N_3591,N_3989);
and U4153 (N_4153,N_3801,N_3072);
xnor U4154 (N_4154,N_3313,N_3425);
nor U4155 (N_4155,N_3385,N_3971);
and U4156 (N_4156,N_3520,N_3308);
or U4157 (N_4157,N_3467,N_3551);
xor U4158 (N_4158,N_3898,N_3312);
xnor U4159 (N_4159,N_3704,N_3397);
xnor U4160 (N_4160,N_3053,N_3555);
nand U4161 (N_4161,N_3095,N_3994);
nor U4162 (N_4162,N_3937,N_3986);
nand U4163 (N_4163,N_3176,N_3239);
or U4164 (N_4164,N_3310,N_3620);
xnor U4165 (N_4165,N_3687,N_3566);
or U4166 (N_4166,N_3398,N_3142);
nor U4167 (N_4167,N_3027,N_3345);
nand U4168 (N_4168,N_3459,N_3104);
and U4169 (N_4169,N_3146,N_3542);
nand U4170 (N_4170,N_3823,N_3024);
nor U4171 (N_4171,N_3368,N_3906);
or U4172 (N_4172,N_3384,N_3715);
and U4173 (N_4173,N_3363,N_3122);
and U4174 (N_4174,N_3129,N_3335);
nor U4175 (N_4175,N_3857,N_3893);
xor U4176 (N_4176,N_3892,N_3464);
xor U4177 (N_4177,N_3903,N_3987);
and U4178 (N_4178,N_3943,N_3878);
and U4179 (N_4179,N_3547,N_3051);
nand U4180 (N_4180,N_3655,N_3802);
xor U4181 (N_4181,N_3120,N_3938);
nor U4182 (N_4182,N_3835,N_3125);
nor U4183 (N_4183,N_3790,N_3488);
xnor U4184 (N_4184,N_3653,N_3037);
and U4185 (N_4185,N_3493,N_3163);
and U4186 (N_4186,N_3145,N_3523);
xor U4187 (N_4187,N_3048,N_3016);
nand U4188 (N_4188,N_3183,N_3325);
or U4189 (N_4189,N_3109,N_3900);
xor U4190 (N_4190,N_3610,N_3394);
nand U4191 (N_4191,N_3367,N_3022);
nor U4192 (N_4192,N_3659,N_3831);
or U4193 (N_4193,N_3876,N_3121);
nor U4194 (N_4194,N_3559,N_3750);
and U4195 (N_4195,N_3211,N_3881);
xnor U4196 (N_4196,N_3597,N_3327);
nand U4197 (N_4197,N_3777,N_3705);
xor U4198 (N_4198,N_3849,N_3203);
or U4199 (N_4199,N_3294,N_3237);
nand U4200 (N_4200,N_3379,N_3050);
and U4201 (N_4201,N_3035,N_3945);
nand U4202 (N_4202,N_3560,N_3915);
nor U4203 (N_4203,N_3357,N_3437);
xnor U4204 (N_4204,N_3861,N_3623);
or U4205 (N_4205,N_3124,N_3711);
nand U4206 (N_4206,N_3963,N_3859);
nand U4207 (N_4207,N_3652,N_3216);
nand U4208 (N_4208,N_3723,N_3789);
xnor U4209 (N_4209,N_3998,N_3433);
or U4210 (N_4210,N_3995,N_3481);
nand U4211 (N_4211,N_3974,N_3541);
or U4212 (N_4212,N_3960,N_3115);
or U4213 (N_4213,N_3592,N_3784);
nor U4214 (N_4214,N_3965,N_3510);
xor U4215 (N_4215,N_3113,N_3810);
nand U4216 (N_4216,N_3599,N_3854);
xnor U4217 (N_4217,N_3296,N_3263);
or U4218 (N_4218,N_3434,N_3184);
nor U4219 (N_4219,N_3648,N_3518);
nand U4220 (N_4220,N_3292,N_3044);
or U4221 (N_4221,N_3851,N_3250);
xnor U4222 (N_4222,N_3604,N_3519);
nor U4223 (N_4223,N_3380,N_3132);
nand U4224 (N_4224,N_3769,N_3155);
and U4225 (N_4225,N_3351,N_3422);
xor U4226 (N_4226,N_3200,N_3491);
or U4227 (N_4227,N_3333,N_3949);
xnor U4228 (N_4228,N_3058,N_3070);
xor U4229 (N_4229,N_3262,N_3014);
xnor U4230 (N_4230,N_3240,N_3847);
nor U4231 (N_4231,N_3013,N_3060);
or U4232 (N_4232,N_3021,N_3117);
and U4233 (N_4233,N_3015,N_3720);
and U4234 (N_4234,N_3679,N_3522);
nand U4235 (N_4235,N_3116,N_3699);
and U4236 (N_4236,N_3382,N_3402);
nand U4237 (N_4237,N_3441,N_3207);
or U4238 (N_4238,N_3372,N_3545);
nand U4239 (N_4239,N_3968,N_3816);
nand U4240 (N_4240,N_3317,N_3209);
xnor U4241 (N_4241,N_3661,N_3800);
or U4242 (N_4242,N_3133,N_3793);
xnor U4243 (N_4243,N_3191,N_3756);
nor U4244 (N_4244,N_3639,N_3895);
nand U4245 (N_4245,N_3512,N_3850);
and U4246 (N_4246,N_3803,N_3299);
nor U4247 (N_4247,N_3297,N_3611);
and U4248 (N_4248,N_3923,N_3305);
and U4249 (N_4249,N_3295,N_3589);
xor U4250 (N_4250,N_3219,N_3068);
or U4251 (N_4251,N_3885,N_3277);
nor U4252 (N_4252,N_3166,N_3185);
xnor U4253 (N_4253,N_3347,N_3992);
and U4254 (N_4254,N_3925,N_3808);
xor U4255 (N_4255,N_3234,N_3408);
or U4256 (N_4256,N_3118,N_3453);
nor U4257 (N_4257,N_3621,N_3167);
or U4258 (N_4258,N_3549,N_3863);
nand U4259 (N_4259,N_3990,N_3126);
or U4260 (N_4260,N_3267,N_3759);
nand U4261 (N_4261,N_3727,N_3583);
or U4262 (N_4262,N_3931,N_3872);
nand U4263 (N_4263,N_3642,N_3712);
nand U4264 (N_4264,N_3100,N_3283);
xnor U4265 (N_4265,N_3405,N_3663);
xnor U4266 (N_4266,N_3097,N_3501);
or U4267 (N_4267,N_3680,N_3543);
and U4268 (N_4268,N_3159,N_3997);
xnor U4269 (N_4269,N_3376,N_3587);
nand U4270 (N_4270,N_3841,N_3274);
or U4271 (N_4271,N_3614,N_3617);
nor U4272 (N_4272,N_3291,N_3460);
nor U4273 (N_4273,N_3381,N_3834);
and U4274 (N_4274,N_3694,N_3565);
xnor U4275 (N_4275,N_3973,N_3515);
nor U4276 (N_4276,N_3550,N_3075);
and U4277 (N_4277,N_3575,N_3985);
nor U4278 (N_4278,N_3980,N_3082);
and U4279 (N_4279,N_3210,N_3404);
and U4280 (N_4280,N_3701,N_3314);
xnor U4281 (N_4281,N_3982,N_3243);
nor U4282 (N_4282,N_3707,N_3174);
or U4283 (N_4283,N_3654,N_3431);
or U4284 (N_4284,N_3603,N_3377);
or U4285 (N_4285,N_3531,N_3779);
nor U4286 (N_4286,N_3584,N_3138);
xnor U4287 (N_4287,N_3698,N_3201);
nor U4288 (N_4288,N_3089,N_3961);
nand U4289 (N_4289,N_3006,N_3039);
nand U4290 (N_4290,N_3278,N_3579);
and U4291 (N_4291,N_3690,N_3868);
or U4292 (N_4292,N_3839,N_3606);
or U4293 (N_4293,N_3691,N_3683);
xnor U4294 (N_4294,N_3890,N_3218);
nand U4295 (N_4295,N_3137,N_3817);
nor U4296 (N_4296,N_3703,N_3667);
and U4297 (N_4297,N_3427,N_3323);
or U4298 (N_4298,N_3914,N_3871);
nand U4299 (N_4299,N_3972,N_3689);
or U4300 (N_4300,N_3647,N_3957);
xor U4301 (N_4301,N_3590,N_3782);
nor U4302 (N_4302,N_3054,N_3952);
nor U4303 (N_4303,N_3188,N_3202);
and U4304 (N_4304,N_3476,N_3848);
nor U4305 (N_4305,N_3181,N_3242);
and U4306 (N_4306,N_3083,N_3485);
nand U4307 (N_4307,N_3025,N_3719);
nand U4308 (N_4308,N_3725,N_3066);
nand U4309 (N_4309,N_3950,N_3456);
or U4310 (N_4310,N_3052,N_3554);
xnor U4311 (N_4311,N_3046,N_3772);
and U4312 (N_4312,N_3254,N_3910);
and U4313 (N_4313,N_3484,N_3999);
or U4314 (N_4314,N_3407,N_3061);
or U4315 (N_4315,N_3771,N_3001);
nor U4316 (N_4316,N_3838,N_3332);
nor U4317 (N_4317,N_3067,N_3752);
or U4318 (N_4318,N_3532,N_3042);
nand U4319 (N_4319,N_3213,N_3471);
or U4320 (N_4320,N_3258,N_3899);
and U4321 (N_4321,N_3533,N_3526);
nor U4322 (N_4322,N_3954,N_3684);
xnor U4323 (N_4323,N_3032,N_3511);
and U4324 (N_4324,N_3673,N_3217);
nand U4325 (N_4325,N_3641,N_3766);
nand U4326 (N_4326,N_3888,N_3282);
nor U4327 (N_4327,N_3879,N_3908);
xor U4328 (N_4328,N_3593,N_3572);
nor U4329 (N_4329,N_3093,N_3740);
xnor U4330 (N_4330,N_3905,N_3265);
xnor U4331 (N_4331,N_3805,N_3939);
nand U4332 (N_4332,N_3154,N_3509);
nor U4333 (N_4333,N_3360,N_3414);
xnor U4334 (N_4334,N_3324,N_3348);
nand U4335 (N_4335,N_3101,N_3958);
nor U4336 (N_4336,N_3737,N_3728);
xnor U4337 (N_4337,N_3472,N_3713);
nor U4338 (N_4338,N_3469,N_3530);
nor U4339 (N_4339,N_3664,N_3416);
xor U4340 (N_4340,N_3036,N_3651);
or U4341 (N_4341,N_3173,N_3660);
and U4342 (N_4342,N_3401,N_3877);
and U4343 (N_4343,N_3361,N_3818);
nor U4344 (N_4344,N_3556,N_3529);
nor U4345 (N_4345,N_3757,N_3633);
nand U4346 (N_4346,N_3688,N_3320);
nand U4347 (N_4347,N_3570,N_3729);
and U4348 (N_4348,N_3731,N_3497);
and U4349 (N_4349,N_3977,N_3969);
and U4350 (N_4350,N_3257,N_3461);
and U4351 (N_4351,N_3107,N_3546);
or U4352 (N_4352,N_3883,N_3749);
or U4353 (N_4353,N_3657,N_3860);
and U4354 (N_4354,N_3420,N_3455);
nor U4355 (N_4355,N_3328,N_3927);
nor U4356 (N_4356,N_3920,N_3521);
or U4357 (N_4357,N_3681,N_3432);
xor U4358 (N_4358,N_3445,N_3073);
or U4359 (N_4359,N_3991,N_3375);
nand U4360 (N_4360,N_3685,N_3875);
and U4361 (N_4361,N_3670,N_3412);
nand U4362 (N_4362,N_3824,N_3979);
nand U4363 (N_4363,N_3091,N_3674);
and U4364 (N_4364,N_3844,N_3423);
or U4365 (N_4365,N_3438,N_3430);
or U4366 (N_4366,N_3192,N_3692);
and U4367 (N_4367,N_3944,N_3388);
nand U4368 (N_4368,N_3253,N_3366);
and U4369 (N_4369,N_3912,N_3315);
or U4370 (N_4370,N_3829,N_3302);
or U4371 (N_4371,N_3622,N_3962);
xnor U4372 (N_4372,N_3874,N_3220);
or U4373 (N_4373,N_3507,N_3112);
and U4374 (N_4374,N_3693,N_3760);
and U4375 (N_4375,N_3208,N_3002);
or U4376 (N_4376,N_3186,N_3840);
and U4377 (N_4377,N_3378,N_3354);
or U4378 (N_4378,N_3076,N_3147);
xnor U4379 (N_4379,N_3411,N_3504);
xnor U4380 (N_4380,N_3252,N_3577);
nor U4381 (N_4381,N_3738,N_3307);
nand U4382 (N_4382,N_3341,N_3319);
nor U4383 (N_4383,N_3475,N_3478);
nand U4384 (N_4384,N_3144,N_3812);
or U4385 (N_4385,N_3182,N_3662);
or U4386 (N_4386,N_3466,N_3710);
nor U4387 (N_4387,N_3197,N_3284);
nor U4388 (N_4388,N_3708,N_3228);
nand U4389 (N_4389,N_3821,N_3108);
nand U4390 (N_4390,N_3189,N_3764);
nor U4391 (N_4391,N_3092,N_3340);
nor U4392 (N_4392,N_3256,N_3178);
nand U4393 (N_4393,N_3988,N_3309);
and U4394 (N_4394,N_3527,N_3856);
and U4395 (N_4395,N_3415,N_3119);
or U4396 (N_4396,N_3008,N_3524);
or U4397 (N_4397,N_3247,N_3628);
xnor U4398 (N_4398,N_3537,N_3564);
nand U4399 (N_4399,N_3807,N_3468);
or U4400 (N_4400,N_3864,N_3102);
nand U4401 (N_4401,N_3932,N_3718);
or U4402 (N_4402,N_3280,N_3458);
nor U4403 (N_4403,N_3561,N_3666);
xnor U4404 (N_4404,N_3204,N_3005);
nand U4405 (N_4405,N_3983,N_3034);
nor U4406 (N_4406,N_3330,N_3742);
and U4407 (N_4407,N_3251,N_3055);
nor U4408 (N_4408,N_3078,N_3457);
nor U4409 (N_4409,N_3975,N_3334);
xnor U4410 (N_4410,N_3004,N_3758);
nor U4411 (N_4411,N_3223,N_3418);
nand U4412 (N_4412,N_3056,N_3233);
nand U4413 (N_4413,N_3141,N_3775);
nor U4414 (N_4414,N_3763,N_3436);
nand U4415 (N_4415,N_3003,N_3269);
nand U4416 (N_4416,N_3776,N_3761);
nand U4417 (N_4417,N_3618,N_3574);
and U4418 (N_4418,N_3922,N_3452);
nor U4419 (N_4419,N_3449,N_3355);
or U4420 (N_4420,N_3636,N_3940);
and U4421 (N_4421,N_3736,N_3158);
and U4422 (N_4422,N_3706,N_3832);
or U4423 (N_4423,N_3249,N_3600);
nor U4424 (N_4424,N_3901,N_3094);
nand U4425 (N_4425,N_3946,N_3601);
nand U4426 (N_4426,N_3077,N_3768);
xnor U4427 (N_4427,N_3383,N_3486);
nand U4428 (N_4428,N_3017,N_3374);
or U4429 (N_4429,N_3645,N_3148);
and U4430 (N_4430,N_3781,N_3837);
or U4431 (N_4431,N_3918,N_3175);
xor U4432 (N_4432,N_3029,N_3717);
or U4433 (N_4433,N_3038,N_3338);
and U4434 (N_4434,N_3063,N_3235);
xor U4435 (N_4435,N_3984,N_3212);
and U4436 (N_4436,N_3298,N_3502);
nand U4437 (N_4437,N_3289,N_3492);
xor U4438 (N_4438,N_3062,N_3956);
or U4439 (N_4439,N_3487,N_3755);
nand U4440 (N_4440,N_3926,N_3586);
nand U4441 (N_4441,N_3450,N_3153);
xor U4442 (N_4442,N_3447,N_3321);
or U4443 (N_4443,N_3028,N_3198);
or U4444 (N_4444,N_3087,N_3585);
xnor U4445 (N_4445,N_3260,N_3594);
nand U4446 (N_4446,N_3765,N_3483);
and U4447 (N_4447,N_3395,N_3582);
xnor U4448 (N_4448,N_3677,N_3123);
or U4449 (N_4449,N_3735,N_3224);
xor U4450 (N_4450,N_3797,N_3306);
xnor U4451 (N_4451,N_3369,N_3161);
nor U4452 (N_4452,N_3352,N_3350);
xnor U4453 (N_4453,N_3907,N_3047);
nor U4454 (N_4454,N_3896,N_3616);
xnor U4455 (N_4455,N_3150,N_3346);
xor U4456 (N_4456,N_3682,N_3399);
and U4457 (N_4457,N_3356,N_3151);
nand U4458 (N_4458,N_3165,N_3318);
or U4459 (N_4459,N_3792,N_3941);
nand U4460 (N_4460,N_3043,N_3238);
nand U4461 (N_4461,N_3846,N_3638);
nand U4462 (N_4462,N_3417,N_3273);
and U4463 (N_4463,N_3678,N_3819);
or U4464 (N_4464,N_3074,N_3571);
and U4465 (N_4465,N_3248,N_3576);
nand U4466 (N_4466,N_3833,N_3935);
nor U4467 (N_4467,N_3873,N_3716);
or U4468 (N_4468,N_3494,N_3897);
xor U4469 (N_4469,N_3080,N_3271);
nand U4470 (N_4470,N_3442,N_3787);
xnor U4471 (N_4471,N_3970,N_3796);
and U4472 (N_4472,N_3084,N_3275);
nand U4473 (N_4473,N_3751,N_3370);
xor U4474 (N_4474,N_3246,N_3733);
xor U4475 (N_4475,N_3539,N_3721);
xnor U4476 (N_4476,N_3770,N_3339);
nor U4477 (N_4477,N_3714,N_3624);
and U4478 (N_4478,N_3858,N_3702);
xnor U4479 (N_4479,N_3040,N_3057);
and U4480 (N_4480,N_3286,N_3889);
or U4481 (N_4481,N_3942,N_3489);
nor U4482 (N_4482,N_3753,N_3517);
or U4483 (N_4483,N_3064,N_3090);
xor U4484 (N_4484,N_3686,N_3630);
or U4485 (N_4485,N_3232,N_3536);
or U4486 (N_4486,N_3826,N_3743);
and U4487 (N_4487,N_3499,N_3964);
nor U4488 (N_4488,N_3149,N_3065);
nand U4489 (N_4489,N_3359,N_3675);
xnor U4490 (N_4490,N_3443,N_3951);
or U4491 (N_4491,N_3891,N_3110);
and U4492 (N_4492,N_3157,N_3836);
or U4493 (N_4493,N_3538,N_3231);
nand U4494 (N_4494,N_3226,N_3573);
xor U4495 (N_4495,N_3419,N_3886);
nor U4496 (N_4496,N_3809,N_3732);
xnor U4497 (N_4497,N_3331,N_3635);
nand U4498 (N_4498,N_3700,N_3508);
nor U4499 (N_4499,N_3293,N_3773);
nand U4500 (N_4500,N_3364,N_3381);
nor U4501 (N_4501,N_3021,N_3267);
xnor U4502 (N_4502,N_3554,N_3756);
nand U4503 (N_4503,N_3012,N_3971);
or U4504 (N_4504,N_3697,N_3457);
and U4505 (N_4505,N_3649,N_3267);
or U4506 (N_4506,N_3330,N_3693);
and U4507 (N_4507,N_3830,N_3587);
or U4508 (N_4508,N_3654,N_3645);
or U4509 (N_4509,N_3022,N_3678);
xor U4510 (N_4510,N_3868,N_3791);
and U4511 (N_4511,N_3315,N_3443);
nand U4512 (N_4512,N_3776,N_3974);
and U4513 (N_4513,N_3995,N_3417);
nor U4514 (N_4514,N_3630,N_3648);
and U4515 (N_4515,N_3658,N_3961);
nor U4516 (N_4516,N_3441,N_3695);
nor U4517 (N_4517,N_3825,N_3421);
xnor U4518 (N_4518,N_3229,N_3027);
nand U4519 (N_4519,N_3755,N_3375);
and U4520 (N_4520,N_3172,N_3837);
or U4521 (N_4521,N_3640,N_3834);
xnor U4522 (N_4522,N_3472,N_3402);
xor U4523 (N_4523,N_3732,N_3257);
or U4524 (N_4524,N_3224,N_3929);
nor U4525 (N_4525,N_3067,N_3827);
nor U4526 (N_4526,N_3178,N_3199);
or U4527 (N_4527,N_3969,N_3689);
xor U4528 (N_4528,N_3683,N_3519);
or U4529 (N_4529,N_3774,N_3686);
or U4530 (N_4530,N_3525,N_3985);
nand U4531 (N_4531,N_3214,N_3855);
xnor U4532 (N_4532,N_3086,N_3061);
and U4533 (N_4533,N_3604,N_3223);
and U4534 (N_4534,N_3165,N_3591);
nand U4535 (N_4535,N_3720,N_3545);
and U4536 (N_4536,N_3497,N_3675);
or U4537 (N_4537,N_3984,N_3543);
nand U4538 (N_4538,N_3482,N_3881);
or U4539 (N_4539,N_3921,N_3609);
xnor U4540 (N_4540,N_3604,N_3348);
xor U4541 (N_4541,N_3178,N_3681);
nand U4542 (N_4542,N_3792,N_3843);
nand U4543 (N_4543,N_3266,N_3685);
nor U4544 (N_4544,N_3857,N_3065);
and U4545 (N_4545,N_3917,N_3506);
xor U4546 (N_4546,N_3392,N_3792);
nor U4547 (N_4547,N_3115,N_3027);
nor U4548 (N_4548,N_3949,N_3891);
xor U4549 (N_4549,N_3862,N_3399);
xor U4550 (N_4550,N_3100,N_3711);
nor U4551 (N_4551,N_3153,N_3760);
nand U4552 (N_4552,N_3668,N_3959);
nor U4553 (N_4553,N_3020,N_3921);
and U4554 (N_4554,N_3629,N_3933);
xnor U4555 (N_4555,N_3060,N_3707);
xnor U4556 (N_4556,N_3283,N_3370);
nor U4557 (N_4557,N_3175,N_3627);
xnor U4558 (N_4558,N_3764,N_3875);
nand U4559 (N_4559,N_3423,N_3706);
nand U4560 (N_4560,N_3107,N_3692);
and U4561 (N_4561,N_3779,N_3807);
xnor U4562 (N_4562,N_3202,N_3561);
nor U4563 (N_4563,N_3163,N_3510);
nand U4564 (N_4564,N_3245,N_3873);
nand U4565 (N_4565,N_3498,N_3041);
nand U4566 (N_4566,N_3120,N_3180);
or U4567 (N_4567,N_3446,N_3920);
xnor U4568 (N_4568,N_3284,N_3139);
nand U4569 (N_4569,N_3502,N_3458);
xor U4570 (N_4570,N_3113,N_3945);
nor U4571 (N_4571,N_3996,N_3867);
or U4572 (N_4572,N_3280,N_3603);
nand U4573 (N_4573,N_3444,N_3119);
nor U4574 (N_4574,N_3308,N_3923);
or U4575 (N_4575,N_3018,N_3579);
or U4576 (N_4576,N_3940,N_3356);
and U4577 (N_4577,N_3838,N_3385);
and U4578 (N_4578,N_3201,N_3857);
and U4579 (N_4579,N_3260,N_3513);
nor U4580 (N_4580,N_3928,N_3855);
or U4581 (N_4581,N_3827,N_3280);
nor U4582 (N_4582,N_3955,N_3832);
nor U4583 (N_4583,N_3380,N_3600);
nand U4584 (N_4584,N_3328,N_3893);
or U4585 (N_4585,N_3982,N_3092);
and U4586 (N_4586,N_3736,N_3589);
and U4587 (N_4587,N_3891,N_3314);
and U4588 (N_4588,N_3882,N_3085);
xor U4589 (N_4589,N_3971,N_3634);
xnor U4590 (N_4590,N_3777,N_3277);
or U4591 (N_4591,N_3452,N_3870);
nor U4592 (N_4592,N_3230,N_3590);
xnor U4593 (N_4593,N_3965,N_3767);
or U4594 (N_4594,N_3652,N_3082);
and U4595 (N_4595,N_3752,N_3647);
and U4596 (N_4596,N_3107,N_3269);
nand U4597 (N_4597,N_3131,N_3598);
and U4598 (N_4598,N_3392,N_3621);
nand U4599 (N_4599,N_3035,N_3517);
xor U4600 (N_4600,N_3679,N_3265);
and U4601 (N_4601,N_3124,N_3339);
or U4602 (N_4602,N_3372,N_3530);
xor U4603 (N_4603,N_3725,N_3193);
or U4604 (N_4604,N_3162,N_3001);
xnor U4605 (N_4605,N_3964,N_3514);
or U4606 (N_4606,N_3001,N_3370);
xnor U4607 (N_4607,N_3390,N_3341);
or U4608 (N_4608,N_3783,N_3900);
nand U4609 (N_4609,N_3347,N_3693);
nor U4610 (N_4610,N_3237,N_3043);
or U4611 (N_4611,N_3274,N_3705);
or U4612 (N_4612,N_3357,N_3978);
and U4613 (N_4613,N_3765,N_3833);
or U4614 (N_4614,N_3880,N_3682);
xor U4615 (N_4615,N_3656,N_3068);
nand U4616 (N_4616,N_3789,N_3065);
nand U4617 (N_4617,N_3754,N_3948);
xor U4618 (N_4618,N_3325,N_3667);
nor U4619 (N_4619,N_3421,N_3122);
xnor U4620 (N_4620,N_3118,N_3590);
and U4621 (N_4621,N_3465,N_3060);
nand U4622 (N_4622,N_3810,N_3432);
xor U4623 (N_4623,N_3470,N_3874);
nand U4624 (N_4624,N_3662,N_3716);
or U4625 (N_4625,N_3704,N_3738);
xnor U4626 (N_4626,N_3876,N_3535);
and U4627 (N_4627,N_3266,N_3299);
xnor U4628 (N_4628,N_3461,N_3298);
and U4629 (N_4629,N_3832,N_3769);
and U4630 (N_4630,N_3838,N_3761);
or U4631 (N_4631,N_3324,N_3074);
nand U4632 (N_4632,N_3236,N_3988);
nor U4633 (N_4633,N_3858,N_3641);
and U4634 (N_4634,N_3260,N_3075);
or U4635 (N_4635,N_3000,N_3152);
xnor U4636 (N_4636,N_3755,N_3284);
or U4637 (N_4637,N_3822,N_3536);
and U4638 (N_4638,N_3110,N_3197);
nand U4639 (N_4639,N_3191,N_3930);
and U4640 (N_4640,N_3289,N_3713);
and U4641 (N_4641,N_3313,N_3584);
and U4642 (N_4642,N_3602,N_3368);
or U4643 (N_4643,N_3941,N_3524);
and U4644 (N_4644,N_3337,N_3238);
nor U4645 (N_4645,N_3208,N_3757);
nor U4646 (N_4646,N_3511,N_3691);
nand U4647 (N_4647,N_3099,N_3201);
and U4648 (N_4648,N_3731,N_3207);
and U4649 (N_4649,N_3142,N_3821);
nor U4650 (N_4650,N_3402,N_3792);
or U4651 (N_4651,N_3877,N_3954);
nor U4652 (N_4652,N_3612,N_3526);
nor U4653 (N_4653,N_3917,N_3346);
xnor U4654 (N_4654,N_3545,N_3873);
nor U4655 (N_4655,N_3444,N_3752);
nand U4656 (N_4656,N_3732,N_3433);
or U4657 (N_4657,N_3166,N_3779);
nand U4658 (N_4658,N_3149,N_3162);
or U4659 (N_4659,N_3730,N_3675);
nand U4660 (N_4660,N_3663,N_3566);
nor U4661 (N_4661,N_3281,N_3735);
and U4662 (N_4662,N_3729,N_3107);
and U4663 (N_4663,N_3357,N_3065);
nand U4664 (N_4664,N_3592,N_3263);
and U4665 (N_4665,N_3380,N_3652);
xnor U4666 (N_4666,N_3864,N_3646);
or U4667 (N_4667,N_3660,N_3281);
nor U4668 (N_4668,N_3207,N_3092);
nor U4669 (N_4669,N_3252,N_3519);
xor U4670 (N_4670,N_3757,N_3439);
nor U4671 (N_4671,N_3535,N_3307);
xor U4672 (N_4672,N_3301,N_3917);
xnor U4673 (N_4673,N_3210,N_3974);
nor U4674 (N_4674,N_3500,N_3210);
xnor U4675 (N_4675,N_3494,N_3701);
xor U4676 (N_4676,N_3615,N_3732);
nand U4677 (N_4677,N_3993,N_3816);
nand U4678 (N_4678,N_3149,N_3113);
and U4679 (N_4679,N_3959,N_3260);
xor U4680 (N_4680,N_3734,N_3001);
or U4681 (N_4681,N_3137,N_3341);
xor U4682 (N_4682,N_3999,N_3979);
nand U4683 (N_4683,N_3231,N_3354);
xnor U4684 (N_4684,N_3042,N_3633);
xnor U4685 (N_4685,N_3765,N_3314);
nand U4686 (N_4686,N_3249,N_3740);
nand U4687 (N_4687,N_3819,N_3817);
or U4688 (N_4688,N_3397,N_3804);
xnor U4689 (N_4689,N_3255,N_3862);
xor U4690 (N_4690,N_3479,N_3666);
and U4691 (N_4691,N_3810,N_3635);
and U4692 (N_4692,N_3572,N_3111);
or U4693 (N_4693,N_3853,N_3903);
nor U4694 (N_4694,N_3085,N_3858);
xor U4695 (N_4695,N_3424,N_3915);
or U4696 (N_4696,N_3558,N_3339);
and U4697 (N_4697,N_3337,N_3593);
xor U4698 (N_4698,N_3500,N_3063);
nor U4699 (N_4699,N_3089,N_3524);
nor U4700 (N_4700,N_3894,N_3016);
and U4701 (N_4701,N_3351,N_3263);
nand U4702 (N_4702,N_3729,N_3086);
and U4703 (N_4703,N_3575,N_3384);
and U4704 (N_4704,N_3895,N_3960);
xnor U4705 (N_4705,N_3294,N_3901);
or U4706 (N_4706,N_3050,N_3211);
nor U4707 (N_4707,N_3850,N_3293);
xor U4708 (N_4708,N_3019,N_3937);
and U4709 (N_4709,N_3124,N_3720);
or U4710 (N_4710,N_3717,N_3133);
and U4711 (N_4711,N_3200,N_3232);
xnor U4712 (N_4712,N_3582,N_3908);
and U4713 (N_4713,N_3414,N_3875);
and U4714 (N_4714,N_3860,N_3506);
nand U4715 (N_4715,N_3945,N_3422);
nand U4716 (N_4716,N_3604,N_3871);
nor U4717 (N_4717,N_3807,N_3017);
xor U4718 (N_4718,N_3543,N_3306);
nor U4719 (N_4719,N_3147,N_3358);
and U4720 (N_4720,N_3677,N_3492);
nor U4721 (N_4721,N_3324,N_3768);
or U4722 (N_4722,N_3425,N_3192);
nand U4723 (N_4723,N_3176,N_3796);
xnor U4724 (N_4724,N_3979,N_3300);
or U4725 (N_4725,N_3703,N_3097);
or U4726 (N_4726,N_3646,N_3500);
nor U4727 (N_4727,N_3989,N_3231);
and U4728 (N_4728,N_3649,N_3910);
nor U4729 (N_4729,N_3975,N_3790);
and U4730 (N_4730,N_3208,N_3589);
and U4731 (N_4731,N_3219,N_3530);
nor U4732 (N_4732,N_3139,N_3799);
xor U4733 (N_4733,N_3942,N_3742);
and U4734 (N_4734,N_3685,N_3779);
and U4735 (N_4735,N_3825,N_3261);
and U4736 (N_4736,N_3134,N_3705);
nand U4737 (N_4737,N_3234,N_3341);
or U4738 (N_4738,N_3058,N_3450);
and U4739 (N_4739,N_3167,N_3610);
and U4740 (N_4740,N_3769,N_3204);
nand U4741 (N_4741,N_3297,N_3853);
nor U4742 (N_4742,N_3920,N_3739);
nand U4743 (N_4743,N_3192,N_3888);
xnor U4744 (N_4744,N_3824,N_3330);
nor U4745 (N_4745,N_3297,N_3330);
or U4746 (N_4746,N_3109,N_3486);
and U4747 (N_4747,N_3343,N_3946);
nand U4748 (N_4748,N_3128,N_3186);
nor U4749 (N_4749,N_3964,N_3149);
and U4750 (N_4750,N_3963,N_3515);
nand U4751 (N_4751,N_3298,N_3286);
nor U4752 (N_4752,N_3322,N_3747);
and U4753 (N_4753,N_3895,N_3498);
or U4754 (N_4754,N_3968,N_3138);
nand U4755 (N_4755,N_3717,N_3596);
nand U4756 (N_4756,N_3834,N_3326);
or U4757 (N_4757,N_3338,N_3341);
nor U4758 (N_4758,N_3429,N_3638);
and U4759 (N_4759,N_3438,N_3594);
nor U4760 (N_4760,N_3673,N_3708);
xnor U4761 (N_4761,N_3752,N_3874);
and U4762 (N_4762,N_3308,N_3825);
nand U4763 (N_4763,N_3611,N_3740);
or U4764 (N_4764,N_3526,N_3928);
nand U4765 (N_4765,N_3349,N_3944);
xor U4766 (N_4766,N_3437,N_3717);
xnor U4767 (N_4767,N_3971,N_3762);
and U4768 (N_4768,N_3114,N_3010);
nor U4769 (N_4769,N_3539,N_3839);
xnor U4770 (N_4770,N_3820,N_3067);
xnor U4771 (N_4771,N_3785,N_3584);
nand U4772 (N_4772,N_3624,N_3311);
nor U4773 (N_4773,N_3825,N_3243);
nand U4774 (N_4774,N_3275,N_3755);
nand U4775 (N_4775,N_3209,N_3467);
xor U4776 (N_4776,N_3016,N_3773);
xnor U4777 (N_4777,N_3829,N_3105);
or U4778 (N_4778,N_3184,N_3812);
xor U4779 (N_4779,N_3585,N_3111);
nand U4780 (N_4780,N_3055,N_3644);
nor U4781 (N_4781,N_3000,N_3316);
nor U4782 (N_4782,N_3144,N_3180);
and U4783 (N_4783,N_3125,N_3872);
nor U4784 (N_4784,N_3153,N_3118);
or U4785 (N_4785,N_3838,N_3871);
and U4786 (N_4786,N_3634,N_3454);
or U4787 (N_4787,N_3756,N_3170);
and U4788 (N_4788,N_3157,N_3979);
and U4789 (N_4789,N_3483,N_3409);
nand U4790 (N_4790,N_3371,N_3671);
or U4791 (N_4791,N_3820,N_3360);
nand U4792 (N_4792,N_3620,N_3082);
or U4793 (N_4793,N_3995,N_3404);
and U4794 (N_4794,N_3968,N_3723);
xnor U4795 (N_4795,N_3497,N_3444);
and U4796 (N_4796,N_3192,N_3691);
nor U4797 (N_4797,N_3936,N_3190);
or U4798 (N_4798,N_3865,N_3132);
nor U4799 (N_4799,N_3351,N_3250);
nor U4800 (N_4800,N_3591,N_3854);
nor U4801 (N_4801,N_3765,N_3104);
nor U4802 (N_4802,N_3912,N_3152);
nor U4803 (N_4803,N_3535,N_3063);
nand U4804 (N_4804,N_3780,N_3899);
xnor U4805 (N_4805,N_3614,N_3647);
xor U4806 (N_4806,N_3356,N_3427);
nor U4807 (N_4807,N_3401,N_3625);
nor U4808 (N_4808,N_3969,N_3842);
and U4809 (N_4809,N_3535,N_3316);
nand U4810 (N_4810,N_3482,N_3552);
nor U4811 (N_4811,N_3748,N_3046);
or U4812 (N_4812,N_3869,N_3921);
nand U4813 (N_4813,N_3322,N_3534);
nand U4814 (N_4814,N_3458,N_3915);
nor U4815 (N_4815,N_3291,N_3514);
and U4816 (N_4816,N_3627,N_3032);
and U4817 (N_4817,N_3763,N_3977);
nor U4818 (N_4818,N_3797,N_3798);
and U4819 (N_4819,N_3384,N_3604);
nor U4820 (N_4820,N_3608,N_3598);
nand U4821 (N_4821,N_3007,N_3410);
and U4822 (N_4822,N_3223,N_3587);
or U4823 (N_4823,N_3359,N_3942);
or U4824 (N_4824,N_3077,N_3872);
nand U4825 (N_4825,N_3521,N_3566);
or U4826 (N_4826,N_3065,N_3196);
xnor U4827 (N_4827,N_3284,N_3208);
nor U4828 (N_4828,N_3271,N_3441);
and U4829 (N_4829,N_3517,N_3611);
nand U4830 (N_4830,N_3605,N_3178);
and U4831 (N_4831,N_3415,N_3291);
nand U4832 (N_4832,N_3773,N_3388);
xor U4833 (N_4833,N_3683,N_3571);
and U4834 (N_4834,N_3029,N_3078);
xor U4835 (N_4835,N_3344,N_3202);
xnor U4836 (N_4836,N_3654,N_3169);
nand U4837 (N_4837,N_3671,N_3903);
nand U4838 (N_4838,N_3715,N_3333);
and U4839 (N_4839,N_3869,N_3884);
nor U4840 (N_4840,N_3400,N_3379);
and U4841 (N_4841,N_3621,N_3021);
and U4842 (N_4842,N_3934,N_3655);
and U4843 (N_4843,N_3277,N_3801);
nor U4844 (N_4844,N_3482,N_3111);
or U4845 (N_4845,N_3410,N_3032);
or U4846 (N_4846,N_3376,N_3043);
nand U4847 (N_4847,N_3012,N_3862);
nor U4848 (N_4848,N_3844,N_3323);
or U4849 (N_4849,N_3353,N_3104);
nand U4850 (N_4850,N_3562,N_3549);
and U4851 (N_4851,N_3391,N_3859);
nor U4852 (N_4852,N_3587,N_3157);
nor U4853 (N_4853,N_3380,N_3814);
or U4854 (N_4854,N_3345,N_3248);
xor U4855 (N_4855,N_3326,N_3508);
and U4856 (N_4856,N_3319,N_3755);
nor U4857 (N_4857,N_3739,N_3586);
and U4858 (N_4858,N_3544,N_3401);
nor U4859 (N_4859,N_3836,N_3628);
nor U4860 (N_4860,N_3424,N_3396);
xnor U4861 (N_4861,N_3187,N_3131);
or U4862 (N_4862,N_3497,N_3994);
xor U4863 (N_4863,N_3194,N_3333);
nand U4864 (N_4864,N_3976,N_3908);
nor U4865 (N_4865,N_3482,N_3560);
or U4866 (N_4866,N_3060,N_3101);
or U4867 (N_4867,N_3123,N_3965);
and U4868 (N_4868,N_3095,N_3043);
or U4869 (N_4869,N_3474,N_3706);
nand U4870 (N_4870,N_3607,N_3664);
nand U4871 (N_4871,N_3184,N_3843);
xor U4872 (N_4872,N_3563,N_3631);
xor U4873 (N_4873,N_3623,N_3876);
nand U4874 (N_4874,N_3268,N_3953);
xnor U4875 (N_4875,N_3150,N_3919);
and U4876 (N_4876,N_3289,N_3967);
and U4877 (N_4877,N_3180,N_3519);
xor U4878 (N_4878,N_3666,N_3037);
and U4879 (N_4879,N_3948,N_3342);
and U4880 (N_4880,N_3873,N_3957);
nand U4881 (N_4881,N_3973,N_3872);
nand U4882 (N_4882,N_3866,N_3402);
nor U4883 (N_4883,N_3697,N_3414);
or U4884 (N_4884,N_3903,N_3460);
and U4885 (N_4885,N_3553,N_3270);
nor U4886 (N_4886,N_3867,N_3288);
nand U4887 (N_4887,N_3940,N_3280);
xor U4888 (N_4888,N_3214,N_3244);
nor U4889 (N_4889,N_3390,N_3744);
nand U4890 (N_4890,N_3458,N_3671);
nor U4891 (N_4891,N_3250,N_3246);
nand U4892 (N_4892,N_3050,N_3751);
or U4893 (N_4893,N_3416,N_3645);
xnor U4894 (N_4894,N_3746,N_3964);
and U4895 (N_4895,N_3407,N_3726);
nand U4896 (N_4896,N_3579,N_3674);
nor U4897 (N_4897,N_3503,N_3610);
and U4898 (N_4898,N_3563,N_3869);
or U4899 (N_4899,N_3019,N_3492);
and U4900 (N_4900,N_3782,N_3238);
nand U4901 (N_4901,N_3309,N_3771);
and U4902 (N_4902,N_3353,N_3792);
nand U4903 (N_4903,N_3436,N_3289);
nor U4904 (N_4904,N_3583,N_3979);
nor U4905 (N_4905,N_3896,N_3192);
or U4906 (N_4906,N_3503,N_3672);
nand U4907 (N_4907,N_3852,N_3579);
or U4908 (N_4908,N_3208,N_3009);
nor U4909 (N_4909,N_3163,N_3661);
and U4910 (N_4910,N_3898,N_3600);
xor U4911 (N_4911,N_3737,N_3611);
or U4912 (N_4912,N_3313,N_3551);
nor U4913 (N_4913,N_3282,N_3658);
xor U4914 (N_4914,N_3975,N_3909);
xnor U4915 (N_4915,N_3116,N_3111);
and U4916 (N_4916,N_3131,N_3271);
nand U4917 (N_4917,N_3666,N_3256);
nor U4918 (N_4918,N_3683,N_3255);
nand U4919 (N_4919,N_3261,N_3487);
nand U4920 (N_4920,N_3141,N_3871);
or U4921 (N_4921,N_3218,N_3851);
nor U4922 (N_4922,N_3120,N_3621);
nand U4923 (N_4923,N_3415,N_3029);
nor U4924 (N_4924,N_3566,N_3979);
nor U4925 (N_4925,N_3131,N_3721);
and U4926 (N_4926,N_3440,N_3724);
nand U4927 (N_4927,N_3510,N_3891);
xnor U4928 (N_4928,N_3202,N_3882);
or U4929 (N_4929,N_3244,N_3040);
nor U4930 (N_4930,N_3705,N_3852);
nand U4931 (N_4931,N_3912,N_3336);
nor U4932 (N_4932,N_3372,N_3989);
and U4933 (N_4933,N_3916,N_3839);
or U4934 (N_4934,N_3451,N_3773);
xor U4935 (N_4935,N_3048,N_3298);
or U4936 (N_4936,N_3764,N_3112);
nor U4937 (N_4937,N_3063,N_3870);
nand U4938 (N_4938,N_3939,N_3086);
xnor U4939 (N_4939,N_3998,N_3293);
and U4940 (N_4940,N_3949,N_3925);
nand U4941 (N_4941,N_3165,N_3285);
nand U4942 (N_4942,N_3938,N_3318);
or U4943 (N_4943,N_3393,N_3308);
and U4944 (N_4944,N_3464,N_3039);
xor U4945 (N_4945,N_3059,N_3310);
nor U4946 (N_4946,N_3212,N_3638);
or U4947 (N_4947,N_3255,N_3122);
or U4948 (N_4948,N_3130,N_3113);
xor U4949 (N_4949,N_3213,N_3414);
nand U4950 (N_4950,N_3598,N_3795);
nor U4951 (N_4951,N_3813,N_3127);
nand U4952 (N_4952,N_3184,N_3634);
nand U4953 (N_4953,N_3048,N_3498);
xnor U4954 (N_4954,N_3785,N_3996);
nor U4955 (N_4955,N_3909,N_3400);
nor U4956 (N_4956,N_3128,N_3941);
and U4957 (N_4957,N_3649,N_3332);
nand U4958 (N_4958,N_3963,N_3040);
nor U4959 (N_4959,N_3538,N_3302);
nor U4960 (N_4960,N_3596,N_3476);
nor U4961 (N_4961,N_3944,N_3519);
nand U4962 (N_4962,N_3858,N_3771);
xnor U4963 (N_4963,N_3166,N_3741);
nor U4964 (N_4964,N_3184,N_3348);
nor U4965 (N_4965,N_3128,N_3095);
or U4966 (N_4966,N_3526,N_3634);
nand U4967 (N_4967,N_3164,N_3022);
nor U4968 (N_4968,N_3289,N_3991);
nand U4969 (N_4969,N_3473,N_3547);
and U4970 (N_4970,N_3229,N_3231);
nand U4971 (N_4971,N_3287,N_3675);
nor U4972 (N_4972,N_3145,N_3245);
xnor U4973 (N_4973,N_3672,N_3482);
and U4974 (N_4974,N_3627,N_3927);
nor U4975 (N_4975,N_3951,N_3852);
nor U4976 (N_4976,N_3363,N_3248);
xnor U4977 (N_4977,N_3626,N_3512);
xor U4978 (N_4978,N_3236,N_3595);
nor U4979 (N_4979,N_3226,N_3921);
nor U4980 (N_4980,N_3486,N_3174);
and U4981 (N_4981,N_3380,N_3281);
or U4982 (N_4982,N_3784,N_3734);
or U4983 (N_4983,N_3015,N_3858);
and U4984 (N_4984,N_3632,N_3052);
and U4985 (N_4985,N_3076,N_3203);
and U4986 (N_4986,N_3988,N_3185);
xnor U4987 (N_4987,N_3047,N_3894);
nand U4988 (N_4988,N_3324,N_3079);
nand U4989 (N_4989,N_3478,N_3357);
or U4990 (N_4990,N_3295,N_3704);
or U4991 (N_4991,N_3647,N_3057);
xnor U4992 (N_4992,N_3812,N_3133);
xnor U4993 (N_4993,N_3662,N_3945);
and U4994 (N_4994,N_3895,N_3033);
nor U4995 (N_4995,N_3633,N_3520);
xor U4996 (N_4996,N_3884,N_3805);
xnor U4997 (N_4997,N_3162,N_3415);
and U4998 (N_4998,N_3565,N_3437);
nor U4999 (N_4999,N_3588,N_3956);
xor UO_0 (O_0,N_4263,N_4277);
xnor UO_1 (O_1,N_4102,N_4326);
and UO_2 (O_2,N_4231,N_4363);
nand UO_3 (O_3,N_4530,N_4626);
xor UO_4 (O_4,N_4307,N_4010);
or UO_5 (O_5,N_4364,N_4367);
nand UO_6 (O_6,N_4953,N_4808);
nand UO_7 (O_7,N_4924,N_4210);
nor UO_8 (O_8,N_4393,N_4731);
nand UO_9 (O_9,N_4400,N_4944);
or UO_10 (O_10,N_4700,N_4373);
or UO_11 (O_11,N_4289,N_4264);
nand UO_12 (O_12,N_4122,N_4043);
xor UO_13 (O_13,N_4872,N_4813);
and UO_14 (O_14,N_4539,N_4323);
xnor UO_15 (O_15,N_4517,N_4108);
xor UO_16 (O_16,N_4151,N_4800);
or UO_17 (O_17,N_4505,N_4491);
xnor UO_18 (O_18,N_4474,N_4062);
xor UO_19 (O_19,N_4567,N_4015);
or UO_20 (O_20,N_4658,N_4466);
nor UO_21 (O_21,N_4313,N_4476);
and UO_22 (O_22,N_4071,N_4411);
and UO_23 (O_23,N_4493,N_4919);
xor UO_24 (O_24,N_4424,N_4926);
xor UO_25 (O_25,N_4041,N_4128);
and UO_26 (O_26,N_4633,N_4627);
nor UO_27 (O_27,N_4479,N_4905);
or UO_28 (O_28,N_4136,N_4087);
nand UO_29 (O_29,N_4114,N_4003);
or UO_30 (O_30,N_4065,N_4645);
xnor UO_31 (O_31,N_4646,N_4399);
nor UO_32 (O_32,N_4750,N_4053);
and UO_33 (O_33,N_4341,N_4511);
xor UO_34 (O_34,N_4427,N_4788);
or UO_35 (O_35,N_4469,N_4647);
xor UO_36 (O_36,N_4580,N_4274);
nor UO_37 (O_37,N_4724,N_4258);
xnor UO_38 (O_38,N_4142,N_4625);
nor UO_39 (O_39,N_4239,N_4999);
or UO_40 (O_40,N_4134,N_4764);
nand UO_41 (O_41,N_4890,N_4506);
nand UO_42 (O_42,N_4771,N_4542);
and UO_43 (O_43,N_4013,N_4722);
nand UO_44 (O_44,N_4310,N_4358);
nor UO_45 (O_45,N_4643,N_4443);
nand UO_46 (O_46,N_4002,N_4436);
nand UO_47 (O_47,N_4862,N_4751);
xnor UO_48 (O_48,N_4713,N_4587);
xor UO_49 (O_49,N_4175,N_4182);
nand UO_50 (O_50,N_4908,N_4100);
or UO_51 (O_51,N_4604,N_4670);
and UO_52 (O_52,N_4847,N_4284);
or UO_53 (O_53,N_4932,N_4941);
nand UO_54 (O_54,N_4064,N_4471);
or UO_55 (O_55,N_4818,N_4060);
nor UO_56 (O_56,N_4662,N_4702);
xnor UO_57 (O_57,N_4431,N_4532);
and UO_58 (O_58,N_4291,N_4714);
and UO_59 (O_59,N_4778,N_4718);
or UO_60 (O_60,N_4189,N_4287);
and UO_61 (O_61,N_4195,N_4732);
or UO_62 (O_62,N_4972,N_4820);
and UO_63 (O_63,N_4384,N_4918);
or UO_64 (O_64,N_4009,N_4024);
nor UO_65 (O_65,N_4769,N_4947);
nand UO_66 (O_66,N_4655,N_4765);
xor UO_67 (O_67,N_4744,N_4472);
and UO_68 (O_68,N_4028,N_4331);
and UO_69 (O_69,N_4164,N_4935);
or UO_70 (O_70,N_4343,N_4279);
nor UO_71 (O_71,N_4300,N_4321);
and UO_72 (O_72,N_4611,N_4385);
nand UO_73 (O_73,N_4698,N_4753);
nand UO_74 (O_74,N_4792,N_4586);
xnor UO_75 (O_75,N_4169,N_4172);
or UO_76 (O_76,N_4735,N_4861);
or UO_77 (O_77,N_4401,N_4336);
and UO_78 (O_78,N_4149,N_4676);
nand UO_79 (O_79,N_4990,N_4319);
nor UO_80 (O_80,N_4799,N_4420);
nand UO_81 (O_81,N_4152,N_4333);
nand UO_82 (O_82,N_4717,N_4876);
nand UO_83 (O_83,N_4679,N_4807);
nand UO_84 (O_84,N_4602,N_4844);
and UO_85 (O_85,N_4892,N_4803);
or UO_86 (O_86,N_4683,N_4170);
xor UO_87 (O_87,N_4330,N_4523);
or UO_88 (O_88,N_4407,N_4081);
or UO_89 (O_89,N_4388,N_4755);
or UO_90 (O_90,N_4644,N_4229);
or UO_91 (O_91,N_4456,N_4797);
nor UO_92 (O_92,N_4337,N_4144);
xnor UO_93 (O_93,N_4954,N_4695);
xnor UO_94 (O_94,N_4510,N_4020);
or UO_95 (O_95,N_4158,N_4641);
or UO_96 (O_96,N_4680,N_4311);
nor UO_97 (O_97,N_4501,N_4775);
or UO_98 (O_98,N_4250,N_4459);
nor UO_99 (O_99,N_4889,N_4334);
or UO_100 (O_100,N_4933,N_4078);
and UO_101 (O_101,N_4458,N_4034);
xor UO_102 (O_102,N_4119,N_4225);
nand UO_103 (O_103,N_4368,N_4162);
and UO_104 (O_104,N_4871,N_4867);
xnor UO_105 (O_105,N_4904,N_4594);
and UO_106 (O_106,N_4754,N_4256);
and UO_107 (O_107,N_4568,N_4187);
nand UO_108 (O_108,N_4138,N_4135);
nor UO_109 (O_109,N_4906,N_4661);
nor UO_110 (O_110,N_4032,N_4885);
nand UO_111 (O_111,N_4692,N_4677);
and UO_112 (O_112,N_4910,N_4981);
xor UO_113 (O_113,N_4579,N_4622);
nor UO_114 (O_114,N_4619,N_4812);
and UO_115 (O_115,N_4605,N_4133);
and UO_116 (O_116,N_4541,N_4371);
and UO_117 (O_117,N_4545,N_4345);
or UO_118 (O_118,N_4632,N_4252);
xor UO_119 (O_119,N_4507,N_4917);
nor UO_120 (O_120,N_4283,N_4016);
or UO_121 (O_121,N_4033,N_4980);
or UO_122 (O_122,N_4901,N_4050);
and UO_123 (O_123,N_4883,N_4590);
and UO_124 (O_124,N_4729,N_4488);
nand UO_125 (O_125,N_4730,N_4747);
and UO_126 (O_126,N_4261,N_4983);
or UO_127 (O_127,N_4249,N_4809);
and UO_128 (O_128,N_4720,N_4549);
or UO_129 (O_129,N_4091,N_4352);
xor UO_130 (O_130,N_4949,N_4092);
and UO_131 (O_131,N_4963,N_4217);
xnor UO_132 (O_132,N_4780,N_4811);
nor UO_133 (O_133,N_4665,N_4094);
nand UO_134 (O_134,N_4098,N_4601);
nand UO_135 (O_135,N_4925,N_4849);
xnor UO_136 (O_136,N_4379,N_4804);
nand UO_137 (O_137,N_4841,N_4327);
xor UO_138 (O_138,N_4259,N_4794);
and UO_139 (O_139,N_4609,N_4445);
or UO_140 (O_140,N_4685,N_4502);
or UO_141 (O_141,N_4913,N_4543);
or UO_142 (O_142,N_4518,N_4682);
and UO_143 (O_143,N_4173,N_4597);
xor UO_144 (O_144,N_4442,N_4974);
nand UO_145 (O_145,N_4691,N_4801);
and UO_146 (O_146,N_4705,N_4104);
or UO_147 (O_147,N_4988,N_4834);
or UO_148 (O_148,N_4779,N_4783);
xnor UO_149 (O_149,N_4480,N_4752);
nor UO_150 (O_150,N_4821,N_4948);
and UO_151 (O_151,N_4846,N_4884);
nor UO_152 (O_152,N_4235,N_4638);
xor UO_153 (O_153,N_4276,N_4045);
nand UO_154 (O_154,N_4435,N_4600);
nand UO_155 (O_155,N_4085,N_4127);
nand UO_156 (O_156,N_4054,N_4631);
or UO_157 (O_157,N_4278,N_4194);
xor UO_158 (O_158,N_4453,N_4332);
nor UO_159 (O_159,N_4951,N_4810);
and UO_160 (O_160,N_4030,N_4011);
or UO_161 (O_161,N_4186,N_4761);
xnor UO_162 (O_162,N_4112,N_4558);
or UO_163 (O_163,N_4725,N_4666);
xor UO_164 (O_164,N_4879,N_4140);
nand UO_165 (O_165,N_4690,N_4095);
or UO_166 (O_166,N_4154,N_4025);
xnor UO_167 (O_167,N_4618,N_4969);
or UO_168 (O_168,N_4124,N_4840);
nand UO_169 (O_169,N_4971,N_4262);
or UO_170 (O_170,N_4483,N_4975);
or UO_171 (O_171,N_4056,N_4433);
and UO_172 (O_172,N_4342,N_4293);
nand UO_173 (O_173,N_4396,N_4001);
xor UO_174 (O_174,N_4785,N_4719);
nor UO_175 (O_175,N_4147,N_4939);
nor UO_176 (O_176,N_4961,N_4909);
or UO_177 (O_177,N_4674,N_4688);
nor UO_178 (O_178,N_4606,N_4891);
and UO_179 (O_179,N_4759,N_4096);
or UO_180 (O_180,N_4425,N_4773);
nand UO_181 (O_181,N_4268,N_4648);
and UO_182 (O_182,N_4495,N_4377);
nand UO_183 (O_183,N_4426,N_4937);
and UO_184 (O_184,N_4607,N_4205);
or UO_185 (O_185,N_4856,N_4072);
or UO_186 (O_186,N_4160,N_4074);
nand UO_187 (O_187,N_4477,N_4304);
xor UO_188 (O_188,N_4843,N_4726);
or UO_189 (O_189,N_4075,N_4766);
nor UO_190 (O_190,N_4624,N_4599);
nand UO_191 (O_191,N_4533,N_4382);
or UO_192 (O_192,N_4418,N_4111);
nand UO_193 (O_193,N_4475,N_4208);
nor UO_194 (O_194,N_4903,N_4563);
and UO_195 (O_195,N_4450,N_4895);
nand UO_196 (O_196,N_4850,N_4389);
or UO_197 (O_197,N_4012,N_4070);
nand UO_198 (O_198,N_4802,N_4328);
nand UO_199 (O_199,N_4593,N_4109);
nor UO_200 (O_200,N_4569,N_4203);
nor UO_201 (O_201,N_4415,N_4965);
and UO_202 (O_202,N_4733,N_4077);
or UO_203 (O_203,N_4831,N_4936);
xnor UO_204 (O_204,N_4893,N_4318);
nand UO_205 (O_205,N_4608,N_4955);
xor UO_206 (O_206,N_4874,N_4575);
and UO_207 (O_207,N_4694,N_4171);
or UO_208 (O_208,N_4985,N_4537);
or UO_209 (O_209,N_4762,N_4551);
nor UO_210 (O_210,N_4260,N_4206);
nand UO_211 (O_211,N_4219,N_4784);
and UO_212 (O_212,N_4930,N_4487);
xor UO_213 (O_213,N_4166,N_4176);
xor UO_214 (O_214,N_4413,N_4434);
xnor UO_215 (O_215,N_4828,N_4522);
nand UO_216 (O_216,N_4022,N_4979);
and UO_217 (O_217,N_4723,N_4196);
nor UO_218 (O_218,N_4430,N_4216);
and UO_219 (O_219,N_4736,N_4423);
and UO_220 (O_220,N_4390,N_4052);
or UO_221 (O_221,N_4929,N_4148);
nor UO_222 (O_222,N_4994,N_4496);
xor UO_223 (O_223,N_4370,N_4295);
nand UO_224 (O_224,N_4155,N_4806);
and UO_225 (O_225,N_4848,N_4888);
nand UO_226 (O_226,N_4129,N_4870);
xnor UO_227 (O_227,N_4721,N_4978);
and UO_228 (O_228,N_4439,N_4226);
or UO_229 (O_229,N_4598,N_4675);
or UO_230 (O_230,N_4687,N_4153);
and UO_231 (O_231,N_4592,N_4869);
xor UO_232 (O_232,N_4966,N_4835);
xnor UO_233 (O_233,N_4512,N_4576);
or UO_234 (O_234,N_4416,N_4707);
and UO_235 (O_235,N_4743,N_4654);
or UO_236 (O_236,N_4465,N_4494);
or UO_237 (O_237,N_4406,N_4902);
xnor UO_238 (O_238,N_4193,N_4000);
nor UO_239 (O_239,N_4757,N_4945);
xor UO_240 (O_240,N_4452,N_4642);
and UO_241 (O_241,N_4199,N_4218);
xor UO_242 (O_242,N_4402,N_4612);
nor UO_243 (O_243,N_4791,N_4673);
or UO_244 (O_244,N_4531,N_4460);
and UO_245 (O_245,N_4760,N_4019);
xor UO_246 (O_246,N_4224,N_4991);
nand UO_247 (O_247,N_4823,N_4438);
nand UO_248 (O_248,N_4696,N_4536);
and UO_249 (O_249,N_4281,N_4865);
and UO_250 (O_250,N_4860,N_4179);
and UO_251 (O_251,N_4042,N_4005);
or UO_252 (O_252,N_4497,N_4286);
xnor UO_253 (O_253,N_4516,N_4786);
nor UO_254 (O_254,N_4697,N_4348);
xor UO_255 (O_255,N_4417,N_4527);
and UO_256 (O_256,N_4428,N_4623);
and UO_257 (O_257,N_4858,N_4710);
nor UO_258 (O_258,N_4620,N_4851);
and UO_259 (O_259,N_4741,N_4316);
xnor UO_260 (O_260,N_4664,N_4204);
and UO_261 (O_261,N_4080,N_4827);
xnor UO_262 (O_262,N_4392,N_4589);
or UO_263 (O_263,N_4198,N_4559);
nor UO_264 (O_264,N_4068,N_4447);
or UO_265 (O_265,N_4163,N_4270);
nor UO_266 (O_266,N_4237,N_4560);
nor UO_267 (O_267,N_4920,N_4635);
nor UO_268 (O_268,N_4120,N_4649);
nand UO_269 (O_269,N_4395,N_4184);
and UO_270 (O_270,N_4581,N_4035);
nand UO_271 (O_271,N_4150,N_4269);
and UO_272 (O_272,N_4046,N_4914);
nand UO_273 (O_273,N_4353,N_4457);
or UO_274 (O_274,N_4728,N_4448);
and UO_275 (O_275,N_4044,N_4329);
nand UO_276 (O_276,N_4830,N_4790);
nand UO_277 (O_277,N_4950,N_4976);
nand UO_278 (O_278,N_4738,N_4898);
nand UO_279 (O_279,N_4796,N_4873);
nand UO_280 (O_280,N_4115,N_4704);
and UO_281 (O_281,N_4473,N_4272);
or UO_282 (O_282,N_4900,N_4181);
or UO_283 (O_283,N_4386,N_4230);
nand UO_284 (O_284,N_4995,N_4526);
xor UO_285 (O_285,N_4959,N_4273);
xnor UO_286 (O_286,N_4361,N_4894);
nor UO_287 (O_287,N_4238,N_4912);
xnor UO_288 (O_288,N_4763,N_4659);
or UO_289 (O_289,N_4556,N_4992);
or UO_290 (O_290,N_4957,N_4322);
xnor UO_291 (O_291,N_4324,N_4774);
nor UO_292 (O_292,N_4756,N_4868);
xnor UO_293 (O_293,N_4500,N_4671);
or UO_294 (O_294,N_4212,N_4076);
nor UO_295 (O_295,N_4440,N_4907);
nand UO_296 (O_296,N_4201,N_4699);
or UO_297 (O_297,N_4528,N_4777);
nor UO_298 (O_298,N_4574,N_4615);
and UO_299 (O_299,N_4737,N_4478);
nor UO_300 (O_300,N_4183,N_4236);
nand UO_301 (O_301,N_4770,N_4651);
xnor UO_302 (O_302,N_4202,N_4866);
nor UO_303 (O_303,N_4234,N_4798);
xnor UO_304 (O_304,N_4577,N_4668);
or UO_305 (O_305,N_4294,N_4829);
nand UO_306 (O_306,N_4842,N_4547);
xnor UO_307 (O_307,N_4548,N_4781);
nand UO_308 (O_308,N_4339,N_4958);
nand UO_309 (O_309,N_4421,N_4561);
xor UO_310 (O_310,N_4837,N_4652);
and UO_311 (O_311,N_4964,N_4365);
nand UO_312 (O_312,N_4970,N_4446);
or UO_313 (O_313,N_4582,N_4657);
and UO_314 (O_314,N_4701,N_4603);
or UO_315 (O_315,N_4055,N_4555);
or UO_316 (O_316,N_4525,N_4931);
nand UO_317 (O_317,N_4093,N_4303);
and UO_318 (O_318,N_4793,N_4513);
nand UO_319 (O_319,N_4610,N_4159);
nor UO_320 (O_320,N_4485,N_4854);
nand UO_321 (O_321,N_4667,N_4090);
or UO_322 (O_322,N_4228,N_4137);
nand UO_323 (O_323,N_4956,N_4708);
and UO_324 (O_324,N_4314,N_4853);
and UO_325 (O_325,N_4767,N_4038);
nor UO_326 (O_326,N_4117,N_4372);
nand UO_327 (O_327,N_4629,N_4529);
xnor UO_328 (O_328,N_4296,N_4110);
nand UO_329 (O_329,N_4192,N_4508);
or UO_330 (O_330,N_4029,N_4143);
xor UO_331 (O_331,N_4486,N_4063);
xnor UO_332 (O_332,N_4214,N_4245);
nand UO_333 (O_333,N_4463,N_4107);
or UO_334 (O_334,N_4165,N_4489);
nor UO_335 (O_335,N_4878,N_4940);
nand UO_336 (O_336,N_4244,N_4742);
nand UO_337 (O_337,N_4213,N_4839);
or UO_338 (O_338,N_4405,N_4515);
nand UO_339 (O_339,N_4734,N_4131);
xnor UO_340 (O_340,N_4130,N_4023);
nor UO_341 (O_341,N_4061,N_4394);
nand UO_342 (O_342,N_4359,N_4583);
or UO_343 (O_343,N_4350,N_4344);
or UO_344 (O_344,N_4161,N_4437);
and UO_345 (O_345,N_4309,N_4200);
nand UO_346 (O_346,N_4007,N_4266);
nand UO_347 (O_347,N_4106,N_4265);
and UO_348 (O_348,N_4197,N_4375);
or UO_349 (O_349,N_4188,N_4887);
xor UO_350 (O_350,N_4922,N_4544);
nand UO_351 (O_351,N_4103,N_4538);
nor UO_352 (O_352,N_4403,N_4715);
or UO_353 (O_353,N_4565,N_4257);
or UO_354 (O_354,N_4315,N_4146);
nand UO_355 (O_355,N_4740,N_4566);
nor UO_356 (O_356,N_4338,N_4468);
or UO_357 (O_357,N_4317,N_4768);
nor UO_358 (O_358,N_4996,N_4748);
or UO_359 (O_359,N_4557,N_4251);
xnor UO_360 (O_360,N_4628,N_4335);
xnor UO_361 (O_361,N_4099,N_4380);
and UO_362 (O_362,N_4121,N_4241);
or UO_363 (O_363,N_4145,N_4464);
and UO_364 (O_364,N_4306,N_4772);
xor UO_365 (O_365,N_4058,N_4596);
nand UO_366 (O_366,N_4320,N_4490);
xor UO_367 (O_367,N_4968,N_4614);
or UO_368 (O_368,N_4573,N_4636);
xor UO_369 (O_369,N_4031,N_4967);
nor UO_370 (O_370,N_4126,N_4116);
xor UO_371 (O_371,N_4066,N_4223);
nor UO_372 (O_372,N_4190,N_4378);
and UO_373 (O_373,N_4745,N_4938);
and UO_374 (O_374,N_4073,N_4180);
nor UO_375 (O_375,N_4298,N_4832);
nor UO_376 (O_376,N_4191,N_4355);
and UO_377 (O_377,N_4470,N_4585);
nor UO_378 (O_378,N_4101,N_4057);
nand UO_379 (O_379,N_4449,N_4037);
xnor UO_380 (O_380,N_4141,N_4357);
nor UO_381 (O_381,N_4362,N_4749);
nor UO_382 (O_382,N_4982,N_4292);
or UO_383 (O_383,N_4816,N_4776);
nand UO_384 (O_384,N_4082,N_4617);
and UO_385 (O_385,N_4211,N_4481);
nand UO_386 (O_386,N_4014,N_4552);
nor UO_387 (O_387,N_4845,N_4681);
or UO_388 (O_388,N_4863,N_4634);
nand UO_389 (O_389,N_4578,N_4167);
and UO_390 (O_390,N_4410,N_4021);
nor UO_391 (O_391,N_4215,N_4899);
nand UO_392 (O_392,N_4267,N_4534);
nor UO_393 (O_393,N_4039,N_4650);
or UO_394 (O_394,N_4026,N_4584);
nand UO_395 (O_395,N_4067,N_4360);
nand UO_396 (O_396,N_4498,N_4275);
xor UO_397 (O_397,N_4989,N_4672);
and UO_398 (O_398,N_4562,N_4059);
or UO_399 (O_399,N_4817,N_4168);
and UO_400 (O_400,N_4325,N_4514);
nor UO_401 (O_401,N_4739,N_4875);
nand UO_402 (O_402,N_4069,N_4911);
xor UO_403 (O_403,N_4962,N_4018);
nand UO_404 (O_404,N_4571,N_4105);
nand UO_405 (O_405,N_4444,N_4916);
xnor UO_406 (O_406,N_4942,N_4977);
xor UO_407 (O_407,N_4369,N_4987);
nand UO_408 (O_408,N_4553,N_4246);
nand UO_409 (O_409,N_4441,N_4630);
nand UO_410 (O_410,N_4248,N_4254);
nor UO_411 (O_411,N_4383,N_4880);
nand UO_412 (O_412,N_4222,N_4637);
and UO_413 (O_413,N_4660,N_4882);
or UO_414 (O_414,N_4156,N_4946);
nor UO_415 (O_415,N_4684,N_4240);
and UO_416 (O_416,N_4591,N_4290);
nor UO_417 (O_417,N_4125,N_4716);
nor UO_418 (O_418,N_4815,N_4006);
or UO_419 (O_419,N_4340,N_4669);
and UO_420 (O_420,N_4712,N_4419);
xnor UO_421 (O_421,N_4540,N_4524);
xnor UO_422 (O_422,N_4454,N_4086);
and UO_423 (O_423,N_4404,N_4787);
nor UO_424 (O_424,N_4049,N_4795);
nor UO_425 (O_425,N_4381,N_4952);
nor UO_426 (O_426,N_4588,N_4079);
xnor UO_427 (O_427,N_4209,N_4689);
and UO_428 (O_428,N_4288,N_4709);
or UO_429 (O_429,N_4960,N_4758);
nand UO_430 (O_430,N_4233,N_4178);
and UO_431 (O_431,N_4550,N_4047);
and UO_432 (O_432,N_4451,N_4927);
nand UO_433 (O_433,N_4509,N_4822);
and UO_434 (O_434,N_4247,N_4613);
or UO_435 (O_435,N_4727,N_4857);
nor UO_436 (O_436,N_4639,N_4703);
xor UO_437 (O_437,N_4896,N_4461);
and UO_438 (O_438,N_4414,N_4640);
or UO_439 (O_439,N_4123,N_4432);
or UO_440 (O_440,N_4521,N_4928);
and UO_441 (O_441,N_4484,N_4897);
nor UO_442 (O_442,N_4299,N_4409);
nor UO_443 (O_443,N_4242,N_4356);
nor UO_444 (O_444,N_4805,N_4572);
or UO_445 (O_445,N_4221,N_4746);
or UO_446 (O_446,N_4852,N_4789);
xnor UO_447 (O_447,N_4998,N_4881);
nand UO_448 (O_448,N_4921,N_4301);
and UO_449 (O_449,N_4084,N_4017);
nand UO_450 (O_450,N_4297,N_4398);
and UO_451 (O_451,N_4243,N_4285);
xor UO_452 (O_452,N_4376,N_4455);
or UO_453 (O_453,N_4412,N_4185);
nand UO_454 (O_454,N_4374,N_4482);
or UO_455 (O_455,N_4554,N_4113);
or UO_456 (O_456,N_4253,N_4864);
nand UO_457 (O_457,N_4915,N_4351);
nor UO_458 (O_458,N_4347,N_4826);
xor UO_459 (O_459,N_4877,N_4220);
and UO_460 (O_460,N_4305,N_4346);
nand UO_461 (O_461,N_4693,N_4535);
nor UO_462 (O_462,N_4711,N_4656);
nand UO_463 (O_463,N_4255,N_4923);
and UO_464 (O_464,N_4973,N_4984);
or UO_465 (O_465,N_4051,N_4934);
nand UO_466 (O_466,N_4036,N_4177);
xnor UO_467 (O_467,N_4422,N_4408);
or UO_468 (O_468,N_4997,N_4004);
nor UO_469 (O_469,N_4782,N_4349);
nor UO_470 (O_470,N_4616,N_4089);
nand UO_471 (O_471,N_4040,N_4097);
nand UO_472 (O_472,N_4519,N_4083);
xnor UO_473 (O_473,N_4621,N_4008);
xor UO_474 (O_474,N_4271,N_4663);
and UO_475 (O_475,N_4429,N_4227);
nand UO_476 (O_476,N_4492,N_4088);
nor UO_477 (O_477,N_4387,N_4157);
xor UO_478 (O_478,N_4819,N_4118);
nand UO_479 (O_479,N_4503,N_4836);
nand UO_480 (O_480,N_4366,N_4993);
nand UO_481 (O_481,N_4855,N_4678);
or UO_482 (O_482,N_4467,N_4706);
and UO_483 (O_483,N_4838,N_4280);
nand UO_484 (O_484,N_4354,N_4139);
nand UO_485 (O_485,N_4825,N_4520);
or UO_486 (O_486,N_4986,N_4686);
xor UO_487 (O_487,N_4174,N_4833);
nor UO_488 (O_488,N_4546,N_4595);
nor UO_489 (O_489,N_4391,N_4462);
or UO_490 (O_490,N_4859,N_4302);
and UO_491 (O_491,N_4653,N_4564);
nand UO_492 (O_492,N_4814,N_4570);
nand UO_493 (O_493,N_4282,N_4886);
and UO_494 (O_494,N_4048,N_4943);
nor UO_495 (O_495,N_4499,N_4397);
and UO_496 (O_496,N_4308,N_4132);
nor UO_497 (O_497,N_4824,N_4504);
nand UO_498 (O_498,N_4027,N_4232);
nand UO_499 (O_499,N_4312,N_4207);
or UO_500 (O_500,N_4821,N_4638);
nor UO_501 (O_501,N_4253,N_4507);
nand UO_502 (O_502,N_4133,N_4527);
and UO_503 (O_503,N_4813,N_4153);
or UO_504 (O_504,N_4433,N_4257);
or UO_505 (O_505,N_4882,N_4308);
nor UO_506 (O_506,N_4432,N_4009);
xnor UO_507 (O_507,N_4630,N_4046);
xnor UO_508 (O_508,N_4650,N_4730);
nand UO_509 (O_509,N_4989,N_4847);
nand UO_510 (O_510,N_4586,N_4159);
nand UO_511 (O_511,N_4332,N_4283);
xnor UO_512 (O_512,N_4240,N_4617);
or UO_513 (O_513,N_4882,N_4387);
and UO_514 (O_514,N_4618,N_4928);
xnor UO_515 (O_515,N_4503,N_4778);
nand UO_516 (O_516,N_4801,N_4376);
nor UO_517 (O_517,N_4774,N_4488);
and UO_518 (O_518,N_4623,N_4456);
nand UO_519 (O_519,N_4230,N_4579);
or UO_520 (O_520,N_4484,N_4299);
nor UO_521 (O_521,N_4615,N_4929);
and UO_522 (O_522,N_4854,N_4582);
and UO_523 (O_523,N_4478,N_4340);
nor UO_524 (O_524,N_4868,N_4477);
or UO_525 (O_525,N_4462,N_4081);
or UO_526 (O_526,N_4487,N_4268);
nor UO_527 (O_527,N_4984,N_4544);
and UO_528 (O_528,N_4156,N_4420);
nor UO_529 (O_529,N_4063,N_4787);
or UO_530 (O_530,N_4192,N_4642);
or UO_531 (O_531,N_4310,N_4143);
xnor UO_532 (O_532,N_4424,N_4005);
and UO_533 (O_533,N_4810,N_4610);
or UO_534 (O_534,N_4171,N_4659);
or UO_535 (O_535,N_4591,N_4187);
xnor UO_536 (O_536,N_4267,N_4079);
xnor UO_537 (O_537,N_4610,N_4442);
and UO_538 (O_538,N_4704,N_4306);
xor UO_539 (O_539,N_4325,N_4874);
nand UO_540 (O_540,N_4216,N_4497);
nor UO_541 (O_541,N_4890,N_4911);
or UO_542 (O_542,N_4242,N_4534);
and UO_543 (O_543,N_4185,N_4688);
and UO_544 (O_544,N_4544,N_4026);
nor UO_545 (O_545,N_4298,N_4003);
nor UO_546 (O_546,N_4737,N_4809);
nand UO_547 (O_547,N_4361,N_4387);
and UO_548 (O_548,N_4979,N_4507);
or UO_549 (O_549,N_4582,N_4991);
nand UO_550 (O_550,N_4012,N_4044);
xor UO_551 (O_551,N_4967,N_4716);
nand UO_552 (O_552,N_4601,N_4529);
nor UO_553 (O_553,N_4040,N_4268);
nand UO_554 (O_554,N_4285,N_4266);
and UO_555 (O_555,N_4978,N_4997);
xor UO_556 (O_556,N_4220,N_4285);
xor UO_557 (O_557,N_4294,N_4754);
xnor UO_558 (O_558,N_4582,N_4407);
and UO_559 (O_559,N_4107,N_4801);
xnor UO_560 (O_560,N_4289,N_4736);
nor UO_561 (O_561,N_4692,N_4192);
or UO_562 (O_562,N_4940,N_4232);
xnor UO_563 (O_563,N_4812,N_4313);
xnor UO_564 (O_564,N_4691,N_4704);
and UO_565 (O_565,N_4400,N_4379);
nor UO_566 (O_566,N_4130,N_4011);
nand UO_567 (O_567,N_4797,N_4006);
or UO_568 (O_568,N_4330,N_4640);
or UO_569 (O_569,N_4958,N_4867);
and UO_570 (O_570,N_4879,N_4062);
and UO_571 (O_571,N_4910,N_4455);
and UO_572 (O_572,N_4293,N_4348);
and UO_573 (O_573,N_4615,N_4579);
nor UO_574 (O_574,N_4147,N_4608);
and UO_575 (O_575,N_4014,N_4750);
nand UO_576 (O_576,N_4765,N_4809);
or UO_577 (O_577,N_4309,N_4053);
xnor UO_578 (O_578,N_4434,N_4004);
xor UO_579 (O_579,N_4101,N_4823);
xor UO_580 (O_580,N_4087,N_4956);
or UO_581 (O_581,N_4239,N_4225);
and UO_582 (O_582,N_4890,N_4257);
nand UO_583 (O_583,N_4897,N_4906);
nand UO_584 (O_584,N_4661,N_4212);
or UO_585 (O_585,N_4384,N_4454);
nand UO_586 (O_586,N_4349,N_4076);
nor UO_587 (O_587,N_4665,N_4147);
or UO_588 (O_588,N_4559,N_4450);
and UO_589 (O_589,N_4154,N_4196);
xor UO_590 (O_590,N_4883,N_4460);
nor UO_591 (O_591,N_4828,N_4127);
nor UO_592 (O_592,N_4454,N_4192);
nand UO_593 (O_593,N_4416,N_4895);
nor UO_594 (O_594,N_4794,N_4387);
nand UO_595 (O_595,N_4360,N_4235);
xnor UO_596 (O_596,N_4893,N_4176);
and UO_597 (O_597,N_4303,N_4554);
nand UO_598 (O_598,N_4221,N_4664);
nand UO_599 (O_599,N_4597,N_4133);
nand UO_600 (O_600,N_4483,N_4079);
nand UO_601 (O_601,N_4137,N_4510);
nand UO_602 (O_602,N_4182,N_4300);
and UO_603 (O_603,N_4109,N_4280);
and UO_604 (O_604,N_4457,N_4459);
nand UO_605 (O_605,N_4448,N_4618);
xor UO_606 (O_606,N_4145,N_4992);
nor UO_607 (O_607,N_4195,N_4340);
xor UO_608 (O_608,N_4771,N_4633);
nor UO_609 (O_609,N_4768,N_4398);
or UO_610 (O_610,N_4538,N_4382);
xnor UO_611 (O_611,N_4043,N_4005);
nor UO_612 (O_612,N_4334,N_4532);
nand UO_613 (O_613,N_4973,N_4889);
xor UO_614 (O_614,N_4557,N_4519);
xor UO_615 (O_615,N_4987,N_4554);
nand UO_616 (O_616,N_4042,N_4030);
nand UO_617 (O_617,N_4427,N_4181);
xnor UO_618 (O_618,N_4117,N_4714);
or UO_619 (O_619,N_4921,N_4345);
xnor UO_620 (O_620,N_4984,N_4350);
nand UO_621 (O_621,N_4359,N_4082);
or UO_622 (O_622,N_4354,N_4134);
or UO_623 (O_623,N_4129,N_4815);
and UO_624 (O_624,N_4514,N_4353);
nor UO_625 (O_625,N_4000,N_4006);
nand UO_626 (O_626,N_4605,N_4494);
or UO_627 (O_627,N_4585,N_4478);
or UO_628 (O_628,N_4320,N_4369);
nor UO_629 (O_629,N_4696,N_4745);
nand UO_630 (O_630,N_4086,N_4336);
nand UO_631 (O_631,N_4113,N_4395);
nand UO_632 (O_632,N_4185,N_4074);
xnor UO_633 (O_633,N_4231,N_4006);
and UO_634 (O_634,N_4891,N_4946);
and UO_635 (O_635,N_4035,N_4260);
and UO_636 (O_636,N_4552,N_4759);
nor UO_637 (O_637,N_4241,N_4302);
nor UO_638 (O_638,N_4943,N_4538);
and UO_639 (O_639,N_4529,N_4536);
or UO_640 (O_640,N_4462,N_4496);
nor UO_641 (O_641,N_4579,N_4684);
xor UO_642 (O_642,N_4589,N_4444);
xor UO_643 (O_643,N_4329,N_4832);
xor UO_644 (O_644,N_4351,N_4204);
or UO_645 (O_645,N_4573,N_4001);
and UO_646 (O_646,N_4493,N_4087);
or UO_647 (O_647,N_4883,N_4014);
nand UO_648 (O_648,N_4630,N_4563);
nand UO_649 (O_649,N_4764,N_4324);
nor UO_650 (O_650,N_4206,N_4419);
nand UO_651 (O_651,N_4196,N_4340);
xnor UO_652 (O_652,N_4234,N_4587);
nor UO_653 (O_653,N_4370,N_4952);
xnor UO_654 (O_654,N_4374,N_4319);
and UO_655 (O_655,N_4661,N_4889);
and UO_656 (O_656,N_4239,N_4017);
xnor UO_657 (O_657,N_4036,N_4725);
nor UO_658 (O_658,N_4351,N_4063);
or UO_659 (O_659,N_4722,N_4249);
or UO_660 (O_660,N_4639,N_4276);
nor UO_661 (O_661,N_4833,N_4128);
nor UO_662 (O_662,N_4182,N_4896);
nor UO_663 (O_663,N_4145,N_4572);
or UO_664 (O_664,N_4054,N_4149);
or UO_665 (O_665,N_4983,N_4819);
and UO_666 (O_666,N_4120,N_4284);
and UO_667 (O_667,N_4754,N_4775);
xnor UO_668 (O_668,N_4797,N_4784);
or UO_669 (O_669,N_4540,N_4924);
xor UO_670 (O_670,N_4130,N_4132);
and UO_671 (O_671,N_4801,N_4308);
xor UO_672 (O_672,N_4774,N_4416);
nand UO_673 (O_673,N_4888,N_4309);
and UO_674 (O_674,N_4787,N_4999);
or UO_675 (O_675,N_4081,N_4233);
and UO_676 (O_676,N_4961,N_4383);
nand UO_677 (O_677,N_4326,N_4805);
and UO_678 (O_678,N_4734,N_4280);
nor UO_679 (O_679,N_4092,N_4268);
nand UO_680 (O_680,N_4239,N_4562);
nand UO_681 (O_681,N_4615,N_4459);
xnor UO_682 (O_682,N_4789,N_4592);
xor UO_683 (O_683,N_4267,N_4912);
nand UO_684 (O_684,N_4296,N_4723);
nand UO_685 (O_685,N_4655,N_4501);
xor UO_686 (O_686,N_4930,N_4086);
or UO_687 (O_687,N_4063,N_4271);
nand UO_688 (O_688,N_4792,N_4973);
nand UO_689 (O_689,N_4975,N_4699);
xor UO_690 (O_690,N_4500,N_4599);
nor UO_691 (O_691,N_4260,N_4203);
or UO_692 (O_692,N_4757,N_4991);
xnor UO_693 (O_693,N_4718,N_4189);
nand UO_694 (O_694,N_4238,N_4558);
and UO_695 (O_695,N_4127,N_4300);
and UO_696 (O_696,N_4710,N_4446);
xnor UO_697 (O_697,N_4749,N_4326);
nand UO_698 (O_698,N_4547,N_4467);
xor UO_699 (O_699,N_4713,N_4807);
or UO_700 (O_700,N_4342,N_4873);
nor UO_701 (O_701,N_4302,N_4012);
and UO_702 (O_702,N_4057,N_4989);
nand UO_703 (O_703,N_4275,N_4705);
nor UO_704 (O_704,N_4318,N_4130);
xor UO_705 (O_705,N_4748,N_4408);
xnor UO_706 (O_706,N_4266,N_4012);
and UO_707 (O_707,N_4894,N_4923);
xor UO_708 (O_708,N_4549,N_4369);
and UO_709 (O_709,N_4656,N_4858);
or UO_710 (O_710,N_4063,N_4517);
or UO_711 (O_711,N_4559,N_4707);
nor UO_712 (O_712,N_4032,N_4539);
nand UO_713 (O_713,N_4838,N_4525);
and UO_714 (O_714,N_4498,N_4733);
nand UO_715 (O_715,N_4111,N_4134);
and UO_716 (O_716,N_4454,N_4672);
or UO_717 (O_717,N_4869,N_4922);
nand UO_718 (O_718,N_4371,N_4162);
xor UO_719 (O_719,N_4566,N_4965);
nand UO_720 (O_720,N_4223,N_4754);
nor UO_721 (O_721,N_4462,N_4164);
or UO_722 (O_722,N_4575,N_4596);
nand UO_723 (O_723,N_4626,N_4087);
nor UO_724 (O_724,N_4763,N_4072);
or UO_725 (O_725,N_4349,N_4309);
nand UO_726 (O_726,N_4331,N_4346);
nor UO_727 (O_727,N_4595,N_4527);
or UO_728 (O_728,N_4056,N_4304);
or UO_729 (O_729,N_4623,N_4577);
xor UO_730 (O_730,N_4865,N_4022);
nor UO_731 (O_731,N_4441,N_4895);
or UO_732 (O_732,N_4839,N_4456);
and UO_733 (O_733,N_4596,N_4886);
or UO_734 (O_734,N_4438,N_4833);
xor UO_735 (O_735,N_4757,N_4356);
and UO_736 (O_736,N_4247,N_4282);
or UO_737 (O_737,N_4281,N_4921);
xnor UO_738 (O_738,N_4451,N_4949);
xnor UO_739 (O_739,N_4151,N_4593);
and UO_740 (O_740,N_4519,N_4748);
and UO_741 (O_741,N_4937,N_4348);
nand UO_742 (O_742,N_4875,N_4135);
xor UO_743 (O_743,N_4228,N_4386);
nor UO_744 (O_744,N_4943,N_4557);
and UO_745 (O_745,N_4377,N_4482);
xnor UO_746 (O_746,N_4660,N_4240);
or UO_747 (O_747,N_4731,N_4411);
nor UO_748 (O_748,N_4953,N_4732);
xor UO_749 (O_749,N_4505,N_4826);
and UO_750 (O_750,N_4769,N_4047);
or UO_751 (O_751,N_4948,N_4550);
or UO_752 (O_752,N_4517,N_4591);
or UO_753 (O_753,N_4012,N_4906);
nor UO_754 (O_754,N_4246,N_4806);
xor UO_755 (O_755,N_4085,N_4797);
nand UO_756 (O_756,N_4865,N_4351);
and UO_757 (O_757,N_4620,N_4253);
or UO_758 (O_758,N_4749,N_4470);
nand UO_759 (O_759,N_4532,N_4859);
or UO_760 (O_760,N_4380,N_4419);
nand UO_761 (O_761,N_4578,N_4120);
and UO_762 (O_762,N_4400,N_4195);
or UO_763 (O_763,N_4582,N_4325);
nand UO_764 (O_764,N_4333,N_4047);
nand UO_765 (O_765,N_4601,N_4117);
or UO_766 (O_766,N_4015,N_4735);
and UO_767 (O_767,N_4700,N_4428);
and UO_768 (O_768,N_4841,N_4501);
and UO_769 (O_769,N_4504,N_4474);
xor UO_770 (O_770,N_4805,N_4538);
or UO_771 (O_771,N_4041,N_4766);
nor UO_772 (O_772,N_4322,N_4519);
and UO_773 (O_773,N_4410,N_4891);
and UO_774 (O_774,N_4928,N_4920);
or UO_775 (O_775,N_4011,N_4876);
xor UO_776 (O_776,N_4724,N_4042);
or UO_777 (O_777,N_4559,N_4890);
or UO_778 (O_778,N_4753,N_4294);
and UO_779 (O_779,N_4565,N_4044);
nand UO_780 (O_780,N_4756,N_4997);
nor UO_781 (O_781,N_4732,N_4377);
nor UO_782 (O_782,N_4833,N_4151);
or UO_783 (O_783,N_4601,N_4306);
and UO_784 (O_784,N_4961,N_4239);
or UO_785 (O_785,N_4961,N_4035);
or UO_786 (O_786,N_4303,N_4117);
and UO_787 (O_787,N_4593,N_4673);
xnor UO_788 (O_788,N_4632,N_4973);
xor UO_789 (O_789,N_4687,N_4391);
or UO_790 (O_790,N_4027,N_4935);
and UO_791 (O_791,N_4716,N_4731);
nor UO_792 (O_792,N_4392,N_4312);
or UO_793 (O_793,N_4294,N_4301);
xor UO_794 (O_794,N_4585,N_4830);
nand UO_795 (O_795,N_4440,N_4656);
nor UO_796 (O_796,N_4019,N_4136);
and UO_797 (O_797,N_4335,N_4448);
nor UO_798 (O_798,N_4841,N_4174);
nand UO_799 (O_799,N_4373,N_4030);
xor UO_800 (O_800,N_4351,N_4954);
nand UO_801 (O_801,N_4049,N_4430);
or UO_802 (O_802,N_4354,N_4743);
nand UO_803 (O_803,N_4344,N_4975);
nor UO_804 (O_804,N_4434,N_4177);
or UO_805 (O_805,N_4518,N_4926);
or UO_806 (O_806,N_4623,N_4962);
nor UO_807 (O_807,N_4054,N_4243);
or UO_808 (O_808,N_4986,N_4533);
nor UO_809 (O_809,N_4392,N_4845);
and UO_810 (O_810,N_4643,N_4456);
and UO_811 (O_811,N_4677,N_4776);
and UO_812 (O_812,N_4349,N_4860);
or UO_813 (O_813,N_4170,N_4926);
xor UO_814 (O_814,N_4492,N_4093);
nor UO_815 (O_815,N_4956,N_4110);
nand UO_816 (O_816,N_4778,N_4365);
xor UO_817 (O_817,N_4267,N_4892);
and UO_818 (O_818,N_4090,N_4384);
nor UO_819 (O_819,N_4716,N_4271);
nor UO_820 (O_820,N_4407,N_4591);
or UO_821 (O_821,N_4006,N_4747);
xnor UO_822 (O_822,N_4795,N_4430);
nor UO_823 (O_823,N_4941,N_4872);
or UO_824 (O_824,N_4985,N_4134);
and UO_825 (O_825,N_4289,N_4356);
nand UO_826 (O_826,N_4888,N_4710);
nor UO_827 (O_827,N_4793,N_4187);
or UO_828 (O_828,N_4354,N_4457);
nand UO_829 (O_829,N_4888,N_4029);
nand UO_830 (O_830,N_4918,N_4061);
nor UO_831 (O_831,N_4927,N_4405);
xnor UO_832 (O_832,N_4890,N_4549);
or UO_833 (O_833,N_4156,N_4085);
and UO_834 (O_834,N_4720,N_4868);
and UO_835 (O_835,N_4486,N_4644);
nor UO_836 (O_836,N_4656,N_4541);
or UO_837 (O_837,N_4294,N_4631);
xnor UO_838 (O_838,N_4743,N_4783);
or UO_839 (O_839,N_4986,N_4303);
or UO_840 (O_840,N_4203,N_4933);
and UO_841 (O_841,N_4063,N_4194);
nor UO_842 (O_842,N_4540,N_4056);
xnor UO_843 (O_843,N_4406,N_4041);
or UO_844 (O_844,N_4756,N_4156);
nor UO_845 (O_845,N_4350,N_4604);
nand UO_846 (O_846,N_4279,N_4191);
nor UO_847 (O_847,N_4182,N_4485);
and UO_848 (O_848,N_4460,N_4898);
nor UO_849 (O_849,N_4661,N_4964);
nand UO_850 (O_850,N_4463,N_4997);
or UO_851 (O_851,N_4528,N_4044);
xor UO_852 (O_852,N_4604,N_4681);
nand UO_853 (O_853,N_4688,N_4666);
xnor UO_854 (O_854,N_4160,N_4116);
xnor UO_855 (O_855,N_4329,N_4127);
nor UO_856 (O_856,N_4056,N_4843);
xnor UO_857 (O_857,N_4519,N_4115);
nand UO_858 (O_858,N_4908,N_4460);
nor UO_859 (O_859,N_4466,N_4532);
or UO_860 (O_860,N_4379,N_4982);
and UO_861 (O_861,N_4831,N_4446);
and UO_862 (O_862,N_4636,N_4756);
or UO_863 (O_863,N_4114,N_4853);
nand UO_864 (O_864,N_4327,N_4367);
and UO_865 (O_865,N_4521,N_4827);
or UO_866 (O_866,N_4760,N_4856);
or UO_867 (O_867,N_4799,N_4061);
xnor UO_868 (O_868,N_4028,N_4069);
xor UO_869 (O_869,N_4581,N_4634);
xnor UO_870 (O_870,N_4105,N_4306);
or UO_871 (O_871,N_4712,N_4865);
and UO_872 (O_872,N_4637,N_4356);
xnor UO_873 (O_873,N_4646,N_4461);
nand UO_874 (O_874,N_4682,N_4223);
xnor UO_875 (O_875,N_4185,N_4438);
nand UO_876 (O_876,N_4156,N_4574);
or UO_877 (O_877,N_4723,N_4923);
nor UO_878 (O_878,N_4163,N_4833);
nand UO_879 (O_879,N_4211,N_4000);
nand UO_880 (O_880,N_4180,N_4924);
xnor UO_881 (O_881,N_4748,N_4005);
nand UO_882 (O_882,N_4098,N_4930);
nand UO_883 (O_883,N_4766,N_4713);
and UO_884 (O_884,N_4851,N_4326);
nand UO_885 (O_885,N_4071,N_4824);
nor UO_886 (O_886,N_4091,N_4545);
or UO_887 (O_887,N_4339,N_4525);
nand UO_888 (O_888,N_4161,N_4349);
nand UO_889 (O_889,N_4440,N_4885);
and UO_890 (O_890,N_4174,N_4750);
or UO_891 (O_891,N_4276,N_4950);
nor UO_892 (O_892,N_4416,N_4591);
and UO_893 (O_893,N_4111,N_4280);
or UO_894 (O_894,N_4714,N_4433);
and UO_895 (O_895,N_4128,N_4122);
nor UO_896 (O_896,N_4127,N_4174);
xnor UO_897 (O_897,N_4761,N_4786);
nor UO_898 (O_898,N_4404,N_4879);
nor UO_899 (O_899,N_4850,N_4884);
xor UO_900 (O_900,N_4552,N_4536);
or UO_901 (O_901,N_4755,N_4500);
nand UO_902 (O_902,N_4181,N_4859);
xnor UO_903 (O_903,N_4603,N_4864);
nor UO_904 (O_904,N_4635,N_4731);
xor UO_905 (O_905,N_4116,N_4010);
xnor UO_906 (O_906,N_4534,N_4643);
nand UO_907 (O_907,N_4624,N_4790);
nor UO_908 (O_908,N_4526,N_4613);
nor UO_909 (O_909,N_4543,N_4407);
xnor UO_910 (O_910,N_4629,N_4458);
xor UO_911 (O_911,N_4986,N_4907);
nor UO_912 (O_912,N_4563,N_4183);
nand UO_913 (O_913,N_4498,N_4085);
xor UO_914 (O_914,N_4952,N_4111);
or UO_915 (O_915,N_4502,N_4677);
nor UO_916 (O_916,N_4689,N_4278);
and UO_917 (O_917,N_4014,N_4489);
or UO_918 (O_918,N_4876,N_4228);
or UO_919 (O_919,N_4727,N_4711);
nand UO_920 (O_920,N_4593,N_4886);
nand UO_921 (O_921,N_4497,N_4652);
nor UO_922 (O_922,N_4149,N_4269);
nand UO_923 (O_923,N_4098,N_4203);
xor UO_924 (O_924,N_4312,N_4703);
and UO_925 (O_925,N_4828,N_4302);
nand UO_926 (O_926,N_4994,N_4121);
nand UO_927 (O_927,N_4856,N_4177);
and UO_928 (O_928,N_4245,N_4537);
or UO_929 (O_929,N_4513,N_4822);
nand UO_930 (O_930,N_4207,N_4978);
or UO_931 (O_931,N_4357,N_4719);
xnor UO_932 (O_932,N_4311,N_4225);
nand UO_933 (O_933,N_4493,N_4548);
xor UO_934 (O_934,N_4710,N_4687);
and UO_935 (O_935,N_4329,N_4931);
or UO_936 (O_936,N_4132,N_4747);
or UO_937 (O_937,N_4110,N_4416);
xnor UO_938 (O_938,N_4384,N_4983);
and UO_939 (O_939,N_4105,N_4620);
xor UO_940 (O_940,N_4329,N_4290);
nand UO_941 (O_941,N_4485,N_4666);
nand UO_942 (O_942,N_4428,N_4415);
nor UO_943 (O_943,N_4384,N_4408);
xnor UO_944 (O_944,N_4256,N_4558);
or UO_945 (O_945,N_4632,N_4961);
nand UO_946 (O_946,N_4988,N_4987);
nand UO_947 (O_947,N_4671,N_4680);
xor UO_948 (O_948,N_4489,N_4567);
or UO_949 (O_949,N_4635,N_4689);
xnor UO_950 (O_950,N_4427,N_4274);
nor UO_951 (O_951,N_4571,N_4102);
nor UO_952 (O_952,N_4665,N_4783);
or UO_953 (O_953,N_4767,N_4992);
nor UO_954 (O_954,N_4294,N_4309);
nand UO_955 (O_955,N_4081,N_4354);
xor UO_956 (O_956,N_4002,N_4823);
nor UO_957 (O_957,N_4626,N_4961);
or UO_958 (O_958,N_4732,N_4234);
xnor UO_959 (O_959,N_4521,N_4494);
or UO_960 (O_960,N_4350,N_4738);
xor UO_961 (O_961,N_4568,N_4201);
xor UO_962 (O_962,N_4773,N_4892);
and UO_963 (O_963,N_4245,N_4434);
and UO_964 (O_964,N_4473,N_4431);
xor UO_965 (O_965,N_4056,N_4712);
xnor UO_966 (O_966,N_4719,N_4847);
nand UO_967 (O_967,N_4745,N_4609);
or UO_968 (O_968,N_4500,N_4472);
and UO_969 (O_969,N_4497,N_4918);
or UO_970 (O_970,N_4211,N_4312);
or UO_971 (O_971,N_4496,N_4805);
xnor UO_972 (O_972,N_4191,N_4682);
xor UO_973 (O_973,N_4229,N_4322);
xnor UO_974 (O_974,N_4789,N_4942);
or UO_975 (O_975,N_4667,N_4303);
nor UO_976 (O_976,N_4340,N_4543);
or UO_977 (O_977,N_4421,N_4203);
and UO_978 (O_978,N_4815,N_4132);
nand UO_979 (O_979,N_4206,N_4053);
or UO_980 (O_980,N_4774,N_4015);
nand UO_981 (O_981,N_4220,N_4979);
nand UO_982 (O_982,N_4805,N_4734);
and UO_983 (O_983,N_4124,N_4143);
nand UO_984 (O_984,N_4793,N_4718);
and UO_985 (O_985,N_4162,N_4599);
nor UO_986 (O_986,N_4528,N_4927);
nor UO_987 (O_987,N_4024,N_4246);
nand UO_988 (O_988,N_4329,N_4203);
nor UO_989 (O_989,N_4560,N_4866);
xor UO_990 (O_990,N_4961,N_4576);
nand UO_991 (O_991,N_4498,N_4904);
xor UO_992 (O_992,N_4387,N_4234);
xnor UO_993 (O_993,N_4411,N_4755);
or UO_994 (O_994,N_4503,N_4957);
nand UO_995 (O_995,N_4746,N_4606);
and UO_996 (O_996,N_4807,N_4736);
nor UO_997 (O_997,N_4656,N_4929);
or UO_998 (O_998,N_4437,N_4460);
nand UO_999 (O_999,N_4382,N_4957);
endmodule