module basic_2000_20000_2500_5_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_326,In_246);
or U1 (N_1,In_1662,In_863);
or U2 (N_2,In_1367,In_192);
and U3 (N_3,In_1928,In_1444);
and U4 (N_4,In_378,In_1863);
or U5 (N_5,In_617,In_696);
nor U6 (N_6,In_751,In_970);
and U7 (N_7,In_972,In_1113);
and U8 (N_8,In_1800,In_1703);
or U9 (N_9,In_1165,In_1514);
nor U10 (N_10,In_231,In_1116);
and U11 (N_11,In_221,In_372);
or U12 (N_12,In_758,In_1555);
nand U13 (N_13,In_155,In_44);
nor U14 (N_14,In_8,In_195);
and U15 (N_15,In_1437,In_1280);
nor U16 (N_16,In_1756,In_1550);
nor U17 (N_17,In_1733,In_1343);
nor U18 (N_18,In_1978,In_1193);
nand U19 (N_19,In_1168,In_214);
nand U20 (N_20,In_1472,In_1545);
nor U21 (N_21,In_1719,In_295);
nor U22 (N_22,In_1519,In_1335);
and U23 (N_23,In_936,In_1096);
and U24 (N_24,In_518,In_1005);
and U25 (N_25,In_1143,In_289);
and U26 (N_26,In_1612,In_942);
or U27 (N_27,In_62,In_1638);
and U28 (N_28,In_186,In_1288);
and U29 (N_29,In_1021,In_908);
and U30 (N_30,In_179,In_678);
nand U31 (N_31,In_69,In_1776);
and U32 (N_32,In_1236,In_947);
or U33 (N_33,In_495,In_755);
or U34 (N_34,In_309,In_1407);
nor U35 (N_35,In_1643,In_1907);
or U36 (N_36,In_375,In_1506);
nand U37 (N_37,In_240,In_361);
and U38 (N_38,In_586,In_172);
or U39 (N_39,In_565,In_549);
or U40 (N_40,In_1974,In_409);
and U41 (N_41,In_774,In_1516);
nand U42 (N_42,In_508,In_1380);
nand U43 (N_43,In_94,In_1793);
or U44 (N_44,In_1631,In_184);
nand U45 (N_45,In_1402,In_1255);
and U46 (N_46,In_1805,In_122);
and U47 (N_47,In_1994,In_895);
nor U48 (N_48,In_1853,In_502);
and U49 (N_49,In_1215,In_1948);
or U50 (N_50,In_29,In_1028);
nand U51 (N_51,In_350,In_1169);
and U52 (N_52,In_1995,In_1956);
nand U53 (N_53,In_1504,In_1349);
and U54 (N_54,In_1518,In_1358);
or U55 (N_55,In_1864,In_120);
and U56 (N_56,In_1850,In_864);
nand U57 (N_57,In_1441,In_399);
nor U58 (N_58,In_1770,In_852);
and U59 (N_59,In_4,In_695);
nor U60 (N_60,In_1617,In_1909);
nor U61 (N_61,In_1466,In_1321);
nor U62 (N_62,In_445,In_1557);
nor U63 (N_63,In_486,In_880);
or U64 (N_64,In_1831,In_1128);
or U65 (N_65,In_1526,In_1977);
or U66 (N_66,In_888,In_435);
nand U67 (N_67,In_89,In_1999);
nand U68 (N_68,In_848,In_1090);
nor U69 (N_69,In_1099,In_1212);
and U70 (N_70,In_1010,In_1339);
nand U71 (N_71,In_446,In_278);
nand U72 (N_72,In_1286,In_1320);
nor U73 (N_73,In_1283,In_635);
nand U74 (N_74,In_836,In_690);
nor U75 (N_75,In_557,In_978);
and U76 (N_76,In_1947,In_649);
or U77 (N_77,In_1972,In_272);
and U78 (N_78,In_1211,In_979);
nor U79 (N_79,In_1259,In_1884);
and U80 (N_80,In_1826,In_337);
nand U81 (N_81,In_780,In_1369);
or U82 (N_82,In_1779,In_1690);
nor U83 (N_83,In_1936,In_1993);
or U84 (N_84,In_311,In_1803);
and U85 (N_85,In_788,In_753);
and U86 (N_86,In_775,In_870);
and U87 (N_87,In_664,In_607);
and U88 (N_88,In_1250,In_1591);
nor U89 (N_89,In_1051,In_1954);
nand U90 (N_90,In_815,In_1757);
or U91 (N_91,In_450,In_702);
nand U92 (N_92,In_1448,In_1158);
and U93 (N_93,In_1953,In_1450);
and U94 (N_94,In_532,In_1091);
nand U95 (N_95,In_1934,In_1804);
and U96 (N_96,In_21,In_488);
and U97 (N_97,In_1963,In_1474);
nand U98 (N_98,In_1299,In_73);
and U99 (N_99,In_1938,In_1937);
nand U100 (N_100,In_1132,In_1063);
nor U101 (N_101,In_505,In_338);
nor U102 (N_102,In_945,In_657);
nand U103 (N_103,In_735,In_687);
nor U104 (N_104,In_1411,In_193);
and U105 (N_105,In_1133,In_1812);
nor U106 (N_106,In_354,In_397);
or U107 (N_107,In_1911,In_1011);
and U108 (N_108,In_468,In_307);
and U109 (N_109,In_1950,In_1538);
and U110 (N_110,In_1752,In_1943);
or U111 (N_111,In_1007,In_1510);
or U112 (N_112,In_1528,In_628);
nor U113 (N_113,In_248,In_1404);
or U114 (N_114,In_1961,In_982);
and U115 (N_115,In_1082,In_1723);
or U116 (N_116,In_1058,In_566);
nand U117 (N_117,In_779,In_1055);
or U118 (N_118,In_226,In_1279);
nor U119 (N_119,In_104,In_1302);
nor U120 (N_120,In_238,In_697);
xor U121 (N_121,In_1983,In_1262);
and U122 (N_122,In_991,In_1544);
nor U123 (N_123,In_1768,In_749);
nand U124 (N_124,In_453,In_461);
or U125 (N_125,In_595,In_829);
and U126 (N_126,In_646,In_669);
or U127 (N_127,In_1126,In_1080);
nor U128 (N_128,In_538,In_904);
or U129 (N_129,In_1606,In_777);
or U130 (N_130,In_475,In_1248);
nor U131 (N_131,In_1728,In_1289);
nand U132 (N_132,In_1013,In_1271);
nand U133 (N_133,In_1334,In_675);
or U134 (N_134,In_773,In_1137);
or U135 (N_135,In_82,In_1340);
nand U136 (N_136,In_203,In_1316);
nor U137 (N_137,In_1813,In_212);
nor U138 (N_138,In_1773,In_443);
nor U139 (N_139,In_1613,In_529);
nor U140 (N_140,In_583,In_1049);
or U141 (N_141,In_16,In_898);
nor U142 (N_142,In_858,In_1186);
or U143 (N_143,In_1342,In_1527);
nor U144 (N_144,In_1741,In_199);
or U145 (N_145,In_967,In_401);
nand U146 (N_146,In_403,In_1681);
nor U147 (N_147,In_466,In_712);
or U148 (N_148,In_1529,In_660);
nor U149 (N_149,In_1860,In_1691);
nand U150 (N_150,In_499,In_624);
or U151 (N_151,In_1246,In_1724);
nor U152 (N_152,In_1144,In_1692);
nand U153 (N_153,In_1251,In_490);
and U154 (N_154,In_1480,In_759);
or U155 (N_155,In_1446,In_1136);
or U156 (N_156,In_421,In_1878);
or U157 (N_157,In_1365,In_1890);
nand U158 (N_158,In_988,In_556);
nand U159 (N_159,In_1685,In_54);
and U160 (N_160,In_1118,In_1241);
or U161 (N_161,In_1354,In_1688);
and U162 (N_162,In_658,In_1743);
or U163 (N_163,In_1027,In_1540);
nor U164 (N_164,In_1849,In_390);
nor U165 (N_165,In_552,In_318);
or U166 (N_166,In_1541,In_921);
nor U167 (N_167,In_140,In_23);
nand U168 (N_168,In_129,In_1440);
nor U169 (N_169,In_816,In_1451);
or U170 (N_170,In_564,In_335);
nor U171 (N_171,In_1227,In_1081);
nand U172 (N_172,In_1755,In_1357);
or U173 (N_173,In_30,In_533);
nand U174 (N_174,In_1257,In_285);
or U175 (N_175,In_1157,In_1314);
nor U176 (N_176,In_1231,In_507);
nand U177 (N_177,In_1270,In_463);
nor U178 (N_178,In_183,In_720);
nand U179 (N_179,In_290,In_1984);
and U180 (N_180,In_596,In_1356);
nor U181 (N_181,In_1325,In_721);
nand U182 (N_182,In_1817,In_1846);
or U183 (N_183,In_43,In_756);
nor U184 (N_184,In_344,In_456);
and U185 (N_185,In_688,In_1892);
or U186 (N_186,In_914,In_1115);
nand U187 (N_187,In_86,In_416);
nand U188 (N_188,In_1195,In_1475);
nor U189 (N_189,In_739,In_151);
nor U190 (N_190,In_177,In_276);
nor U191 (N_191,In_1677,In_75);
nand U192 (N_192,In_1558,In_95);
or U193 (N_193,In_152,In_431);
or U194 (N_194,In_230,In_1597);
nor U195 (N_195,In_1203,In_1525);
nand U196 (N_196,In_180,In_1881);
nand U197 (N_197,In_189,In_31);
or U198 (N_198,In_1867,In_157);
nor U199 (N_199,In_1784,In_642);
and U200 (N_200,In_1180,In_551);
and U201 (N_201,In_725,In_1245);
and U202 (N_202,In_1263,In_79);
and U203 (N_203,In_724,In_1431);
or U204 (N_204,In_971,In_1998);
nor U205 (N_205,In_1019,In_249);
and U206 (N_206,In_958,In_1744);
and U207 (N_207,In_1652,In_1228);
and U208 (N_208,In_1734,In_1276);
or U209 (N_209,In_763,In_1389);
nor U210 (N_210,In_578,In_822);
and U211 (N_211,In_1832,In_917);
nor U212 (N_212,In_1306,In_55);
or U213 (N_213,In_118,In_1700);
and U214 (N_214,In_821,In_101);
nor U215 (N_215,In_804,In_1249);
nor U216 (N_216,In_209,In_339);
nand U217 (N_217,In_1374,In_317);
and U218 (N_218,In_679,In_1513);
and U219 (N_219,In_1587,In_1442);
nand U220 (N_220,In_1584,In_374);
nor U221 (N_221,In_392,In_433);
and U222 (N_222,In_1798,In_977);
nor U223 (N_223,In_1054,In_410);
or U224 (N_224,In_668,In_1789);
nor U225 (N_225,In_1877,In_14);
nand U226 (N_226,In_1064,In_1347);
nand U227 (N_227,In_300,In_90);
nand U228 (N_228,In_1478,In_1944);
and U229 (N_229,In_912,In_99);
nand U230 (N_230,In_386,In_1346);
nand U231 (N_231,In_1646,In_1657);
nor U232 (N_232,In_893,In_950);
or U233 (N_233,In_1712,In_402);
nor U234 (N_234,In_676,In_1223);
or U235 (N_235,In_555,In_1778);
nor U236 (N_236,In_1102,In_1199);
nand U237 (N_237,In_1598,In_839);
nor U238 (N_238,In_1722,In_652);
and U239 (N_239,In_1,In_185);
nor U240 (N_240,In_49,In_757);
nand U241 (N_241,In_851,In_1517);
and U242 (N_242,In_738,In_1568);
nor U243 (N_243,In_1390,In_857);
nor U244 (N_244,In_1239,In_1261);
nand U245 (N_245,In_287,In_1185);
or U246 (N_246,In_274,In_585);
nand U247 (N_247,In_283,In_1145);
nor U248 (N_248,In_778,In_472);
xor U249 (N_249,In_277,In_1704);
or U250 (N_250,In_281,In_449);
nand U251 (N_251,In_517,In_1611);
nand U252 (N_252,In_882,In_535);
nand U253 (N_253,In_813,In_754);
or U254 (N_254,In_1196,In_1275);
and U255 (N_255,In_1505,In_1896);
and U256 (N_256,In_1014,In_327);
nand U257 (N_257,In_1273,In_783);
and U258 (N_258,In_236,In_1083);
nand U259 (N_259,In_35,In_553);
nand U260 (N_260,In_770,In_726);
nor U261 (N_261,In_37,In_953);
and U262 (N_262,In_1312,In_530);
nand U263 (N_263,In_1731,In_1674);
or U264 (N_264,In_342,In_1658);
nor U265 (N_265,In_1848,In_875);
and U266 (N_266,In_131,In_1109);
nor U267 (N_267,In_1492,In_1368);
nor U268 (N_268,In_503,In_1176);
or U269 (N_269,In_1989,In_667);
nand U270 (N_270,In_868,In_434);
or U271 (N_271,In_1701,In_407);
and U272 (N_272,In_1040,In_292);
nand U273 (N_273,In_1809,In_1351);
or U274 (N_274,In_1205,In_1840);
nand U275 (N_275,In_588,In_1426);
or U276 (N_276,In_1112,In_860);
or U277 (N_277,In_218,In_174);
or U278 (N_278,In_1588,In_641);
and U279 (N_279,In_1471,In_576);
nand U280 (N_280,In_216,In_371);
and U281 (N_281,In_1775,In_792);
nand U282 (N_282,In_250,In_1068);
or U283 (N_283,In_634,In_1315);
or U284 (N_284,In_1060,In_1511);
and U285 (N_285,In_786,In_886);
nor U286 (N_286,In_1037,In_969);
nand U287 (N_287,In_1069,In_485);
nand U288 (N_288,In_1659,In_255);
nor U289 (N_289,In_1094,In_332);
or U290 (N_290,In_1689,In_1332);
and U291 (N_291,In_519,In_479);
nor U292 (N_292,In_437,In_1379);
nor U293 (N_293,In_1981,In_981);
or U294 (N_294,In_427,In_510);
nand U295 (N_295,In_831,In_1206);
or U296 (N_296,In_1683,In_1162);
and U297 (N_297,In_1650,In_18);
nor U298 (N_298,In_191,In_671);
nand U299 (N_299,In_484,In_1164);
nor U300 (N_300,In_1484,In_208);
and U301 (N_301,In_83,In_1243);
nor U302 (N_302,In_1745,In_1030);
and U303 (N_303,In_415,In_683);
nor U304 (N_304,In_280,In_1819);
nand U305 (N_305,In_1429,In_1012);
and U306 (N_306,In_1695,In_1059);
nor U307 (N_307,In_353,In_1119);
nor U308 (N_308,In_308,In_973);
nor U309 (N_309,In_1560,In_1464);
nand U310 (N_310,In_1496,In_493);
nor U311 (N_311,In_347,In_1101);
nand U312 (N_312,In_1194,In_232);
or U313 (N_313,In_1421,In_1352);
nor U314 (N_314,In_1532,In_1048);
and U315 (N_315,In_355,In_938);
nand U316 (N_316,In_284,In_1171);
xor U317 (N_317,In_570,In_1163);
nand U318 (N_318,In_1238,In_1990);
nor U319 (N_319,In_1893,In_213);
and U320 (N_320,In_1216,In_1763);
and U321 (N_321,In_1406,In_614);
and U322 (N_322,In_1190,In_1057);
nand U323 (N_323,In_1660,In_672);
nor U324 (N_324,In_699,In_1876);
and U325 (N_325,In_264,In_1781);
or U326 (N_326,In_3,In_1873);
nor U327 (N_327,In_247,In_733);
nand U328 (N_328,In_793,In_1417);
nor U329 (N_329,In_491,In_1183);
and U330 (N_330,In_741,In_1601);
nand U331 (N_331,In_316,In_1648);
nor U332 (N_332,In_542,In_1891);
or U333 (N_333,In_647,In_748);
nand U334 (N_334,In_418,In_385);
or U335 (N_335,In_1655,In_873);
or U336 (N_336,In_306,In_1329);
nor U337 (N_337,In_1780,In_653);
and U338 (N_338,In_275,In_145);
or U339 (N_339,In_245,In_1868);
nor U340 (N_340,In_1430,In_698);
and U341 (N_341,In_1697,In_258);
nand U342 (N_342,In_92,In_1327);
nand U343 (N_343,In_1495,In_1710);
nand U344 (N_344,In_1543,In_382);
nand U345 (N_345,In_1201,In_1220);
xor U346 (N_346,In_834,In_1488);
xor U347 (N_347,In_896,In_1034);
and U348 (N_348,In_1303,In_1684);
xor U349 (N_349,In_124,In_293);
nand U350 (N_350,In_1419,In_525);
or U351 (N_351,In_1285,In_128);
nand U352 (N_352,In_1139,In_1141);
nor U353 (N_353,In_271,In_1151);
or U354 (N_354,In_810,In_643);
nor U355 (N_355,In_1622,In_1375);
or U356 (N_356,In_1160,In_1820);
nor U357 (N_357,In_581,In_1318);
and U358 (N_358,In_1284,In_1341);
nor U359 (N_359,In_1535,In_1859);
and U360 (N_360,In_1256,In_462);
nor U361 (N_361,In_1487,In_1654);
or U362 (N_362,In_1815,In_1782);
or U363 (N_363,In_539,In_1788);
nor U364 (N_364,In_1265,In_476);
and U365 (N_365,In_1297,In_1260);
or U366 (N_366,In_865,In_1138);
nor U367 (N_367,In_1629,In_1479);
nor U368 (N_368,In_637,In_655);
or U369 (N_369,In_575,In_910);
and U370 (N_370,In_454,In_706);
and U371 (N_371,In_1642,In_1580);
or U372 (N_372,In_808,In_891);
and U373 (N_373,In_1906,In_200);
and U374 (N_374,In_1415,In_1175);
or U375 (N_375,In_1627,In_1089);
nand U376 (N_376,In_425,In_36);
nand U377 (N_377,In_951,In_32);
nand U378 (N_378,In_871,In_964);
nor U379 (N_379,In_1301,In_1494);
nand U380 (N_380,In_522,In_1720);
nor U381 (N_381,In_1777,In_1871);
or U382 (N_382,In_805,In_1004);
or U383 (N_383,In_494,In_176);
nand U384 (N_384,In_546,In_13);
or U385 (N_385,In_88,In_639);
nor U386 (N_386,In_794,In_405);
and U387 (N_387,In_1264,In_610);
xor U388 (N_388,In_253,In_998);
and U389 (N_389,In_141,In_2);
nand U390 (N_390,In_601,In_1951);
nand U391 (N_391,In_1836,In_1213);
and U392 (N_392,In_1581,In_1845);
xnor U393 (N_393,In_789,In_963);
nand U394 (N_394,In_561,In_1470);
or U395 (N_395,In_1072,In_1465);
and U396 (N_396,In_666,In_1758);
or U397 (N_397,In_46,In_1575);
or U398 (N_398,In_1108,In_1949);
nor U399 (N_399,In_121,In_638);
and U400 (N_400,In_708,In_731);
or U401 (N_401,In_844,In_1338);
nor U402 (N_402,In_1491,In_112);
xor U403 (N_403,In_67,In_1856);
nand U404 (N_404,In_340,In_1025);
nor U405 (N_405,In_931,In_243);
nor U406 (N_406,In_1387,In_1436);
nor U407 (N_407,In_1905,In_147);
or U408 (N_408,In_1097,In_1708);
nand U409 (N_409,In_826,In_1459);
and U410 (N_410,In_1915,In_824);
or U411 (N_411,In_1399,In_1336);
nand U412 (N_412,In_1134,In_1563);
nor U413 (N_413,In_1391,In_33);
and U414 (N_414,In_881,In_1578);
nor U415 (N_415,In_441,In_336);
or U416 (N_416,In_1556,In_182);
nand U417 (N_417,In_1149,In_9);
and U418 (N_418,In_1490,In_1571);
or U419 (N_419,In_215,In_84);
nor U420 (N_420,In_1585,In_1696);
nand U421 (N_421,In_1140,In_159);
or U422 (N_422,In_384,In_1620);
nand U423 (N_423,In_1110,In_1530);
nand U424 (N_424,In_734,In_932);
or U425 (N_425,In_1675,In_1707);
and U426 (N_426,In_659,In_1500);
and U427 (N_427,In_1353,In_1566);
or U428 (N_428,In_990,In_1308);
or U429 (N_429,In_1412,In_1795);
and U430 (N_430,In_288,In_1326);
nand U431 (N_431,In_220,In_961);
nand U432 (N_432,In_1278,In_985);
and U433 (N_433,In_1766,In_1769);
nand U434 (N_434,In_577,In_388);
or U435 (N_435,In_429,In_1502);
xor U436 (N_436,In_1449,In_887);
nor U437 (N_437,In_1420,In_345);
and U438 (N_438,In_1287,In_438);
nor U439 (N_439,In_878,In_791);
nand U440 (N_440,In_470,In_618);
nand U441 (N_441,In_228,In_1957);
or U442 (N_442,In_1632,In_1754);
nand U443 (N_443,In_1737,In_1862);
nand U444 (N_444,In_1425,In_569);
nor U445 (N_445,In_714,In_1837);
or U446 (N_446,In_1125,In_732);
xnor U447 (N_447,In_352,In_1123);
nor U448 (N_448,In_291,In_1384);
nor U449 (N_449,In_536,In_843);
and U450 (N_450,In_795,In_1046);
nand U451 (N_451,In_611,In_477);
and U452 (N_452,In_1774,In_259);
nand U453 (N_453,In_541,In_136);
nand U454 (N_454,In_498,In_682);
nand U455 (N_455,In_605,In_930);
or U456 (N_456,In_521,In_820);
and U457 (N_457,In_323,In_959);
and U458 (N_458,In_1574,In_704);
nor U459 (N_459,In_1047,In_1053);
xor U460 (N_460,In_919,In_509);
nand U461 (N_461,In_1033,In_833);
nor U462 (N_462,In_640,In_606);
and U463 (N_463,In_856,In_513);
nand U464 (N_464,In_764,In_1237);
and U465 (N_465,In_1266,In_1965);
or U466 (N_466,In_1960,In_1721);
and U467 (N_467,In_257,In_114);
and U468 (N_468,In_1608,In_568);
and U469 (N_469,In_1344,In_52);
nand U470 (N_470,In_1888,In_1570);
or U471 (N_471,In_548,In_853);
or U472 (N_472,In_346,In_673);
nand U473 (N_473,In_97,In_139);
nand U474 (N_474,In_1135,In_162);
and U475 (N_475,In_1427,In_370);
or U476 (N_476,In_400,In_394);
nand U477 (N_477,In_1386,In_1857);
or U478 (N_478,In_330,In_1935);
nand U479 (N_479,In_650,In_357);
nor U480 (N_480,In_782,In_1640);
nand U481 (N_481,In_432,In_273);
nor U482 (N_482,In_527,In_1976);
or U483 (N_483,In_1087,In_913);
and U484 (N_484,In_1618,In_436);
nor U485 (N_485,In_567,In_572);
nand U486 (N_486,In_1489,In_1067);
xnor U487 (N_487,In_497,In_861);
nor U488 (N_488,In_482,In_1866);
nand U489 (N_489,In_1838,In_1825);
nand U490 (N_490,In_906,In_71);
and U491 (N_491,In_1727,In_1467);
nor U492 (N_492,In_1032,In_1003);
nor U493 (N_493,In_730,In_1673);
nor U494 (N_494,In_107,In_173);
nor U495 (N_495,In_1894,In_1930);
or U496 (N_496,In_465,In_1071);
and U497 (N_497,In_1039,In_1625);
or U498 (N_498,In_1373,In_1503);
nor U499 (N_499,In_1483,In_1024);
nor U500 (N_500,In_1207,In_1967);
nand U501 (N_501,In_1572,In_1305);
and U502 (N_502,In_902,In_1932);
nor U503 (N_503,In_181,In_1940);
nand U504 (N_504,In_1322,In_1875);
nor U505 (N_505,In_1523,In_262);
or U506 (N_506,In_677,In_1969);
and U507 (N_507,In_812,In_1605);
or U508 (N_508,In_1586,In_686);
or U509 (N_509,In_458,In_1253);
or U510 (N_510,In_1594,In_711);
and U511 (N_511,In_137,In_1787);
nand U512 (N_512,In_1188,In_1056);
and U513 (N_513,In_1913,In_1740);
nand U514 (N_514,In_545,In_223);
nand U515 (N_515,In_106,In_68);
and U516 (N_516,In_1653,In_85);
nand U517 (N_517,In_1309,In_268);
nand U518 (N_518,In_662,In_0);
or U519 (N_519,In_1124,In_1668);
nand U520 (N_520,In_1822,In_827);
nand U521 (N_521,In_471,In_1214);
and U522 (N_522,In_1699,In_1360);
or U523 (N_523,In_705,In_1786);
nand U524 (N_524,In_1022,In_1564);
nand U525 (N_525,In_322,In_1942);
and U526 (N_526,In_1394,In_623);
and U527 (N_527,In_1918,In_558);
nor U528 (N_528,In_64,In_1310);
nand U529 (N_529,In_1762,In_781);
nand U530 (N_530,In_1747,In_1842);
nor U531 (N_531,In_630,In_1924);
nand U532 (N_532,In_1222,In_1240);
nor U533 (N_533,In_138,In_772);
and U534 (N_534,In_1290,In_63);
and U535 (N_535,In_983,In_1554);
and U536 (N_536,In_1463,In_1392);
nor U537 (N_537,In_603,In_362);
nand U538 (N_538,In_1403,In_524);
and U539 (N_539,In_1593,In_1882);
nor U540 (N_540,In_1590,In_966);
or U541 (N_541,In_1709,In_1964);
and U542 (N_542,In_765,In_1823);
and U543 (N_543,In_1732,In_1679);
and U544 (N_544,In_1084,In_574);
or U545 (N_545,In_747,In_1439);
and U546 (N_546,In_211,In_1966);
or U547 (N_547,In_1282,In_965);
and U548 (N_548,In_1105,In_997);
and U549 (N_549,In_260,In_837);
nor U550 (N_550,In_1904,In_100);
nand U551 (N_551,In_252,In_360);
nand U552 (N_552,In_158,In_602);
nor U553 (N_553,In_1562,In_1899);
nor U554 (N_554,In_313,In_1066);
nand U555 (N_555,In_133,In_1567);
nor U556 (N_556,In_34,In_1268);
or U557 (N_557,In_1742,In_1725);
nand U558 (N_558,In_263,In_866);
nor U559 (N_559,In_654,In_1156);
nor U560 (N_560,In_1885,In_742);
or U561 (N_561,In_1476,In_80);
nor U562 (N_562,In_188,In_10);
or U563 (N_563,In_1453,In_796);
nand U564 (N_564,In_1897,In_661);
nor U565 (N_565,In_1687,In_366);
nor U566 (N_566,In_1117,In_743);
and U567 (N_567,In_1916,In_1274);
or U568 (N_568,In_903,In_1985);
or U569 (N_569,In_455,In_1433);
nand U570 (N_570,In_976,In_343);
nor U571 (N_571,In_113,In_633);
nor U572 (N_572,In_60,In_1962);
nand U573 (N_573,In_164,In_1364);
xor U574 (N_574,In_1718,In_1008);
or U575 (N_575,In_1045,In_1801);
nand U576 (N_576,In_1493,In_1317);
or U577 (N_577,In_1661,In_66);
nor U578 (N_578,In_1676,In_1456);
xor U579 (N_579,In_1414,In_1621);
or U580 (N_580,In_412,In_1189);
and U581 (N_581,In_1077,In_430);
nand U582 (N_582,In_1179,In_924);
and U583 (N_583,In_1736,In_1559);
and U584 (N_584,In_1361,In_1706);
or U585 (N_585,In_1172,In_1912);
nand U586 (N_586,In_1079,In_261);
or U587 (N_587,In_1821,In_1095);
or U588 (N_588,In_1150,In_175);
nand U589 (N_589,In_1771,In_562);
nand U590 (N_590,In_1886,In_1292);
or U591 (N_591,In_876,In_1148);
or U592 (N_592,In_954,In_1383);
nand U593 (N_593,In_198,In_61);
and U594 (N_594,In_1738,In_229);
or U595 (N_595,In_1184,In_1536);
nor U596 (N_596,In_1802,In_986);
nand U597 (N_597,In_644,In_1553);
or U598 (N_598,In_480,In_1486);
nor U599 (N_599,In_819,In_1350);
nand U600 (N_600,In_1166,In_1997);
nand U601 (N_601,In_636,In_25);
nor U602 (N_602,In_593,In_920);
nand U603 (N_603,In_626,In_879);
and U604 (N_604,In_874,In_1577);
and U605 (N_605,In_1042,In_803);
and U606 (N_606,In_41,In_1705);
nor U607 (N_607,In_1036,In_1626);
nand U608 (N_608,In_1120,In_892);
or U609 (N_609,In_943,In_974);
or U610 (N_610,In_608,In_926);
or U611 (N_611,In_356,In_1889);
nand U612 (N_612,In_840,In_42);
nand U613 (N_613,In_1232,In_1376);
nor U614 (N_614,In_933,In_1931);
and U615 (N_615,In_785,In_526);
nand U616 (N_616,In_674,In_980);
nand U617 (N_617,In_984,In_1619);
or U618 (N_618,In_1362,In_1711);
and U619 (N_619,In_1573,In_841);
nor U620 (N_620,In_1542,In_1610);
and U621 (N_621,In_110,In_1378);
and U622 (N_622,In_269,In_367);
nand U623 (N_623,In_1816,In_1609);
and U624 (N_624,In_1923,In_1469);
nand U625 (N_625,In_1018,In_1854);
nor U626 (N_626,In_116,In_736);
nand U627 (N_627,In_414,In_65);
or U628 (N_628,In_1630,In_492);
or U629 (N_629,In_1405,In_149);
nand U630 (N_630,In_74,In_1423);
nand U631 (N_631,In_349,In_227);
nor U632 (N_632,In_1127,In_1624);
nor U633 (N_633,In_1921,In_7);
nand U634 (N_634,In_746,In_718);
nor U635 (N_635,In_537,In_762);
nor U636 (N_636,In_1507,In_1726);
nand U637 (N_637,In_469,In_1749);
nand U638 (N_638,In_365,In_1114);
and U639 (N_639,In_1035,In_1395);
nand U640 (N_640,In_1254,In_160);
and U641 (N_641,In_50,In_222);
or U642 (N_642,In_1398,In_1422);
nand U643 (N_643,In_302,In_444);
and U644 (N_644,In_776,In_1167);
or U645 (N_645,In_811,In_1551);
and U646 (N_646,In_1945,In_1682);
nor U647 (N_647,In_1808,In_1970);
and U648 (N_648,In_1473,In_251);
nand U649 (N_649,In_1225,In_1767);
or U650 (N_650,In_1869,In_1130);
nor U651 (N_651,In_1901,In_1015);
nand U652 (N_652,In_922,In_1764);
or U653 (N_653,In_719,In_1634);
nor U654 (N_654,In_1293,In_1900);
nand U655 (N_655,In_171,In_1669);
nand U656 (N_656,In_125,In_885);
nor U657 (N_657,In_1359,In_800);
nor U658 (N_658,In_1111,In_478);
nor U659 (N_659,In_391,In_1050);
or U660 (N_660,In_729,In_506);
nor U661 (N_661,In_1182,In_379);
nor U662 (N_662,In_167,In_286);
nand U663 (N_663,In_481,In_1192);
nand U664 (N_664,In_684,In_341);
or U665 (N_665,In_1649,In_814);
and U666 (N_666,In_752,In_123);
or U667 (N_667,In_1922,In_225);
or U668 (N_668,In_111,In_282);
nand U669 (N_669,In_761,In_1461);
and U670 (N_670,In_1370,In_426);
nand U671 (N_671,In_832,In_501);
and U672 (N_672,In_767,In_884);
nor U673 (N_673,In_383,In_1714);
nor U674 (N_674,In_559,In_1468);
nor U675 (N_675,In_1142,In_1129);
or U676 (N_676,In_897,In_1765);
or U677 (N_677,In_1281,In_534);
and U678 (N_678,In_621,In_314);
and U679 (N_679,In_146,In_1515);
and U680 (N_680,In_398,In_1843);
nand U681 (N_681,In_1497,In_1397);
and U682 (N_682,In_1818,In_1103);
nand U683 (N_683,In_905,In_87);
nor U684 (N_684,In_1267,In_1746);
nand U685 (N_685,In_952,In_1509);
nor U686 (N_686,In_740,In_1001);
nand U687 (N_687,In_1547,In_1686);
or U688 (N_688,In_81,In_1191);
nand U689 (N_689,In_594,In_1908);
and U690 (N_690,In_1592,In_1952);
or U691 (N_691,In_1366,In_119);
or U692 (N_692,In_270,In_1671);
nor U693 (N_693,In_487,In_520);
nor U694 (N_694,In_1107,In_150);
nand U695 (N_695,In_835,In_987);
and U696 (N_696,In_395,In_1226);
and U697 (N_697,In_1477,In_1017);
and U698 (N_698,In_1992,In_818);
nor U699 (N_699,In_1428,In_1987);
nand U700 (N_700,In_911,In_651);
or U701 (N_701,In_1811,In_1539);
or U702 (N_702,In_992,In_955);
nand U703 (N_703,In_937,In_1796);
nor U704 (N_704,In_1919,In_877);
nor U705 (N_705,In_1401,In_294);
or U706 (N_706,In_528,In_242);
nand U707 (N_707,In_103,In_364);
nand U708 (N_708,In_154,In_523);
nand U709 (N_709,In_927,In_1152);
nor U710 (N_710,In_1807,In_889);
or U711 (N_711,In_254,In_1667);
and U712 (N_712,In_1300,In_1061);
nor U713 (N_713,In_801,In_1865);
and U714 (N_714,In_516,In_700);
and U715 (N_715,In_1929,In_807);
xnor U716 (N_716,In_709,In_612);
and U717 (N_717,In_194,In_1044);
or U718 (N_718,In_98,In_694);
nand U719 (N_719,In_115,In_1104);
or U720 (N_720,In_929,In_217);
nor U721 (N_721,In_631,In_1644);
nand U722 (N_722,In_1603,In_210);
nor U723 (N_723,In_1973,In_1324);
or U724 (N_724,In_27,In_1920);
or U725 (N_725,In_417,In_11);
nand U726 (N_726,In_615,In_1672);
or U727 (N_727,In_1533,In_1159);
nor U728 (N_728,In_797,In_1154);
and U729 (N_729,In_554,In_685);
nand U730 (N_730,In_867,In_197);
nor U731 (N_731,In_142,In_1155);
nand U732 (N_732,In_1218,In_1382);
and U733 (N_733,In_419,In_1330);
nor U734 (N_734,In_1841,In_1521);
nor U735 (N_735,In_204,In_1418);
and U736 (N_736,In_483,In_6);
or U737 (N_737,In_842,In_1772);
and U738 (N_738,In_424,In_219);
nor U739 (N_739,In_1910,In_380);
and U740 (N_740,In_1628,In_1941);
nand U741 (N_741,In_1006,In_1792);
or U742 (N_742,In_1311,In_935);
nor U743 (N_743,In_127,In_38);
nor U744 (N_744,In_1760,In_543);
nor U745 (N_745,In_56,In_838);
nand U746 (N_746,In_1883,In_1835);
nand U747 (N_747,In_77,In_512);
nand U748 (N_748,In_1197,In_165);
and U749 (N_749,In_1258,In_604);
or U750 (N_750,In_1131,In_909);
or U751 (N_751,In_1698,In_1298);
or U752 (N_752,In_727,In_358);
or U753 (N_753,In_1093,In_1852);
or U754 (N_754,In_328,In_1693);
or U755 (N_755,In_849,In_1078);
nand U756 (N_756,In_1294,In_563);
or U757 (N_757,In_244,In_1844);
nor U758 (N_758,In_303,In_1016);
nor U759 (N_759,In_408,In_301);
nand U760 (N_760,In_703,In_1847);
nand U761 (N_761,In_590,In_1520);
or U762 (N_762,In_1946,In_1307);
nand U763 (N_763,In_1729,In_802);
nor U764 (N_764,In_1546,In_72);
or U765 (N_765,In_1903,In_310);
and U766 (N_766,In_592,In_1208);
and U767 (N_767,In_1029,In_1252);
nand U768 (N_768,In_846,In_737);
or U769 (N_769,In_716,In_1026);
nand U770 (N_770,In_442,In_143);
and U771 (N_771,In_613,In_744);
and U772 (N_772,In_968,In_1170);
nor U773 (N_773,In_790,In_266);
nor U774 (N_774,In_1561,In_489);
and U775 (N_775,In_663,In_620);
or U776 (N_776,In_1291,In_580);
nand U777 (N_777,In_170,In_1579);
or U778 (N_778,In_1455,In_1730);
and U779 (N_779,In_1173,In_547);
nor U780 (N_780,In_40,In_1272);
and U781 (N_781,In_560,In_359);
and U782 (N_782,In_619,In_1443);
or U783 (N_783,In_1009,In_597);
nor U784 (N_784,In_1244,In_132);
and U785 (N_785,In_17,In_1187);
xor U786 (N_786,In_1161,In_1880);
and U787 (N_787,In_817,In_1925);
nor U788 (N_788,In_1988,In_1534);
and U789 (N_789,In_798,In_1432);
and U790 (N_790,In_1198,In_117);
and U791 (N_791,In_768,In_830);
nor U792 (N_792,In_1230,In_1914);
nand U793 (N_793,In_47,In_1153);
and U794 (N_794,In_928,In_514);
or U795 (N_795,In_57,In_1002);
or U796 (N_796,In_315,In_404);
and U797 (N_797,In_1345,In_769);
nor U798 (N_798,In_1242,In_956);
nor U799 (N_799,In_1319,In_1522);
nor U800 (N_800,In_1971,In_1851);
nand U801 (N_801,In_1181,In_396);
nor U802 (N_802,In_899,In_591);
and U803 (N_803,In_1702,In_1827);
and U804 (N_804,In_319,In_809);
and U805 (N_805,In_48,In_1337);
nand U806 (N_806,In_1552,In_1599);
and U807 (N_807,In_1235,In_859);
nand U808 (N_808,In_1616,In_1680);
and U809 (N_809,In_321,In_1968);
nor U810 (N_810,In_108,In_460);
nor U811 (N_811,In_1269,In_918);
nor U812 (N_812,In_1694,In_1121);
nor U813 (N_813,In_1986,In_1482);
or U814 (N_814,In_1927,In_939);
and U815 (N_815,In_722,In_995);
nand U816 (N_816,In_1106,In_1219);
nand U817 (N_817,In_1939,In_1926);
nand U818 (N_818,In_787,In_627);
xnor U819 (N_819,In_1531,In_1445);
or U820 (N_820,In_1209,In_728);
and U821 (N_821,In_1834,In_1991);
nor U822 (N_822,In_504,In_1512);
or U823 (N_823,In_201,In_916);
nand U824 (N_824,In_1855,In_233);
nand U825 (N_825,In_422,In_872);
and U826 (N_826,In_1313,In_1664);
or U827 (N_827,In_1565,In_440);
nand U828 (N_828,In_946,In_1799);
or U829 (N_829,In_1582,In_1065);
or U830 (N_830,In_944,In_1748);
nand U831 (N_831,In_692,In_680);
nand U832 (N_832,In_1499,In_70);
and U833 (N_833,In_1635,In_1204);
nand U834 (N_834,In_1604,In_1447);
nand U835 (N_835,In_701,In_331);
or U836 (N_836,In_854,In_144);
nand U837 (N_837,In_1385,In_582);
nand U838 (N_838,In_1409,In_609);
and U839 (N_839,In_915,In_544);
nor U840 (N_840,In_1000,In_589);
nand U841 (N_841,In_1348,In_1829);
nor U842 (N_842,In_957,In_1569);
or U843 (N_843,In_1607,In_1791);
nor U844 (N_844,In_178,In_806);
nor U845 (N_845,In_1381,In_161);
and U846 (N_846,In_1839,In_1716);
or U847 (N_847,In_850,In_1713);
nor U848 (N_848,In_1085,In_1958);
and U849 (N_849,In_207,In_665);
and U850 (N_850,In_1872,In_298);
or U851 (N_851,In_723,In_616);
and U852 (N_852,In_1636,In_1735);
nor U853 (N_853,In_925,In_1434);
nand U854 (N_854,In_1031,In_439);
nor U855 (N_855,In_348,In_500);
nor U856 (N_856,In_413,In_202);
xnor U857 (N_857,In_1959,In_102);
nor U858 (N_858,In_1092,In_940);
nor U859 (N_859,In_1098,In_126);
nand U860 (N_860,In_473,In_901);
or U861 (N_861,In_717,In_369);
xnor U862 (N_862,In_296,In_828);
or U863 (N_863,In_457,In_377);
or U864 (N_864,In_320,In_1020);
and U865 (N_865,In_825,In_989);
and U866 (N_866,In_710,In_241);
nand U867 (N_867,In_823,In_153);
and U868 (N_868,In_1895,In_750);
nand U869 (N_869,In_1177,In_1122);
nor U870 (N_870,In_12,In_1996);
nor U871 (N_871,In_1074,In_1979);
xnor U872 (N_872,In_76,In_1073);
or U873 (N_873,In_1898,In_1295);
and U874 (N_874,In_363,In_571);
nor U875 (N_875,In_1043,In_1224);
and U876 (N_876,In_452,In_156);
or U877 (N_877,In_1917,In_1323);
nand U878 (N_878,In_53,In_1596);
nor U879 (N_879,In_1221,In_190);
and U880 (N_880,In_847,In_39);
nand U881 (N_881,In_1933,In_1656);
or U882 (N_882,In_1062,In_376);
nand U883 (N_883,In_1174,In_1070);
and U884 (N_884,In_745,In_1615);
or U885 (N_885,In_279,In_1623);
and U886 (N_886,In_1537,In_26);
or U887 (N_887,In_1416,In_890);
nand U888 (N_888,In_883,In_1783);
or U889 (N_889,In_206,In_305);
nor U890 (N_890,In_1462,In_600);
and U891 (N_891,In_1388,In_297);
and U892 (N_892,In_1396,In_1549);
nor U893 (N_893,In_373,In_670);
or U894 (N_894,In_467,In_15);
nand U895 (N_895,In_1508,In_693);
nor U896 (N_896,In_1902,In_689);
nor U897 (N_897,In_423,In_855);
and U898 (N_898,In_351,In_496);
nor U899 (N_899,In_1806,In_1955);
nor U900 (N_900,In_1810,In_771);
nor U901 (N_901,In_1761,In_45);
nor U902 (N_902,In_1498,In_148);
nand U903 (N_903,In_1602,In_1641);
or U904 (N_904,In_325,In_1637);
and U905 (N_905,In_1797,In_428);
nand U906 (N_906,In_1595,In_1355);
nand U907 (N_907,In_20,In_1887);
or U908 (N_908,In_1870,In_1830);
and U909 (N_909,In_93,In_474);
and U910 (N_910,In_1828,In_1086);
nand U911 (N_911,In_130,In_707);
nand U912 (N_912,In_51,In_1331);
nand U913 (N_913,In_573,In_598);
nor U914 (N_914,In_1234,In_1076);
nand U915 (N_915,In_1633,In_1982);
nor U916 (N_916,In_1576,In_900);
and U917 (N_917,In_629,In_515);
and U918 (N_918,In_1600,In_163);
or U919 (N_919,In_59,In_799);
or U920 (N_920,In_948,In_1146);
nand U921 (N_921,In_135,In_1408);
or U922 (N_922,In_584,In_1833);
or U923 (N_923,In_996,In_993);
nor U924 (N_924,In_540,In_1217);
and U925 (N_925,In_267,In_166);
and U926 (N_926,In_312,In_420);
or U927 (N_927,In_1790,In_1328);
or U928 (N_928,In_1739,In_1861);
and U929 (N_929,In_760,In_329);
nor U930 (N_930,In_1645,In_187);
nand U931 (N_931,In_265,In_1715);
nand U932 (N_932,In_393,In_78);
or U933 (N_933,In_894,In_531);
nand U934 (N_934,In_58,In_234);
nor U935 (N_935,In_22,In_1363);
nand U936 (N_936,In_24,In_1583);
nor U937 (N_937,In_1589,In_715);
nor U938 (N_938,In_1277,In_1333);
or U939 (N_939,In_299,In_622);
and U940 (N_940,In_1485,In_237);
and U941 (N_941,In_1750,In_1874);
and U942 (N_942,In_1088,In_907);
and U943 (N_943,In_1371,In_19);
nand U944 (N_944,In_387,In_1975);
nand U945 (N_945,In_368,In_784);
nor U946 (N_946,In_224,In_411);
nand U947 (N_947,In_1824,In_235);
nand U948 (N_948,In_448,In_632);
and U949 (N_949,In_1663,In_28);
or U950 (N_950,In_389,In_550);
or U951 (N_951,In_1678,In_324);
nor U952 (N_952,In_1210,In_1178);
and U953 (N_953,In_205,In_239);
nand U954 (N_954,In_962,In_1377);
nor U955 (N_955,In_96,In_862);
nand U956 (N_956,In_334,In_1980);
or U957 (N_957,In_1481,In_1759);
or U958 (N_958,In_1751,In_1501);
nand U959 (N_959,In_1639,In_1393);
or U960 (N_960,In_168,In_134);
and U961 (N_961,In_960,In_1372);
and U962 (N_962,In_923,In_579);
or U963 (N_963,In_304,In_845);
or U964 (N_964,In_1200,In_975);
and U965 (N_965,In_949,In_1452);
or U966 (N_966,In_91,In_1052);
and U967 (N_967,In_1858,In_1614);
or U968 (N_968,In_464,In_1548);
nand U969 (N_969,In_459,In_1666);
or U970 (N_970,In_645,In_1454);
nand U971 (N_971,In_1794,In_406);
or U972 (N_972,In_587,In_1651);
or U973 (N_973,In_599,In_1435);
or U974 (N_974,In_1023,In_941);
or U975 (N_975,In_447,In_1075);
nor U976 (N_976,In_5,In_625);
and U977 (N_977,In_109,In_1147);
nand U978 (N_978,In_1413,In_451);
and U979 (N_979,In_1524,In_381);
and U980 (N_980,In_1665,In_1879);
nor U981 (N_981,In_1670,In_1438);
or U982 (N_982,In_1041,In_1785);
and U983 (N_983,In_994,In_196);
or U984 (N_984,In_1100,In_1296);
or U985 (N_985,In_1458,In_648);
nor U986 (N_986,In_1753,In_1233);
and U987 (N_987,In_105,In_656);
nand U988 (N_988,In_1460,In_1424);
nor U989 (N_989,In_1304,In_256);
nand U990 (N_990,In_691,In_333);
or U991 (N_991,In_169,In_1457);
nor U992 (N_992,In_1202,In_511);
nor U993 (N_993,In_1647,In_766);
xnor U994 (N_994,In_869,In_1814);
or U995 (N_995,In_1400,In_999);
and U996 (N_996,In_681,In_1229);
and U997 (N_997,In_1247,In_1717);
nand U998 (N_998,In_934,In_1038);
nand U999 (N_999,In_1410,In_713);
and U1000 (N_1000,In_196,In_1107);
nor U1001 (N_1001,In_787,In_213);
and U1002 (N_1002,In_598,In_1620);
nor U1003 (N_1003,In_706,In_1971);
and U1004 (N_1004,In_64,In_1705);
or U1005 (N_1005,In_725,In_1874);
and U1006 (N_1006,In_613,In_1289);
nand U1007 (N_1007,In_1943,In_926);
and U1008 (N_1008,In_967,In_1314);
and U1009 (N_1009,In_152,In_1073);
nand U1010 (N_1010,In_1407,In_1663);
or U1011 (N_1011,In_1926,In_1704);
nor U1012 (N_1012,In_1381,In_292);
or U1013 (N_1013,In_923,In_1793);
or U1014 (N_1014,In_1026,In_215);
nor U1015 (N_1015,In_629,In_676);
and U1016 (N_1016,In_923,In_51);
nor U1017 (N_1017,In_1033,In_875);
and U1018 (N_1018,In_271,In_380);
nor U1019 (N_1019,In_1169,In_1111);
and U1020 (N_1020,In_196,In_1984);
and U1021 (N_1021,In_568,In_35);
nor U1022 (N_1022,In_959,In_617);
nand U1023 (N_1023,In_1644,In_1629);
or U1024 (N_1024,In_1959,In_1001);
or U1025 (N_1025,In_1282,In_829);
nand U1026 (N_1026,In_718,In_1194);
nand U1027 (N_1027,In_1321,In_1935);
nor U1028 (N_1028,In_1347,In_1441);
and U1029 (N_1029,In_1026,In_984);
nand U1030 (N_1030,In_855,In_1487);
nor U1031 (N_1031,In_1857,In_1498);
nand U1032 (N_1032,In_1160,In_573);
nand U1033 (N_1033,In_652,In_405);
and U1034 (N_1034,In_854,In_1507);
or U1035 (N_1035,In_1300,In_1965);
or U1036 (N_1036,In_1123,In_448);
and U1037 (N_1037,In_378,In_1514);
and U1038 (N_1038,In_1000,In_205);
nand U1039 (N_1039,In_1690,In_557);
nor U1040 (N_1040,In_728,In_1232);
nand U1041 (N_1041,In_1704,In_1667);
and U1042 (N_1042,In_823,In_849);
nor U1043 (N_1043,In_798,In_78);
and U1044 (N_1044,In_1290,In_264);
nor U1045 (N_1045,In_1884,In_52);
xor U1046 (N_1046,In_700,In_179);
nand U1047 (N_1047,In_98,In_243);
nor U1048 (N_1048,In_1272,In_135);
nor U1049 (N_1049,In_1758,In_865);
nand U1050 (N_1050,In_1009,In_1190);
or U1051 (N_1051,In_1995,In_94);
nor U1052 (N_1052,In_1848,In_898);
and U1053 (N_1053,In_69,In_1608);
nand U1054 (N_1054,In_114,In_412);
and U1055 (N_1055,In_312,In_1285);
nor U1056 (N_1056,In_188,In_1400);
or U1057 (N_1057,In_1775,In_610);
nor U1058 (N_1058,In_1399,In_353);
or U1059 (N_1059,In_1516,In_777);
nor U1060 (N_1060,In_1894,In_969);
nor U1061 (N_1061,In_858,In_103);
nand U1062 (N_1062,In_457,In_1877);
nand U1063 (N_1063,In_1744,In_603);
nand U1064 (N_1064,In_1532,In_390);
nand U1065 (N_1065,In_807,In_750);
or U1066 (N_1066,In_1364,In_1166);
and U1067 (N_1067,In_269,In_254);
or U1068 (N_1068,In_1750,In_1345);
nor U1069 (N_1069,In_376,In_73);
nor U1070 (N_1070,In_3,In_1411);
or U1071 (N_1071,In_268,In_1110);
nand U1072 (N_1072,In_321,In_1079);
or U1073 (N_1073,In_867,In_1338);
and U1074 (N_1074,In_846,In_1775);
nand U1075 (N_1075,In_465,In_549);
and U1076 (N_1076,In_675,In_755);
nand U1077 (N_1077,In_536,In_1447);
nor U1078 (N_1078,In_1982,In_1540);
and U1079 (N_1079,In_1816,In_572);
and U1080 (N_1080,In_342,In_1244);
and U1081 (N_1081,In_677,In_1413);
and U1082 (N_1082,In_54,In_1205);
and U1083 (N_1083,In_1250,In_783);
nand U1084 (N_1084,In_948,In_1088);
and U1085 (N_1085,In_141,In_1700);
or U1086 (N_1086,In_860,In_948);
or U1087 (N_1087,In_434,In_200);
nand U1088 (N_1088,In_1064,In_1831);
or U1089 (N_1089,In_1747,In_243);
nand U1090 (N_1090,In_1388,In_233);
nor U1091 (N_1091,In_241,In_1561);
or U1092 (N_1092,In_329,In_1850);
and U1093 (N_1093,In_1887,In_1442);
and U1094 (N_1094,In_801,In_17);
nand U1095 (N_1095,In_1208,In_1120);
or U1096 (N_1096,In_387,In_406);
and U1097 (N_1097,In_1059,In_1483);
and U1098 (N_1098,In_1850,In_1530);
nand U1099 (N_1099,In_20,In_1370);
nand U1100 (N_1100,In_1193,In_1662);
or U1101 (N_1101,In_260,In_737);
and U1102 (N_1102,In_842,In_832);
and U1103 (N_1103,In_1258,In_269);
nor U1104 (N_1104,In_903,In_509);
nand U1105 (N_1105,In_795,In_1208);
or U1106 (N_1106,In_1641,In_1955);
nor U1107 (N_1107,In_1937,In_1945);
or U1108 (N_1108,In_159,In_1923);
nand U1109 (N_1109,In_1077,In_1896);
nand U1110 (N_1110,In_675,In_867);
and U1111 (N_1111,In_800,In_1412);
or U1112 (N_1112,In_616,In_1544);
and U1113 (N_1113,In_353,In_1451);
and U1114 (N_1114,In_1344,In_1300);
nand U1115 (N_1115,In_1098,In_480);
nand U1116 (N_1116,In_723,In_1461);
and U1117 (N_1117,In_1037,In_458);
or U1118 (N_1118,In_355,In_807);
and U1119 (N_1119,In_986,In_1401);
xnor U1120 (N_1120,In_1132,In_1375);
nor U1121 (N_1121,In_1387,In_999);
nor U1122 (N_1122,In_412,In_865);
nand U1123 (N_1123,In_1426,In_1787);
or U1124 (N_1124,In_1246,In_333);
or U1125 (N_1125,In_1919,In_941);
nor U1126 (N_1126,In_329,In_1443);
or U1127 (N_1127,In_448,In_1998);
nor U1128 (N_1128,In_1410,In_324);
nand U1129 (N_1129,In_1364,In_1506);
or U1130 (N_1130,In_1764,In_963);
nand U1131 (N_1131,In_1697,In_295);
nand U1132 (N_1132,In_677,In_1103);
or U1133 (N_1133,In_1949,In_165);
nor U1134 (N_1134,In_493,In_601);
and U1135 (N_1135,In_1706,In_478);
nand U1136 (N_1136,In_186,In_1359);
and U1137 (N_1137,In_473,In_1315);
or U1138 (N_1138,In_1239,In_99);
or U1139 (N_1139,In_790,In_1889);
nor U1140 (N_1140,In_1073,In_63);
nor U1141 (N_1141,In_1314,In_470);
nor U1142 (N_1142,In_634,In_1131);
nand U1143 (N_1143,In_1016,In_1432);
nor U1144 (N_1144,In_1597,In_1277);
nor U1145 (N_1145,In_305,In_527);
or U1146 (N_1146,In_231,In_1426);
nor U1147 (N_1147,In_1457,In_1228);
or U1148 (N_1148,In_320,In_1725);
nand U1149 (N_1149,In_1360,In_613);
nor U1150 (N_1150,In_1696,In_810);
or U1151 (N_1151,In_251,In_1008);
nor U1152 (N_1152,In_840,In_842);
or U1153 (N_1153,In_1297,In_197);
nor U1154 (N_1154,In_476,In_1018);
nor U1155 (N_1155,In_42,In_998);
nand U1156 (N_1156,In_1678,In_176);
nor U1157 (N_1157,In_1256,In_730);
xnor U1158 (N_1158,In_691,In_1964);
and U1159 (N_1159,In_233,In_1534);
and U1160 (N_1160,In_1312,In_1753);
nand U1161 (N_1161,In_107,In_774);
nand U1162 (N_1162,In_638,In_1415);
nand U1163 (N_1163,In_755,In_730);
or U1164 (N_1164,In_1974,In_639);
or U1165 (N_1165,In_1230,In_386);
and U1166 (N_1166,In_469,In_1302);
nand U1167 (N_1167,In_742,In_1302);
nor U1168 (N_1168,In_1708,In_1679);
or U1169 (N_1169,In_941,In_558);
nand U1170 (N_1170,In_1776,In_165);
or U1171 (N_1171,In_314,In_1135);
and U1172 (N_1172,In_1894,In_1652);
nor U1173 (N_1173,In_1674,In_401);
nor U1174 (N_1174,In_127,In_236);
or U1175 (N_1175,In_1498,In_84);
nand U1176 (N_1176,In_919,In_1322);
nor U1177 (N_1177,In_1693,In_1111);
nand U1178 (N_1178,In_1570,In_715);
nor U1179 (N_1179,In_1904,In_896);
and U1180 (N_1180,In_1915,In_220);
and U1181 (N_1181,In_1669,In_1181);
or U1182 (N_1182,In_1784,In_1133);
and U1183 (N_1183,In_1138,In_1854);
and U1184 (N_1184,In_199,In_1548);
and U1185 (N_1185,In_1180,In_989);
nor U1186 (N_1186,In_602,In_1304);
or U1187 (N_1187,In_1725,In_417);
nor U1188 (N_1188,In_1323,In_1037);
and U1189 (N_1189,In_516,In_581);
and U1190 (N_1190,In_683,In_1657);
nor U1191 (N_1191,In_990,In_323);
nor U1192 (N_1192,In_1240,In_201);
or U1193 (N_1193,In_52,In_1367);
nor U1194 (N_1194,In_1642,In_1182);
or U1195 (N_1195,In_1022,In_571);
and U1196 (N_1196,In_1442,In_1560);
or U1197 (N_1197,In_1464,In_1740);
or U1198 (N_1198,In_1936,In_792);
or U1199 (N_1199,In_854,In_1982);
nor U1200 (N_1200,In_1606,In_994);
or U1201 (N_1201,In_311,In_640);
nor U1202 (N_1202,In_1720,In_1197);
or U1203 (N_1203,In_831,In_1323);
and U1204 (N_1204,In_760,In_579);
nand U1205 (N_1205,In_1346,In_183);
or U1206 (N_1206,In_610,In_1377);
nor U1207 (N_1207,In_76,In_25);
and U1208 (N_1208,In_389,In_710);
and U1209 (N_1209,In_180,In_90);
nand U1210 (N_1210,In_434,In_39);
or U1211 (N_1211,In_1965,In_810);
and U1212 (N_1212,In_487,In_1008);
and U1213 (N_1213,In_1707,In_1812);
or U1214 (N_1214,In_1591,In_1068);
nand U1215 (N_1215,In_299,In_1257);
nand U1216 (N_1216,In_1475,In_125);
nand U1217 (N_1217,In_518,In_1326);
nor U1218 (N_1218,In_716,In_393);
nand U1219 (N_1219,In_567,In_529);
nand U1220 (N_1220,In_651,In_491);
and U1221 (N_1221,In_1420,In_1223);
nand U1222 (N_1222,In_1937,In_1981);
and U1223 (N_1223,In_1403,In_1963);
and U1224 (N_1224,In_989,In_436);
and U1225 (N_1225,In_878,In_112);
nand U1226 (N_1226,In_1997,In_731);
and U1227 (N_1227,In_863,In_1649);
nor U1228 (N_1228,In_357,In_232);
or U1229 (N_1229,In_766,In_541);
and U1230 (N_1230,In_542,In_1598);
or U1231 (N_1231,In_1120,In_448);
or U1232 (N_1232,In_970,In_623);
or U1233 (N_1233,In_1151,In_1970);
nor U1234 (N_1234,In_1697,In_1934);
nor U1235 (N_1235,In_967,In_1981);
and U1236 (N_1236,In_366,In_370);
or U1237 (N_1237,In_1180,In_1830);
nor U1238 (N_1238,In_757,In_605);
nor U1239 (N_1239,In_534,In_1113);
nor U1240 (N_1240,In_1839,In_1276);
and U1241 (N_1241,In_457,In_1232);
or U1242 (N_1242,In_1594,In_435);
nand U1243 (N_1243,In_850,In_1488);
and U1244 (N_1244,In_1396,In_838);
and U1245 (N_1245,In_831,In_1090);
or U1246 (N_1246,In_812,In_213);
nor U1247 (N_1247,In_464,In_351);
or U1248 (N_1248,In_1288,In_510);
or U1249 (N_1249,In_1537,In_1062);
nand U1250 (N_1250,In_1986,In_1207);
and U1251 (N_1251,In_577,In_1096);
nor U1252 (N_1252,In_1207,In_1578);
nand U1253 (N_1253,In_1652,In_1386);
and U1254 (N_1254,In_587,In_347);
and U1255 (N_1255,In_1038,In_1677);
or U1256 (N_1256,In_885,In_28);
and U1257 (N_1257,In_284,In_1743);
or U1258 (N_1258,In_1583,In_216);
and U1259 (N_1259,In_756,In_931);
or U1260 (N_1260,In_1810,In_1046);
or U1261 (N_1261,In_1932,In_358);
and U1262 (N_1262,In_1131,In_1520);
and U1263 (N_1263,In_574,In_1802);
nor U1264 (N_1264,In_430,In_1389);
and U1265 (N_1265,In_1465,In_1544);
xnor U1266 (N_1266,In_1536,In_1693);
or U1267 (N_1267,In_578,In_166);
nor U1268 (N_1268,In_266,In_1617);
and U1269 (N_1269,In_914,In_945);
nand U1270 (N_1270,In_1520,In_814);
nand U1271 (N_1271,In_1493,In_804);
or U1272 (N_1272,In_143,In_487);
and U1273 (N_1273,In_739,In_669);
nand U1274 (N_1274,In_1562,In_1691);
nand U1275 (N_1275,In_385,In_618);
nand U1276 (N_1276,In_182,In_928);
nor U1277 (N_1277,In_484,In_804);
nor U1278 (N_1278,In_594,In_94);
nor U1279 (N_1279,In_829,In_192);
nor U1280 (N_1280,In_1858,In_1258);
nand U1281 (N_1281,In_531,In_518);
or U1282 (N_1282,In_1425,In_1858);
and U1283 (N_1283,In_1572,In_897);
or U1284 (N_1284,In_1954,In_180);
nand U1285 (N_1285,In_1961,In_1356);
and U1286 (N_1286,In_692,In_1055);
or U1287 (N_1287,In_958,In_1478);
nand U1288 (N_1288,In_1079,In_1366);
and U1289 (N_1289,In_1630,In_807);
or U1290 (N_1290,In_467,In_1745);
or U1291 (N_1291,In_420,In_1973);
nand U1292 (N_1292,In_173,In_1330);
or U1293 (N_1293,In_228,In_651);
nand U1294 (N_1294,In_1957,In_1824);
nand U1295 (N_1295,In_209,In_1286);
nand U1296 (N_1296,In_1612,In_623);
and U1297 (N_1297,In_652,In_1202);
nand U1298 (N_1298,In_840,In_1081);
nand U1299 (N_1299,In_1753,In_209);
nand U1300 (N_1300,In_897,In_892);
nand U1301 (N_1301,In_1631,In_51);
nand U1302 (N_1302,In_589,In_1815);
and U1303 (N_1303,In_34,In_644);
nand U1304 (N_1304,In_1746,In_1180);
and U1305 (N_1305,In_1599,In_1076);
and U1306 (N_1306,In_1109,In_1339);
or U1307 (N_1307,In_1528,In_1469);
nand U1308 (N_1308,In_560,In_1840);
or U1309 (N_1309,In_469,In_1473);
nand U1310 (N_1310,In_842,In_1527);
nor U1311 (N_1311,In_1176,In_1190);
nand U1312 (N_1312,In_1264,In_580);
nand U1313 (N_1313,In_444,In_278);
xor U1314 (N_1314,In_163,In_387);
or U1315 (N_1315,In_1026,In_571);
nand U1316 (N_1316,In_754,In_1734);
and U1317 (N_1317,In_1553,In_576);
nor U1318 (N_1318,In_1940,In_676);
and U1319 (N_1319,In_19,In_117);
or U1320 (N_1320,In_1086,In_1420);
nand U1321 (N_1321,In_485,In_1400);
nand U1322 (N_1322,In_832,In_748);
nand U1323 (N_1323,In_1765,In_1500);
nand U1324 (N_1324,In_1801,In_1363);
nand U1325 (N_1325,In_760,In_948);
and U1326 (N_1326,In_1295,In_1716);
nor U1327 (N_1327,In_181,In_507);
nor U1328 (N_1328,In_1947,In_97);
nand U1329 (N_1329,In_25,In_294);
or U1330 (N_1330,In_85,In_1822);
nand U1331 (N_1331,In_1065,In_1589);
nand U1332 (N_1332,In_423,In_436);
nand U1333 (N_1333,In_388,In_295);
and U1334 (N_1334,In_19,In_1394);
nand U1335 (N_1335,In_1469,In_158);
and U1336 (N_1336,In_105,In_1496);
nor U1337 (N_1337,In_1328,In_90);
and U1338 (N_1338,In_1400,In_216);
nor U1339 (N_1339,In_1637,In_1124);
and U1340 (N_1340,In_964,In_1593);
and U1341 (N_1341,In_1681,In_349);
nand U1342 (N_1342,In_1527,In_1109);
nor U1343 (N_1343,In_345,In_1965);
nor U1344 (N_1344,In_1765,In_1137);
nor U1345 (N_1345,In_851,In_1552);
and U1346 (N_1346,In_157,In_1931);
nand U1347 (N_1347,In_1323,In_1427);
and U1348 (N_1348,In_487,In_1916);
nand U1349 (N_1349,In_271,In_284);
nor U1350 (N_1350,In_593,In_1546);
and U1351 (N_1351,In_1338,In_47);
nor U1352 (N_1352,In_1860,In_1733);
or U1353 (N_1353,In_1153,In_983);
nand U1354 (N_1354,In_922,In_441);
and U1355 (N_1355,In_565,In_1082);
and U1356 (N_1356,In_1541,In_1231);
and U1357 (N_1357,In_87,In_585);
and U1358 (N_1358,In_1544,In_803);
or U1359 (N_1359,In_436,In_1790);
and U1360 (N_1360,In_575,In_646);
nand U1361 (N_1361,In_1748,In_479);
nor U1362 (N_1362,In_1531,In_631);
nor U1363 (N_1363,In_1512,In_720);
or U1364 (N_1364,In_34,In_1624);
nand U1365 (N_1365,In_384,In_1225);
and U1366 (N_1366,In_319,In_1792);
nand U1367 (N_1367,In_1975,In_568);
or U1368 (N_1368,In_423,In_144);
nor U1369 (N_1369,In_942,In_1098);
nand U1370 (N_1370,In_3,In_1730);
or U1371 (N_1371,In_713,In_820);
nor U1372 (N_1372,In_147,In_507);
or U1373 (N_1373,In_514,In_1593);
and U1374 (N_1374,In_50,In_815);
nor U1375 (N_1375,In_1202,In_52);
nor U1376 (N_1376,In_1232,In_1603);
and U1377 (N_1377,In_798,In_951);
and U1378 (N_1378,In_342,In_1885);
or U1379 (N_1379,In_1377,In_387);
or U1380 (N_1380,In_1397,In_1840);
nand U1381 (N_1381,In_1022,In_1164);
and U1382 (N_1382,In_394,In_1304);
or U1383 (N_1383,In_388,In_48);
nor U1384 (N_1384,In_161,In_213);
xor U1385 (N_1385,In_689,In_1229);
nand U1386 (N_1386,In_1709,In_884);
nand U1387 (N_1387,In_550,In_129);
nand U1388 (N_1388,In_1553,In_1504);
or U1389 (N_1389,In_325,In_882);
nand U1390 (N_1390,In_1778,In_1354);
nor U1391 (N_1391,In_1570,In_397);
nor U1392 (N_1392,In_627,In_60);
nor U1393 (N_1393,In_219,In_1960);
nor U1394 (N_1394,In_1622,In_432);
nor U1395 (N_1395,In_109,In_1823);
or U1396 (N_1396,In_1159,In_472);
nand U1397 (N_1397,In_401,In_1825);
nor U1398 (N_1398,In_1578,In_427);
or U1399 (N_1399,In_1840,In_974);
or U1400 (N_1400,In_1366,In_1013);
and U1401 (N_1401,In_646,In_1073);
nor U1402 (N_1402,In_411,In_1843);
nor U1403 (N_1403,In_98,In_1745);
xnor U1404 (N_1404,In_1501,In_1375);
nor U1405 (N_1405,In_1884,In_129);
xor U1406 (N_1406,In_72,In_1063);
nand U1407 (N_1407,In_1189,In_23);
and U1408 (N_1408,In_248,In_553);
and U1409 (N_1409,In_821,In_937);
nand U1410 (N_1410,In_492,In_895);
or U1411 (N_1411,In_332,In_727);
or U1412 (N_1412,In_1387,In_4);
and U1413 (N_1413,In_1508,In_683);
nand U1414 (N_1414,In_1547,In_340);
or U1415 (N_1415,In_615,In_38);
nor U1416 (N_1416,In_663,In_1094);
or U1417 (N_1417,In_1263,In_23);
nor U1418 (N_1418,In_958,In_550);
or U1419 (N_1419,In_302,In_1074);
and U1420 (N_1420,In_720,In_1374);
nor U1421 (N_1421,In_944,In_1076);
nor U1422 (N_1422,In_563,In_1728);
and U1423 (N_1423,In_1132,In_1801);
nor U1424 (N_1424,In_1380,In_1179);
nand U1425 (N_1425,In_1299,In_761);
nor U1426 (N_1426,In_1313,In_787);
nor U1427 (N_1427,In_613,In_1376);
nand U1428 (N_1428,In_1842,In_1445);
or U1429 (N_1429,In_524,In_1454);
nand U1430 (N_1430,In_1685,In_1523);
nor U1431 (N_1431,In_761,In_846);
or U1432 (N_1432,In_1422,In_1666);
nor U1433 (N_1433,In_545,In_28);
nor U1434 (N_1434,In_878,In_1415);
nand U1435 (N_1435,In_439,In_60);
or U1436 (N_1436,In_1141,In_929);
nor U1437 (N_1437,In_1779,In_1701);
nand U1438 (N_1438,In_1218,In_642);
nor U1439 (N_1439,In_487,In_672);
and U1440 (N_1440,In_1640,In_606);
nor U1441 (N_1441,In_683,In_1995);
nand U1442 (N_1442,In_1501,In_363);
nor U1443 (N_1443,In_953,In_1259);
and U1444 (N_1444,In_1490,In_296);
or U1445 (N_1445,In_269,In_686);
nand U1446 (N_1446,In_782,In_733);
nor U1447 (N_1447,In_945,In_751);
and U1448 (N_1448,In_1670,In_131);
nand U1449 (N_1449,In_840,In_1690);
and U1450 (N_1450,In_522,In_528);
or U1451 (N_1451,In_634,In_731);
or U1452 (N_1452,In_897,In_97);
nor U1453 (N_1453,In_854,In_1734);
nand U1454 (N_1454,In_1378,In_1115);
or U1455 (N_1455,In_750,In_1252);
nand U1456 (N_1456,In_1676,In_449);
or U1457 (N_1457,In_1313,In_155);
and U1458 (N_1458,In_179,In_1479);
nand U1459 (N_1459,In_969,In_928);
or U1460 (N_1460,In_224,In_1815);
and U1461 (N_1461,In_1226,In_131);
and U1462 (N_1462,In_1338,In_1401);
or U1463 (N_1463,In_464,In_1317);
nor U1464 (N_1464,In_1424,In_1726);
nor U1465 (N_1465,In_27,In_724);
and U1466 (N_1466,In_206,In_804);
nor U1467 (N_1467,In_839,In_1247);
and U1468 (N_1468,In_396,In_1123);
or U1469 (N_1469,In_493,In_1252);
and U1470 (N_1470,In_1632,In_822);
or U1471 (N_1471,In_211,In_48);
nand U1472 (N_1472,In_665,In_416);
nand U1473 (N_1473,In_1639,In_1390);
and U1474 (N_1474,In_820,In_212);
and U1475 (N_1475,In_1193,In_1135);
or U1476 (N_1476,In_539,In_1420);
and U1477 (N_1477,In_177,In_308);
and U1478 (N_1478,In_1673,In_1628);
and U1479 (N_1479,In_1245,In_1316);
nand U1480 (N_1480,In_298,In_856);
nand U1481 (N_1481,In_672,In_740);
or U1482 (N_1482,In_772,In_767);
and U1483 (N_1483,In_1734,In_1505);
nand U1484 (N_1484,In_396,In_61);
nor U1485 (N_1485,In_1150,In_898);
and U1486 (N_1486,In_1775,In_1919);
or U1487 (N_1487,In_368,In_1972);
or U1488 (N_1488,In_268,In_890);
or U1489 (N_1489,In_931,In_903);
nand U1490 (N_1490,In_1852,In_312);
and U1491 (N_1491,In_212,In_1689);
and U1492 (N_1492,In_72,In_807);
nand U1493 (N_1493,In_156,In_434);
nand U1494 (N_1494,In_952,In_1612);
nand U1495 (N_1495,In_1709,In_1867);
or U1496 (N_1496,In_1286,In_1459);
or U1497 (N_1497,In_1387,In_84);
or U1498 (N_1498,In_1236,In_357);
nor U1499 (N_1499,In_934,In_544);
or U1500 (N_1500,In_98,In_1004);
xor U1501 (N_1501,In_67,In_1563);
nand U1502 (N_1502,In_446,In_246);
or U1503 (N_1503,In_1493,In_1124);
and U1504 (N_1504,In_192,In_854);
or U1505 (N_1505,In_1520,In_457);
nor U1506 (N_1506,In_1419,In_802);
nand U1507 (N_1507,In_1917,In_34);
or U1508 (N_1508,In_1662,In_87);
nand U1509 (N_1509,In_515,In_273);
nand U1510 (N_1510,In_1467,In_379);
nor U1511 (N_1511,In_1391,In_1030);
and U1512 (N_1512,In_1089,In_204);
and U1513 (N_1513,In_1654,In_1674);
nand U1514 (N_1514,In_679,In_1969);
or U1515 (N_1515,In_1663,In_772);
or U1516 (N_1516,In_1868,In_1620);
and U1517 (N_1517,In_482,In_1431);
and U1518 (N_1518,In_1520,In_1840);
and U1519 (N_1519,In_465,In_1152);
or U1520 (N_1520,In_491,In_1792);
nor U1521 (N_1521,In_561,In_167);
nand U1522 (N_1522,In_1388,In_1357);
nor U1523 (N_1523,In_1197,In_276);
or U1524 (N_1524,In_875,In_1514);
or U1525 (N_1525,In_1345,In_1087);
nor U1526 (N_1526,In_1514,In_890);
or U1527 (N_1527,In_114,In_118);
nor U1528 (N_1528,In_593,In_1897);
and U1529 (N_1529,In_290,In_1280);
and U1530 (N_1530,In_1383,In_1746);
nor U1531 (N_1531,In_339,In_952);
nand U1532 (N_1532,In_754,In_289);
nand U1533 (N_1533,In_1640,In_568);
xnor U1534 (N_1534,In_1224,In_623);
or U1535 (N_1535,In_1612,In_1632);
and U1536 (N_1536,In_927,In_1838);
nand U1537 (N_1537,In_546,In_728);
xor U1538 (N_1538,In_1252,In_652);
and U1539 (N_1539,In_182,In_1272);
and U1540 (N_1540,In_1817,In_1149);
nor U1541 (N_1541,In_459,In_1509);
or U1542 (N_1542,In_1446,In_1957);
xor U1543 (N_1543,In_65,In_1305);
and U1544 (N_1544,In_1607,In_1771);
or U1545 (N_1545,In_969,In_1107);
or U1546 (N_1546,In_1506,In_1408);
and U1547 (N_1547,In_886,In_609);
nand U1548 (N_1548,In_1137,In_1754);
or U1549 (N_1549,In_1073,In_1117);
nand U1550 (N_1550,In_1414,In_480);
or U1551 (N_1551,In_1239,In_321);
nor U1552 (N_1552,In_119,In_1586);
nand U1553 (N_1553,In_978,In_1904);
nor U1554 (N_1554,In_774,In_1622);
nor U1555 (N_1555,In_250,In_1163);
and U1556 (N_1556,In_1323,In_690);
or U1557 (N_1557,In_1045,In_1224);
or U1558 (N_1558,In_1041,In_856);
or U1559 (N_1559,In_1336,In_1322);
nand U1560 (N_1560,In_304,In_112);
nand U1561 (N_1561,In_672,In_1366);
or U1562 (N_1562,In_1054,In_887);
and U1563 (N_1563,In_522,In_1254);
or U1564 (N_1564,In_1806,In_1947);
nand U1565 (N_1565,In_712,In_145);
or U1566 (N_1566,In_253,In_559);
nor U1567 (N_1567,In_1942,In_328);
nand U1568 (N_1568,In_779,In_1707);
nor U1569 (N_1569,In_1812,In_1534);
and U1570 (N_1570,In_701,In_927);
or U1571 (N_1571,In_1644,In_442);
nor U1572 (N_1572,In_505,In_1614);
and U1573 (N_1573,In_1376,In_1592);
and U1574 (N_1574,In_1130,In_1528);
nor U1575 (N_1575,In_382,In_1315);
and U1576 (N_1576,In_1768,In_1060);
and U1577 (N_1577,In_1210,In_763);
nand U1578 (N_1578,In_583,In_1681);
nor U1579 (N_1579,In_1658,In_650);
and U1580 (N_1580,In_514,In_156);
and U1581 (N_1581,In_1951,In_897);
or U1582 (N_1582,In_1121,In_223);
or U1583 (N_1583,In_1948,In_263);
and U1584 (N_1584,In_882,In_1919);
or U1585 (N_1585,In_405,In_193);
nand U1586 (N_1586,In_67,In_1839);
and U1587 (N_1587,In_907,In_661);
nand U1588 (N_1588,In_1323,In_1897);
and U1589 (N_1589,In_1521,In_1853);
nor U1590 (N_1590,In_1129,In_193);
and U1591 (N_1591,In_194,In_803);
or U1592 (N_1592,In_551,In_944);
and U1593 (N_1593,In_869,In_207);
nand U1594 (N_1594,In_99,In_537);
and U1595 (N_1595,In_1177,In_1345);
or U1596 (N_1596,In_484,In_71);
nor U1597 (N_1597,In_1992,In_110);
and U1598 (N_1598,In_1307,In_653);
or U1599 (N_1599,In_1336,In_1450);
and U1600 (N_1600,In_21,In_470);
nand U1601 (N_1601,In_1071,In_335);
nand U1602 (N_1602,In_2,In_423);
and U1603 (N_1603,In_1022,In_1914);
and U1604 (N_1604,In_745,In_430);
or U1605 (N_1605,In_831,In_1917);
nand U1606 (N_1606,In_1326,In_1151);
nor U1607 (N_1607,In_930,In_69);
and U1608 (N_1608,In_404,In_1834);
or U1609 (N_1609,In_1552,In_1153);
nand U1610 (N_1610,In_757,In_1140);
or U1611 (N_1611,In_1350,In_1256);
and U1612 (N_1612,In_501,In_1510);
nor U1613 (N_1613,In_534,In_239);
and U1614 (N_1614,In_59,In_1625);
nand U1615 (N_1615,In_1122,In_1830);
or U1616 (N_1616,In_194,In_1982);
or U1617 (N_1617,In_1007,In_1783);
nor U1618 (N_1618,In_1023,In_596);
or U1619 (N_1619,In_1511,In_1295);
or U1620 (N_1620,In_1612,In_874);
nand U1621 (N_1621,In_849,In_1268);
nor U1622 (N_1622,In_654,In_1666);
or U1623 (N_1623,In_1707,In_1524);
or U1624 (N_1624,In_515,In_628);
or U1625 (N_1625,In_1841,In_1454);
and U1626 (N_1626,In_384,In_910);
nand U1627 (N_1627,In_1728,In_452);
nor U1628 (N_1628,In_1211,In_1421);
nor U1629 (N_1629,In_162,In_541);
and U1630 (N_1630,In_230,In_1431);
or U1631 (N_1631,In_1758,In_993);
or U1632 (N_1632,In_379,In_31);
nor U1633 (N_1633,In_1335,In_1885);
and U1634 (N_1634,In_841,In_242);
nor U1635 (N_1635,In_1490,In_749);
and U1636 (N_1636,In_537,In_1285);
nor U1637 (N_1637,In_326,In_1249);
nor U1638 (N_1638,In_1106,In_888);
or U1639 (N_1639,In_1888,In_239);
or U1640 (N_1640,In_1906,In_1272);
and U1641 (N_1641,In_356,In_1376);
and U1642 (N_1642,In_1039,In_559);
nor U1643 (N_1643,In_484,In_1424);
or U1644 (N_1644,In_1109,In_569);
and U1645 (N_1645,In_1335,In_1217);
or U1646 (N_1646,In_328,In_428);
or U1647 (N_1647,In_1346,In_909);
nand U1648 (N_1648,In_706,In_1783);
nand U1649 (N_1649,In_1048,In_1718);
or U1650 (N_1650,In_240,In_339);
nand U1651 (N_1651,In_1487,In_160);
or U1652 (N_1652,In_1283,In_1293);
and U1653 (N_1653,In_1368,In_940);
nor U1654 (N_1654,In_921,In_1723);
nand U1655 (N_1655,In_1714,In_79);
and U1656 (N_1656,In_575,In_364);
xor U1657 (N_1657,In_69,In_463);
nor U1658 (N_1658,In_993,In_794);
nor U1659 (N_1659,In_45,In_587);
nor U1660 (N_1660,In_725,In_675);
nand U1661 (N_1661,In_1858,In_924);
nor U1662 (N_1662,In_1594,In_574);
nor U1663 (N_1663,In_1007,In_648);
and U1664 (N_1664,In_129,In_1607);
nor U1665 (N_1665,In_685,In_1120);
nor U1666 (N_1666,In_1621,In_1357);
nor U1667 (N_1667,In_43,In_604);
or U1668 (N_1668,In_168,In_330);
or U1669 (N_1669,In_263,In_1607);
nand U1670 (N_1670,In_320,In_528);
xor U1671 (N_1671,In_1272,In_1504);
and U1672 (N_1672,In_1840,In_975);
nand U1673 (N_1673,In_89,In_1561);
and U1674 (N_1674,In_422,In_1554);
nand U1675 (N_1675,In_364,In_1352);
or U1676 (N_1676,In_890,In_424);
or U1677 (N_1677,In_1180,In_525);
and U1678 (N_1678,In_1700,In_62);
or U1679 (N_1679,In_1930,In_818);
and U1680 (N_1680,In_572,In_1026);
nor U1681 (N_1681,In_1371,In_1367);
and U1682 (N_1682,In_899,In_695);
nand U1683 (N_1683,In_1365,In_599);
nand U1684 (N_1684,In_812,In_349);
nor U1685 (N_1685,In_1122,In_1267);
xnor U1686 (N_1686,In_1685,In_343);
nand U1687 (N_1687,In_493,In_704);
nor U1688 (N_1688,In_1557,In_566);
nand U1689 (N_1689,In_701,In_1635);
nand U1690 (N_1690,In_1721,In_835);
or U1691 (N_1691,In_1483,In_1300);
or U1692 (N_1692,In_1658,In_1021);
or U1693 (N_1693,In_953,In_1479);
or U1694 (N_1694,In_367,In_1535);
nand U1695 (N_1695,In_1031,In_1951);
or U1696 (N_1696,In_1821,In_1444);
or U1697 (N_1697,In_1854,In_665);
nor U1698 (N_1698,In_1239,In_1376);
or U1699 (N_1699,In_646,In_747);
nor U1700 (N_1700,In_1676,In_1178);
and U1701 (N_1701,In_151,In_1988);
nand U1702 (N_1702,In_370,In_199);
or U1703 (N_1703,In_1067,In_1052);
and U1704 (N_1704,In_1329,In_286);
nand U1705 (N_1705,In_709,In_1924);
or U1706 (N_1706,In_537,In_1804);
nand U1707 (N_1707,In_338,In_345);
nand U1708 (N_1708,In_820,In_1381);
nor U1709 (N_1709,In_1802,In_1524);
and U1710 (N_1710,In_46,In_34);
or U1711 (N_1711,In_1431,In_848);
and U1712 (N_1712,In_1171,In_659);
or U1713 (N_1713,In_130,In_923);
nor U1714 (N_1714,In_1929,In_792);
and U1715 (N_1715,In_1086,In_1657);
nand U1716 (N_1716,In_389,In_653);
nor U1717 (N_1717,In_421,In_494);
nand U1718 (N_1718,In_1821,In_204);
and U1719 (N_1719,In_790,In_1049);
nand U1720 (N_1720,In_815,In_506);
nand U1721 (N_1721,In_1724,In_1137);
and U1722 (N_1722,In_1086,In_944);
nand U1723 (N_1723,In_1184,In_1037);
nor U1724 (N_1724,In_282,In_1005);
nor U1725 (N_1725,In_344,In_37);
nand U1726 (N_1726,In_165,In_172);
and U1727 (N_1727,In_1417,In_1486);
and U1728 (N_1728,In_313,In_1413);
nand U1729 (N_1729,In_13,In_1448);
nor U1730 (N_1730,In_618,In_1083);
nand U1731 (N_1731,In_63,In_1563);
and U1732 (N_1732,In_1870,In_708);
nand U1733 (N_1733,In_915,In_837);
nand U1734 (N_1734,In_520,In_1490);
xor U1735 (N_1735,In_103,In_1738);
nand U1736 (N_1736,In_1603,In_1855);
nor U1737 (N_1737,In_1130,In_961);
nor U1738 (N_1738,In_1239,In_707);
or U1739 (N_1739,In_124,In_1425);
and U1740 (N_1740,In_1325,In_561);
or U1741 (N_1741,In_612,In_1462);
xnor U1742 (N_1742,In_1717,In_727);
nand U1743 (N_1743,In_1139,In_378);
nand U1744 (N_1744,In_1959,In_530);
and U1745 (N_1745,In_1381,In_959);
and U1746 (N_1746,In_158,In_1689);
nor U1747 (N_1747,In_1942,In_72);
or U1748 (N_1748,In_1873,In_716);
nand U1749 (N_1749,In_523,In_466);
nand U1750 (N_1750,In_337,In_1465);
nand U1751 (N_1751,In_1365,In_385);
nor U1752 (N_1752,In_257,In_1717);
or U1753 (N_1753,In_1405,In_215);
nand U1754 (N_1754,In_39,In_429);
nor U1755 (N_1755,In_1534,In_373);
and U1756 (N_1756,In_1840,In_1052);
and U1757 (N_1757,In_1464,In_1584);
nand U1758 (N_1758,In_844,In_1562);
and U1759 (N_1759,In_1455,In_12);
xnor U1760 (N_1760,In_1393,In_1811);
nor U1761 (N_1761,In_656,In_208);
nand U1762 (N_1762,In_694,In_181);
and U1763 (N_1763,In_1562,In_1903);
nor U1764 (N_1764,In_1881,In_730);
nand U1765 (N_1765,In_545,In_405);
nand U1766 (N_1766,In_60,In_1055);
nor U1767 (N_1767,In_402,In_877);
and U1768 (N_1768,In_1337,In_1278);
nor U1769 (N_1769,In_367,In_237);
nand U1770 (N_1770,In_837,In_899);
nand U1771 (N_1771,In_1295,In_1391);
nor U1772 (N_1772,In_558,In_447);
nand U1773 (N_1773,In_302,In_1934);
and U1774 (N_1774,In_1745,In_1956);
or U1775 (N_1775,In_332,In_180);
nor U1776 (N_1776,In_968,In_1005);
nor U1777 (N_1777,In_437,In_169);
nor U1778 (N_1778,In_804,In_158);
nand U1779 (N_1779,In_436,In_756);
or U1780 (N_1780,In_1096,In_520);
or U1781 (N_1781,In_1516,In_1106);
nand U1782 (N_1782,In_1187,In_56);
nor U1783 (N_1783,In_375,In_1719);
and U1784 (N_1784,In_1150,In_672);
nand U1785 (N_1785,In_436,In_1645);
or U1786 (N_1786,In_491,In_968);
and U1787 (N_1787,In_1485,In_990);
xor U1788 (N_1788,In_1217,In_1550);
or U1789 (N_1789,In_1136,In_737);
or U1790 (N_1790,In_725,In_1146);
or U1791 (N_1791,In_1608,In_1584);
nor U1792 (N_1792,In_904,In_1351);
and U1793 (N_1793,In_1433,In_1370);
and U1794 (N_1794,In_430,In_321);
nor U1795 (N_1795,In_1120,In_1522);
nor U1796 (N_1796,In_1494,In_1784);
nand U1797 (N_1797,In_1684,In_1702);
or U1798 (N_1798,In_1430,In_517);
or U1799 (N_1799,In_1350,In_658);
and U1800 (N_1800,In_1987,In_1105);
nor U1801 (N_1801,In_3,In_713);
or U1802 (N_1802,In_180,In_1133);
nand U1803 (N_1803,In_543,In_547);
or U1804 (N_1804,In_1493,In_1318);
xnor U1805 (N_1805,In_920,In_1696);
nand U1806 (N_1806,In_932,In_1317);
and U1807 (N_1807,In_777,In_855);
nor U1808 (N_1808,In_499,In_1753);
nand U1809 (N_1809,In_1153,In_547);
and U1810 (N_1810,In_914,In_934);
nand U1811 (N_1811,In_1712,In_106);
or U1812 (N_1812,In_178,In_925);
and U1813 (N_1813,In_842,In_1646);
and U1814 (N_1814,In_1299,In_831);
nand U1815 (N_1815,In_1827,In_819);
nor U1816 (N_1816,In_450,In_789);
nor U1817 (N_1817,In_1400,In_1538);
nor U1818 (N_1818,In_1194,In_1735);
or U1819 (N_1819,In_426,In_1111);
or U1820 (N_1820,In_1704,In_1253);
and U1821 (N_1821,In_1652,In_1115);
and U1822 (N_1822,In_167,In_1446);
nand U1823 (N_1823,In_136,In_1116);
nand U1824 (N_1824,In_1515,In_1683);
or U1825 (N_1825,In_701,In_931);
or U1826 (N_1826,In_565,In_531);
nor U1827 (N_1827,In_48,In_1592);
or U1828 (N_1828,In_529,In_858);
nor U1829 (N_1829,In_1695,In_1827);
nor U1830 (N_1830,In_1095,In_1242);
and U1831 (N_1831,In_1840,In_215);
and U1832 (N_1832,In_189,In_1332);
nand U1833 (N_1833,In_1874,In_1643);
nor U1834 (N_1834,In_1149,In_215);
or U1835 (N_1835,In_1191,In_555);
or U1836 (N_1836,In_1394,In_1184);
nand U1837 (N_1837,In_1919,In_1585);
nand U1838 (N_1838,In_865,In_839);
and U1839 (N_1839,In_914,In_4);
or U1840 (N_1840,In_1571,In_1097);
or U1841 (N_1841,In_431,In_1333);
nand U1842 (N_1842,In_859,In_494);
and U1843 (N_1843,In_848,In_1862);
or U1844 (N_1844,In_755,In_519);
and U1845 (N_1845,In_1817,In_841);
nor U1846 (N_1846,In_72,In_226);
nor U1847 (N_1847,In_259,In_657);
nor U1848 (N_1848,In_1728,In_140);
and U1849 (N_1849,In_1659,In_836);
nand U1850 (N_1850,In_782,In_1621);
or U1851 (N_1851,In_1540,In_1372);
nand U1852 (N_1852,In_766,In_956);
nor U1853 (N_1853,In_1053,In_1238);
and U1854 (N_1854,In_1646,In_452);
and U1855 (N_1855,In_1031,In_733);
or U1856 (N_1856,In_885,In_1895);
and U1857 (N_1857,In_1172,In_1670);
nand U1858 (N_1858,In_1598,In_1870);
or U1859 (N_1859,In_903,In_950);
or U1860 (N_1860,In_1508,In_699);
nand U1861 (N_1861,In_1654,In_1984);
nand U1862 (N_1862,In_1598,In_1025);
and U1863 (N_1863,In_635,In_764);
and U1864 (N_1864,In_104,In_1419);
nand U1865 (N_1865,In_783,In_1614);
nor U1866 (N_1866,In_729,In_1751);
nand U1867 (N_1867,In_1935,In_1409);
nand U1868 (N_1868,In_1501,In_869);
xnor U1869 (N_1869,In_679,In_1351);
or U1870 (N_1870,In_1425,In_872);
nand U1871 (N_1871,In_682,In_243);
nor U1872 (N_1872,In_545,In_1174);
or U1873 (N_1873,In_1015,In_1550);
or U1874 (N_1874,In_1437,In_814);
and U1875 (N_1875,In_56,In_1099);
or U1876 (N_1876,In_48,In_1042);
xnor U1877 (N_1877,In_856,In_497);
or U1878 (N_1878,In_507,In_1271);
or U1879 (N_1879,In_1382,In_264);
or U1880 (N_1880,In_1405,In_1879);
nand U1881 (N_1881,In_590,In_259);
nand U1882 (N_1882,In_293,In_1719);
nor U1883 (N_1883,In_1360,In_989);
and U1884 (N_1884,In_1330,In_1094);
and U1885 (N_1885,In_1479,In_1876);
or U1886 (N_1886,In_1713,In_947);
or U1887 (N_1887,In_800,In_1873);
or U1888 (N_1888,In_1482,In_640);
or U1889 (N_1889,In_315,In_1900);
nor U1890 (N_1890,In_608,In_434);
nand U1891 (N_1891,In_64,In_1002);
nand U1892 (N_1892,In_1863,In_155);
and U1893 (N_1893,In_706,In_1478);
nand U1894 (N_1894,In_1855,In_479);
and U1895 (N_1895,In_1023,In_1283);
and U1896 (N_1896,In_580,In_281);
or U1897 (N_1897,In_779,In_170);
nor U1898 (N_1898,In_1423,In_1703);
nor U1899 (N_1899,In_1411,In_244);
nand U1900 (N_1900,In_18,In_141);
or U1901 (N_1901,In_1287,In_1892);
or U1902 (N_1902,In_1641,In_1259);
nand U1903 (N_1903,In_657,In_1162);
nand U1904 (N_1904,In_1894,In_918);
nand U1905 (N_1905,In_682,In_1646);
nand U1906 (N_1906,In_720,In_1098);
nand U1907 (N_1907,In_901,In_1051);
or U1908 (N_1908,In_1707,In_604);
or U1909 (N_1909,In_888,In_541);
nor U1910 (N_1910,In_205,In_4);
nand U1911 (N_1911,In_1455,In_379);
xnor U1912 (N_1912,In_65,In_1350);
nor U1913 (N_1913,In_984,In_1665);
or U1914 (N_1914,In_961,In_1538);
or U1915 (N_1915,In_537,In_368);
and U1916 (N_1916,In_930,In_1328);
nand U1917 (N_1917,In_1673,In_118);
or U1918 (N_1918,In_1896,In_1513);
and U1919 (N_1919,In_1400,In_1321);
and U1920 (N_1920,In_1826,In_1238);
nand U1921 (N_1921,In_330,In_226);
or U1922 (N_1922,In_899,In_1468);
and U1923 (N_1923,In_569,In_1686);
nor U1924 (N_1924,In_1793,In_920);
nand U1925 (N_1925,In_496,In_787);
nor U1926 (N_1926,In_401,In_192);
or U1927 (N_1927,In_1815,In_809);
and U1928 (N_1928,In_1422,In_1869);
nand U1929 (N_1929,In_1567,In_686);
nor U1930 (N_1930,In_1105,In_585);
or U1931 (N_1931,In_1050,In_545);
or U1932 (N_1932,In_763,In_469);
and U1933 (N_1933,In_551,In_1294);
nand U1934 (N_1934,In_720,In_725);
or U1935 (N_1935,In_1282,In_1443);
or U1936 (N_1936,In_1475,In_776);
or U1937 (N_1937,In_1876,In_1757);
nand U1938 (N_1938,In_1539,In_628);
nor U1939 (N_1939,In_1493,In_593);
nor U1940 (N_1940,In_1066,In_1840);
nand U1941 (N_1941,In_115,In_1248);
nor U1942 (N_1942,In_640,In_391);
or U1943 (N_1943,In_606,In_1327);
or U1944 (N_1944,In_1030,In_1998);
and U1945 (N_1945,In_1613,In_290);
and U1946 (N_1946,In_990,In_1145);
xnor U1947 (N_1947,In_67,In_1823);
nor U1948 (N_1948,In_667,In_763);
nand U1949 (N_1949,In_1806,In_31);
and U1950 (N_1950,In_127,In_1303);
nand U1951 (N_1951,In_817,In_1457);
nor U1952 (N_1952,In_910,In_1119);
nor U1953 (N_1953,In_1661,In_1657);
or U1954 (N_1954,In_1286,In_1964);
or U1955 (N_1955,In_690,In_645);
or U1956 (N_1956,In_774,In_1439);
or U1957 (N_1957,In_1066,In_852);
nand U1958 (N_1958,In_1142,In_1590);
nor U1959 (N_1959,In_1024,In_233);
nand U1960 (N_1960,In_1869,In_1972);
nand U1961 (N_1961,In_781,In_845);
nand U1962 (N_1962,In_1800,In_562);
nand U1963 (N_1963,In_573,In_468);
or U1964 (N_1964,In_673,In_1584);
and U1965 (N_1965,In_251,In_154);
and U1966 (N_1966,In_1392,In_1720);
nand U1967 (N_1967,In_1229,In_841);
and U1968 (N_1968,In_1249,In_1882);
and U1969 (N_1969,In_742,In_606);
nor U1970 (N_1970,In_735,In_1847);
nor U1971 (N_1971,In_1122,In_360);
and U1972 (N_1972,In_1024,In_1502);
and U1973 (N_1973,In_327,In_1747);
nand U1974 (N_1974,In_1388,In_1011);
nor U1975 (N_1975,In_193,In_1621);
nand U1976 (N_1976,In_318,In_1270);
and U1977 (N_1977,In_276,In_253);
nor U1978 (N_1978,In_427,In_1508);
and U1979 (N_1979,In_691,In_268);
nand U1980 (N_1980,In_1801,In_1819);
and U1981 (N_1981,In_1136,In_1584);
or U1982 (N_1982,In_1995,In_841);
and U1983 (N_1983,In_311,In_1105);
or U1984 (N_1984,In_933,In_875);
or U1985 (N_1985,In_1026,In_221);
and U1986 (N_1986,In_1614,In_910);
and U1987 (N_1987,In_915,In_1243);
nor U1988 (N_1988,In_924,In_1978);
or U1989 (N_1989,In_1696,In_144);
nand U1990 (N_1990,In_1226,In_592);
nand U1991 (N_1991,In_912,In_1845);
nand U1992 (N_1992,In_1554,In_956);
and U1993 (N_1993,In_1500,In_1339);
and U1994 (N_1994,In_1697,In_113);
nand U1995 (N_1995,In_158,In_1461);
and U1996 (N_1996,In_1074,In_1734);
or U1997 (N_1997,In_973,In_1079);
nor U1998 (N_1998,In_1418,In_1971);
and U1999 (N_1999,In_1675,In_939);
and U2000 (N_2000,In_1902,In_13);
nand U2001 (N_2001,In_1116,In_1605);
and U2002 (N_2002,In_1162,In_1754);
nor U2003 (N_2003,In_349,In_350);
nor U2004 (N_2004,In_645,In_1349);
nand U2005 (N_2005,In_446,In_1848);
nor U2006 (N_2006,In_1217,In_116);
and U2007 (N_2007,In_1052,In_1810);
nand U2008 (N_2008,In_563,In_0);
and U2009 (N_2009,In_438,In_195);
and U2010 (N_2010,In_679,In_1216);
nor U2011 (N_2011,In_271,In_1321);
or U2012 (N_2012,In_1334,In_1481);
or U2013 (N_2013,In_1992,In_18);
or U2014 (N_2014,In_396,In_1569);
or U2015 (N_2015,In_1860,In_817);
or U2016 (N_2016,In_496,In_1447);
nand U2017 (N_2017,In_1056,In_1507);
nor U2018 (N_2018,In_1135,In_933);
or U2019 (N_2019,In_1879,In_584);
and U2020 (N_2020,In_479,In_1572);
or U2021 (N_2021,In_366,In_747);
and U2022 (N_2022,In_1622,In_334);
or U2023 (N_2023,In_1169,In_1237);
nor U2024 (N_2024,In_29,In_961);
nand U2025 (N_2025,In_736,In_692);
nand U2026 (N_2026,In_478,In_1759);
nand U2027 (N_2027,In_579,In_1517);
nand U2028 (N_2028,In_1911,In_1976);
or U2029 (N_2029,In_324,In_633);
or U2030 (N_2030,In_720,In_128);
nor U2031 (N_2031,In_710,In_1842);
nand U2032 (N_2032,In_321,In_1058);
nand U2033 (N_2033,In_1443,In_194);
or U2034 (N_2034,In_14,In_749);
or U2035 (N_2035,In_819,In_743);
nand U2036 (N_2036,In_608,In_1045);
nor U2037 (N_2037,In_1206,In_229);
or U2038 (N_2038,In_667,In_1283);
or U2039 (N_2039,In_1167,In_1919);
nand U2040 (N_2040,In_1822,In_1808);
and U2041 (N_2041,In_1240,In_396);
and U2042 (N_2042,In_686,In_697);
nor U2043 (N_2043,In_592,In_1930);
nor U2044 (N_2044,In_963,In_580);
nand U2045 (N_2045,In_1861,In_1113);
nor U2046 (N_2046,In_1529,In_258);
nand U2047 (N_2047,In_73,In_1621);
nand U2048 (N_2048,In_812,In_834);
nor U2049 (N_2049,In_1036,In_499);
nor U2050 (N_2050,In_932,In_754);
nand U2051 (N_2051,In_179,In_1771);
and U2052 (N_2052,In_878,In_1500);
or U2053 (N_2053,In_1538,In_1383);
nor U2054 (N_2054,In_1474,In_1551);
or U2055 (N_2055,In_299,In_1634);
nand U2056 (N_2056,In_1830,In_1364);
and U2057 (N_2057,In_773,In_1654);
nor U2058 (N_2058,In_1595,In_1286);
or U2059 (N_2059,In_1167,In_1079);
or U2060 (N_2060,In_1672,In_1747);
nor U2061 (N_2061,In_1028,In_1607);
or U2062 (N_2062,In_454,In_996);
or U2063 (N_2063,In_1877,In_1661);
and U2064 (N_2064,In_1434,In_666);
or U2065 (N_2065,In_708,In_1338);
nand U2066 (N_2066,In_833,In_358);
or U2067 (N_2067,In_1104,In_1971);
nor U2068 (N_2068,In_425,In_323);
nor U2069 (N_2069,In_718,In_297);
nor U2070 (N_2070,In_868,In_1855);
and U2071 (N_2071,In_392,In_1036);
nand U2072 (N_2072,In_136,In_1099);
or U2073 (N_2073,In_1608,In_444);
nand U2074 (N_2074,In_1175,In_546);
nor U2075 (N_2075,In_1950,In_1220);
nor U2076 (N_2076,In_954,In_1155);
or U2077 (N_2077,In_1274,In_84);
nor U2078 (N_2078,In_1615,In_62);
and U2079 (N_2079,In_971,In_1962);
and U2080 (N_2080,In_1091,In_1150);
or U2081 (N_2081,In_1380,In_304);
nand U2082 (N_2082,In_1170,In_959);
and U2083 (N_2083,In_376,In_1732);
nor U2084 (N_2084,In_1048,In_502);
and U2085 (N_2085,In_1080,In_1730);
or U2086 (N_2086,In_38,In_592);
nor U2087 (N_2087,In_1178,In_1637);
nand U2088 (N_2088,In_1528,In_1691);
nand U2089 (N_2089,In_971,In_238);
nor U2090 (N_2090,In_514,In_263);
nor U2091 (N_2091,In_617,In_1280);
nand U2092 (N_2092,In_1911,In_1949);
nor U2093 (N_2093,In_1444,In_1634);
and U2094 (N_2094,In_83,In_1461);
and U2095 (N_2095,In_675,In_1838);
xor U2096 (N_2096,In_746,In_862);
or U2097 (N_2097,In_1017,In_585);
nor U2098 (N_2098,In_443,In_1627);
nand U2099 (N_2099,In_871,In_246);
or U2100 (N_2100,In_435,In_294);
or U2101 (N_2101,In_549,In_1992);
nor U2102 (N_2102,In_1061,In_196);
nand U2103 (N_2103,In_1853,In_986);
nand U2104 (N_2104,In_271,In_324);
nand U2105 (N_2105,In_863,In_1695);
nor U2106 (N_2106,In_1433,In_689);
nor U2107 (N_2107,In_1646,In_599);
nand U2108 (N_2108,In_1083,In_1278);
nand U2109 (N_2109,In_102,In_1817);
and U2110 (N_2110,In_1847,In_94);
nand U2111 (N_2111,In_1827,In_529);
and U2112 (N_2112,In_906,In_1642);
and U2113 (N_2113,In_1313,In_1377);
and U2114 (N_2114,In_1163,In_98);
nand U2115 (N_2115,In_871,In_1196);
or U2116 (N_2116,In_988,In_308);
and U2117 (N_2117,In_1792,In_869);
or U2118 (N_2118,In_1766,In_959);
nor U2119 (N_2119,In_1608,In_785);
or U2120 (N_2120,In_571,In_1942);
and U2121 (N_2121,In_1651,In_666);
nand U2122 (N_2122,In_1828,In_1262);
and U2123 (N_2123,In_1186,In_633);
nor U2124 (N_2124,In_1831,In_616);
and U2125 (N_2125,In_1212,In_548);
and U2126 (N_2126,In_1478,In_1507);
and U2127 (N_2127,In_447,In_560);
nand U2128 (N_2128,In_1159,In_121);
nor U2129 (N_2129,In_36,In_55);
and U2130 (N_2130,In_1932,In_491);
and U2131 (N_2131,In_922,In_1512);
nor U2132 (N_2132,In_1158,In_1837);
nor U2133 (N_2133,In_858,In_1106);
or U2134 (N_2134,In_1828,In_698);
or U2135 (N_2135,In_1424,In_1011);
nor U2136 (N_2136,In_1395,In_69);
nor U2137 (N_2137,In_1612,In_810);
nor U2138 (N_2138,In_277,In_491);
nor U2139 (N_2139,In_1258,In_1648);
and U2140 (N_2140,In_1613,In_385);
nor U2141 (N_2141,In_1790,In_271);
xnor U2142 (N_2142,In_1033,In_1944);
nand U2143 (N_2143,In_727,In_477);
and U2144 (N_2144,In_806,In_686);
or U2145 (N_2145,In_460,In_1405);
nor U2146 (N_2146,In_1414,In_1410);
or U2147 (N_2147,In_1156,In_1231);
nand U2148 (N_2148,In_1882,In_929);
nor U2149 (N_2149,In_1651,In_836);
and U2150 (N_2150,In_238,In_96);
or U2151 (N_2151,In_1124,In_135);
and U2152 (N_2152,In_1505,In_836);
nand U2153 (N_2153,In_1148,In_488);
nand U2154 (N_2154,In_1964,In_1411);
or U2155 (N_2155,In_44,In_346);
and U2156 (N_2156,In_1556,In_216);
nor U2157 (N_2157,In_1558,In_1281);
or U2158 (N_2158,In_968,In_1218);
nand U2159 (N_2159,In_1407,In_1372);
or U2160 (N_2160,In_1442,In_1411);
nand U2161 (N_2161,In_796,In_1533);
or U2162 (N_2162,In_1789,In_1564);
nand U2163 (N_2163,In_1245,In_958);
nand U2164 (N_2164,In_1849,In_888);
nand U2165 (N_2165,In_383,In_863);
nor U2166 (N_2166,In_737,In_1851);
or U2167 (N_2167,In_637,In_1770);
nand U2168 (N_2168,In_1061,In_1560);
nand U2169 (N_2169,In_12,In_1463);
and U2170 (N_2170,In_189,In_1473);
nor U2171 (N_2171,In_821,In_405);
and U2172 (N_2172,In_1115,In_1967);
and U2173 (N_2173,In_904,In_1077);
nor U2174 (N_2174,In_1495,In_679);
nor U2175 (N_2175,In_1781,In_276);
or U2176 (N_2176,In_112,In_1125);
and U2177 (N_2177,In_1053,In_1298);
or U2178 (N_2178,In_1327,In_1602);
or U2179 (N_2179,In_1367,In_1057);
nand U2180 (N_2180,In_1399,In_868);
nand U2181 (N_2181,In_49,In_1099);
nand U2182 (N_2182,In_42,In_1568);
or U2183 (N_2183,In_779,In_920);
or U2184 (N_2184,In_1397,In_550);
or U2185 (N_2185,In_6,In_531);
xor U2186 (N_2186,In_1527,In_1587);
and U2187 (N_2187,In_1040,In_636);
nor U2188 (N_2188,In_1935,In_410);
nor U2189 (N_2189,In_534,In_1203);
or U2190 (N_2190,In_643,In_1220);
or U2191 (N_2191,In_1307,In_448);
nand U2192 (N_2192,In_931,In_1318);
and U2193 (N_2193,In_450,In_463);
and U2194 (N_2194,In_237,In_592);
or U2195 (N_2195,In_264,In_480);
or U2196 (N_2196,In_415,In_788);
nand U2197 (N_2197,In_137,In_338);
nand U2198 (N_2198,In_1666,In_416);
nand U2199 (N_2199,In_1045,In_1103);
and U2200 (N_2200,In_733,In_357);
and U2201 (N_2201,In_51,In_1949);
nand U2202 (N_2202,In_288,In_582);
nor U2203 (N_2203,In_656,In_1826);
nor U2204 (N_2204,In_1764,In_21);
or U2205 (N_2205,In_1816,In_1584);
and U2206 (N_2206,In_152,In_1938);
or U2207 (N_2207,In_728,In_1589);
nor U2208 (N_2208,In_1846,In_541);
or U2209 (N_2209,In_1584,In_1514);
nor U2210 (N_2210,In_78,In_1107);
nor U2211 (N_2211,In_1364,In_1844);
or U2212 (N_2212,In_749,In_1846);
nor U2213 (N_2213,In_1232,In_1863);
and U2214 (N_2214,In_586,In_1301);
nor U2215 (N_2215,In_900,In_205);
or U2216 (N_2216,In_1216,In_1093);
and U2217 (N_2217,In_1931,In_657);
or U2218 (N_2218,In_1435,In_523);
nand U2219 (N_2219,In_1781,In_734);
or U2220 (N_2220,In_1175,In_758);
and U2221 (N_2221,In_1342,In_359);
nor U2222 (N_2222,In_194,In_1225);
nor U2223 (N_2223,In_919,In_413);
and U2224 (N_2224,In_993,In_1728);
and U2225 (N_2225,In_283,In_643);
nor U2226 (N_2226,In_1884,In_326);
nor U2227 (N_2227,In_216,In_1553);
nor U2228 (N_2228,In_289,In_140);
or U2229 (N_2229,In_945,In_859);
or U2230 (N_2230,In_240,In_1826);
and U2231 (N_2231,In_280,In_1605);
and U2232 (N_2232,In_1504,In_332);
nand U2233 (N_2233,In_329,In_1075);
and U2234 (N_2234,In_1895,In_1020);
nor U2235 (N_2235,In_239,In_1783);
or U2236 (N_2236,In_918,In_1194);
nor U2237 (N_2237,In_970,In_683);
nor U2238 (N_2238,In_1154,In_160);
or U2239 (N_2239,In_643,In_1078);
and U2240 (N_2240,In_584,In_1388);
and U2241 (N_2241,In_149,In_406);
or U2242 (N_2242,In_792,In_1605);
xnor U2243 (N_2243,In_1798,In_1487);
nor U2244 (N_2244,In_331,In_698);
and U2245 (N_2245,In_1367,In_1456);
and U2246 (N_2246,In_1691,In_1765);
or U2247 (N_2247,In_1505,In_592);
nand U2248 (N_2248,In_13,In_1973);
or U2249 (N_2249,In_936,In_614);
nand U2250 (N_2250,In_724,In_561);
nand U2251 (N_2251,In_994,In_360);
nor U2252 (N_2252,In_1737,In_198);
and U2253 (N_2253,In_1295,In_150);
or U2254 (N_2254,In_1307,In_979);
nand U2255 (N_2255,In_1978,In_172);
nand U2256 (N_2256,In_7,In_1917);
and U2257 (N_2257,In_187,In_737);
or U2258 (N_2258,In_450,In_1353);
nand U2259 (N_2259,In_1737,In_1423);
and U2260 (N_2260,In_1660,In_1858);
or U2261 (N_2261,In_1297,In_1911);
or U2262 (N_2262,In_410,In_662);
nand U2263 (N_2263,In_1517,In_1460);
nand U2264 (N_2264,In_406,In_874);
nand U2265 (N_2265,In_1355,In_1898);
xor U2266 (N_2266,In_844,In_763);
or U2267 (N_2267,In_674,In_232);
nand U2268 (N_2268,In_1502,In_337);
nand U2269 (N_2269,In_1739,In_1205);
or U2270 (N_2270,In_1406,In_516);
nand U2271 (N_2271,In_193,In_631);
nand U2272 (N_2272,In_661,In_80);
nor U2273 (N_2273,In_1189,In_1057);
nor U2274 (N_2274,In_231,In_1024);
nor U2275 (N_2275,In_640,In_230);
or U2276 (N_2276,In_1208,In_1641);
or U2277 (N_2277,In_1241,In_1839);
nand U2278 (N_2278,In_1297,In_499);
nand U2279 (N_2279,In_201,In_1520);
nor U2280 (N_2280,In_410,In_1261);
nand U2281 (N_2281,In_1714,In_826);
nor U2282 (N_2282,In_181,In_642);
nor U2283 (N_2283,In_991,In_1377);
nor U2284 (N_2284,In_1448,In_497);
nand U2285 (N_2285,In_64,In_1633);
nand U2286 (N_2286,In_234,In_1173);
nor U2287 (N_2287,In_1799,In_1139);
nor U2288 (N_2288,In_1921,In_152);
and U2289 (N_2289,In_694,In_1813);
or U2290 (N_2290,In_21,In_607);
nand U2291 (N_2291,In_1088,In_406);
and U2292 (N_2292,In_1951,In_980);
and U2293 (N_2293,In_259,In_650);
nand U2294 (N_2294,In_394,In_1652);
nand U2295 (N_2295,In_281,In_180);
nand U2296 (N_2296,In_1519,In_1180);
nand U2297 (N_2297,In_797,In_756);
or U2298 (N_2298,In_638,In_731);
and U2299 (N_2299,In_1525,In_435);
or U2300 (N_2300,In_1851,In_698);
and U2301 (N_2301,In_1346,In_1964);
nor U2302 (N_2302,In_1610,In_1804);
nor U2303 (N_2303,In_1784,In_1461);
and U2304 (N_2304,In_1262,In_1016);
nor U2305 (N_2305,In_1588,In_1460);
nand U2306 (N_2306,In_665,In_1888);
or U2307 (N_2307,In_1691,In_313);
nor U2308 (N_2308,In_1971,In_1351);
nor U2309 (N_2309,In_1046,In_696);
nand U2310 (N_2310,In_1724,In_1589);
nor U2311 (N_2311,In_1774,In_1168);
nand U2312 (N_2312,In_1264,In_150);
nand U2313 (N_2313,In_352,In_953);
nand U2314 (N_2314,In_951,In_913);
and U2315 (N_2315,In_1758,In_477);
nor U2316 (N_2316,In_74,In_733);
nand U2317 (N_2317,In_509,In_430);
nand U2318 (N_2318,In_1639,In_332);
nand U2319 (N_2319,In_1527,In_734);
or U2320 (N_2320,In_1499,In_1416);
or U2321 (N_2321,In_1459,In_979);
or U2322 (N_2322,In_328,In_876);
and U2323 (N_2323,In_1058,In_130);
nand U2324 (N_2324,In_1088,In_295);
nor U2325 (N_2325,In_1373,In_7);
nor U2326 (N_2326,In_355,In_1939);
and U2327 (N_2327,In_1533,In_1822);
nand U2328 (N_2328,In_1624,In_1230);
or U2329 (N_2329,In_197,In_1009);
and U2330 (N_2330,In_425,In_370);
nand U2331 (N_2331,In_417,In_808);
or U2332 (N_2332,In_259,In_93);
nor U2333 (N_2333,In_35,In_135);
nand U2334 (N_2334,In_386,In_51);
or U2335 (N_2335,In_712,In_1781);
nor U2336 (N_2336,In_1374,In_744);
nor U2337 (N_2337,In_775,In_744);
or U2338 (N_2338,In_1540,In_253);
nand U2339 (N_2339,In_1478,In_1140);
nor U2340 (N_2340,In_1790,In_158);
and U2341 (N_2341,In_865,In_1526);
nor U2342 (N_2342,In_679,In_1279);
nand U2343 (N_2343,In_96,In_1666);
or U2344 (N_2344,In_307,In_898);
or U2345 (N_2345,In_715,In_362);
or U2346 (N_2346,In_520,In_146);
xor U2347 (N_2347,In_1492,In_511);
or U2348 (N_2348,In_971,In_1567);
or U2349 (N_2349,In_1247,In_314);
nand U2350 (N_2350,In_463,In_1230);
or U2351 (N_2351,In_919,In_1233);
and U2352 (N_2352,In_1436,In_659);
and U2353 (N_2353,In_1304,In_282);
or U2354 (N_2354,In_87,In_30);
and U2355 (N_2355,In_153,In_605);
or U2356 (N_2356,In_1245,In_972);
nand U2357 (N_2357,In_362,In_1387);
nor U2358 (N_2358,In_1756,In_1804);
nor U2359 (N_2359,In_1196,In_254);
and U2360 (N_2360,In_129,In_1905);
or U2361 (N_2361,In_1259,In_365);
and U2362 (N_2362,In_1273,In_865);
or U2363 (N_2363,In_301,In_44);
nand U2364 (N_2364,In_53,In_1876);
and U2365 (N_2365,In_843,In_824);
and U2366 (N_2366,In_833,In_753);
and U2367 (N_2367,In_1211,In_1550);
nand U2368 (N_2368,In_15,In_69);
or U2369 (N_2369,In_546,In_4);
nor U2370 (N_2370,In_1779,In_258);
or U2371 (N_2371,In_1050,In_88);
and U2372 (N_2372,In_1010,In_424);
nand U2373 (N_2373,In_1953,In_1502);
and U2374 (N_2374,In_1060,In_737);
nand U2375 (N_2375,In_892,In_67);
or U2376 (N_2376,In_712,In_1145);
nor U2377 (N_2377,In_896,In_602);
or U2378 (N_2378,In_44,In_1017);
or U2379 (N_2379,In_1483,In_734);
and U2380 (N_2380,In_1129,In_259);
nand U2381 (N_2381,In_548,In_120);
or U2382 (N_2382,In_621,In_1361);
and U2383 (N_2383,In_477,In_770);
nor U2384 (N_2384,In_745,In_1083);
and U2385 (N_2385,In_1460,In_179);
and U2386 (N_2386,In_725,In_59);
nor U2387 (N_2387,In_1766,In_1712);
or U2388 (N_2388,In_1436,In_1731);
nor U2389 (N_2389,In_1940,In_1942);
nor U2390 (N_2390,In_1754,In_12);
and U2391 (N_2391,In_398,In_1365);
or U2392 (N_2392,In_1119,In_971);
or U2393 (N_2393,In_1382,In_120);
nand U2394 (N_2394,In_1745,In_1496);
or U2395 (N_2395,In_1189,In_237);
and U2396 (N_2396,In_694,In_1902);
or U2397 (N_2397,In_1842,In_1681);
nor U2398 (N_2398,In_1073,In_1287);
or U2399 (N_2399,In_839,In_231);
nand U2400 (N_2400,In_831,In_1919);
nor U2401 (N_2401,In_662,In_813);
nor U2402 (N_2402,In_1941,In_239);
nand U2403 (N_2403,In_1369,In_436);
nand U2404 (N_2404,In_564,In_245);
nand U2405 (N_2405,In_1979,In_959);
nor U2406 (N_2406,In_1964,In_64);
xor U2407 (N_2407,In_532,In_1304);
nand U2408 (N_2408,In_1486,In_1535);
or U2409 (N_2409,In_1996,In_371);
or U2410 (N_2410,In_1002,In_492);
nand U2411 (N_2411,In_118,In_1376);
and U2412 (N_2412,In_1389,In_784);
and U2413 (N_2413,In_1313,In_85);
nor U2414 (N_2414,In_1039,In_1559);
or U2415 (N_2415,In_742,In_957);
or U2416 (N_2416,In_526,In_1853);
and U2417 (N_2417,In_1952,In_694);
nand U2418 (N_2418,In_711,In_49);
nand U2419 (N_2419,In_813,In_147);
nor U2420 (N_2420,In_154,In_744);
nand U2421 (N_2421,In_876,In_1870);
and U2422 (N_2422,In_636,In_1701);
or U2423 (N_2423,In_841,In_379);
nor U2424 (N_2424,In_29,In_1690);
nor U2425 (N_2425,In_1148,In_1278);
nand U2426 (N_2426,In_189,In_1281);
and U2427 (N_2427,In_542,In_571);
nor U2428 (N_2428,In_1748,In_206);
and U2429 (N_2429,In_240,In_682);
nor U2430 (N_2430,In_1284,In_374);
and U2431 (N_2431,In_1705,In_1640);
nor U2432 (N_2432,In_1244,In_1400);
nor U2433 (N_2433,In_1679,In_404);
and U2434 (N_2434,In_213,In_1244);
and U2435 (N_2435,In_395,In_363);
and U2436 (N_2436,In_1354,In_1396);
and U2437 (N_2437,In_1624,In_945);
nor U2438 (N_2438,In_1149,In_18);
nor U2439 (N_2439,In_115,In_699);
nor U2440 (N_2440,In_1349,In_1786);
nand U2441 (N_2441,In_59,In_27);
and U2442 (N_2442,In_24,In_1313);
and U2443 (N_2443,In_1563,In_141);
nand U2444 (N_2444,In_380,In_1129);
or U2445 (N_2445,In_446,In_885);
or U2446 (N_2446,In_1373,In_225);
nor U2447 (N_2447,In_198,In_1606);
nand U2448 (N_2448,In_1746,In_1108);
or U2449 (N_2449,In_756,In_1144);
nand U2450 (N_2450,In_863,In_1492);
and U2451 (N_2451,In_1442,In_1071);
xor U2452 (N_2452,In_1027,In_30);
and U2453 (N_2453,In_1091,In_358);
nand U2454 (N_2454,In_412,In_1830);
nor U2455 (N_2455,In_277,In_518);
nor U2456 (N_2456,In_346,In_41);
nand U2457 (N_2457,In_242,In_1850);
or U2458 (N_2458,In_1809,In_1718);
or U2459 (N_2459,In_954,In_1069);
nand U2460 (N_2460,In_887,In_493);
nand U2461 (N_2461,In_695,In_10);
and U2462 (N_2462,In_1185,In_1122);
nor U2463 (N_2463,In_521,In_1445);
nor U2464 (N_2464,In_1432,In_252);
or U2465 (N_2465,In_1392,In_891);
nor U2466 (N_2466,In_1306,In_1950);
nor U2467 (N_2467,In_458,In_1328);
or U2468 (N_2468,In_1679,In_1449);
and U2469 (N_2469,In_911,In_1065);
nor U2470 (N_2470,In_1872,In_65);
nand U2471 (N_2471,In_1576,In_1224);
nor U2472 (N_2472,In_1774,In_1293);
nand U2473 (N_2473,In_1158,In_1804);
or U2474 (N_2474,In_769,In_1259);
or U2475 (N_2475,In_791,In_1282);
nand U2476 (N_2476,In_361,In_72);
nand U2477 (N_2477,In_668,In_601);
or U2478 (N_2478,In_120,In_386);
nand U2479 (N_2479,In_1377,In_838);
nand U2480 (N_2480,In_1955,In_453);
nand U2481 (N_2481,In_1675,In_1374);
and U2482 (N_2482,In_309,In_970);
or U2483 (N_2483,In_700,In_1170);
or U2484 (N_2484,In_1253,In_1453);
or U2485 (N_2485,In_622,In_1536);
or U2486 (N_2486,In_888,In_135);
and U2487 (N_2487,In_475,In_1854);
and U2488 (N_2488,In_1995,In_1344);
nand U2489 (N_2489,In_186,In_268);
nor U2490 (N_2490,In_238,In_1733);
nor U2491 (N_2491,In_1450,In_1962);
nor U2492 (N_2492,In_555,In_1753);
or U2493 (N_2493,In_1222,In_340);
nor U2494 (N_2494,In_1233,In_1768);
nor U2495 (N_2495,In_1441,In_1478);
and U2496 (N_2496,In_626,In_279);
nor U2497 (N_2497,In_301,In_1712);
and U2498 (N_2498,In_134,In_1635);
xnor U2499 (N_2499,In_52,In_1743);
or U2500 (N_2500,In_1983,In_96);
nand U2501 (N_2501,In_1099,In_1818);
and U2502 (N_2502,In_1101,In_1693);
and U2503 (N_2503,In_168,In_1983);
nand U2504 (N_2504,In_1643,In_1930);
nor U2505 (N_2505,In_1853,In_1888);
and U2506 (N_2506,In_269,In_308);
or U2507 (N_2507,In_75,In_1236);
and U2508 (N_2508,In_583,In_494);
or U2509 (N_2509,In_463,In_549);
or U2510 (N_2510,In_321,In_1782);
nand U2511 (N_2511,In_460,In_348);
or U2512 (N_2512,In_873,In_292);
nor U2513 (N_2513,In_859,In_1821);
nand U2514 (N_2514,In_1566,In_1616);
nor U2515 (N_2515,In_225,In_1567);
nor U2516 (N_2516,In_1560,In_1432);
nor U2517 (N_2517,In_10,In_547);
nor U2518 (N_2518,In_527,In_656);
nand U2519 (N_2519,In_832,In_438);
or U2520 (N_2520,In_921,In_728);
nor U2521 (N_2521,In_377,In_954);
or U2522 (N_2522,In_417,In_881);
and U2523 (N_2523,In_1984,In_1300);
and U2524 (N_2524,In_57,In_88);
and U2525 (N_2525,In_175,In_747);
and U2526 (N_2526,In_302,In_1803);
nor U2527 (N_2527,In_1298,In_1744);
or U2528 (N_2528,In_1640,In_1798);
nand U2529 (N_2529,In_830,In_1319);
and U2530 (N_2530,In_29,In_794);
or U2531 (N_2531,In_1770,In_1738);
and U2532 (N_2532,In_727,In_363);
and U2533 (N_2533,In_622,In_172);
nor U2534 (N_2534,In_366,In_876);
and U2535 (N_2535,In_458,In_1936);
nor U2536 (N_2536,In_1549,In_723);
or U2537 (N_2537,In_1764,In_1637);
nor U2538 (N_2538,In_1182,In_1068);
nand U2539 (N_2539,In_1416,In_1648);
nor U2540 (N_2540,In_643,In_1393);
and U2541 (N_2541,In_852,In_111);
or U2542 (N_2542,In_124,In_1286);
nand U2543 (N_2543,In_1919,In_1109);
nor U2544 (N_2544,In_1394,In_168);
nor U2545 (N_2545,In_1607,In_1012);
or U2546 (N_2546,In_1437,In_1120);
and U2547 (N_2547,In_829,In_1583);
nand U2548 (N_2548,In_1,In_1110);
nand U2549 (N_2549,In_765,In_583);
or U2550 (N_2550,In_609,In_849);
and U2551 (N_2551,In_1407,In_1006);
and U2552 (N_2552,In_1314,In_300);
and U2553 (N_2553,In_286,In_1068);
and U2554 (N_2554,In_37,In_1135);
nor U2555 (N_2555,In_1092,In_1317);
or U2556 (N_2556,In_1314,In_765);
and U2557 (N_2557,In_563,In_1997);
and U2558 (N_2558,In_1812,In_1681);
or U2559 (N_2559,In_1223,In_1053);
nor U2560 (N_2560,In_1601,In_514);
nor U2561 (N_2561,In_493,In_126);
and U2562 (N_2562,In_849,In_405);
and U2563 (N_2563,In_1210,In_1658);
or U2564 (N_2564,In_1165,In_1746);
or U2565 (N_2565,In_979,In_1591);
nand U2566 (N_2566,In_96,In_1718);
and U2567 (N_2567,In_153,In_1404);
nor U2568 (N_2568,In_1283,In_69);
nand U2569 (N_2569,In_1794,In_499);
or U2570 (N_2570,In_361,In_379);
nor U2571 (N_2571,In_747,In_1765);
and U2572 (N_2572,In_1181,In_485);
nand U2573 (N_2573,In_328,In_1345);
nand U2574 (N_2574,In_636,In_310);
nand U2575 (N_2575,In_1846,In_987);
nor U2576 (N_2576,In_1007,In_708);
xnor U2577 (N_2577,In_805,In_281);
nand U2578 (N_2578,In_261,In_1261);
or U2579 (N_2579,In_332,In_1968);
nand U2580 (N_2580,In_1082,In_1417);
and U2581 (N_2581,In_379,In_606);
or U2582 (N_2582,In_1951,In_152);
nand U2583 (N_2583,In_1724,In_236);
and U2584 (N_2584,In_1396,In_191);
nor U2585 (N_2585,In_1768,In_843);
nand U2586 (N_2586,In_504,In_659);
and U2587 (N_2587,In_85,In_815);
and U2588 (N_2588,In_1361,In_1854);
or U2589 (N_2589,In_1143,In_416);
nor U2590 (N_2590,In_962,In_209);
and U2591 (N_2591,In_984,In_1589);
and U2592 (N_2592,In_727,In_284);
nor U2593 (N_2593,In_1954,In_769);
and U2594 (N_2594,In_959,In_79);
xnor U2595 (N_2595,In_620,In_1127);
and U2596 (N_2596,In_37,In_794);
nor U2597 (N_2597,In_1536,In_1782);
nor U2598 (N_2598,In_1291,In_1365);
and U2599 (N_2599,In_1663,In_1660);
and U2600 (N_2600,In_599,In_1060);
nor U2601 (N_2601,In_1411,In_505);
nand U2602 (N_2602,In_1498,In_673);
xnor U2603 (N_2603,In_1724,In_1733);
nand U2604 (N_2604,In_583,In_437);
nand U2605 (N_2605,In_241,In_1988);
or U2606 (N_2606,In_11,In_1997);
and U2607 (N_2607,In_511,In_621);
and U2608 (N_2608,In_57,In_1283);
or U2609 (N_2609,In_1004,In_1019);
or U2610 (N_2610,In_1592,In_1891);
and U2611 (N_2611,In_255,In_117);
and U2612 (N_2612,In_1705,In_197);
nand U2613 (N_2613,In_1938,In_1920);
nor U2614 (N_2614,In_341,In_1636);
or U2615 (N_2615,In_619,In_1761);
and U2616 (N_2616,In_1411,In_1210);
or U2617 (N_2617,In_1099,In_1421);
nor U2618 (N_2618,In_1354,In_1465);
or U2619 (N_2619,In_1955,In_1112);
nor U2620 (N_2620,In_905,In_1220);
and U2621 (N_2621,In_208,In_666);
and U2622 (N_2622,In_856,In_855);
xnor U2623 (N_2623,In_341,In_647);
nor U2624 (N_2624,In_315,In_717);
and U2625 (N_2625,In_1713,In_1774);
and U2626 (N_2626,In_1700,In_993);
nor U2627 (N_2627,In_1049,In_378);
or U2628 (N_2628,In_1577,In_400);
and U2629 (N_2629,In_970,In_1034);
or U2630 (N_2630,In_808,In_327);
nor U2631 (N_2631,In_1230,In_654);
and U2632 (N_2632,In_1705,In_989);
nor U2633 (N_2633,In_1293,In_268);
and U2634 (N_2634,In_1039,In_487);
and U2635 (N_2635,In_1536,In_305);
nand U2636 (N_2636,In_498,In_298);
and U2637 (N_2637,In_265,In_164);
and U2638 (N_2638,In_827,In_1232);
nand U2639 (N_2639,In_904,In_1208);
nor U2640 (N_2640,In_542,In_234);
nor U2641 (N_2641,In_81,In_1084);
nor U2642 (N_2642,In_1570,In_1673);
nand U2643 (N_2643,In_60,In_1000);
nor U2644 (N_2644,In_1836,In_1695);
nand U2645 (N_2645,In_938,In_745);
and U2646 (N_2646,In_1247,In_933);
nor U2647 (N_2647,In_866,In_1196);
and U2648 (N_2648,In_1539,In_845);
or U2649 (N_2649,In_1168,In_1713);
nor U2650 (N_2650,In_1828,In_812);
and U2651 (N_2651,In_1326,In_372);
nand U2652 (N_2652,In_1641,In_1457);
and U2653 (N_2653,In_205,In_115);
or U2654 (N_2654,In_1767,In_1917);
and U2655 (N_2655,In_619,In_86);
nand U2656 (N_2656,In_683,In_1932);
and U2657 (N_2657,In_555,In_631);
nor U2658 (N_2658,In_58,In_716);
or U2659 (N_2659,In_1772,In_810);
and U2660 (N_2660,In_696,In_1876);
or U2661 (N_2661,In_175,In_1126);
or U2662 (N_2662,In_562,In_691);
xnor U2663 (N_2663,In_1846,In_685);
or U2664 (N_2664,In_1212,In_517);
or U2665 (N_2665,In_1530,In_1094);
or U2666 (N_2666,In_1171,In_1119);
nor U2667 (N_2667,In_1998,In_1412);
nor U2668 (N_2668,In_1060,In_626);
or U2669 (N_2669,In_161,In_1041);
or U2670 (N_2670,In_1364,In_15);
or U2671 (N_2671,In_117,In_857);
nand U2672 (N_2672,In_129,In_1810);
nor U2673 (N_2673,In_1216,In_1103);
and U2674 (N_2674,In_406,In_1126);
nand U2675 (N_2675,In_1417,In_1240);
and U2676 (N_2676,In_1986,In_204);
or U2677 (N_2677,In_1201,In_80);
nand U2678 (N_2678,In_600,In_379);
and U2679 (N_2679,In_58,In_245);
or U2680 (N_2680,In_110,In_1012);
nor U2681 (N_2681,In_37,In_311);
and U2682 (N_2682,In_88,In_1328);
or U2683 (N_2683,In_465,In_340);
and U2684 (N_2684,In_1840,In_834);
or U2685 (N_2685,In_248,In_1072);
nand U2686 (N_2686,In_1283,In_611);
nand U2687 (N_2687,In_282,In_1256);
nor U2688 (N_2688,In_1590,In_1527);
nand U2689 (N_2689,In_139,In_90);
nor U2690 (N_2690,In_618,In_1441);
nand U2691 (N_2691,In_1713,In_407);
and U2692 (N_2692,In_748,In_497);
or U2693 (N_2693,In_1565,In_881);
nand U2694 (N_2694,In_1631,In_1738);
and U2695 (N_2695,In_1784,In_926);
or U2696 (N_2696,In_837,In_1941);
and U2697 (N_2697,In_1189,In_1684);
nor U2698 (N_2698,In_1903,In_407);
and U2699 (N_2699,In_272,In_1755);
nand U2700 (N_2700,In_1717,In_265);
nand U2701 (N_2701,In_940,In_1522);
or U2702 (N_2702,In_1328,In_649);
nor U2703 (N_2703,In_1380,In_860);
or U2704 (N_2704,In_1258,In_651);
xnor U2705 (N_2705,In_1553,In_1107);
nor U2706 (N_2706,In_801,In_368);
nor U2707 (N_2707,In_899,In_1516);
and U2708 (N_2708,In_1243,In_275);
nand U2709 (N_2709,In_448,In_1309);
and U2710 (N_2710,In_642,In_40);
and U2711 (N_2711,In_268,In_1360);
and U2712 (N_2712,In_835,In_1585);
nand U2713 (N_2713,In_677,In_1214);
and U2714 (N_2714,In_811,In_1855);
and U2715 (N_2715,In_912,In_1814);
nand U2716 (N_2716,In_1181,In_304);
xnor U2717 (N_2717,In_1445,In_475);
or U2718 (N_2718,In_126,In_1681);
or U2719 (N_2719,In_1998,In_1085);
and U2720 (N_2720,In_182,In_155);
xnor U2721 (N_2721,In_136,In_1401);
nand U2722 (N_2722,In_1246,In_1958);
nand U2723 (N_2723,In_320,In_268);
or U2724 (N_2724,In_974,In_801);
or U2725 (N_2725,In_1243,In_322);
nand U2726 (N_2726,In_1500,In_643);
nor U2727 (N_2727,In_615,In_1181);
nand U2728 (N_2728,In_1113,In_42);
and U2729 (N_2729,In_1304,In_224);
nor U2730 (N_2730,In_1617,In_925);
or U2731 (N_2731,In_1406,In_1778);
nand U2732 (N_2732,In_386,In_1076);
nand U2733 (N_2733,In_206,In_1252);
and U2734 (N_2734,In_1066,In_1876);
nor U2735 (N_2735,In_219,In_1248);
and U2736 (N_2736,In_1029,In_347);
nor U2737 (N_2737,In_1753,In_1982);
xnor U2738 (N_2738,In_1311,In_1318);
nand U2739 (N_2739,In_1271,In_1817);
and U2740 (N_2740,In_1862,In_428);
and U2741 (N_2741,In_1374,In_1268);
nor U2742 (N_2742,In_1851,In_807);
nor U2743 (N_2743,In_1008,In_1871);
nand U2744 (N_2744,In_798,In_762);
nor U2745 (N_2745,In_1939,In_281);
nor U2746 (N_2746,In_479,In_837);
nor U2747 (N_2747,In_1552,In_1732);
or U2748 (N_2748,In_516,In_1470);
and U2749 (N_2749,In_794,In_945);
nor U2750 (N_2750,In_311,In_3);
and U2751 (N_2751,In_890,In_980);
nor U2752 (N_2752,In_694,In_1946);
and U2753 (N_2753,In_468,In_922);
nand U2754 (N_2754,In_539,In_974);
nand U2755 (N_2755,In_19,In_1620);
nor U2756 (N_2756,In_261,In_744);
or U2757 (N_2757,In_618,In_1774);
nor U2758 (N_2758,In_1244,In_910);
nand U2759 (N_2759,In_1335,In_1976);
nor U2760 (N_2760,In_954,In_1470);
nand U2761 (N_2761,In_1979,In_1748);
nand U2762 (N_2762,In_289,In_1736);
nand U2763 (N_2763,In_1373,In_27);
and U2764 (N_2764,In_197,In_1145);
and U2765 (N_2765,In_452,In_1180);
nand U2766 (N_2766,In_169,In_586);
or U2767 (N_2767,In_1764,In_295);
or U2768 (N_2768,In_1927,In_190);
and U2769 (N_2769,In_1841,In_1379);
or U2770 (N_2770,In_53,In_96);
or U2771 (N_2771,In_903,In_176);
or U2772 (N_2772,In_1160,In_1215);
or U2773 (N_2773,In_1426,In_953);
or U2774 (N_2774,In_421,In_194);
or U2775 (N_2775,In_1824,In_1600);
nor U2776 (N_2776,In_1437,In_1031);
nor U2777 (N_2777,In_1774,In_1413);
and U2778 (N_2778,In_1246,In_273);
nor U2779 (N_2779,In_1837,In_114);
or U2780 (N_2780,In_1230,In_567);
nand U2781 (N_2781,In_1193,In_330);
or U2782 (N_2782,In_1214,In_1655);
nor U2783 (N_2783,In_1238,In_1252);
nand U2784 (N_2784,In_704,In_43);
or U2785 (N_2785,In_764,In_1095);
and U2786 (N_2786,In_1745,In_239);
nand U2787 (N_2787,In_1014,In_1538);
nor U2788 (N_2788,In_358,In_1786);
nand U2789 (N_2789,In_705,In_627);
nand U2790 (N_2790,In_1568,In_1514);
or U2791 (N_2791,In_1484,In_403);
nor U2792 (N_2792,In_1592,In_1447);
and U2793 (N_2793,In_1531,In_191);
nor U2794 (N_2794,In_1835,In_1546);
or U2795 (N_2795,In_107,In_1);
nand U2796 (N_2796,In_1894,In_1219);
nor U2797 (N_2797,In_1790,In_598);
and U2798 (N_2798,In_1787,In_845);
or U2799 (N_2799,In_147,In_256);
nand U2800 (N_2800,In_1629,In_1493);
and U2801 (N_2801,In_1942,In_448);
nand U2802 (N_2802,In_106,In_1058);
nor U2803 (N_2803,In_1107,In_258);
or U2804 (N_2804,In_972,In_1667);
nor U2805 (N_2805,In_1392,In_933);
and U2806 (N_2806,In_1437,In_1989);
or U2807 (N_2807,In_790,In_1071);
or U2808 (N_2808,In_374,In_122);
and U2809 (N_2809,In_939,In_146);
or U2810 (N_2810,In_1115,In_1132);
nor U2811 (N_2811,In_530,In_344);
nor U2812 (N_2812,In_1294,In_1323);
and U2813 (N_2813,In_91,In_1631);
nor U2814 (N_2814,In_242,In_599);
and U2815 (N_2815,In_1135,In_675);
and U2816 (N_2816,In_1375,In_1272);
and U2817 (N_2817,In_1279,In_726);
and U2818 (N_2818,In_616,In_511);
nor U2819 (N_2819,In_738,In_1417);
or U2820 (N_2820,In_1089,In_1781);
nand U2821 (N_2821,In_1752,In_1541);
and U2822 (N_2822,In_143,In_1347);
nand U2823 (N_2823,In_730,In_302);
nor U2824 (N_2824,In_939,In_425);
nor U2825 (N_2825,In_1445,In_834);
or U2826 (N_2826,In_429,In_1204);
nor U2827 (N_2827,In_683,In_1369);
nor U2828 (N_2828,In_1689,In_264);
nor U2829 (N_2829,In_707,In_176);
nand U2830 (N_2830,In_714,In_203);
nor U2831 (N_2831,In_1526,In_602);
nand U2832 (N_2832,In_885,In_1481);
nand U2833 (N_2833,In_516,In_1936);
and U2834 (N_2834,In_919,In_678);
nand U2835 (N_2835,In_353,In_1131);
and U2836 (N_2836,In_1397,In_1630);
and U2837 (N_2837,In_699,In_5);
nor U2838 (N_2838,In_1879,In_412);
nand U2839 (N_2839,In_1054,In_1214);
or U2840 (N_2840,In_1930,In_109);
nor U2841 (N_2841,In_1166,In_1295);
nor U2842 (N_2842,In_670,In_1840);
and U2843 (N_2843,In_1495,In_53);
nor U2844 (N_2844,In_1397,In_1902);
or U2845 (N_2845,In_701,In_1619);
nand U2846 (N_2846,In_1480,In_102);
and U2847 (N_2847,In_1727,In_1687);
nand U2848 (N_2848,In_751,In_948);
nor U2849 (N_2849,In_1188,In_970);
and U2850 (N_2850,In_1408,In_1153);
and U2851 (N_2851,In_543,In_643);
and U2852 (N_2852,In_1901,In_1767);
nor U2853 (N_2853,In_1090,In_1206);
and U2854 (N_2854,In_1476,In_179);
nand U2855 (N_2855,In_1055,In_199);
and U2856 (N_2856,In_1997,In_278);
or U2857 (N_2857,In_149,In_1447);
nand U2858 (N_2858,In_1161,In_1865);
and U2859 (N_2859,In_20,In_1575);
nor U2860 (N_2860,In_364,In_1782);
nand U2861 (N_2861,In_433,In_874);
nor U2862 (N_2862,In_956,In_362);
nor U2863 (N_2863,In_1403,In_1417);
or U2864 (N_2864,In_787,In_809);
nand U2865 (N_2865,In_1215,In_1156);
and U2866 (N_2866,In_386,In_1877);
or U2867 (N_2867,In_280,In_462);
and U2868 (N_2868,In_619,In_958);
nand U2869 (N_2869,In_1090,In_463);
and U2870 (N_2870,In_1167,In_1787);
and U2871 (N_2871,In_810,In_292);
nor U2872 (N_2872,In_1983,In_1950);
and U2873 (N_2873,In_1340,In_1442);
nor U2874 (N_2874,In_74,In_896);
nand U2875 (N_2875,In_364,In_1129);
and U2876 (N_2876,In_1967,In_290);
nor U2877 (N_2877,In_1970,In_771);
nor U2878 (N_2878,In_162,In_207);
nand U2879 (N_2879,In_1637,In_1231);
or U2880 (N_2880,In_1631,In_291);
or U2881 (N_2881,In_1904,In_358);
and U2882 (N_2882,In_1533,In_106);
nand U2883 (N_2883,In_1965,In_1505);
or U2884 (N_2884,In_1816,In_402);
nand U2885 (N_2885,In_1494,In_1407);
or U2886 (N_2886,In_1608,In_1092);
or U2887 (N_2887,In_1536,In_988);
and U2888 (N_2888,In_1518,In_1831);
nor U2889 (N_2889,In_294,In_1600);
nor U2890 (N_2890,In_1607,In_1279);
or U2891 (N_2891,In_918,In_1978);
nor U2892 (N_2892,In_764,In_1980);
nand U2893 (N_2893,In_1154,In_464);
nand U2894 (N_2894,In_564,In_1254);
nand U2895 (N_2895,In_1356,In_197);
or U2896 (N_2896,In_1871,In_673);
nand U2897 (N_2897,In_870,In_433);
nand U2898 (N_2898,In_1386,In_406);
and U2899 (N_2899,In_195,In_1874);
nor U2900 (N_2900,In_1419,In_275);
nor U2901 (N_2901,In_1202,In_829);
and U2902 (N_2902,In_562,In_458);
nand U2903 (N_2903,In_127,In_880);
nand U2904 (N_2904,In_1325,In_1327);
nor U2905 (N_2905,In_1929,In_1490);
nor U2906 (N_2906,In_1449,In_593);
and U2907 (N_2907,In_1615,In_1179);
and U2908 (N_2908,In_1342,In_477);
nand U2909 (N_2909,In_1780,In_1230);
and U2910 (N_2910,In_1404,In_1064);
nand U2911 (N_2911,In_1307,In_1922);
and U2912 (N_2912,In_386,In_306);
nor U2913 (N_2913,In_1617,In_1482);
and U2914 (N_2914,In_1797,In_866);
nand U2915 (N_2915,In_1079,In_308);
nand U2916 (N_2916,In_1845,In_1344);
nor U2917 (N_2917,In_926,In_567);
nand U2918 (N_2918,In_1302,In_543);
and U2919 (N_2919,In_1778,In_771);
and U2920 (N_2920,In_723,In_286);
or U2921 (N_2921,In_941,In_534);
nor U2922 (N_2922,In_475,In_870);
or U2923 (N_2923,In_1564,In_1231);
nand U2924 (N_2924,In_987,In_1762);
or U2925 (N_2925,In_63,In_184);
and U2926 (N_2926,In_599,In_1335);
or U2927 (N_2927,In_628,In_24);
nand U2928 (N_2928,In_132,In_148);
nor U2929 (N_2929,In_1011,In_863);
or U2930 (N_2930,In_924,In_837);
or U2931 (N_2931,In_47,In_958);
nand U2932 (N_2932,In_1513,In_547);
or U2933 (N_2933,In_464,In_432);
and U2934 (N_2934,In_101,In_1781);
nor U2935 (N_2935,In_20,In_1185);
nand U2936 (N_2936,In_92,In_967);
or U2937 (N_2937,In_141,In_540);
nand U2938 (N_2938,In_583,In_983);
nand U2939 (N_2939,In_1898,In_1835);
nor U2940 (N_2940,In_1245,In_399);
and U2941 (N_2941,In_1553,In_1803);
or U2942 (N_2942,In_312,In_715);
and U2943 (N_2943,In_594,In_1268);
and U2944 (N_2944,In_554,In_1936);
and U2945 (N_2945,In_132,In_1132);
or U2946 (N_2946,In_1725,In_985);
or U2947 (N_2947,In_449,In_1717);
or U2948 (N_2948,In_581,In_804);
or U2949 (N_2949,In_586,In_88);
nand U2950 (N_2950,In_756,In_1808);
nor U2951 (N_2951,In_276,In_1375);
nor U2952 (N_2952,In_641,In_1014);
and U2953 (N_2953,In_312,In_280);
nand U2954 (N_2954,In_1645,In_327);
xor U2955 (N_2955,In_1128,In_1158);
and U2956 (N_2956,In_411,In_878);
nand U2957 (N_2957,In_1977,In_347);
nand U2958 (N_2958,In_1083,In_150);
nor U2959 (N_2959,In_1724,In_881);
nor U2960 (N_2960,In_1543,In_94);
or U2961 (N_2961,In_503,In_701);
and U2962 (N_2962,In_1363,In_97);
and U2963 (N_2963,In_1456,In_1670);
nand U2964 (N_2964,In_300,In_680);
and U2965 (N_2965,In_964,In_1465);
nor U2966 (N_2966,In_171,In_690);
nand U2967 (N_2967,In_1567,In_43);
nand U2968 (N_2968,In_1143,In_626);
nand U2969 (N_2969,In_867,In_828);
or U2970 (N_2970,In_1175,In_924);
nor U2971 (N_2971,In_100,In_1220);
nand U2972 (N_2972,In_1725,In_1987);
nand U2973 (N_2973,In_1829,In_125);
or U2974 (N_2974,In_1926,In_1996);
and U2975 (N_2975,In_1902,In_1525);
or U2976 (N_2976,In_1273,In_615);
and U2977 (N_2977,In_306,In_35);
nand U2978 (N_2978,In_1497,In_1133);
or U2979 (N_2979,In_573,In_622);
or U2980 (N_2980,In_1650,In_959);
nor U2981 (N_2981,In_1105,In_1447);
and U2982 (N_2982,In_1337,In_521);
nor U2983 (N_2983,In_640,In_1985);
nor U2984 (N_2984,In_1336,In_167);
or U2985 (N_2985,In_961,In_1492);
nand U2986 (N_2986,In_89,In_1285);
nor U2987 (N_2987,In_1860,In_15);
nor U2988 (N_2988,In_1146,In_418);
nor U2989 (N_2989,In_1337,In_1741);
nor U2990 (N_2990,In_800,In_442);
and U2991 (N_2991,In_1979,In_1355);
or U2992 (N_2992,In_647,In_885);
or U2993 (N_2993,In_524,In_74);
nor U2994 (N_2994,In_303,In_1498);
and U2995 (N_2995,In_537,In_581);
and U2996 (N_2996,In_874,In_890);
nand U2997 (N_2997,In_510,In_509);
nor U2998 (N_2998,In_521,In_483);
nand U2999 (N_2999,In_1902,In_139);
and U3000 (N_3000,In_1290,In_1300);
nand U3001 (N_3001,In_1859,In_1228);
xnor U3002 (N_3002,In_1545,In_1834);
nor U3003 (N_3003,In_909,In_955);
nor U3004 (N_3004,In_451,In_203);
or U3005 (N_3005,In_161,In_354);
and U3006 (N_3006,In_1651,In_576);
and U3007 (N_3007,In_80,In_448);
or U3008 (N_3008,In_423,In_1943);
nand U3009 (N_3009,In_527,In_485);
nand U3010 (N_3010,In_771,In_1444);
and U3011 (N_3011,In_1349,In_789);
nor U3012 (N_3012,In_1555,In_797);
nor U3013 (N_3013,In_1378,In_839);
nor U3014 (N_3014,In_1248,In_1979);
nand U3015 (N_3015,In_1512,In_1794);
nand U3016 (N_3016,In_553,In_1112);
nand U3017 (N_3017,In_615,In_880);
xnor U3018 (N_3018,In_288,In_1123);
nor U3019 (N_3019,In_848,In_1375);
nand U3020 (N_3020,In_277,In_1408);
nor U3021 (N_3021,In_1294,In_649);
nand U3022 (N_3022,In_1506,In_302);
nor U3023 (N_3023,In_1351,In_1615);
nor U3024 (N_3024,In_1359,In_1113);
nor U3025 (N_3025,In_575,In_1642);
or U3026 (N_3026,In_1082,In_1353);
nand U3027 (N_3027,In_59,In_1273);
nor U3028 (N_3028,In_1877,In_235);
and U3029 (N_3029,In_1872,In_1873);
and U3030 (N_3030,In_490,In_1297);
nand U3031 (N_3031,In_480,In_1450);
nand U3032 (N_3032,In_1407,In_209);
and U3033 (N_3033,In_1228,In_1489);
nand U3034 (N_3034,In_814,In_1641);
nand U3035 (N_3035,In_270,In_1153);
nand U3036 (N_3036,In_1409,In_1639);
nand U3037 (N_3037,In_1173,In_672);
nor U3038 (N_3038,In_1072,In_308);
nand U3039 (N_3039,In_276,In_403);
or U3040 (N_3040,In_846,In_1829);
nand U3041 (N_3041,In_280,In_122);
nor U3042 (N_3042,In_1453,In_640);
nor U3043 (N_3043,In_287,In_1119);
nand U3044 (N_3044,In_857,In_964);
nor U3045 (N_3045,In_120,In_1542);
nor U3046 (N_3046,In_1304,In_278);
and U3047 (N_3047,In_923,In_1761);
nor U3048 (N_3048,In_850,In_1033);
and U3049 (N_3049,In_230,In_1372);
and U3050 (N_3050,In_1925,In_87);
or U3051 (N_3051,In_1012,In_1311);
nand U3052 (N_3052,In_1728,In_1473);
and U3053 (N_3053,In_946,In_163);
and U3054 (N_3054,In_1911,In_1408);
nand U3055 (N_3055,In_1396,In_1881);
and U3056 (N_3056,In_384,In_1388);
nor U3057 (N_3057,In_532,In_732);
or U3058 (N_3058,In_475,In_1423);
xor U3059 (N_3059,In_1708,In_865);
nor U3060 (N_3060,In_1111,In_1793);
nor U3061 (N_3061,In_113,In_1872);
nand U3062 (N_3062,In_499,In_732);
and U3063 (N_3063,In_1554,In_862);
nor U3064 (N_3064,In_14,In_1632);
and U3065 (N_3065,In_1739,In_514);
nand U3066 (N_3066,In_384,In_1329);
nand U3067 (N_3067,In_865,In_1892);
and U3068 (N_3068,In_746,In_1457);
or U3069 (N_3069,In_1452,In_1054);
and U3070 (N_3070,In_382,In_1660);
nand U3071 (N_3071,In_1272,In_859);
or U3072 (N_3072,In_1365,In_1397);
nor U3073 (N_3073,In_224,In_1303);
or U3074 (N_3074,In_667,In_974);
or U3075 (N_3075,In_729,In_1512);
nor U3076 (N_3076,In_363,In_1781);
nor U3077 (N_3077,In_1475,In_1499);
and U3078 (N_3078,In_1897,In_169);
or U3079 (N_3079,In_1960,In_68);
nand U3080 (N_3080,In_1695,In_1401);
and U3081 (N_3081,In_1643,In_1689);
and U3082 (N_3082,In_1232,In_1943);
nor U3083 (N_3083,In_1061,In_1058);
and U3084 (N_3084,In_530,In_1676);
nor U3085 (N_3085,In_1128,In_1166);
and U3086 (N_3086,In_1165,In_968);
nor U3087 (N_3087,In_166,In_1347);
nand U3088 (N_3088,In_1829,In_1843);
and U3089 (N_3089,In_475,In_56);
nand U3090 (N_3090,In_688,In_1183);
nand U3091 (N_3091,In_897,In_719);
or U3092 (N_3092,In_884,In_1481);
and U3093 (N_3093,In_380,In_417);
or U3094 (N_3094,In_415,In_368);
and U3095 (N_3095,In_1657,In_627);
and U3096 (N_3096,In_709,In_1941);
nor U3097 (N_3097,In_53,In_1510);
or U3098 (N_3098,In_1335,In_1177);
nand U3099 (N_3099,In_1969,In_1597);
nor U3100 (N_3100,In_330,In_1208);
nand U3101 (N_3101,In_1190,In_229);
and U3102 (N_3102,In_583,In_1558);
nand U3103 (N_3103,In_1559,In_230);
nand U3104 (N_3104,In_1992,In_1289);
and U3105 (N_3105,In_1176,In_168);
and U3106 (N_3106,In_691,In_757);
nor U3107 (N_3107,In_1470,In_120);
nand U3108 (N_3108,In_461,In_1236);
nand U3109 (N_3109,In_1004,In_856);
and U3110 (N_3110,In_1791,In_1546);
nor U3111 (N_3111,In_310,In_832);
or U3112 (N_3112,In_1409,In_1957);
xnor U3113 (N_3113,In_1937,In_788);
nor U3114 (N_3114,In_1385,In_1293);
and U3115 (N_3115,In_387,In_876);
nor U3116 (N_3116,In_769,In_1649);
and U3117 (N_3117,In_680,In_92);
xor U3118 (N_3118,In_225,In_862);
nor U3119 (N_3119,In_143,In_51);
and U3120 (N_3120,In_564,In_584);
or U3121 (N_3121,In_776,In_1036);
or U3122 (N_3122,In_987,In_1750);
nand U3123 (N_3123,In_1989,In_241);
nand U3124 (N_3124,In_1175,In_94);
nand U3125 (N_3125,In_1371,In_1806);
or U3126 (N_3126,In_522,In_765);
nor U3127 (N_3127,In_695,In_1251);
nand U3128 (N_3128,In_1040,In_1867);
nor U3129 (N_3129,In_1173,In_993);
nor U3130 (N_3130,In_347,In_322);
nor U3131 (N_3131,In_706,In_1254);
and U3132 (N_3132,In_856,In_1090);
nor U3133 (N_3133,In_1295,In_1871);
nor U3134 (N_3134,In_1741,In_1540);
nor U3135 (N_3135,In_1209,In_1557);
and U3136 (N_3136,In_1119,In_269);
nor U3137 (N_3137,In_1300,In_284);
or U3138 (N_3138,In_1650,In_714);
and U3139 (N_3139,In_729,In_1866);
or U3140 (N_3140,In_182,In_1618);
and U3141 (N_3141,In_871,In_851);
and U3142 (N_3142,In_1909,In_1342);
or U3143 (N_3143,In_495,In_611);
and U3144 (N_3144,In_1812,In_85);
and U3145 (N_3145,In_1680,In_409);
or U3146 (N_3146,In_1160,In_57);
and U3147 (N_3147,In_456,In_1692);
and U3148 (N_3148,In_1115,In_948);
and U3149 (N_3149,In_1915,In_1606);
nor U3150 (N_3150,In_1453,In_1282);
or U3151 (N_3151,In_896,In_954);
nand U3152 (N_3152,In_36,In_253);
and U3153 (N_3153,In_162,In_1219);
and U3154 (N_3154,In_579,In_1410);
nor U3155 (N_3155,In_1458,In_1282);
nor U3156 (N_3156,In_1561,In_289);
nor U3157 (N_3157,In_337,In_1732);
or U3158 (N_3158,In_237,In_1082);
or U3159 (N_3159,In_824,In_1864);
nor U3160 (N_3160,In_1972,In_1655);
and U3161 (N_3161,In_1557,In_1115);
or U3162 (N_3162,In_689,In_201);
nand U3163 (N_3163,In_1780,In_211);
nor U3164 (N_3164,In_451,In_1528);
or U3165 (N_3165,In_1407,In_1887);
nand U3166 (N_3166,In_131,In_425);
or U3167 (N_3167,In_73,In_519);
and U3168 (N_3168,In_1580,In_672);
nor U3169 (N_3169,In_376,In_885);
or U3170 (N_3170,In_265,In_1853);
xnor U3171 (N_3171,In_1758,In_656);
nand U3172 (N_3172,In_1204,In_895);
or U3173 (N_3173,In_731,In_1896);
nor U3174 (N_3174,In_202,In_116);
and U3175 (N_3175,In_762,In_210);
and U3176 (N_3176,In_402,In_427);
nand U3177 (N_3177,In_1430,In_8);
and U3178 (N_3178,In_1254,In_1335);
and U3179 (N_3179,In_214,In_412);
nor U3180 (N_3180,In_1125,In_1842);
or U3181 (N_3181,In_21,In_1894);
and U3182 (N_3182,In_812,In_1371);
nand U3183 (N_3183,In_1915,In_1281);
nor U3184 (N_3184,In_1350,In_172);
nor U3185 (N_3185,In_1415,In_1661);
nand U3186 (N_3186,In_180,In_950);
nor U3187 (N_3187,In_1586,In_363);
nand U3188 (N_3188,In_824,In_197);
or U3189 (N_3189,In_242,In_1567);
nor U3190 (N_3190,In_239,In_1256);
nand U3191 (N_3191,In_992,In_661);
or U3192 (N_3192,In_363,In_366);
nand U3193 (N_3193,In_1575,In_1757);
nor U3194 (N_3194,In_1517,In_1891);
or U3195 (N_3195,In_764,In_69);
nand U3196 (N_3196,In_219,In_675);
and U3197 (N_3197,In_1422,In_501);
nor U3198 (N_3198,In_1967,In_1119);
nor U3199 (N_3199,In_1773,In_1829);
or U3200 (N_3200,In_684,In_1677);
nor U3201 (N_3201,In_612,In_1662);
and U3202 (N_3202,In_1037,In_1842);
or U3203 (N_3203,In_74,In_1469);
nand U3204 (N_3204,In_1223,In_1132);
nand U3205 (N_3205,In_1826,In_430);
or U3206 (N_3206,In_1088,In_194);
nand U3207 (N_3207,In_1626,In_1964);
nand U3208 (N_3208,In_431,In_1530);
or U3209 (N_3209,In_1061,In_1750);
and U3210 (N_3210,In_1255,In_1406);
and U3211 (N_3211,In_1334,In_691);
or U3212 (N_3212,In_1933,In_1889);
and U3213 (N_3213,In_430,In_127);
nand U3214 (N_3214,In_1859,In_1006);
nor U3215 (N_3215,In_292,In_995);
nor U3216 (N_3216,In_585,In_975);
nand U3217 (N_3217,In_1429,In_1049);
or U3218 (N_3218,In_755,In_467);
or U3219 (N_3219,In_103,In_852);
nor U3220 (N_3220,In_1859,In_1811);
nand U3221 (N_3221,In_355,In_873);
nor U3222 (N_3222,In_1699,In_1415);
nand U3223 (N_3223,In_939,In_517);
nor U3224 (N_3224,In_1015,In_1916);
nand U3225 (N_3225,In_877,In_86);
or U3226 (N_3226,In_127,In_1946);
and U3227 (N_3227,In_1813,In_1983);
and U3228 (N_3228,In_1323,In_1014);
nand U3229 (N_3229,In_1607,In_1921);
nor U3230 (N_3230,In_1629,In_1262);
or U3231 (N_3231,In_68,In_551);
nor U3232 (N_3232,In_362,In_667);
nand U3233 (N_3233,In_462,In_147);
nand U3234 (N_3234,In_1066,In_529);
nor U3235 (N_3235,In_1718,In_777);
or U3236 (N_3236,In_395,In_890);
nor U3237 (N_3237,In_1497,In_1484);
or U3238 (N_3238,In_1043,In_238);
xor U3239 (N_3239,In_1120,In_1217);
nand U3240 (N_3240,In_875,In_1529);
nand U3241 (N_3241,In_391,In_1958);
and U3242 (N_3242,In_1256,In_1705);
nor U3243 (N_3243,In_635,In_1627);
nand U3244 (N_3244,In_727,In_1748);
nor U3245 (N_3245,In_1992,In_943);
nand U3246 (N_3246,In_1569,In_125);
or U3247 (N_3247,In_860,In_1598);
or U3248 (N_3248,In_854,In_1388);
nor U3249 (N_3249,In_443,In_1769);
nor U3250 (N_3250,In_1994,In_1233);
nor U3251 (N_3251,In_765,In_105);
nand U3252 (N_3252,In_1886,In_545);
or U3253 (N_3253,In_425,In_775);
and U3254 (N_3254,In_1504,In_389);
or U3255 (N_3255,In_1106,In_1524);
or U3256 (N_3256,In_919,In_1140);
or U3257 (N_3257,In_1761,In_841);
or U3258 (N_3258,In_47,In_1787);
and U3259 (N_3259,In_1203,In_1321);
and U3260 (N_3260,In_851,In_1120);
and U3261 (N_3261,In_1183,In_56);
nor U3262 (N_3262,In_863,In_1187);
nand U3263 (N_3263,In_1590,In_1888);
nor U3264 (N_3264,In_1359,In_93);
nor U3265 (N_3265,In_1719,In_844);
xnor U3266 (N_3266,In_1132,In_428);
and U3267 (N_3267,In_1660,In_109);
or U3268 (N_3268,In_375,In_1463);
and U3269 (N_3269,In_1417,In_1691);
nand U3270 (N_3270,In_67,In_1363);
and U3271 (N_3271,In_584,In_1658);
nor U3272 (N_3272,In_717,In_1281);
or U3273 (N_3273,In_423,In_1466);
and U3274 (N_3274,In_1851,In_945);
or U3275 (N_3275,In_1311,In_522);
nand U3276 (N_3276,In_1986,In_307);
and U3277 (N_3277,In_765,In_177);
nand U3278 (N_3278,In_396,In_1588);
and U3279 (N_3279,In_1176,In_1416);
nor U3280 (N_3280,In_1967,In_800);
nand U3281 (N_3281,In_1622,In_1850);
nor U3282 (N_3282,In_1869,In_797);
nand U3283 (N_3283,In_412,In_1689);
nor U3284 (N_3284,In_202,In_872);
nor U3285 (N_3285,In_1620,In_985);
nand U3286 (N_3286,In_451,In_855);
nor U3287 (N_3287,In_411,In_681);
or U3288 (N_3288,In_1117,In_369);
and U3289 (N_3289,In_1334,In_845);
or U3290 (N_3290,In_812,In_910);
nand U3291 (N_3291,In_748,In_236);
nor U3292 (N_3292,In_4,In_1234);
nand U3293 (N_3293,In_623,In_612);
or U3294 (N_3294,In_1192,In_672);
or U3295 (N_3295,In_1122,In_1996);
or U3296 (N_3296,In_1844,In_1345);
nor U3297 (N_3297,In_1962,In_1245);
nor U3298 (N_3298,In_1114,In_1055);
or U3299 (N_3299,In_1664,In_1237);
or U3300 (N_3300,In_1532,In_357);
nor U3301 (N_3301,In_71,In_1173);
and U3302 (N_3302,In_90,In_1565);
or U3303 (N_3303,In_1383,In_1418);
and U3304 (N_3304,In_130,In_1200);
and U3305 (N_3305,In_959,In_449);
or U3306 (N_3306,In_211,In_1316);
or U3307 (N_3307,In_1306,In_1662);
or U3308 (N_3308,In_1164,In_1734);
nand U3309 (N_3309,In_708,In_360);
or U3310 (N_3310,In_1780,In_842);
or U3311 (N_3311,In_0,In_859);
or U3312 (N_3312,In_1433,In_629);
nor U3313 (N_3313,In_1155,In_346);
nor U3314 (N_3314,In_462,In_1561);
or U3315 (N_3315,In_1226,In_1228);
nand U3316 (N_3316,In_1009,In_1040);
nand U3317 (N_3317,In_1073,In_860);
or U3318 (N_3318,In_829,In_945);
nor U3319 (N_3319,In_1834,In_1613);
or U3320 (N_3320,In_1682,In_1398);
or U3321 (N_3321,In_816,In_387);
nor U3322 (N_3322,In_216,In_984);
nand U3323 (N_3323,In_670,In_911);
xnor U3324 (N_3324,In_782,In_1534);
or U3325 (N_3325,In_78,In_941);
nor U3326 (N_3326,In_59,In_315);
nor U3327 (N_3327,In_738,In_682);
nor U3328 (N_3328,In_1057,In_455);
or U3329 (N_3329,In_1399,In_1215);
and U3330 (N_3330,In_886,In_1085);
and U3331 (N_3331,In_1612,In_1188);
nand U3332 (N_3332,In_1772,In_502);
nor U3333 (N_3333,In_1609,In_752);
and U3334 (N_3334,In_567,In_528);
and U3335 (N_3335,In_865,In_1491);
nand U3336 (N_3336,In_115,In_263);
or U3337 (N_3337,In_1846,In_1670);
and U3338 (N_3338,In_776,In_55);
nor U3339 (N_3339,In_421,In_1488);
nor U3340 (N_3340,In_364,In_68);
nand U3341 (N_3341,In_414,In_836);
or U3342 (N_3342,In_1013,In_1001);
nand U3343 (N_3343,In_503,In_1679);
nand U3344 (N_3344,In_738,In_186);
nand U3345 (N_3345,In_670,In_879);
and U3346 (N_3346,In_24,In_880);
and U3347 (N_3347,In_250,In_1934);
and U3348 (N_3348,In_273,In_78);
or U3349 (N_3349,In_290,In_1939);
or U3350 (N_3350,In_1747,In_49);
and U3351 (N_3351,In_951,In_592);
nor U3352 (N_3352,In_385,In_1397);
and U3353 (N_3353,In_1726,In_157);
and U3354 (N_3354,In_1381,In_1440);
nor U3355 (N_3355,In_446,In_88);
nand U3356 (N_3356,In_666,In_1648);
nand U3357 (N_3357,In_1148,In_1940);
nor U3358 (N_3358,In_1322,In_1946);
nand U3359 (N_3359,In_1621,In_275);
nor U3360 (N_3360,In_1864,In_664);
and U3361 (N_3361,In_1144,In_527);
xnor U3362 (N_3362,In_1456,In_378);
nor U3363 (N_3363,In_299,In_137);
or U3364 (N_3364,In_232,In_658);
nand U3365 (N_3365,In_47,In_612);
nor U3366 (N_3366,In_1990,In_752);
or U3367 (N_3367,In_1804,In_1735);
nand U3368 (N_3368,In_1334,In_384);
and U3369 (N_3369,In_1849,In_827);
nand U3370 (N_3370,In_1805,In_1834);
nand U3371 (N_3371,In_841,In_1392);
nand U3372 (N_3372,In_686,In_1249);
or U3373 (N_3373,In_338,In_1638);
and U3374 (N_3374,In_524,In_1831);
or U3375 (N_3375,In_738,In_1321);
or U3376 (N_3376,In_616,In_1531);
or U3377 (N_3377,In_374,In_425);
nand U3378 (N_3378,In_1818,In_1558);
or U3379 (N_3379,In_1334,In_1281);
nor U3380 (N_3380,In_416,In_1114);
nand U3381 (N_3381,In_227,In_1338);
nand U3382 (N_3382,In_1154,In_799);
or U3383 (N_3383,In_1574,In_1470);
nand U3384 (N_3384,In_1806,In_1128);
and U3385 (N_3385,In_1181,In_0);
nand U3386 (N_3386,In_131,In_1793);
and U3387 (N_3387,In_1663,In_1819);
nor U3388 (N_3388,In_799,In_339);
nand U3389 (N_3389,In_1514,In_252);
nand U3390 (N_3390,In_1823,In_887);
and U3391 (N_3391,In_626,In_857);
nand U3392 (N_3392,In_620,In_1206);
or U3393 (N_3393,In_1275,In_692);
and U3394 (N_3394,In_918,In_898);
and U3395 (N_3395,In_1874,In_1282);
and U3396 (N_3396,In_798,In_1210);
nand U3397 (N_3397,In_192,In_39);
nor U3398 (N_3398,In_56,In_1157);
and U3399 (N_3399,In_1737,In_1976);
nand U3400 (N_3400,In_819,In_1415);
nand U3401 (N_3401,In_1646,In_670);
or U3402 (N_3402,In_402,In_1197);
or U3403 (N_3403,In_452,In_1152);
or U3404 (N_3404,In_1034,In_732);
nand U3405 (N_3405,In_709,In_120);
nor U3406 (N_3406,In_1006,In_1992);
or U3407 (N_3407,In_1365,In_1342);
nor U3408 (N_3408,In_1060,In_550);
nand U3409 (N_3409,In_1401,In_12);
or U3410 (N_3410,In_1276,In_372);
or U3411 (N_3411,In_1199,In_1830);
and U3412 (N_3412,In_1602,In_1028);
nand U3413 (N_3413,In_916,In_71);
nor U3414 (N_3414,In_694,In_1818);
nand U3415 (N_3415,In_18,In_97);
xnor U3416 (N_3416,In_1086,In_1225);
or U3417 (N_3417,In_1178,In_793);
nand U3418 (N_3418,In_330,In_1074);
nor U3419 (N_3419,In_250,In_478);
nand U3420 (N_3420,In_759,In_629);
or U3421 (N_3421,In_1212,In_1666);
and U3422 (N_3422,In_958,In_1734);
nand U3423 (N_3423,In_66,In_1396);
nor U3424 (N_3424,In_936,In_1983);
nor U3425 (N_3425,In_707,In_193);
or U3426 (N_3426,In_1006,In_891);
and U3427 (N_3427,In_1002,In_1003);
or U3428 (N_3428,In_498,In_242);
nor U3429 (N_3429,In_1256,In_834);
and U3430 (N_3430,In_838,In_1836);
and U3431 (N_3431,In_11,In_661);
nor U3432 (N_3432,In_362,In_1500);
and U3433 (N_3433,In_622,In_935);
or U3434 (N_3434,In_938,In_283);
or U3435 (N_3435,In_661,In_912);
and U3436 (N_3436,In_1024,In_928);
nand U3437 (N_3437,In_1123,In_355);
and U3438 (N_3438,In_641,In_1840);
nand U3439 (N_3439,In_1784,In_202);
and U3440 (N_3440,In_1405,In_1224);
and U3441 (N_3441,In_1901,In_865);
and U3442 (N_3442,In_1603,In_482);
and U3443 (N_3443,In_569,In_1462);
and U3444 (N_3444,In_1852,In_1203);
nand U3445 (N_3445,In_39,In_1915);
nand U3446 (N_3446,In_1286,In_1288);
and U3447 (N_3447,In_1378,In_344);
nor U3448 (N_3448,In_345,In_848);
and U3449 (N_3449,In_1831,In_1745);
nor U3450 (N_3450,In_1236,In_963);
nor U3451 (N_3451,In_742,In_1035);
nor U3452 (N_3452,In_1039,In_1908);
nand U3453 (N_3453,In_1033,In_1850);
or U3454 (N_3454,In_1110,In_1991);
or U3455 (N_3455,In_1033,In_665);
or U3456 (N_3456,In_1906,In_669);
nand U3457 (N_3457,In_937,In_763);
nor U3458 (N_3458,In_807,In_851);
nor U3459 (N_3459,In_140,In_1416);
nand U3460 (N_3460,In_1045,In_909);
or U3461 (N_3461,In_1281,In_1715);
nor U3462 (N_3462,In_1388,In_1591);
nand U3463 (N_3463,In_1059,In_1772);
and U3464 (N_3464,In_1647,In_475);
nand U3465 (N_3465,In_1429,In_933);
or U3466 (N_3466,In_614,In_1466);
nor U3467 (N_3467,In_47,In_549);
nor U3468 (N_3468,In_1224,In_1695);
or U3469 (N_3469,In_124,In_1852);
nand U3470 (N_3470,In_1670,In_228);
nor U3471 (N_3471,In_1402,In_154);
and U3472 (N_3472,In_0,In_2);
or U3473 (N_3473,In_1705,In_783);
nor U3474 (N_3474,In_485,In_768);
nand U3475 (N_3475,In_1887,In_792);
and U3476 (N_3476,In_29,In_972);
nand U3477 (N_3477,In_1293,In_1626);
and U3478 (N_3478,In_599,In_686);
or U3479 (N_3479,In_450,In_1349);
or U3480 (N_3480,In_1190,In_921);
nand U3481 (N_3481,In_277,In_1690);
nor U3482 (N_3482,In_1326,In_385);
and U3483 (N_3483,In_1818,In_1157);
or U3484 (N_3484,In_1088,In_687);
nor U3485 (N_3485,In_9,In_1475);
nor U3486 (N_3486,In_9,In_408);
and U3487 (N_3487,In_1875,In_1823);
and U3488 (N_3488,In_272,In_760);
nor U3489 (N_3489,In_1497,In_945);
and U3490 (N_3490,In_160,In_864);
and U3491 (N_3491,In_1878,In_1323);
nand U3492 (N_3492,In_1363,In_1929);
and U3493 (N_3493,In_1450,In_1536);
nor U3494 (N_3494,In_1290,In_441);
or U3495 (N_3495,In_676,In_520);
nand U3496 (N_3496,In_1438,In_629);
and U3497 (N_3497,In_1358,In_250);
nor U3498 (N_3498,In_1739,In_259);
nand U3499 (N_3499,In_640,In_609);
or U3500 (N_3500,In_1885,In_1365);
nand U3501 (N_3501,In_1665,In_1311);
nor U3502 (N_3502,In_1919,In_63);
or U3503 (N_3503,In_1864,In_885);
or U3504 (N_3504,In_1158,In_778);
nand U3505 (N_3505,In_1715,In_1015);
nand U3506 (N_3506,In_1393,In_1861);
nor U3507 (N_3507,In_1416,In_1158);
nand U3508 (N_3508,In_1529,In_1388);
nand U3509 (N_3509,In_1865,In_1962);
or U3510 (N_3510,In_554,In_1102);
nor U3511 (N_3511,In_1502,In_1893);
and U3512 (N_3512,In_371,In_646);
nor U3513 (N_3513,In_563,In_1808);
nor U3514 (N_3514,In_1589,In_502);
and U3515 (N_3515,In_835,In_826);
and U3516 (N_3516,In_1102,In_625);
or U3517 (N_3517,In_303,In_221);
or U3518 (N_3518,In_1107,In_1539);
nor U3519 (N_3519,In_310,In_1223);
and U3520 (N_3520,In_1362,In_130);
nand U3521 (N_3521,In_1839,In_1662);
nor U3522 (N_3522,In_529,In_1043);
nor U3523 (N_3523,In_117,In_397);
and U3524 (N_3524,In_967,In_1265);
nand U3525 (N_3525,In_819,In_1176);
nand U3526 (N_3526,In_802,In_33);
and U3527 (N_3527,In_1114,In_865);
nor U3528 (N_3528,In_1564,In_369);
and U3529 (N_3529,In_489,In_361);
nand U3530 (N_3530,In_1345,In_1181);
and U3531 (N_3531,In_490,In_1482);
nand U3532 (N_3532,In_1757,In_414);
nand U3533 (N_3533,In_8,In_1102);
nand U3534 (N_3534,In_891,In_324);
nor U3535 (N_3535,In_1778,In_109);
and U3536 (N_3536,In_1800,In_427);
or U3537 (N_3537,In_595,In_696);
nor U3538 (N_3538,In_1919,In_1927);
nand U3539 (N_3539,In_1035,In_1777);
or U3540 (N_3540,In_1526,In_270);
and U3541 (N_3541,In_1493,In_1671);
nand U3542 (N_3542,In_915,In_1831);
or U3543 (N_3543,In_725,In_1127);
nor U3544 (N_3544,In_1018,In_1839);
or U3545 (N_3545,In_1570,In_1794);
and U3546 (N_3546,In_1945,In_898);
and U3547 (N_3547,In_1303,In_104);
and U3548 (N_3548,In_851,In_265);
or U3549 (N_3549,In_307,In_873);
nor U3550 (N_3550,In_1875,In_460);
and U3551 (N_3551,In_1079,In_772);
nor U3552 (N_3552,In_441,In_310);
nand U3553 (N_3553,In_797,In_315);
nand U3554 (N_3554,In_426,In_320);
or U3555 (N_3555,In_724,In_1865);
nand U3556 (N_3556,In_1509,In_1860);
and U3557 (N_3557,In_1881,In_1218);
and U3558 (N_3558,In_1196,In_1435);
nand U3559 (N_3559,In_1729,In_822);
and U3560 (N_3560,In_1212,In_627);
and U3561 (N_3561,In_1601,In_1314);
or U3562 (N_3562,In_1646,In_178);
nand U3563 (N_3563,In_1900,In_301);
or U3564 (N_3564,In_151,In_523);
or U3565 (N_3565,In_1770,In_812);
and U3566 (N_3566,In_1587,In_1031);
or U3567 (N_3567,In_951,In_1590);
nor U3568 (N_3568,In_1174,In_687);
nand U3569 (N_3569,In_1397,In_1205);
nor U3570 (N_3570,In_1185,In_903);
nor U3571 (N_3571,In_648,In_202);
and U3572 (N_3572,In_419,In_1230);
and U3573 (N_3573,In_1758,In_1227);
nor U3574 (N_3574,In_1079,In_320);
nor U3575 (N_3575,In_129,In_1420);
or U3576 (N_3576,In_1383,In_349);
and U3577 (N_3577,In_1345,In_896);
or U3578 (N_3578,In_1909,In_854);
and U3579 (N_3579,In_1308,In_940);
nor U3580 (N_3580,In_591,In_674);
or U3581 (N_3581,In_1550,In_1545);
and U3582 (N_3582,In_1630,In_738);
nand U3583 (N_3583,In_844,In_1771);
or U3584 (N_3584,In_832,In_742);
nor U3585 (N_3585,In_445,In_363);
nand U3586 (N_3586,In_1367,In_1052);
and U3587 (N_3587,In_1870,In_1770);
nand U3588 (N_3588,In_216,In_1806);
and U3589 (N_3589,In_1571,In_1141);
nor U3590 (N_3590,In_932,In_777);
or U3591 (N_3591,In_172,In_6);
and U3592 (N_3592,In_713,In_1061);
and U3593 (N_3593,In_1497,In_851);
nor U3594 (N_3594,In_368,In_659);
or U3595 (N_3595,In_1407,In_1872);
nor U3596 (N_3596,In_694,In_1014);
nand U3597 (N_3597,In_77,In_1117);
and U3598 (N_3598,In_379,In_1933);
or U3599 (N_3599,In_1118,In_1710);
and U3600 (N_3600,In_653,In_301);
and U3601 (N_3601,In_157,In_1753);
nand U3602 (N_3602,In_1250,In_1813);
nand U3603 (N_3603,In_561,In_297);
nor U3604 (N_3604,In_700,In_955);
or U3605 (N_3605,In_1077,In_963);
and U3606 (N_3606,In_1121,In_1720);
xnor U3607 (N_3607,In_534,In_626);
and U3608 (N_3608,In_1895,In_1386);
nor U3609 (N_3609,In_1990,In_123);
nand U3610 (N_3610,In_1677,In_405);
or U3611 (N_3611,In_1606,In_329);
or U3612 (N_3612,In_1643,In_1371);
or U3613 (N_3613,In_1492,In_561);
or U3614 (N_3614,In_85,In_555);
nor U3615 (N_3615,In_1469,In_1483);
nor U3616 (N_3616,In_766,In_442);
nor U3617 (N_3617,In_1944,In_1863);
nor U3618 (N_3618,In_182,In_647);
nor U3619 (N_3619,In_1419,In_963);
nand U3620 (N_3620,In_1274,In_1361);
nand U3621 (N_3621,In_1336,In_765);
or U3622 (N_3622,In_1870,In_525);
nor U3623 (N_3623,In_537,In_1400);
and U3624 (N_3624,In_1653,In_1356);
nand U3625 (N_3625,In_385,In_801);
or U3626 (N_3626,In_446,In_1797);
nor U3627 (N_3627,In_1403,In_1128);
or U3628 (N_3628,In_614,In_689);
or U3629 (N_3629,In_1571,In_771);
and U3630 (N_3630,In_1663,In_225);
nor U3631 (N_3631,In_1500,In_447);
or U3632 (N_3632,In_61,In_304);
or U3633 (N_3633,In_1134,In_826);
nor U3634 (N_3634,In_119,In_1777);
xnor U3635 (N_3635,In_478,In_637);
nor U3636 (N_3636,In_1184,In_1565);
nor U3637 (N_3637,In_270,In_1769);
nor U3638 (N_3638,In_1088,In_357);
and U3639 (N_3639,In_1213,In_1);
nor U3640 (N_3640,In_1189,In_401);
and U3641 (N_3641,In_816,In_1898);
and U3642 (N_3642,In_1299,In_355);
xor U3643 (N_3643,In_1826,In_985);
nand U3644 (N_3644,In_1798,In_1486);
or U3645 (N_3645,In_503,In_1042);
nand U3646 (N_3646,In_495,In_1833);
or U3647 (N_3647,In_1564,In_1659);
or U3648 (N_3648,In_1120,In_1927);
nor U3649 (N_3649,In_1930,In_752);
nor U3650 (N_3650,In_1614,In_954);
and U3651 (N_3651,In_762,In_267);
or U3652 (N_3652,In_338,In_744);
nor U3653 (N_3653,In_480,In_1711);
nand U3654 (N_3654,In_22,In_71);
nor U3655 (N_3655,In_138,In_1875);
or U3656 (N_3656,In_538,In_970);
nor U3657 (N_3657,In_1936,In_1912);
nor U3658 (N_3658,In_160,In_193);
or U3659 (N_3659,In_1422,In_989);
or U3660 (N_3660,In_1062,In_1615);
or U3661 (N_3661,In_167,In_91);
and U3662 (N_3662,In_737,In_1321);
nor U3663 (N_3663,In_1198,In_817);
nor U3664 (N_3664,In_339,In_933);
or U3665 (N_3665,In_1691,In_1910);
nand U3666 (N_3666,In_1047,In_433);
xnor U3667 (N_3667,In_966,In_1239);
or U3668 (N_3668,In_1845,In_485);
and U3669 (N_3669,In_1429,In_1131);
and U3670 (N_3670,In_1632,In_1928);
nor U3671 (N_3671,In_1993,In_1041);
nor U3672 (N_3672,In_1202,In_1814);
or U3673 (N_3673,In_1431,In_9);
and U3674 (N_3674,In_768,In_164);
nor U3675 (N_3675,In_592,In_587);
and U3676 (N_3676,In_876,In_752);
and U3677 (N_3677,In_1539,In_386);
nand U3678 (N_3678,In_1966,In_277);
nand U3679 (N_3679,In_1616,In_1609);
nor U3680 (N_3680,In_1985,In_1129);
and U3681 (N_3681,In_213,In_1270);
nand U3682 (N_3682,In_113,In_431);
nor U3683 (N_3683,In_1218,In_624);
or U3684 (N_3684,In_495,In_109);
and U3685 (N_3685,In_1721,In_627);
nand U3686 (N_3686,In_702,In_366);
nand U3687 (N_3687,In_1290,In_988);
and U3688 (N_3688,In_126,In_1501);
nor U3689 (N_3689,In_1301,In_313);
and U3690 (N_3690,In_1663,In_1268);
and U3691 (N_3691,In_604,In_1384);
nor U3692 (N_3692,In_560,In_1086);
nand U3693 (N_3693,In_532,In_1758);
nand U3694 (N_3694,In_662,In_1693);
nor U3695 (N_3695,In_872,In_1118);
nand U3696 (N_3696,In_1584,In_1952);
or U3697 (N_3697,In_309,In_1431);
or U3698 (N_3698,In_866,In_1375);
and U3699 (N_3699,In_1231,In_325);
or U3700 (N_3700,In_1632,In_887);
nand U3701 (N_3701,In_1303,In_107);
nand U3702 (N_3702,In_530,In_608);
or U3703 (N_3703,In_1535,In_1069);
nand U3704 (N_3704,In_344,In_206);
and U3705 (N_3705,In_668,In_1343);
nand U3706 (N_3706,In_351,In_202);
or U3707 (N_3707,In_1161,In_952);
or U3708 (N_3708,In_220,In_1);
nand U3709 (N_3709,In_221,In_614);
nor U3710 (N_3710,In_1218,In_390);
and U3711 (N_3711,In_1677,In_1305);
or U3712 (N_3712,In_1924,In_1871);
and U3713 (N_3713,In_1535,In_1916);
and U3714 (N_3714,In_586,In_450);
nand U3715 (N_3715,In_500,In_1108);
nor U3716 (N_3716,In_498,In_1243);
and U3717 (N_3717,In_1844,In_69);
or U3718 (N_3718,In_1526,In_305);
and U3719 (N_3719,In_828,In_1245);
or U3720 (N_3720,In_524,In_781);
nand U3721 (N_3721,In_883,In_1871);
nor U3722 (N_3722,In_1635,In_966);
nand U3723 (N_3723,In_1925,In_1920);
or U3724 (N_3724,In_1906,In_1996);
and U3725 (N_3725,In_1157,In_535);
xnor U3726 (N_3726,In_48,In_288);
nand U3727 (N_3727,In_0,In_1445);
and U3728 (N_3728,In_1977,In_1253);
nor U3729 (N_3729,In_1448,In_644);
and U3730 (N_3730,In_295,In_1563);
and U3731 (N_3731,In_374,In_1560);
and U3732 (N_3732,In_417,In_818);
and U3733 (N_3733,In_1606,In_516);
and U3734 (N_3734,In_1460,In_434);
or U3735 (N_3735,In_560,In_1877);
nor U3736 (N_3736,In_1119,In_1907);
nor U3737 (N_3737,In_1453,In_1859);
or U3738 (N_3738,In_394,In_169);
or U3739 (N_3739,In_381,In_781);
or U3740 (N_3740,In_1185,In_1196);
and U3741 (N_3741,In_1991,In_361);
or U3742 (N_3742,In_1773,In_1531);
or U3743 (N_3743,In_938,In_1148);
nor U3744 (N_3744,In_206,In_540);
nor U3745 (N_3745,In_495,In_1653);
nand U3746 (N_3746,In_1006,In_1563);
and U3747 (N_3747,In_1775,In_759);
or U3748 (N_3748,In_1830,In_572);
nand U3749 (N_3749,In_584,In_1961);
and U3750 (N_3750,In_1286,In_1878);
and U3751 (N_3751,In_1467,In_1265);
and U3752 (N_3752,In_1934,In_1626);
nor U3753 (N_3753,In_1055,In_894);
nor U3754 (N_3754,In_788,In_1064);
nand U3755 (N_3755,In_1214,In_1331);
or U3756 (N_3756,In_879,In_1032);
nor U3757 (N_3757,In_395,In_782);
nor U3758 (N_3758,In_701,In_1787);
or U3759 (N_3759,In_563,In_1246);
and U3760 (N_3760,In_749,In_559);
nor U3761 (N_3761,In_497,In_1838);
and U3762 (N_3762,In_286,In_1927);
nor U3763 (N_3763,In_1988,In_804);
or U3764 (N_3764,In_1341,In_651);
or U3765 (N_3765,In_624,In_1417);
nand U3766 (N_3766,In_1471,In_968);
nand U3767 (N_3767,In_1989,In_33);
nand U3768 (N_3768,In_15,In_369);
nor U3769 (N_3769,In_1166,In_1900);
or U3770 (N_3770,In_1421,In_55);
nor U3771 (N_3771,In_145,In_1649);
nor U3772 (N_3772,In_1559,In_699);
xnor U3773 (N_3773,In_1271,In_969);
nor U3774 (N_3774,In_1443,In_999);
nor U3775 (N_3775,In_512,In_1627);
and U3776 (N_3776,In_1053,In_440);
nor U3777 (N_3777,In_834,In_1913);
nand U3778 (N_3778,In_1880,In_1033);
or U3779 (N_3779,In_140,In_736);
and U3780 (N_3780,In_1548,In_1484);
nand U3781 (N_3781,In_770,In_18);
nand U3782 (N_3782,In_1722,In_590);
nand U3783 (N_3783,In_3,In_449);
xnor U3784 (N_3784,In_678,In_490);
and U3785 (N_3785,In_1462,In_233);
and U3786 (N_3786,In_1422,In_1573);
and U3787 (N_3787,In_833,In_331);
nand U3788 (N_3788,In_877,In_1696);
nor U3789 (N_3789,In_197,In_1081);
nor U3790 (N_3790,In_1047,In_199);
nor U3791 (N_3791,In_1294,In_1523);
or U3792 (N_3792,In_409,In_1285);
and U3793 (N_3793,In_619,In_1227);
nand U3794 (N_3794,In_23,In_1974);
nor U3795 (N_3795,In_836,In_1449);
nand U3796 (N_3796,In_1424,In_824);
nor U3797 (N_3797,In_213,In_281);
nor U3798 (N_3798,In_1532,In_1912);
nand U3799 (N_3799,In_814,In_1967);
or U3800 (N_3800,In_1082,In_386);
and U3801 (N_3801,In_941,In_62);
nor U3802 (N_3802,In_1709,In_1453);
nor U3803 (N_3803,In_867,In_1142);
and U3804 (N_3804,In_1005,In_1032);
nor U3805 (N_3805,In_1879,In_1681);
or U3806 (N_3806,In_1338,In_517);
nand U3807 (N_3807,In_881,In_367);
or U3808 (N_3808,In_756,In_1244);
nor U3809 (N_3809,In_704,In_1183);
nand U3810 (N_3810,In_1042,In_899);
or U3811 (N_3811,In_1082,In_1963);
or U3812 (N_3812,In_1037,In_1514);
or U3813 (N_3813,In_194,In_1196);
or U3814 (N_3814,In_373,In_487);
nand U3815 (N_3815,In_288,In_1580);
nor U3816 (N_3816,In_732,In_81);
or U3817 (N_3817,In_157,In_1290);
nor U3818 (N_3818,In_1699,In_1289);
nor U3819 (N_3819,In_1805,In_1352);
nand U3820 (N_3820,In_758,In_714);
nor U3821 (N_3821,In_829,In_1019);
nand U3822 (N_3822,In_1368,In_1837);
and U3823 (N_3823,In_1020,In_1752);
or U3824 (N_3824,In_283,In_1281);
nor U3825 (N_3825,In_1464,In_46);
nor U3826 (N_3826,In_1421,In_1026);
nand U3827 (N_3827,In_570,In_1842);
nand U3828 (N_3828,In_1286,In_199);
nand U3829 (N_3829,In_1146,In_126);
nand U3830 (N_3830,In_1407,In_431);
nand U3831 (N_3831,In_1139,In_394);
nor U3832 (N_3832,In_501,In_1978);
nor U3833 (N_3833,In_1892,In_1481);
nor U3834 (N_3834,In_573,In_352);
nand U3835 (N_3835,In_1439,In_1954);
and U3836 (N_3836,In_214,In_1563);
and U3837 (N_3837,In_1209,In_1715);
and U3838 (N_3838,In_739,In_218);
nor U3839 (N_3839,In_236,In_495);
and U3840 (N_3840,In_275,In_492);
and U3841 (N_3841,In_1560,In_100);
nor U3842 (N_3842,In_1256,In_1369);
or U3843 (N_3843,In_1232,In_1983);
nor U3844 (N_3844,In_1803,In_709);
or U3845 (N_3845,In_1352,In_1656);
or U3846 (N_3846,In_1300,In_1096);
nor U3847 (N_3847,In_1086,In_87);
and U3848 (N_3848,In_208,In_876);
nor U3849 (N_3849,In_798,In_730);
nor U3850 (N_3850,In_1365,In_1585);
nor U3851 (N_3851,In_1946,In_637);
nor U3852 (N_3852,In_794,In_388);
nand U3853 (N_3853,In_1527,In_1019);
or U3854 (N_3854,In_1678,In_1716);
nor U3855 (N_3855,In_1478,In_641);
or U3856 (N_3856,In_908,In_1998);
nand U3857 (N_3857,In_617,In_674);
nor U3858 (N_3858,In_1925,In_380);
and U3859 (N_3859,In_1574,In_1583);
nand U3860 (N_3860,In_29,In_1379);
nor U3861 (N_3861,In_77,In_1793);
or U3862 (N_3862,In_403,In_1109);
nand U3863 (N_3863,In_228,In_1461);
nand U3864 (N_3864,In_562,In_26);
nor U3865 (N_3865,In_1603,In_1992);
nor U3866 (N_3866,In_1599,In_251);
and U3867 (N_3867,In_1379,In_195);
nand U3868 (N_3868,In_149,In_858);
nor U3869 (N_3869,In_289,In_1740);
or U3870 (N_3870,In_1645,In_9);
or U3871 (N_3871,In_774,In_1276);
nor U3872 (N_3872,In_1938,In_691);
nand U3873 (N_3873,In_270,In_1889);
nand U3874 (N_3874,In_1854,In_880);
nand U3875 (N_3875,In_112,In_1674);
and U3876 (N_3876,In_799,In_1058);
nand U3877 (N_3877,In_1616,In_1426);
or U3878 (N_3878,In_797,In_287);
nand U3879 (N_3879,In_1479,In_1705);
or U3880 (N_3880,In_1414,In_159);
nor U3881 (N_3881,In_178,In_325);
or U3882 (N_3882,In_756,In_248);
nand U3883 (N_3883,In_1482,In_1336);
and U3884 (N_3884,In_462,In_1566);
or U3885 (N_3885,In_726,In_352);
nand U3886 (N_3886,In_1920,In_1310);
and U3887 (N_3887,In_1613,In_771);
nand U3888 (N_3888,In_209,In_170);
nand U3889 (N_3889,In_962,In_1433);
xnor U3890 (N_3890,In_516,In_1105);
or U3891 (N_3891,In_1131,In_1606);
xor U3892 (N_3892,In_1129,In_1717);
nor U3893 (N_3893,In_1183,In_1005);
nand U3894 (N_3894,In_129,In_1004);
or U3895 (N_3895,In_544,In_1136);
nor U3896 (N_3896,In_50,In_569);
or U3897 (N_3897,In_508,In_781);
nor U3898 (N_3898,In_1509,In_1828);
nor U3899 (N_3899,In_741,In_1175);
nor U3900 (N_3900,In_1488,In_1776);
or U3901 (N_3901,In_1242,In_731);
and U3902 (N_3902,In_1372,In_1471);
and U3903 (N_3903,In_1196,In_580);
or U3904 (N_3904,In_1829,In_1455);
or U3905 (N_3905,In_1294,In_369);
nand U3906 (N_3906,In_396,In_1854);
nor U3907 (N_3907,In_728,In_1260);
nand U3908 (N_3908,In_942,In_541);
nand U3909 (N_3909,In_1423,In_1103);
nand U3910 (N_3910,In_1337,In_236);
nor U3911 (N_3911,In_17,In_1607);
nand U3912 (N_3912,In_920,In_1870);
nor U3913 (N_3913,In_985,In_59);
nor U3914 (N_3914,In_1784,In_603);
nand U3915 (N_3915,In_297,In_1808);
and U3916 (N_3916,In_1829,In_52);
nor U3917 (N_3917,In_767,In_96);
and U3918 (N_3918,In_1956,In_1962);
nor U3919 (N_3919,In_1066,In_1225);
nand U3920 (N_3920,In_462,In_1257);
nor U3921 (N_3921,In_877,In_100);
or U3922 (N_3922,In_662,In_1336);
nand U3923 (N_3923,In_215,In_415);
and U3924 (N_3924,In_43,In_1786);
or U3925 (N_3925,In_1102,In_101);
nand U3926 (N_3926,In_1241,In_1212);
or U3927 (N_3927,In_452,In_848);
and U3928 (N_3928,In_1956,In_349);
and U3929 (N_3929,In_940,In_394);
nand U3930 (N_3930,In_1931,In_1366);
nand U3931 (N_3931,In_578,In_612);
nand U3932 (N_3932,In_1795,In_598);
or U3933 (N_3933,In_95,In_337);
nand U3934 (N_3934,In_1317,In_1855);
nand U3935 (N_3935,In_1448,In_513);
or U3936 (N_3936,In_1641,In_1757);
or U3937 (N_3937,In_479,In_749);
and U3938 (N_3938,In_1413,In_1266);
or U3939 (N_3939,In_312,In_1810);
nand U3940 (N_3940,In_303,In_1005);
and U3941 (N_3941,In_865,In_1376);
or U3942 (N_3942,In_1881,In_1090);
nand U3943 (N_3943,In_1526,In_256);
or U3944 (N_3944,In_1674,In_1414);
and U3945 (N_3945,In_693,In_48);
nor U3946 (N_3946,In_501,In_1015);
nand U3947 (N_3947,In_239,In_389);
or U3948 (N_3948,In_1675,In_1281);
nand U3949 (N_3949,In_78,In_1453);
or U3950 (N_3950,In_895,In_913);
and U3951 (N_3951,In_396,In_1304);
nor U3952 (N_3952,In_290,In_517);
xor U3953 (N_3953,In_220,In_1009);
and U3954 (N_3954,In_563,In_91);
or U3955 (N_3955,In_878,In_1063);
nor U3956 (N_3956,In_240,In_1186);
nand U3957 (N_3957,In_1669,In_883);
and U3958 (N_3958,In_977,In_1486);
nand U3959 (N_3959,In_425,In_905);
nor U3960 (N_3960,In_1729,In_1715);
xnor U3961 (N_3961,In_317,In_969);
nand U3962 (N_3962,In_815,In_1706);
or U3963 (N_3963,In_1477,In_1819);
or U3964 (N_3964,In_1980,In_1173);
and U3965 (N_3965,In_497,In_1780);
and U3966 (N_3966,In_103,In_242);
nor U3967 (N_3967,In_1124,In_21);
nor U3968 (N_3968,In_527,In_1389);
and U3969 (N_3969,In_1579,In_755);
or U3970 (N_3970,In_293,In_1563);
or U3971 (N_3971,In_1206,In_869);
nand U3972 (N_3972,In_431,In_3);
nand U3973 (N_3973,In_1749,In_827);
or U3974 (N_3974,In_617,In_561);
nand U3975 (N_3975,In_232,In_1741);
nand U3976 (N_3976,In_1476,In_92);
nor U3977 (N_3977,In_1583,In_186);
and U3978 (N_3978,In_1503,In_1561);
nor U3979 (N_3979,In_894,In_327);
and U3980 (N_3980,In_122,In_922);
nand U3981 (N_3981,In_809,In_1264);
nand U3982 (N_3982,In_1385,In_1852);
nand U3983 (N_3983,In_1880,In_129);
nor U3984 (N_3984,In_691,In_1402);
or U3985 (N_3985,In_997,In_272);
nor U3986 (N_3986,In_827,In_1371);
and U3987 (N_3987,In_1936,In_1556);
or U3988 (N_3988,In_1696,In_79);
and U3989 (N_3989,In_1009,In_958);
nor U3990 (N_3990,In_170,In_1292);
or U3991 (N_3991,In_515,In_344);
and U3992 (N_3992,In_1839,In_906);
nor U3993 (N_3993,In_1192,In_1750);
or U3994 (N_3994,In_986,In_1098);
or U3995 (N_3995,In_1323,In_1813);
or U3996 (N_3996,In_1961,In_1440);
and U3997 (N_3997,In_1691,In_961);
and U3998 (N_3998,In_443,In_220);
nand U3999 (N_3999,In_753,In_1929);
nor U4000 (N_4000,N_3432,N_397);
nand U4001 (N_4001,N_3858,N_3528);
nand U4002 (N_4002,N_3225,N_2585);
nor U4003 (N_4003,N_1842,N_1799);
nand U4004 (N_4004,N_3940,N_3288);
nand U4005 (N_4005,N_1927,N_1600);
nand U4006 (N_4006,N_1581,N_947);
nor U4007 (N_4007,N_645,N_3354);
nand U4008 (N_4008,N_3058,N_1249);
nor U4009 (N_4009,N_3601,N_2308);
and U4010 (N_4010,N_2555,N_211);
or U4011 (N_4011,N_2867,N_898);
nand U4012 (N_4012,N_3254,N_3325);
nand U4013 (N_4013,N_3807,N_689);
nor U4014 (N_4014,N_3054,N_3646);
and U4015 (N_4015,N_3320,N_2068);
nor U4016 (N_4016,N_2352,N_3821);
nand U4017 (N_4017,N_2069,N_2616);
and U4018 (N_4018,N_3545,N_701);
or U4019 (N_4019,N_1533,N_493);
nand U4020 (N_4020,N_2674,N_1528);
nor U4021 (N_4021,N_3275,N_3612);
nand U4022 (N_4022,N_2956,N_86);
nand U4023 (N_4023,N_776,N_954);
nand U4024 (N_4024,N_2666,N_2770);
xor U4025 (N_4025,N_2428,N_2905);
nor U4026 (N_4026,N_404,N_1452);
nor U4027 (N_4027,N_2763,N_2544);
nand U4028 (N_4028,N_1252,N_3376);
nand U4029 (N_4029,N_1714,N_2590);
or U4030 (N_4030,N_3274,N_160);
nor U4031 (N_4031,N_639,N_2321);
or U4032 (N_4032,N_666,N_1626);
or U4033 (N_4033,N_1510,N_1782);
or U4034 (N_4034,N_909,N_1113);
nor U4035 (N_4035,N_1073,N_2021);
or U4036 (N_4036,N_1443,N_3890);
nand U4037 (N_4037,N_3947,N_3389);
nor U4038 (N_4038,N_3170,N_1145);
and U4039 (N_4039,N_519,N_2503);
nor U4040 (N_4040,N_1667,N_2841);
nor U4041 (N_4041,N_353,N_1502);
nor U4042 (N_4042,N_2105,N_3820);
and U4043 (N_4043,N_2496,N_158);
nor U4044 (N_4044,N_844,N_1181);
nor U4045 (N_4045,N_92,N_3514);
or U4046 (N_4046,N_2515,N_3798);
or U4047 (N_4047,N_656,N_2708);
or U4048 (N_4048,N_1102,N_3238);
and U4049 (N_4049,N_3206,N_2917);
nand U4050 (N_4050,N_3950,N_2764);
nand U4051 (N_4051,N_1817,N_213);
nand U4052 (N_4052,N_1119,N_3040);
nand U4053 (N_4053,N_769,N_2406);
and U4054 (N_4054,N_3508,N_2276);
nor U4055 (N_4055,N_2865,N_1050);
xnor U4056 (N_4056,N_531,N_1676);
and U4057 (N_4057,N_37,N_1549);
or U4058 (N_4058,N_376,N_1472);
xnor U4059 (N_4059,N_1248,N_1154);
nor U4060 (N_4060,N_3989,N_1614);
nor U4061 (N_4061,N_3405,N_252);
nand U4062 (N_4062,N_386,N_346);
nor U4063 (N_4063,N_2676,N_927);
or U4064 (N_4064,N_1469,N_2003);
nand U4065 (N_4065,N_1790,N_3833);
and U4066 (N_4066,N_1384,N_1173);
nand U4067 (N_4067,N_1881,N_2045);
nor U4068 (N_4068,N_895,N_1142);
nor U4069 (N_4069,N_3655,N_3417);
nand U4070 (N_4070,N_1243,N_3961);
nand U4071 (N_4071,N_815,N_3390);
nand U4072 (N_4072,N_2540,N_2692);
nand U4073 (N_4073,N_621,N_2620);
or U4074 (N_4074,N_2507,N_3914);
and U4075 (N_4075,N_3067,N_662);
nand U4076 (N_4076,N_1024,N_1986);
nor U4077 (N_4077,N_2939,N_3181);
nor U4078 (N_4078,N_2118,N_3231);
nor U4079 (N_4079,N_2579,N_1048);
nand U4080 (N_4080,N_3461,N_3036);
and U4081 (N_4081,N_2619,N_2982);
nand U4082 (N_4082,N_3358,N_2145);
and U4083 (N_4083,N_2638,N_1327);
and U4084 (N_4084,N_1786,N_2583);
and U4085 (N_4085,N_2106,N_1390);
nor U4086 (N_4086,N_2618,N_3623);
and U4087 (N_4087,N_587,N_2307);
xor U4088 (N_4088,N_192,N_2312);
nor U4089 (N_4089,N_2209,N_72);
nor U4090 (N_4090,N_2463,N_1075);
nand U4091 (N_4091,N_1435,N_2965);
nand U4092 (N_4092,N_2732,N_3816);
and U4093 (N_4093,N_3971,N_281);
or U4094 (N_4094,N_3537,N_2809);
and U4095 (N_4095,N_2851,N_2942);
and U4096 (N_4096,N_565,N_3769);
and U4097 (N_4097,N_969,N_2044);
nor U4098 (N_4098,N_2998,N_789);
or U4099 (N_4099,N_1076,N_2015);
nand U4100 (N_4100,N_216,N_3122);
nor U4101 (N_4101,N_742,N_2854);
or U4102 (N_4102,N_3504,N_84);
xnor U4103 (N_4103,N_1771,N_1876);
xor U4104 (N_4104,N_2701,N_140);
or U4105 (N_4105,N_3626,N_3538);
or U4106 (N_4106,N_1266,N_3199);
xnor U4107 (N_4107,N_294,N_3263);
nand U4108 (N_4108,N_1787,N_177);
or U4109 (N_4109,N_5,N_1002);
and U4110 (N_4110,N_1943,N_311);
nand U4111 (N_4111,N_3886,N_2240);
nand U4112 (N_4112,N_1211,N_2143);
nand U4113 (N_4113,N_713,N_3450);
nand U4114 (N_4114,N_1983,N_758);
and U4115 (N_4115,N_1360,N_3859);
or U4116 (N_4116,N_1847,N_3611);
nor U4117 (N_4117,N_1634,N_755);
nor U4118 (N_4118,N_3806,N_411);
or U4119 (N_4119,N_1853,N_2421);
and U4120 (N_4120,N_1740,N_1064);
or U4121 (N_4121,N_786,N_374);
and U4122 (N_4122,N_609,N_1172);
and U4123 (N_4123,N_2869,N_310);
nand U4124 (N_4124,N_2191,N_1030);
nand U4125 (N_4125,N_1926,N_3330);
nand U4126 (N_4126,N_467,N_726);
and U4127 (N_4127,N_2458,N_1246);
nand U4128 (N_4128,N_823,N_176);
and U4129 (N_4129,N_558,N_2800);
or U4130 (N_4130,N_3352,N_191);
or U4131 (N_4131,N_2804,N_2990);
nor U4132 (N_4132,N_2474,N_3804);
or U4133 (N_4133,N_3047,N_591);
and U4134 (N_4134,N_1987,N_472);
and U4135 (N_4135,N_3369,N_2975);
and U4136 (N_4136,N_1499,N_1020);
or U4137 (N_4137,N_2761,N_2399);
or U4138 (N_4138,N_3053,N_1284);
and U4139 (N_4139,N_3644,N_2637);
nor U4140 (N_4140,N_2491,N_2667);
and U4141 (N_4141,N_836,N_3282);
nor U4142 (N_4142,N_214,N_3789);
and U4143 (N_4143,N_1929,N_3709);
nor U4144 (N_4144,N_517,N_2280);
nor U4145 (N_4145,N_167,N_3215);
nand U4146 (N_4146,N_741,N_3915);
nor U4147 (N_4147,N_3883,N_2823);
nand U4148 (N_4148,N_2197,N_1099);
or U4149 (N_4149,N_3479,N_2325);
nor U4150 (N_4150,N_1796,N_2632);
nand U4151 (N_4151,N_3312,N_1091);
or U4152 (N_4152,N_2745,N_284);
and U4153 (N_4153,N_3147,N_3281);
or U4154 (N_4154,N_2393,N_141);
and U4155 (N_4155,N_246,N_1868);
and U4156 (N_4156,N_2996,N_2895);
and U4157 (N_4157,N_2392,N_876);
and U4158 (N_4158,N_2034,N_1255);
and U4159 (N_4159,N_3924,N_1925);
or U4160 (N_4160,N_2441,N_2612);
or U4161 (N_4161,N_2592,N_3808);
nand U4162 (N_4162,N_1705,N_401);
nand U4163 (N_4163,N_321,N_2987);
nand U4164 (N_4164,N_1296,N_2379);
or U4165 (N_4165,N_2156,N_1857);
nand U4166 (N_4166,N_1163,N_3790);
and U4167 (N_4167,N_2363,N_3518);
nand U4168 (N_4168,N_2545,N_2094);
and U4169 (N_4169,N_1316,N_611);
and U4170 (N_4170,N_724,N_3861);
or U4171 (N_4171,N_2232,N_87);
or U4172 (N_4172,N_2670,N_2086);
nor U4173 (N_4173,N_1712,N_1649);
nor U4174 (N_4174,N_199,N_2214);
and U4175 (N_4175,N_1395,N_1950);
nor U4176 (N_4176,N_1354,N_157);
and U4177 (N_4177,N_3388,N_3673);
and U4178 (N_4178,N_3427,N_2556);
or U4179 (N_4179,N_2346,N_627);
and U4180 (N_4180,N_226,N_1170);
and U4181 (N_4181,N_3933,N_2944);
and U4182 (N_4182,N_682,N_1486);
nand U4183 (N_4183,N_1222,N_3318);
and U4184 (N_4184,N_3822,N_548);
or U4185 (N_4185,N_3097,N_3640);
nor U4186 (N_4186,N_714,N_215);
or U4187 (N_4187,N_1961,N_2631);
and U4188 (N_4188,N_1368,N_447);
or U4189 (N_4189,N_2261,N_3243);
nor U4190 (N_4190,N_3250,N_2832);
nand U4191 (N_4191,N_750,N_1412);
or U4192 (N_4192,N_845,N_2260);
and U4193 (N_4193,N_1399,N_3973);
nor U4194 (N_4194,N_1948,N_2012);
or U4195 (N_4195,N_2582,N_283);
nor U4196 (N_4196,N_3013,N_3594);
and U4197 (N_4197,N_2215,N_2160);
and U4198 (N_4198,N_2054,N_2085);
nor U4199 (N_4199,N_1497,N_429);
or U4200 (N_4200,N_2932,N_291);
or U4201 (N_4201,N_2812,N_3339);
nand U4202 (N_4202,N_3912,N_59);
or U4203 (N_4203,N_392,N_985);
nor U4204 (N_4204,N_2903,N_520);
nor U4205 (N_4205,N_1468,N_3355);
nor U4206 (N_4206,N_3314,N_1358);
and U4207 (N_4207,N_2575,N_2977);
nand U4208 (N_4208,N_911,N_1232);
or U4209 (N_4209,N_608,N_3090);
nand U4210 (N_4210,N_2537,N_1436);
nand U4211 (N_4211,N_1561,N_389);
or U4212 (N_4212,N_3697,N_1205);
nand U4213 (N_4213,N_3313,N_388);
and U4214 (N_4214,N_2359,N_1032);
nand U4215 (N_4215,N_3847,N_3412);
nor U4216 (N_4216,N_1861,N_2166);
and U4217 (N_4217,N_2641,N_2614);
nor U4218 (N_4218,N_2084,N_1837);
or U4219 (N_4219,N_628,N_2347);
and U4220 (N_4220,N_3927,N_1540);
nand U4221 (N_4221,N_3023,N_1335);
nor U4222 (N_4222,N_450,N_1426);
or U4223 (N_4223,N_859,N_3459);
and U4224 (N_4224,N_2642,N_827);
nor U4225 (N_4225,N_2175,N_1450);
or U4226 (N_4226,N_3160,N_3345);
and U4227 (N_4227,N_858,N_534);
nand U4228 (N_4228,N_1956,N_1845);
and U4229 (N_4229,N_715,N_322);
nand U4230 (N_4230,N_495,N_3609);
nand U4231 (N_4231,N_1548,N_2465);
and U4232 (N_4232,N_2114,N_2457);
or U4233 (N_4233,N_699,N_1116);
xnor U4234 (N_4234,N_3509,N_3616);
nand U4235 (N_4235,N_3418,N_907);
or U4236 (N_4236,N_1150,N_794);
and U4237 (N_4237,N_173,N_1201);
nor U4238 (N_4238,N_1897,N_2373);
nand U4239 (N_4239,N_2025,N_422);
or U4240 (N_4240,N_1781,N_210);
nand U4241 (N_4241,N_1671,N_3571);
nand U4242 (N_4242,N_3303,N_555);
or U4243 (N_4243,N_3460,N_2731);
and U4244 (N_4244,N_542,N_335);
nor U4245 (N_4245,N_613,N_2512);
and U4246 (N_4246,N_3172,N_1813);
and U4247 (N_4247,N_3502,N_2032);
or U4248 (N_4248,N_733,N_865);
nand U4249 (N_4249,N_1285,N_2274);
and U4250 (N_4250,N_3109,N_2001);
nand U4251 (N_4251,N_1613,N_552);
nand U4252 (N_4252,N_3127,N_3424);
nor U4253 (N_4253,N_2570,N_1108);
nand U4254 (N_4254,N_3069,N_2394);
nand U4255 (N_4255,N_1337,N_2439);
xnor U4256 (N_4256,N_148,N_345);
nand U4257 (N_4257,N_498,N_2508);
or U4258 (N_4258,N_1098,N_1212);
or U4259 (N_4259,N_988,N_2607);
nor U4260 (N_4260,N_2466,N_1250);
or U4261 (N_4261,N_1543,N_2133);
nor U4262 (N_4262,N_2759,N_1953);
or U4263 (N_4263,N_2283,N_2908);
nand U4264 (N_4264,N_953,N_2679);
nor U4265 (N_4265,N_3123,N_2268);
nor U4266 (N_4266,N_2332,N_3286);
nor U4267 (N_4267,N_3041,N_2838);
or U4268 (N_4268,N_2391,N_2991);
nor U4269 (N_4269,N_2729,N_1514);
and U4270 (N_4270,N_1911,N_1605);
nor U4271 (N_4271,N_2088,N_1701);
and U4272 (N_4272,N_3399,N_3873);
or U4273 (N_4273,N_2342,N_3695);
and U4274 (N_4274,N_1001,N_69);
and U4275 (N_4275,N_333,N_1158);
nor U4276 (N_4276,N_3081,N_2891);
nor U4277 (N_4277,N_2901,N_3809);
nor U4278 (N_4278,N_839,N_1726);
nand U4279 (N_4279,N_759,N_1578);
nor U4280 (N_4280,N_1374,N_1785);
nand U4281 (N_4281,N_1833,N_1109);
and U4282 (N_4282,N_143,N_350);
or U4283 (N_4283,N_1094,N_2422);
and U4284 (N_4284,N_3050,N_2092);
nor U4285 (N_4285,N_3637,N_1446);
or U4286 (N_4286,N_1805,N_3319);
and U4287 (N_4287,N_810,N_723);
or U4288 (N_4288,N_830,N_3756);
and U4289 (N_4289,N_1488,N_359);
nor U4290 (N_4290,N_993,N_1177);
and U4291 (N_4291,N_3665,N_1905);
or U4292 (N_4292,N_501,N_1820);
nand U4293 (N_4293,N_1276,N_3393);
and U4294 (N_4294,N_2236,N_2714);
xnor U4295 (N_4295,N_7,N_1070);
and U4296 (N_4296,N_3641,N_3624);
and U4297 (N_4297,N_233,N_2884);
nor U4298 (N_4298,N_3784,N_972);
and U4299 (N_4299,N_2010,N_181);
nor U4300 (N_4300,N_28,N_3576);
and U4301 (N_4301,N_2665,N_2625);
nand U4302 (N_4302,N_249,N_1373);
or U4303 (N_4303,N_1668,N_2778);
nand U4304 (N_4304,N_3876,N_1542);
and U4305 (N_4305,N_289,N_115);
nor U4306 (N_4306,N_2213,N_1277);
or U4307 (N_4307,N_2622,N_1924);
nor U4308 (N_4308,N_1536,N_362);
and U4309 (N_4309,N_491,N_1229);
nor U4310 (N_4310,N_3370,N_3150);
and U4311 (N_4311,N_3797,N_2485);
or U4312 (N_4312,N_2773,N_3902);
xor U4313 (N_4313,N_207,N_3585);
or U4314 (N_4314,N_3516,N_2824);
nand U4315 (N_4315,N_1451,N_938);
and U4316 (N_4316,N_1982,N_847);
or U4317 (N_4317,N_2302,N_530);
nand U4318 (N_4318,N_336,N_3691);
nor U4319 (N_4319,N_400,N_636);
nand U4320 (N_4320,N_2447,N_2935);
or U4321 (N_4321,N_3503,N_300);
and U4322 (N_4322,N_966,N_3965);
nand U4323 (N_4323,N_888,N_722);
nand U4324 (N_4324,N_2289,N_2000);
nor U4325 (N_4325,N_3670,N_340);
or U4326 (N_4326,N_2652,N_2456);
nand U4327 (N_4327,N_3497,N_272);
or U4328 (N_4328,N_2877,N_2488);
and U4329 (N_4329,N_3982,N_3746);
and U4330 (N_4330,N_3828,N_3278);
or U4331 (N_4331,N_983,N_3378);
and U4332 (N_4332,N_202,N_2052);
nand U4333 (N_4333,N_1706,N_108);
nand U4334 (N_4334,N_3002,N_1015);
and U4335 (N_4335,N_1101,N_78);
nor U4336 (N_4336,N_385,N_549);
or U4337 (N_4337,N_3791,N_51);
nor U4338 (N_4338,N_1164,N_1361);
nor U4339 (N_4339,N_1573,N_3802);
or U4340 (N_4340,N_1046,N_1028);
nor U4341 (N_4341,N_546,N_3373);
nor U4342 (N_4342,N_1466,N_3224);
and U4343 (N_4343,N_3778,N_2089);
and U4344 (N_4344,N_624,N_1603);
or U4345 (N_4345,N_1657,N_169);
nand U4346 (N_4346,N_3510,N_2097);
or U4347 (N_4347,N_2962,N_1630);
or U4348 (N_4348,N_3544,N_3614);
nor U4349 (N_4349,N_3635,N_2041);
or U4350 (N_4350,N_2574,N_1455);
or U4351 (N_4351,N_1520,N_2573);
and U4352 (N_4352,N_439,N_2974);
or U4353 (N_4353,N_971,N_431);
and U4354 (N_4354,N_3327,N_194);
and U4355 (N_4355,N_171,N_3685);
and U4356 (N_4356,N_751,N_974);
and U4357 (N_4357,N_1690,N_2475);
and U4358 (N_4358,N_132,N_1544);
nand U4359 (N_4359,N_1505,N_27);
and U4360 (N_4360,N_81,N_1131);
or U4361 (N_4361,N_874,N_3546);
or U4362 (N_4362,N_1081,N_3027);
nand U4363 (N_4363,N_2292,N_2914);
and U4364 (N_4364,N_1580,N_2563);
or U4365 (N_4365,N_2953,N_965);
nor U4366 (N_4366,N_700,N_153);
and U4367 (N_4367,N_2370,N_672);
or U4368 (N_4368,N_3867,N_75);
nor U4369 (N_4369,N_835,N_2892);
and U4370 (N_4370,N_3668,N_1406);
or U4371 (N_4371,N_170,N_1538);
and U4372 (N_4372,N_2983,N_3719);
nand U4373 (N_4373,N_1144,N_1971);
nand U4374 (N_4374,N_3954,N_3863);
nand U4375 (N_4375,N_3938,N_36);
and U4376 (N_4376,N_3092,N_2022);
and U4377 (N_4377,N_277,N_1223);
or U4378 (N_4378,N_2769,N_3857);
or U4379 (N_4379,N_3870,N_2397);
and U4380 (N_4380,N_1749,N_649);
and U4381 (N_4381,N_2718,N_239);
or U4382 (N_4382,N_2385,N_2141);
nand U4383 (N_4383,N_106,N_1003);
and U4384 (N_4384,N_550,N_3005);
nor U4385 (N_4385,N_3483,N_3760);
nand U4386 (N_4386,N_3513,N_963);
nand U4387 (N_4387,N_2358,N_3070);
and U4388 (N_4388,N_1840,N_1954);
nor U4389 (N_4389,N_3855,N_1934);
or U4390 (N_4390,N_1969,N_3073);
and U4391 (N_4391,N_309,N_1097);
nor U4392 (N_4392,N_2921,N_514);
or U4393 (N_4393,N_2569,N_1898);
or U4394 (N_4394,N_973,N_1496);
xor U4395 (N_4395,N_2155,N_688);
or U4396 (N_4396,N_1106,N_1000);
and U4397 (N_4397,N_113,N_1661);
or U4398 (N_4398,N_2418,N_3446);
nor U4399 (N_4399,N_3022,N_2187);
and U4400 (N_4400,N_2472,N_1739);
nor U4401 (N_4401,N_2549,N_1587);
or U4402 (N_4402,N_1289,N_3521);
and U4403 (N_4403,N_222,N_1319);
nor U4404 (N_4404,N_2890,N_3977);
nand U4405 (N_4405,N_2915,N_3185);
or U4406 (N_4406,N_332,N_509);
nand U4407 (N_4407,N_2311,N_1936);
nor U4408 (N_4408,N_1365,N_2431);
or U4409 (N_4409,N_2937,N_2366);
nand U4410 (N_4410,N_2300,N_571);
nand U4411 (N_4411,N_1751,N_1441);
or U4412 (N_4412,N_3106,N_2314);
nor U4413 (N_4413,N_2539,N_2597);
nor U4414 (N_4414,N_2117,N_2427);
nand U4415 (N_4415,N_1914,N_161);
and U4416 (N_4416,N_1460,N_260);
or U4417 (N_4417,N_744,N_2423);
and U4418 (N_4418,N_3400,N_1732);
xor U4419 (N_4419,N_2425,N_1184);
nand U4420 (N_4420,N_3118,N_391);
nand U4421 (N_4421,N_2684,N_1856);
nor U4422 (N_4422,N_2171,N_1968);
nor U4423 (N_4423,N_1299,N_45);
nand U4424 (N_4424,N_1060,N_1362);
or U4425 (N_4425,N_2779,N_1976);
xnor U4426 (N_4426,N_760,N_2478);
nand U4427 (N_4427,N_1409,N_484);
nor U4428 (N_4428,N_1039,N_853);
or U4429 (N_4429,N_370,N_2231);
nor U4430 (N_4430,N_3703,N_2560);
and U4431 (N_4431,N_3734,N_2789);
nand U4432 (N_4432,N_99,N_990);
or U4433 (N_4433,N_2700,N_2390);
and U4434 (N_4434,N_2857,N_808);
or U4435 (N_4435,N_761,N_2698);
or U4436 (N_4436,N_100,N_1874);
or U4437 (N_4437,N_3885,N_1909);
nand U4438 (N_4438,N_3395,N_3204);
or U4439 (N_4439,N_469,N_1579);
nor U4440 (N_4440,N_2100,N_3737);
nand U4441 (N_4441,N_1673,N_803);
or U4442 (N_4442,N_2295,N_2303);
or U4443 (N_4443,N_1599,N_2081);
or U4444 (N_4444,N_3362,N_2202);
or U4445 (N_4445,N_2972,N_3311);
xnor U4446 (N_4446,N_3553,N_1104);
and U4447 (N_4447,N_299,N_1883);
nor U4448 (N_4448,N_298,N_364);
nor U4449 (N_4449,N_3711,N_2664);
or U4450 (N_4450,N_1919,N_468);
nand U4451 (N_4451,N_2695,N_1746);
xnor U4452 (N_4452,N_1597,N_3203);
nand U4453 (N_4453,N_220,N_2879);
and U4454 (N_4454,N_1918,N_164);
or U4455 (N_4455,N_1566,N_2310);
nand U4456 (N_4456,N_18,N_579);
nor U4457 (N_4457,N_1999,N_2495);
or U4458 (N_4458,N_3452,N_3377);
nand U4459 (N_4459,N_1584,N_1652);
or U4460 (N_4460,N_269,N_1005);
and U4461 (N_4461,N_2492,N_114);
and U4462 (N_4462,N_1941,N_149);
nand U4463 (N_4463,N_1294,N_1917);
nor U4464 (N_4464,N_2756,N_2238);
nor U4465 (N_4465,N_3615,N_897);
or U4466 (N_4466,N_1779,N_1816);
nor U4467 (N_4467,N_3182,N_2705);
nor U4468 (N_4468,N_105,N_2257);
nor U4469 (N_4469,N_1031,N_708);
nand U4470 (N_4470,N_127,N_3580);
or U4471 (N_4471,N_1939,N_2180);
and U4472 (N_4472,N_956,N_461);
nand U4473 (N_4473,N_3943,N_1998);
nand U4474 (N_4474,N_1858,N_2926);
or U4475 (N_4475,N_1831,N_2079);
or U4476 (N_4476,N_2790,N_3687);
and U4477 (N_4477,N_3466,N_3721);
or U4478 (N_4478,N_3743,N_620);
and U4479 (N_4479,N_1312,N_449);
or U4480 (N_4480,N_1423,N_2324);
nor U4481 (N_4481,N_3884,N_1829);
nand U4482 (N_4482,N_976,N_1565);
or U4483 (N_4483,N_3819,N_3402);
or U4484 (N_4484,N_1162,N_251);
nand U4485 (N_4485,N_707,N_1722);
or U4486 (N_4486,N_2339,N_748);
nor U4487 (N_4487,N_2852,N_2699);
nor U4488 (N_4488,N_2997,N_1723);
or U4489 (N_4489,N_2429,N_3841);
nand U4490 (N_4490,N_465,N_1662);
nand U4491 (N_4491,N_1892,N_2934);
nand U4492 (N_4492,N_3492,N_3679);
and U4493 (N_4493,N_3138,N_3666);
or U4494 (N_4494,N_3184,N_2609);
nor U4495 (N_4495,N_650,N_3477);
and U4496 (N_4496,N_3941,N_1363);
or U4497 (N_4497,N_308,N_2357);
nor U4498 (N_4498,N_1347,N_1459);
and U4499 (N_4499,N_1916,N_2361);
or U4500 (N_4500,N_1259,N_1241);
nand U4501 (N_4501,N_1612,N_702);
nand U4502 (N_4502,N_580,N_1860);
nand U4503 (N_4503,N_3284,N_1679);
and U4504 (N_4504,N_635,N_3012);
nand U4505 (N_4505,N_399,N_3948);
nor U4506 (N_4506,N_2109,N_1962);
xnor U4507 (N_4507,N_1080,N_2072);
or U4508 (N_4508,N_1607,N_1058);
nor U4509 (N_4509,N_80,N_1063);
and U4510 (N_4510,N_1841,N_1424);
or U4511 (N_4511,N_518,N_2577);
and U4512 (N_4512,N_2711,N_3920);
or U4513 (N_4513,N_1823,N_1655);
nand U4514 (N_4514,N_920,N_3636);
nor U4515 (N_4515,N_3632,N_2152);
nand U4516 (N_4516,N_2053,N_667);
nor U4517 (N_4517,N_3304,N_670);
nor U4518 (N_4518,N_3102,N_2564);
nor U4519 (N_4519,N_2968,N_313);
nor U4520 (N_4520,N_57,N_1410);
nand U4521 (N_4521,N_2875,N_1237);
nand U4522 (N_4522,N_379,N_1736);
nor U4523 (N_4523,N_3096,N_2706);
nand U4524 (N_4524,N_2494,N_3917);
nor U4525 (N_4525,N_1372,N_899);
nand U4526 (N_4526,N_594,N_848);
nor U4527 (N_4527,N_851,N_2120);
or U4528 (N_4528,N_3613,N_1700);
nand U4529 (N_4529,N_2107,N_201);
and U4530 (N_4530,N_3763,N_1513);
and U4531 (N_4531,N_3931,N_2476);
nand U4532 (N_4532,N_2020,N_2103);
nand U4533 (N_4533,N_2636,N_3328);
nor U4534 (N_4534,N_3741,N_1526);
and U4535 (N_4535,N_243,N_445);
nand U4536 (N_4536,N_997,N_3500);
and U4537 (N_4537,N_1345,N_478);
and U4538 (N_4538,N_22,N_2629);
nand U4539 (N_4539,N_902,N_1735);
nor U4540 (N_4540,N_3045,N_2330);
nand U4541 (N_4541,N_2896,N_2727);
and U4542 (N_4542,N_1991,N_2412);
and U4543 (N_4543,N_3485,N_3151);
and U4544 (N_4544,N_819,N_1651);
nand U4545 (N_4545,N_599,N_3869);
nand U4546 (N_4546,N_1313,N_486);
and U4547 (N_4547,N_2002,N_2653);
nand U4548 (N_4548,N_1778,N_3126);
and U4549 (N_4549,N_2814,N_2046);
and U4550 (N_4550,N_2493,N_2519);
nor U4551 (N_4551,N_2828,N_434);
and U4552 (N_4552,N_3753,N_3331);
or U4553 (N_4553,N_230,N_3878);
and U4554 (N_4554,N_991,N_1351);
or U4555 (N_4555,N_360,N_104);
and U4556 (N_4556,N_1773,N_193);
nor U4557 (N_4557,N_1966,N_3764);
or U4558 (N_4558,N_3678,N_903);
and U4559 (N_4559,N_305,N_1586);
and U4560 (N_4560,N_1215,N_183);
nor U4561 (N_4561,N_1346,N_3921);
and U4562 (N_4562,N_1886,N_3785);
and U4563 (N_4563,N_982,N_3153);
or U4564 (N_4564,N_1733,N_1308);
or U4565 (N_4565,N_3063,N_3829);
or U4566 (N_4566,N_3071,N_2479);
nand U4567 (N_4567,N_814,N_2608);
nor U4568 (N_4568,N_3925,N_2254);
and U4569 (N_4569,N_453,N_1204);
nor U4570 (N_4570,N_1096,N_2252);
and U4571 (N_4571,N_1067,N_2659);
nand U4572 (N_4572,N_483,N_1849);
or U4573 (N_4573,N_2846,N_2075);
nand U4574 (N_4574,N_200,N_2955);
or U4575 (N_4575,N_3849,N_3531);
nand U4576 (N_4576,N_919,N_3030);
or U4577 (N_4577,N_2149,N_1465);
and U4578 (N_4578,N_1342,N_2192);
nand U4579 (N_4579,N_0,N_655);
or U4580 (N_4580,N_1413,N_3391);
and U4581 (N_4581,N_24,N_1198);
or U4582 (N_4582,N_3332,N_3083);
and U4583 (N_4583,N_3396,N_3413);
nor U4584 (N_4584,N_2199,N_1492);
and U4585 (N_4585,N_2989,N_1642);
and U4586 (N_4586,N_616,N_20);
nor U4587 (N_4587,N_3228,N_435);
nand U4588 (N_4588,N_3653,N_1509);
nor U4589 (N_4589,N_3928,N_3280);
xnor U4590 (N_4590,N_879,N_2565);
or U4591 (N_4591,N_999,N_1103);
and U4592 (N_4592,N_3720,N_2402);
and U4593 (N_4593,N_433,N_1758);
and U4594 (N_4594,N_1155,N_2432);
nand U4595 (N_4595,N_1325,N_159);
or U4596 (N_4596,N_49,N_1100);
nor U4597 (N_4597,N_1694,N_756);
nand U4598 (N_4598,N_3568,N_3684);
nor U4599 (N_4599,N_2285,N_1891);
or U4600 (N_4600,N_968,N_3253);
nand U4601 (N_4601,N_3028,N_1873);
nor U4602 (N_4602,N_2749,N_1234);
nand U4603 (N_4603,N_2396,N_3359);
nor U4604 (N_4604,N_3864,N_889);
nand U4605 (N_4605,N_1295,N_1774);
or U4606 (N_4606,N_2306,N_3487);
and U4607 (N_4607,N_622,N_2703);
and U4608 (N_4608,N_2923,N_1394);
nor U4609 (N_4609,N_2567,N_3796);
nor U4610 (N_4610,N_893,N_451);
nand U4611 (N_4611,N_1656,N_932);
nand U4612 (N_4612,N_3046,N_2216);
or U4613 (N_4613,N_2558,N_3813);
and U4614 (N_4614,N_1795,N_2999);
or U4615 (N_4615,N_2076,N_2126);
nor U4616 (N_4616,N_3562,N_2532);
nor U4617 (N_4617,N_2516,N_1583);
nor U4618 (N_4618,N_3482,N_3175);
and U4619 (N_4619,N_266,N_94);
nor U4620 (N_4620,N_2723,N_665);
and U4621 (N_4621,N_1625,N_1559);
and U4622 (N_4622,N_516,N_454);
nor U4623 (N_4623,N_3946,N_2606);
or U4624 (N_4624,N_1767,N_3979);
and U4625 (N_4625,N_3718,N_3269);
or U4626 (N_4626,N_2042,N_2945);
nor U4627 (N_4627,N_2461,N_754);
nor U4628 (N_4628,N_2801,N_2027);
and U4629 (N_4629,N_675,N_256);
and U4630 (N_4630,N_1129,N_3077);
nor U4631 (N_4631,N_1852,N_145);
or U4632 (N_4632,N_1594,N_208);
or U4633 (N_4633,N_1660,N_3052);
or U4634 (N_4634,N_2985,N_1920);
and U4635 (N_4635,N_3659,N_1721);
nor U4636 (N_4636,N_1955,N_3932);
nand U4637 (N_4637,N_3549,N_26);
or U4638 (N_4638,N_85,N_1022);
nor U4639 (N_4639,N_1398,N_1978);
or U4640 (N_4640,N_1882,N_809);
nor U4641 (N_4641,N_780,N_3208);
nor U4642 (N_4642,N_1665,N_3608);
nor U4643 (N_4643,N_1072,N_3094);
and U4644 (N_4644,N_3366,N_2660);
nor U4645 (N_4645,N_96,N_3672);
nor U4646 (N_4646,N_2951,N_921);
and U4647 (N_4647,N_838,N_1404);
nor U4648 (N_4648,N_1609,N_2204);
or U4649 (N_4649,N_438,N_111);
and U4650 (N_4650,N_1750,N_1290);
nor U4651 (N_4651,N_234,N_152);
nor U4652 (N_4652,N_3134,N_1608);
or U4653 (N_4653,N_2320,N_1938);
and U4654 (N_4654,N_1843,N_791);
nand U4655 (N_4655,N_1684,N_2211);
and U4656 (N_4656,N_1391,N_492);
nand U4657 (N_4657,N_2777,N_1960);
nor U4658 (N_4658,N_2112,N_1945);
nor U4659 (N_4659,N_68,N_2058);
and U4660 (N_4660,N_885,N_1629);
nor U4661 (N_4661,N_1762,N_1904);
nand U4662 (N_4662,N_1017,N_1377);
nor U4663 (N_4663,N_3519,N_3229);
and U4664 (N_4664,N_992,N_1697);
and U4665 (N_4665,N_3104,N_3507);
or U4666 (N_4666,N_2671,N_3962);
or U4667 (N_4667,N_1054,N_3363);
or U4668 (N_4668,N_2028,N_3474);
nor U4669 (N_4669,N_2771,N_2061);
xor U4670 (N_4670,N_3146,N_3599);
nor U4671 (N_4671,N_934,N_3267);
nand U4672 (N_4672,N_373,N_2500);
and U4673 (N_4673,N_926,N_1552);
and U4674 (N_4674,N_1194,N_275);
nand U4675 (N_4675,N_2460,N_1025);
nor U4676 (N_4676,N_1648,N_2818);
or U4677 (N_4677,N_344,N_2369);
nand U4678 (N_4678,N_3029,N_3079);
and U4679 (N_4679,N_1126,N_186);
and U4680 (N_4680,N_717,N_3290);
and U4681 (N_4681,N_731,N_2870);
xnor U4682 (N_4682,N_2994,N_1228);
or U4683 (N_4683,N_2016,N_653);
and U4684 (N_4684,N_2628,N_2430);
or U4685 (N_4685,N_1680,N_866);
and U4686 (N_4686,N_2350,N_1071);
nand U4687 (N_4687,N_2543,N_618);
nor U4688 (N_4688,N_1146,N_1678);
and U4689 (N_4689,N_2848,N_678);
or U4690 (N_4690,N_1167,N_1291);
nor U4691 (N_4691,N_1429,N_262);
or U4692 (N_4692,N_1233,N_3055);
or U4693 (N_4693,N_1970,N_1719);
or U4694 (N_4694,N_3425,N_139);
xnor U4695 (N_4695,N_2101,N_3677);
nand U4696 (N_4696,N_1636,N_1417);
or U4697 (N_4697,N_1944,N_2147);
or U4698 (N_4698,N_728,N_2134);
and U4699 (N_4699,N_1851,N_121);
nor U4700 (N_4700,N_3565,N_1425);
nand U4701 (N_4701,N_3439,N_2263);
nand U4702 (N_4702,N_2341,N_3227);
and U4703 (N_4703,N_1688,N_418);
and U4704 (N_4704,N_270,N_527);
nor U4705 (N_4705,N_76,N_2063);
or U4706 (N_4706,N_1988,N_2343);
nor U4707 (N_4707,N_65,N_1725);
and U4708 (N_4708,N_1434,N_1231);
nand U4709 (N_4709,N_1972,N_3866);
or U4710 (N_4710,N_779,N_3992);
or U4711 (N_4711,N_1367,N_3660);
nand U4712 (N_4712,N_3713,N_2602);
nand U4713 (N_4713,N_1822,N_2517);
or U4714 (N_4714,N_3019,N_2651);
nand U4715 (N_4715,N_2668,N_3794);
and U4716 (N_4716,N_43,N_1870);
nor U4717 (N_4717,N_2444,N_1832);
and U4718 (N_4718,N_629,N_1045);
or U4719 (N_4719,N_109,N_2521);
or U4720 (N_4720,N_2596,N_832);
and U4721 (N_4721,N_1534,N_1900);
or U4722 (N_4722,N_592,N_3072);
or U4723 (N_4723,N_2530,N_3716);
and U4724 (N_4724,N_3105,N_771);
nor U4725 (N_4725,N_3468,N_2525);
and U4726 (N_4726,N_2704,N_567);
nor U4727 (N_4727,N_1899,N_40);
or U4728 (N_4728,N_767,N_1355);
nand U4729 (N_4729,N_512,N_150);
nand U4730 (N_4730,N_408,N_3360);
nand U4731 (N_4731,N_1623,N_2821);
or U4732 (N_4732,N_1677,N_21);
nor U4733 (N_4733,N_1507,N_3738);
and U4734 (N_4734,N_358,N_526);
nand U4735 (N_4735,N_198,N_2864);
nand U4736 (N_4736,N_1692,N_3952);
nor U4737 (N_4737,N_2572,N_3475);
or U4738 (N_4738,N_1086,N_380);
and U4739 (N_4739,N_423,N_2388);
and U4740 (N_4740,N_1095,N_540);
or U4741 (N_4741,N_508,N_288);
or U4742 (N_4742,N_642,N_2702);
or U4743 (N_4743,N_2691,N_1035);
nor U4744 (N_4744,N_3783,N_2398);
nand U4745 (N_4745,N_3087,N_2205);
and U4746 (N_4746,N_1029,N_2064);
nor U4747 (N_4747,N_2630,N_1038);
nor U4748 (N_4748,N_673,N_3021);
and U4749 (N_4749,N_2163,N_3066);
nor U4750 (N_4750,N_1523,N_2265);
nor U4751 (N_4751,N_1282,N_282);
nand U4752 (N_4752,N_1165,N_1310);
or U4753 (N_4753,N_2798,N_2847);
xor U4754 (N_4754,N_2963,N_694);
or U4755 (N_4755,N_1947,N_485);
nor U4756 (N_4756,N_3471,N_3244);
and U4757 (N_4757,N_852,N_265);
nand U4758 (N_4758,N_746,N_236);
nor U4759 (N_4759,N_3586,N_2979);
or U4760 (N_4760,N_2743,N_180);
nand U4761 (N_4761,N_574,N_52);
nor U4762 (N_4762,N_2219,N_3772);
nand U4763 (N_4763,N_1023,N_280);
or U4764 (N_4764,N_833,N_1087);
nor U4765 (N_4765,N_807,N_3411);
nor U4766 (N_4766,N_1850,N_2661);
or U4767 (N_4767,N_2278,N_1449);
and U4768 (N_4768,N_3939,N_770);
nor U4769 (N_4769,N_1263,N_2551);
and U4770 (N_4770,N_3985,N_497);
and U4771 (N_4771,N_3279,N_1592);
and U4772 (N_4772,N_395,N_800);
or U4773 (N_4773,N_2542,N_2326);
or U4774 (N_4774,N_3817,N_1550);
or U4775 (N_4775,N_1835,N_2470);
or U4776 (N_4776,N_3414,N_1021);
nand U4777 (N_4777,N_3913,N_1824);
nor U4778 (N_4778,N_10,N_2142);
or U4779 (N_4779,N_2835,N_1068);
nor U4780 (N_4780,N_950,N_425);
or U4781 (N_4781,N_3899,N_3634);
and U4782 (N_4782,N_3664,N_9);
or U4783 (N_4783,N_142,N_2234);
or U4784 (N_4784,N_3498,N_2739);
nand U4785 (N_4785,N_3431,N_2267);
and U4786 (N_4786,N_253,N_1989);
and U4787 (N_4787,N_3744,N_2897);
nand U4788 (N_4788,N_3202,N_1323);
nor U4789 (N_4789,N_2408,N_762);
nor U4790 (N_4790,N_1105,N_205);
nand U4791 (N_4791,N_3223,N_2646);
or U4792 (N_4792,N_1757,N_1946);
nand U4793 (N_4793,N_3152,N_351);
and U4794 (N_4794,N_2794,N_745);
nand U4795 (N_4795,N_1278,N_2448);
nand U4796 (N_4796,N_3076,N_1214);
and U4797 (N_4797,N_2039,N_884);
or U4798 (N_4798,N_2687,N_957);
nor U4799 (N_4799,N_1458,N_146);
or U4800 (N_4800,N_2091,N_816);
nand U4801 (N_4801,N_2533,N_237);
or U4802 (N_4802,N_2277,N_79);
nor U4803 (N_4803,N_129,N_3384);
or U4804 (N_4804,N_1653,N_2894);
or U4805 (N_4805,N_1604,N_864);
nand U4806 (N_4806,N_1033,N_2634);
and U4807 (N_4807,N_2297,N_2906);
and U4808 (N_4808,N_680,N_2272);
nor U4809 (N_4809,N_1261,N_3117);
nor U4810 (N_4810,N_1693,N_1776);
nand U4811 (N_4811,N_357,N_2836);
nand U4812 (N_4812,N_695,N_511);
or U4813 (N_4813,N_302,N_3383);
or U4814 (N_4814,N_3511,N_3780);
nor U4815 (N_4815,N_2050,N_3774);
nor U4816 (N_4816,N_3573,N_647);
nand U4817 (N_4817,N_1089,N_1810);
or U4818 (N_4818,N_2309,N_2450);
nor U4819 (N_4819,N_3524,N_3998);
nor U4820 (N_4820,N_1300,N_38);
nand U4821 (N_4821,N_162,N_1437);
and U4822 (N_4822,N_933,N_2013);
and U4823 (N_4823,N_1937,N_3893);
nand U4824 (N_4824,N_812,N_1515);
nor U4825 (N_4825,N_1432,N_849);
and U4826 (N_4826,N_3526,N_2662);
nor U4827 (N_4827,N_598,N_772);
and U4828 (N_4828,N_892,N_432);
nand U4829 (N_4829,N_904,N_2898);
and U4830 (N_4830,N_1480,N_3239);
or U4831 (N_4831,N_3457,N_1311);
nand U4832 (N_4832,N_940,N_407);
nand U4833 (N_4833,N_184,N_3881);
nand U4834 (N_4834,N_2669,N_2354);
and U4835 (N_4835,N_2561,N_1143);
nand U4836 (N_4836,N_923,N_3909);
or U4837 (N_4837,N_48,N_2228);
or U4838 (N_4838,N_3739,N_1491);
nor U4839 (N_4839,N_3532,N_3401);
or U4840 (N_4840,N_1483,N_3501);
and U4841 (N_4841,N_908,N_533);
and U4842 (N_4842,N_2635,N_584);
nor U4843 (N_4843,N_3522,N_1895);
or U4844 (N_4844,N_2958,N_3701);
nand U4845 (N_4845,N_3722,N_3922);
or U4846 (N_4846,N_1593,N_2925);
or U4847 (N_4847,N_2007,N_2206);
or U4848 (N_4848,N_3639,N_2110);
or U4849 (N_4849,N_637,N_1545);
and U4850 (N_4850,N_3110,N_29);
nand U4851 (N_4851,N_3473,N_165);
nand U4852 (N_4852,N_2176,N_3645);
nand U4853 (N_4853,N_3065,N_1793);
and U4854 (N_4854,N_417,N_834);
nor U4855 (N_4855,N_3845,N_1503);
nor U4856 (N_4856,N_2433,N_2445);
nor U4857 (N_4857,N_2190,N_3618);
nor U4858 (N_4858,N_2335,N_507);
and U4859 (N_4859,N_2621,N_905);
or U4860 (N_4860,N_818,N_765);
nand U4861 (N_4861,N_3101,N_3505);
and U4862 (N_4862,N_2218,N_593);
and U4863 (N_4863,N_244,N_1744);
or U4864 (N_4864,N_545,N_1884);
nor U4865 (N_4865,N_1160,N_1197);
and U4866 (N_4866,N_3983,N_1606);
nand U4867 (N_4867,N_2511,N_2387);
xnor U4868 (N_4868,N_218,N_2266);
and U4869 (N_4869,N_2568,N_1888);
and U4870 (N_4870,N_1415,N_3009);
and U4871 (N_4871,N_47,N_133);
nand U4872 (N_4872,N_692,N_3578);
nand U4873 (N_4873,N_3095,N_134);
and U4874 (N_4874,N_2115,N_1379);
or U4875 (N_4875,N_2986,N_2355);
and U4876 (N_4876,N_138,N_1218);
or U4877 (N_4877,N_3323,N_2807);
or U4878 (N_4878,N_2681,N_2462);
nor U4879 (N_4879,N_3310,N_2023);
or U4880 (N_4880,N_3308,N_2694);
and U4881 (N_4881,N_704,N_1647);
and U4882 (N_4882,N_588,N_2164);
and U4883 (N_4883,N_306,N_2677);
or U4884 (N_4884,N_2073,N_3478);
nand U4885 (N_4885,N_1763,N_3082);
or U4886 (N_4886,N_2799,N_2374);
nor U4887 (N_4887,N_3340,N_2255);
nand U4888 (N_4888,N_2647,N_2148);
nand U4889 (N_4889,N_1709,N_2212);
nor U4890 (N_4890,N_3298,N_2442);
or U4891 (N_4891,N_1431,N_1059);
and U4892 (N_4892,N_2874,N_2725);
nor U4893 (N_4893,N_3945,N_2327);
and U4894 (N_4894,N_906,N_1397);
or U4895 (N_4895,N_1169,N_1788);
nand U4896 (N_4896,N_3037,N_2316);
or U4897 (N_4897,N_2239,N_3682);
or U4898 (N_4898,N_3062,N_981);
nor U4899 (N_4899,N_1624,N_479);
or U4900 (N_4900,N_3814,N_1893);
xnor U4901 (N_4901,N_3249,N_2282);
nand U4902 (N_4902,N_659,N_837);
nor U4903 (N_4903,N_2576,N_3892);
nor U4904 (N_4904,N_3630,N_1008);
nor U4905 (N_4905,N_3189,N_3357);
nor U4906 (N_4906,N_2286,N_326);
and U4907 (N_4907,N_603,N_3119);
nand U4908 (N_4908,N_2113,N_3588);
nand U4909 (N_4909,N_3661,N_440);
nand U4910 (N_4910,N_3493,N_1010);
nor U4911 (N_4911,N_500,N_1332);
and U4912 (N_4912,N_3157,N_1846);
and U4913 (N_4913,N_3300,N_523);
and U4914 (N_4914,N_3906,N_3725);
or U4915 (N_4915,N_2640,N_1137);
or U4916 (N_4916,N_2831,N_55);
nor U4917 (N_4917,N_3559,N_2839);
nor U4918 (N_4918,N_3221,N_3900);
nor U4919 (N_4919,N_1479,N_3128);
nor U4920 (N_4920,N_3730,N_2438);
nor U4921 (N_4921,N_1935,N_1180);
nand U4922 (N_4922,N_352,N_931);
or U4923 (N_4923,N_3201,N_2353);
nand U4924 (N_4924,N_178,N_1092);
nand U4925 (N_4925,N_2615,N_2258);
and U4926 (N_4926,N_414,N_1053);
and U4927 (N_4927,N_3995,N_2970);
and U4928 (N_4928,N_3496,N_1734);
or U4929 (N_4929,N_2179,N_1159);
nor U4930 (N_4930,N_1866,N_1040);
or U4931 (N_4931,N_910,N_1619);
or U4932 (N_4932,N_2786,N_3850);
nor U4933 (N_4933,N_1125,N_984);
or U4934 (N_4934,N_1047,N_1438);
and U4935 (N_4935,N_2554,N_3085);
nand U4936 (N_4936,N_3748,N_456);
and U4937 (N_4937,N_490,N_734);
nand U4938 (N_4938,N_797,N_2473);
nand U4939 (N_4939,N_2882,N_3837);
nand U4940 (N_4940,N_1803,N_1283);
nor U4941 (N_4941,N_2150,N_3043);
and U4942 (N_4942,N_363,N_3560);
nand U4943 (N_4943,N_466,N_3057);
and U4944 (N_4944,N_3163,N_2389);
or U4945 (N_4945,N_2813,N_1784);
nor U4946 (N_4946,N_873,N_2787);
and U4947 (N_4947,N_2144,N_1389);
nand U4948 (N_4948,N_559,N_1301);
nor U4949 (N_4949,N_1286,N_3969);
nor U4950 (N_4950,N_1013,N_1344);
nand U4951 (N_4951,N_3839,N_2376);
nand U4952 (N_4952,N_1079,N_962);
and U4953 (N_4953,N_795,N_405);
nand U4954 (N_4954,N_97,N_3051);
nor U4955 (N_4955,N_1419,N_3168);
or U4956 (N_4956,N_2591,N_1601);
nor U4957 (N_4957,N_1577,N_3444);
or U4958 (N_4958,N_1508,N_174);
or U4959 (N_4959,N_3844,N_994);
and U4960 (N_4960,N_2967,N_2531);
or U4961 (N_4961,N_1830,N_2153);
and U4962 (N_4962,N_914,N_1539);
nand U4963 (N_4963,N_2395,N_3326);
and U4964 (N_4964,N_1085,N_1244);
or U4965 (N_4965,N_2059,N_1187);
or U4966 (N_4966,N_1242,N_98);
or U4967 (N_4967,N_1620,N_325);
nand U4968 (N_4968,N_3633,N_116);
nand U4969 (N_4969,N_3727,N_1383);
nand U4970 (N_4970,N_3074,N_1270);
nand U4971 (N_4971,N_3197,N_70);
or U4972 (N_4972,N_1118,N_3757);
and U4973 (N_4973,N_625,N_3824);
nand U4974 (N_4974,N_2087,N_1885);
or U4975 (N_4975,N_2842,N_2247);
nand U4976 (N_4976,N_2933,N_101);
or U4977 (N_4977,N_3631,N_2026);
or U4978 (N_4978,N_3723,N_3972);
and U4979 (N_4979,N_2182,N_881);
nor U4980 (N_4980,N_2480,N_2534);
nor U4981 (N_4981,N_2753,N_2313);
or U4982 (N_4982,N_3830,N_3120);
or U4983 (N_4983,N_850,N_91);
or U4984 (N_4984,N_2557,N_711);
and U4985 (N_4985,N_1764,N_887);
nand U4986 (N_4986,N_3115,N_195);
or U4987 (N_4987,N_581,N_3652);
nand U4988 (N_4988,N_2524,N_3704);
nand U4989 (N_4989,N_1275,N_307);
or U4990 (N_4990,N_1307,N_1463);
nor U4991 (N_4991,N_3860,N_3663);
nand U4992 (N_4992,N_1770,N_2011);
and U4993 (N_4993,N_2482,N_1836);
nor U4994 (N_4994,N_970,N_3167);
or U4995 (N_4995,N_154,N_1531);
or U4996 (N_4996,N_2269,N_231);
nor U4997 (N_4997,N_2036,N_883);
or U4998 (N_4998,N_696,N_1495);
or U4999 (N_4999,N_387,N_3815);
and U5000 (N_5000,N_3394,N_560);
and U5001 (N_5001,N_151,N_2331);
and U5002 (N_5002,N_811,N_330);
nand U5003 (N_5003,N_3582,N_1348);
and U5004 (N_5004,N_2796,N_3408);
and U5005 (N_5005,N_2693,N_1871);
nor U5006 (N_5006,N_1718,N_658);
and U5007 (N_5007,N_63,N_1975);
nor U5008 (N_5008,N_2290,N_261);
nor U5009 (N_5009,N_928,N_3793);
and U5010 (N_5010,N_2949,N_107);
or U5011 (N_5011,N_554,N_2858);
nand U5012 (N_5012,N_2735,N_3397);
or U5013 (N_5013,N_1317,N_1615);
nand U5014 (N_5014,N_2961,N_462);
nor U5015 (N_5015,N_2116,N_3690);
and U5016 (N_5016,N_3786,N_1052);
and U5017 (N_5017,N_2950,N_2344);
or U5018 (N_5018,N_2673,N_2177);
nor U5019 (N_5019,N_3597,N_296);
and U5020 (N_5020,N_996,N_2710);
nor U5021 (N_5021,N_2603,N_1933);
xor U5022 (N_5022,N_367,N_738);
or U5023 (N_5023,N_3141,N_1589);
or U5024 (N_5024,N_1168,N_420);
or U5025 (N_5025,N_3598,N_784);
and U5026 (N_5026,N_2872,N_19);
nor U5027 (N_5027,N_842,N_2047);
nor U5028 (N_5028,N_1430,N_443);
and U5029 (N_5029,N_1980,N_2562);
or U5030 (N_5030,N_2803,N_3656);
and U5031 (N_5031,N_943,N_1875);
xor U5032 (N_5032,N_1408,N_2030);
nand U5033 (N_5033,N_1268,N_2146);
nand U5034 (N_5034,N_1553,N_476);
nand U5035 (N_5035,N_2688,N_1121);
nand U5036 (N_5036,N_327,N_1675);
and U5037 (N_5037,N_3018,N_3604);
nor U5038 (N_5038,N_1407,N_3307);
nand U5039 (N_5039,N_2960,N_444);
nand U5040 (N_5040,N_3348,N_1111);
nand U5041 (N_5041,N_2850,N_1556);
or U5042 (N_5042,N_2588,N_1161);
nor U5043 (N_5043,N_3173,N_1382);
or U5044 (N_5044,N_287,N_1942);
or U5045 (N_5045,N_1590,N_1756);
or U5046 (N_5046,N_3752,N_187);
or U5047 (N_5047,N_355,N_1801);
nand U5048 (N_5048,N_2683,N_2323);
or U5049 (N_5049,N_56,N_2371);
nor U5050 (N_5050,N_219,N_1153);
nor U5051 (N_5051,N_3874,N_2899);
and U5052 (N_5052,N_64,N_3392);
nand U5053 (N_5053,N_1304,N_2716);
nor U5054 (N_5054,N_1207,N_3981);
or U5055 (N_5055,N_1761,N_1055);
or U5056 (N_5056,N_1132,N_348);
and U5057 (N_5057,N_50,N_3986);
and U5058 (N_5058,N_1405,N_1959);
or U5059 (N_5059,N_730,N_2776);
nor U5060 (N_5060,N_2139,N_3792);
and U5061 (N_5061,N_2645,N_3587);
nand U5062 (N_5062,N_1807,N_1202);
or U5063 (N_5063,N_424,N_2367);
nor U5064 (N_5064,N_841,N_3462);
or U5065 (N_5065,N_2377,N_3364);
nand U5066 (N_5066,N_2400,N_3142);
and U5067 (N_5067,N_31,N_1645);
or U5068 (N_5068,N_929,N_1320);
or U5069 (N_5069,N_1862,N_1427);
and U5070 (N_5070,N_2726,N_915);
or U5071 (N_5071,N_1731,N_1245);
or U5072 (N_5072,N_1128,N_961);
and U5073 (N_5073,N_2440,N_1110);
nor U5074 (N_5074,N_3416,N_2657);
nor U5075 (N_5075,N_3342,N_2382);
nand U5076 (N_5076,N_3669,N_1574);
nor U5077 (N_5077,N_1260,N_641);
nor U5078 (N_5078,N_398,N_562);
nand U5079 (N_5079,N_3338,N_1742);
and U5080 (N_5080,N_292,N_1511);
nand U5081 (N_5081,N_2035,N_1209);
or U5082 (N_5082,N_437,N_242);
or U5083 (N_5083,N_657,N_1418);
nor U5084 (N_5084,N_2766,N_2378);
nand U5085 (N_5085,N_3415,N_2186);
or U5086 (N_5086,N_3283,N_2203);
or U5087 (N_5087,N_2499,N_788);
nor U5088 (N_5088,N_3136,N_441);
and U5089 (N_5089,N_3042,N_1585);
or U5090 (N_5090,N_375,N_1568);
nor U5091 (N_5091,N_3574,N_3149);
and U5092 (N_5092,N_1985,N_1293);
nor U5093 (N_5093,N_2273,N_1506);
nor U5094 (N_5094,N_980,N_2830);
or U5095 (N_5095,N_457,N_1777);
and U5096 (N_5096,N_1907,N_2889);
and U5097 (N_5097,N_768,N_1887);
or U5098 (N_5098,N_2051,N_2060);
or U5099 (N_5099,N_2840,N_3010);
and U5100 (N_5100,N_3277,N_826);
nand U5101 (N_5101,N_556,N_2184);
nor U5102 (N_5102,N_1120,N_3420);
or U5103 (N_5103,N_2587,N_3854);
nand U5104 (N_5104,N_2038,N_3896);
or U5105 (N_5105,N_777,N_1532);
nand U5106 (N_5106,N_3997,N_995);
and U5107 (N_5107,N_1133,N_1112);
nor U5108 (N_5108,N_857,N_1913);
nand U5109 (N_5109,N_1178,N_3894);
nand U5110 (N_5110,N_204,N_2528);
nand U5111 (N_5111,N_2791,N_2888);
nor U5112 (N_5112,N_1747,N_2131);
nand U5113 (N_5113,N_1708,N_886);
and U5114 (N_5114,N_2742,N_1380);
and U5115 (N_5115,N_3762,N_736);
or U5116 (N_5116,N_2121,N_3591);
nor U5117 (N_5117,N_2802,N_3190);
or U5118 (N_5118,N_785,N_1644);
or U5119 (N_5119,N_1084,N_1188);
nand U5120 (N_5120,N_2483,N_3091);
nor U5121 (N_5121,N_1302,N_3441);
nand U5122 (N_5122,N_203,N_3434);
nor U5123 (N_5123,N_3771,N_3438);
nor U5124 (N_5124,N_3166,N_1766);
and U5125 (N_5125,N_2728,N_2686);
nor U5126 (N_5126,N_3593,N_3196);
or U5127 (N_5127,N_2244,N_378);
nand U5128 (N_5128,N_3621,N_1672);
nand U5129 (N_5129,N_3458,N_2029);
or U5130 (N_5130,N_3220,N_824);
or U5131 (N_5131,N_1702,N_1602);
and U5132 (N_5132,N_1922,N_790);
nor U5133 (N_5133,N_3271,N_2919);
or U5134 (N_5134,N_2881,N_543);
nor U5135 (N_5135,N_3025,N_2349);
and U5136 (N_5136,N_607,N_1224);
and U5137 (N_5137,N_3761,N_3879);
nand U5138 (N_5138,N_3853,N_2185);
or U5139 (N_5139,N_3590,N_3433);
or U5140 (N_5140,N_1257,N_3958);
and U5141 (N_5141,N_3088,N_3113);
nand U5142 (N_5142,N_2178,N_3712);
nor U5143 (N_5143,N_475,N_3930);
nand U5144 (N_5144,N_1715,N_1061);
and U5145 (N_5145,N_3139,N_2584);
and U5146 (N_5146,N_2362,N_721);
and U5147 (N_5147,N_1042,N_510);
or U5148 (N_5148,N_421,N_1485);
nor U5149 (N_5149,N_2788,N_119);
or U5150 (N_5150,N_1199,N_1171);
or U5151 (N_5151,N_1090,N_1794);
and U5152 (N_5152,N_2829,N_1403);
or U5153 (N_5153,N_3294,N_3187);
nor U5154 (N_5154,N_3657,N_3536);
and U5155 (N_5155,N_525,N_3161);
nor U5156 (N_5156,N_868,N_2415);
nor U5157 (N_5157,N_3918,N_3923);
nor U5158 (N_5158,N_182,N_2455);
or U5159 (N_5159,N_828,N_544);
nor U5160 (N_5160,N_3305,N_576);
nand U5161 (N_5161,N_3707,N_3596);
and U5162 (N_5162,N_2477,N_2128);
and U5163 (N_5163,N_3671,N_2883);
or U5164 (N_5164,N_2037,N_3124);
and U5165 (N_5165,N_1014,N_3260);
nand U5166 (N_5166,N_2270,N_2644);
and U5167 (N_5167,N_3750,N_1306);
nand U5168 (N_5168,N_1804,N_3154);
nand U5169 (N_5169,N_3731,N_2713);
nand U5170 (N_5170,N_942,N_2843);
or U5171 (N_5171,N_2744,N_1827);
nand U5172 (N_5172,N_3758,N_3686);
nand U5173 (N_5173,N_3843,N_3);
nand U5174 (N_5174,N_3937,N_13);
nand U5175 (N_5175,N_660,N_1949);
and U5176 (N_5176,N_740,N_1251);
and U5177 (N_5177,N_1082,N_3125);
nand U5178 (N_5178,N_390,N_1191);
nor U5179 (N_5179,N_3334,N_1754);
or U5180 (N_5180,N_2817,N_2124);
and U5181 (N_5181,N_2559,N_937);
nor U5182 (N_5182,N_3557,N_1056);
nand U5183 (N_5183,N_3463,N_878);
and U5184 (N_5184,N_2547,N_683);
or U5185 (N_5185,N_2154,N_494);
nor U5186 (N_5186,N_3740,N_1018);
and U5187 (N_5187,N_1664,N_547);
or U5188 (N_5188,N_2077,N_1610);
nand U5189 (N_5189,N_3261,N_648);
or U5190 (N_5190,N_2976,N_1699);
or U5191 (N_5191,N_703,N_1792);
nand U5192 (N_5192,N_1859,N_3385);
and U5193 (N_5193,N_117,N_644);
nor U5194 (N_5194,N_1588,N_1457);
and U5195 (N_5195,N_2471,N_3044);
or U5196 (N_5196,N_2167,N_2356);
and U5197 (N_5197,N_3692,N_1303);
and U5198 (N_5198,N_1225,N_3919);
nand U5199 (N_5199,N_3904,N_3788);
nand U5200 (N_5200,N_3728,N_1471);
and U5201 (N_5201,N_1910,N_505);
and U5202 (N_5202,N_661,N_3114);
nor U5203 (N_5203,N_1716,N_1974);
nor U5204 (N_5204,N_3467,N_802);
nor U5205 (N_5205,N_77,N_2893);
nor U5206 (N_5206,N_3773,N_3386);
nor U5207 (N_5207,N_382,N_459);
nand U5208 (N_5208,N_3387,N_496);
or U5209 (N_5209,N_315,N_3777);
nand U5210 (N_5210,N_3210,N_1271);
nor U5211 (N_5211,N_1281,N_3205);
nor U5212 (N_5212,N_1019,N_3235);
nand U5213 (N_5213,N_3335,N_3426);
or U5214 (N_5214,N_3093,N_595);
or U5215 (N_5215,N_2207,N_2129);
xor U5216 (N_5216,N_1530,N_2057);
or U5217 (N_5217,N_1236,N_3856);
or U5218 (N_5218,N_1527,N_3649);
and U5219 (N_5219,N_2317,N_896);
nor U5220 (N_5220,N_2226,N_3099);
nand U5221 (N_5221,N_3589,N_3237);
and U5222 (N_5222,N_34,N_2538);
nand U5223 (N_5223,N_3540,N_2453);
and U5224 (N_5224,N_747,N_1809);
or U5225 (N_5225,N_3810,N_329);
or U5226 (N_5226,N_2468,N_2497);
or U5227 (N_5227,N_3846,N_2287);
nor U5228 (N_5228,N_2328,N_2993);
and U5229 (N_5229,N_1,N_1682);
or U5230 (N_5230,N_2900,N_3003);
and U5231 (N_5231,N_2639,N_1522);
and U5232 (N_5232,N_372,N_2826);
nand U5233 (N_5233,N_1036,N_640);
and U5234 (N_5234,N_1474,N_2911);
and U5235 (N_5235,N_2067,N_1473);
or U5236 (N_5236,N_2348,N_2338);
nand U5237 (N_5237,N_596,N_3975);
nand U5238 (N_5238,N_2509,N_668);
or U5239 (N_5239,N_2315,N_735);
nor U5240 (N_5240,N_2225,N_1265);
and U5241 (N_5241,N_900,N_569);
nor U5242 (N_5242,N_448,N_3164);
and U5243 (N_5243,N_1611,N_3084);
nand U5244 (N_5244,N_1518,N_1951);
nand U5245 (N_5245,N_958,N_3517);
or U5246 (N_5246,N_1309,N_2952);
nand U5247 (N_5247,N_2336,N_502);
and U5248 (N_5248,N_2819,N_764);
or U5249 (N_5249,N_577,N_2340);
nor U5250 (N_5250,N_2125,N_2623);
nor U5251 (N_5251,N_3765,N_3827);
nor U5252 (N_5252,N_3455,N_1490);
or U5253 (N_5253,N_870,N_1069);
nor U5254 (N_5254,N_2595,N_2426);
and U5255 (N_5255,N_2062,N_3016);
nor U5256 (N_5256,N_301,N_2467);
or U5257 (N_5257,N_3770,N_1114);
and U5258 (N_5258,N_89,N_1315);
and U5259 (N_5259,N_1440,N_3296);
nor U5260 (N_5260,N_964,N_2680);
and U5261 (N_5261,N_1157,N_3619);
nand U5262 (N_5262,N_1262,N_687);
and U5263 (N_5263,N_998,N_2006);
and U5264 (N_5264,N_882,N_1713);
nand U5265 (N_5265,N_1819,N_1546);
and U5266 (N_5266,N_3186,N_2741);
nand U5267 (N_5267,N_3572,N_1814);
and U5268 (N_5268,N_1931,N_2844);
nor U5269 (N_5269,N_3382,N_248);
xnor U5270 (N_5270,N_677,N_240);
nand U5271 (N_5271,N_2815,N_458);
nand U5272 (N_5272,N_632,N_2122);
nor U5273 (N_5273,N_1571,N_2504);
or U5274 (N_5274,N_2360,N_578);
nand U5275 (N_5275,N_3898,N_2924);
nor U5276 (N_5276,N_3907,N_2195);
nor U5277 (N_5277,N_2868,N_1963);
and U5278 (N_5278,N_1200,N_3179);
nand U5279 (N_5279,N_2403,N_817);
nand U5280 (N_5280,N_71,N_3183);
nor U5281 (N_5281,N_136,N_1650);
nor U5282 (N_5282,N_1854,N_1470);
nor U5283 (N_5283,N_3306,N_3984);
or U5284 (N_5284,N_2230,N_3234);
or U5285 (N_5285,N_2066,N_1994);
nand U5286 (N_5286,N_1743,N_412);
nor U5287 (N_5287,N_2837,N_366);
and U5288 (N_5288,N_1815,N_2855);
or U5289 (N_5289,N_2775,N_3955);
and U5290 (N_5290,N_1865,N_3301);
nand U5291 (N_5291,N_2451,N_93);
and U5292 (N_5292,N_258,N_763);
nand U5293 (N_5293,N_3337,N_3024);
or U5294 (N_5294,N_323,N_2368);
or U5295 (N_5295,N_2940,N_46);
nor U5296 (N_5296,N_3889,N_2165);
and U5297 (N_5297,N_3033,N_2296);
nor U5298 (N_5298,N_2943,N_634);
xnor U5299 (N_5299,N_1138,N_206);
or U5300 (N_5300,N_1640,N_82);
or U5301 (N_5301,N_589,N_3675);
nand U5302 (N_5302,N_1009,N_2284);
nand U5303 (N_5303,N_324,N_3529);
and U5304 (N_5304,N_1206,N_271);
nor U5305 (N_5305,N_3676,N_2918);
nor U5306 (N_5306,N_1227,N_1595);
nor U5307 (N_5307,N_825,N_3732);
nand U5308 (N_5308,N_3535,N_2827);
nor U5309 (N_5309,N_3004,N_617);
and U5310 (N_5310,N_2253,N_1476);
nor U5311 (N_5311,N_922,N_3602);
nand U5312 (N_5312,N_1321,N_1912);
and U5313 (N_5313,N_3605,N_2080);
nand U5314 (N_5314,N_3880,N_2245);
nand U5315 (N_5315,N_729,N_3486);
and U5316 (N_5316,N_1965,N_2365);
and U5317 (N_5317,N_930,N_3174);
and U5318 (N_5318,N_912,N_2656);
nor U5319 (N_5319,N_2611,N_2074);
nor U5320 (N_5320,N_3759,N_3729);
nand U5321 (N_5321,N_778,N_123);
and U5322 (N_5322,N_3212,N_3365);
and U5323 (N_5323,N_1428,N_1134);
and U5324 (N_5324,N_1338,N_428);
nor U5325 (N_5325,N_3638,N_225);
or U5326 (N_5326,N_188,N_3782);
nand U5327 (N_5327,N_1728,N_1973);
nor U5328 (N_5328,N_2849,N_131);
nor U5329 (N_5329,N_224,N_1564);
nor U5330 (N_5330,N_3643,N_3031);
nor U5331 (N_5331,N_773,N_1336);
nor U5332 (N_5332,N_945,N_2678);
or U5333 (N_5333,N_743,N_2224);
nand U5334 (N_5334,N_585,N_615);
nor U5335 (N_5335,N_2751,N_1940);
and U5336 (N_5336,N_3825,N_1921);
and U5337 (N_5337,N_3897,N_3561);
nor U5338 (N_5338,N_1932,N_2992);
or U5339 (N_5339,N_3368,N_2434);
nand U5340 (N_5340,N_2720,N_3472);
nor U5341 (N_5341,N_3285,N_532);
nor U5342 (N_5342,N_286,N_2043);
nand U5343 (N_5343,N_3799,N_3647);
nor U5344 (N_5344,N_3715,N_436);
nor U5345 (N_5345,N_2446,N_2329);
and U5346 (N_5346,N_3541,N_3606);
xor U5347 (N_5347,N_2643,N_3130);
and U5348 (N_5348,N_3059,N_2243);
nand U5349 (N_5349,N_1149,N_1256);
nor U5350 (N_5350,N_3523,N_1591);
nand U5351 (N_5351,N_406,N_3443);
nor U5352 (N_5352,N_1772,N_2589);
and U5353 (N_5353,N_2546,N_3265);
or U5354 (N_5354,N_1420,N_774);
or U5355 (N_5355,N_1478,N_1186);
nand U5356 (N_5356,N_3974,N_446);
nor U5357 (N_5357,N_3137,N_3038);
or U5358 (N_5358,N_2381,N_3470);
nand U5359 (N_5359,N_1524,N_477);
and U5360 (N_5360,N_128,N_989);
nand U5361 (N_5361,N_342,N_3419);
or U5362 (N_5362,N_2833,N_2862);
nor U5363 (N_5363,N_2407,N_3410);
nor U5364 (N_5364,N_221,N_3558);
nor U5365 (N_5365,N_1196,N_3272);
or U5366 (N_5366,N_1152,N_2754);
or U5367 (N_5367,N_1272,N_1322);
nor U5368 (N_5368,N_2098,N_245);
nand U5369 (N_5369,N_3035,N_693);
nor U5370 (N_5370,N_3688,N_2095);
nand U5371 (N_5371,N_3926,N_3700);
nor U5372 (N_5372,N_3494,N_651);
or U5373 (N_5373,N_90,N_1741);
nand U5374 (N_5374,N_1541,N_470);
nand U5375 (N_5375,N_2119,N_3207);
nand U5376 (N_5376,N_247,N_3367);
and U5377 (N_5377,N_3803,N_2469);
and U5378 (N_5378,N_1439,N_254);
nand U5379 (N_5379,N_3681,N_2158);
and U5380 (N_5380,N_720,N_3942);
nand U5381 (N_5381,N_612,N_3600);
and U5382 (N_5382,N_1717,N_1674);
nand U5383 (N_5383,N_2876,N_2541);
or U5384 (N_5384,N_229,N_1041);
and U5385 (N_5385,N_1353,N_1253);
xnor U5386 (N_5386,N_255,N_3929);
nand U5387 (N_5387,N_3464,N_1755);
or U5388 (N_5388,N_2200,N_3495);
and U5389 (N_5389,N_2443,N_1995);
and U5390 (N_5390,N_14,N_691);
or U5391 (N_5391,N_341,N_1280);
or U5392 (N_5392,N_403,N_2383);
nor U5393 (N_5393,N_1711,N_1695);
and U5394 (N_5394,N_3871,N_3527);
and U5395 (N_5395,N_2220,N_2172);
nand U5396 (N_5396,N_3556,N_2449);
or U5397 (N_5397,N_1448,N_3567);
and U5398 (N_5398,N_3951,N_2904);
and U5399 (N_5399,N_1730,N_2747);
nor U5400 (N_5400,N_3868,N_752);
nand U5401 (N_5401,N_3714,N_53);
nand U5402 (N_5402,N_916,N_861);
nand U5403 (N_5403,N_471,N_1670);
nand U5404 (N_5404,N_1481,N_371);
nand U5405 (N_5405,N_2613,N_3779);
nor U5406 (N_5406,N_4,N_2301);
nand U5407 (N_5407,N_3295,N_2757);
nand U5408 (N_5408,N_460,N_2737);
nand U5409 (N_5409,N_263,N_1582);
and U5410 (N_5410,N_3959,N_1273);
nand U5411 (N_5411,N_3988,N_2873);
nor U5412 (N_5412,N_3422,N_633);
nand U5413 (N_5413,N_2655,N_1475);
and U5414 (N_5414,N_1698,N_3000);
and U5415 (N_5415,N_2189,N_2885);
or U5416 (N_5416,N_1658,N_1663);
nor U5417 (N_5417,N_1217,N_232);
or U5418 (N_5418,N_1387,N_1130);
and U5419 (N_5419,N_3162,N_8);
or U5420 (N_5420,N_685,N_384);
and U5421 (N_5421,N_1489,N_2169);
or U5422 (N_5422,N_328,N_474);
or U5423 (N_5423,N_1447,N_3966);
or U5424 (N_5424,N_1737,N_2174);
nor U5425 (N_5425,N_1416,N_2750);
and U5426 (N_5426,N_2130,N_782);
or U5427 (N_5427,N_2514,N_3499);
nand U5428 (N_5428,N_2104,N_3144);
nand U5429 (N_5429,N_3916,N_2822);
or U5430 (N_5430,N_3835,N_2333);
nor U5431 (N_5431,N_705,N_1707);
nand U5432 (N_5432,N_419,N_2712);
xor U5433 (N_5433,N_1826,N_600);
nand U5434 (N_5434,N_257,N_1908);
nand U5435 (N_5435,N_223,N_2624);
or U5436 (N_5436,N_2866,N_1123);
or U5437 (N_5437,N_3112,N_1279);
and U5438 (N_5438,N_2964,N_2256);
and U5439 (N_5439,N_2298,N_1537);
or U5440 (N_5440,N_1838,N_2527);
xnor U5441 (N_5441,N_1957,N_1124);
nand U5442 (N_5442,N_3706,N_690);
nand U5443 (N_5443,N_1797,N_3437);
xor U5444 (N_5444,N_3447,N_1643);
nor U5445 (N_5445,N_936,N_62);
or U5446 (N_5446,N_605,N_268);
nand U5447 (N_5447,N_1685,N_529);
or U5448 (N_5448,N_2498,N_196);
nand U5449 (N_5449,N_3032,N_564);
or U5450 (N_5450,N_1517,N_1990);
or U5451 (N_5451,N_2159,N_2162);
nor U5452 (N_5452,N_297,N_3289);
nand U5453 (N_5453,N_3255,N_6);
nand U5454 (N_5454,N_1333,N_3068);
nor U5455 (N_5455,N_862,N_725);
and U5456 (N_5456,N_189,N_3086);
and U5457 (N_5457,N_3406,N_1396);
nand U5458 (N_5458,N_2161,N_1501);
and U5459 (N_5459,N_2413,N_2264);
or U5460 (N_5460,N_804,N_2157);
and U5461 (N_5461,N_2070,N_368);
and U5462 (N_5462,N_1878,N_103);
or U5463 (N_5463,N_1563,N_843);
nor U5464 (N_5464,N_2241,N_365);
nor U5465 (N_5465,N_1093,N_3217);
nand U5466 (N_5466,N_1618,N_3515);
nor U5467 (N_5467,N_955,N_3060);
or U5468 (N_5468,N_3017,N_3169);
and U5469 (N_5469,N_2188,N_2959);
or U5470 (N_5470,N_2738,N_2151);
and U5471 (N_5471,N_872,N_3317);
or U5472 (N_5472,N_3872,N_792);
nor U5473 (N_5473,N_515,N_1477);
and U5474 (N_5474,N_3251,N_775);
and U5475 (N_5475,N_676,N_1562);
nor U5476 (N_5476,N_2648,N_3449);
nor U5477 (N_5477,N_2946,N_1195);
nor U5478 (N_5478,N_3256,N_2765);
nand U5479 (N_5479,N_2229,N_455);
nand U5480 (N_5480,N_2675,N_3191);
or U5481 (N_5481,N_2481,N_1752);
or U5482 (N_5482,N_3901,N_1402);
and U5483 (N_5483,N_3512,N_1780);
and U5484 (N_5484,N_712,N_3226);
and U5485 (N_5485,N_3014,N_1964);
or U5486 (N_5486,N_716,N_2928);
and U5487 (N_5487,N_2774,N_935);
nand U5488 (N_5488,N_551,N_3702);
and U5489 (N_5489,N_1370,N_1906);
or U5490 (N_5490,N_1748,N_3840);
and U5491 (N_5491,N_1760,N_427);
or U5492 (N_5492,N_2345,N_1364);
nor U5493 (N_5493,N_1356,N_2927);
and U5494 (N_5494,N_2600,N_12);
or U5495 (N_5495,N_156,N_939);
nor U5496 (N_5496,N_2416,N_2198);
or U5497 (N_5497,N_2685,N_664);
or U5498 (N_5498,N_513,N_54);
xnor U5499 (N_5499,N_2518,N_1453);
nor U5500 (N_5500,N_3232,N_3768);
nor U5501 (N_5501,N_604,N_2318);
or U5502 (N_5502,N_2452,N_3550);
or U5503 (N_5503,N_2755,N_3242);
or U5504 (N_5504,N_3222,N_3165);
and U5505 (N_5505,N_3145,N_3430);
and U5506 (N_5506,N_1525,N_1669);
or U5507 (N_5507,N_3180,N_3699);
nand U5508 (N_5508,N_856,N_179);
nand U5509 (N_5509,N_1635,N_1993);
or U5510 (N_5510,N_1641,N_2409);
and U5511 (N_5511,N_3956,N_941);
nand U5512 (N_5512,N_3742,N_2808);
nor U5513 (N_5513,N_1867,N_16);
or U5514 (N_5514,N_3554,N_1889);
and U5515 (N_5515,N_499,N_2797);
nor U5516 (N_5516,N_41,N_2008);
and U5517 (N_5517,N_2988,N_172);
nand U5518 (N_5518,N_1378,N_3177);
or U5519 (N_5519,N_1687,N_3219);
and U5520 (N_5520,N_3812,N_2227);
or U5521 (N_5521,N_986,N_3530);
or U5522 (N_5522,N_1529,N_2510);
or U5523 (N_5523,N_67,N_1051);
nor U5524 (N_5524,N_1219,N_684);
or U5525 (N_5525,N_1981,N_2304);
nor U5526 (N_5526,N_2221,N_185);
nor U5527 (N_5527,N_480,N_601);
nor U5528 (N_5528,N_3198,N_3489);
and U5529 (N_5529,N_924,N_3015);
and U5530 (N_5530,N_1375,N_671);
or U5531 (N_5531,N_917,N_1239);
nor U5532 (N_5532,N_3484,N_3584);
nor U5533 (N_5533,N_2419,N_2984);
and U5534 (N_5534,N_1461,N_1632);
nand U5535 (N_5535,N_1576,N_3949);
nand U5536 (N_5536,N_15,N_1122);
nor U5537 (N_5537,N_1724,N_2364);
and U5538 (N_5538,N_3733,N_61);
or U5539 (N_5539,N_820,N_3625);
nand U5540 (N_5540,N_781,N_1798);
nand U5541 (N_5541,N_2168,N_3481);
nand U5542 (N_5542,N_2553,N_2995);
nand U5543 (N_5543,N_1148,N_1247);
nor U5544 (N_5544,N_3887,N_1575);
nand U5545 (N_5545,N_3980,N_319);
nand U5546 (N_5546,N_2795,N_3767);
nand U5547 (N_5547,N_1901,N_2658);
nor U5548 (N_5548,N_228,N_426);
or U5549 (N_5549,N_3297,N_2981);
or U5550 (N_5550,N_2135,N_1768);
nand U5551 (N_5551,N_3934,N_3111);
or U5552 (N_5552,N_2782,N_3781);
nand U5553 (N_5553,N_23,N_1341);
or U5554 (N_5554,N_3241,N_383);
nand U5555 (N_5555,N_2505,N_1074);
nand U5556 (N_5556,N_1512,N_3423);
or U5557 (N_5557,N_863,N_1683);
nand U5558 (N_5558,N_1745,N_2259);
and U5559 (N_5559,N_3453,N_586);
or U5560 (N_5560,N_2210,N_1115);
xnor U5561 (N_5561,N_2196,N_126);
nand U5562 (N_5562,N_1977,N_1696);
nand U5563 (N_5563,N_2424,N_1877);
or U5564 (N_5564,N_718,N_3171);
nor U5565 (N_5565,N_1007,N_1371);
or U5566 (N_5566,N_1343,N_2930);
nand U5567 (N_5567,N_2717,N_875);
or U5568 (N_5568,N_787,N_356);
and U5569 (N_5569,N_766,N_2033);
nand U5570 (N_5570,N_1519,N_3936);
nand U5571 (N_5571,N_1210,N_2137);
and U5572 (N_5572,N_473,N_464);
nor U5573 (N_5573,N_3195,N_1166);
or U5574 (N_5574,N_238,N_2784);
nor U5575 (N_5575,N_3628,N_1808);
or U5576 (N_5576,N_2108,N_829);
and U5577 (N_5577,N_3978,N_2617);
nand U5578 (N_5578,N_3293,N_3534);
and U5579 (N_5579,N_2783,N_2878);
and U5580 (N_5580,N_3129,N_2758);
nand U5581 (N_5581,N_1806,N_2566);
and U5582 (N_5582,N_1958,N_1078);
nand U5583 (N_5583,N_1185,N_737);
nor U5584 (N_5584,N_681,N_2948);
and U5585 (N_5585,N_3131,N_1666);
nor U5586 (N_5586,N_3011,N_813);
nand U5587 (N_5587,N_3108,N_2916);
nand U5588 (N_5588,N_1287,N_2279);
or U5589 (N_5589,N_481,N_2859);
xor U5590 (N_5590,N_1179,N_3888);
nand U5591 (N_5591,N_3273,N_1433);
and U5592 (N_5592,N_3491,N_3440);
nor U5593 (N_5593,N_987,N_3552);
nor U5594 (N_5594,N_144,N_276);
or U5595 (N_5595,N_416,N_118);
or U5596 (N_5596,N_706,N_1811);
and U5597 (N_5597,N_1639,N_1844);
nand U5598 (N_5598,N_39,N_2288);
or U5599 (N_5599,N_3865,N_3380);
nand U5600 (N_5600,N_1729,N_3292);
or U5601 (N_5601,N_1156,N_2947);
xnor U5602 (N_5602,N_1004,N_2242);
and U5603 (N_5603,N_1570,N_3020);
or U5604 (N_5604,N_2536,N_1616);
nand U5605 (N_5605,N_2722,N_2696);
nor U5606 (N_5606,N_2049,N_503);
or U5607 (N_5607,N_946,N_452);
and U5608 (N_5608,N_2513,N_521);
nand U5609 (N_5609,N_488,N_2886);
nand U5610 (N_5610,N_2682,N_410);
and U5611 (N_5611,N_137,N_2410);
and U5612 (N_5612,N_3245,N_2334);
nor U5613 (N_5613,N_709,N_1314);
or U5614 (N_5614,N_3877,N_3193);
nor U5615 (N_5615,N_3176,N_2111);
or U5616 (N_5616,N_3333,N_674);
and U5617 (N_5617,N_2459,N_1789);
nand U5618 (N_5618,N_3963,N_1305);
nor U5619 (N_5619,N_278,N_3724);
and U5620 (N_5620,N_2663,N_489);
or U5621 (N_5621,N_1366,N_2805);
and U5622 (N_5622,N_413,N_2435);
or U5623 (N_5623,N_1621,N_3436);
or U5624 (N_5624,N_3233,N_2724);
and U5625 (N_5625,N_112,N_2132);
nand U5626 (N_5626,N_686,N_831);
nand U5627 (N_5627,N_566,N_2746);
and U5628 (N_5628,N_1330,N_415);
and U5629 (N_5629,N_3579,N_2887);
and U5630 (N_5630,N_1401,N_487);
or U5631 (N_5631,N_2078,N_3257);
or U5632 (N_5632,N_334,N_2626);
or U5633 (N_5633,N_3039,N_1414);
and U5634 (N_5634,N_536,N_2922);
or U5635 (N_5635,N_1659,N_3658);
nand U5636 (N_5636,N_1818,N_122);
or U5637 (N_5637,N_58,N_3717);
nand U5638 (N_5638,N_1915,N_1350);
or U5639 (N_5639,N_2183,N_2138);
or U5640 (N_5640,N_2748,N_2040);
nor U5641 (N_5641,N_3299,N_2);
and U5642 (N_5642,N_3818,N_393);
nand U5643 (N_5643,N_3996,N_2484);
or U5644 (N_5644,N_1880,N_124);
nand U5645 (N_5645,N_3178,N_524);
or U5646 (N_5646,N_698,N_2293);
nor U5647 (N_5647,N_1339,N_3836);
nand U5648 (N_5648,N_66,N_2598);
or U5649 (N_5649,N_1006,N_2305);
and U5650 (N_5650,N_1839,N_1083);
and U5651 (N_5651,N_1828,N_2762);
or U5652 (N_5652,N_3970,N_3148);
nor U5653 (N_5653,N_960,N_877);
and U5654 (N_5654,N_3445,N_2099);
nand U5655 (N_5655,N_1494,N_3642);
and U5656 (N_5656,N_1686,N_2351);
or U5657 (N_5657,N_1516,N_739);
nand U5658 (N_5658,N_303,N_3230);
nor U5659 (N_5659,N_801,N_290);
nor U5660 (N_5660,N_3543,N_949);
nor U5661 (N_5661,N_2437,N_3236);
or U5662 (N_5662,N_2173,N_1928);
nor U5663 (N_5663,N_3064,N_295);
and U5664 (N_5664,N_1254,N_2281);
nand U5665 (N_5665,N_535,N_1637);
nor U5666 (N_5666,N_646,N_3944);
nand U5667 (N_5667,N_2123,N_3547);
and U5668 (N_5668,N_3428,N_2523);
and U5669 (N_5669,N_1551,N_2250);
nand U5670 (N_5670,N_3852,N_3048);
or U5671 (N_5671,N_1340,N_2938);
nor U5672 (N_5672,N_3200,N_3533);
and U5673 (N_5673,N_3008,N_343);
nor U5674 (N_5674,N_2487,N_1633);
xor U5675 (N_5675,N_2571,N_349);
and U5676 (N_5676,N_3726,N_669);
nor U5677 (N_5677,N_2971,N_2633);
or U5678 (N_5678,N_2730,N_3248);
and U5679 (N_5679,N_3156,N_573);
and U5680 (N_5680,N_1445,N_2386);
nor U5681 (N_5681,N_2707,N_274);
and U5682 (N_5682,N_2902,N_3309);
and U5683 (N_5683,N_2090,N_2436);
xnor U5684 (N_5684,N_3322,N_630);
nand U5685 (N_5685,N_2820,N_2201);
nor U5686 (N_5686,N_318,N_3622);
nand U5687 (N_5687,N_285,N_1369);
nand U5688 (N_5688,N_2690,N_3976);
nor U5689 (N_5689,N_1388,N_2384);
nor U5690 (N_5690,N_2420,N_1043);
nor U5691 (N_5691,N_1992,N_3341);
and U5692 (N_5692,N_1802,N_3268);
nor U5693 (N_5693,N_3776,N_3343);
or U5694 (N_5694,N_3451,N_166);
nand U5695 (N_5695,N_944,N_1318);
or U5696 (N_5696,N_537,N_1298);
and U5697 (N_5697,N_506,N_3610);
nand U5698 (N_5698,N_2581,N_619);
nand U5699 (N_5699,N_2065,N_1464);
nand U5700 (N_5700,N_3291,N_1759);
nor U5701 (N_5701,N_2594,N_2856);
nand U5702 (N_5702,N_2734,N_3276);
nor U5703 (N_5703,N_3747,N_1631);
or U5704 (N_5704,N_2969,N_1864);
and U5705 (N_5705,N_582,N_3667);
nor U5706 (N_5706,N_3993,N_663);
or U5707 (N_5707,N_394,N_654);
or U5708 (N_5708,N_2249,N_312);
and U5709 (N_5709,N_3192,N_2417);
nand U5710 (N_5710,N_3247,N_3409);
nand U5711 (N_5711,N_3356,N_3321);
nor U5712 (N_5712,N_2271,N_2767);
and U5713 (N_5713,N_3908,N_3960);
nor U5714 (N_5714,N_3315,N_3749);
and U5715 (N_5715,N_3078,N_979);
and U5716 (N_5716,N_338,N_1627);
and U5717 (N_5717,N_3211,N_2237);
and U5718 (N_5718,N_3266,N_3525);
or U5719 (N_5719,N_1141,N_2586);
nand U5720 (N_5720,N_2715,N_3832);
nand U5721 (N_5721,N_3964,N_3469);
or U5722 (N_5722,N_147,N_2580);
or U5723 (N_5723,N_3838,N_1504);
and U5724 (N_5724,N_1557,N_1107);
or U5725 (N_5725,N_3372,N_2380);
nand U5726 (N_5726,N_1352,N_3539);
or U5727 (N_5727,N_1984,N_610);
and U5728 (N_5728,N_3465,N_3607);
nand U5729 (N_5729,N_2404,N_2501);
or U5730 (N_5730,N_361,N_2578);
or U5731 (N_5731,N_130,N_175);
or U5732 (N_5732,N_2599,N_190);
nand U5733 (N_5733,N_1484,N_871);
or U5734 (N_5734,N_1140,N_967);
or U5735 (N_5735,N_2208,N_3903);
nor U5736 (N_5736,N_1535,N_3891);
nand U5737 (N_5737,N_3569,N_381);
nor U5738 (N_5738,N_2627,N_3214);
or U5739 (N_5739,N_2973,N_568);
nand U5740 (N_5740,N_1288,N_2194);
nand U5741 (N_5741,N_538,N_1896);
and U5742 (N_5742,N_3708,N_2697);
or U5743 (N_5743,N_805,N_463);
xor U5744 (N_5744,N_753,N_2806);
nand U5745 (N_5745,N_3583,N_1800);
and U5746 (N_5746,N_267,N_822);
or U5747 (N_5747,N_3476,N_1894);
nand U5748 (N_5748,N_3994,N_3116);
and U5749 (N_5749,N_1812,N_314);
nand U5750 (N_5750,N_88,N_626);
and U5751 (N_5751,N_42,N_2853);
or U5752 (N_5752,N_1357,N_11);
nand U5753 (N_5753,N_1775,N_102);
nor U5754 (N_5754,N_1646,N_1622);
nand U5755 (N_5755,N_3346,N_3103);
and U5756 (N_5756,N_798,N_2248);
and U5757 (N_5757,N_1500,N_3575);
and U5758 (N_5758,N_2909,N_3935);
and U5759 (N_5759,N_3140,N_2604);
nand U5760 (N_5760,N_1016,N_3213);
or U5761 (N_5761,N_1174,N_110);
or U5762 (N_5762,N_2506,N_3488);
or U5763 (N_5763,N_975,N_2980);
nand U5764 (N_5764,N_3006,N_2920);
and U5765 (N_5765,N_925,N_1691);
nand U5766 (N_5766,N_901,N_1334);
nand U5767 (N_5767,N_3188,N_3795);
nand U5768 (N_5768,N_1230,N_1274);
nor U5769 (N_5769,N_1498,N_1203);
or U5770 (N_5770,N_3805,N_241);
xnor U5771 (N_5771,N_1349,N_1923);
nand U5772 (N_5772,N_1088,N_2772);
nand U5773 (N_5773,N_1689,N_1825);
or U5774 (N_5774,N_293,N_3905);
or U5775 (N_5775,N_3787,N_3651);
nor U5776 (N_5776,N_2860,N_3155);
nor U5777 (N_5777,N_1598,N_402);
xnor U5778 (N_5778,N_3381,N_977);
and U5779 (N_5779,N_3324,N_869);
nor U5780 (N_5780,N_3007,N_1783);
or U5781 (N_5781,N_2816,N_2733);
nand U5782 (N_5782,N_3862,N_1240);
and U5783 (N_5783,N_3107,N_2217);
and U5784 (N_5784,N_3209,N_3968);
nand U5785 (N_5785,N_846,N_3143);
or U5786 (N_5786,N_597,N_2810);
nor U5787 (N_5787,N_3566,N_2082);
or U5788 (N_5788,N_1066,N_2610);
nor U5789 (N_5789,N_482,N_948);
nand U5790 (N_5790,N_430,N_2127);
and U5791 (N_5791,N_442,N_2913);
xnor U5792 (N_5792,N_227,N_2083);
and U5793 (N_5793,N_3617,N_1147);
nor U5794 (N_5794,N_3240,N_570);
and U5795 (N_5795,N_2529,N_602);
or U5796 (N_5796,N_1012,N_2251);
and U5797 (N_5797,N_3194,N_2294);
nand U5798 (N_5798,N_894,N_1703);
nand U5799 (N_5799,N_1558,N_32);
nor U5800 (N_5800,N_1890,N_2535);
or U5801 (N_5801,N_2936,N_2291);
and U5802 (N_5802,N_3218,N_347);
nor U5803 (N_5803,N_951,N_2721);
nand U5804 (N_5804,N_2941,N_3745);
and U5805 (N_5805,N_2785,N_2957);
and U5806 (N_5806,N_2464,N_2780);
and U5807 (N_5807,N_2861,N_1628);
nand U5808 (N_5808,N_1213,N_3693);
and U5809 (N_5809,N_279,N_339);
and U5810 (N_5810,N_3735,N_638);
nand U5811 (N_5811,N_1238,N_2768);
or U5812 (N_5812,N_1037,N_3056);
nor U5813 (N_5813,N_3080,N_2649);
nand U5814 (N_5814,N_727,N_2719);
and U5815 (N_5815,N_1011,N_757);
nand U5816 (N_5816,N_2593,N_3629);
and U5817 (N_5817,N_860,N_2880);
and U5818 (N_5818,N_3823,N_2170);
nor U5819 (N_5819,N_1269,N_3648);
and U5820 (N_5820,N_710,N_867);
and U5821 (N_5821,N_890,N_3135);
nand U5822 (N_5822,N_1208,N_1569);
nor U5823 (N_5823,N_583,N_3564);
or U5824 (N_5824,N_2760,N_3403);
nor U5825 (N_5825,N_3775,N_1226);
or U5826 (N_5826,N_2014,N_806);
and U5827 (N_5827,N_1189,N_1482);
nand U5828 (N_5828,N_3262,N_1411);
or U5829 (N_5829,N_163,N_3800);
or U5830 (N_5830,N_1392,N_749);
nand U5831 (N_5831,N_3875,N_3347);
or U5832 (N_5832,N_2929,N_1376);
or U5833 (N_5833,N_3216,N_2792);
or U5834 (N_5834,N_3034,N_3694);
nand U5835 (N_5835,N_679,N_1421);
and U5836 (N_5836,N_3374,N_3001);
nand U5837 (N_5837,N_250,N_1654);
and U5838 (N_5838,N_33,N_2520);
nor U5839 (N_5839,N_561,N_3264);
nor U5840 (N_5840,N_3811,N_3371);
or U5841 (N_5841,N_1077,N_3696);
and U5842 (N_5842,N_2825,N_3801);
nor U5843 (N_5843,N_2181,N_2262);
or U5844 (N_5844,N_3442,N_3674);
nor U5845 (N_5845,N_1264,N_2490);
nand U5846 (N_5846,N_3990,N_3851);
or U5847 (N_5847,N_1738,N_3490);
nor U5848 (N_5848,N_1769,N_3911);
or U5849 (N_5849,N_125,N_2372);
nand U5850 (N_5850,N_2740,N_3627);
nor U5851 (N_5851,N_3506,N_3520);
and U5852 (N_5852,N_2140,N_209);
xor U5853 (N_5853,N_539,N_3100);
or U5854 (N_5854,N_1462,N_1385);
nand U5855 (N_5855,N_3603,N_1192);
nand U5856 (N_5856,N_652,N_317);
and U5857 (N_5857,N_1444,N_1638);
nor U5858 (N_5858,N_2650,N_3350);
nand U5859 (N_5859,N_1996,N_3595);
and U5860 (N_5860,N_1400,N_3577);
or U5861 (N_5861,N_73,N_3132);
nor U5862 (N_5862,N_3429,N_1381);
nand U5863 (N_5863,N_1547,N_1136);
nand U5864 (N_5864,N_3570,N_1952);
nor U5865 (N_5865,N_2454,N_2414);
and U5866 (N_5866,N_1292,N_3842);
or U5867 (N_5867,N_2689,N_3581);
or U5868 (N_5868,N_3957,N_1704);
nand U5869 (N_5869,N_3834,N_796);
nor U5870 (N_5870,N_3316,N_2736);
or U5871 (N_5871,N_1454,N_3848);
and U5872 (N_5872,N_60,N_1127);
or U5873 (N_5873,N_3361,N_3133);
and U5874 (N_5874,N_1493,N_2548);
xnor U5875 (N_5875,N_522,N_2401);
nor U5876 (N_5876,N_3662,N_3751);
nor U5877 (N_5877,N_1727,N_2966);
or U5878 (N_5878,N_697,N_1869);
nor U5879 (N_5879,N_2811,N_1422);
and U5880 (N_5880,N_3754,N_557);
nor U5881 (N_5881,N_3349,N_3736);
or U5882 (N_5882,N_2102,N_1554);
nand U5883 (N_5883,N_3089,N_35);
or U5884 (N_5884,N_1151,N_1331);
and U5885 (N_5885,N_3252,N_2931);
or U5886 (N_5886,N_1863,N_3689);
or U5887 (N_5887,N_2319,N_913);
or U5888 (N_5888,N_3555,N_2834);
nor U5889 (N_5889,N_959,N_3755);
nor U5890 (N_5890,N_320,N_631);
nor U5891 (N_5891,N_572,N_2233);
or U5892 (N_5892,N_2235,N_563);
or U5893 (N_5893,N_95,N_1190);
nand U5894 (N_5894,N_3991,N_1596);
or U5895 (N_5895,N_821,N_3061);
nor U5896 (N_5896,N_1117,N_1710);
or U5897 (N_5897,N_3826,N_2552);
or U5898 (N_5898,N_1848,N_83);
nand U5899 (N_5899,N_2605,N_2246);
nand U5900 (N_5900,N_783,N_2907);
nand U5901 (N_5901,N_1681,N_880);
or U5902 (N_5902,N_3683,N_1879);
nor U5903 (N_5903,N_3620,N_1572);
nor U5904 (N_5904,N_3158,N_2275);
nor U5905 (N_5905,N_1617,N_2056);
or U5906 (N_5906,N_1834,N_2009);
nand U5907 (N_5907,N_3379,N_2411);
nor U5908 (N_5908,N_2978,N_120);
xnor U5909 (N_5909,N_2526,N_2522);
nand U5910 (N_5910,N_541,N_3654);
and U5911 (N_5911,N_799,N_3398);
nand U5912 (N_5912,N_590,N_1967);
nand U5913 (N_5913,N_3548,N_2910);
or U5914 (N_5914,N_1235,N_1057);
nand U5915 (N_5915,N_1386,N_3258);
nor U5916 (N_5916,N_3098,N_3351);
or U5917 (N_5917,N_409,N_2672);
nor U5918 (N_5918,N_1872,N_891);
nor U5919 (N_5919,N_3448,N_1555);
or U5920 (N_5920,N_235,N_3882);
nand U5921 (N_5921,N_304,N_3407);
or U5922 (N_5922,N_2550,N_3270);
or U5923 (N_5923,N_1359,N_1135);
or U5924 (N_5924,N_1326,N_2954);
nor U5925 (N_5925,N_1765,N_217);
nand U5926 (N_5926,N_396,N_2322);
nand U5927 (N_5927,N_3698,N_1456);
nor U5928 (N_5928,N_3987,N_331);
or U5929 (N_5929,N_30,N_3480);
and U5930 (N_5930,N_1175,N_369);
nand U5931 (N_5931,N_1329,N_3650);
and U5932 (N_5932,N_2654,N_2299);
nor U5933 (N_5933,N_2048,N_1521);
nor U5934 (N_5934,N_2405,N_197);
xor U5935 (N_5935,N_2486,N_3435);
nand U5936 (N_5936,N_2337,N_3075);
nand U5937 (N_5937,N_1062,N_614);
nand U5938 (N_5938,N_2502,N_1176);
nand U5939 (N_5939,N_1567,N_2071);
nor U5940 (N_5940,N_3999,N_623);
nand U5941 (N_5941,N_337,N_1791);
or U5942 (N_5942,N_74,N_854);
and U5943 (N_5943,N_3375,N_3456);
and U5944 (N_5944,N_1026,N_2018);
nor U5945 (N_5945,N_3121,N_2845);
and U5946 (N_5946,N_1183,N_1221);
and U5947 (N_5947,N_1267,N_1297);
or U5948 (N_5948,N_1324,N_2752);
and U5949 (N_5949,N_316,N_354);
nand U5950 (N_5950,N_3049,N_3404);
nand U5951 (N_5951,N_1753,N_793);
nand U5952 (N_5952,N_1902,N_3680);
or U5953 (N_5953,N_259,N_3287);
or U5954 (N_5954,N_1034,N_44);
nor U5955 (N_5955,N_2031,N_168);
or U5956 (N_5956,N_1139,N_1720);
nand U5957 (N_5957,N_840,N_2863);
nor U5958 (N_5958,N_719,N_1328);
and U5959 (N_5959,N_1065,N_1044);
nand U5960 (N_5960,N_3454,N_1049);
nand U5961 (N_5961,N_3910,N_3563);
and U5962 (N_5962,N_606,N_2793);
and U5963 (N_5963,N_918,N_732);
nor U5964 (N_5964,N_3353,N_553);
nand U5965 (N_5965,N_855,N_3026);
nor U5966 (N_5966,N_2912,N_1258);
or U5967 (N_5967,N_528,N_3159);
nand U5968 (N_5968,N_2055,N_2193);
nand U5969 (N_5969,N_273,N_17);
nor U5970 (N_5970,N_2019,N_978);
nand U5971 (N_5971,N_2709,N_1467);
and U5972 (N_5972,N_1855,N_212);
and U5973 (N_5973,N_2781,N_3953);
and U5974 (N_5974,N_3705,N_2004);
and U5975 (N_5975,N_1560,N_3259);
or U5976 (N_5976,N_2136,N_1997);
nand U5977 (N_5977,N_3329,N_3831);
nand U5978 (N_5978,N_2096,N_2489);
nor U5979 (N_5979,N_1487,N_3592);
nand U5980 (N_5980,N_575,N_2017);
nor U5981 (N_5981,N_264,N_377);
and U5982 (N_5982,N_952,N_3895);
or U5983 (N_5983,N_504,N_2223);
nand U5984 (N_5984,N_2005,N_2222);
or U5985 (N_5985,N_2093,N_3421);
or U5986 (N_5986,N_1027,N_3246);
nand U5987 (N_5987,N_3336,N_3551);
nor U5988 (N_5988,N_1821,N_1903);
and U5989 (N_5989,N_135,N_1182);
and U5990 (N_5990,N_2375,N_3710);
and U5991 (N_5991,N_1930,N_1442);
nand U5992 (N_5992,N_1220,N_2601);
and U5993 (N_5993,N_3766,N_1979);
nor U5994 (N_5994,N_3967,N_155);
or U5995 (N_5995,N_25,N_1216);
and U5996 (N_5996,N_1393,N_3542);
and U5997 (N_5997,N_2024,N_3302);
and U5998 (N_5998,N_643,N_1193);
nand U5999 (N_5999,N_3344,N_2871);
and U6000 (N_6000,N_2725,N_3876);
nor U6001 (N_6001,N_113,N_2548);
nand U6002 (N_6002,N_2818,N_2732);
nand U6003 (N_6003,N_3035,N_2716);
nand U6004 (N_6004,N_2006,N_3389);
and U6005 (N_6005,N_213,N_2950);
or U6006 (N_6006,N_2384,N_3942);
nand U6007 (N_6007,N_2421,N_3893);
nor U6008 (N_6008,N_3987,N_3342);
nor U6009 (N_6009,N_1950,N_3945);
nor U6010 (N_6010,N_935,N_3095);
nor U6011 (N_6011,N_599,N_2281);
and U6012 (N_6012,N_101,N_2052);
or U6013 (N_6013,N_1419,N_2576);
nor U6014 (N_6014,N_3329,N_129);
or U6015 (N_6015,N_3294,N_3604);
nand U6016 (N_6016,N_2245,N_3562);
nand U6017 (N_6017,N_3543,N_2801);
and U6018 (N_6018,N_234,N_1698);
nand U6019 (N_6019,N_1500,N_3224);
and U6020 (N_6020,N_1824,N_447);
nor U6021 (N_6021,N_1432,N_471);
and U6022 (N_6022,N_2498,N_90);
or U6023 (N_6023,N_2012,N_363);
nand U6024 (N_6024,N_3580,N_660);
and U6025 (N_6025,N_3183,N_2448);
nand U6026 (N_6026,N_786,N_3606);
nand U6027 (N_6027,N_2592,N_3469);
and U6028 (N_6028,N_2308,N_1093);
nor U6029 (N_6029,N_2458,N_316);
nand U6030 (N_6030,N_3027,N_3275);
nor U6031 (N_6031,N_1019,N_1703);
or U6032 (N_6032,N_2378,N_389);
and U6033 (N_6033,N_3432,N_2678);
nand U6034 (N_6034,N_471,N_2383);
and U6035 (N_6035,N_600,N_3486);
nor U6036 (N_6036,N_2178,N_2245);
or U6037 (N_6037,N_2542,N_1527);
or U6038 (N_6038,N_3239,N_2186);
nor U6039 (N_6039,N_3121,N_3498);
and U6040 (N_6040,N_3855,N_1110);
nand U6041 (N_6041,N_1788,N_1925);
nand U6042 (N_6042,N_1971,N_1569);
or U6043 (N_6043,N_1187,N_570);
and U6044 (N_6044,N_2300,N_3094);
nand U6045 (N_6045,N_1931,N_1158);
and U6046 (N_6046,N_1850,N_3160);
nand U6047 (N_6047,N_1008,N_1348);
and U6048 (N_6048,N_1833,N_2824);
or U6049 (N_6049,N_3361,N_1700);
or U6050 (N_6050,N_2784,N_2131);
nand U6051 (N_6051,N_2839,N_1785);
nor U6052 (N_6052,N_696,N_3516);
or U6053 (N_6053,N_448,N_192);
nand U6054 (N_6054,N_1443,N_2720);
nand U6055 (N_6055,N_217,N_2020);
and U6056 (N_6056,N_840,N_142);
nand U6057 (N_6057,N_2707,N_3645);
and U6058 (N_6058,N_642,N_2976);
nor U6059 (N_6059,N_1646,N_411);
nor U6060 (N_6060,N_2026,N_3640);
and U6061 (N_6061,N_2173,N_757);
nor U6062 (N_6062,N_3374,N_3227);
nor U6063 (N_6063,N_1138,N_1506);
nand U6064 (N_6064,N_2318,N_3342);
or U6065 (N_6065,N_2369,N_1895);
nor U6066 (N_6066,N_3886,N_3594);
nand U6067 (N_6067,N_455,N_3617);
and U6068 (N_6068,N_290,N_3004);
or U6069 (N_6069,N_2420,N_2021);
and U6070 (N_6070,N_2021,N_1637);
and U6071 (N_6071,N_505,N_2433);
and U6072 (N_6072,N_2160,N_2044);
and U6073 (N_6073,N_3600,N_113);
nor U6074 (N_6074,N_3647,N_2756);
nand U6075 (N_6075,N_1895,N_1379);
or U6076 (N_6076,N_870,N_1324);
and U6077 (N_6077,N_1055,N_1617);
nor U6078 (N_6078,N_1147,N_2181);
nand U6079 (N_6079,N_621,N_1623);
and U6080 (N_6080,N_600,N_3988);
or U6081 (N_6081,N_2395,N_2009);
and U6082 (N_6082,N_1564,N_2406);
and U6083 (N_6083,N_2928,N_3907);
nand U6084 (N_6084,N_1262,N_752);
nor U6085 (N_6085,N_3174,N_877);
nand U6086 (N_6086,N_1324,N_3667);
or U6087 (N_6087,N_1607,N_1105);
nor U6088 (N_6088,N_3719,N_524);
and U6089 (N_6089,N_3516,N_1060);
nor U6090 (N_6090,N_3751,N_1413);
nand U6091 (N_6091,N_363,N_2963);
nor U6092 (N_6092,N_1708,N_3020);
and U6093 (N_6093,N_2226,N_1209);
nand U6094 (N_6094,N_11,N_3893);
and U6095 (N_6095,N_3976,N_608);
nor U6096 (N_6096,N_1322,N_3322);
and U6097 (N_6097,N_1872,N_1244);
or U6098 (N_6098,N_3391,N_1846);
and U6099 (N_6099,N_2085,N_1727);
nand U6100 (N_6100,N_1199,N_64);
nor U6101 (N_6101,N_3688,N_60);
and U6102 (N_6102,N_1234,N_931);
or U6103 (N_6103,N_3045,N_605);
nand U6104 (N_6104,N_3708,N_303);
and U6105 (N_6105,N_3839,N_45);
nor U6106 (N_6106,N_1783,N_1239);
and U6107 (N_6107,N_3586,N_3422);
nor U6108 (N_6108,N_2924,N_2480);
nand U6109 (N_6109,N_1424,N_2966);
nand U6110 (N_6110,N_2320,N_3893);
nor U6111 (N_6111,N_2481,N_1704);
or U6112 (N_6112,N_2763,N_2833);
and U6113 (N_6113,N_2926,N_1108);
nand U6114 (N_6114,N_3765,N_796);
or U6115 (N_6115,N_1788,N_3925);
nor U6116 (N_6116,N_1468,N_1915);
and U6117 (N_6117,N_989,N_3369);
or U6118 (N_6118,N_819,N_577);
or U6119 (N_6119,N_2379,N_139);
or U6120 (N_6120,N_2393,N_804);
or U6121 (N_6121,N_553,N_2912);
or U6122 (N_6122,N_3358,N_3246);
nor U6123 (N_6123,N_1430,N_716);
nor U6124 (N_6124,N_3244,N_641);
nand U6125 (N_6125,N_848,N_2602);
or U6126 (N_6126,N_1384,N_852);
and U6127 (N_6127,N_721,N_1471);
and U6128 (N_6128,N_2723,N_1848);
or U6129 (N_6129,N_3664,N_2421);
or U6130 (N_6130,N_1631,N_2703);
or U6131 (N_6131,N_1361,N_2905);
nand U6132 (N_6132,N_32,N_3325);
and U6133 (N_6133,N_714,N_2303);
and U6134 (N_6134,N_1586,N_88);
nand U6135 (N_6135,N_2270,N_2989);
and U6136 (N_6136,N_834,N_2221);
nand U6137 (N_6137,N_2011,N_3347);
xnor U6138 (N_6138,N_1143,N_707);
nand U6139 (N_6139,N_2450,N_496);
nor U6140 (N_6140,N_2002,N_2872);
and U6141 (N_6141,N_2249,N_2963);
and U6142 (N_6142,N_1825,N_2885);
and U6143 (N_6143,N_3944,N_2812);
and U6144 (N_6144,N_3438,N_3062);
and U6145 (N_6145,N_423,N_602);
and U6146 (N_6146,N_3915,N_2400);
nand U6147 (N_6147,N_3547,N_2079);
or U6148 (N_6148,N_3680,N_2713);
nand U6149 (N_6149,N_929,N_1995);
nand U6150 (N_6150,N_26,N_2504);
or U6151 (N_6151,N_464,N_1102);
nor U6152 (N_6152,N_3488,N_162);
and U6153 (N_6153,N_515,N_3541);
nand U6154 (N_6154,N_3667,N_2141);
nand U6155 (N_6155,N_251,N_2728);
or U6156 (N_6156,N_1408,N_3501);
or U6157 (N_6157,N_2625,N_3821);
or U6158 (N_6158,N_3059,N_1312);
or U6159 (N_6159,N_2392,N_814);
or U6160 (N_6160,N_3273,N_1878);
or U6161 (N_6161,N_3290,N_246);
or U6162 (N_6162,N_2312,N_976);
nor U6163 (N_6163,N_225,N_682);
nand U6164 (N_6164,N_1953,N_3465);
nand U6165 (N_6165,N_2021,N_3813);
or U6166 (N_6166,N_1433,N_3274);
nand U6167 (N_6167,N_1217,N_3284);
or U6168 (N_6168,N_2474,N_1444);
and U6169 (N_6169,N_2104,N_2854);
nand U6170 (N_6170,N_2216,N_3436);
nand U6171 (N_6171,N_3094,N_833);
and U6172 (N_6172,N_1685,N_1320);
nor U6173 (N_6173,N_3230,N_3407);
nand U6174 (N_6174,N_2079,N_508);
and U6175 (N_6175,N_1260,N_2126);
and U6176 (N_6176,N_1177,N_3113);
nand U6177 (N_6177,N_692,N_835);
and U6178 (N_6178,N_933,N_1497);
and U6179 (N_6179,N_1666,N_2318);
nor U6180 (N_6180,N_1262,N_1257);
or U6181 (N_6181,N_3647,N_879);
nor U6182 (N_6182,N_2807,N_2881);
nor U6183 (N_6183,N_3014,N_1948);
or U6184 (N_6184,N_2190,N_181);
nor U6185 (N_6185,N_1135,N_3024);
or U6186 (N_6186,N_3082,N_3641);
nor U6187 (N_6187,N_84,N_3149);
and U6188 (N_6188,N_3080,N_2880);
and U6189 (N_6189,N_1853,N_2382);
and U6190 (N_6190,N_2298,N_1707);
or U6191 (N_6191,N_2857,N_2796);
nor U6192 (N_6192,N_1911,N_3297);
nand U6193 (N_6193,N_2210,N_1610);
and U6194 (N_6194,N_821,N_2016);
and U6195 (N_6195,N_817,N_714);
or U6196 (N_6196,N_108,N_184);
and U6197 (N_6197,N_2688,N_397);
nor U6198 (N_6198,N_573,N_1007);
or U6199 (N_6199,N_770,N_2021);
nand U6200 (N_6200,N_1808,N_2142);
or U6201 (N_6201,N_454,N_3069);
nand U6202 (N_6202,N_2259,N_3565);
nand U6203 (N_6203,N_3547,N_1068);
nor U6204 (N_6204,N_3780,N_326);
nor U6205 (N_6205,N_3883,N_2781);
or U6206 (N_6206,N_3199,N_122);
or U6207 (N_6207,N_3453,N_1221);
and U6208 (N_6208,N_615,N_423);
nand U6209 (N_6209,N_300,N_1457);
and U6210 (N_6210,N_1418,N_741);
nand U6211 (N_6211,N_2117,N_3473);
and U6212 (N_6212,N_2295,N_2992);
nor U6213 (N_6213,N_3453,N_2511);
nor U6214 (N_6214,N_2314,N_2501);
or U6215 (N_6215,N_1538,N_2575);
nand U6216 (N_6216,N_715,N_559);
and U6217 (N_6217,N_3636,N_3158);
or U6218 (N_6218,N_2716,N_3205);
nor U6219 (N_6219,N_1661,N_858);
and U6220 (N_6220,N_398,N_602);
nor U6221 (N_6221,N_47,N_3599);
or U6222 (N_6222,N_1907,N_2001);
or U6223 (N_6223,N_3272,N_1270);
nand U6224 (N_6224,N_1850,N_59);
nand U6225 (N_6225,N_1387,N_3664);
nor U6226 (N_6226,N_2797,N_2125);
or U6227 (N_6227,N_1164,N_3373);
nand U6228 (N_6228,N_3197,N_2992);
nor U6229 (N_6229,N_2825,N_3159);
nor U6230 (N_6230,N_2567,N_649);
nor U6231 (N_6231,N_1421,N_1198);
or U6232 (N_6232,N_2982,N_1754);
or U6233 (N_6233,N_1383,N_2403);
nand U6234 (N_6234,N_3803,N_2575);
nand U6235 (N_6235,N_3512,N_1224);
or U6236 (N_6236,N_2430,N_1981);
nor U6237 (N_6237,N_1024,N_870);
nand U6238 (N_6238,N_2110,N_2259);
nor U6239 (N_6239,N_2011,N_1836);
nand U6240 (N_6240,N_3898,N_2876);
nor U6241 (N_6241,N_1898,N_2202);
and U6242 (N_6242,N_2945,N_3755);
nand U6243 (N_6243,N_2094,N_3076);
or U6244 (N_6244,N_3108,N_562);
nor U6245 (N_6245,N_1192,N_2009);
or U6246 (N_6246,N_637,N_3128);
and U6247 (N_6247,N_308,N_2576);
xor U6248 (N_6248,N_976,N_2103);
and U6249 (N_6249,N_2454,N_96);
and U6250 (N_6250,N_3918,N_3668);
and U6251 (N_6251,N_2901,N_3614);
nand U6252 (N_6252,N_386,N_2339);
and U6253 (N_6253,N_2958,N_1102);
and U6254 (N_6254,N_3636,N_3253);
or U6255 (N_6255,N_1605,N_1381);
nand U6256 (N_6256,N_11,N_1005);
and U6257 (N_6257,N_1893,N_2242);
and U6258 (N_6258,N_946,N_2616);
nor U6259 (N_6259,N_2515,N_402);
nor U6260 (N_6260,N_137,N_1340);
and U6261 (N_6261,N_3821,N_2655);
nor U6262 (N_6262,N_2003,N_1897);
or U6263 (N_6263,N_2030,N_129);
nor U6264 (N_6264,N_2682,N_2311);
or U6265 (N_6265,N_728,N_1884);
and U6266 (N_6266,N_3424,N_3775);
nor U6267 (N_6267,N_3420,N_1053);
nor U6268 (N_6268,N_3641,N_3536);
and U6269 (N_6269,N_3936,N_645);
nand U6270 (N_6270,N_479,N_3943);
or U6271 (N_6271,N_1228,N_3867);
nand U6272 (N_6272,N_3720,N_1351);
nand U6273 (N_6273,N_2385,N_204);
nor U6274 (N_6274,N_924,N_94);
nand U6275 (N_6275,N_1518,N_1341);
and U6276 (N_6276,N_2652,N_1064);
nor U6277 (N_6277,N_3792,N_1407);
and U6278 (N_6278,N_3121,N_1576);
nand U6279 (N_6279,N_327,N_3822);
or U6280 (N_6280,N_1267,N_112);
or U6281 (N_6281,N_3937,N_2929);
or U6282 (N_6282,N_1294,N_950);
nand U6283 (N_6283,N_3378,N_369);
or U6284 (N_6284,N_2761,N_3480);
and U6285 (N_6285,N_2954,N_709);
and U6286 (N_6286,N_1445,N_2807);
or U6287 (N_6287,N_1785,N_2491);
or U6288 (N_6288,N_1762,N_1228);
nor U6289 (N_6289,N_1511,N_1950);
and U6290 (N_6290,N_3122,N_604);
nand U6291 (N_6291,N_2955,N_3002);
nor U6292 (N_6292,N_2178,N_183);
or U6293 (N_6293,N_203,N_3254);
nand U6294 (N_6294,N_1753,N_3320);
nand U6295 (N_6295,N_2999,N_3053);
and U6296 (N_6296,N_3791,N_2741);
and U6297 (N_6297,N_350,N_798);
or U6298 (N_6298,N_2243,N_2954);
nand U6299 (N_6299,N_1838,N_3542);
nand U6300 (N_6300,N_2436,N_3038);
and U6301 (N_6301,N_1297,N_3415);
nor U6302 (N_6302,N_3325,N_1157);
or U6303 (N_6303,N_3918,N_2810);
nor U6304 (N_6304,N_1404,N_1857);
nand U6305 (N_6305,N_3832,N_378);
and U6306 (N_6306,N_258,N_826);
and U6307 (N_6307,N_1487,N_2178);
and U6308 (N_6308,N_3019,N_3502);
or U6309 (N_6309,N_3249,N_2512);
or U6310 (N_6310,N_1867,N_3947);
nor U6311 (N_6311,N_1560,N_2663);
and U6312 (N_6312,N_2520,N_1431);
and U6313 (N_6313,N_404,N_3171);
nor U6314 (N_6314,N_3121,N_1387);
or U6315 (N_6315,N_3459,N_1706);
nor U6316 (N_6316,N_1,N_3857);
nand U6317 (N_6317,N_1992,N_2019);
nor U6318 (N_6318,N_1364,N_2480);
or U6319 (N_6319,N_1166,N_560);
nand U6320 (N_6320,N_256,N_520);
and U6321 (N_6321,N_1723,N_846);
nor U6322 (N_6322,N_1833,N_364);
and U6323 (N_6323,N_11,N_2893);
and U6324 (N_6324,N_3274,N_1203);
or U6325 (N_6325,N_729,N_2771);
or U6326 (N_6326,N_2032,N_2489);
nor U6327 (N_6327,N_2450,N_2855);
and U6328 (N_6328,N_3910,N_3077);
and U6329 (N_6329,N_2848,N_2969);
and U6330 (N_6330,N_3154,N_2668);
nand U6331 (N_6331,N_1838,N_3626);
or U6332 (N_6332,N_1005,N_589);
and U6333 (N_6333,N_2517,N_3912);
nand U6334 (N_6334,N_1241,N_1563);
nand U6335 (N_6335,N_84,N_65);
nor U6336 (N_6336,N_2214,N_3028);
nand U6337 (N_6337,N_3922,N_2989);
and U6338 (N_6338,N_3610,N_405);
nand U6339 (N_6339,N_3261,N_2410);
nor U6340 (N_6340,N_545,N_1050);
and U6341 (N_6341,N_3709,N_3624);
nand U6342 (N_6342,N_3455,N_2534);
nand U6343 (N_6343,N_136,N_547);
nor U6344 (N_6344,N_3734,N_3728);
or U6345 (N_6345,N_3270,N_123);
nand U6346 (N_6346,N_3386,N_716);
and U6347 (N_6347,N_1806,N_1439);
or U6348 (N_6348,N_2001,N_292);
nor U6349 (N_6349,N_2365,N_2466);
nor U6350 (N_6350,N_3054,N_3667);
nor U6351 (N_6351,N_3889,N_2987);
nand U6352 (N_6352,N_870,N_3907);
nand U6353 (N_6353,N_2052,N_3848);
nand U6354 (N_6354,N_1346,N_3068);
and U6355 (N_6355,N_2246,N_1607);
nand U6356 (N_6356,N_3911,N_3563);
nand U6357 (N_6357,N_1151,N_2781);
or U6358 (N_6358,N_487,N_3553);
or U6359 (N_6359,N_3210,N_362);
and U6360 (N_6360,N_2605,N_1729);
and U6361 (N_6361,N_1336,N_3191);
or U6362 (N_6362,N_148,N_2041);
and U6363 (N_6363,N_277,N_1829);
or U6364 (N_6364,N_2764,N_777);
or U6365 (N_6365,N_3944,N_3106);
nor U6366 (N_6366,N_2797,N_3843);
and U6367 (N_6367,N_2109,N_1709);
nor U6368 (N_6368,N_1431,N_2060);
or U6369 (N_6369,N_3316,N_2927);
nand U6370 (N_6370,N_3193,N_80);
or U6371 (N_6371,N_2722,N_1048);
nor U6372 (N_6372,N_1170,N_3598);
and U6373 (N_6373,N_2274,N_1042);
or U6374 (N_6374,N_2052,N_3588);
or U6375 (N_6375,N_3697,N_62);
and U6376 (N_6376,N_1188,N_3360);
and U6377 (N_6377,N_3489,N_435);
or U6378 (N_6378,N_1412,N_1562);
nand U6379 (N_6379,N_3003,N_2842);
or U6380 (N_6380,N_617,N_183);
nor U6381 (N_6381,N_1446,N_2306);
and U6382 (N_6382,N_2624,N_1593);
nand U6383 (N_6383,N_272,N_347);
nand U6384 (N_6384,N_1198,N_734);
or U6385 (N_6385,N_3488,N_3129);
or U6386 (N_6386,N_3556,N_2552);
or U6387 (N_6387,N_2568,N_3262);
nand U6388 (N_6388,N_1425,N_7);
and U6389 (N_6389,N_3708,N_3730);
nand U6390 (N_6390,N_967,N_3408);
and U6391 (N_6391,N_1164,N_3258);
and U6392 (N_6392,N_3736,N_1393);
nor U6393 (N_6393,N_1736,N_2886);
or U6394 (N_6394,N_161,N_364);
nand U6395 (N_6395,N_3594,N_2454);
and U6396 (N_6396,N_2855,N_2201);
nand U6397 (N_6397,N_750,N_97);
or U6398 (N_6398,N_199,N_1134);
nand U6399 (N_6399,N_3329,N_2841);
or U6400 (N_6400,N_2659,N_1365);
and U6401 (N_6401,N_3556,N_3495);
and U6402 (N_6402,N_1583,N_830);
or U6403 (N_6403,N_1364,N_1537);
nor U6404 (N_6404,N_468,N_250);
nand U6405 (N_6405,N_1401,N_1002);
nor U6406 (N_6406,N_2210,N_950);
or U6407 (N_6407,N_75,N_754);
and U6408 (N_6408,N_3495,N_2384);
nor U6409 (N_6409,N_3611,N_2600);
or U6410 (N_6410,N_2276,N_1039);
nor U6411 (N_6411,N_3511,N_3813);
and U6412 (N_6412,N_588,N_968);
or U6413 (N_6413,N_1007,N_671);
nor U6414 (N_6414,N_1558,N_339);
nor U6415 (N_6415,N_2289,N_2724);
nor U6416 (N_6416,N_427,N_523);
nor U6417 (N_6417,N_235,N_3535);
and U6418 (N_6418,N_750,N_3492);
nor U6419 (N_6419,N_3764,N_948);
or U6420 (N_6420,N_32,N_411);
nand U6421 (N_6421,N_1263,N_3862);
nor U6422 (N_6422,N_1234,N_2248);
nor U6423 (N_6423,N_725,N_2908);
and U6424 (N_6424,N_252,N_2742);
and U6425 (N_6425,N_3185,N_273);
nor U6426 (N_6426,N_3931,N_328);
nor U6427 (N_6427,N_2055,N_548);
nand U6428 (N_6428,N_3054,N_3231);
and U6429 (N_6429,N_3129,N_2792);
nand U6430 (N_6430,N_770,N_2017);
and U6431 (N_6431,N_1968,N_821);
nor U6432 (N_6432,N_2498,N_3620);
or U6433 (N_6433,N_2744,N_2079);
nor U6434 (N_6434,N_1012,N_3914);
nor U6435 (N_6435,N_1191,N_1133);
nand U6436 (N_6436,N_1080,N_187);
nor U6437 (N_6437,N_3767,N_3534);
nand U6438 (N_6438,N_1365,N_365);
nand U6439 (N_6439,N_2525,N_1940);
nor U6440 (N_6440,N_472,N_1766);
xor U6441 (N_6441,N_2809,N_3785);
nor U6442 (N_6442,N_1163,N_3891);
nand U6443 (N_6443,N_486,N_566);
nand U6444 (N_6444,N_557,N_2857);
nand U6445 (N_6445,N_1301,N_3909);
and U6446 (N_6446,N_844,N_1681);
nand U6447 (N_6447,N_2441,N_1211);
and U6448 (N_6448,N_2912,N_2983);
or U6449 (N_6449,N_3808,N_812);
nor U6450 (N_6450,N_1618,N_773);
xor U6451 (N_6451,N_798,N_1402);
nor U6452 (N_6452,N_2660,N_2700);
or U6453 (N_6453,N_322,N_3635);
nand U6454 (N_6454,N_3393,N_2374);
nor U6455 (N_6455,N_2292,N_2847);
and U6456 (N_6456,N_1336,N_2687);
nor U6457 (N_6457,N_2314,N_2378);
nor U6458 (N_6458,N_2596,N_1785);
nand U6459 (N_6459,N_2872,N_1166);
or U6460 (N_6460,N_2338,N_3125);
or U6461 (N_6461,N_866,N_1634);
nor U6462 (N_6462,N_76,N_2389);
and U6463 (N_6463,N_3204,N_3671);
or U6464 (N_6464,N_1368,N_3306);
or U6465 (N_6465,N_1090,N_196);
nor U6466 (N_6466,N_337,N_1221);
or U6467 (N_6467,N_969,N_3140);
or U6468 (N_6468,N_2039,N_3316);
and U6469 (N_6469,N_822,N_3525);
and U6470 (N_6470,N_3964,N_1027);
and U6471 (N_6471,N_484,N_2062);
and U6472 (N_6472,N_2055,N_1355);
or U6473 (N_6473,N_3267,N_3676);
nand U6474 (N_6474,N_1974,N_2410);
nor U6475 (N_6475,N_558,N_3019);
nor U6476 (N_6476,N_1131,N_3392);
and U6477 (N_6477,N_953,N_3101);
or U6478 (N_6478,N_1470,N_2863);
nand U6479 (N_6479,N_3383,N_975);
and U6480 (N_6480,N_3300,N_1343);
nor U6481 (N_6481,N_2159,N_2809);
and U6482 (N_6482,N_372,N_1184);
and U6483 (N_6483,N_3117,N_19);
or U6484 (N_6484,N_386,N_2608);
and U6485 (N_6485,N_2121,N_3617);
and U6486 (N_6486,N_820,N_677);
or U6487 (N_6487,N_2418,N_2726);
and U6488 (N_6488,N_999,N_2408);
nand U6489 (N_6489,N_3039,N_2830);
and U6490 (N_6490,N_1682,N_2460);
nand U6491 (N_6491,N_1914,N_2946);
nor U6492 (N_6492,N_1360,N_1584);
and U6493 (N_6493,N_3220,N_2341);
xnor U6494 (N_6494,N_2004,N_524);
nor U6495 (N_6495,N_2511,N_3070);
or U6496 (N_6496,N_1304,N_3554);
nand U6497 (N_6497,N_1003,N_997);
nor U6498 (N_6498,N_3053,N_2693);
or U6499 (N_6499,N_495,N_3260);
and U6500 (N_6500,N_1780,N_3997);
nor U6501 (N_6501,N_1741,N_2470);
nand U6502 (N_6502,N_1370,N_1115);
and U6503 (N_6503,N_1917,N_2370);
nor U6504 (N_6504,N_1109,N_2839);
nor U6505 (N_6505,N_1887,N_1158);
nor U6506 (N_6506,N_3909,N_3463);
nor U6507 (N_6507,N_2112,N_429);
nand U6508 (N_6508,N_2056,N_1203);
nand U6509 (N_6509,N_1450,N_1161);
nor U6510 (N_6510,N_2607,N_3414);
or U6511 (N_6511,N_752,N_400);
nand U6512 (N_6512,N_2142,N_2622);
nand U6513 (N_6513,N_3708,N_1625);
or U6514 (N_6514,N_191,N_1919);
or U6515 (N_6515,N_1067,N_100);
or U6516 (N_6516,N_3715,N_1360);
nor U6517 (N_6517,N_1990,N_3299);
or U6518 (N_6518,N_525,N_2587);
nand U6519 (N_6519,N_3436,N_2230);
nor U6520 (N_6520,N_1317,N_320);
nand U6521 (N_6521,N_1457,N_263);
and U6522 (N_6522,N_1840,N_71);
nor U6523 (N_6523,N_1205,N_1762);
and U6524 (N_6524,N_2044,N_3845);
or U6525 (N_6525,N_3669,N_681);
or U6526 (N_6526,N_763,N_638);
nand U6527 (N_6527,N_1742,N_1219);
nor U6528 (N_6528,N_672,N_3813);
nand U6529 (N_6529,N_1239,N_3905);
and U6530 (N_6530,N_1354,N_3508);
nor U6531 (N_6531,N_3800,N_578);
nor U6532 (N_6532,N_2167,N_757);
and U6533 (N_6533,N_3468,N_1071);
and U6534 (N_6534,N_2613,N_2083);
and U6535 (N_6535,N_1818,N_2794);
nor U6536 (N_6536,N_2954,N_3621);
or U6537 (N_6537,N_694,N_2607);
nand U6538 (N_6538,N_936,N_825);
and U6539 (N_6539,N_3256,N_19);
nand U6540 (N_6540,N_2376,N_2460);
nand U6541 (N_6541,N_3993,N_3367);
nand U6542 (N_6542,N_2575,N_2310);
nor U6543 (N_6543,N_1224,N_2245);
nor U6544 (N_6544,N_1470,N_406);
xor U6545 (N_6545,N_3086,N_3470);
or U6546 (N_6546,N_1825,N_1970);
and U6547 (N_6547,N_3551,N_1975);
or U6548 (N_6548,N_1007,N_2790);
or U6549 (N_6549,N_1161,N_1020);
or U6550 (N_6550,N_3101,N_3343);
nand U6551 (N_6551,N_2970,N_2349);
and U6552 (N_6552,N_116,N_678);
nor U6553 (N_6553,N_1803,N_1033);
and U6554 (N_6554,N_634,N_2490);
nor U6555 (N_6555,N_3682,N_2882);
or U6556 (N_6556,N_3517,N_3537);
and U6557 (N_6557,N_3560,N_1959);
or U6558 (N_6558,N_3763,N_596);
or U6559 (N_6559,N_1253,N_1502);
or U6560 (N_6560,N_1117,N_1876);
and U6561 (N_6561,N_3171,N_2797);
nand U6562 (N_6562,N_1001,N_2841);
or U6563 (N_6563,N_3827,N_987);
nand U6564 (N_6564,N_1375,N_2296);
and U6565 (N_6565,N_98,N_351);
or U6566 (N_6566,N_813,N_2380);
and U6567 (N_6567,N_2720,N_290);
and U6568 (N_6568,N_3099,N_3848);
nor U6569 (N_6569,N_208,N_87);
or U6570 (N_6570,N_2595,N_1968);
xor U6571 (N_6571,N_2745,N_3240);
nand U6572 (N_6572,N_2506,N_221);
nand U6573 (N_6573,N_938,N_1128);
and U6574 (N_6574,N_571,N_393);
nor U6575 (N_6575,N_1007,N_3647);
or U6576 (N_6576,N_3872,N_525);
nand U6577 (N_6577,N_2656,N_1972);
and U6578 (N_6578,N_1576,N_1312);
nand U6579 (N_6579,N_336,N_173);
nor U6580 (N_6580,N_775,N_1221);
and U6581 (N_6581,N_3937,N_3121);
or U6582 (N_6582,N_3832,N_1436);
nor U6583 (N_6583,N_3448,N_2189);
nand U6584 (N_6584,N_2752,N_3025);
and U6585 (N_6585,N_1260,N_144);
and U6586 (N_6586,N_103,N_1902);
or U6587 (N_6587,N_2160,N_697);
nand U6588 (N_6588,N_478,N_1327);
nor U6589 (N_6589,N_1704,N_2589);
and U6590 (N_6590,N_1622,N_1813);
or U6591 (N_6591,N_3868,N_1932);
or U6592 (N_6592,N_2579,N_9);
or U6593 (N_6593,N_1836,N_2802);
and U6594 (N_6594,N_14,N_2899);
and U6595 (N_6595,N_2057,N_3946);
or U6596 (N_6596,N_2760,N_790);
nand U6597 (N_6597,N_1933,N_436);
or U6598 (N_6598,N_3564,N_2776);
and U6599 (N_6599,N_683,N_240);
nand U6600 (N_6600,N_3686,N_1174);
or U6601 (N_6601,N_351,N_131);
nand U6602 (N_6602,N_1116,N_2228);
nand U6603 (N_6603,N_1389,N_3109);
or U6604 (N_6604,N_791,N_2707);
or U6605 (N_6605,N_1915,N_837);
or U6606 (N_6606,N_3954,N_2676);
nor U6607 (N_6607,N_1449,N_127);
and U6608 (N_6608,N_1229,N_2363);
nand U6609 (N_6609,N_2815,N_2774);
or U6610 (N_6610,N_2977,N_3750);
nand U6611 (N_6611,N_3761,N_3953);
and U6612 (N_6612,N_1792,N_2999);
nand U6613 (N_6613,N_537,N_1318);
nand U6614 (N_6614,N_541,N_67);
nor U6615 (N_6615,N_2321,N_2958);
nand U6616 (N_6616,N_2500,N_849);
or U6617 (N_6617,N_1496,N_2086);
and U6618 (N_6618,N_2507,N_1202);
and U6619 (N_6619,N_1435,N_2177);
or U6620 (N_6620,N_193,N_2593);
and U6621 (N_6621,N_2116,N_33);
nor U6622 (N_6622,N_2217,N_2910);
and U6623 (N_6623,N_2191,N_3114);
and U6624 (N_6624,N_1914,N_1128);
nand U6625 (N_6625,N_1495,N_233);
or U6626 (N_6626,N_3255,N_356);
nand U6627 (N_6627,N_3731,N_235);
nor U6628 (N_6628,N_211,N_2120);
nand U6629 (N_6629,N_542,N_3370);
xor U6630 (N_6630,N_1443,N_3862);
nand U6631 (N_6631,N_2152,N_628);
nand U6632 (N_6632,N_216,N_2464);
or U6633 (N_6633,N_3159,N_981);
nand U6634 (N_6634,N_3723,N_2151);
nor U6635 (N_6635,N_3260,N_3876);
nor U6636 (N_6636,N_1952,N_2252);
or U6637 (N_6637,N_1059,N_2562);
and U6638 (N_6638,N_1823,N_901);
nor U6639 (N_6639,N_1084,N_781);
or U6640 (N_6640,N_3625,N_2982);
and U6641 (N_6641,N_3566,N_735);
and U6642 (N_6642,N_293,N_2025);
or U6643 (N_6643,N_2840,N_1924);
nand U6644 (N_6644,N_683,N_935);
or U6645 (N_6645,N_2436,N_3851);
or U6646 (N_6646,N_2202,N_1880);
or U6647 (N_6647,N_3767,N_3101);
nand U6648 (N_6648,N_2748,N_13);
or U6649 (N_6649,N_1398,N_2831);
or U6650 (N_6650,N_3861,N_2750);
nor U6651 (N_6651,N_350,N_3128);
nand U6652 (N_6652,N_1672,N_1526);
and U6653 (N_6653,N_1176,N_1119);
or U6654 (N_6654,N_2400,N_1436);
and U6655 (N_6655,N_626,N_230);
nor U6656 (N_6656,N_3372,N_2580);
nor U6657 (N_6657,N_2576,N_2889);
nand U6658 (N_6658,N_1706,N_2170);
or U6659 (N_6659,N_29,N_3778);
or U6660 (N_6660,N_393,N_2341);
and U6661 (N_6661,N_126,N_2912);
nand U6662 (N_6662,N_603,N_3668);
or U6663 (N_6663,N_3877,N_3069);
and U6664 (N_6664,N_1831,N_1853);
nand U6665 (N_6665,N_3739,N_2252);
nand U6666 (N_6666,N_1862,N_2193);
and U6667 (N_6667,N_906,N_1039);
nor U6668 (N_6668,N_3324,N_3485);
nand U6669 (N_6669,N_2788,N_639);
and U6670 (N_6670,N_2567,N_1761);
or U6671 (N_6671,N_1544,N_3014);
or U6672 (N_6672,N_3015,N_1895);
and U6673 (N_6673,N_2273,N_3617);
or U6674 (N_6674,N_969,N_2428);
and U6675 (N_6675,N_282,N_2810);
or U6676 (N_6676,N_537,N_2180);
and U6677 (N_6677,N_3822,N_84);
nand U6678 (N_6678,N_2347,N_1139);
nor U6679 (N_6679,N_272,N_968);
nand U6680 (N_6680,N_3801,N_3180);
and U6681 (N_6681,N_338,N_724);
nand U6682 (N_6682,N_2618,N_1201);
nand U6683 (N_6683,N_1191,N_2775);
nand U6684 (N_6684,N_3290,N_3059);
nor U6685 (N_6685,N_507,N_2729);
and U6686 (N_6686,N_3157,N_3620);
nand U6687 (N_6687,N_442,N_273);
nand U6688 (N_6688,N_3100,N_3765);
and U6689 (N_6689,N_3596,N_635);
nand U6690 (N_6690,N_3732,N_3606);
nor U6691 (N_6691,N_1275,N_2048);
nand U6692 (N_6692,N_1566,N_2834);
and U6693 (N_6693,N_811,N_23);
and U6694 (N_6694,N_2835,N_1899);
and U6695 (N_6695,N_1769,N_2035);
or U6696 (N_6696,N_2936,N_2649);
nor U6697 (N_6697,N_3539,N_1068);
nand U6698 (N_6698,N_1402,N_1103);
or U6699 (N_6699,N_3339,N_3344);
nor U6700 (N_6700,N_2674,N_940);
nand U6701 (N_6701,N_791,N_578);
and U6702 (N_6702,N_1542,N_1929);
or U6703 (N_6703,N_3831,N_163);
nand U6704 (N_6704,N_3368,N_615);
nor U6705 (N_6705,N_488,N_282);
nand U6706 (N_6706,N_2143,N_2122);
xor U6707 (N_6707,N_3140,N_486);
and U6708 (N_6708,N_3884,N_101);
nor U6709 (N_6709,N_863,N_218);
or U6710 (N_6710,N_1387,N_1214);
nand U6711 (N_6711,N_1599,N_1989);
and U6712 (N_6712,N_2271,N_624);
nand U6713 (N_6713,N_451,N_2963);
and U6714 (N_6714,N_3247,N_1168);
nor U6715 (N_6715,N_1078,N_2992);
or U6716 (N_6716,N_598,N_197);
nand U6717 (N_6717,N_1007,N_2750);
nor U6718 (N_6718,N_444,N_925);
and U6719 (N_6719,N_3428,N_3516);
or U6720 (N_6720,N_1583,N_660);
or U6721 (N_6721,N_1999,N_3304);
nor U6722 (N_6722,N_3178,N_1682);
and U6723 (N_6723,N_2508,N_2423);
or U6724 (N_6724,N_1207,N_1246);
or U6725 (N_6725,N_1642,N_3687);
nand U6726 (N_6726,N_3413,N_2075);
or U6727 (N_6727,N_1778,N_3696);
and U6728 (N_6728,N_1682,N_3675);
or U6729 (N_6729,N_1511,N_3033);
or U6730 (N_6730,N_1010,N_1700);
or U6731 (N_6731,N_3225,N_1930);
nand U6732 (N_6732,N_2773,N_1792);
or U6733 (N_6733,N_1327,N_481);
nor U6734 (N_6734,N_3947,N_1419);
nor U6735 (N_6735,N_1261,N_278);
and U6736 (N_6736,N_435,N_1856);
nor U6737 (N_6737,N_1352,N_809);
nand U6738 (N_6738,N_852,N_2670);
and U6739 (N_6739,N_2489,N_1841);
or U6740 (N_6740,N_1444,N_2161);
nand U6741 (N_6741,N_2310,N_3022);
nand U6742 (N_6742,N_3297,N_2286);
and U6743 (N_6743,N_336,N_1858);
or U6744 (N_6744,N_1613,N_3119);
nor U6745 (N_6745,N_1276,N_3568);
or U6746 (N_6746,N_1712,N_760);
nand U6747 (N_6747,N_2316,N_2861);
and U6748 (N_6748,N_2769,N_1658);
or U6749 (N_6749,N_1257,N_369);
and U6750 (N_6750,N_3838,N_2546);
or U6751 (N_6751,N_141,N_2316);
nand U6752 (N_6752,N_1887,N_1521);
nand U6753 (N_6753,N_3240,N_631);
nand U6754 (N_6754,N_3255,N_1086);
nand U6755 (N_6755,N_3159,N_759);
nor U6756 (N_6756,N_324,N_1867);
or U6757 (N_6757,N_2732,N_551);
and U6758 (N_6758,N_2942,N_2864);
nand U6759 (N_6759,N_2075,N_2881);
or U6760 (N_6760,N_1718,N_3504);
and U6761 (N_6761,N_2127,N_3309);
or U6762 (N_6762,N_674,N_2170);
nand U6763 (N_6763,N_532,N_1627);
nand U6764 (N_6764,N_3569,N_745);
nor U6765 (N_6765,N_1631,N_2244);
nor U6766 (N_6766,N_782,N_3227);
nor U6767 (N_6767,N_3215,N_240);
and U6768 (N_6768,N_2963,N_365);
and U6769 (N_6769,N_560,N_1135);
nor U6770 (N_6770,N_1900,N_412);
and U6771 (N_6771,N_3081,N_264);
nand U6772 (N_6772,N_3003,N_1104);
and U6773 (N_6773,N_1057,N_1728);
or U6774 (N_6774,N_698,N_1105);
nor U6775 (N_6775,N_3602,N_2456);
or U6776 (N_6776,N_3616,N_2614);
nor U6777 (N_6777,N_3997,N_3822);
nor U6778 (N_6778,N_3381,N_2013);
and U6779 (N_6779,N_401,N_2939);
nand U6780 (N_6780,N_3372,N_1828);
nand U6781 (N_6781,N_1513,N_229);
nand U6782 (N_6782,N_969,N_1781);
and U6783 (N_6783,N_222,N_2228);
nor U6784 (N_6784,N_985,N_3908);
nor U6785 (N_6785,N_620,N_2973);
nor U6786 (N_6786,N_1197,N_1877);
or U6787 (N_6787,N_638,N_2764);
or U6788 (N_6788,N_1012,N_2968);
nor U6789 (N_6789,N_3897,N_2338);
nor U6790 (N_6790,N_261,N_3923);
nand U6791 (N_6791,N_2770,N_1771);
or U6792 (N_6792,N_3885,N_2335);
or U6793 (N_6793,N_122,N_2427);
nand U6794 (N_6794,N_3191,N_1649);
or U6795 (N_6795,N_1414,N_274);
and U6796 (N_6796,N_84,N_1328);
and U6797 (N_6797,N_3927,N_2694);
nand U6798 (N_6798,N_726,N_2872);
nor U6799 (N_6799,N_2442,N_3305);
or U6800 (N_6800,N_1802,N_2950);
nor U6801 (N_6801,N_3712,N_3847);
nand U6802 (N_6802,N_1026,N_2040);
nand U6803 (N_6803,N_1266,N_1364);
nor U6804 (N_6804,N_3256,N_223);
nor U6805 (N_6805,N_1333,N_387);
nand U6806 (N_6806,N_954,N_2837);
nand U6807 (N_6807,N_3612,N_2600);
nand U6808 (N_6808,N_150,N_1029);
or U6809 (N_6809,N_1853,N_3852);
nor U6810 (N_6810,N_837,N_3814);
or U6811 (N_6811,N_1676,N_108);
or U6812 (N_6812,N_2491,N_273);
and U6813 (N_6813,N_3852,N_2831);
or U6814 (N_6814,N_2346,N_639);
nand U6815 (N_6815,N_1613,N_1383);
nor U6816 (N_6816,N_2110,N_1198);
or U6817 (N_6817,N_37,N_2235);
nor U6818 (N_6818,N_2838,N_227);
or U6819 (N_6819,N_3253,N_3582);
nor U6820 (N_6820,N_3649,N_3594);
nand U6821 (N_6821,N_200,N_1451);
nor U6822 (N_6822,N_3407,N_199);
or U6823 (N_6823,N_1173,N_2553);
and U6824 (N_6824,N_431,N_1484);
nand U6825 (N_6825,N_3795,N_94);
and U6826 (N_6826,N_463,N_58);
nor U6827 (N_6827,N_287,N_1294);
nor U6828 (N_6828,N_948,N_428);
nand U6829 (N_6829,N_839,N_1156);
or U6830 (N_6830,N_3425,N_1745);
nor U6831 (N_6831,N_3767,N_128);
nand U6832 (N_6832,N_714,N_902);
and U6833 (N_6833,N_1572,N_190);
or U6834 (N_6834,N_418,N_2626);
nand U6835 (N_6835,N_1743,N_1771);
or U6836 (N_6836,N_2667,N_3922);
nand U6837 (N_6837,N_3981,N_1577);
nor U6838 (N_6838,N_3997,N_2224);
or U6839 (N_6839,N_2712,N_281);
and U6840 (N_6840,N_212,N_3333);
and U6841 (N_6841,N_1322,N_985);
nand U6842 (N_6842,N_2138,N_2791);
and U6843 (N_6843,N_3101,N_1201);
nor U6844 (N_6844,N_400,N_1739);
or U6845 (N_6845,N_3676,N_467);
nand U6846 (N_6846,N_1941,N_220);
nand U6847 (N_6847,N_775,N_1854);
nand U6848 (N_6848,N_290,N_1260);
nand U6849 (N_6849,N_3147,N_1290);
nand U6850 (N_6850,N_2136,N_3680);
and U6851 (N_6851,N_1766,N_752);
nor U6852 (N_6852,N_1849,N_1002);
or U6853 (N_6853,N_1973,N_3442);
nor U6854 (N_6854,N_2915,N_2525);
nor U6855 (N_6855,N_1531,N_1844);
nand U6856 (N_6856,N_532,N_3582);
and U6857 (N_6857,N_2057,N_424);
nand U6858 (N_6858,N_531,N_1351);
or U6859 (N_6859,N_1230,N_2799);
or U6860 (N_6860,N_1885,N_3797);
and U6861 (N_6861,N_2199,N_3806);
or U6862 (N_6862,N_3867,N_163);
nor U6863 (N_6863,N_554,N_1535);
or U6864 (N_6864,N_295,N_93);
nand U6865 (N_6865,N_1380,N_3309);
and U6866 (N_6866,N_1060,N_1008);
and U6867 (N_6867,N_3146,N_468);
nand U6868 (N_6868,N_2918,N_1591);
and U6869 (N_6869,N_130,N_1631);
or U6870 (N_6870,N_3272,N_3464);
or U6871 (N_6871,N_3659,N_1513);
nor U6872 (N_6872,N_1419,N_1352);
nand U6873 (N_6873,N_2580,N_3237);
nand U6874 (N_6874,N_3153,N_1196);
nand U6875 (N_6875,N_2067,N_938);
nor U6876 (N_6876,N_598,N_808);
nor U6877 (N_6877,N_652,N_1443);
or U6878 (N_6878,N_493,N_1068);
or U6879 (N_6879,N_1759,N_742);
nor U6880 (N_6880,N_991,N_1979);
nand U6881 (N_6881,N_788,N_2057);
xor U6882 (N_6882,N_2166,N_1415);
nor U6883 (N_6883,N_2327,N_3301);
nor U6884 (N_6884,N_1861,N_1723);
nand U6885 (N_6885,N_2603,N_3438);
nor U6886 (N_6886,N_2662,N_291);
nand U6887 (N_6887,N_978,N_414);
nand U6888 (N_6888,N_1568,N_2979);
nand U6889 (N_6889,N_3949,N_2444);
or U6890 (N_6890,N_3343,N_954);
nand U6891 (N_6891,N_3523,N_3862);
and U6892 (N_6892,N_3426,N_3300);
nand U6893 (N_6893,N_3703,N_3529);
nor U6894 (N_6894,N_3024,N_734);
or U6895 (N_6895,N_1624,N_499);
nand U6896 (N_6896,N_3768,N_1065);
nand U6897 (N_6897,N_3550,N_617);
or U6898 (N_6898,N_2008,N_1762);
nand U6899 (N_6899,N_991,N_3226);
nand U6900 (N_6900,N_3593,N_437);
nor U6901 (N_6901,N_3932,N_1308);
or U6902 (N_6902,N_2891,N_3593);
and U6903 (N_6903,N_737,N_2067);
nand U6904 (N_6904,N_0,N_1080);
and U6905 (N_6905,N_482,N_1641);
or U6906 (N_6906,N_1165,N_1442);
nand U6907 (N_6907,N_1498,N_2770);
nand U6908 (N_6908,N_1478,N_1549);
or U6909 (N_6909,N_2925,N_187);
and U6910 (N_6910,N_401,N_3115);
nand U6911 (N_6911,N_3182,N_2758);
or U6912 (N_6912,N_1877,N_1184);
nor U6913 (N_6913,N_2561,N_1457);
or U6914 (N_6914,N_1022,N_940);
nand U6915 (N_6915,N_769,N_1680);
or U6916 (N_6916,N_3911,N_3593);
nand U6917 (N_6917,N_3191,N_1589);
nor U6918 (N_6918,N_751,N_3594);
or U6919 (N_6919,N_3812,N_610);
nand U6920 (N_6920,N_488,N_3022);
or U6921 (N_6921,N_3087,N_3390);
and U6922 (N_6922,N_2089,N_3520);
or U6923 (N_6923,N_3992,N_3285);
or U6924 (N_6924,N_3314,N_3353);
xor U6925 (N_6925,N_731,N_3771);
nand U6926 (N_6926,N_400,N_3774);
nand U6927 (N_6927,N_3237,N_1154);
nor U6928 (N_6928,N_1373,N_617);
nor U6929 (N_6929,N_2599,N_3681);
and U6930 (N_6930,N_610,N_3454);
or U6931 (N_6931,N_846,N_510);
nor U6932 (N_6932,N_581,N_694);
and U6933 (N_6933,N_2942,N_1833);
or U6934 (N_6934,N_29,N_3738);
nand U6935 (N_6935,N_453,N_1460);
or U6936 (N_6936,N_1131,N_1285);
nand U6937 (N_6937,N_713,N_571);
and U6938 (N_6938,N_177,N_1837);
nand U6939 (N_6939,N_1257,N_1155);
and U6940 (N_6940,N_3772,N_1632);
nor U6941 (N_6941,N_375,N_1730);
or U6942 (N_6942,N_231,N_393);
and U6943 (N_6943,N_2902,N_1931);
or U6944 (N_6944,N_3662,N_919);
nor U6945 (N_6945,N_3816,N_2989);
or U6946 (N_6946,N_2206,N_293);
and U6947 (N_6947,N_3981,N_495);
or U6948 (N_6948,N_403,N_927);
or U6949 (N_6949,N_3442,N_2194);
nor U6950 (N_6950,N_2514,N_1004);
or U6951 (N_6951,N_587,N_2073);
or U6952 (N_6952,N_2445,N_1435);
and U6953 (N_6953,N_1594,N_1598);
nand U6954 (N_6954,N_3788,N_171);
or U6955 (N_6955,N_975,N_3887);
or U6956 (N_6956,N_3896,N_63);
nand U6957 (N_6957,N_3174,N_213);
nand U6958 (N_6958,N_2307,N_880);
nand U6959 (N_6959,N_817,N_1337);
or U6960 (N_6960,N_827,N_2835);
xor U6961 (N_6961,N_1244,N_651);
nand U6962 (N_6962,N_3910,N_2881);
or U6963 (N_6963,N_2166,N_2804);
or U6964 (N_6964,N_2899,N_132);
nand U6965 (N_6965,N_1171,N_2381);
nand U6966 (N_6966,N_1655,N_759);
nor U6967 (N_6967,N_185,N_915);
or U6968 (N_6968,N_2890,N_2705);
and U6969 (N_6969,N_3075,N_3317);
and U6970 (N_6970,N_1985,N_3444);
nand U6971 (N_6971,N_808,N_2416);
or U6972 (N_6972,N_1801,N_3271);
and U6973 (N_6973,N_3825,N_3741);
or U6974 (N_6974,N_3551,N_871);
nand U6975 (N_6975,N_2790,N_1878);
nand U6976 (N_6976,N_3131,N_2244);
xor U6977 (N_6977,N_3477,N_2100);
nor U6978 (N_6978,N_2152,N_576);
nor U6979 (N_6979,N_202,N_3264);
nor U6980 (N_6980,N_283,N_1780);
and U6981 (N_6981,N_3969,N_2646);
or U6982 (N_6982,N_2899,N_3081);
and U6983 (N_6983,N_684,N_2052);
and U6984 (N_6984,N_2769,N_881);
and U6985 (N_6985,N_641,N_2583);
nand U6986 (N_6986,N_700,N_2216);
nor U6987 (N_6987,N_1934,N_2342);
or U6988 (N_6988,N_908,N_3524);
or U6989 (N_6989,N_699,N_2024);
and U6990 (N_6990,N_160,N_2788);
nand U6991 (N_6991,N_1685,N_1738);
nor U6992 (N_6992,N_2460,N_839);
nor U6993 (N_6993,N_2932,N_1871);
nand U6994 (N_6994,N_2492,N_1514);
nor U6995 (N_6995,N_187,N_3125);
or U6996 (N_6996,N_2772,N_1302);
or U6997 (N_6997,N_2744,N_1430);
nor U6998 (N_6998,N_2705,N_3710);
nor U6999 (N_6999,N_2578,N_3339);
nand U7000 (N_7000,N_1720,N_2840);
nor U7001 (N_7001,N_2596,N_2511);
and U7002 (N_7002,N_2430,N_2044);
and U7003 (N_7003,N_1084,N_1252);
nor U7004 (N_7004,N_2426,N_1320);
nand U7005 (N_7005,N_3540,N_2932);
or U7006 (N_7006,N_2275,N_2860);
nand U7007 (N_7007,N_1159,N_310);
nor U7008 (N_7008,N_2388,N_2797);
or U7009 (N_7009,N_2781,N_2566);
or U7010 (N_7010,N_510,N_786);
nor U7011 (N_7011,N_1301,N_2091);
nand U7012 (N_7012,N_217,N_3315);
and U7013 (N_7013,N_1605,N_1648);
nand U7014 (N_7014,N_297,N_3314);
and U7015 (N_7015,N_1564,N_2607);
or U7016 (N_7016,N_2055,N_1416);
or U7017 (N_7017,N_714,N_241);
or U7018 (N_7018,N_2529,N_12);
and U7019 (N_7019,N_3265,N_1054);
and U7020 (N_7020,N_3774,N_1171);
nor U7021 (N_7021,N_2419,N_2860);
nand U7022 (N_7022,N_2553,N_2562);
and U7023 (N_7023,N_3042,N_2669);
or U7024 (N_7024,N_2405,N_1533);
or U7025 (N_7025,N_2774,N_1575);
nand U7026 (N_7026,N_2069,N_2664);
or U7027 (N_7027,N_37,N_62);
or U7028 (N_7028,N_2220,N_3654);
and U7029 (N_7029,N_542,N_1555);
and U7030 (N_7030,N_3279,N_1799);
or U7031 (N_7031,N_2760,N_2987);
or U7032 (N_7032,N_2226,N_460);
and U7033 (N_7033,N_598,N_1363);
nor U7034 (N_7034,N_1514,N_2043);
or U7035 (N_7035,N_3013,N_868);
or U7036 (N_7036,N_1863,N_3687);
nand U7037 (N_7037,N_1067,N_3339);
or U7038 (N_7038,N_417,N_1951);
nand U7039 (N_7039,N_2697,N_3244);
nor U7040 (N_7040,N_3842,N_1534);
nand U7041 (N_7041,N_2554,N_237);
or U7042 (N_7042,N_2269,N_837);
nor U7043 (N_7043,N_1180,N_1862);
or U7044 (N_7044,N_2792,N_2361);
or U7045 (N_7045,N_2591,N_2695);
or U7046 (N_7046,N_1715,N_2304);
nor U7047 (N_7047,N_2014,N_9);
nor U7048 (N_7048,N_1359,N_881);
nor U7049 (N_7049,N_181,N_258);
and U7050 (N_7050,N_2922,N_52);
nand U7051 (N_7051,N_1559,N_1492);
nand U7052 (N_7052,N_2154,N_2044);
and U7053 (N_7053,N_3714,N_2216);
nand U7054 (N_7054,N_736,N_1290);
xor U7055 (N_7055,N_788,N_329);
or U7056 (N_7056,N_1792,N_2629);
or U7057 (N_7057,N_1874,N_2328);
nor U7058 (N_7058,N_3518,N_2907);
nor U7059 (N_7059,N_338,N_1969);
nand U7060 (N_7060,N_71,N_3976);
nand U7061 (N_7061,N_2063,N_549);
and U7062 (N_7062,N_2869,N_2305);
nor U7063 (N_7063,N_1636,N_3026);
nand U7064 (N_7064,N_1625,N_2240);
nand U7065 (N_7065,N_3165,N_644);
and U7066 (N_7066,N_3225,N_1171);
or U7067 (N_7067,N_3211,N_2238);
or U7068 (N_7068,N_2848,N_1039);
or U7069 (N_7069,N_1204,N_342);
nand U7070 (N_7070,N_3533,N_1343);
nor U7071 (N_7071,N_117,N_2792);
nor U7072 (N_7072,N_2355,N_526);
nor U7073 (N_7073,N_1372,N_3255);
nand U7074 (N_7074,N_805,N_2147);
nand U7075 (N_7075,N_1476,N_1359);
nand U7076 (N_7076,N_1537,N_1264);
nand U7077 (N_7077,N_3826,N_1594);
or U7078 (N_7078,N_2619,N_1816);
nand U7079 (N_7079,N_2201,N_2357);
and U7080 (N_7080,N_785,N_1177);
and U7081 (N_7081,N_1098,N_1842);
and U7082 (N_7082,N_1688,N_693);
nor U7083 (N_7083,N_2009,N_632);
and U7084 (N_7084,N_2178,N_2305);
nand U7085 (N_7085,N_1806,N_1576);
and U7086 (N_7086,N_2476,N_3619);
and U7087 (N_7087,N_420,N_636);
nand U7088 (N_7088,N_652,N_3134);
nand U7089 (N_7089,N_2495,N_2676);
nor U7090 (N_7090,N_2368,N_1653);
and U7091 (N_7091,N_2303,N_1877);
and U7092 (N_7092,N_655,N_552);
and U7093 (N_7093,N_3075,N_3387);
nand U7094 (N_7094,N_3769,N_2412);
nor U7095 (N_7095,N_27,N_182);
or U7096 (N_7096,N_1002,N_3750);
and U7097 (N_7097,N_2369,N_2837);
or U7098 (N_7098,N_297,N_758);
nor U7099 (N_7099,N_458,N_2299);
nand U7100 (N_7100,N_360,N_2220);
and U7101 (N_7101,N_3316,N_2710);
nand U7102 (N_7102,N_844,N_3254);
nor U7103 (N_7103,N_677,N_2830);
and U7104 (N_7104,N_2125,N_3856);
or U7105 (N_7105,N_2142,N_3092);
nand U7106 (N_7106,N_1068,N_3598);
or U7107 (N_7107,N_273,N_1715);
nor U7108 (N_7108,N_2059,N_2696);
and U7109 (N_7109,N_346,N_3467);
and U7110 (N_7110,N_3313,N_2381);
or U7111 (N_7111,N_3544,N_669);
nand U7112 (N_7112,N_2269,N_2040);
or U7113 (N_7113,N_894,N_1622);
and U7114 (N_7114,N_82,N_1621);
nor U7115 (N_7115,N_2407,N_107);
or U7116 (N_7116,N_2315,N_123);
and U7117 (N_7117,N_3511,N_1728);
nor U7118 (N_7118,N_784,N_1750);
nand U7119 (N_7119,N_345,N_1582);
xnor U7120 (N_7120,N_2250,N_2298);
or U7121 (N_7121,N_888,N_3532);
and U7122 (N_7122,N_1030,N_279);
nor U7123 (N_7123,N_2042,N_2076);
nand U7124 (N_7124,N_3930,N_190);
nand U7125 (N_7125,N_3382,N_1673);
nor U7126 (N_7126,N_3582,N_1953);
or U7127 (N_7127,N_3545,N_1786);
nand U7128 (N_7128,N_2597,N_1430);
nand U7129 (N_7129,N_116,N_897);
nand U7130 (N_7130,N_3181,N_1695);
nor U7131 (N_7131,N_1106,N_1893);
or U7132 (N_7132,N_2360,N_1188);
or U7133 (N_7133,N_1350,N_3906);
nand U7134 (N_7134,N_1997,N_130);
nand U7135 (N_7135,N_3056,N_1570);
and U7136 (N_7136,N_366,N_1379);
nor U7137 (N_7137,N_1349,N_933);
or U7138 (N_7138,N_2702,N_986);
or U7139 (N_7139,N_2321,N_1938);
nor U7140 (N_7140,N_820,N_1233);
nand U7141 (N_7141,N_379,N_2621);
nand U7142 (N_7142,N_3256,N_3018);
nand U7143 (N_7143,N_3269,N_2912);
nand U7144 (N_7144,N_1540,N_1658);
nand U7145 (N_7145,N_3720,N_3228);
and U7146 (N_7146,N_3949,N_3245);
nor U7147 (N_7147,N_474,N_1972);
and U7148 (N_7148,N_1961,N_2480);
nand U7149 (N_7149,N_2340,N_697);
and U7150 (N_7150,N_3075,N_3158);
nand U7151 (N_7151,N_1784,N_2677);
or U7152 (N_7152,N_2614,N_2512);
nand U7153 (N_7153,N_2365,N_3637);
nand U7154 (N_7154,N_78,N_1059);
and U7155 (N_7155,N_3047,N_1456);
xnor U7156 (N_7156,N_2525,N_1256);
or U7157 (N_7157,N_2331,N_623);
xor U7158 (N_7158,N_1016,N_2354);
or U7159 (N_7159,N_1001,N_3591);
or U7160 (N_7160,N_3826,N_3005);
or U7161 (N_7161,N_2420,N_2761);
nand U7162 (N_7162,N_1975,N_2324);
nand U7163 (N_7163,N_1230,N_1092);
nand U7164 (N_7164,N_1451,N_95);
and U7165 (N_7165,N_3195,N_2820);
nor U7166 (N_7166,N_1415,N_2794);
nand U7167 (N_7167,N_2175,N_3057);
or U7168 (N_7168,N_2336,N_70);
nor U7169 (N_7169,N_2001,N_1719);
nor U7170 (N_7170,N_1407,N_1054);
and U7171 (N_7171,N_2156,N_3088);
nor U7172 (N_7172,N_2533,N_23);
and U7173 (N_7173,N_1347,N_3382);
nor U7174 (N_7174,N_1866,N_2800);
and U7175 (N_7175,N_834,N_2881);
and U7176 (N_7176,N_582,N_408);
and U7177 (N_7177,N_895,N_1705);
nor U7178 (N_7178,N_24,N_204);
and U7179 (N_7179,N_3149,N_2595);
or U7180 (N_7180,N_3953,N_802);
or U7181 (N_7181,N_2830,N_1685);
or U7182 (N_7182,N_1702,N_3352);
nor U7183 (N_7183,N_3896,N_2394);
nor U7184 (N_7184,N_1531,N_3484);
nand U7185 (N_7185,N_5,N_2221);
nor U7186 (N_7186,N_3627,N_1186);
and U7187 (N_7187,N_1588,N_799);
nor U7188 (N_7188,N_300,N_1913);
and U7189 (N_7189,N_1399,N_299);
and U7190 (N_7190,N_2720,N_3777);
nand U7191 (N_7191,N_945,N_1174);
nor U7192 (N_7192,N_1016,N_2365);
or U7193 (N_7193,N_2312,N_1150);
nor U7194 (N_7194,N_1226,N_2008);
nor U7195 (N_7195,N_3047,N_960);
and U7196 (N_7196,N_1688,N_97);
nand U7197 (N_7197,N_1645,N_576);
and U7198 (N_7198,N_737,N_3912);
or U7199 (N_7199,N_3846,N_3761);
and U7200 (N_7200,N_633,N_297);
or U7201 (N_7201,N_867,N_3931);
and U7202 (N_7202,N_2765,N_724);
nand U7203 (N_7203,N_3603,N_2199);
nand U7204 (N_7204,N_2447,N_521);
and U7205 (N_7205,N_2565,N_522);
or U7206 (N_7206,N_2152,N_3393);
nor U7207 (N_7207,N_1327,N_2857);
nand U7208 (N_7208,N_2561,N_441);
or U7209 (N_7209,N_929,N_921);
and U7210 (N_7210,N_2168,N_1538);
nand U7211 (N_7211,N_3044,N_2125);
nor U7212 (N_7212,N_2124,N_1195);
or U7213 (N_7213,N_1011,N_1919);
or U7214 (N_7214,N_2436,N_978);
nand U7215 (N_7215,N_1169,N_253);
nand U7216 (N_7216,N_818,N_3232);
nand U7217 (N_7217,N_3130,N_3410);
or U7218 (N_7218,N_1496,N_709);
nor U7219 (N_7219,N_1406,N_3093);
or U7220 (N_7220,N_801,N_1795);
or U7221 (N_7221,N_3490,N_672);
nand U7222 (N_7222,N_2108,N_1460);
or U7223 (N_7223,N_867,N_106);
nand U7224 (N_7224,N_827,N_588);
or U7225 (N_7225,N_504,N_1972);
or U7226 (N_7226,N_2247,N_3726);
or U7227 (N_7227,N_3967,N_85);
xnor U7228 (N_7228,N_3751,N_2208);
nor U7229 (N_7229,N_566,N_3820);
nand U7230 (N_7230,N_2147,N_3070);
nor U7231 (N_7231,N_264,N_804);
and U7232 (N_7232,N_2382,N_1124);
xor U7233 (N_7233,N_3245,N_2927);
and U7234 (N_7234,N_1128,N_1038);
or U7235 (N_7235,N_1302,N_1426);
and U7236 (N_7236,N_3721,N_3066);
or U7237 (N_7237,N_1665,N_3717);
and U7238 (N_7238,N_1087,N_3308);
nand U7239 (N_7239,N_2103,N_1440);
and U7240 (N_7240,N_3037,N_2422);
and U7241 (N_7241,N_2327,N_1490);
nand U7242 (N_7242,N_1191,N_3302);
or U7243 (N_7243,N_2848,N_2935);
xor U7244 (N_7244,N_3098,N_2204);
nor U7245 (N_7245,N_3514,N_3883);
nor U7246 (N_7246,N_448,N_775);
or U7247 (N_7247,N_616,N_2245);
or U7248 (N_7248,N_1369,N_3348);
nand U7249 (N_7249,N_1792,N_315);
nand U7250 (N_7250,N_3661,N_2355);
and U7251 (N_7251,N_2802,N_2781);
nand U7252 (N_7252,N_617,N_2709);
nor U7253 (N_7253,N_3829,N_3705);
or U7254 (N_7254,N_2599,N_1307);
or U7255 (N_7255,N_1820,N_3406);
xnor U7256 (N_7256,N_1071,N_458);
or U7257 (N_7257,N_3849,N_2957);
nor U7258 (N_7258,N_1908,N_3874);
nor U7259 (N_7259,N_1750,N_2996);
nor U7260 (N_7260,N_1198,N_3324);
or U7261 (N_7261,N_3834,N_262);
and U7262 (N_7262,N_407,N_1288);
and U7263 (N_7263,N_610,N_3587);
and U7264 (N_7264,N_2401,N_1054);
nand U7265 (N_7265,N_350,N_3323);
and U7266 (N_7266,N_2702,N_3656);
or U7267 (N_7267,N_3514,N_2059);
or U7268 (N_7268,N_1605,N_2500);
or U7269 (N_7269,N_346,N_1808);
nand U7270 (N_7270,N_3616,N_1188);
or U7271 (N_7271,N_3505,N_3717);
nor U7272 (N_7272,N_3935,N_285);
nand U7273 (N_7273,N_3995,N_3008);
nand U7274 (N_7274,N_3727,N_2944);
or U7275 (N_7275,N_3798,N_3018);
nand U7276 (N_7276,N_1785,N_3739);
nor U7277 (N_7277,N_17,N_517);
or U7278 (N_7278,N_2760,N_1505);
and U7279 (N_7279,N_823,N_2814);
nand U7280 (N_7280,N_2547,N_1237);
nand U7281 (N_7281,N_1301,N_1203);
nor U7282 (N_7282,N_3576,N_2962);
nand U7283 (N_7283,N_3672,N_143);
or U7284 (N_7284,N_3990,N_2781);
or U7285 (N_7285,N_3052,N_847);
xnor U7286 (N_7286,N_2726,N_1110);
nor U7287 (N_7287,N_731,N_1164);
nand U7288 (N_7288,N_3148,N_3100);
and U7289 (N_7289,N_144,N_3687);
and U7290 (N_7290,N_2298,N_2829);
or U7291 (N_7291,N_2087,N_3947);
or U7292 (N_7292,N_3813,N_565);
nand U7293 (N_7293,N_1346,N_1789);
nor U7294 (N_7294,N_1201,N_251);
nor U7295 (N_7295,N_201,N_209);
and U7296 (N_7296,N_936,N_2781);
nand U7297 (N_7297,N_2189,N_1124);
or U7298 (N_7298,N_3536,N_2591);
and U7299 (N_7299,N_1207,N_2394);
and U7300 (N_7300,N_3998,N_1479);
nor U7301 (N_7301,N_3289,N_1774);
nor U7302 (N_7302,N_1624,N_2518);
or U7303 (N_7303,N_1127,N_2338);
and U7304 (N_7304,N_2981,N_212);
nor U7305 (N_7305,N_3760,N_3843);
or U7306 (N_7306,N_3248,N_414);
and U7307 (N_7307,N_1903,N_2645);
nor U7308 (N_7308,N_2413,N_2242);
or U7309 (N_7309,N_1913,N_2732);
nand U7310 (N_7310,N_1363,N_2438);
nand U7311 (N_7311,N_3303,N_9);
nor U7312 (N_7312,N_1547,N_99);
nor U7313 (N_7313,N_3641,N_1767);
or U7314 (N_7314,N_324,N_3300);
xor U7315 (N_7315,N_873,N_1532);
nor U7316 (N_7316,N_2949,N_2138);
nor U7317 (N_7317,N_119,N_935);
nand U7318 (N_7318,N_856,N_3279);
nand U7319 (N_7319,N_3353,N_1480);
or U7320 (N_7320,N_3904,N_1128);
nand U7321 (N_7321,N_546,N_330);
nor U7322 (N_7322,N_3232,N_3733);
nand U7323 (N_7323,N_785,N_1896);
and U7324 (N_7324,N_2030,N_3397);
nand U7325 (N_7325,N_1177,N_3899);
nand U7326 (N_7326,N_1995,N_2380);
or U7327 (N_7327,N_473,N_1102);
xnor U7328 (N_7328,N_1729,N_1880);
and U7329 (N_7329,N_228,N_3452);
or U7330 (N_7330,N_2958,N_2823);
or U7331 (N_7331,N_3148,N_289);
and U7332 (N_7332,N_1127,N_3259);
and U7333 (N_7333,N_1856,N_2037);
nand U7334 (N_7334,N_601,N_2614);
or U7335 (N_7335,N_2948,N_1798);
or U7336 (N_7336,N_2107,N_3598);
nand U7337 (N_7337,N_3322,N_903);
nor U7338 (N_7338,N_2980,N_3557);
xnor U7339 (N_7339,N_313,N_1663);
nand U7340 (N_7340,N_3401,N_711);
or U7341 (N_7341,N_805,N_2724);
nor U7342 (N_7342,N_3465,N_3561);
or U7343 (N_7343,N_3341,N_381);
nand U7344 (N_7344,N_1108,N_911);
and U7345 (N_7345,N_3,N_1270);
or U7346 (N_7346,N_1891,N_1376);
or U7347 (N_7347,N_346,N_3199);
or U7348 (N_7348,N_1218,N_1839);
or U7349 (N_7349,N_1157,N_350);
or U7350 (N_7350,N_1009,N_2684);
or U7351 (N_7351,N_139,N_2435);
and U7352 (N_7352,N_2176,N_1622);
or U7353 (N_7353,N_747,N_62);
nand U7354 (N_7354,N_2813,N_2071);
or U7355 (N_7355,N_1389,N_636);
nor U7356 (N_7356,N_3646,N_1942);
nor U7357 (N_7357,N_308,N_1810);
nand U7358 (N_7358,N_1838,N_2704);
or U7359 (N_7359,N_1308,N_2774);
or U7360 (N_7360,N_3494,N_1906);
nand U7361 (N_7361,N_2529,N_2057);
nor U7362 (N_7362,N_2703,N_3123);
nand U7363 (N_7363,N_2229,N_2663);
or U7364 (N_7364,N_2133,N_2566);
and U7365 (N_7365,N_2835,N_3998);
nand U7366 (N_7366,N_808,N_2065);
or U7367 (N_7367,N_1223,N_1698);
and U7368 (N_7368,N_1009,N_3588);
and U7369 (N_7369,N_3148,N_871);
nor U7370 (N_7370,N_3627,N_2179);
or U7371 (N_7371,N_3264,N_3753);
or U7372 (N_7372,N_3401,N_3876);
and U7373 (N_7373,N_1907,N_1470);
nand U7374 (N_7374,N_2728,N_2175);
and U7375 (N_7375,N_2766,N_481);
and U7376 (N_7376,N_3359,N_3236);
nand U7377 (N_7377,N_512,N_481);
and U7378 (N_7378,N_1605,N_3959);
nand U7379 (N_7379,N_1142,N_3108);
or U7380 (N_7380,N_1641,N_1962);
or U7381 (N_7381,N_3629,N_3331);
nor U7382 (N_7382,N_1225,N_1085);
or U7383 (N_7383,N_1856,N_3908);
and U7384 (N_7384,N_677,N_2971);
xor U7385 (N_7385,N_333,N_2709);
and U7386 (N_7386,N_701,N_3322);
or U7387 (N_7387,N_3476,N_3798);
and U7388 (N_7388,N_711,N_3045);
or U7389 (N_7389,N_221,N_1001);
nor U7390 (N_7390,N_882,N_3760);
and U7391 (N_7391,N_409,N_2363);
and U7392 (N_7392,N_3652,N_351);
and U7393 (N_7393,N_1385,N_3362);
or U7394 (N_7394,N_479,N_3565);
nand U7395 (N_7395,N_3699,N_964);
and U7396 (N_7396,N_612,N_2418);
nor U7397 (N_7397,N_621,N_3178);
and U7398 (N_7398,N_184,N_2599);
or U7399 (N_7399,N_3367,N_1243);
nor U7400 (N_7400,N_3738,N_2038);
nand U7401 (N_7401,N_3671,N_2428);
or U7402 (N_7402,N_1337,N_3850);
and U7403 (N_7403,N_3920,N_1138);
nor U7404 (N_7404,N_29,N_3439);
nor U7405 (N_7405,N_3316,N_636);
nor U7406 (N_7406,N_2246,N_3298);
and U7407 (N_7407,N_1946,N_406);
or U7408 (N_7408,N_181,N_1803);
or U7409 (N_7409,N_3101,N_2096);
nand U7410 (N_7410,N_3819,N_37);
and U7411 (N_7411,N_329,N_3734);
or U7412 (N_7412,N_3946,N_3282);
or U7413 (N_7413,N_739,N_1980);
or U7414 (N_7414,N_1858,N_2984);
and U7415 (N_7415,N_3210,N_2837);
nor U7416 (N_7416,N_1483,N_2308);
or U7417 (N_7417,N_3491,N_2891);
nand U7418 (N_7418,N_3978,N_1146);
or U7419 (N_7419,N_3958,N_3879);
and U7420 (N_7420,N_1392,N_2004);
nand U7421 (N_7421,N_3490,N_3803);
and U7422 (N_7422,N_3280,N_847);
nand U7423 (N_7423,N_773,N_2834);
nor U7424 (N_7424,N_259,N_3770);
and U7425 (N_7425,N_1002,N_814);
or U7426 (N_7426,N_1516,N_3837);
nor U7427 (N_7427,N_2248,N_3024);
nand U7428 (N_7428,N_3178,N_2721);
nand U7429 (N_7429,N_2238,N_3421);
nor U7430 (N_7430,N_458,N_1894);
and U7431 (N_7431,N_1511,N_3775);
nand U7432 (N_7432,N_3376,N_2632);
nand U7433 (N_7433,N_2813,N_1803);
or U7434 (N_7434,N_1435,N_3382);
or U7435 (N_7435,N_1023,N_1794);
and U7436 (N_7436,N_640,N_2599);
nand U7437 (N_7437,N_53,N_3951);
nand U7438 (N_7438,N_2685,N_3231);
and U7439 (N_7439,N_206,N_1346);
or U7440 (N_7440,N_2166,N_3719);
or U7441 (N_7441,N_2168,N_2207);
nand U7442 (N_7442,N_2958,N_2928);
or U7443 (N_7443,N_2257,N_962);
and U7444 (N_7444,N_2910,N_1610);
nand U7445 (N_7445,N_699,N_386);
nor U7446 (N_7446,N_1908,N_1530);
and U7447 (N_7447,N_2013,N_1624);
and U7448 (N_7448,N_1081,N_3420);
nor U7449 (N_7449,N_3011,N_1161);
or U7450 (N_7450,N_577,N_231);
or U7451 (N_7451,N_1243,N_2403);
and U7452 (N_7452,N_2679,N_2635);
nand U7453 (N_7453,N_2081,N_472);
nand U7454 (N_7454,N_2853,N_3218);
nand U7455 (N_7455,N_3815,N_1567);
or U7456 (N_7456,N_292,N_521);
nand U7457 (N_7457,N_914,N_3402);
nor U7458 (N_7458,N_442,N_2172);
or U7459 (N_7459,N_3615,N_184);
nor U7460 (N_7460,N_1987,N_3862);
and U7461 (N_7461,N_2240,N_2265);
nor U7462 (N_7462,N_638,N_415);
and U7463 (N_7463,N_2456,N_1551);
and U7464 (N_7464,N_3071,N_866);
nand U7465 (N_7465,N_1133,N_68);
and U7466 (N_7466,N_1478,N_2345);
nand U7467 (N_7467,N_3904,N_1709);
nor U7468 (N_7468,N_1077,N_2460);
xor U7469 (N_7469,N_3067,N_3134);
or U7470 (N_7470,N_1918,N_1083);
or U7471 (N_7471,N_387,N_3530);
nand U7472 (N_7472,N_2623,N_1263);
nand U7473 (N_7473,N_3433,N_2666);
nand U7474 (N_7474,N_3195,N_3111);
and U7475 (N_7475,N_1581,N_769);
and U7476 (N_7476,N_2080,N_1885);
or U7477 (N_7477,N_2817,N_2130);
nor U7478 (N_7478,N_404,N_2686);
nand U7479 (N_7479,N_1995,N_3545);
and U7480 (N_7480,N_2450,N_2896);
and U7481 (N_7481,N_1432,N_3883);
and U7482 (N_7482,N_595,N_950);
nand U7483 (N_7483,N_2016,N_835);
nor U7484 (N_7484,N_2537,N_1665);
and U7485 (N_7485,N_331,N_600);
nand U7486 (N_7486,N_3516,N_3057);
and U7487 (N_7487,N_1643,N_1335);
and U7488 (N_7488,N_1852,N_2831);
or U7489 (N_7489,N_2522,N_1833);
nand U7490 (N_7490,N_3318,N_3882);
and U7491 (N_7491,N_2868,N_589);
and U7492 (N_7492,N_528,N_2955);
nand U7493 (N_7493,N_3956,N_3529);
and U7494 (N_7494,N_2256,N_3425);
or U7495 (N_7495,N_3447,N_2228);
nand U7496 (N_7496,N_410,N_2806);
nand U7497 (N_7497,N_3366,N_3879);
or U7498 (N_7498,N_49,N_3441);
and U7499 (N_7499,N_760,N_2468);
xor U7500 (N_7500,N_2259,N_2636);
nor U7501 (N_7501,N_3052,N_1033);
nor U7502 (N_7502,N_883,N_1335);
and U7503 (N_7503,N_229,N_3084);
xor U7504 (N_7504,N_2094,N_3568);
and U7505 (N_7505,N_277,N_1534);
and U7506 (N_7506,N_1993,N_226);
and U7507 (N_7507,N_3880,N_3121);
and U7508 (N_7508,N_92,N_3722);
and U7509 (N_7509,N_1073,N_1854);
nand U7510 (N_7510,N_3468,N_1467);
and U7511 (N_7511,N_41,N_3989);
or U7512 (N_7512,N_1393,N_3069);
nor U7513 (N_7513,N_2266,N_646);
nand U7514 (N_7514,N_3228,N_1723);
or U7515 (N_7515,N_105,N_1193);
nand U7516 (N_7516,N_382,N_2493);
and U7517 (N_7517,N_3346,N_2242);
nand U7518 (N_7518,N_778,N_1672);
and U7519 (N_7519,N_3257,N_590);
nand U7520 (N_7520,N_2238,N_3821);
nand U7521 (N_7521,N_3636,N_1797);
nor U7522 (N_7522,N_1230,N_2846);
or U7523 (N_7523,N_78,N_1674);
nor U7524 (N_7524,N_1179,N_3957);
and U7525 (N_7525,N_2958,N_3291);
and U7526 (N_7526,N_2338,N_2339);
or U7527 (N_7527,N_628,N_115);
and U7528 (N_7528,N_3068,N_2614);
or U7529 (N_7529,N_3989,N_3250);
and U7530 (N_7530,N_2109,N_2740);
nor U7531 (N_7531,N_3492,N_3884);
nor U7532 (N_7532,N_1589,N_2031);
nand U7533 (N_7533,N_1747,N_1340);
nand U7534 (N_7534,N_3993,N_2143);
nor U7535 (N_7535,N_3291,N_2232);
or U7536 (N_7536,N_1190,N_3646);
nor U7537 (N_7537,N_2517,N_989);
nor U7538 (N_7538,N_3212,N_1164);
or U7539 (N_7539,N_3836,N_1365);
nor U7540 (N_7540,N_2034,N_1305);
and U7541 (N_7541,N_116,N_3409);
nand U7542 (N_7542,N_3834,N_3595);
nor U7543 (N_7543,N_1001,N_167);
and U7544 (N_7544,N_3297,N_959);
nand U7545 (N_7545,N_703,N_956);
nor U7546 (N_7546,N_1915,N_3509);
nor U7547 (N_7547,N_592,N_3883);
or U7548 (N_7548,N_2376,N_2932);
and U7549 (N_7549,N_960,N_3787);
nor U7550 (N_7550,N_2367,N_3431);
nor U7551 (N_7551,N_2840,N_2567);
nand U7552 (N_7552,N_2538,N_1588);
or U7553 (N_7553,N_2126,N_3941);
and U7554 (N_7554,N_1792,N_121);
and U7555 (N_7555,N_630,N_23);
nor U7556 (N_7556,N_3523,N_3051);
nand U7557 (N_7557,N_261,N_1387);
nand U7558 (N_7558,N_3222,N_572);
and U7559 (N_7559,N_3787,N_1649);
nor U7560 (N_7560,N_1129,N_1917);
or U7561 (N_7561,N_949,N_3605);
or U7562 (N_7562,N_249,N_3371);
nand U7563 (N_7563,N_1263,N_786);
and U7564 (N_7564,N_1056,N_2908);
or U7565 (N_7565,N_3782,N_2369);
nor U7566 (N_7566,N_2067,N_1075);
nand U7567 (N_7567,N_1523,N_2519);
nor U7568 (N_7568,N_2965,N_1488);
or U7569 (N_7569,N_457,N_15);
nand U7570 (N_7570,N_2826,N_1962);
nor U7571 (N_7571,N_2133,N_1081);
and U7572 (N_7572,N_3579,N_428);
nand U7573 (N_7573,N_1924,N_2855);
nor U7574 (N_7574,N_664,N_2108);
and U7575 (N_7575,N_1585,N_1856);
nor U7576 (N_7576,N_259,N_2561);
and U7577 (N_7577,N_1357,N_3385);
nand U7578 (N_7578,N_757,N_930);
nand U7579 (N_7579,N_437,N_3470);
or U7580 (N_7580,N_1689,N_497);
nand U7581 (N_7581,N_638,N_1250);
and U7582 (N_7582,N_2964,N_2768);
and U7583 (N_7583,N_1613,N_1664);
nand U7584 (N_7584,N_2986,N_1195);
xnor U7585 (N_7585,N_1908,N_670);
and U7586 (N_7586,N_1267,N_2313);
xnor U7587 (N_7587,N_2512,N_1243);
nor U7588 (N_7588,N_1616,N_3105);
and U7589 (N_7589,N_524,N_79);
nand U7590 (N_7590,N_2520,N_227);
nor U7591 (N_7591,N_522,N_3283);
and U7592 (N_7592,N_2296,N_874);
and U7593 (N_7593,N_3542,N_361);
nor U7594 (N_7594,N_1909,N_3946);
and U7595 (N_7595,N_2612,N_507);
nor U7596 (N_7596,N_1609,N_3504);
nand U7597 (N_7597,N_280,N_2887);
or U7598 (N_7598,N_464,N_1739);
or U7599 (N_7599,N_725,N_1482);
or U7600 (N_7600,N_2782,N_2950);
nor U7601 (N_7601,N_3347,N_447);
and U7602 (N_7602,N_1764,N_754);
or U7603 (N_7603,N_171,N_2523);
and U7604 (N_7604,N_2329,N_2914);
or U7605 (N_7605,N_3646,N_1304);
or U7606 (N_7606,N_2764,N_2839);
nand U7607 (N_7607,N_212,N_2879);
nor U7608 (N_7608,N_3858,N_1491);
nor U7609 (N_7609,N_2853,N_3235);
nand U7610 (N_7610,N_303,N_698);
nand U7611 (N_7611,N_1911,N_3312);
or U7612 (N_7612,N_678,N_3851);
nor U7613 (N_7613,N_432,N_388);
and U7614 (N_7614,N_1452,N_1942);
nor U7615 (N_7615,N_769,N_674);
nor U7616 (N_7616,N_1656,N_1382);
nand U7617 (N_7617,N_2794,N_495);
or U7618 (N_7618,N_1409,N_489);
nor U7619 (N_7619,N_2491,N_1204);
nor U7620 (N_7620,N_1504,N_2528);
nand U7621 (N_7621,N_3486,N_848);
or U7622 (N_7622,N_1596,N_1483);
and U7623 (N_7623,N_3625,N_2275);
nand U7624 (N_7624,N_3410,N_2444);
nor U7625 (N_7625,N_3112,N_1040);
nor U7626 (N_7626,N_3404,N_3905);
or U7627 (N_7627,N_1350,N_1879);
nand U7628 (N_7628,N_427,N_2349);
and U7629 (N_7629,N_1352,N_1131);
and U7630 (N_7630,N_1070,N_2378);
and U7631 (N_7631,N_2612,N_617);
nand U7632 (N_7632,N_2282,N_1502);
nand U7633 (N_7633,N_189,N_1806);
nor U7634 (N_7634,N_2415,N_3331);
and U7635 (N_7635,N_3879,N_1484);
nor U7636 (N_7636,N_2081,N_2897);
nand U7637 (N_7637,N_1473,N_3790);
nor U7638 (N_7638,N_3725,N_1871);
or U7639 (N_7639,N_1835,N_2170);
nand U7640 (N_7640,N_205,N_2464);
and U7641 (N_7641,N_376,N_3824);
or U7642 (N_7642,N_3912,N_3981);
and U7643 (N_7643,N_2576,N_2649);
nor U7644 (N_7644,N_3985,N_3728);
and U7645 (N_7645,N_2518,N_3851);
nand U7646 (N_7646,N_1110,N_3507);
nor U7647 (N_7647,N_2188,N_1807);
nand U7648 (N_7648,N_1656,N_84);
nor U7649 (N_7649,N_3461,N_1786);
and U7650 (N_7650,N_1382,N_3949);
nor U7651 (N_7651,N_911,N_2159);
and U7652 (N_7652,N_2692,N_3463);
nor U7653 (N_7653,N_3336,N_2616);
nor U7654 (N_7654,N_932,N_605);
or U7655 (N_7655,N_1326,N_326);
or U7656 (N_7656,N_1036,N_412);
and U7657 (N_7657,N_2092,N_1038);
and U7658 (N_7658,N_2331,N_794);
nor U7659 (N_7659,N_3568,N_2813);
or U7660 (N_7660,N_1911,N_2227);
and U7661 (N_7661,N_1631,N_1523);
nand U7662 (N_7662,N_1406,N_3466);
and U7663 (N_7663,N_1281,N_3607);
nor U7664 (N_7664,N_988,N_164);
or U7665 (N_7665,N_207,N_3004);
or U7666 (N_7666,N_1871,N_1837);
nand U7667 (N_7667,N_1882,N_2917);
or U7668 (N_7668,N_3290,N_2015);
nand U7669 (N_7669,N_614,N_2809);
nand U7670 (N_7670,N_3510,N_1191);
nor U7671 (N_7671,N_2873,N_13);
nand U7672 (N_7672,N_3021,N_688);
nand U7673 (N_7673,N_2651,N_65);
nand U7674 (N_7674,N_3411,N_3294);
xnor U7675 (N_7675,N_1107,N_1506);
nor U7676 (N_7676,N_3193,N_3960);
nand U7677 (N_7677,N_3439,N_2725);
nor U7678 (N_7678,N_74,N_966);
xor U7679 (N_7679,N_793,N_3007);
or U7680 (N_7680,N_1532,N_1370);
or U7681 (N_7681,N_2515,N_990);
nand U7682 (N_7682,N_3276,N_2238);
nor U7683 (N_7683,N_3707,N_3386);
nand U7684 (N_7684,N_3447,N_1142);
and U7685 (N_7685,N_756,N_1045);
or U7686 (N_7686,N_3298,N_3730);
and U7687 (N_7687,N_1764,N_1726);
nand U7688 (N_7688,N_2774,N_3571);
nand U7689 (N_7689,N_3743,N_3108);
nor U7690 (N_7690,N_292,N_2399);
nand U7691 (N_7691,N_911,N_1617);
or U7692 (N_7692,N_1894,N_1588);
nand U7693 (N_7693,N_29,N_1110);
nand U7694 (N_7694,N_3669,N_1203);
or U7695 (N_7695,N_2015,N_498);
and U7696 (N_7696,N_3742,N_511);
and U7697 (N_7697,N_2575,N_3847);
nor U7698 (N_7698,N_3795,N_2162);
and U7699 (N_7699,N_3793,N_3774);
nand U7700 (N_7700,N_80,N_1953);
nand U7701 (N_7701,N_772,N_1338);
nand U7702 (N_7702,N_842,N_525);
nor U7703 (N_7703,N_3265,N_3862);
nor U7704 (N_7704,N_2812,N_418);
nand U7705 (N_7705,N_1293,N_2707);
nand U7706 (N_7706,N_1683,N_1889);
or U7707 (N_7707,N_767,N_366);
or U7708 (N_7708,N_1688,N_590);
and U7709 (N_7709,N_1829,N_1462);
nand U7710 (N_7710,N_1552,N_10);
nand U7711 (N_7711,N_627,N_3863);
nand U7712 (N_7712,N_721,N_151);
or U7713 (N_7713,N_2792,N_1292);
or U7714 (N_7714,N_1859,N_3629);
and U7715 (N_7715,N_717,N_1436);
nor U7716 (N_7716,N_640,N_958);
nor U7717 (N_7717,N_2375,N_3559);
or U7718 (N_7718,N_1637,N_575);
or U7719 (N_7719,N_3082,N_3612);
and U7720 (N_7720,N_3137,N_360);
and U7721 (N_7721,N_140,N_2338);
and U7722 (N_7722,N_1943,N_1872);
or U7723 (N_7723,N_1729,N_1383);
or U7724 (N_7724,N_2977,N_3901);
or U7725 (N_7725,N_3239,N_337);
or U7726 (N_7726,N_1644,N_3355);
and U7727 (N_7727,N_1219,N_1216);
nand U7728 (N_7728,N_3583,N_659);
and U7729 (N_7729,N_3129,N_3500);
and U7730 (N_7730,N_1568,N_756);
and U7731 (N_7731,N_375,N_2443);
nand U7732 (N_7732,N_1392,N_1671);
and U7733 (N_7733,N_1220,N_1675);
or U7734 (N_7734,N_1983,N_2074);
nor U7735 (N_7735,N_329,N_120);
nor U7736 (N_7736,N_712,N_1410);
nor U7737 (N_7737,N_3923,N_3799);
nor U7738 (N_7738,N_2550,N_277);
nand U7739 (N_7739,N_1490,N_1335);
nor U7740 (N_7740,N_2209,N_2009);
nor U7741 (N_7741,N_3372,N_2696);
nor U7742 (N_7742,N_2759,N_1038);
nand U7743 (N_7743,N_1509,N_3257);
nand U7744 (N_7744,N_2816,N_1647);
or U7745 (N_7745,N_3757,N_800);
and U7746 (N_7746,N_1690,N_1218);
nand U7747 (N_7747,N_3328,N_3155);
nor U7748 (N_7748,N_2799,N_2943);
nand U7749 (N_7749,N_3948,N_3571);
nor U7750 (N_7750,N_2861,N_3050);
or U7751 (N_7751,N_1774,N_2048);
or U7752 (N_7752,N_44,N_2121);
nor U7753 (N_7753,N_3225,N_125);
and U7754 (N_7754,N_3431,N_635);
or U7755 (N_7755,N_2566,N_621);
nand U7756 (N_7756,N_332,N_459);
nor U7757 (N_7757,N_1511,N_418);
nand U7758 (N_7758,N_1738,N_2487);
or U7759 (N_7759,N_1895,N_713);
and U7760 (N_7760,N_2199,N_764);
and U7761 (N_7761,N_1686,N_3000);
or U7762 (N_7762,N_2522,N_2627);
nand U7763 (N_7763,N_575,N_1859);
nand U7764 (N_7764,N_1456,N_1981);
and U7765 (N_7765,N_1944,N_1540);
or U7766 (N_7766,N_221,N_3713);
nor U7767 (N_7767,N_123,N_3966);
and U7768 (N_7768,N_2167,N_615);
and U7769 (N_7769,N_510,N_3267);
or U7770 (N_7770,N_1263,N_2201);
or U7771 (N_7771,N_11,N_3136);
nand U7772 (N_7772,N_1475,N_171);
nor U7773 (N_7773,N_1894,N_2368);
or U7774 (N_7774,N_2645,N_3568);
nor U7775 (N_7775,N_3002,N_2204);
and U7776 (N_7776,N_2501,N_640);
and U7777 (N_7777,N_2578,N_455);
nand U7778 (N_7778,N_782,N_2346);
or U7779 (N_7779,N_2329,N_2946);
and U7780 (N_7780,N_2021,N_1726);
nand U7781 (N_7781,N_1722,N_2886);
and U7782 (N_7782,N_2434,N_2800);
or U7783 (N_7783,N_2526,N_1236);
nand U7784 (N_7784,N_2660,N_2574);
and U7785 (N_7785,N_1459,N_2937);
or U7786 (N_7786,N_3232,N_1537);
nand U7787 (N_7787,N_492,N_3603);
and U7788 (N_7788,N_562,N_3078);
nand U7789 (N_7789,N_2638,N_2744);
nand U7790 (N_7790,N_1280,N_2436);
or U7791 (N_7791,N_2558,N_1036);
nor U7792 (N_7792,N_235,N_3600);
nor U7793 (N_7793,N_1337,N_1526);
or U7794 (N_7794,N_1234,N_452);
or U7795 (N_7795,N_3171,N_3227);
and U7796 (N_7796,N_10,N_2641);
nand U7797 (N_7797,N_1161,N_3888);
nand U7798 (N_7798,N_2256,N_464);
nor U7799 (N_7799,N_580,N_2535);
nor U7800 (N_7800,N_2385,N_3321);
and U7801 (N_7801,N_1925,N_3227);
nor U7802 (N_7802,N_292,N_3161);
nor U7803 (N_7803,N_2328,N_2217);
or U7804 (N_7804,N_1693,N_2283);
and U7805 (N_7805,N_3399,N_457);
and U7806 (N_7806,N_1231,N_2950);
nor U7807 (N_7807,N_2796,N_3784);
and U7808 (N_7808,N_1102,N_58);
or U7809 (N_7809,N_3096,N_379);
nand U7810 (N_7810,N_1807,N_2453);
or U7811 (N_7811,N_3694,N_3062);
nor U7812 (N_7812,N_2735,N_1118);
nor U7813 (N_7813,N_3691,N_2465);
and U7814 (N_7814,N_734,N_946);
or U7815 (N_7815,N_611,N_2795);
nor U7816 (N_7816,N_3089,N_627);
nand U7817 (N_7817,N_2539,N_663);
nand U7818 (N_7818,N_3001,N_3142);
nand U7819 (N_7819,N_3965,N_3574);
nor U7820 (N_7820,N_2775,N_1324);
nand U7821 (N_7821,N_3621,N_2556);
nand U7822 (N_7822,N_2082,N_1366);
or U7823 (N_7823,N_2242,N_394);
nand U7824 (N_7824,N_2861,N_58);
nor U7825 (N_7825,N_2473,N_1238);
nand U7826 (N_7826,N_137,N_645);
nand U7827 (N_7827,N_3761,N_250);
nor U7828 (N_7828,N_3136,N_2688);
nor U7829 (N_7829,N_1550,N_1699);
and U7830 (N_7830,N_2234,N_1471);
or U7831 (N_7831,N_594,N_188);
or U7832 (N_7832,N_3214,N_2455);
nor U7833 (N_7833,N_3862,N_624);
or U7834 (N_7834,N_2720,N_2841);
nor U7835 (N_7835,N_232,N_526);
nand U7836 (N_7836,N_241,N_1237);
nor U7837 (N_7837,N_2976,N_2432);
or U7838 (N_7838,N_707,N_3870);
nor U7839 (N_7839,N_2168,N_370);
and U7840 (N_7840,N_3822,N_181);
nand U7841 (N_7841,N_848,N_1853);
xor U7842 (N_7842,N_2640,N_1462);
or U7843 (N_7843,N_908,N_3637);
nand U7844 (N_7844,N_2904,N_749);
nor U7845 (N_7845,N_1254,N_1515);
nand U7846 (N_7846,N_1026,N_163);
and U7847 (N_7847,N_1396,N_3031);
or U7848 (N_7848,N_815,N_2603);
nand U7849 (N_7849,N_3772,N_3102);
nand U7850 (N_7850,N_3944,N_3042);
and U7851 (N_7851,N_3530,N_634);
and U7852 (N_7852,N_3034,N_282);
or U7853 (N_7853,N_1116,N_576);
or U7854 (N_7854,N_3735,N_353);
nand U7855 (N_7855,N_3941,N_3933);
or U7856 (N_7856,N_119,N_2941);
and U7857 (N_7857,N_991,N_3925);
or U7858 (N_7858,N_310,N_132);
or U7859 (N_7859,N_3646,N_2631);
and U7860 (N_7860,N_819,N_2231);
nand U7861 (N_7861,N_1578,N_1369);
and U7862 (N_7862,N_3277,N_126);
or U7863 (N_7863,N_3010,N_3187);
nor U7864 (N_7864,N_3276,N_1390);
nor U7865 (N_7865,N_2811,N_2758);
nand U7866 (N_7866,N_2763,N_2489);
xnor U7867 (N_7867,N_3272,N_43);
nand U7868 (N_7868,N_2537,N_3798);
or U7869 (N_7869,N_3254,N_3223);
or U7870 (N_7870,N_2733,N_2601);
and U7871 (N_7871,N_1574,N_196);
and U7872 (N_7872,N_3266,N_1791);
nor U7873 (N_7873,N_2563,N_849);
nand U7874 (N_7874,N_1060,N_433);
nand U7875 (N_7875,N_3939,N_592);
nand U7876 (N_7876,N_3895,N_2178);
xor U7877 (N_7877,N_1347,N_3747);
or U7878 (N_7878,N_958,N_1843);
or U7879 (N_7879,N_1663,N_1096);
and U7880 (N_7880,N_1511,N_2321);
and U7881 (N_7881,N_851,N_841);
nor U7882 (N_7882,N_1076,N_1384);
and U7883 (N_7883,N_2387,N_2283);
or U7884 (N_7884,N_522,N_2363);
nor U7885 (N_7885,N_2364,N_1825);
or U7886 (N_7886,N_1349,N_2284);
or U7887 (N_7887,N_165,N_2955);
or U7888 (N_7888,N_3671,N_3963);
nand U7889 (N_7889,N_185,N_2489);
and U7890 (N_7890,N_726,N_1675);
nand U7891 (N_7891,N_3282,N_3018);
nand U7892 (N_7892,N_909,N_281);
or U7893 (N_7893,N_3064,N_1058);
and U7894 (N_7894,N_625,N_1984);
nor U7895 (N_7895,N_2190,N_3335);
and U7896 (N_7896,N_1769,N_3456);
nor U7897 (N_7897,N_2196,N_191);
nor U7898 (N_7898,N_3635,N_943);
or U7899 (N_7899,N_1627,N_273);
and U7900 (N_7900,N_3145,N_1464);
nand U7901 (N_7901,N_775,N_3715);
or U7902 (N_7902,N_1905,N_1666);
nor U7903 (N_7903,N_536,N_3035);
and U7904 (N_7904,N_795,N_3845);
or U7905 (N_7905,N_1930,N_3685);
or U7906 (N_7906,N_2744,N_3678);
xnor U7907 (N_7907,N_3081,N_717);
or U7908 (N_7908,N_3573,N_2175);
and U7909 (N_7909,N_2877,N_2438);
nor U7910 (N_7910,N_572,N_1312);
or U7911 (N_7911,N_3863,N_2347);
nor U7912 (N_7912,N_3677,N_813);
nor U7913 (N_7913,N_1136,N_3687);
nand U7914 (N_7914,N_1855,N_194);
and U7915 (N_7915,N_3830,N_166);
and U7916 (N_7916,N_1718,N_3393);
nor U7917 (N_7917,N_3921,N_1176);
and U7918 (N_7918,N_771,N_3712);
or U7919 (N_7919,N_3974,N_3581);
or U7920 (N_7920,N_3051,N_1840);
or U7921 (N_7921,N_3708,N_2328);
xor U7922 (N_7922,N_2357,N_435);
and U7923 (N_7923,N_852,N_1579);
or U7924 (N_7924,N_3030,N_3415);
nand U7925 (N_7925,N_992,N_1651);
and U7926 (N_7926,N_3951,N_1602);
nand U7927 (N_7927,N_3486,N_3968);
nand U7928 (N_7928,N_1419,N_1124);
or U7929 (N_7929,N_119,N_2949);
nand U7930 (N_7930,N_154,N_281);
and U7931 (N_7931,N_3490,N_2876);
nor U7932 (N_7932,N_2533,N_728);
nand U7933 (N_7933,N_684,N_3500);
and U7934 (N_7934,N_2363,N_1174);
or U7935 (N_7935,N_1784,N_290);
nand U7936 (N_7936,N_3635,N_3544);
nand U7937 (N_7937,N_2026,N_1279);
or U7938 (N_7938,N_2088,N_2777);
nand U7939 (N_7939,N_3440,N_1286);
or U7940 (N_7940,N_2622,N_2672);
and U7941 (N_7941,N_1807,N_1635);
nand U7942 (N_7942,N_2926,N_2413);
nand U7943 (N_7943,N_3342,N_2963);
nand U7944 (N_7944,N_1663,N_2015);
or U7945 (N_7945,N_3201,N_3815);
nor U7946 (N_7946,N_3855,N_1351);
or U7947 (N_7947,N_3341,N_146);
nor U7948 (N_7948,N_3552,N_3251);
or U7949 (N_7949,N_2003,N_870);
or U7950 (N_7950,N_3331,N_3119);
nand U7951 (N_7951,N_2217,N_176);
or U7952 (N_7952,N_3902,N_3804);
nand U7953 (N_7953,N_851,N_328);
nor U7954 (N_7954,N_3554,N_2642);
or U7955 (N_7955,N_481,N_165);
and U7956 (N_7956,N_1202,N_1239);
or U7957 (N_7957,N_512,N_1553);
nand U7958 (N_7958,N_1534,N_1163);
or U7959 (N_7959,N_584,N_1925);
nand U7960 (N_7960,N_1508,N_3867);
nor U7961 (N_7961,N_643,N_1097);
and U7962 (N_7962,N_371,N_1127);
and U7963 (N_7963,N_3218,N_2068);
nor U7964 (N_7964,N_1221,N_2354);
or U7965 (N_7965,N_654,N_840);
and U7966 (N_7966,N_3159,N_422);
nand U7967 (N_7967,N_3250,N_3678);
nand U7968 (N_7968,N_1203,N_79);
nand U7969 (N_7969,N_2545,N_2919);
nand U7970 (N_7970,N_1548,N_2476);
nand U7971 (N_7971,N_2015,N_1834);
nand U7972 (N_7972,N_419,N_2780);
nor U7973 (N_7973,N_3386,N_3118);
xnor U7974 (N_7974,N_2,N_948);
or U7975 (N_7975,N_2386,N_2212);
and U7976 (N_7976,N_1774,N_1869);
nor U7977 (N_7977,N_137,N_3189);
nand U7978 (N_7978,N_1090,N_236);
and U7979 (N_7979,N_3298,N_1243);
nand U7980 (N_7980,N_3973,N_1156);
nand U7981 (N_7981,N_3736,N_901);
or U7982 (N_7982,N_513,N_1811);
or U7983 (N_7983,N_1371,N_1572);
xor U7984 (N_7984,N_1136,N_299);
nand U7985 (N_7985,N_2897,N_3100);
xor U7986 (N_7986,N_417,N_2186);
nand U7987 (N_7987,N_2475,N_308);
nor U7988 (N_7988,N_403,N_1219);
or U7989 (N_7989,N_1044,N_640);
or U7990 (N_7990,N_2120,N_3013);
and U7991 (N_7991,N_2403,N_1904);
nor U7992 (N_7992,N_536,N_1141);
nor U7993 (N_7993,N_3953,N_1325);
and U7994 (N_7994,N_3943,N_1273);
nand U7995 (N_7995,N_2341,N_3645);
and U7996 (N_7996,N_1557,N_3983);
nand U7997 (N_7997,N_2314,N_3007);
nor U7998 (N_7998,N_3221,N_1289);
nor U7999 (N_7999,N_429,N_807);
and U8000 (N_8000,N_6977,N_4365);
nor U8001 (N_8001,N_6546,N_5343);
xor U8002 (N_8002,N_4481,N_4716);
nand U8003 (N_8003,N_6012,N_6614);
nor U8004 (N_8004,N_6602,N_5612);
nor U8005 (N_8005,N_4047,N_4097);
nor U8006 (N_8006,N_5147,N_5222);
nor U8007 (N_8007,N_5620,N_4052);
nand U8008 (N_8008,N_5616,N_4703);
and U8009 (N_8009,N_6383,N_4066);
nand U8010 (N_8010,N_4137,N_4876);
xnor U8011 (N_8011,N_7888,N_4962);
and U8012 (N_8012,N_6644,N_7398);
and U8013 (N_8013,N_6010,N_7996);
or U8014 (N_8014,N_7341,N_5779);
or U8015 (N_8015,N_5424,N_5210);
and U8016 (N_8016,N_6405,N_7503);
nor U8017 (N_8017,N_7671,N_7316);
nand U8018 (N_8018,N_7758,N_7878);
and U8019 (N_8019,N_4808,N_5171);
nand U8020 (N_8020,N_5765,N_5964);
or U8021 (N_8021,N_4651,N_6757);
and U8022 (N_8022,N_7274,N_4616);
nor U8023 (N_8023,N_7505,N_5339);
or U8024 (N_8024,N_6563,N_4114);
or U8025 (N_8025,N_7824,N_7013);
nor U8026 (N_8026,N_6776,N_7492);
or U8027 (N_8027,N_6105,N_6719);
or U8028 (N_8028,N_6975,N_5662);
or U8029 (N_8029,N_4514,N_5911);
nand U8030 (N_8030,N_7283,N_6525);
or U8031 (N_8031,N_4430,N_5609);
or U8032 (N_8032,N_4099,N_4232);
or U8033 (N_8033,N_7899,N_4136);
or U8034 (N_8034,N_4402,N_4834);
or U8035 (N_8035,N_5017,N_7884);
nor U8036 (N_8036,N_6324,N_5512);
nor U8037 (N_8037,N_5149,N_5225);
or U8038 (N_8038,N_4112,N_5992);
and U8039 (N_8039,N_6223,N_4253);
and U8040 (N_8040,N_4625,N_5728);
nor U8041 (N_8041,N_6378,N_7975);
or U8042 (N_8042,N_4568,N_6842);
and U8043 (N_8043,N_6565,N_7006);
xnor U8044 (N_8044,N_4918,N_5414);
and U8045 (N_8045,N_7711,N_4060);
nand U8046 (N_8046,N_4351,N_5570);
or U8047 (N_8047,N_5094,N_7998);
nand U8048 (N_8048,N_6856,N_6081);
nand U8049 (N_8049,N_7203,N_7208);
nor U8050 (N_8050,N_7488,N_5143);
or U8051 (N_8051,N_6964,N_4658);
and U8052 (N_8052,N_4222,N_4970);
nor U8053 (N_8053,N_5279,N_6168);
nor U8054 (N_8054,N_4171,N_6976);
and U8055 (N_8055,N_7877,N_4030);
or U8056 (N_8056,N_7388,N_7469);
nand U8057 (N_8057,N_7734,N_4815);
and U8058 (N_8058,N_7618,N_4337);
and U8059 (N_8059,N_4077,N_7875);
and U8060 (N_8060,N_6543,N_6103);
and U8061 (N_8061,N_5234,N_4446);
nor U8062 (N_8062,N_7217,N_4290);
nor U8063 (N_8063,N_4592,N_4374);
nand U8064 (N_8064,N_4497,N_4566);
and U8065 (N_8065,N_7893,N_7150);
or U8066 (N_8066,N_5795,N_5580);
nand U8067 (N_8067,N_6998,N_5514);
nor U8068 (N_8068,N_5075,N_4118);
nor U8069 (N_8069,N_4740,N_7243);
nor U8070 (N_8070,N_4323,N_5454);
and U8071 (N_8071,N_6247,N_4184);
nand U8072 (N_8072,N_6309,N_5833);
nor U8073 (N_8073,N_7856,N_4668);
or U8074 (N_8074,N_5655,N_6731);
or U8075 (N_8075,N_5719,N_6456);
nor U8076 (N_8076,N_5398,N_5155);
nand U8077 (N_8077,N_7801,N_6888);
and U8078 (N_8078,N_6735,N_7206);
or U8079 (N_8079,N_7119,N_5578);
or U8080 (N_8080,N_7154,N_4547);
nor U8081 (N_8081,N_6067,N_4724);
and U8082 (N_8082,N_5531,N_4513);
nor U8083 (N_8083,N_7866,N_4665);
xor U8084 (N_8084,N_7832,N_4996);
nor U8085 (N_8085,N_5688,N_7481);
nand U8086 (N_8086,N_6285,N_5749);
nand U8087 (N_8087,N_6327,N_5340);
or U8088 (N_8088,N_6689,N_5634);
nand U8089 (N_8089,N_5261,N_4604);
nand U8090 (N_8090,N_7635,N_5389);
or U8091 (N_8091,N_4781,N_4937);
nand U8092 (N_8092,N_7923,N_6155);
nand U8093 (N_8093,N_4154,N_6165);
and U8094 (N_8094,N_7743,N_4847);
or U8095 (N_8095,N_7068,N_4960);
and U8096 (N_8096,N_6000,N_5381);
nand U8097 (N_8097,N_7615,N_7708);
or U8098 (N_8098,N_6225,N_5484);
and U8099 (N_8099,N_7805,N_4257);
or U8100 (N_8100,N_5955,N_5456);
and U8101 (N_8101,N_6711,N_5378);
and U8102 (N_8102,N_5518,N_7415);
and U8103 (N_8103,N_4848,N_5027);
or U8104 (N_8104,N_6679,N_5581);
and U8105 (N_8105,N_6462,N_5387);
and U8106 (N_8106,N_4428,N_5707);
nor U8107 (N_8107,N_6003,N_7352);
nand U8108 (N_8108,N_5879,N_4585);
or U8109 (N_8109,N_5376,N_7261);
and U8110 (N_8110,N_5540,N_5863);
or U8111 (N_8111,N_7192,N_7683);
and U8112 (N_8112,N_5851,N_6379);
nor U8113 (N_8113,N_7187,N_5917);
nand U8114 (N_8114,N_4571,N_6001);
and U8115 (N_8115,N_7370,N_7616);
and U8116 (N_8116,N_4537,N_5295);
and U8117 (N_8117,N_7174,N_7291);
and U8118 (N_8118,N_4810,N_5706);
nor U8119 (N_8119,N_7416,N_5517);
nand U8120 (N_8120,N_7531,N_4559);
nand U8121 (N_8121,N_7762,N_6006);
and U8122 (N_8122,N_4051,N_6049);
nand U8123 (N_8123,N_7788,N_6903);
nand U8124 (N_8124,N_5754,N_7599);
or U8125 (N_8125,N_7993,N_4973);
and U8126 (N_8126,N_7922,N_4965);
and U8127 (N_8127,N_5941,N_5011);
nand U8128 (N_8128,N_6276,N_7081);
nand U8129 (N_8129,N_5752,N_6152);
or U8130 (N_8130,N_7581,N_7628);
and U8131 (N_8131,N_5912,N_7949);
nor U8132 (N_8132,N_4587,N_7904);
nand U8133 (N_8133,N_5346,N_6552);
nor U8134 (N_8134,N_4684,N_7770);
and U8135 (N_8135,N_5298,N_7980);
and U8136 (N_8136,N_5862,N_5588);
nand U8137 (N_8137,N_4264,N_5076);
nor U8138 (N_8138,N_4491,N_7061);
and U8139 (N_8139,N_4338,N_4227);
nand U8140 (N_8140,N_7432,N_6827);
or U8141 (N_8141,N_7631,N_6040);
nand U8142 (N_8142,N_5335,N_6085);
and U8143 (N_8143,N_5247,N_4265);
nor U8144 (N_8144,N_4818,N_6897);
nor U8145 (N_8145,N_7300,N_6253);
nand U8146 (N_8146,N_4316,N_6920);
nand U8147 (N_8147,N_7556,N_6883);
nor U8148 (N_8148,N_4450,N_7759);
or U8149 (N_8149,N_5781,N_5922);
nand U8150 (N_8150,N_4336,N_4427);
and U8151 (N_8151,N_5152,N_6516);
nor U8152 (N_8152,N_7059,N_6541);
or U8153 (N_8153,N_7016,N_4468);
nor U8154 (N_8154,N_7236,N_7390);
xnor U8155 (N_8155,N_6186,N_6385);
nor U8156 (N_8156,N_7771,N_4618);
nor U8157 (N_8157,N_7333,N_5939);
and U8158 (N_8158,N_7664,N_7799);
and U8159 (N_8159,N_6956,N_7368);
nor U8160 (N_8160,N_7158,N_6609);
or U8161 (N_8161,N_4378,N_4441);
nand U8162 (N_8162,N_4649,N_4675);
nand U8163 (N_8163,N_5057,N_5640);
or U8164 (N_8164,N_5235,N_4659);
or U8165 (N_8165,N_4904,N_4076);
or U8166 (N_8166,N_5552,N_7041);
nor U8167 (N_8167,N_6039,N_4555);
or U8168 (N_8168,N_7858,N_7905);
or U8169 (N_8169,N_5994,N_5743);
nand U8170 (N_8170,N_4729,N_4622);
nor U8171 (N_8171,N_7662,N_7427);
nand U8172 (N_8172,N_4536,N_4170);
and U8173 (N_8173,N_6620,N_4862);
nand U8174 (N_8174,N_6863,N_4237);
xor U8175 (N_8175,N_7062,N_5563);
or U8176 (N_8176,N_6844,N_5052);
and U8177 (N_8177,N_7789,N_5604);
or U8178 (N_8178,N_7241,N_4967);
nand U8179 (N_8179,N_6498,N_7981);
and U8180 (N_8180,N_4643,N_4899);
and U8181 (N_8181,N_7324,N_4755);
nand U8182 (N_8182,N_4550,N_4499);
and U8183 (N_8183,N_6292,N_4433);
and U8184 (N_8184,N_4489,N_6058);
nand U8185 (N_8185,N_5538,N_6947);
and U8186 (N_8186,N_6053,N_4844);
and U8187 (N_8187,N_4326,N_5003);
nor U8188 (N_8188,N_5033,N_4209);
nor U8189 (N_8189,N_5287,N_4062);
nor U8190 (N_8190,N_6572,N_5560);
or U8191 (N_8191,N_4760,N_5985);
nor U8192 (N_8192,N_5436,N_4576);
nand U8193 (N_8193,N_5893,N_7667);
nand U8194 (N_8194,N_7304,N_4455);
or U8195 (N_8195,N_7967,N_6944);
nor U8196 (N_8196,N_4804,N_4994);
or U8197 (N_8197,N_7846,N_5480);
nand U8198 (N_8198,N_6872,N_4508);
and U8199 (N_8199,N_5957,N_6570);
and U8200 (N_8200,N_5180,N_6547);
nor U8201 (N_8201,N_6435,N_6569);
or U8202 (N_8202,N_6054,N_7529);
and U8203 (N_8203,N_5021,N_6079);
nor U8204 (N_8204,N_4917,N_4059);
or U8205 (N_8205,N_5363,N_5887);
nand U8206 (N_8206,N_4878,N_6090);
or U8207 (N_8207,N_4602,N_5747);
nor U8208 (N_8208,N_7885,N_5472);
nor U8209 (N_8209,N_5972,N_6720);
nand U8210 (N_8210,N_5019,N_6019);
nor U8211 (N_8211,N_7590,N_7937);
nand U8212 (N_8212,N_4768,N_7753);
or U8213 (N_8213,N_7471,N_6232);
or U8214 (N_8214,N_5723,N_7600);
nor U8215 (N_8215,N_5768,N_7647);
or U8216 (N_8216,N_4950,N_4382);
and U8217 (N_8217,N_7686,N_5993);
nor U8218 (N_8218,N_6297,N_5115);
and U8219 (N_8219,N_5755,N_5798);
nor U8220 (N_8220,N_6521,N_4942);
nor U8221 (N_8221,N_4371,N_7165);
or U8222 (N_8222,N_6597,N_5354);
and U8223 (N_8223,N_5285,N_6156);
nand U8224 (N_8224,N_6650,N_7802);
and U8225 (N_8225,N_4863,N_4836);
or U8226 (N_8226,N_7038,N_4458);
and U8227 (N_8227,N_7682,N_7983);
and U8228 (N_8228,N_4400,N_7850);
nand U8229 (N_8229,N_5047,N_7032);
nand U8230 (N_8230,N_7500,N_6931);
or U8231 (N_8231,N_5528,N_4191);
or U8232 (N_8232,N_6765,N_6916);
nor U8233 (N_8233,N_4483,N_4838);
nor U8234 (N_8234,N_4551,N_4064);
or U8235 (N_8235,N_4269,N_6634);
or U8236 (N_8236,N_6995,N_6902);
or U8237 (N_8237,N_5063,N_7112);
nor U8238 (N_8238,N_4163,N_4035);
nand U8239 (N_8239,N_5797,N_5214);
or U8240 (N_8240,N_4463,N_4903);
or U8241 (N_8241,N_6640,N_7396);
nor U8242 (N_8242,N_6335,N_7195);
and U8243 (N_8243,N_7498,N_4248);
nand U8244 (N_8244,N_5297,N_6918);
nor U8245 (N_8245,N_7385,N_7308);
or U8246 (N_8246,N_4355,N_6014);
and U8247 (N_8247,N_6434,N_4005);
or U8248 (N_8248,N_4500,N_5827);
or U8249 (N_8249,N_4849,N_6958);
nand U8250 (N_8250,N_7051,N_6716);
and U8251 (N_8251,N_4833,N_4343);
nor U8252 (N_8252,N_5413,N_5093);
and U8253 (N_8253,N_7421,N_4368);
nor U8254 (N_8254,N_7760,N_5839);
nor U8255 (N_8255,N_5445,N_4695);
and U8256 (N_8256,N_6542,N_6063);
nand U8257 (N_8257,N_4484,N_5394);
and U8258 (N_8258,N_7325,N_7144);
nor U8259 (N_8259,N_7249,N_4404);
or U8260 (N_8260,N_7157,N_7185);
xor U8261 (N_8261,N_7568,N_7124);
nand U8262 (N_8262,N_5883,N_6112);
or U8263 (N_8263,N_4669,N_5539);
or U8264 (N_8264,N_6382,N_4666);
xor U8265 (N_8265,N_5561,N_7467);
and U8266 (N_8266,N_5159,N_6811);
nand U8267 (N_8267,N_7530,N_4936);
and U8268 (N_8268,N_4293,N_5429);
xor U8269 (N_8269,N_5949,N_7544);
nand U8270 (N_8270,N_6415,N_5191);
or U8271 (N_8271,N_5004,N_7228);
or U8272 (N_8272,N_4068,N_4133);
nor U8273 (N_8273,N_7257,N_6320);
or U8274 (N_8274,N_4792,N_5774);
and U8275 (N_8275,N_4652,N_5181);
nand U8276 (N_8276,N_6207,N_5983);
or U8277 (N_8277,N_7794,N_5963);
and U8278 (N_8278,N_4270,N_5355);
nor U8279 (N_8279,N_6924,N_4283);
and U8280 (N_8280,N_6807,N_7527);
and U8281 (N_8281,N_5090,N_7588);
nor U8282 (N_8282,N_6219,N_6914);
or U8283 (N_8283,N_4423,N_4310);
nor U8284 (N_8284,N_4190,N_6159);
and U8285 (N_8285,N_5325,N_5170);
nor U8286 (N_8286,N_6102,N_5694);
and U8287 (N_8287,N_7458,N_6305);
nor U8288 (N_8288,N_4243,N_5043);
nor U8289 (N_8289,N_6884,N_4690);
and U8290 (N_8290,N_5569,N_7831);
nor U8291 (N_8291,N_7409,N_7841);
or U8292 (N_8292,N_6352,N_5049);
nand U8293 (N_8293,N_6927,N_5468);
and U8294 (N_8294,N_4174,N_5260);
nor U8295 (N_8295,N_6493,N_5525);
nor U8296 (N_8296,N_4084,N_6700);
nor U8297 (N_8297,N_5022,N_4582);
nand U8298 (N_8298,N_7610,N_7879);
nand U8299 (N_8299,N_4138,N_5145);
nand U8300 (N_8300,N_7189,N_6694);
nand U8301 (N_8301,N_7811,N_6233);
and U8302 (N_8302,N_5137,N_5970);
nand U8303 (N_8303,N_6221,N_7080);
nand U8304 (N_8304,N_7571,N_6970);
or U8305 (N_8305,N_6973,N_7696);
and U8306 (N_8306,N_7982,N_5741);
nor U8307 (N_8307,N_5365,N_6616);
nor U8308 (N_8308,N_4158,N_7479);
nor U8309 (N_8309,N_6440,N_5397);
or U8310 (N_8310,N_6710,N_5679);
and U8311 (N_8311,N_5522,N_7435);
nand U8312 (N_8312,N_4603,N_7029);
nor U8313 (N_8313,N_7161,N_5751);
nand U8314 (N_8314,N_5324,N_5844);
and U8315 (N_8315,N_4661,N_6727);
nand U8316 (N_8316,N_4839,N_6092);
nor U8317 (N_8317,N_7644,N_7950);
nor U8318 (N_8318,N_7972,N_7392);
nor U8319 (N_8319,N_5165,N_4869);
nor U8320 (N_8320,N_7230,N_5031);
nor U8321 (N_8321,N_6060,N_6454);
nor U8322 (N_8322,N_4535,N_4939);
nand U8323 (N_8323,N_7046,N_4247);
or U8324 (N_8324,N_5379,N_7483);
nand U8325 (N_8325,N_4002,N_7219);
nand U8326 (N_8326,N_5668,N_7512);
nand U8327 (N_8327,N_4977,N_7736);
nor U8328 (N_8328,N_5998,N_4864);
or U8329 (N_8329,N_4286,N_4296);
nand U8330 (N_8330,N_5733,N_4771);
and U8331 (N_8331,N_4153,N_4182);
or U8332 (N_8332,N_5979,N_6419);
and U8333 (N_8333,N_6312,N_7861);
nor U8334 (N_8334,N_7844,N_7619);
nand U8335 (N_8335,N_6586,N_4884);
nor U8336 (N_8336,N_7699,N_5085);
nand U8337 (N_8337,N_6124,N_6707);
nor U8338 (N_8338,N_7847,N_7023);
and U8339 (N_8339,N_7188,N_6751);
nor U8340 (N_8340,N_5866,N_5737);
nor U8341 (N_8341,N_5626,N_6699);
or U8342 (N_8342,N_6741,N_5184);
and U8343 (N_8343,N_4895,N_4858);
or U8344 (N_8344,N_7545,N_5881);
nor U8345 (N_8345,N_7726,N_5693);
nor U8346 (N_8346,N_4746,N_7606);
nand U8347 (N_8347,N_4453,N_4277);
and U8348 (N_8348,N_4206,N_6862);
or U8349 (N_8349,N_7924,N_7716);
and U8350 (N_8350,N_6619,N_7223);
and U8351 (N_8351,N_5266,N_5273);
and U8352 (N_8352,N_7166,N_5508);
nor U8353 (N_8353,N_6553,N_7477);
nand U8354 (N_8354,N_5607,N_6917);
nor U8355 (N_8355,N_6409,N_7456);
and U8356 (N_8356,N_6339,N_5106);
nor U8357 (N_8357,N_4092,N_6633);
nor U8358 (N_8358,N_4805,N_4313);
nor U8359 (N_8359,N_5520,N_4008);
nor U8360 (N_8360,N_5220,N_5189);
nor U8361 (N_8361,N_7499,N_7547);
and U8362 (N_8362,N_7168,N_5259);
or U8363 (N_8363,N_5161,N_4681);
and U8364 (N_8364,N_6627,N_7690);
or U8365 (N_8365,N_5943,N_7874);
xor U8366 (N_8366,N_4027,N_4831);
nor U8367 (N_8367,N_4633,N_6835);
or U8368 (N_8368,N_5932,N_7087);
and U8369 (N_8369,N_5914,N_4593);
and U8370 (N_8370,N_6398,N_7473);
nand U8371 (N_8371,N_6281,N_5054);
nand U8372 (N_8372,N_6740,N_6898);
or U8373 (N_8373,N_7826,N_7707);
nand U8374 (N_8374,N_5132,N_5483);
or U8375 (N_8375,N_4640,N_4783);
nand U8376 (N_8376,N_4944,N_5848);
nand U8377 (N_8377,N_5564,N_4811);
or U8378 (N_8378,N_4436,N_7795);
and U8379 (N_8379,N_5956,N_5038);
and U8380 (N_8380,N_7084,N_4572);
nor U8381 (N_8381,N_4554,N_5989);
or U8382 (N_8382,N_7720,N_5614);
nor U8383 (N_8383,N_7160,N_6306);
or U8384 (N_8384,N_6915,N_7868);
nand U8385 (N_8385,N_4888,N_6851);
nand U8386 (N_8386,N_7709,N_6100);
nor U8387 (N_8387,N_6638,N_4242);
nor U8388 (N_8388,N_5853,N_5889);
nand U8389 (N_8389,N_6148,N_5740);
nand U8390 (N_8390,N_7817,N_4702);
nor U8391 (N_8391,N_4615,N_4325);
nand U8392 (N_8392,N_4766,N_6522);
and U8393 (N_8393,N_6133,N_5621);
nand U8394 (N_8394,N_6110,N_4330);
nor U8395 (N_8395,N_4410,N_5029);
and U8396 (N_8396,N_5111,N_4495);
nor U8397 (N_8397,N_7540,N_6023);
and U8398 (N_8398,N_5537,N_5867);
or U8399 (N_8399,N_7738,N_7303);
and U8400 (N_8400,N_4879,N_6037);
nand U8401 (N_8401,N_4333,N_6826);
or U8402 (N_8402,N_6736,N_4982);
and U8403 (N_8403,N_6904,N_6198);
nand U8404 (N_8404,N_7963,N_6367);
and U8405 (N_8405,N_4505,N_6676);
and U8406 (N_8406,N_4686,N_7073);
nor U8407 (N_8407,N_5982,N_5884);
and U8408 (N_8408,N_6401,N_7069);
nand U8409 (N_8409,N_7263,N_7395);
or U8410 (N_8410,N_7431,N_4910);
nand U8411 (N_8411,N_5493,N_7040);
and U8412 (N_8412,N_7194,N_6480);
nand U8413 (N_8413,N_6236,N_4177);
and U8414 (N_8414,N_4122,N_6366);
nand U8415 (N_8415,N_5645,N_7697);
nor U8416 (N_8416,N_5223,N_6226);
and U8417 (N_8417,N_6467,N_7202);
nor U8418 (N_8418,N_4580,N_6137);
or U8419 (N_8419,N_7889,N_6158);
and U8420 (N_8420,N_4266,N_6746);
nand U8421 (N_8421,N_5083,N_7476);
or U8422 (N_8422,N_5254,N_7244);
and U8423 (N_8423,N_5700,N_5854);
and U8424 (N_8424,N_4629,N_4348);
and U8425 (N_8425,N_7079,N_7323);
nor U8426 (N_8426,N_5330,N_6176);
nor U8427 (N_8427,N_7509,N_5128);
xnor U8428 (N_8428,N_7089,N_5933);
or U8429 (N_8429,N_5055,N_4743);
and U8430 (N_8430,N_6457,N_5948);
nand U8431 (N_8431,N_7896,N_7918);
or U8432 (N_8432,N_4197,N_7227);
nand U8433 (N_8433,N_7391,N_4600);
nand U8434 (N_8434,N_7714,N_7179);
nand U8435 (N_8435,N_7141,N_4258);
and U8436 (N_8436,N_4851,N_6353);
nand U8437 (N_8437,N_5486,N_4656);
or U8438 (N_8438,N_7163,N_5623);
and U8439 (N_8439,N_4714,N_5925);
nand U8440 (N_8440,N_6317,N_7248);
and U8441 (N_8441,N_6296,N_5713);
and U8442 (N_8442,N_4817,N_5608);
nor U8443 (N_8443,N_5382,N_7380);
nand U8444 (N_8444,N_7781,N_7541);
or U8445 (N_8445,N_6730,N_4473);
and U8446 (N_8446,N_5120,N_5407);
and U8447 (N_8447,N_7293,N_5658);
or U8448 (N_8448,N_6071,N_4853);
nor U8449 (N_8449,N_5630,N_5504);
and U8450 (N_8450,N_7554,N_7193);
and U8451 (N_8451,N_6768,N_6518);
and U8452 (N_8452,N_7442,N_6867);
nand U8453 (N_8453,N_4352,N_7894);
nand U8454 (N_8454,N_7024,N_4462);
nand U8455 (N_8455,N_5691,N_5975);
and U8456 (N_8456,N_6798,N_6013);
and U8457 (N_8457,N_4751,N_5712);
nand U8458 (N_8458,N_4108,N_7692);
or U8459 (N_8459,N_4900,N_5406);
or U8460 (N_8460,N_7070,N_5399);
nor U8461 (N_8461,N_4812,N_6980);
nor U8462 (N_8462,N_5250,N_4388);
nand U8463 (N_8463,N_6938,N_4947);
nand U8464 (N_8464,N_6592,N_6362);
nor U8465 (N_8465,N_7804,N_4802);
or U8466 (N_8466,N_7774,N_6406);
and U8467 (N_8467,N_7676,N_6408);
and U8468 (N_8468,N_4019,N_7110);
and U8469 (N_8469,N_5678,N_5232);
or U8470 (N_8470,N_4314,N_7613);
nand U8471 (N_8471,N_4413,N_4653);
nand U8472 (N_8472,N_7927,N_4055);
nor U8473 (N_8473,N_6266,N_7020);
or U8474 (N_8474,N_4992,N_6463);
and U8475 (N_8475,N_4034,N_6659);
and U8476 (N_8476,N_5039,N_7819);
nor U8477 (N_8477,N_7576,N_5221);
or U8478 (N_8478,N_4215,N_5665);
nand U8479 (N_8479,N_7104,N_6300);
xor U8480 (N_8480,N_6585,N_5028);
or U8481 (N_8481,N_5196,N_6376);
nand U8482 (N_8482,N_5776,N_4121);
or U8483 (N_8483,N_4850,N_6857);
nor U8484 (N_8484,N_4475,N_5434);
nor U8485 (N_8485,N_6796,N_6988);
or U8486 (N_8486,N_7872,N_5711);
and U8487 (N_8487,N_5168,N_5818);
nand U8488 (N_8488,N_4376,N_4534);
or U8489 (N_8489,N_7765,N_6802);
nor U8490 (N_8490,N_6870,N_4435);
nand U8491 (N_8491,N_6359,N_4529);
nand U8492 (N_8492,N_4161,N_6374);
nand U8493 (N_8493,N_7663,N_5492);
and U8494 (N_8494,N_5329,N_6330);
nand U8495 (N_8495,N_4416,N_6709);
and U8496 (N_8496,N_6438,N_5507);
nor U8497 (N_8497,N_4078,N_6178);
or U8498 (N_8498,N_7951,N_6635);
nor U8499 (N_8499,N_6706,N_5858);
and U8500 (N_8500,N_5727,N_4272);
and U8501 (N_8501,N_5659,N_7865);
and U8502 (N_8502,N_4408,N_5940);
or U8503 (N_8503,N_4015,N_5341);
nand U8504 (N_8504,N_7941,N_7630);
xnor U8505 (N_8505,N_7966,N_7121);
and U8506 (N_8506,N_7065,N_7286);
nor U8507 (N_8507,N_5453,N_6879);
and U8508 (N_8508,N_4762,N_7484);
nand U8509 (N_8509,N_5760,N_4173);
nand U8510 (N_8510,N_6196,N_5323);
and U8511 (N_8511,N_7852,N_6475);
or U8512 (N_8512,N_4492,N_4662);
nor U8513 (N_8513,N_4682,N_6043);
nand U8514 (N_8514,N_7353,N_5637);
or U8515 (N_8515,N_7510,N_7252);
or U8516 (N_8516,N_4498,N_6969);
nor U8517 (N_8517,N_4860,N_6590);
nand U8518 (N_8518,N_5116,N_7902);
or U8519 (N_8519,N_7790,N_6083);
nor U8520 (N_8520,N_6605,N_7317);
nor U8521 (N_8521,N_6630,N_5140);
nor U8522 (N_8522,N_6906,N_4557);
and U8523 (N_8523,N_4152,N_5515);
and U8524 (N_8524,N_6132,N_6645);
or U8525 (N_8525,N_4968,N_6781);
nor U8526 (N_8526,N_7221,N_7047);
nor U8527 (N_8527,N_4943,N_6118);
and U8528 (N_8528,N_6116,N_4617);
and U8529 (N_8529,N_5714,N_7015);
and U8530 (N_8530,N_6468,N_7355);
nand U8531 (N_8531,N_7632,N_4929);
nor U8532 (N_8532,N_7984,N_4958);
nor U8533 (N_8533,N_4938,N_6446);
nand U8534 (N_8534,N_6831,N_6414);
and U8535 (N_8535,N_7710,N_7744);
nand U8536 (N_8536,N_4909,N_7642);
and U8537 (N_8537,N_6965,N_6495);
nand U8538 (N_8538,N_6392,N_5309);
nor U8539 (N_8539,N_7880,N_7127);
and U8540 (N_8540,N_5158,N_6758);
and U8541 (N_8541,N_4892,N_5162);
or U8542 (N_8542,N_7204,N_4645);
or U8543 (N_8543,N_4680,N_6651);
nand U8544 (N_8544,N_7139,N_4109);
and U8545 (N_8545,N_5762,N_7214);
and U8546 (N_8546,N_5997,N_4309);
nor U8547 (N_8547,N_7132,N_4082);
nor U8548 (N_8548,N_4124,N_4216);
nand U8549 (N_8549,N_5891,N_5268);
xnor U8550 (N_8550,N_6728,N_7049);
or U8551 (N_8551,N_5510,N_6416);
nand U8552 (N_8552,N_5473,N_7180);
and U8553 (N_8553,N_7489,N_4688);
or U8554 (N_8554,N_5421,N_7653);
nor U8555 (N_8555,N_4210,N_4887);
and U8556 (N_8556,N_5864,N_5316);
nand U8557 (N_8557,N_7198,N_7256);
nor U8558 (N_8558,N_6786,N_4459);
nand U8559 (N_8559,N_5353,N_4945);
and U8560 (N_8560,N_5065,N_4380);
nor U8561 (N_8561,N_7601,N_6509);
or U8562 (N_8562,N_5815,N_6974);
or U8563 (N_8563,N_4318,N_5173);
nand U8564 (N_8564,N_6595,N_7152);
nand U8565 (N_8565,N_6443,N_4721);
nor U8566 (N_8566,N_5104,N_5372);
nor U8567 (N_8567,N_4883,N_4788);
or U8568 (N_8568,N_4281,N_7118);
or U8569 (N_8569,N_6667,N_5650);
and U8570 (N_8570,N_7183,N_7809);
and U8571 (N_8571,N_5785,N_5828);
or U8572 (N_8572,N_7533,N_4605);
nor U8573 (N_8573,N_4321,N_5241);
or U8574 (N_8574,N_7408,N_6424);
nor U8575 (N_8575,N_4997,N_4111);
or U8576 (N_8576,N_7403,N_5689);
nor U8577 (N_8577,N_7005,N_5635);
nor U8578 (N_8578,N_6611,N_5822);
or U8579 (N_8579,N_6042,N_5841);
and U8580 (N_8580,N_4431,N_5269);
nor U8581 (N_8581,N_7749,N_4699);
nand U8582 (N_8582,N_5834,N_6838);
and U8583 (N_8583,N_7701,N_5882);
nand U8584 (N_8584,N_5984,N_5058);
and U8585 (N_8585,N_4785,N_7964);
or U8586 (N_8586,N_6500,N_4650);
and U8587 (N_8587,N_6878,N_5988);
or U8588 (N_8588,N_7665,N_7251);
nand U8589 (N_8589,N_4981,N_6608);
nor U8590 (N_8590,N_5248,N_6648);
nor U8591 (N_8591,N_4579,N_7420);
and U8592 (N_8592,N_6853,N_7715);
and U8593 (N_8593,N_7974,N_5331);
and U8594 (N_8594,N_6749,N_5805);
nand U8595 (N_8595,N_7987,N_7107);
or U8596 (N_8596,N_7305,N_7806);
or U8597 (N_8597,N_7357,N_7050);
and U8598 (N_8598,N_4827,N_5304);
and U8599 (N_8599,N_4971,N_6941);
or U8600 (N_8600,N_6808,N_5016);
and U8601 (N_8601,N_7609,N_4089);
xor U8602 (N_8602,N_5257,N_4198);
or U8603 (N_8603,N_4159,N_4398);
nand U8604 (N_8604,N_6905,N_4143);
nor U8605 (N_8605,N_7250,N_5199);
and U8606 (N_8606,N_6190,N_4327);
nor U8607 (N_8607,N_4395,N_7836);
nand U8608 (N_8608,N_6830,N_4588);
and U8609 (N_8609,N_6269,N_6624);
nand U8610 (N_8610,N_4178,N_5095);
or U8611 (N_8611,N_6469,N_4252);
nand U8612 (N_8612,N_6246,N_7414);
nor U8613 (N_8613,N_6164,N_6593);
nor U8614 (N_8614,N_6274,N_5908);
and U8615 (N_8615,N_5605,N_7232);
nand U8616 (N_8616,N_6578,N_4134);
nand U8617 (N_8617,N_6643,N_6987);
or U8618 (N_8618,N_6251,N_7910);
or U8619 (N_8619,N_5175,N_6819);
or U8620 (N_8620,N_6119,N_6180);
and U8621 (N_8621,N_6909,N_6823);
nor U8622 (N_8622,N_6812,N_7869);
and U8623 (N_8623,N_5701,N_7561);
and U8624 (N_8624,N_7882,N_4297);
nand U8625 (N_8625,N_7233,N_4636);
nor U8626 (N_8626,N_5880,N_5041);
nand U8627 (N_8627,N_7350,N_4208);
nand U8628 (N_8628,N_7345,N_4487);
nor U8629 (N_8629,N_5796,N_7890);
nor U8630 (N_8630,N_4504,N_4478);
and U8631 (N_8631,N_5320,N_6785);
nor U8632 (N_8632,N_6673,N_6436);
or U8633 (N_8633,N_4707,N_6080);
or U8634 (N_8634,N_7071,N_5201);
nor U8635 (N_8635,N_7855,N_4957);
or U8636 (N_8636,N_4670,N_5651);
nand U8637 (N_8637,N_6591,N_7021);
or U8638 (N_8638,N_4698,N_4448);
nand U8639 (N_8639,N_5290,N_6782);
xor U8640 (N_8640,N_7362,N_6205);
nor U8641 (N_8641,N_5690,N_4001);
nand U8642 (N_8642,N_6078,N_6664);
or U8643 (N_8643,N_7534,N_5550);
xnor U8644 (N_8644,N_6504,N_6537);
and U8645 (N_8645,N_4287,N_6182);
nor U8646 (N_8646,N_5218,N_4168);
and U8647 (N_8647,N_4339,N_7793);
nor U8648 (N_8648,N_7506,N_7406);
or U8649 (N_8649,N_4289,N_4245);
or U8650 (N_8650,N_5885,N_4586);
or U8651 (N_8651,N_4193,N_7063);
and U8652 (N_8652,N_6653,N_7444);
nor U8653 (N_8653,N_5824,N_4386);
nand U8654 (N_8654,N_4229,N_5905);
or U8655 (N_8655,N_4753,N_5649);
nand U8656 (N_8656,N_5838,N_7526);
and U8657 (N_8657,N_7747,N_7105);
or U8658 (N_8658,N_6871,N_5366);
and U8659 (N_8659,N_4744,N_6323);
or U8660 (N_8660,N_6818,N_4581);
nand U8661 (N_8661,N_7400,N_5784);
or U8662 (N_8662,N_5860,N_7298);
and U8663 (N_8663,N_6877,N_4379);
and U8664 (N_8664,N_5739,N_6698);
or U8665 (N_8665,N_4516,N_5025);
and U8666 (N_8666,N_7045,N_5253);
and U8667 (N_8667,N_5386,N_6800);
and U8668 (N_8668,N_5367,N_7359);
nor U8669 (N_8669,N_4719,N_4449);
nand U8670 (N_8670,N_7260,N_7807);
nor U8671 (N_8671,N_6663,N_6231);
and U8672 (N_8672,N_7128,N_4199);
or U8673 (N_8673,N_6160,N_6508);
nand U8674 (N_8674,N_7853,N_5420);
or U8675 (N_8675,N_6589,N_7528);
xnor U8676 (N_8676,N_4362,N_4342);
and U8677 (N_8677,N_6747,N_4186);
nor U8678 (N_8678,N_4250,N_7319);
or U8679 (N_8679,N_5591,N_5392);
nand U8680 (N_8680,N_4345,N_6135);
or U8681 (N_8681,N_6070,N_5627);
and U8682 (N_8682,N_4787,N_7786);
nand U8683 (N_8683,N_4948,N_7482);
nor U8684 (N_8684,N_4843,N_5121);
nor U8685 (N_8685,N_4842,N_4482);
nor U8686 (N_8686,N_5333,N_4790);
nor U8687 (N_8687,N_4986,N_6479);
and U8688 (N_8688,N_5597,N_4584);
and U8689 (N_8689,N_6465,N_6459);
or U8690 (N_8690,N_5361,N_7829);
and U8691 (N_8691,N_7375,N_4974);
nand U8692 (N_8692,N_5442,N_7349);
nand U8693 (N_8693,N_7958,N_5023);
nand U8694 (N_8694,N_6145,N_5373);
nor U8695 (N_8695,N_5947,N_5289);
or U8696 (N_8696,N_4029,N_4043);
or U8697 (N_8697,N_5401,N_4873);
nor U8698 (N_8698,N_7487,N_4037);
and U8699 (N_8699,N_7562,N_4344);
and U8700 (N_8700,N_6555,N_6674);
and U8701 (N_8701,N_4822,N_5802);
and U8702 (N_8702,N_7386,N_6109);
and U8703 (N_8703,N_7881,N_6564);
and U8704 (N_8704,N_7182,N_7424);
or U8705 (N_8705,N_7999,N_5459);
and U8706 (N_8706,N_7101,N_6095);
or U8707 (N_8707,N_7318,N_6803);
and U8708 (N_8708,N_4704,N_6417);
and U8709 (N_8709,N_4837,N_4069);
or U8710 (N_8710,N_7146,N_7712);
nand U8711 (N_8711,N_4175,N_7018);
and U8712 (N_8712,N_5729,N_5009);
and U8713 (N_8713,N_7670,N_6992);
or U8714 (N_8714,N_7597,N_7901);
nand U8715 (N_8715,N_6052,N_5439);
nor U8716 (N_8716,N_5562,N_4926);
or U8717 (N_8717,N_4101,N_7093);
or U8718 (N_8718,N_5763,N_6245);
nand U8719 (N_8719,N_5748,N_4407);
or U8720 (N_8720,N_5980,N_7468);
and U8721 (N_8721,N_4647,N_6512);
nor U8722 (N_8722,N_4601,N_6813);
nor U8723 (N_8723,N_6429,N_7125);
nor U8724 (N_8724,N_7933,N_6759);
and U8725 (N_8725,N_4120,N_6349);
nand U8726 (N_8726,N_4608,N_7803);
nand U8727 (N_8727,N_4429,N_4856);
or U8728 (N_8728,N_5586,N_6091);
or U8729 (N_8729,N_5611,N_4306);
and U8730 (N_8730,N_7213,N_4610);
nand U8731 (N_8731,N_5037,N_5084);
or U8732 (N_8732,N_6325,N_5954);
and U8733 (N_8733,N_7205,N_6955);
nand U8734 (N_8734,N_7675,N_4747);
and U8735 (N_8735,N_4891,N_6936);
nand U8736 (N_8736,N_4793,N_4855);
and U8737 (N_8737,N_6804,N_5347);
nand U8738 (N_8738,N_7116,N_5319);
nand U8739 (N_8739,N_5177,N_4901);
and U8740 (N_8740,N_4543,N_5138);
nor U8741 (N_8741,N_7863,N_5877);
nor U8742 (N_8742,N_6099,N_7315);
nor U8743 (N_8743,N_4574,N_5996);
nand U8744 (N_8744,N_6501,N_6750);
nor U8745 (N_8745,N_6045,N_4711);
nand U8746 (N_8746,N_4194,N_4411);
or U8747 (N_8747,N_5150,N_7151);
nor U8748 (N_8748,N_4540,N_4528);
nor U8749 (N_8749,N_7462,N_4870);
or U8750 (N_8750,N_6248,N_7265);
xor U8751 (N_8751,N_4759,N_6510);
nand U8752 (N_8752,N_5046,N_4147);
or U8753 (N_8753,N_7563,N_7077);
or U8754 (N_8754,N_6901,N_6397);
and U8755 (N_8755,N_7076,N_7384);
nand U8756 (N_8756,N_5731,N_5995);
nor U8757 (N_8757,N_6549,N_5962);
nand U8758 (N_8758,N_4390,N_7604);
or U8759 (N_8759,N_6028,N_4117);
nor U8760 (N_8760,N_4447,N_5265);
and U8761 (N_8761,N_5764,N_5458);
or U8762 (N_8762,N_5308,N_7099);
nand U8763 (N_8763,N_7558,N_7511);
nand U8764 (N_8764,N_7518,N_5928);
or U8765 (N_8765,N_7524,N_4530);
nand U8766 (N_8766,N_7279,N_6793);
and U8767 (N_8767,N_6725,N_6952);
and U8768 (N_8768,N_6657,N_5545);
or U8769 (N_8769,N_5292,N_4477);
nor U8770 (N_8770,N_4360,N_7623);
or U8771 (N_8771,N_4367,N_7946);
nand U8772 (N_8772,N_4094,N_6217);
nand U8773 (N_8773,N_5636,N_4456);
and U8774 (N_8774,N_5973,N_4192);
nand U8775 (N_8775,N_4160,N_4807);
nand U8776 (N_8776,N_7461,N_7014);
or U8777 (N_8777,N_4291,N_6007);
and U8778 (N_8778,N_6675,N_5722);
and U8779 (N_8779,N_4115,N_4185);
nand U8780 (N_8780,N_4331,N_5521);
nor U8781 (N_8781,N_7155,N_6487);
and U8782 (N_8782,N_6939,N_6448);
nor U8783 (N_8783,N_4820,N_7777);
nand U8784 (N_8784,N_4312,N_7959);
or U8785 (N_8785,N_7989,N_4457);
nand U8786 (N_8786,N_4525,N_5641);
nand U8787 (N_8787,N_6218,N_6418);
and U8788 (N_8788,N_6388,N_7448);
and U8789 (N_8789,N_7437,N_7641);
nor U8790 (N_8790,N_4526,N_7677);
xnor U8791 (N_8791,N_4020,N_7754);
nand U8792 (N_8792,N_5005,N_4692);
nor U8793 (N_8793,N_6687,N_5080);
or U8794 (N_8794,N_6195,N_5415);
nor U8795 (N_8795,N_6492,N_6966);
or U8796 (N_8796,N_4070,N_5557);
nor U8797 (N_8797,N_5618,N_6455);
and U8798 (N_8798,N_7117,N_5919);
and U8799 (N_8799,N_5568,N_7331);
and U8800 (N_8800,N_5359,N_5408);
or U8801 (N_8801,N_5000,N_5444);
or U8802 (N_8802,N_6460,N_4474);
and U8803 (N_8803,N_5725,N_7169);
nand U8804 (N_8804,N_4925,N_7130);
and U8805 (N_8805,N_5129,N_6647);
xnor U8806 (N_8806,N_7238,N_7247);
or U8807 (N_8807,N_5969,N_6268);
and U8808 (N_8808,N_7862,N_4260);
or U8809 (N_8809,N_6858,N_6254);
nand U8810 (N_8810,N_4179,N_6183);
or U8811 (N_8811,N_5907,N_7940);
and U8812 (N_8812,N_7135,N_7867);
or U8813 (N_8813,N_7566,N_6074);
nor U8814 (N_8814,N_6282,N_6437);
nand U8815 (N_8815,N_4292,N_7242);
nor U8816 (N_8816,N_5108,N_4466);
nand U8817 (N_8817,N_5499,N_4667);
or U8818 (N_8818,N_7792,N_6250);
nor U8819 (N_8819,N_4784,N_5067);
nor U8820 (N_8820,N_7091,N_6234);
and U8821 (N_8821,N_6332,N_5275);
and U8822 (N_8822,N_5816,N_7943);
xnor U8823 (N_8823,N_7008,N_6291);
xor U8824 (N_8824,N_7695,N_5185);
or U8825 (N_8825,N_5471,N_4969);
and U8826 (N_8826,N_7727,N_4238);
or U8827 (N_8827,N_4119,N_4146);
or U8828 (N_8828,N_4169,N_4391);
and U8829 (N_8829,N_5909,N_6373);
nor U8830 (N_8830,N_6715,N_5642);
and U8831 (N_8831,N_5619,N_6950);
or U8832 (N_8832,N_6840,N_7648);
nor U8833 (N_8833,N_4598,N_4696);
or U8834 (N_8834,N_6756,N_5263);
nor U8835 (N_8835,N_7054,N_6056);
and U8836 (N_8836,N_5873,N_4302);
and U8837 (N_8837,N_4772,N_4244);
xor U8838 (N_8838,N_6151,N_6272);
or U8839 (N_8839,N_4745,N_6990);
and U8840 (N_8840,N_5443,N_6930);
nor U8841 (N_8841,N_6724,N_4727);
nor U8842 (N_8842,N_7608,N_6485);
nor U8843 (N_8843,N_7689,N_5432);
or U8844 (N_8844,N_5345,N_7295);
nor U8845 (N_8845,N_5300,N_6351);
and U8846 (N_8846,N_5481,N_7285);
and U8847 (N_8847,N_4132,N_5195);
and U8848 (N_8848,N_5470,N_5053);
and U8849 (N_8849,N_5417,N_7605);
nand U8850 (N_8850,N_5426,N_7679);
and U8851 (N_8851,N_7994,N_6855);
nor U8852 (N_8852,N_5639,N_5318);
nand U8853 (N_8853,N_4956,N_4042);
and U8854 (N_8854,N_6294,N_7570);
or U8855 (N_8855,N_7092,N_5718);
or U8856 (N_8856,N_7626,N_6141);
nand U8857 (N_8857,N_5758,N_4162);
nor U8858 (N_8858,N_6310,N_6764);
and U8859 (N_8859,N_7027,N_6900);
nand U8860 (N_8860,N_4268,N_4279);
nand U8861 (N_8861,N_7515,N_6483);
or U8862 (N_8862,N_5534,N_5847);
and U8863 (N_8863,N_7553,N_6846);
and U8864 (N_8864,N_7725,N_5427);
or U8865 (N_8865,N_6963,N_6948);
or U8866 (N_8866,N_4426,N_4523);
and U8867 (N_8867,N_6228,N_5464);
nor U8868 (N_8868,N_6940,N_6471);
or U8869 (N_8869,N_5348,N_4626);
nand U8870 (N_8870,N_7453,N_4796);
nand U8871 (N_8871,N_6954,N_4731);
and U8872 (N_8872,N_6123,N_5474);
nand U8873 (N_8873,N_5643,N_6584);
or U8874 (N_8874,N_7596,N_4777);
nand U8875 (N_8875,N_4641,N_6044);
or U8876 (N_8876,N_7313,N_6032);
or U8877 (N_8877,N_6345,N_5553);
nand U8878 (N_8878,N_6770,N_6072);
and U8879 (N_8879,N_6202,N_4471);
nor U8880 (N_8880,N_6163,N_6810);
or U8881 (N_8881,N_4091,N_6693);
nand U8882 (N_8882,N_6432,N_7009);
nor U8883 (N_8883,N_5656,N_5242);
nor U8884 (N_8884,N_5082,N_5936);
nand U8885 (N_8885,N_4789,N_4452);
and U8886 (N_8886,N_6169,N_7129);
nand U8887 (N_8887,N_6682,N_7929);
nor U8888 (N_8888,N_7197,N_6742);
or U8889 (N_8889,N_4569,N_6441);
nor U8890 (N_8890,N_4387,N_5131);
nor U8891 (N_8891,N_4125,N_4518);
and U8892 (N_8892,N_5513,N_7848);
nand U8893 (N_8893,N_7851,N_7328);
or U8894 (N_8894,N_5117,N_7486);
and U8895 (N_8895,N_7678,N_7463);
nor U8896 (N_8896,N_7474,N_5479);
nor U8897 (N_8897,N_5209,N_7821);
nand U8898 (N_8898,N_4709,N_5892);
or U8899 (N_8899,N_4733,N_6734);
and U8900 (N_8900,N_5466,N_6117);
and U8901 (N_8901,N_6801,N_7657);
nor U8902 (N_8902,N_7309,N_7772);
nand U8903 (N_8903,N_6111,N_5288);
nand U8904 (N_8904,N_5174,N_5368);
nand U8905 (N_8905,N_7871,N_4975);
and U8906 (N_8906,N_5766,N_7731);
or U8907 (N_8907,N_7870,N_6833);
and U8908 (N_8908,N_5886,N_6881);
or U8909 (N_8909,N_7985,N_6656);
nor U8910 (N_8910,N_5380,N_7342);
xnor U8911 (N_8911,N_6496,N_7742);
or U8912 (N_8912,N_4304,N_7153);
or U8913 (N_8913,N_5079,N_6131);
nor U8914 (N_8914,N_6722,N_6828);
xnor U8915 (N_8915,N_7582,N_5981);
nand U8916 (N_8916,N_5091,N_5087);
and U8917 (N_8917,N_6779,N_4894);
nand U8918 (N_8918,N_4334,N_5648);
nand U8919 (N_8919,N_4234,N_5423);
and U8920 (N_8920,N_7083,N_6660);
nand U8921 (N_8921,N_6193,N_6249);
and U8922 (N_8922,N_7572,N_7404);
nor U8923 (N_8923,N_6913,N_5388);
nand U8924 (N_8924,N_4677,N_7685);
nor U8925 (N_8925,N_5900,N_7485);
nor U8926 (N_8926,N_5192,N_7134);
and U8927 (N_8927,N_5204,N_5390);
or U8928 (N_8928,N_4738,N_5460);
and U8929 (N_8929,N_4966,N_6009);
nor U8930 (N_8930,N_6322,N_5753);
nor U8931 (N_8931,N_5904,N_6945);
nor U8932 (N_8932,N_6557,N_5670);
nand U8933 (N_8933,N_5412,N_5579);
nand U8934 (N_8934,N_6777,N_7897);
or U8935 (N_8935,N_7520,N_6302);
nand U8936 (N_8936,N_6911,N_7906);
or U8937 (N_8937,N_6355,N_5868);
nand U8938 (N_8938,N_6021,N_4442);
nand U8939 (N_8939,N_4219,N_7109);
and U8940 (N_8940,N_4757,N_6017);
nand U8941 (N_8941,N_5946,N_6298);
nor U8942 (N_8942,N_4107,N_4424);
nand U8943 (N_8943,N_5820,N_4425);
or U8944 (N_8944,N_6077,N_5780);
nor U8945 (N_8945,N_6815,N_4741);
nor U8946 (N_8946,N_7056,N_6536);
and U8947 (N_8947,N_5228,N_7297);
or U8948 (N_8948,N_4949,N_7335);
and U8949 (N_8949,N_4213,N_4419);
and U8950 (N_8950,N_5435,N_6174);
or U8951 (N_8951,N_4924,N_6420);
and U8952 (N_8952,N_4556,N_5487);
nand U8953 (N_8953,N_7909,N_6106);
and U8954 (N_8954,N_7968,N_6554);
nand U8955 (N_8955,N_6670,N_5602);
or U8956 (N_8956,N_6821,N_6887);
nor U8957 (N_8957,N_5062,N_7658);
and U8958 (N_8958,N_4921,N_7917);
nand U8959 (N_8959,N_5543,N_7892);
nor U8960 (N_8960,N_6685,N_6532);
nand U8961 (N_8961,N_7812,N_4742);
and U8962 (N_8962,N_7607,N_6303);
or U8963 (N_8963,N_7557,N_4826);
or U8964 (N_8964,N_4432,N_6989);
nand U8965 (N_8965,N_7336,N_7186);
nor U8966 (N_8966,N_6147,N_4539);
nand U8967 (N_8967,N_5042,N_4350);
and U8968 (N_8968,N_4346,N_6662);
or U8969 (N_8969,N_6041,N_4985);
and U8970 (N_8970,N_7706,N_7995);
or U8971 (N_8971,N_6170,N_5461);
and U8972 (N_8972,N_4403,N_5968);
and U8973 (N_8973,N_4612,N_5945);
nand U8974 (N_8974,N_4349,N_5628);
and U8975 (N_8975,N_4676,N_7986);
and U8976 (N_8976,N_5478,N_7044);
nor U8977 (N_8977,N_7339,N_7948);
nor U8978 (N_8978,N_6907,N_4401);
or U8979 (N_8979,N_6717,N_6410);
nor U8980 (N_8980,N_5585,N_6149);
and U8981 (N_8981,N_4867,N_6641);
nor U8982 (N_8982,N_7748,N_6488);
nor U8983 (N_8983,N_4683,N_4775);
nor U8984 (N_8984,N_7508,N_5495);
nand U8985 (N_8985,N_6370,N_5809);
and U8986 (N_8986,N_6933,N_5991);
or U8987 (N_8987,N_4284,N_6427);
nand U8988 (N_8988,N_5450,N_6050);
or U8989 (N_8989,N_7327,N_5449);
or U8990 (N_8990,N_6646,N_7767);
or U8991 (N_8991,N_4819,N_7962);
nor U8992 (N_8992,N_4357,N_5153);
nor U8993 (N_8993,N_5788,N_4657);
nor U8994 (N_8994,N_4857,N_5629);
nor U8995 (N_8995,N_6445,N_6087);
or U8996 (N_8996,N_5574,N_7307);
and U8997 (N_8997,N_7886,N_6790);
or U8998 (N_8998,N_6594,N_6113);
nor U8999 (N_8999,N_4607,N_4778);
nand U9000 (N_9000,N_5178,N_6258);
nor U9001 (N_9001,N_7550,N_6157);
nand U9002 (N_9002,N_5669,N_7569);
and U9003 (N_9003,N_6968,N_5411);
nand U9004 (N_9004,N_4825,N_4749);
nor U9005 (N_9005,N_6925,N_6197);
nand U9006 (N_9006,N_6450,N_6882);
or U9007 (N_9007,N_5542,N_6257);
and U9008 (N_9008,N_7410,N_6743);
nor U9009 (N_9009,N_7970,N_7302);
nor U9010 (N_9010,N_7532,N_6789);
nand U9011 (N_9011,N_5830,N_6984);
nor U9012 (N_9012,N_4022,N_6753);
nor U9013 (N_9013,N_6604,N_5535);
or U9014 (N_9014,N_4693,N_6175);
and U9015 (N_9015,N_6561,N_5227);
and U9016 (N_9016,N_5806,N_7517);
nor U9017 (N_9017,N_5596,N_5186);
nor U9018 (N_9018,N_5952,N_4079);
and U9019 (N_9019,N_7565,N_5572);
nand U9020 (N_9020,N_5567,N_7654);
or U9021 (N_9021,N_5457,N_7235);
or U9022 (N_9022,N_6125,N_7239);
nor U9023 (N_9023,N_5601,N_7322);
nor U9024 (N_9024,N_6334,N_6996);
nor U9025 (N_9025,N_7376,N_4510);
or U9026 (N_9026,N_4916,N_4003);
nand U9027 (N_9027,N_6559,N_5910);
nor U9028 (N_9028,N_7181,N_7513);
nor U9029 (N_9029,N_7614,N_7646);
nor U9030 (N_9030,N_7270,N_4485);
nand U9031 (N_9031,N_5606,N_4180);
or U9032 (N_9032,N_7167,N_7361);
nand U9033 (N_9033,N_4166,N_5182);
nor U9034 (N_9034,N_7100,N_4830);
or U9035 (N_9035,N_6466,N_7947);
or U9036 (N_9036,N_6439,N_6286);
and U9037 (N_9037,N_7907,N_7288);
and U9038 (N_9038,N_6896,N_6375);
and U9039 (N_9039,N_4317,N_4941);
and U9040 (N_9040,N_5249,N_5734);
and U9041 (N_9041,N_7019,N_4689);
and U9042 (N_9042,N_7311,N_7343);
and U9043 (N_9043,N_4596,N_4980);
nand U9044 (N_9044,N_7773,N_4288);
or U9045 (N_9045,N_4126,N_6912);
nor U9046 (N_9046,N_6979,N_7495);
or U9047 (N_9047,N_6545,N_7443);
nand U9048 (N_9048,N_5446,N_4646);
or U9049 (N_9049,N_6200,N_4723);
or U9050 (N_9050,N_5987,N_7521);
nor U9051 (N_9051,N_6729,N_4479);
nand U9052 (N_9052,N_5160,N_7457);
nand U9053 (N_9053,N_7439,N_6688);
and U9054 (N_9054,N_7207,N_6311);
nor U9055 (N_9055,N_4552,N_7751);
or U9056 (N_9056,N_7891,N_5505);
and U9057 (N_9057,N_5819,N_6326);
and U9058 (N_9058,N_5270,N_7969);
and U9059 (N_9059,N_7859,N_7816);
and U9060 (N_9060,N_4940,N_7464);
nand U9061 (N_9061,N_4737,N_7312);
nand U9062 (N_9062,N_7365,N_4493);
or U9063 (N_9063,N_7064,N_6610);
nand U9064 (N_9064,N_6035,N_5559);
and U9065 (N_9065,N_7478,N_6395);
nor U9066 (N_9066,N_6739,N_6921);
nor U9067 (N_9067,N_7001,N_7066);
nand U9068 (N_9068,N_7594,N_4865);
or U9069 (N_9069,N_4225,N_7548);
nand U9070 (N_9070,N_4732,N_4189);
nand U9071 (N_9071,N_4039,N_5594);
nand U9072 (N_9072,N_5098,N_7264);
or U9073 (N_9073,N_4221,N_6890);
nand U9074 (N_9074,N_5894,N_6574);
nor U9075 (N_9075,N_6771,N_6772);
nand U9076 (N_9076,N_5548,N_6097);
and U9077 (N_9077,N_6599,N_7764);
nand U9078 (N_9078,N_7411,N_5541);
and U9079 (N_9079,N_4828,N_7267);
or U9080 (N_9080,N_6201,N_7808);
nor U9081 (N_9081,N_4671,N_6929);
nor U9082 (N_9082,N_7231,N_4040);
and U9083 (N_9083,N_7234,N_6402);
or U9084 (N_9084,N_7334,N_4295);
or U9085 (N_9085,N_4274,N_5448);
and U9086 (N_9086,N_5385,N_7688);
nand U9087 (N_9087,N_5720,N_7405);
nor U9088 (N_9088,N_7425,N_7916);
and U9089 (N_9089,N_4999,N_4085);
nand U9090 (N_9090,N_7843,N_7072);
nor U9091 (N_9091,N_6255,N_7222);
xor U9092 (N_9092,N_6372,N_7412);
nand U9093 (N_9093,N_7680,N_6562);
or U9094 (N_9094,N_4728,N_7586);
nor U9095 (N_9095,N_7900,N_6399);
and U9096 (N_9096,N_4486,N_5002);
or U9097 (N_9097,N_7971,N_6026);
and U9098 (N_9098,N_5447,N_5826);
and U9099 (N_9099,N_6817,N_4261);
and U9100 (N_9100,N_7082,N_7201);
and U9101 (N_9101,N_4983,N_7272);
nor U9102 (N_9102,N_7717,N_6464);
nand U9103 (N_9103,N_6096,N_4509);
and U9104 (N_9104,N_7280,N_6428);
or U9105 (N_9105,N_7269,N_4663);
or U9106 (N_9106,N_4103,N_5852);
or U9107 (N_9107,N_6744,N_6384);
nand U9108 (N_9108,N_4445,N_4567);
or U9109 (N_9109,N_5203,N_7693);
and U9110 (N_9110,N_7413,N_4128);
or U9111 (N_9111,N_4861,N_4063);
and U9112 (N_9112,N_7684,N_4521);
and U9113 (N_9113,N_6868,N_4434);
or U9114 (N_9114,N_4545,N_6393);
or U9115 (N_9115,N_7301,N_4025);
or U9116 (N_9116,N_6120,N_4156);
nor U9117 (N_9117,N_4106,N_5013);
or U9118 (N_9118,N_4127,N_5393);
nor U9119 (N_9119,N_6062,N_7800);
and U9120 (N_9120,N_6144,N_4480);
nand U9121 (N_9121,N_6762,N_7625);
and U9122 (N_9122,N_7603,N_6059);
nor U9123 (N_9123,N_6377,N_6865);
and U9124 (N_9124,N_7034,N_6654);
and U9125 (N_9125,N_6568,N_6637);
or U9126 (N_9126,N_7497,N_4074);
nand U9127 (N_9127,N_5913,N_7672);
nand U9128 (N_9128,N_4624,N_6166);
nor U9129 (N_9129,N_4875,N_6162);
and U9130 (N_9130,N_5617,N_6607);
or U9131 (N_9131,N_7348,N_5281);
and U9132 (N_9132,N_7827,N_4955);
or U9133 (N_9133,N_4672,N_7952);
nand U9134 (N_9134,N_5589,N_4575);
nand U9135 (N_9135,N_4715,N_4353);
nand U9136 (N_9136,N_7745,N_7915);
or U9137 (N_9137,N_7162,N_5035);
or U9138 (N_9138,N_7200,N_7939);
or U9139 (N_9139,N_7407,N_6240);
nor U9140 (N_9140,N_7796,N_4621);
or U9141 (N_9141,N_7645,N_5583);
and U9142 (N_9142,N_7737,N_5967);
nor U9143 (N_9143,N_6962,N_7028);
nor U9144 (N_9144,N_5770,N_6652);
and U9145 (N_9145,N_7928,N_6982);
and U9146 (N_9146,N_6961,N_5267);
or U9147 (N_9147,N_7373,N_4782);
nand U9148 (N_9148,N_6697,N_4299);
nand U9149 (N_9149,N_6983,N_4150);
and U9150 (N_9150,N_4897,N_4630);
and U9151 (N_9151,N_7732,N_5306);
nor U9152 (N_9152,N_5924,N_6507);
or U9153 (N_9153,N_6034,N_4071);
and U9154 (N_9154,N_6098,N_6520);
nor U9155 (N_9155,N_4212,N_6566);
and U9156 (N_9156,N_4761,N_7096);
nand U9157 (N_9157,N_6220,N_5855);
or U9158 (N_9158,N_7965,N_5166);
and U9159 (N_9159,N_4578,N_4987);
and U9160 (N_9160,N_6655,N_7037);
nand U9161 (N_9161,N_5322,N_6452);
or U9162 (N_9162,N_7430,N_7074);
or U9163 (N_9163,N_6677,N_6922);
or U9164 (N_9164,N_7452,N_5377);
nor U9165 (N_9165,N_5271,N_5715);
nor U9166 (N_9166,N_5831,N_4823);
and U9167 (N_9167,N_4722,N_7393);
nor U9168 (N_9168,N_4705,N_5400);
nand U9169 (N_9169,N_5920,N_5211);
nand U9170 (N_9170,N_5927,N_5342);
nor U9171 (N_9171,N_5144,N_6031);
nand U9172 (N_9172,N_5305,N_4750);
nor U9173 (N_9173,N_4880,N_5313);
and U9174 (N_9174,N_4383,N_6265);
nand U9175 (N_9175,N_6845,N_7276);
and U9176 (N_9176,N_7698,N_7579);
nand U9177 (N_9177,N_4460,N_5813);
nor U9178 (N_9178,N_7724,N_6967);
nand U9179 (N_9179,N_6484,N_6068);
and U9180 (N_9180,N_7022,N_4841);
and U9181 (N_9181,N_7137,N_4809);
nor U9182 (N_9182,N_7055,N_5657);
or U9183 (N_9183,N_6919,N_4273);
nor U9184 (N_9184,N_4016,N_6763);
nor U9185 (N_9185,N_5810,N_4558);
or U9186 (N_9186,N_4654,N_7401);
and U9187 (N_9187,N_5245,N_7122);
or U9188 (N_9188,N_7525,N_6866);
nor U9189 (N_9189,N_6140,N_6055);
nor U9190 (N_9190,N_4767,N_6528);
and U9191 (N_9191,N_5615,N_5451);
nor U9192 (N_9192,N_6277,N_5761);
nand U9193 (N_9193,N_5901,N_7289);
or U9194 (N_9194,N_5593,N_7577);
nor U9195 (N_9195,N_7048,N_5068);
nand U9196 (N_9196,N_4606,N_7224);
nor U9197 (N_9197,N_7656,N_7822);
or U9198 (N_9198,N_7542,N_4438);
and U9199 (N_9199,N_4096,N_4263);
nor U9200 (N_9200,N_4923,N_4057);
and U9201 (N_9201,N_4620,N_5717);
and U9202 (N_9202,N_6535,N_5296);
nor U9203 (N_9203,N_7813,N_7067);
nor U9204 (N_9204,N_6755,N_7011);
nand U9205 (N_9205,N_6761,N_4511);
nor U9206 (N_9206,N_5775,N_5644);
nand U9207 (N_9207,N_6061,N_7031);
nand U9208 (N_9208,N_5516,N_4151);
nor U9209 (N_9209,N_7992,N_7147);
nor U9210 (N_9210,N_5176,N_7176);
and U9211 (N_9211,N_7374,N_7583);
or U9212 (N_9212,N_5119,N_6780);
nand U9213 (N_9213,N_6531,N_5081);
or U9214 (N_9214,N_5974,N_7535);
nor U9215 (N_9215,N_6337,N_5571);
and U9216 (N_9216,N_4300,N_5666);
nand U9217 (N_9217,N_7979,N_7337);
nand U9218 (N_9218,N_4359,N_5843);
nand U9219 (N_9219,N_4130,N_7229);
nand U9220 (N_9220,N_5030,N_5929);
and U9221 (N_9221,N_6404,N_6210);
nor U9222 (N_9222,N_5744,N_7470);
nand U9223 (N_9223,N_6864,N_6413);
or U9224 (N_9224,N_7493,N_5898);
nand U9225 (N_9225,N_6101,N_6859);
nor U9226 (N_9226,N_7460,N_4533);
and U9227 (N_9227,N_7783,N_6283);
or U9228 (N_9228,N_5663,N_6577);
nor U9229 (N_9229,N_5350,N_5207);
nand U9230 (N_9230,N_4920,N_4794);
or U9231 (N_9231,N_7649,N_5633);
nor U9232 (N_9232,N_7496,N_7379);
nand U9233 (N_9233,N_4801,N_4613);
nand U9234 (N_9234,N_6308,N_5476);
and U9235 (N_9235,N_5832,N_6177);
and U9236 (N_9236,N_7945,N_6261);
and U9237 (N_9237,N_6482,N_5890);
or U9238 (N_9238,N_6104,N_4679);
nand U9239 (N_9239,N_7090,N_7585);
and U9240 (N_9240,N_7551,N_6423);
and U9241 (N_9241,N_4890,N_6288);
nor U9242 (N_9242,N_5239,N_4406);
nand U9243 (N_9243,N_6505,N_7290);
and U9244 (N_9244,N_7857,N_6684);
nor U9245 (N_9245,N_6986,N_4631);
nor U9246 (N_9246,N_6391,N_7120);
nor U9247 (N_9247,N_4218,N_5530);
nand U9248 (N_9248,N_5032,N_6669);
or U9249 (N_9249,N_6632,N_4080);
and U9250 (N_9250,N_6262,N_5078);
and U9251 (N_9251,N_4187,N_7114);
or U9252 (N_9252,N_6082,N_6628);
or U9253 (N_9253,N_6481,N_4991);
nor U9254 (N_9254,N_6239,N_7275);
xnor U9255 (N_9255,N_5503,N_4928);
nand U9256 (N_9256,N_4541,N_6179);
xor U9257 (N_9257,N_7912,N_6412);
or U9258 (N_9258,N_5951,N_6018);
or U9259 (N_9259,N_5113,N_5167);
nor U9260 (N_9260,N_5437,N_4341);
nor U9261 (N_9261,N_5859,N_7417);
or U9262 (N_9262,N_6093,N_4638);
and U9263 (N_9263,N_7058,N_7700);
nand U9264 (N_9264,N_7253,N_5647);
or U9265 (N_9265,N_7172,N_6343);
or U9266 (N_9266,N_4597,N_7957);
nand U9267 (N_9267,N_4786,N_7218);
nand U9268 (N_9268,N_5573,N_6161);
or U9269 (N_9269,N_7258,N_6551);
nor U9270 (N_9270,N_7216,N_5736);
nand U9271 (N_9271,N_4226,N_7277);
nand U9272 (N_9272,N_7519,N_7761);
or U9273 (N_9273,N_6895,N_7268);
or U9274 (N_9274,N_4231,N_6271);
nor U9275 (N_9275,N_5899,N_7739);
or U9276 (N_9276,N_4797,N_4240);
and U9277 (N_9277,N_4532,N_7196);
or U9278 (N_9278,N_7143,N_6932);
or U9279 (N_9279,N_7351,N_6613);
nor U9280 (N_9280,N_5066,N_5551);
and U9281 (N_9281,N_5582,N_4795);
nor U9282 (N_9282,N_6295,N_7637);
xnor U9283 (N_9283,N_4148,N_4821);
or U9284 (N_9284,N_6396,N_7330);
nand U9285 (N_9285,N_4549,N_6368);
and U9286 (N_9286,N_7284,N_4469);
nor U9287 (N_9287,N_4660,N_4553);
or U9288 (N_9288,N_6626,N_4315);
or U9289 (N_9289,N_4563,N_7347);
or U9290 (N_9290,N_5018,N_7455);
xnor U9291 (N_9291,N_5219,N_4211);
nand U9292 (N_9292,N_6690,N_4251);
and U9293 (N_9293,N_7573,N_5358);
or U9294 (N_9294,N_5759,N_4565);
nand U9295 (N_9295,N_7292,N_6350);
or U9296 (N_9296,N_6713,N_7057);
and U9297 (N_9297,N_7669,N_6030);
and U9298 (N_9298,N_7687,N_7782);
nand U9299 (N_9299,N_6046,N_4405);
nand U9300 (N_9300,N_6544,N_6702);
and U9301 (N_9301,N_5793,N_5125);
nor U9302 (N_9302,N_4422,N_7281);
and U9303 (N_9303,N_5416,N_6928);
and U9304 (N_9304,N_4239,N_5498);
or U9305 (N_9305,N_6390,N_6150);
or U9306 (N_9306,N_5014,N_6036);
or U9307 (N_9307,N_6403,N_7043);
nand U9308 (N_9308,N_4363,N_5746);
nor U9309 (N_9309,N_6567,N_5653);
or U9310 (N_9310,N_4905,N_4758);
nor U9311 (N_9311,N_4814,N_4262);
nand U9312 (N_9312,N_7587,N_6127);
nand U9313 (N_9313,N_7367,N_4000);
and U9314 (N_9314,N_7620,N_5575);
nor U9315 (N_9315,N_7175,N_5206);
nor U9316 (N_9316,N_5240,N_5790);
or U9317 (N_9317,N_6603,N_4706);
nor U9318 (N_9318,N_7012,N_6703);
nor U9319 (N_9319,N_7956,N_5229);
nand U9320 (N_9320,N_6153,N_6486);
or U9321 (N_9321,N_6313,N_6029);
nor U9322 (N_9322,N_5362,N_7842);
or U9323 (N_9323,N_4583,N_4832);
or U9324 (N_9324,N_7445,N_6860);
nor U9325 (N_9325,N_5931,N_6230);
or U9326 (N_9326,N_4840,N_4673);
and U9327 (N_9327,N_7925,N_6526);
nor U9328 (N_9328,N_6666,N_4440);
and U9329 (N_9329,N_7103,N_6787);
or U9330 (N_9330,N_6216,N_5986);
nor U9331 (N_9331,N_7454,N_6832);
nand U9332 (N_9332,N_6792,N_7115);
and U9333 (N_9333,N_4594,N_4720);
or U9334 (N_9334,N_6491,N_4140);
nand U9335 (N_9335,N_5506,N_4320);
or U9336 (N_9336,N_5613,N_7769);
nand U9337 (N_9337,N_6733,N_5024);
and U9338 (N_9338,N_5126,N_5337);
or U9339 (N_9339,N_6338,N_6256);
nor U9340 (N_9340,N_5311,N_5302);
and U9341 (N_9341,N_6328,N_7643);
nor U9342 (N_9342,N_7638,N_7828);
or U9343 (N_9343,N_7713,N_4561);
and U9344 (N_9344,N_5244,N_7559);
or U9345 (N_9345,N_4116,N_7935);
nand U9346 (N_9346,N_7960,N_4026);
nor U9347 (N_9347,N_6981,N_4235);
nand U9348 (N_9348,N_4155,N_7921);
nor U9349 (N_9349,N_5624,N_5769);
nor U9350 (N_9350,N_6016,N_6529);
nand U9351 (N_9351,N_7820,N_7382);
and U9352 (N_9352,N_6154,N_4417);
or U9353 (N_9353,N_6712,N_4725);
or U9354 (N_9354,N_6738,N_6033);
and U9355 (N_9355,N_7830,N_4619);
and U9356 (N_9356,N_5825,N_5704);
and U9357 (N_9357,N_5875,N_6084);
nand U9358 (N_9358,N_6027,N_4953);
and U9359 (N_9359,N_4908,N_7004);
nand U9360 (N_9360,N_5523,N_4054);
nand U9361 (N_9361,N_6088,N_6665);
nand U9362 (N_9362,N_6754,N_6214);
and U9363 (N_9363,N_5328,N_6206);
nor U9364 (N_9364,N_7344,N_6421);
and U9365 (N_9365,N_4087,N_4507);
nor U9366 (N_9366,N_7978,N_5756);
nor U9367 (N_9367,N_5804,N_4444);
and U9368 (N_9368,N_5870,N_5148);
or U9369 (N_9369,N_5215,N_6426);
nand U9370 (N_9370,N_4765,N_6329);
or U9371 (N_9371,N_5808,N_6293);
xor U9372 (N_9372,N_4735,N_5441);
or U9373 (N_9373,N_5930,N_5008);
or U9374 (N_9374,N_7126,N_5433);
or U9375 (N_9375,N_6203,N_4004);
nor U9376 (N_9376,N_5127,N_7053);
and U9377 (N_9377,N_7814,N_4527);
or U9378 (N_9378,N_7266,N_5684);
or U9379 (N_9379,N_5837,N_4591);
or U9380 (N_9380,N_6073,N_6066);
nand U9381 (N_9381,N_4642,N_7555);
nand U9382 (N_9382,N_6714,N_6820);
nand U9383 (N_9383,N_5710,N_5778);
nand U9384 (N_9384,N_6601,N_6273);
and U9385 (N_9385,N_4139,N_5738);
or U9386 (N_9386,N_7627,N_4932);
nand U9387 (N_9387,N_6573,N_6708);
or U9388 (N_9388,N_7366,N_6517);
and U9389 (N_9389,N_7475,N_7422);
nor U9390 (N_9390,N_6511,N_6461);
nor U9391 (N_9391,N_7681,N_7932);
or U9392 (N_9392,N_4167,N_7721);
nor U9393 (N_9393,N_7310,N_6126);
and U9394 (N_9394,N_6235,N_6065);
nor U9395 (N_9395,N_6726,N_4083);
and U9396 (N_9396,N_7611,N_5105);
or U9397 (N_9397,N_5274,N_7919);
or U9398 (N_9398,N_4674,N_4053);
nand U9399 (N_9399,N_5801,N_4129);
or U9400 (N_9400,N_6957,N_6278);
or U9401 (N_9401,N_5103,N_7030);
or U9402 (N_9402,N_6188,N_6639);
or U9403 (N_9403,N_5692,N_4081);
or U9404 (N_9404,N_7991,N_6222);
or U9405 (N_9405,N_7580,N_6696);
nand U9406 (N_9406,N_6184,N_5001);
nand U9407 (N_9407,N_7086,N_4075);
nor U9408 (N_9408,N_6209,N_5961);
or U9409 (N_9409,N_6649,N_5654);
and U9410 (N_9410,N_6191,N_5151);
and U9411 (N_9411,N_5789,N_7930);
nand U9412 (N_9412,N_7472,N_6004);
nand U9413 (N_9413,N_7360,N_4010);
or U9414 (N_9414,N_4816,N_4246);
nand U9415 (N_9415,N_4984,N_5906);
nand U9416 (N_9416,N_6477,N_4183);
and U9417 (N_9417,N_6365,N_4451);
nand U9418 (N_9418,N_6893,N_7602);
and U9419 (N_9419,N_5490,N_4241);
or U9420 (N_9420,N_5283,N_6558);
nand U9421 (N_9421,N_7934,N_4377);
and U9422 (N_9422,N_7145,N_7639);
nand U9423 (N_9423,N_7164,N_6494);
nand U9424 (N_9424,N_6290,N_4049);
nor U9425 (N_9425,N_5101,N_7490);
and U9426 (N_9426,N_5418,N_7133);
nand U9427 (N_9427,N_5937,N_7539);
nor U9428 (N_9428,N_7402,N_4503);
nor U9429 (N_9429,N_4033,N_7763);
nand U9430 (N_9430,N_7042,N_5475);
and U9431 (N_9431,N_7564,N_6523);
nor U9432 (N_9432,N_6315,N_5566);
or U9433 (N_9433,N_5142,N_6244);
nand U9434 (N_9434,N_5187,N_4259);
and U9435 (N_9435,N_4564,N_6576);
nand U9436 (N_9436,N_6299,N_7287);
nor U9437 (N_9437,N_7666,N_6224);
and U9438 (N_9438,N_6138,N_7592);
nand U9439 (N_9439,N_5698,N_7033);
and U9440 (N_9440,N_5303,N_7598);
nor U9441 (N_9441,N_7504,N_7039);
and U9442 (N_9442,N_4824,N_7502);
and U9443 (N_9443,N_6580,N_4188);
nand U9444 (N_9444,N_5364,N_7138);
and U9445 (N_9445,N_7876,N_5255);
nand U9446 (N_9446,N_7358,N_5338);
nand U9447 (N_9447,N_6341,N_4763);
or U9448 (N_9448,N_4637,N_5246);
nand U9449 (N_9449,N_6347,N_4868);
nor U9450 (N_9450,N_7381,N_6121);
or U9451 (N_9451,N_6143,N_6515);
nand U9452 (N_9452,N_4271,N_7245);
nor U9453 (N_9453,N_5040,N_6444);
nand U9454 (N_9454,N_4919,N_5703);
nand U9455 (N_9455,N_5431,N_4976);
or U9456 (N_9456,N_6692,N_4871);
nor U9457 (N_9457,N_5360,N_5236);
nor U9458 (N_9458,N_6824,N_6022);
nand U9459 (N_9459,N_4098,N_5205);
or U9460 (N_9460,N_4614,N_7449);
nor U9461 (N_9461,N_4322,N_6908);
nor U9462 (N_9462,N_5202,N_4934);
and U9463 (N_9463,N_7633,N_7094);
nand U9464 (N_9464,N_5357,N_5849);
nor U9465 (N_9465,N_5496,N_4384);
or U9466 (N_9466,N_7254,N_5687);
nor U9467 (N_9467,N_7815,N_6008);
or U9468 (N_9468,N_4852,N_6213);
nor U9469 (N_9469,N_4951,N_7387);
nor U9470 (N_9470,N_7729,N_7017);
nand U9471 (N_9471,N_5183,N_7944);
nand U9472 (N_9472,N_4628,N_5829);
and U9473 (N_9473,N_4995,N_5840);
nor U9474 (N_9474,N_7883,N_5048);
and U9475 (N_9475,N_5403,N_6671);
nor U9476 (N_9476,N_4396,N_5061);
or U9477 (N_9477,N_6400,N_5807);
and U9478 (N_9478,N_5558,N_4048);
or U9479 (N_9479,N_4846,N_6571);
or U9480 (N_9480,N_4394,N_6873);
nor U9481 (N_9481,N_5050,N_6048);
nor U9482 (N_9482,N_5977,N_6173);
or U9483 (N_9483,N_5794,N_4736);
nand U9484 (N_9484,N_6212,N_7673);
nor U9485 (N_9485,N_4734,N_4233);
and U9486 (N_9486,N_7271,N_4655);
or U9487 (N_9487,N_5294,N_5842);
nand U9488 (N_9488,N_7516,N_5599);
nand U9489 (N_9489,N_7791,N_5592);
and U9490 (N_9490,N_4439,N_5069);
nor U9491 (N_9491,N_5861,N_7895);
and U9492 (N_9492,N_5321,N_6854);
nor U9493 (N_9493,N_6767,N_6267);
nand U9494 (N_9494,N_6791,N_5959);
and U9495 (N_9495,N_5370,N_6336);
nand U9496 (N_9496,N_4538,N_6242);
or U9497 (N_9497,N_7088,N_4893);
or U9498 (N_9498,N_5264,N_6499);
nand U9499 (N_9499,N_6661,N_5020);
and U9500 (N_9500,N_7755,N_6636);
or U9501 (N_9501,N_4718,N_6839);
nor U9502 (N_9502,N_5404,N_7911);
nand U9503 (N_9503,N_4627,N_7320);
nand U9504 (N_9504,N_5465,N_4014);
nand U9505 (N_9505,N_4964,N_6011);
or U9506 (N_9506,N_4935,N_4978);
nor U9507 (N_9507,N_6880,N_4217);
or U9508 (N_9508,N_4335,N_7988);
nand U9509 (N_9509,N_5109,N_7190);
nor U9510 (N_9510,N_7215,N_5193);
nand U9511 (N_9511,N_7612,N_7798);
nand U9512 (N_9512,N_4803,N_4249);
or U9513 (N_9513,N_4214,N_5419);
and U9514 (N_9514,N_5156,N_6560);
nor U9515 (N_9515,N_4635,N_5251);
nand U9516 (N_9516,N_6502,N_7255);
or U9517 (N_9517,N_7436,N_5256);
nand U9518 (N_9518,N_7780,N_7321);
or U9519 (N_9519,N_5402,N_6869);
or U9520 (N_9520,N_5965,N_7306);
nand U9521 (N_9521,N_5395,N_5494);
nand U9522 (N_9522,N_6002,N_4093);
nand U9523 (N_9523,N_7111,N_4866);
or U9524 (N_9524,N_4308,N_6047);
xor U9525 (N_9525,N_6513,N_4364);
nand U9526 (N_9526,N_7536,N_5817);
or U9527 (N_9527,N_5124,N_7954);
nand U9528 (N_9528,N_7591,N_5238);
nor U9529 (N_9529,N_4697,N_4280);
or U9530 (N_9530,N_5682,N_4712);
or U9531 (N_9531,N_4267,N_4632);
nand U9532 (N_9532,N_6745,N_5071);
and U9533 (N_9533,N_7426,N_6241);
nor U9534 (N_9534,N_5467,N_6951);
nand U9535 (N_9535,N_7567,N_4319);
nand U9536 (N_9536,N_5114,N_5865);
or U9537 (N_9537,N_7920,N_5230);
nand U9538 (N_9538,N_7102,N_6357);
nor U9539 (N_9539,N_4708,N_5903);
and U9540 (N_9540,N_5438,N_5112);
nor U9541 (N_9541,N_5383,N_7778);
nand U9542 (N_9542,N_6136,N_4044);
nand U9543 (N_9543,N_7078,N_6530);
nor U9544 (N_9544,N_5934,N_4813);
nand U9545 (N_9545,N_4393,N_6596);
nand U9546 (N_9546,N_7429,N_6425);
nand U9547 (N_9547,N_5164,N_7839);
or U9548 (N_9548,N_7294,N_6994);
nand U9549 (N_9549,N_6540,N_4165);
or U9550 (N_9550,N_5622,N_4881);
nand U9551 (N_9551,N_5587,N_7131);
xor U9552 (N_9552,N_4687,N_4046);
nand U9553 (N_9553,N_6024,N_4275);
or U9554 (N_9554,N_5477,N_7705);
nor U9555 (N_9555,N_5356,N_5696);
and U9556 (N_9556,N_4038,N_7329);
nor U9557 (N_9557,N_4931,N_6588);
nor U9558 (N_9558,N_6935,N_6185);
and U9559 (N_9559,N_4522,N_4882);
or U9560 (N_9560,N_5312,N_6752);
nor U9561 (N_9561,N_5918,N_7451);
and U9562 (N_9562,N_5595,N_7538);
xnor U9563 (N_9563,N_7178,N_6942);
and U9564 (N_9564,N_7507,N_5501);
nor U9565 (N_9565,N_4332,N_5576);
nor U9566 (N_9566,N_5524,N_4570);
nand U9567 (N_9567,N_4123,N_7750);
and U9568 (N_9568,N_5978,N_4412);
or U9569 (N_9569,N_4877,N_5139);
and U9570 (N_9570,N_4685,N_5064);
nand U9571 (N_9571,N_6889,N_5374);
or U9572 (N_9572,N_7926,N_4490);
or U9573 (N_9573,N_6020,N_6683);
nor U9574 (N_9574,N_7903,N_6167);
or U9575 (N_9575,N_5286,N_7494);
or U9576 (N_9576,N_5527,N_7447);
and U9577 (N_9577,N_5652,N_5771);
nand U9578 (N_9578,N_6721,N_4011);
nand U9579 (N_9579,N_7860,N_7873);
nor U9580 (N_9580,N_4067,N_5154);
nor U9581 (N_9581,N_6923,N_7651);
and U9582 (N_9582,N_5745,N_7942);
and U9583 (N_9583,N_4889,N_6181);
nand U9584 (N_9584,N_5172,N_4515);
nand U9585 (N_9585,N_4609,N_5811);
and U9586 (N_9586,N_6737,N_6259);
nor U9587 (N_9587,N_6788,N_7574);
nor U9588 (N_9588,N_6142,N_5896);
nor U9589 (N_9589,N_4145,N_6316);
or U9590 (N_9590,N_7210,N_4748);
nand U9591 (N_9591,N_4018,N_5497);
nand U9592 (N_9592,N_7694,N_4061);
and U9593 (N_9593,N_4294,N_7142);
nor U9594 (N_9594,N_4036,N_4990);
and U9595 (N_9595,N_5226,N_5369);
or U9596 (N_9596,N_6875,N_4954);
nor U9597 (N_9597,N_7340,N_6497);
or U9598 (N_9598,N_5869,N_4476);
and U9599 (N_9599,N_6850,N_7378);
nand U9600 (N_9600,N_6891,N_5845);
or U9601 (N_9601,N_6678,N_4577);
and U9602 (N_9602,N_4713,N_6943);
nor U9603 (N_9603,N_6204,N_5216);
nand U9604 (N_9604,N_5110,N_4144);
or U9605 (N_9605,N_7973,N_5874);
or U9606 (N_9606,N_5772,N_4056);
nor U9607 (N_9607,N_6874,N_4806);
xnor U9608 (N_9608,N_4989,N_5660);
and U9609 (N_9609,N_4779,N_5352);
or U9610 (N_9610,N_6617,N_4726);
or U9611 (N_9611,N_5491,N_5141);
or U9612 (N_9612,N_5757,N_7326);
nor U9613 (N_9613,N_4912,N_7719);
nor U9614 (N_9614,N_5391,N_6229);
or U9615 (N_9615,N_4090,N_4546);
nor U9616 (N_9616,N_5821,N_4113);
nand U9617 (N_9617,N_4520,N_5773);
and U9618 (N_9618,N_6057,N_4050);
nand U9619 (N_9619,N_4328,N_5371);
or U9620 (N_9620,N_5675,N_7768);
and U9621 (N_9621,N_4358,N_4164);
nand U9622 (N_9622,N_5123,N_5073);
or U9623 (N_9623,N_7389,N_5938);
or U9624 (N_9624,N_7757,N_7898);
nor U9625 (N_9625,N_5547,N_5405);
or U9626 (N_9626,N_6623,N_4517);
or U9627 (N_9627,N_4993,N_5782);
and U9628 (N_9628,N_7784,N_6431);
or U9629 (N_9629,N_4385,N_7332);
nor U9630 (N_9630,N_7514,N_4361);
nor U9631 (N_9631,N_5334,N_6519);
nor U9632 (N_9632,N_6556,N_7560);
nand U9633 (N_9633,N_5198,N_6668);
nand U9634 (N_9634,N_7668,N_7746);
nand U9635 (N_9635,N_5469,N_6122);
or U9636 (N_9636,N_4142,N_7740);
or U9637 (N_9637,N_5555,N_5336);
and U9638 (N_9638,N_5133,N_5077);
nand U9639 (N_9639,N_5999,N_6795);
xor U9640 (N_9640,N_6360,N_4835);
or U9641 (N_9641,N_4589,N_6524);
and U9642 (N_9642,N_7177,N_7537);
nand U9643 (N_9643,N_5803,N_4906);
or U9644 (N_9644,N_5878,N_6263);
nand U9645 (N_9645,N_4885,N_4104);
nand U9646 (N_9646,N_4542,N_7446);
nand U9647 (N_9647,N_4017,N_7976);
and U9648 (N_9648,N_6129,N_7730);
nand U9649 (N_9649,N_5632,N_6340);
and U9650 (N_9650,N_5051,N_4896);
xor U9651 (N_9651,N_4664,N_7299);
nand U9652 (N_9652,N_4278,N_5440);
nand U9653 (N_9653,N_7240,N_4979);
or U9654 (N_9654,N_6876,N_5726);
nand U9655 (N_9655,N_6134,N_4236);
and U9656 (N_9656,N_7652,N_4009);
nor U9657 (N_9657,N_5966,N_6187);
nand U9658 (N_9658,N_7961,N_6354);
nand U9659 (N_9659,N_5724,N_5059);
nand U9660 (N_9660,N_7025,N_6364);
nand U9661 (N_9661,N_7938,N_6394);
nor U9662 (N_9662,N_4102,N_5282);
nand U9663 (N_9663,N_7199,N_6849);
nand U9664 (N_9664,N_5799,N_5237);
or U9665 (N_9665,N_4340,N_7212);
and U9666 (N_9666,N_6681,N_5200);
or U9667 (N_9667,N_7624,N_6622);
or U9668 (N_9668,N_4356,N_5529);
nor U9669 (N_9669,N_7372,N_5598);
nor U9670 (N_9670,N_7589,N_4519);
nor U9671 (N_9671,N_6280,N_4512);
nor U9672 (N_9672,N_4105,N_4073);
or U9673 (N_9673,N_5895,N_5208);
nor U9674 (N_9674,N_4414,N_5284);
or U9675 (N_9675,N_6575,N_7977);
nor U9676 (N_9676,N_7703,N_5258);
and U9677 (N_9677,N_7636,N_5332);
and U9678 (N_9678,N_5488,N_6387);
or U9679 (N_9679,N_7438,N_6342);
nor U9680 (N_9680,N_4730,N_5384);
nor U9681 (N_9681,N_4691,N_6841);
nand U9682 (N_9682,N_6894,N_7552);
nor U9683 (N_9683,N_7418,N_4149);
or U9684 (N_9684,N_4041,N_6361);
nand U9685 (N_9685,N_7578,N_6199);
or U9686 (N_9686,N_5425,N_5074);
or U9687 (N_9687,N_4028,N_4898);
or U9688 (N_9688,N_5430,N_4560);
or U9689 (N_9689,N_4952,N_4370);
nor U9690 (N_9690,N_4381,N_5278);
nor U9691 (N_9691,N_6934,N_4780);
and U9692 (N_9692,N_4095,N_4739);
nand U9693 (N_9693,N_6064,N_4228);
or U9694 (N_9694,N_5857,N_7262);
or U9695 (N_9695,N_4203,N_6051);
or U9696 (N_9696,N_6581,N_6797);
and U9697 (N_9697,N_4392,N_6848);
or U9698 (N_9698,N_6075,N_4065);
and U9699 (N_9699,N_5277,N_4933);
nor U9700 (N_9700,N_4701,N_6344);
nand U9701 (N_9701,N_7779,N_5565);
and U9702 (N_9702,N_4770,N_6108);
or U9703 (N_9703,N_6453,N_6038);
or U9704 (N_9704,N_7931,N_5683);
or U9705 (N_9705,N_4354,N_5950);
nor U9706 (N_9706,N_7003,N_4131);
nor U9707 (N_9707,N_4366,N_4494);
or U9708 (N_9708,N_4639,N_6629);
nor U9709 (N_9709,N_7864,N_4946);
nand U9710 (N_9710,N_4196,N_5603);
and U9711 (N_9711,N_4230,N_5902);
nand U9712 (N_9712,N_4998,N_6279);
nand U9713 (N_9713,N_5519,N_6642);
or U9714 (N_9714,N_4045,N_4012);
nand U9715 (N_9715,N_6583,N_4201);
or U9716 (N_9716,N_6886,N_7466);
nor U9717 (N_9717,N_7785,N_6348);
and U9718 (N_9718,N_5428,N_4464);
nor U9719 (N_9719,N_6238,N_7026);
or U9720 (N_9720,N_5146,N_5958);
nor U9721 (N_9721,N_5314,N_5463);
nand U9722 (N_9722,N_6806,N_5088);
or U9723 (N_9723,N_6548,N_7787);
or U9724 (N_9724,N_5791,N_4488);
nand U9725 (N_9725,N_5584,N_4399);
nand U9726 (N_9726,N_7837,N_7434);
and U9727 (N_9727,N_6015,N_4172);
or U9728 (N_9728,N_6704,N_4421);
and U9729 (N_9729,N_6686,N_5280);
and U9730 (N_9730,N_7170,N_7097);
nand U9731 (N_9731,N_7650,N_4930);
and U9732 (N_9732,N_7621,N_4461);
nor U9733 (N_9733,N_6825,N_7595);
and U9734 (N_9734,N_5272,N_6778);
nor U9735 (N_9735,N_5921,N_4285);
or U9736 (N_9736,N_5097,N_7423);
and U9737 (N_9737,N_6451,N_7854);
and U9738 (N_9738,N_7914,N_6473);
nor U9739 (N_9739,N_7523,N_6318);
nor U9740 (N_9740,N_6680,N_6836);
nor U9741 (N_9741,N_7756,N_6985);
nor U9742 (N_9742,N_4678,N_4223);
nor U9743 (N_9743,N_4470,N_6380);
or U9744 (N_9744,N_6926,N_7936);
nand U9745 (N_9745,N_5452,N_6506);
nand U9746 (N_9746,N_6723,N_6430);
nand U9747 (N_9747,N_6346,N_4176);
nand U9748 (N_9748,N_5212,N_6809);
nor U9749 (N_9749,N_6146,N_6978);
and U9750 (N_9750,N_6534,N_4195);
or U9751 (N_9751,N_5096,N_6732);
nor U9752 (N_9752,N_5135,N_4774);
xnor U9753 (N_9753,N_5100,N_6760);
and U9754 (N_9754,N_7371,N_7273);
nand U9755 (N_9755,N_5836,N_7887);
nand U9756 (N_9756,N_4590,N_5787);
or U9757 (N_9757,N_5422,N_4524);
nor U9758 (N_9758,N_7098,N_5012);
nor U9759 (N_9759,N_4305,N_5888);
or U9760 (N_9760,N_4791,N_6769);
or U9761 (N_9761,N_5102,N_6115);
and U9762 (N_9762,N_4907,N_7383);
or U9763 (N_9763,N_4644,N_6208);
and U9764 (N_9764,N_6407,N_5695);
and U9765 (N_9765,N_6538,N_7674);
nand U9766 (N_9766,N_6363,N_7060);
or U9767 (N_9767,N_6775,N_6171);
and U9768 (N_9768,N_5072,N_6422);
or U9769 (N_9769,N_4634,N_6264);
nor U9770 (N_9770,N_5546,N_5500);
nand U9771 (N_9771,N_6476,N_4157);
nand U9772 (N_9772,N_7108,N_6527);
nor U9773 (N_9773,N_6946,N_5455);
or U9774 (N_9774,N_5375,N_6025);
or U9775 (N_9775,N_5301,N_7106);
nand U9776 (N_9776,N_5233,N_6705);
nand U9777 (N_9777,N_6718,N_5482);
nand U9778 (N_9778,N_5485,N_6899);
and U9779 (N_9779,N_6192,N_6701);
and U9780 (N_9780,N_6783,N_7356);
nor U9781 (N_9781,N_4694,N_7835);
xnor U9782 (N_9782,N_5344,N_5876);
or U9783 (N_9783,N_7159,N_5777);
nor U9784 (N_9784,N_6579,N_5686);
nand U9785 (N_9785,N_5976,N_7314);
nand U9786 (N_9786,N_4006,N_4329);
nor U9787 (N_9787,N_7171,N_4373);
nor U9788 (N_9788,N_7733,N_5702);
or U9789 (N_9789,N_5026,N_4769);
nand U9790 (N_9790,N_7575,N_6356);
nand U9791 (N_9791,N_5194,N_4922);
nand U9792 (N_9792,N_6937,N_4874);
or U9793 (N_9793,N_7501,N_5872);
xor U9794 (N_9794,N_6861,N_7593);
nand U9795 (N_9795,N_5786,N_4915);
nand U9796 (N_9796,N_5163,N_7840);
nand U9797 (N_9797,N_4135,N_4007);
and U9798 (N_9798,N_4307,N_4369);
nor U9799 (N_9799,N_4911,N_5243);
or U9800 (N_9800,N_6275,N_4752);
and U9801 (N_9801,N_4472,N_4254);
nand U9802 (N_9802,N_6949,N_7728);
nand U9803 (N_9803,N_6442,N_5317);
nand U9804 (N_9804,N_6600,N_6369);
or U9805 (N_9805,N_7634,N_5916);
or U9806 (N_9806,N_5680,N_6843);
nand U9807 (N_9807,N_4829,N_5532);
and U9808 (N_9808,N_7465,N_7052);
or U9809 (N_9809,N_5672,N_5835);
or U9810 (N_9810,N_5577,N_4454);
nor U9811 (N_9811,N_4496,N_6672);
nand U9812 (N_9812,N_5089,N_4845);
nor U9813 (N_9813,N_6478,N_5489);
and U9814 (N_9814,N_4301,N_7010);
nand U9815 (N_9815,N_5092,N_7655);
and U9816 (N_9816,N_5122,N_5823);
and U9817 (N_9817,N_7704,N_5971);
nand U9818 (N_9818,N_7480,N_7399);
nand U9819 (N_9819,N_7123,N_7640);
nand U9820 (N_9820,N_6227,N_4872);
or U9821 (N_9821,N_5045,N_4088);
or U9822 (N_9822,N_5631,N_5638);
nor U9823 (N_9823,N_5006,N_7953);
nand U9824 (N_9824,N_5953,N_4800);
and U9825 (N_9825,N_6094,N_5179);
or U9826 (N_9826,N_7818,N_4764);
or U9827 (N_9827,N_6997,N_5677);
and U9828 (N_9828,N_5750,N_5846);
nor U9829 (N_9829,N_6885,N_7838);
nand U9830 (N_9830,N_4324,N_4282);
and U9831 (N_9831,N_4024,N_5130);
or U9832 (N_9832,N_7661,N_5767);
and U9833 (N_9833,N_5118,N_5926);
nor U9834 (N_9834,N_4181,N_7296);
nand U9835 (N_9835,N_6999,N_7441);
nand U9836 (N_9836,N_4311,N_4963);
nor U9837 (N_9837,N_7075,N_7702);
and U9838 (N_9838,N_6799,N_7211);
and U9839 (N_9839,N_7085,N_6612);
or U9840 (N_9840,N_5509,N_7450);
nand U9841 (N_9841,N_6503,N_7419);
nand U9842 (N_9842,N_5661,N_4072);
nand U9843 (N_9843,N_5099,N_7226);
and U9844 (N_9844,N_5231,N_6389);
nand U9845 (N_9845,N_6386,N_5673);
and U9846 (N_9846,N_4031,N_5742);
nor U9847 (N_9847,N_7775,N_6691);
nor U9848 (N_9848,N_4754,N_6953);
nor U9849 (N_9849,N_5697,N_6252);
or U9850 (N_9850,N_5169,N_6107);
or U9851 (N_9851,N_5396,N_5667);
nor U9852 (N_9852,N_4375,N_5015);
and U9853 (N_9853,N_5060,N_7191);
nor U9854 (N_9854,N_5190,N_7491);
nand U9855 (N_9855,N_4418,N_5034);
nand U9856 (N_9856,N_6489,N_6314);
nand U9857 (N_9857,N_5276,N_7225);
or U9858 (N_9858,N_6816,N_6358);
or U9859 (N_9859,N_6076,N_7220);
or U9860 (N_9860,N_7776,N_7209);
and U9861 (N_9861,N_4437,N_4397);
or U9862 (N_9862,N_4959,N_7113);
nor U9863 (N_9863,N_7394,N_5705);
nor U9864 (N_9864,N_7908,N_7149);
and U9865 (N_9865,N_5134,N_5871);
or U9866 (N_9866,N_7629,N_5850);
nor U9867 (N_9867,N_4202,N_7428);
or U9868 (N_9868,N_4506,N_7173);
and U9869 (N_9869,N_5915,N_5800);
nor U9870 (N_9870,N_7823,N_5610);
nor U9871 (N_9871,N_5685,N_5136);
and U9872 (N_9872,N_7834,N_4389);
and U9873 (N_9873,N_6814,N_5213);
or U9874 (N_9874,N_4859,N_7990);
nor U9875 (N_9875,N_4595,N_5549);
nand U9876 (N_9876,N_5600,N_7718);
or U9877 (N_9877,N_4502,N_5942);
nor U9878 (N_9878,N_5010,N_5217);
and U9879 (N_9879,N_4611,N_6621);
or U9880 (N_9880,N_5536,N_6539);
nor U9881 (N_9881,N_4032,N_4372);
or U9882 (N_9882,N_5681,N_6331);
and U9883 (N_9883,N_7440,N_5646);
nor U9884 (N_9884,N_5960,N_5197);
or U9885 (N_9885,N_7000,N_6470);
nor U9886 (N_9886,N_6971,N_5410);
nand U9887 (N_9887,N_4756,N_6321);
or U9888 (N_9888,N_7184,N_6837);
nor U9889 (N_9889,N_5070,N_4562);
nor U9890 (N_9890,N_6615,N_4303);
nand U9891 (N_9891,N_6972,N_6447);
and U9892 (N_9892,N_4023,N_5671);
or U9893 (N_9893,N_4207,N_7810);
nand U9894 (N_9894,N_6910,N_4773);
or U9895 (N_9895,N_6587,N_7363);
or U9896 (N_9896,N_4415,N_7259);
or U9897 (N_9897,N_6490,N_4100);
nor U9898 (N_9898,N_7833,N_6130);
and U9899 (N_9899,N_5056,N_4914);
nand U9900 (N_9900,N_4204,N_5349);
nor U9901 (N_9901,N_5990,N_7549);
or U9902 (N_9902,N_5792,N_7007);
and U9903 (N_9903,N_4086,N_4467);
nand U9904 (N_9904,N_7797,N_7584);
or U9905 (N_9905,N_6695,N_7459);
and U9906 (N_9906,N_5676,N_4913);
or U9907 (N_9907,N_7741,N_4058);
nor U9908 (N_9908,N_4599,N_6189);
or U9909 (N_9909,N_5699,N_6991);
and U9910 (N_9910,N_6304,N_5462);
nand U9911 (N_9911,N_5544,N_6172);
nor U9912 (N_9912,N_6822,N_5732);
and U9913 (N_9913,N_7282,N_6114);
and U9914 (N_9914,N_6458,N_7156);
and U9915 (N_9915,N_5735,N_7136);
and U9916 (N_9916,N_5086,N_5533);
or U9917 (N_9917,N_6089,N_7095);
nand U9918 (N_9918,N_5315,N_6474);
nor U9919 (N_9919,N_6215,N_7002);
or U9920 (N_9920,N_6631,N_7849);
or U9921 (N_9921,N_5625,N_5007);
nor U9922 (N_9922,N_5326,N_5590);
or U9923 (N_9923,N_6301,N_5556);
and U9924 (N_9924,N_6829,N_4347);
or U9925 (N_9925,N_6892,N_5299);
nand U9926 (N_9926,N_7825,N_5307);
and U9927 (N_9927,N_5721,N_6005);
or U9928 (N_9928,N_7543,N_4276);
nor U9929 (N_9929,N_5856,N_4409);
or U9930 (N_9930,N_4255,N_7691);
nor U9931 (N_9931,N_5923,N_5157);
or U9932 (N_9932,N_6618,N_5526);
or U9933 (N_9933,N_6211,N_5674);
or U9934 (N_9934,N_6243,N_6748);
nand U9935 (N_9935,N_5044,N_7338);
nor U9936 (N_9936,N_4927,N_7546);
nand U9937 (N_9937,N_4972,N_4854);
and U9938 (N_9938,N_6449,N_5783);
or U9939 (N_9939,N_6260,N_6794);
or U9940 (N_9940,N_7140,N_7660);
or U9941 (N_9941,N_6139,N_6852);
or U9942 (N_9942,N_7036,N_6086);
or U9943 (N_9943,N_7955,N_6433);
nor U9944 (N_9944,N_6550,N_5944);
nor U9945 (N_9945,N_4799,N_6606);
nand U9946 (N_9946,N_7617,N_4776);
and U9947 (N_9947,N_4256,N_5511);
nand U9948 (N_9948,N_7364,N_4141);
or U9949 (N_9949,N_5351,N_5293);
or U9950 (N_9950,N_4465,N_7522);
xor U9951 (N_9951,N_5708,N_6993);
nor U9952 (N_9952,N_6774,N_7622);
or U9953 (N_9953,N_6411,N_7346);
nand U9954 (N_9954,N_5502,N_6658);
nand U9955 (N_9955,N_4200,N_6333);
nor U9956 (N_9956,N_7397,N_7237);
nor U9957 (N_9957,N_6834,N_6472);
and U9958 (N_9958,N_5327,N_4110);
and U9959 (N_9959,N_6284,N_7722);
and U9960 (N_9960,N_6289,N_6805);
nor U9961 (N_9961,N_5935,N_7735);
nand U9962 (N_9962,N_7148,N_7659);
nand U9963 (N_9963,N_4700,N_6381);
and U9964 (N_9964,N_6582,N_5554);
and U9965 (N_9965,N_4648,N_6069);
nand U9966 (N_9966,N_6319,N_7246);
nand U9967 (N_9967,N_7035,N_6625);
or U9968 (N_9968,N_4573,N_4544);
or U9969 (N_9969,N_5036,N_4717);
nand U9970 (N_9970,N_5252,N_4623);
or U9971 (N_9971,N_7433,N_4021);
and U9972 (N_9972,N_5814,N_4420);
and U9973 (N_9973,N_5897,N_4220);
nor U9974 (N_9974,N_4501,N_7752);
nand U9975 (N_9975,N_4443,N_7369);
nand U9976 (N_9976,N_4224,N_5224);
or U9977 (N_9977,N_6307,N_6514);
nand U9978 (N_9978,N_5262,N_7278);
nand U9979 (N_9979,N_6960,N_6371);
nand U9980 (N_9980,N_6270,N_6237);
and U9981 (N_9981,N_4710,N_6784);
nor U9982 (N_9982,N_4961,N_7354);
or U9983 (N_9983,N_6766,N_5409);
or U9984 (N_9984,N_4988,N_6598);
nor U9985 (N_9985,N_7723,N_4298);
nand U9986 (N_9986,N_5709,N_4013);
nand U9987 (N_9987,N_4886,N_6533);
and U9988 (N_9988,N_6773,N_7766);
nand U9989 (N_9989,N_4798,N_5310);
or U9990 (N_9990,N_7377,N_6847);
nor U9991 (N_9991,N_5107,N_4548);
and U9992 (N_9992,N_6128,N_6959);
and U9993 (N_9993,N_6287,N_7913);
nand U9994 (N_9994,N_5716,N_5188);
nor U9995 (N_9995,N_5730,N_7997);
nor U9996 (N_9996,N_4205,N_6194);
or U9997 (N_9997,N_5812,N_4531);
or U9998 (N_9998,N_7845,N_5291);
nand U9999 (N_9999,N_4902,N_5664);
or U10000 (N_10000,N_4517,N_4238);
nand U10001 (N_10001,N_5356,N_7858);
nor U10002 (N_10002,N_7661,N_4984);
nand U10003 (N_10003,N_4327,N_5604);
nor U10004 (N_10004,N_5946,N_5657);
and U10005 (N_10005,N_5014,N_5365);
nor U10006 (N_10006,N_6533,N_5148);
nand U10007 (N_10007,N_5220,N_5437);
nand U10008 (N_10008,N_7049,N_5820);
nand U10009 (N_10009,N_7598,N_6833);
nand U10010 (N_10010,N_4453,N_7733);
nor U10011 (N_10011,N_7863,N_6529);
nand U10012 (N_10012,N_5092,N_4330);
and U10013 (N_10013,N_6998,N_6697);
and U10014 (N_10014,N_4265,N_7164);
or U10015 (N_10015,N_5898,N_7490);
nand U10016 (N_10016,N_5579,N_6260);
nor U10017 (N_10017,N_4127,N_5477);
or U10018 (N_10018,N_4125,N_6990);
and U10019 (N_10019,N_6049,N_5066);
and U10020 (N_10020,N_7134,N_4454);
and U10021 (N_10021,N_4086,N_4260);
and U10022 (N_10022,N_4578,N_6353);
or U10023 (N_10023,N_4686,N_5717);
nand U10024 (N_10024,N_4307,N_7150);
nand U10025 (N_10025,N_4080,N_5498);
or U10026 (N_10026,N_6573,N_5805);
or U10027 (N_10027,N_5839,N_4807);
or U10028 (N_10028,N_6018,N_7257);
nand U10029 (N_10029,N_6195,N_7214);
nor U10030 (N_10030,N_6599,N_5754);
nor U10031 (N_10031,N_7472,N_7261);
nor U10032 (N_10032,N_7502,N_4677);
or U10033 (N_10033,N_7021,N_4064);
nand U10034 (N_10034,N_7420,N_4567);
nand U10035 (N_10035,N_4048,N_6566);
nand U10036 (N_10036,N_5413,N_6215);
or U10037 (N_10037,N_6956,N_5750);
nor U10038 (N_10038,N_6664,N_4945);
or U10039 (N_10039,N_6252,N_6158);
nor U10040 (N_10040,N_4116,N_5022);
and U10041 (N_10041,N_4115,N_4311);
or U10042 (N_10042,N_6289,N_4284);
and U10043 (N_10043,N_6431,N_6343);
or U10044 (N_10044,N_4133,N_5234);
or U10045 (N_10045,N_5806,N_6152);
nor U10046 (N_10046,N_6891,N_4779);
nand U10047 (N_10047,N_4254,N_4933);
and U10048 (N_10048,N_4828,N_6130);
nor U10049 (N_10049,N_4750,N_5901);
and U10050 (N_10050,N_4410,N_6440);
nand U10051 (N_10051,N_7928,N_5351);
and U10052 (N_10052,N_7842,N_7889);
nand U10053 (N_10053,N_6794,N_6456);
and U10054 (N_10054,N_6259,N_6763);
nand U10055 (N_10055,N_7099,N_6962);
or U10056 (N_10056,N_6754,N_7590);
or U10057 (N_10057,N_5021,N_7938);
or U10058 (N_10058,N_7936,N_5852);
nor U10059 (N_10059,N_4411,N_4717);
nand U10060 (N_10060,N_4948,N_6753);
and U10061 (N_10061,N_5460,N_7964);
and U10062 (N_10062,N_7706,N_7264);
nor U10063 (N_10063,N_4826,N_4013);
and U10064 (N_10064,N_6624,N_7861);
or U10065 (N_10065,N_6780,N_7199);
and U10066 (N_10066,N_7025,N_4641);
or U10067 (N_10067,N_6500,N_5363);
nor U10068 (N_10068,N_6626,N_5378);
and U10069 (N_10069,N_5493,N_4974);
or U10070 (N_10070,N_6273,N_4679);
and U10071 (N_10071,N_6569,N_6846);
and U10072 (N_10072,N_4147,N_7274);
and U10073 (N_10073,N_5807,N_7208);
and U10074 (N_10074,N_4333,N_7382);
nand U10075 (N_10075,N_7999,N_5340);
nand U10076 (N_10076,N_6195,N_7735);
nand U10077 (N_10077,N_6887,N_4942);
or U10078 (N_10078,N_7422,N_4426);
nor U10079 (N_10079,N_7581,N_5636);
nand U10080 (N_10080,N_6552,N_7151);
nand U10081 (N_10081,N_4707,N_5684);
or U10082 (N_10082,N_4345,N_4364);
nand U10083 (N_10083,N_4372,N_5130);
or U10084 (N_10084,N_4838,N_5074);
or U10085 (N_10085,N_6569,N_7987);
and U10086 (N_10086,N_7894,N_6220);
nand U10087 (N_10087,N_4322,N_4134);
and U10088 (N_10088,N_4715,N_6660);
nor U10089 (N_10089,N_4990,N_6039);
or U10090 (N_10090,N_5684,N_5840);
and U10091 (N_10091,N_6502,N_7933);
nand U10092 (N_10092,N_7106,N_7805);
nor U10093 (N_10093,N_4242,N_7042);
nor U10094 (N_10094,N_5794,N_4499);
nand U10095 (N_10095,N_7598,N_4924);
and U10096 (N_10096,N_7569,N_6482);
and U10097 (N_10097,N_6337,N_5978);
nand U10098 (N_10098,N_4699,N_4918);
and U10099 (N_10099,N_7309,N_5371);
nand U10100 (N_10100,N_6073,N_7422);
nor U10101 (N_10101,N_4228,N_6017);
or U10102 (N_10102,N_6090,N_5634);
nor U10103 (N_10103,N_4740,N_5693);
nor U10104 (N_10104,N_5789,N_6690);
nor U10105 (N_10105,N_4773,N_4744);
and U10106 (N_10106,N_6439,N_5070);
and U10107 (N_10107,N_5490,N_5134);
or U10108 (N_10108,N_5195,N_4512);
nor U10109 (N_10109,N_4240,N_4229);
and U10110 (N_10110,N_7897,N_7723);
and U10111 (N_10111,N_5943,N_4600);
nand U10112 (N_10112,N_4665,N_4251);
nor U10113 (N_10113,N_4950,N_7313);
nor U10114 (N_10114,N_7659,N_5406);
nor U10115 (N_10115,N_5068,N_5924);
xor U10116 (N_10116,N_6679,N_5900);
nand U10117 (N_10117,N_7921,N_6726);
or U10118 (N_10118,N_5676,N_5154);
or U10119 (N_10119,N_4157,N_6431);
nand U10120 (N_10120,N_5009,N_4504);
nor U10121 (N_10121,N_7543,N_6703);
nor U10122 (N_10122,N_4493,N_7974);
nor U10123 (N_10123,N_4843,N_5183);
or U10124 (N_10124,N_6458,N_7628);
nand U10125 (N_10125,N_4236,N_6252);
nor U10126 (N_10126,N_5755,N_6165);
and U10127 (N_10127,N_5578,N_6957);
nor U10128 (N_10128,N_6667,N_5973);
nor U10129 (N_10129,N_6345,N_4230);
or U10130 (N_10130,N_7459,N_6497);
and U10131 (N_10131,N_7448,N_6183);
nor U10132 (N_10132,N_6253,N_5228);
or U10133 (N_10133,N_5863,N_5128);
and U10134 (N_10134,N_5307,N_5408);
nand U10135 (N_10135,N_6086,N_5442);
nand U10136 (N_10136,N_4910,N_5455);
or U10137 (N_10137,N_5798,N_7292);
xor U10138 (N_10138,N_5178,N_4798);
nor U10139 (N_10139,N_4063,N_4161);
nand U10140 (N_10140,N_5745,N_7252);
nor U10141 (N_10141,N_4515,N_5426);
nand U10142 (N_10142,N_4543,N_6117);
and U10143 (N_10143,N_5609,N_5687);
and U10144 (N_10144,N_4321,N_5074);
and U10145 (N_10145,N_6354,N_6189);
nor U10146 (N_10146,N_7601,N_6122);
nand U10147 (N_10147,N_4968,N_4455);
or U10148 (N_10148,N_5457,N_7982);
and U10149 (N_10149,N_4304,N_7418);
and U10150 (N_10150,N_6892,N_5961);
nand U10151 (N_10151,N_7793,N_7233);
nor U10152 (N_10152,N_6412,N_7436);
or U10153 (N_10153,N_5721,N_5620);
and U10154 (N_10154,N_5944,N_5872);
nor U10155 (N_10155,N_7470,N_7737);
or U10156 (N_10156,N_5551,N_4695);
nand U10157 (N_10157,N_5554,N_5699);
xnor U10158 (N_10158,N_4753,N_6466);
and U10159 (N_10159,N_7201,N_5450);
or U10160 (N_10160,N_4810,N_7288);
nand U10161 (N_10161,N_6690,N_5501);
or U10162 (N_10162,N_6268,N_7912);
nand U10163 (N_10163,N_7525,N_6124);
nor U10164 (N_10164,N_5614,N_4772);
and U10165 (N_10165,N_7788,N_5137);
nor U10166 (N_10166,N_7383,N_6779);
nand U10167 (N_10167,N_7745,N_5513);
nand U10168 (N_10168,N_6186,N_5831);
and U10169 (N_10169,N_7098,N_7532);
or U10170 (N_10170,N_4770,N_4005);
nand U10171 (N_10171,N_7418,N_6539);
nand U10172 (N_10172,N_7524,N_5000);
nand U10173 (N_10173,N_5747,N_6986);
or U10174 (N_10174,N_7815,N_6889);
and U10175 (N_10175,N_4408,N_4485);
or U10176 (N_10176,N_5891,N_6074);
nor U10177 (N_10177,N_5119,N_4770);
or U10178 (N_10178,N_6896,N_6985);
and U10179 (N_10179,N_7575,N_5336);
nand U10180 (N_10180,N_6503,N_7069);
or U10181 (N_10181,N_5337,N_4361);
nand U10182 (N_10182,N_4554,N_5222);
nand U10183 (N_10183,N_7842,N_5079);
nand U10184 (N_10184,N_5981,N_5360);
or U10185 (N_10185,N_5168,N_7258);
nand U10186 (N_10186,N_7099,N_4407);
or U10187 (N_10187,N_4540,N_7921);
or U10188 (N_10188,N_7454,N_6697);
and U10189 (N_10189,N_7930,N_6094);
nor U10190 (N_10190,N_7460,N_4456);
nand U10191 (N_10191,N_7491,N_4747);
and U10192 (N_10192,N_7480,N_7171);
or U10193 (N_10193,N_5315,N_7668);
and U10194 (N_10194,N_4875,N_5804);
and U10195 (N_10195,N_4577,N_6547);
and U10196 (N_10196,N_7475,N_4759);
or U10197 (N_10197,N_7537,N_7308);
nand U10198 (N_10198,N_6286,N_7483);
nand U10199 (N_10199,N_6678,N_5007);
or U10200 (N_10200,N_5469,N_5738);
and U10201 (N_10201,N_4005,N_7694);
nor U10202 (N_10202,N_6052,N_6096);
and U10203 (N_10203,N_5955,N_7424);
and U10204 (N_10204,N_5969,N_5188);
nand U10205 (N_10205,N_4583,N_7716);
nand U10206 (N_10206,N_4490,N_6027);
or U10207 (N_10207,N_4348,N_4766);
and U10208 (N_10208,N_6201,N_7291);
and U10209 (N_10209,N_7289,N_4926);
or U10210 (N_10210,N_4892,N_4938);
or U10211 (N_10211,N_6925,N_4493);
and U10212 (N_10212,N_5177,N_4869);
nand U10213 (N_10213,N_7101,N_4847);
nor U10214 (N_10214,N_5616,N_5251);
and U10215 (N_10215,N_7703,N_4587);
nor U10216 (N_10216,N_7120,N_5679);
or U10217 (N_10217,N_5685,N_6640);
or U10218 (N_10218,N_7106,N_5275);
nor U10219 (N_10219,N_6628,N_6087);
and U10220 (N_10220,N_4643,N_4121);
or U10221 (N_10221,N_4988,N_4868);
nor U10222 (N_10222,N_7606,N_5510);
nand U10223 (N_10223,N_6065,N_6570);
and U10224 (N_10224,N_4282,N_4400);
and U10225 (N_10225,N_7044,N_5577);
or U10226 (N_10226,N_5090,N_5552);
nor U10227 (N_10227,N_4769,N_7439);
or U10228 (N_10228,N_7717,N_5304);
or U10229 (N_10229,N_4696,N_7388);
or U10230 (N_10230,N_6483,N_4345);
nor U10231 (N_10231,N_6175,N_6242);
nand U10232 (N_10232,N_6004,N_6894);
nand U10233 (N_10233,N_4078,N_6637);
or U10234 (N_10234,N_7048,N_4702);
or U10235 (N_10235,N_5424,N_5954);
nor U10236 (N_10236,N_7109,N_5267);
or U10237 (N_10237,N_7947,N_5723);
or U10238 (N_10238,N_5430,N_5516);
or U10239 (N_10239,N_5030,N_6552);
or U10240 (N_10240,N_6113,N_4413);
and U10241 (N_10241,N_4787,N_5780);
and U10242 (N_10242,N_6838,N_6925);
and U10243 (N_10243,N_5821,N_5092);
and U10244 (N_10244,N_4384,N_5393);
nand U10245 (N_10245,N_7168,N_4925);
nor U10246 (N_10246,N_4523,N_6393);
and U10247 (N_10247,N_5955,N_4966);
nor U10248 (N_10248,N_6128,N_4890);
or U10249 (N_10249,N_5486,N_7844);
nand U10250 (N_10250,N_4249,N_4751);
and U10251 (N_10251,N_6175,N_6008);
nand U10252 (N_10252,N_6395,N_5605);
nor U10253 (N_10253,N_7431,N_5589);
and U10254 (N_10254,N_5253,N_5769);
nor U10255 (N_10255,N_6676,N_5124);
nand U10256 (N_10256,N_6405,N_7618);
nand U10257 (N_10257,N_6038,N_7344);
and U10258 (N_10258,N_6183,N_7912);
nand U10259 (N_10259,N_7616,N_7891);
or U10260 (N_10260,N_6652,N_5938);
nand U10261 (N_10261,N_6372,N_5165);
nand U10262 (N_10262,N_7172,N_4347);
nor U10263 (N_10263,N_4426,N_6519);
and U10264 (N_10264,N_6744,N_6300);
nor U10265 (N_10265,N_5985,N_6200);
or U10266 (N_10266,N_6036,N_4135);
nor U10267 (N_10267,N_6990,N_4285);
or U10268 (N_10268,N_7482,N_7663);
nand U10269 (N_10269,N_7313,N_5526);
nor U10270 (N_10270,N_5323,N_5905);
nand U10271 (N_10271,N_6762,N_6139);
or U10272 (N_10272,N_4425,N_4147);
nor U10273 (N_10273,N_6552,N_5601);
or U10274 (N_10274,N_6038,N_6905);
and U10275 (N_10275,N_7400,N_7600);
and U10276 (N_10276,N_6327,N_6792);
nor U10277 (N_10277,N_5864,N_6032);
and U10278 (N_10278,N_5090,N_5906);
xor U10279 (N_10279,N_4171,N_4985);
and U10280 (N_10280,N_6025,N_6469);
nand U10281 (N_10281,N_7953,N_6256);
or U10282 (N_10282,N_5314,N_6878);
nor U10283 (N_10283,N_6029,N_6607);
and U10284 (N_10284,N_6121,N_6257);
or U10285 (N_10285,N_7036,N_6791);
nor U10286 (N_10286,N_4196,N_4172);
or U10287 (N_10287,N_4545,N_6201);
nor U10288 (N_10288,N_6083,N_5145);
xor U10289 (N_10289,N_6705,N_5161);
and U10290 (N_10290,N_5111,N_6374);
xnor U10291 (N_10291,N_6084,N_4029);
or U10292 (N_10292,N_5817,N_5183);
nand U10293 (N_10293,N_4315,N_7528);
nand U10294 (N_10294,N_4899,N_7310);
nor U10295 (N_10295,N_7410,N_7554);
and U10296 (N_10296,N_4673,N_6479);
nor U10297 (N_10297,N_4105,N_5451);
nand U10298 (N_10298,N_7994,N_7149);
nor U10299 (N_10299,N_7012,N_5165);
or U10300 (N_10300,N_6181,N_6071);
or U10301 (N_10301,N_4474,N_5222);
nand U10302 (N_10302,N_6330,N_4700);
nand U10303 (N_10303,N_6172,N_6472);
and U10304 (N_10304,N_6953,N_6544);
and U10305 (N_10305,N_7576,N_5024);
or U10306 (N_10306,N_4520,N_6462);
nor U10307 (N_10307,N_6387,N_4207);
and U10308 (N_10308,N_4864,N_6192);
nor U10309 (N_10309,N_6444,N_5647);
and U10310 (N_10310,N_6984,N_6616);
or U10311 (N_10311,N_5903,N_5321);
and U10312 (N_10312,N_4129,N_4118);
nand U10313 (N_10313,N_4749,N_6116);
nand U10314 (N_10314,N_5460,N_5268);
or U10315 (N_10315,N_4228,N_6074);
or U10316 (N_10316,N_6251,N_6213);
nand U10317 (N_10317,N_7522,N_6486);
and U10318 (N_10318,N_7915,N_4385);
nand U10319 (N_10319,N_4741,N_4395);
nor U10320 (N_10320,N_4079,N_4048);
and U10321 (N_10321,N_7475,N_5943);
and U10322 (N_10322,N_4492,N_7488);
and U10323 (N_10323,N_6500,N_6841);
and U10324 (N_10324,N_6186,N_5079);
or U10325 (N_10325,N_7139,N_6987);
nand U10326 (N_10326,N_6243,N_4058);
or U10327 (N_10327,N_7979,N_4913);
nand U10328 (N_10328,N_4829,N_4816);
and U10329 (N_10329,N_4844,N_4366);
nor U10330 (N_10330,N_6103,N_4498);
and U10331 (N_10331,N_7127,N_4494);
and U10332 (N_10332,N_4060,N_5803);
nand U10333 (N_10333,N_4288,N_4641);
and U10334 (N_10334,N_7979,N_7989);
nor U10335 (N_10335,N_4848,N_6015);
nand U10336 (N_10336,N_7167,N_4774);
nor U10337 (N_10337,N_6893,N_5801);
or U10338 (N_10338,N_7554,N_7933);
or U10339 (N_10339,N_5096,N_7848);
nand U10340 (N_10340,N_5567,N_5624);
or U10341 (N_10341,N_5067,N_4997);
or U10342 (N_10342,N_4250,N_6411);
and U10343 (N_10343,N_5391,N_5685);
and U10344 (N_10344,N_4682,N_4950);
or U10345 (N_10345,N_5242,N_6789);
nand U10346 (N_10346,N_4081,N_7491);
and U10347 (N_10347,N_5850,N_4537);
or U10348 (N_10348,N_5287,N_4783);
or U10349 (N_10349,N_5052,N_6370);
or U10350 (N_10350,N_7934,N_6390);
nand U10351 (N_10351,N_6711,N_4125);
nand U10352 (N_10352,N_6204,N_7738);
nand U10353 (N_10353,N_4119,N_6299);
nor U10354 (N_10354,N_5026,N_5440);
nand U10355 (N_10355,N_4946,N_5072);
nand U10356 (N_10356,N_7425,N_5438);
nor U10357 (N_10357,N_4323,N_7562);
or U10358 (N_10358,N_7696,N_6122);
nand U10359 (N_10359,N_6552,N_4851);
and U10360 (N_10360,N_7416,N_6043);
nor U10361 (N_10361,N_6851,N_4566);
nand U10362 (N_10362,N_5847,N_4516);
nor U10363 (N_10363,N_6224,N_5370);
and U10364 (N_10364,N_7227,N_7426);
and U10365 (N_10365,N_4027,N_4646);
nor U10366 (N_10366,N_7295,N_7430);
or U10367 (N_10367,N_5173,N_4693);
nor U10368 (N_10368,N_7133,N_5019);
nand U10369 (N_10369,N_5032,N_4824);
nor U10370 (N_10370,N_5385,N_7908);
nand U10371 (N_10371,N_5700,N_4754);
or U10372 (N_10372,N_5029,N_7114);
and U10373 (N_10373,N_5935,N_5640);
nor U10374 (N_10374,N_5038,N_6564);
nand U10375 (N_10375,N_4275,N_7381);
and U10376 (N_10376,N_6246,N_4245);
and U10377 (N_10377,N_4629,N_4317);
nor U10378 (N_10378,N_7235,N_6656);
or U10379 (N_10379,N_4807,N_5528);
nand U10380 (N_10380,N_7728,N_6824);
nor U10381 (N_10381,N_6348,N_6774);
and U10382 (N_10382,N_7086,N_5275);
nand U10383 (N_10383,N_5665,N_5810);
nand U10384 (N_10384,N_7773,N_7188);
or U10385 (N_10385,N_4977,N_6769);
nor U10386 (N_10386,N_7729,N_4334);
nor U10387 (N_10387,N_7615,N_6756);
or U10388 (N_10388,N_5265,N_4822);
and U10389 (N_10389,N_7509,N_5327);
nand U10390 (N_10390,N_4127,N_7939);
nand U10391 (N_10391,N_4310,N_4583);
and U10392 (N_10392,N_5343,N_5101);
nand U10393 (N_10393,N_5648,N_6421);
nand U10394 (N_10394,N_7379,N_5636);
nand U10395 (N_10395,N_6778,N_7697);
or U10396 (N_10396,N_6326,N_4377);
nor U10397 (N_10397,N_5009,N_4591);
nor U10398 (N_10398,N_5044,N_7198);
nor U10399 (N_10399,N_7472,N_7492);
and U10400 (N_10400,N_7871,N_5434);
nand U10401 (N_10401,N_5266,N_6456);
nor U10402 (N_10402,N_6763,N_4127);
and U10403 (N_10403,N_6172,N_5411);
and U10404 (N_10404,N_4078,N_4523);
or U10405 (N_10405,N_4982,N_7547);
or U10406 (N_10406,N_6283,N_6036);
or U10407 (N_10407,N_5280,N_6491);
or U10408 (N_10408,N_6723,N_6234);
or U10409 (N_10409,N_4727,N_7850);
nand U10410 (N_10410,N_5343,N_4308);
nor U10411 (N_10411,N_5979,N_5971);
nand U10412 (N_10412,N_7389,N_4631);
nand U10413 (N_10413,N_4615,N_7376);
or U10414 (N_10414,N_7956,N_5909);
nand U10415 (N_10415,N_7084,N_7703);
or U10416 (N_10416,N_7259,N_5423);
nand U10417 (N_10417,N_4860,N_4396);
nor U10418 (N_10418,N_6680,N_5814);
or U10419 (N_10419,N_7088,N_5417);
or U10420 (N_10420,N_5083,N_4305);
nor U10421 (N_10421,N_5959,N_5968);
nor U10422 (N_10422,N_4103,N_7553);
nand U10423 (N_10423,N_4156,N_5247);
and U10424 (N_10424,N_7181,N_7920);
and U10425 (N_10425,N_5401,N_5613);
or U10426 (N_10426,N_5028,N_7692);
and U10427 (N_10427,N_6132,N_7427);
and U10428 (N_10428,N_4661,N_7586);
or U10429 (N_10429,N_6412,N_6989);
nor U10430 (N_10430,N_7780,N_5742);
and U10431 (N_10431,N_7083,N_7952);
and U10432 (N_10432,N_4887,N_6124);
nand U10433 (N_10433,N_7673,N_7048);
nor U10434 (N_10434,N_4185,N_5952);
nand U10435 (N_10435,N_4377,N_5335);
nor U10436 (N_10436,N_6413,N_7634);
nand U10437 (N_10437,N_6440,N_4207);
and U10438 (N_10438,N_6854,N_4975);
nand U10439 (N_10439,N_4284,N_5540);
and U10440 (N_10440,N_5015,N_4290);
nand U10441 (N_10441,N_6297,N_6759);
nand U10442 (N_10442,N_5822,N_7121);
nor U10443 (N_10443,N_4314,N_6918);
nor U10444 (N_10444,N_6306,N_4858);
or U10445 (N_10445,N_5064,N_7217);
and U10446 (N_10446,N_5214,N_4079);
or U10447 (N_10447,N_6334,N_4325);
and U10448 (N_10448,N_5389,N_5422);
and U10449 (N_10449,N_4773,N_6995);
nor U10450 (N_10450,N_4483,N_6540);
or U10451 (N_10451,N_7787,N_4078);
nor U10452 (N_10452,N_7545,N_6513);
nand U10453 (N_10453,N_7735,N_6792);
nor U10454 (N_10454,N_5703,N_7106);
or U10455 (N_10455,N_7900,N_5756);
nor U10456 (N_10456,N_4318,N_6034);
nor U10457 (N_10457,N_5356,N_5261);
nand U10458 (N_10458,N_7708,N_5911);
nand U10459 (N_10459,N_6976,N_7346);
or U10460 (N_10460,N_4971,N_6836);
nor U10461 (N_10461,N_4119,N_5127);
nand U10462 (N_10462,N_6079,N_7915);
and U10463 (N_10463,N_7560,N_7408);
nor U10464 (N_10464,N_5931,N_6791);
or U10465 (N_10465,N_4915,N_5938);
nor U10466 (N_10466,N_7789,N_6844);
or U10467 (N_10467,N_5918,N_5767);
and U10468 (N_10468,N_5557,N_6497);
nand U10469 (N_10469,N_6883,N_6866);
nand U10470 (N_10470,N_4569,N_6970);
and U10471 (N_10471,N_6219,N_7773);
nand U10472 (N_10472,N_6118,N_7285);
nor U10473 (N_10473,N_7174,N_5430);
nor U10474 (N_10474,N_5587,N_4739);
nand U10475 (N_10475,N_5992,N_6152);
nand U10476 (N_10476,N_6142,N_5490);
nor U10477 (N_10477,N_5406,N_6770);
nand U10478 (N_10478,N_7898,N_7387);
and U10479 (N_10479,N_4672,N_4584);
nand U10480 (N_10480,N_5926,N_4944);
nand U10481 (N_10481,N_6449,N_7281);
and U10482 (N_10482,N_6987,N_4846);
nor U10483 (N_10483,N_4333,N_4585);
xor U10484 (N_10484,N_7822,N_4156);
and U10485 (N_10485,N_4930,N_5506);
and U10486 (N_10486,N_6153,N_7526);
nor U10487 (N_10487,N_7289,N_7415);
and U10488 (N_10488,N_7719,N_7369);
and U10489 (N_10489,N_6456,N_4194);
nor U10490 (N_10490,N_5956,N_4128);
nor U10491 (N_10491,N_7889,N_5978);
or U10492 (N_10492,N_5085,N_4582);
and U10493 (N_10493,N_7972,N_6925);
or U10494 (N_10494,N_5064,N_4452);
or U10495 (N_10495,N_4508,N_5976);
or U10496 (N_10496,N_5002,N_6444);
or U10497 (N_10497,N_4036,N_6718);
and U10498 (N_10498,N_4685,N_4921);
nand U10499 (N_10499,N_4575,N_6197);
nand U10500 (N_10500,N_5389,N_4863);
nor U10501 (N_10501,N_6679,N_6062);
nor U10502 (N_10502,N_6030,N_4881);
nand U10503 (N_10503,N_6866,N_4264);
and U10504 (N_10504,N_4359,N_4707);
nand U10505 (N_10505,N_7839,N_7045);
or U10506 (N_10506,N_7204,N_6783);
and U10507 (N_10507,N_7366,N_5372);
nor U10508 (N_10508,N_4265,N_5281);
or U10509 (N_10509,N_5945,N_4119);
or U10510 (N_10510,N_4473,N_5793);
and U10511 (N_10511,N_6516,N_4175);
nand U10512 (N_10512,N_4239,N_7082);
nor U10513 (N_10513,N_7010,N_5560);
nor U10514 (N_10514,N_7953,N_7733);
nand U10515 (N_10515,N_4867,N_6563);
nand U10516 (N_10516,N_7982,N_7045);
or U10517 (N_10517,N_5310,N_4194);
or U10518 (N_10518,N_7012,N_5534);
xnor U10519 (N_10519,N_7125,N_5537);
or U10520 (N_10520,N_7779,N_7401);
and U10521 (N_10521,N_5624,N_4306);
or U10522 (N_10522,N_7795,N_4756);
or U10523 (N_10523,N_4774,N_5895);
nand U10524 (N_10524,N_7733,N_6807);
nor U10525 (N_10525,N_7435,N_4073);
nand U10526 (N_10526,N_4520,N_4786);
or U10527 (N_10527,N_7257,N_5189);
nor U10528 (N_10528,N_6714,N_7393);
nand U10529 (N_10529,N_7633,N_6079);
and U10530 (N_10530,N_6358,N_5268);
nand U10531 (N_10531,N_7969,N_7878);
nor U10532 (N_10532,N_4844,N_4442);
nor U10533 (N_10533,N_6148,N_5150);
nand U10534 (N_10534,N_7711,N_6391);
nor U10535 (N_10535,N_5951,N_7223);
nand U10536 (N_10536,N_4722,N_6904);
and U10537 (N_10537,N_4089,N_6031);
nor U10538 (N_10538,N_7417,N_5044);
or U10539 (N_10539,N_6851,N_7025);
and U10540 (N_10540,N_5981,N_7011);
nor U10541 (N_10541,N_4277,N_5555);
and U10542 (N_10542,N_7564,N_7327);
and U10543 (N_10543,N_5616,N_5534);
nand U10544 (N_10544,N_4791,N_6676);
nor U10545 (N_10545,N_4315,N_5297);
and U10546 (N_10546,N_5805,N_7502);
nor U10547 (N_10547,N_4950,N_4244);
nor U10548 (N_10548,N_5776,N_6801);
and U10549 (N_10549,N_6008,N_4240);
and U10550 (N_10550,N_5150,N_5370);
or U10551 (N_10551,N_7094,N_7307);
nor U10552 (N_10552,N_5355,N_4431);
nor U10553 (N_10553,N_7236,N_5904);
nand U10554 (N_10554,N_5262,N_5427);
or U10555 (N_10555,N_4005,N_7705);
nor U10556 (N_10556,N_5233,N_7242);
nor U10557 (N_10557,N_7482,N_5984);
nand U10558 (N_10558,N_5439,N_6871);
or U10559 (N_10559,N_7924,N_5210);
nand U10560 (N_10560,N_7184,N_7419);
or U10561 (N_10561,N_4259,N_5732);
or U10562 (N_10562,N_5111,N_4439);
and U10563 (N_10563,N_6773,N_6668);
nand U10564 (N_10564,N_7371,N_7731);
nor U10565 (N_10565,N_6589,N_5106);
nor U10566 (N_10566,N_4322,N_6708);
or U10567 (N_10567,N_5083,N_4281);
or U10568 (N_10568,N_4947,N_5575);
nor U10569 (N_10569,N_4226,N_7658);
or U10570 (N_10570,N_4389,N_7493);
nand U10571 (N_10571,N_4422,N_7075);
nor U10572 (N_10572,N_7935,N_4216);
nand U10573 (N_10573,N_5564,N_7389);
nor U10574 (N_10574,N_7651,N_7354);
nand U10575 (N_10575,N_6247,N_6972);
nand U10576 (N_10576,N_7940,N_4617);
nor U10577 (N_10577,N_4409,N_4331);
or U10578 (N_10578,N_4208,N_5520);
or U10579 (N_10579,N_7666,N_4198);
nor U10580 (N_10580,N_4118,N_5872);
nand U10581 (N_10581,N_4552,N_5790);
nand U10582 (N_10582,N_5888,N_7610);
nor U10583 (N_10583,N_7658,N_5568);
nand U10584 (N_10584,N_5212,N_7364);
nor U10585 (N_10585,N_7481,N_7294);
nor U10586 (N_10586,N_5381,N_4537);
or U10587 (N_10587,N_6140,N_5896);
or U10588 (N_10588,N_6813,N_5414);
nand U10589 (N_10589,N_5865,N_6199);
nor U10590 (N_10590,N_4595,N_6243);
or U10591 (N_10591,N_4699,N_6419);
nor U10592 (N_10592,N_4953,N_6462);
or U10593 (N_10593,N_7679,N_4945);
or U10594 (N_10594,N_4707,N_7503);
and U10595 (N_10595,N_5309,N_5623);
and U10596 (N_10596,N_5797,N_7870);
or U10597 (N_10597,N_6791,N_7093);
nor U10598 (N_10598,N_6669,N_7926);
or U10599 (N_10599,N_7297,N_7010);
and U10600 (N_10600,N_4591,N_4552);
or U10601 (N_10601,N_5118,N_4143);
or U10602 (N_10602,N_6968,N_5376);
and U10603 (N_10603,N_5367,N_4091);
and U10604 (N_10604,N_5785,N_5450);
or U10605 (N_10605,N_7628,N_6535);
nor U10606 (N_10606,N_7130,N_7413);
nand U10607 (N_10607,N_4414,N_6068);
nor U10608 (N_10608,N_5076,N_6759);
and U10609 (N_10609,N_4762,N_5180);
or U10610 (N_10610,N_7382,N_7333);
or U10611 (N_10611,N_4618,N_7376);
and U10612 (N_10612,N_7154,N_5881);
nor U10613 (N_10613,N_4888,N_5837);
or U10614 (N_10614,N_7410,N_4575);
or U10615 (N_10615,N_6531,N_6766);
and U10616 (N_10616,N_4708,N_5290);
nor U10617 (N_10617,N_7099,N_7968);
or U10618 (N_10618,N_4784,N_6295);
nor U10619 (N_10619,N_6706,N_6424);
nor U10620 (N_10620,N_7285,N_4068);
or U10621 (N_10621,N_4391,N_6671);
nand U10622 (N_10622,N_4282,N_5070);
and U10623 (N_10623,N_5407,N_7668);
or U10624 (N_10624,N_5616,N_4934);
nand U10625 (N_10625,N_6784,N_6254);
or U10626 (N_10626,N_7098,N_7576);
or U10627 (N_10627,N_4051,N_7146);
and U10628 (N_10628,N_4985,N_5280);
nor U10629 (N_10629,N_4289,N_6662);
nor U10630 (N_10630,N_4667,N_7213);
nand U10631 (N_10631,N_4187,N_5750);
nand U10632 (N_10632,N_5429,N_4735);
nor U10633 (N_10633,N_6782,N_6396);
nand U10634 (N_10634,N_6847,N_5849);
and U10635 (N_10635,N_7286,N_4188);
nand U10636 (N_10636,N_7106,N_7463);
nand U10637 (N_10637,N_4927,N_6269);
and U10638 (N_10638,N_7667,N_7812);
and U10639 (N_10639,N_7944,N_7184);
or U10640 (N_10640,N_6301,N_5238);
and U10641 (N_10641,N_7200,N_5901);
and U10642 (N_10642,N_7158,N_6954);
nand U10643 (N_10643,N_7530,N_5023);
or U10644 (N_10644,N_7875,N_4922);
nor U10645 (N_10645,N_4591,N_4770);
nand U10646 (N_10646,N_5737,N_4190);
or U10647 (N_10647,N_7694,N_6129);
and U10648 (N_10648,N_5987,N_6024);
nand U10649 (N_10649,N_7846,N_7917);
nor U10650 (N_10650,N_7395,N_4924);
nand U10651 (N_10651,N_7824,N_6524);
or U10652 (N_10652,N_5986,N_4423);
nor U10653 (N_10653,N_7902,N_6269);
or U10654 (N_10654,N_4832,N_7831);
and U10655 (N_10655,N_7540,N_6395);
nor U10656 (N_10656,N_5242,N_6931);
nor U10657 (N_10657,N_7796,N_6911);
or U10658 (N_10658,N_4020,N_6577);
or U10659 (N_10659,N_4553,N_7527);
or U10660 (N_10660,N_7662,N_7859);
and U10661 (N_10661,N_7919,N_4713);
or U10662 (N_10662,N_7247,N_5370);
nand U10663 (N_10663,N_7076,N_6178);
nand U10664 (N_10664,N_6997,N_7195);
and U10665 (N_10665,N_4308,N_6413);
nand U10666 (N_10666,N_7291,N_5001);
nand U10667 (N_10667,N_7505,N_7589);
nor U10668 (N_10668,N_5870,N_6242);
nand U10669 (N_10669,N_7775,N_7794);
or U10670 (N_10670,N_5226,N_7973);
nor U10671 (N_10671,N_6337,N_4320);
nor U10672 (N_10672,N_6966,N_4385);
or U10673 (N_10673,N_6254,N_6807);
or U10674 (N_10674,N_4290,N_4640);
nor U10675 (N_10675,N_5839,N_6530);
nand U10676 (N_10676,N_5267,N_4546);
nor U10677 (N_10677,N_4563,N_7782);
nor U10678 (N_10678,N_6808,N_4242);
nand U10679 (N_10679,N_5967,N_5348);
nor U10680 (N_10680,N_4468,N_4187);
or U10681 (N_10681,N_5152,N_7093);
nor U10682 (N_10682,N_4433,N_6304);
and U10683 (N_10683,N_6352,N_7304);
nor U10684 (N_10684,N_7271,N_6542);
nand U10685 (N_10685,N_6565,N_6096);
or U10686 (N_10686,N_7789,N_5894);
nor U10687 (N_10687,N_6408,N_5436);
or U10688 (N_10688,N_7948,N_5666);
nand U10689 (N_10689,N_7324,N_6090);
nor U10690 (N_10690,N_5860,N_4767);
nor U10691 (N_10691,N_4247,N_4874);
or U10692 (N_10692,N_7241,N_7951);
nand U10693 (N_10693,N_4624,N_4941);
nand U10694 (N_10694,N_6377,N_5514);
and U10695 (N_10695,N_6111,N_4006);
and U10696 (N_10696,N_7466,N_6269);
or U10697 (N_10697,N_6789,N_6727);
nor U10698 (N_10698,N_7601,N_7877);
and U10699 (N_10699,N_7931,N_4520);
nor U10700 (N_10700,N_7424,N_5597);
nand U10701 (N_10701,N_6740,N_6050);
and U10702 (N_10702,N_5873,N_5506);
nor U10703 (N_10703,N_6108,N_5019);
nor U10704 (N_10704,N_6516,N_5609);
and U10705 (N_10705,N_6102,N_6918);
nor U10706 (N_10706,N_7724,N_6633);
and U10707 (N_10707,N_4245,N_5101);
and U10708 (N_10708,N_5732,N_4590);
nor U10709 (N_10709,N_5633,N_5797);
nor U10710 (N_10710,N_7461,N_5010);
nand U10711 (N_10711,N_6761,N_5090);
and U10712 (N_10712,N_6423,N_4757);
or U10713 (N_10713,N_4993,N_4070);
nor U10714 (N_10714,N_7770,N_6291);
and U10715 (N_10715,N_4364,N_4097);
and U10716 (N_10716,N_5372,N_7998);
nand U10717 (N_10717,N_5076,N_6586);
and U10718 (N_10718,N_4978,N_7389);
and U10719 (N_10719,N_7257,N_4352);
or U10720 (N_10720,N_4259,N_6036);
or U10721 (N_10721,N_6128,N_5834);
and U10722 (N_10722,N_5457,N_4014);
nand U10723 (N_10723,N_6153,N_5396);
or U10724 (N_10724,N_4793,N_4890);
or U10725 (N_10725,N_4638,N_7711);
nand U10726 (N_10726,N_5994,N_5376);
and U10727 (N_10727,N_7203,N_7492);
or U10728 (N_10728,N_6993,N_5430);
nand U10729 (N_10729,N_6454,N_4778);
or U10730 (N_10730,N_7425,N_7137);
nor U10731 (N_10731,N_5276,N_6298);
and U10732 (N_10732,N_7648,N_7426);
and U10733 (N_10733,N_4153,N_4137);
nand U10734 (N_10734,N_5899,N_7102);
nand U10735 (N_10735,N_5361,N_5614);
or U10736 (N_10736,N_4195,N_7409);
and U10737 (N_10737,N_7487,N_6675);
or U10738 (N_10738,N_5009,N_4564);
and U10739 (N_10739,N_4409,N_6982);
nor U10740 (N_10740,N_7507,N_5596);
or U10741 (N_10741,N_7783,N_5022);
or U10742 (N_10742,N_5811,N_5485);
or U10743 (N_10743,N_7826,N_4985);
nor U10744 (N_10744,N_7734,N_6145);
and U10745 (N_10745,N_4235,N_6983);
nor U10746 (N_10746,N_4405,N_7298);
nor U10747 (N_10747,N_7854,N_6615);
or U10748 (N_10748,N_7625,N_7097);
and U10749 (N_10749,N_4193,N_7218);
nand U10750 (N_10750,N_5960,N_4845);
xor U10751 (N_10751,N_4962,N_4190);
or U10752 (N_10752,N_5957,N_6150);
nor U10753 (N_10753,N_6016,N_6449);
or U10754 (N_10754,N_5781,N_5254);
and U10755 (N_10755,N_5720,N_6346);
xnor U10756 (N_10756,N_5461,N_4618);
nand U10757 (N_10757,N_4405,N_6785);
or U10758 (N_10758,N_4286,N_5270);
and U10759 (N_10759,N_4427,N_7489);
and U10760 (N_10760,N_7836,N_6701);
nand U10761 (N_10761,N_5698,N_5169);
or U10762 (N_10762,N_4881,N_7699);
nor U10763 (N_10763,N_5469,N_7660);
or U10764 (N_10764,N_5006,N_6011);
nor U10765 (N_10765,N_7214,N_7639);
and U10766 (N_10766,N_7353,N_7260);
or U10767 (N_10767,N_4988,N_4698);
and U10768 (N_10768,N_6696,N_7015);
xor U10769 (N_10769,N_7281,N_5246);
xor U10770 (N_10770,N_4044,N_6386);
nand U10771 (N_10771,N_7128,N_7102);
nor U10772 (N_10772,N_5157,N_4654);
and U10773 (N_10773,N_5985,N_7963);
or U10774 (N_10774,N_6410,N_4984);
or U10775 (N_10775,N_4866,N_4868);
or U10776 (N_10776,N_6025,N_6624);
or U10777 (N_10777,N_5167,N_7910);
or U10778 (N_10778,N_7987,N_4884);
and U10779 (N_10779,N_7889,N_7678);
nand U10780 (N_10780,N_5508,N_4493);
nor U10781 (N_10781,N_7825,N_4549);
and U10782 (N_10782,N_4477,N_4888);
nand U10783 (N_10783,N_6483,N_6724);
or U10784 (N_10784,N_5512,N_6751);
nor U10785 (N_10785,N_4805,N_4992);
nand U10786 (N_10786,N_7231,N_7962);
nor U10787 (N_10787,N_5544,N_5890);
and U10788 (N_10788,N_5043,N_7133);
nand U10789 (N_10789,N_4370,N_7271);
nor U10790 (N_10790,N_6225,N_7384);
nand U10791 (N_10791,N_7882,N_4930);
or U10792 (N_10792,N_6036,N_5251);
and U10793 (N_10793,N_6018,N_7568);
and U10794 (N_10794,N_7741,N_5137);
or U10795 (N_10795,N_7609,N_5476);
or U10796 (N_10796,N_5638,N_5756);
or U10797 (N_10797,N_7324,N_5670);
nor U10798 (N_10798,N_6216,N_4667);
and U10799 (N_10799,N_6120,N_5145);
nor U10800 (N_10800,N_7475,N_4139);
or U10801 (N_10801,N_5306,N_5168);
and U10802 (N_10802,N_7740,N_5232);
nand U10803 (N_10803,N_6469,N_4728);
and U10804 (N_10804,N_5428,N_4012);
or U10805 (N_10805,N_5803,N_5850);
nand U10806 (N_10806,N_6559,N_5278);
nand U10807 (N_10807,N_4665,N_5800);
nand U10808 (N_10808,N_7680,N_5171);
nor U10809 (N_10809,N_7918,N_7339);
or U10810 (N_10810,N_7991,N_7719);
nor U10811 (N_10811,N_7489,N_5824);
and U10812 (N_10812,N_5521,N_6705);
nor U10813 (N_10813,N_5740,N_4223);
nor U10814 (N_10814,N_4853,N_5464);
nand U10815 (N_10815,N_5686,N_6692);
xor U10816 (N_10816,N_4859,N_7178);
nand U10817 (N_10817,N_4624,N_6101);
and U10818 (N_10818,N_4408,N_5983);
nand U10819 (N_10819,N_6492,N_5639);
or U10820 (N_10820,N_6422,N_5477);
nand U10821 (N_10821,N_7819,N_7705);
and U10822 (N_10822,N_6319,N_6570);
nand U10823 (N_10823,N_7169,N_7424);
and U10824 (N_10824,N_5957,N_4899);
or U10825 (N_10825,N_7364,N_5803);
nand U10826 (N_10826,N_7537,N_5277);
and U10827 (N_10827,N_5671,N_5623);
nor U10828 (N_10828,N_6807,N_5885);
nor U10829 (N_10829,N_6271,N_7642);
nand U10830 (N_10830,N_6724,N_6791);
or U10831 (N_10831,N_5772,N_7417);
nand U10832 (N_10832,N_4018,N_6442);
and U10833 (N_10833,N_7166,N_6129);
nor U10834 (N_10834,N_7886,N_5775);
and U10835 (N_10835,N_7877,N_6741);
and U10836 (N_10836,N_6905,N_7817);
nor U10837 (N_10837,N_4789,N_6681);
nor U10838 (N_10838,N_7754,N_4344);
nand U10839 (N_10839,N_7435,N_5197);
nand U10840 (N_10840,N_4818,N_6589);
or U10841 (N_10841,N_4719,N_5412);
and U10842 (N_10842,N_7249,N_5049);
or U10843 (N_10843,N_7198,N_7678);
or U10844 (N_10844,N_5818,N_5552);
or U10845 (N_10845,N_7294,N_4719);
nand U10846 (N_10846,N_4998,N_6220);
nor U10847 (N_10847,N_4613,N_4160);
nand U10848 (N_10848,N_5728,N_5045);
nor U10849 (N_10849,N_7933,N_5945);
nor U10850 (N_10850,N_5405,N_7356);
nor U10851 (N_10851,N_4758,N_4210);
nand U10852 (N_10852,N_4566,N_5024);
nor U10853 (N_10853,N_5671,N_4130);
and U10854 (N_10854,N_6258,N_7672);
and U10855 (N_10855,N_4210,N_6654);
or U10856 (N_10856,N_5054,N_4954);
nand U10857 (N_10857,N_6418,N_7917);
nand U10858 (N_10858,N_6254,N_6184);
or U10859 (N_10859,N_5931,N_6893);
nor U10860 (N_10860,N_6837,N_4671);
nor U10861 (N_10861,N_6490,N_7298);
or U10862 (N_10862,N_4528,N_7927);
nand U10863 (N_10863,N_6837,N_4889);
and U10864 (N_10864,N_7830,N_7684);
and U10865 (N_10865,N_4930,N_5847);
or U10866 (N_10866,N_4760,N_7379);
or U10867 (N_10867,N_6328,N_6152);
nand U10868 (N_10868,N_6354,N_5898);
or U10869 (N_10869,N_4948,N_5286);
nor U10870 (N_10870,N_6787,N_4276);
or U10871 (N_10871,N_4447,N_5436);
and U10872 (N_10872,N_6560,N_4502);
and U10873 (N_10873,N_7926,N_4750);
and U10874 (N_10874,N_4385,N_4176);
nand U10875 (N_10875,N_4246,N_5008);
nor U10876 (N_10876,N_4326,N_4957);
or U10877 (N_10877,N_5868,N_5161);
or U10878 (N_10878,N_4817,N_5917);
and U10879 (N_10879,N_5554,N_5991);
and U10880 (N_10880,N_4536,N_6085);
nor U10881 (N_10881,N_5271,N_7455);
nor U10882 (N_10882,N_4471,N_6654);
or U10883 (N_10883,N_5859,N_4111);
and U10884 (N_10884,N_5875,N_7319);
or U10885 (N_10885,N_4937,N_5401);
and U10886 (N_10886,N_7294,N_6121);
nor U10887 (N_10887,N_4559,N_4869);
or U10888 (N_10888,N_6890,N_4003);
nor U10889 (N_10889,N_6226,N_5080);
nand U10890 (N_10890,N_7950,N_7521);
nor U10891 (N_10891,N_7341,N_4825);
nor U10892 (N_10892,N_4176,N_6241);
and U10893 (N_10893,N_7115,N_7478);
nand U10894 (N_10894,N_4768,N_4661);
or U10895 (N_10895,N_5058,N_6496);
and U10896 (N_10896,N_4459,N_4109);
nor U10897 (N_10897,N_5772,N_7394);
or U10898 (N_10898,N_5363,N_5747);
nor U10899 (N_10899,N_5297,N_6723);
nor U10900 (N_10900,N_5167,N_7604);
or U10901 (N_10901,N_5087,N_5104);
nand U10902 (N_10902,N_7881,N_4708);
or U10903 (N_10903,N_7551,N_5984);
nor U10904 (N_10904,N_5207,N_5683);
and U10905 (N_10905,N_6240,N_4812);
or U10906 (N_10906,N_7983,N_4305);
nand U10907 (N_10907,N_7787,N_7943);
nor U10908 (N_10908,N_5139,N_4418);
or U10909 (N_10909,N_6934,N_7177);
nand U10910 (N_10910,N_7762,N_4623);
and U10911 (N_10911,N_6899,N_5899);
or U10912 (N_10912,N_7763,N_5253);
nor U10913 (N_10913,N_6577,N_7019);
or U10914 (N_10914,N_5052,N_7117);
nand U10915 (N_10915,N_5946,N_4361);
or U10916 (N_10916,N_5517,N_4051);
and U10917 (N_10917,N_6942,N_5108);
and U10918 (N_10918,N_7429,N_5169);
or U10919 (N_10919,N_5942,N_7253);
nand U10920 (N_10920,N_5651,N_5509);
or U10921 (N_10921,N_5996,N_7670);
or U10922 (N_10922,N_5891,N_7584);
and U10923 (N_10923,N_4070,N_6875);
and U10924 (N_10924,N_6999,N_7826);
and U10925 (N_10925,N_7306,N_7344);
nand U10926 (N_10926,N_6954,N_5869);
nand U10927 (N_10927,N_7758,N_4902);
nor U10928 (N_10928,N_4553,N_4158);
or U10929 (N_10929,N_4715,N_4634);
nand U10930 (N_10930,N_7015,N_6712);
and U10931 (N_10931,N_5579,N_6174);
nand U10932 (N_10932,N_7297,N_7693);
nand U10933 (N_10933,N_4700,N_7124);
or U10934 (N_10934,N_4709,N_6056);
and U10935 (N_10935,N_4334,N_4226);
and U10936 (N_10936,N_4238,N_5187);
nand U10937 (N_10937,N_5430,N_5103);
nand U10938 (N_10938,N_5850,N_5614);
nor U10939 (N_10939,N_6298,N_5272);
nor U10940 (N_10940,N_7986,N_4934);
nor U10941 (N_10941,N_5251,N_7760);
nand U10942 (N_10942,N_4920,N_7249);
and U10943 (N_10943,N_5837,N_4977);
nor U10944 (N_10944,N_5034,N_5378);
nor U10945 (N_10945,N_4731,N_4056);
nand U10946 (N_10946,N_4608,N_4677);
nor U10947 (N_10947,N_7642,N_7955);
or U10948 (N_10948,N_4817,N_6722);
nand U10949 (N_10949,N_7301,N_7676);
nor U10950 (N_10950,N_4924,N_6300);
and U10951 (N_10951,N_7056,N_5159);
and U10952 (N_10952,N_7117,N_6090);
nand U10953 (N_10953,N_4801,N_7086);
or U10954 (N_10954,N_4764,N_6250);
nand U10955 (N_10955,N_6187,N_7858);
and U10956 (N_10956,N_4292,N_4890);
nand U10957 (N_10957,N_6033,N_7006);
or U10958 (N_10958,N_5044,N_4348);
and U10959 (N_10959,N_4515,N_7801);
and U10960 (N_10960,N_5203,N_5581);
and U10961 (N_10961,N_5082,N_7988);
nand U10962 (N_10962,N_7977,N_5820);
nor U10963 (N_10963,N_5437,N_6420);
xnor U10964 (N_10964,N_6872,N_4841);
and U10965 (N_10965,N_6866,N_5592);
and U10966 (N_10966,N_7721,N_7449);
nor U10967 (N_10967,N_6452,N_5136);
or U10968 (N_10968,N_7844,N_4865);
or U10969 (N_10969,N_7780,N_7133);
nor U10970 (N_10970,N_6485,N_7200);
nor U10971 (N_10971,N_5742,N_5414);
nor U10972 (N_10972,N_6555,N_6671);
and U10973 (N_10973,N_6613,N_4066);
nand U10974 (N_10974,N_4559,N_6486);
nand U10975 (N_10975,N_7397,N_4250);
or U10976 (N_10976,N_7545,N_5546);
and U10977 (N_10977,N_4926,N_7641);
and U10978 (N_10978,N_5078,N_5985);
or U10979 (N_10979,N_5134,N_4988);
and U10980 (N_10980,N_5937,N_7168);
nand U10981 (N_10981,N_7602,N_6447);
xnor U10982 (N_10982,N_4363,N_5263);
nand U10983 (N_10983,N_6076,N_4459);
or U10984 (N_10984,N_5934,N_4501);
nand U10985 (N_10985,N_5023,N_5998);
or U10986 (N_10986,N_5034,N_4917);
or U10987 (N_10987,N_6622,N_7158);
nand U10988 (N_10988,N_5378,N_5558);
or U10989 (N_10989,N_5981,N_5407);
nor U10990 (N_10990,N_6288,N_6130);
nand U10991 (N_10991,N_5279,N_7004);
nand U10992 (N_10992,N_7973,N_5658);
and U10993 (N_10993,N_5729,N_7377);
nor U10994 (N_10994,N_6890,N_5528);
nand U10995 (N_10995,N_6036,N_6496);
nor U10996 (N_10996,N_5187,N_6640);
nor U10997 (N_10997,N_5373,N_5818);
nor U10998 (N_10998,N_6306,N_7619);
or U10999 (N_10999,N_6454,N_5956);
xor U11000 (N_11000,N_5624,N_7580);
and U11001 (N_11001,N_7180,N_5550);
or U11002 (N_11002,N_5321,N_4296);
or U11003 (N_11003,N_4650,N_5964);
or U11004 (N_11004,N_5206,N_4904);
and U11005 (N_11005,N_4016,N_7977);
or U11006 (N_11006,N_6416,N_5902);
or U11007 (N_11007,N_5446,N_6166);
and U11008 (N_11008,N_7130,N_5964);
nor U11009 (N_11009,N_4532,N_7120);
and U11010 (N_11010,N_6616,N_6264);
nor U11011 (N_11011,N_6119,N_5527);
or U11012 (N_11012,N_7612,N_6569);
nor U11013 (N_11013,N_6625,N_7690);
nand U11014 (N_11014,N_6159,N_4428);
nand U11015 (N_11015,N_4211,N_4947);
nand U11016 (N_11016,N_5169,N_6617);
nor U11017 (N_11017,N_6502,N_5592);
and U11018 (N_11018,N_6192,N_5509);
nor U11019 (N_11019,N_6736,N_6624);
nor U11020 (N_11020,N_5544,N_6634);
or U11021 (N_11021,N_5006,N_7182);
nand U11022 (N_11022,N_7825,N_7212);
or U11023 (N_11023,N_6326,N_6596);
and U11024 (N_11024,N_6195,N_7597);
nor U11025 (N_11025,N_5391,N_6917);
nor U11026 (N_11026,N_4305,N_7368);
or U11027 (N_11027,N_6547,N_5370);
nor U11028 (N_11028,N_7883,N_5510);
nor U11029 (N_11029,N_4937,N_7743);
nor U11030 (N_11030,N_7588,N_7558);
and U11031 (N_11031,N_6313,N_5253);
or U11032 (N_11032,N_5579,N_6962);
nor U11033 (N_11033,N_4727,N_6905);
or U11034 (N_11034,N_5769,N_4969);
nor U11035 (N_11035,N_4612,N_7129);
or U11036 (N_11036,N_4864,N_7935);
nor U11037 (N_11037,N_5235,N_5526);
or U11038 (N_11038,N_7293,N_7070);
or U11039 (N_11039,N_6606,N_7981);
nor U11040 (N_11040,N_5291,N_7524);
and U11041 (N_11041,N_6478,N_6297);
nor U11042 (N_11042,N_5837,N_4172);
nor U11043 (N_11043,N_5599,N_4070);
nand U11044 (N_11044,N_7299,N_6503);
nor U11045 (N_11045,N_7445,N_4963);
and U11046 (N_11046,N_7325,N_4421);
and U11047 (N_11047,N_4330,N_5591);
nor U11048 (N_11048,N_4705,N_7399);
or U11049 (N_11049,N_7398,N_4622);
nand U11050 (N_11050,N_4749,N_5282);
and U11051 (N_11051,N_7430,N_5754);
nand U11052 (N_11052,N_6369,N_6380);
nor U11053 (N_11053,N_6992,N_6479);
or U11054 (N_11054,N_6514,N_7466);
nor U11055 (N_11055,N_4491,N_6286);
and U11056 (N_11056,N_5181,N_5180);
and U11057 (N_11057,N_4127,N_4337);
nand U11058 (N_11058,N_6030,N_6050);
or U11059 (N_11059,N_6263,N_5214);
or U11060 (N_11060,N_5530,N_6112);
nand U11061 (N_11061,N_7998,N_5718);
and U11062 (N_11062,N_6010,N_7932);
and U11063 (N_11063,N_5063,N_7824);
nand U11064 (N_11064,N_4736,N_7870);
or U11065 (N_11065,N_5993,N_4058);
nand U11066 (N_11066,N_6083,N_5955);
nand U11067 (N_11067,N_4582,N_6578);
xnor U11068 (N_11068,N_4694,N_4712);
and U11069 (N_11069,N_5555,N_7922);
nand U11070 (N_11070,N_5475,N_7555);
nand U11071 (N_11071,N_7865,N_5857);
nor U11072 (N_11072,N_6649,N_6180);
nand U11073 (N_11073,N_4960,N_7367);
nor U11074 (N_11074,N_6638,N_6315);
or U11075 (N_11075,N_6899,N_5961);
nor U11076 (N_11076,N_7136,N_7892);
and U11077 (N_11077,N_5491,N_6188);
nor U11078 (N_11078,N_5872,N_7061);
or U11079 (N_11079,N_4664,N_4623);
or U11080 (N_11080,N_7658,N_7845);
nor U11081 (N_11081,N_7450,N_7799);
and U11082 (N_11082,N_7162,N_7824);
or U11083 (N_11083,N_5757,N_5639);
nor U11084 (N_11084,N_5861,N_4948);
or U11085 (N_11085,N_6517,N_5297);
nand U11086 (N_11086,N_7410,N_6918);
and U11087 (N_11087,N_5803,N_7132);
nand U11088 (N_11088,N_7200,N_7983);
nand U11089 (N_11089,N_6647,N_7992);
or U11090 (N_11090,N_5743,N_7030);
nand U11091 (N_11091,N_5351,N_6786);
or U11092 (N_11092,N_5267,N_6069);
nor U11093 (N_11093,N_4677,N_6920);
and U11094 (N_11094,N_4569,N_5629);
nor U11095 (N_11095,N_7974,N_4657);
nor U11096 (N_11096,N_7736,N_7572);
and U11097 (N_11097,N_5752,N_5220);
or U11098 (N_11098,N_7925,N_4482);
nand U11099 (N_11099,N_6051,N_6174);
and U11100 (N_11100,N_6805,N_7428);
nand U11101 (N_11101,N_6014,N_5252);
or U11102 (N_11102,N_4886,N_5970);
nand U11103 (N_11103,N_5832,N_5732);
and U11104 (N_11104,N_7840,N_6420);
xnor U11105 (N_11105,N_4511,N_7819);
nand U11106 (N_11106,N_4007,N_5419);
or U11107 (N_11107,N_6073,N_7818);
or U11108 (N_11108,N_4541,N_6189);
and U11109 (N_11109,N_6101,N_7259);
nand U11110 (N_11110,N_7522,N_4272);
nand U11111 (N_11111,N_6605,N_6324);
nor U11112 (N_11112,N_5859,N_6214);
nor U11113 (N_11113,N_5560,N_4188);
nand U11114 (N_11114,N_4214,N_7754);
nand U11115 (N_11115,N_6980,N_5067);
nor U11116 (N_11116,N_5552,N_5556);
or U11117 (N_11117,N_6228,N_6567);
and U11118 (N_11118,N_5512,N_7986);
nand U11119 (N_11119,N_4698,N_5981);
nand U11120 (N_11120,N_4793,N_5987);
and U11121 (N_11121,N_5637,N_4906);
nand U11122 (N_11122,N_7555,N_5098);
nand U11123 (N_11123,N_4094,N_5742);
nor U11124 (N_11124,N_5548,N_4756);
nor U11125 (N_11125,N_5817,N_6907);
and U11126 (N_11126,N_7905,N_5018);
and U11127 (N_11127,N_7634,N_5867);
and U11128 (N_11128,N_5651,N_6649);
xnor U11129 (N_11129,N_6880,N_6821);
nor U11130 (N_11130,N_5647,N_5047);
and U11131 (N_11131,N_5496,N_4788);
nand U11132 (N_11132,N_4320,N_6180);
or U11133 (N_11133,N_4750,N_5872);
nand U11134 (N_11134,N_6700,N_4369);
and U11135 (N_11135,N_7590,N_4307);
and U11136 (N_11136,N_7666,N_6466);
or U11137 (N_11137,N_5324,N_4533);
or U11138 (N_11138,N_6536,N_6210);
nand U11139 (N_11139,N_7321,N_5328);
or U11140 (N_11140,N_4813,N_4758);
or U11141 (N_11141,N_6948,N_6602);
nor U11142 (N_11142,N_6206,N_5380);
nand U11143 (N_11143,N_5840,N_7632);
nand U11144 (N_11144,N_6973,N_7259);
or U11145 (N_11145,N_7980,N_4978);
nand U11146 (N_11146,N_5589,N_7740);
nor U11147 (N_11147,N_7306,N_4756);
nand U11148 (N_11148,N_4559,N_4036);
or U11149 (N_11149,N_7394,N_4494);
or U11150 (N_11150,N_6541,N_4752);
and U11151 (N_11151,N_5983,N_5024);
nand U11152 (N_11152,N_6409,N_5896);
or U11153 (N_11153,N_7682,N_4948);
and U11154 (N_11154,N_7490,N_7807);
nand U11155 (N_11155,N_5251,N_4927);
nand U11156 (N_11156,N_6538,N_4754);
and U11157 (N_11157,N_7373,N_5690);
or U11158 (N_11158,N_5540,N_7235);
nand U11159 (N_11159,N_7028,N_4641);
and U11160 (N_11160,N_5814,N_4860);
and U11161 (N_11161,N_6407,N_4288);
and U11162 (N_11162,N_5919,N_6018);
or U11163 (N_11163,N_6437,N_4016);
or U11164 (N_11164,N_5872,N_7696);
and U11165 (N_11165,N_6988,N_4212);
and U11166 (N_11166,N_4186,N_7662);
or U11167 (N_11167,N_4100,N_5861);
nor U11168 (N_11168,N_7601,N_7791);
nand U11169 (N_11169,N_6091,N_4834);
nand U11170 (N_11170,N_4168,N_7047);
or U11171 (N_11171,N_4155,N_4761);
nand U11172 (N_11172,N_4610,N_4659);
or U11173 (N_11173,N_4129,N_4560);
and U11174 (N_11174,N_7381,N_6018);
nor U11175 (N_11175,N_7602,N_7212);
or U11176 (N_11176,N_5903,N_6212);
nor U11177 (N_11177,N_5264,N_6069);
or U11178 (N_11178,N_7746,N_6156);
xor U11179 (N_11179,N_6321,N_6381);
nand U11180 (N_11180,N_5285,N_4855);
nor U11181 (N_11181,N_7919,N_5319);
nor U11182 (N_11182,N_7477,N_4167);
or U11183 (N_11183,N_6924,N_4025);
nor U11184 (N_11184,N_6978,N_6912);
nand U11185 (N_11185,N_5449,N_5957);
and U11186 (N_11186,N_6774,N_4966);
nor U11187 (N_11187,N_7762,N_7277);
or U11188 (N_11188,N_5197,N_5162);
or U11189 (N_11189,N_6455,N_6125);
or U11190 (N_11190,N_7965,N_4692);
nor U11191 (N_11191,N_7867,N_4913);
and U11192 (N_11192,N_4205,N_5670);
or U11193 (N_11193,N_6430,N_6892);
and U11194 (N_11194,N_5400,N_5397);
nand U11195 (N_11195,N_7735,N_5300);
or U11196 (N_11196,N_6058,N_7055);
and U11197 (N_11197,N_4790,N_4455);
and U11198 (N_11198,N_4533,N_4207);
nor U11199 (N_11199,N_7056,N_6425);
nor U11200 (N_11200,N_6924,N_7778);
or U11201 (N_11201,N_5993,N_4771);
and U11202 (N_11202,N_6762,N_7796);
or U11203 (N_11203,N_7626,N_7982);
nor U11204 (N_11204,N_4715,N_6203);
nor U11205 (N_11205,N_5881,N_7534);
or U11206 (N_11206,N_4318,N_7460);
nand U11207 (N_11207,N_4983,N_7277);
nor U11208 (N_11208,N_6457,N_6801);
and U11209 (N_11209,N_5027,N_7912);
and U11210 (N_11210,N_4127,N_7753);
nand U11211 (N_11211,N_7706,N_5698);
nor U11212 (N_11212,N_7826,N_6632);
nor U11213 (N_11213,N_5892,N_4551);
nor U11214 (N_11214,N_4506,N_6456);
nor U11215 (N_11215,N_4547,N_4724);
nand U11216 (N_11216,N_5787,N_6602);
nand U11217 (N_11217,N_7018,N_7651);
nand U11218 (N_11218,N_6777,N_6369);
nand U11219 (N_11219,N_5355,N_5079);
nand U11220 (N_11220,N_4019,N_4841);
nor U11221 (N_11221,N_6704,N_5715);
nor U11222 (N_11222,N_5303,N_4729);
nor U11223 (N_11223,N_4282,N_4749);
nand U11224 (N_11224,N_7277,N_7211);
or U11225 (N_11225,N_6158,N_4516);
or U11226 (N_11226,N_4643,N_4100);
or U11227 (N_11227,N_7566,N_6097);
nor U11228 (N_11228,N_4392,N_6831);
and U11229 (N_11229,N_4677,N_7350);
nor U11230 (N_11230,N_4533,N_4741);
and U11231 (N_11231,N_5437,N_5562);
or U11232 (N_11232,N_4297,N_6876);
or U11233 (N_11233,N_7689,N_7894);
nand U11234 (N_11234,N_4351,N_7349);
or U11235 (N_11235,N_4115,N_6832);
nor U11236 (N_11236,N_4800,N_6851);
nor U11237 (N_11237,N_7315,N_7809);
nor U11238 (N_11238,N_5419,N_5862);
nand U11239 (N_11239,N_5953,N_5126);
and U11240 (N_11240,N_5669,N_5007);
and U11241 (N_11241,N_7931,N_7776);
nand U11242 (N_11242,N_6426,N_7924);
nor U11243 (N_11243,N_5138,N_6790);
nor U11244 (N_11244,N_4120,N_4966);
nand U11245 (N_11245,N_5077,N_6137);
nand U11246 (N_11246,N_7099,N_5929);
and U11247 (N_11247,N_4988,N_6731);
or U11248 (N_11248,N_7477,N_7160);
nand U11249 (N_11249,N_6063,N_6159);
nor U11250 (N_11250,N_6069,N_6599);
and U11251 (N_11251,N_5824,N_4353);
nor U11252 (N_11252,N_5488,N_6087);
nand U11253 (N_11253,N_5659,N_7915);
nand U11254 (N_11254,N_4047,N_7051);
nand U11255 (N_11255,N_4963,N_5338);
nor U11256 (N_11256,N_6968,N_6812);
and U11257 (N_11257,N_6466,N_4184);
and U11258 (N_11258,N_4752,N_6123);
nand U11259 (N_11259,N_6783,N_5911);
nor U11260 (N_11260,N_7298,N_4299);
and U11261 (N_11261,N_6715,N_4469);
nor U11262 (N_11262,N_4014,N_7768);
nor U11263 (N_11263,N_4905,N_7923);
or U11264 (N_11264,N_5850,N_6194);
or U11265 (N_11265,N_4120,N_4282);
nand U11266 (N_11266,N_4614,N_7016);
nor U11267 (N_11267,N_5554,N_7224);
nor U11268 (N_11268,N_7150,N_7203);
or U11269 (N_11269,N_4262,N_5123);
nor U11270 (N_11270,N_5055,N_5735);
or U11271 (N_11271,N_5470,N_6658);
nand U11272 (N_11272,N_6394,N_5255);
nand U11273 (N_11273,N_5497,N_5701);
or U11274 (N_11274,N_6000,N_4340);
or U11275 (N_11275,N_7356,N_6884);
and U11276 (N_11276,N_7804,N_4233);
and U11277 (N_11277,N_4029,N_4993);
or U11278 (N_11278,N_4322,N_4077);
nor U11279 (N_11279,N_7161,N_4609);
or U11280 (N_11280,N_6460,N_5664);
nor U11281 (N_11281,N_6128,N_7525);
nor U11282 (N_11282,N_7258,N_6681);
and U11283 (N_11283,N_4442,N_6558);
or U11284 (N_11284,N_6776,N_5902);
and U11285 (N_11285,N_6864,N_6001);
nor U11286 (N_11286,N_5390,N_4161);
and U11287 (N_11287,N_7413,N_7124);
and U11288 (N_11288,N_6282,N_6255);
or U11289 (N_11289,N_4110,N_6584);
nand U11290 (N_11290,N_4935,N_6774);
and U11291 (N_11291,N_7839,N_4159);
nor U11292 (N_11292,N_5849,N_7204);
nand U11293 (N_11293,N_5989,N_6785);
nand U11294 (N_11294,N_6825,N_4438);
or U11295 (N_11295,N_7789,N_6371);
nor U11296 (N_11296,N_6521,N_6102);
nor U11297 (N_11297,N_4936,N_4199);
nand U11298 (N_11298,N_4645,N_6005);
nor U11299 (N_11299,N_5159,N_6523);
nor U11300 (N_11300,N_5471,N_4304);
and U11301 (N_11301,N_6421,N_4916);
or U11302 (N_11302,N_7711,N_7866);
nand U11303 (N_11303,N_4893,N_6472);
nand U11304 (N_11304,N_5626,N_6095);
nand U11305 (N_11305,N_4512,N_5016);
or U11306 (N_11306,N_4894,N_7588);
nand U11307 (N_11307,N_5272,N_4854);
nor U11308 (N_11308,N_4365,N_4639);
and U11309 (N_11309,N_5319,N_7895);
nor U11310 (N_11310,N_5294,N_7916);
and U11311 (N_11311,N_7762,N_6383);
nor U11312 (N_11312,N_4617,N_5736);
or U11313 (N_11313,N_7217,N_4233);
and U11314 (N_11314,N_7720,N_7180);
nand U11315 (N_11315,N_7485,N_5889);
or U11316 (N_11316,N_4667,N_7019);
nor U11317 (N_11317,N_4899,N_5670);
nor U11318 (N_11318,N_4931,N_5890);
nand U11319 (N_11319,N_5136,N_5097);
and U11320 (N_11320,N_7286,N_6153);
or U11321 (N_11321,N_7646,N_4606);
or U11322 (N_11322,N_6982,N_6295);
and U11323 (N_11323,N_7675,N_7587);
nand U11324 (N_11324,N_4389,N_6093);
nor U11325 (N_11325,N_6143,N_7873);
xnor U11326 (N_11326,N_5435,N_4746);
nor U11327 (N_11327,N_6160,N_7502);
nand U11328 (N_11328,N_4911,N_4030);
and U11329 (N_11329,N_6625,N_5295);
nand U11330 (N_11330,N_5067,N_7148);
or U11331 (N_11331,N_7946,N_4933);
nand U11332 (N_11332,N_6028,N_5694);
nor U11333 (N_11333,N_5524,N_6150);
or U11334 (N_11334,N_7871,N_4028);
or U11335 (N_11335,N_5258,N_4086);
and U11336 (N_11336,N_7895,N_5450);
nor U11337 (N_11337,N_4523,N_6043);
and U11338 (N_11338,N_5776,N_4011);
nor U11339 (N_11339,N_6612,N_6316);
nand U11340 (N_11340,N_5283,N_6330);
nor U11341 (N_11341,N_6354,N_4798);
nand U11342 (N_11342,N_5958,N_5179);
nor U11343 (N_11343,N_7156,N_7154);
and U11344 (N_11344,N_6538,N_5260);
and U11345 (N_11345,N_6311,N_5370);
or U11346 (N_11346,N_4803,N_5210);
nand U11347 (N_11347,N_6601,N_4416);
nand U11348 (N_11348,N_4180,N_6737);
and U11349 (N_11349,N_6932,N_4380);
nor U11350 (N_11350,N_7506,N_4748);
or U11351 (N_11351,N_5432,N_5836);
nand U11352 (N_11352,N_7551,N_7094);
nand U11353 (N_11353,N_6760,N_4457);
and U11354 (N_11354,N_4152,N_6796);
and U11355 (N_11355,N_6385,N_5542);
or U11356 (N_11356,N_7704,N_6316);
nor U11357 (N_11357,N_6745,N_7451);
nand U11358 (N_11358,N_5483,N_4037);
nand U11359 (N_11359,N_4726,N_7908);
and U11360 (N_11360,N_7893,N_5753);
and U11361 (N_11361,N_4471,N_7345);
nor U11362 (N_11362,N_6928,N_6458);
nor U11363 (N_11363,N_7075,N_5757);
nor U11364 (N_11364,N_7359,N_6498);
xor U11365 (N_11365,N_5601,N_5464);
nand U11366 (N_11366,N_6445,N_6073);
and U11367 (N_11367,N_4564,N_4588);
or U11368 (N_11368,N_6056,N_7924);
and U11369 (N_11369,N_7026,N_6328);
or U11370 (N_11370,N_4738,N_6637);
or U11371 (N_11371,N_6265,N_6926);
or U11372 (N_11372,N_7571,N_5971);
nand U11373 (N_11373,N_5176,N_5103);
and U11374 (N_11374,N_5426,N_6431);
nand U11375 (N_11375,N_4352,N_4071);
nor U11376 (N_11376,N_5685,N_4847);
or U11377 (N_11377,N_7315,N_6230);
nor U11378 (N_11378,N_4251,N_7619);
and U11379 (N_11379,N_7805,N_7105);
and U11380 (N_11380,N_4659,N_5722);
nand U11381 (N_11381,N_6053,N_5550);
nor U11382 (N_11382,N_5700,N_7383);
or U11383 (N_11383,N_7742,N_5914);
or U11384 (N_11384,N_6495,N_5283);
nor U11385 (N_11385,N_5906,N_6749);
nor U11386 (N_11386,N_6910,N_6691);
or U11387 (N_11387,N_5159,N_6118);
nor U11388 (N_11388,N_4737,N_6824);
and U11389 (N_11389,N_5145,N_7365);
or U11390 (N_11390,N_7196,N_7227);
and U11391 (N_11391,N_5441,N_7391);
nor U11392 (N_11392,N_6453,N_7008);
and U11393 (N_11393,N_6804,N_7086);
nand U11394 (N_11394,N_7436,N_6372);
and U11395 (N_11395,N_5632,N_7483);
nand U11396 (N_11396,N_6873,N_5877);
nand U11397 (N_11397,N_7012,N_4523);
nor U11398 (N_11398,N_6533,N_6682);
nand U11399 (N_11399,N_6093,N_6510);
nor U11400 (N_11400,N_4016,N_7385);
and U11401 (N_11401,N_7336,N_5379);
or U11402 (N_11402,N_6550,N_4347);
nor U11403 (N_11403,N_7492,N_7443);
nor U11404 (N_11404,N_6124,N_5287);
nor U11405 (N_11405,N_4612,N_5928);
or U11406 (N_11406,N_4320,N_5409);
or U11407 (N_11407,N_6519,N_4826);
or U11408 (N_11408,N_5273,N_5061);
or U11409 (N_11409,N_4482,N_6118);
or U11410 (N_11410,N_5583,N_7569);
or U11411 (N_11411,N_6296,N_7810);
nand U11412 (N_11412,N_7930,N_4089);
nor U11413 (N_11413,N_7612,N_4765);
nor U11414 (N_11414,N_5962,N_5309);
and U11415 (N_11415,N_4283,N_7178);
nor U11416 (N_11416,N_4080,N_5658);
nand U11417 (N_11417,N_6455,N_4299);
or U11418 (N_11418,N_7585,N_7845);
or U11419 (N_11419,N_6709,N_6906);
or U11420 (N_11420,N_7811,N_6508);
nand U11421 (N_11421,N_5949,N_6067);
nand U11422 (N_11422,N_7483,N_6495);
nand U11423 (N_11423,N_7869,N_5280);
nand U11424 (N_11424,N_4796,N_7994);
and U11425 (N_11425,N_7758,N_5181);
and U11426 (N_11426,N_5572,N_7931);
nor U11427 (N_11427,N_6782,N_4334);
nand U11428 (N_11428,N_5522,N_5427);
or U11429 (N_11429,N_7660,N_7850);
nor U11430 (N_11430,N_7296,N_4448);
or U11431 (N_11431,N_4525,N_5786);
nor U11432 (N_11432,N_6506,N_4915);
and U11433 (N_11433,N_4153,N_6004);
and U11434 (N_11434,N_5115,N_5082);
or U11435 (N_11435,N_5979,N_7295);
or U11436 (N_11436,N_4940,N_6351);
xnor U11437 (N_11437,N_6396,N_4345);
nand U11438 (N_11438,N_4087,N_6698);
nor U11439 (N_11439,N_4855,N_4174);
nand U11440 (N_11440,N_6664,N_7132);
or U11441 (N_11441,N_4266,N_7766);
nand U11442 (N_11442,N_4102,N_6534);
and U11443 (N_11443,N_5463,N_6830);
nor U11444 (N_11444,N_7968,N_4822);
nand U11445 (N_11445,N_5768,N_4471);
nor U11446 (N_11446,N_6412,N_4108);
or U11447 (N_11447,N_6002,N_6632);
and U11448 (N_11448,N_6093,N_6943);
nor U11449 (N_11449,N_4767,N_5461);
and U11450 (N_11450,N_4929,N_6862);
nand U11451 (N_11451,N_5576,N_6146);
nor U11452 (N_11452,N_5478,N_5594);
or U11453 (N_11453,N_5199,N_7093);
or U11454 (N_11454,N_6386,N_6625);
or U11455 (N_11455,N_4923,N_6731);
nand U11456 (N_11456,N_6661,N_4139);
nor U11457 (N_11457,N_6473,N_5014);
nor U11458 (N_11458,N_6960,N_4694);
nand U11459 (N_11459,N_6264,N_5979);
nand U11460 (N_11460,N_5926,N_5073);
and U11461 (N_11461,N_5635,N_4913);
nand U11462 (N_11462,N_5130,N_7769);
nor U11463 (N_11463,N_4268,N_7551);
or U11464 (N_11464,N_4414,N_4783);
and U11465 (N_11465,N_4661,N_7121);
nand U11466 (N_11466,N_5344,N_5499);
xnor U11467 (N_11467,N_5439,N_6017);
or U11468 (N_11468,N_5807,N_4924);
or U11469 (N_11469,N_6075,N_7649);
xnor U11470 (N_11470,N_4694,N_6583);
or U11471 (N_11471,N_6933,N_5913);
nand U11472 (N_11472,N_6742,N_5424);
nand U11473 (N_11473,N_4589,N_6800);
nor U11474 (N_11474,N_6732,N_7789);
nor U11475 (N_11475,N_5257,N_7819);
or U11476 (N_11476,N_7690,N_7444);
or U11477 (N_11477,N_5803,N_6890);
and U11478 (N_11478,N_5368,N_5502);
nor U11479 (N_11479,N_5838,N_6167);
nor U11480 (N_11480,N_6761,N_7854);
nor U11481 (N_11481,N_7800,N_6094);
or U11482 (N_11482,N_4794,N_4467);
and U11483 (N_11483,N_5173,N_5849);
and U11484 (N_11484,N_4628,N_6444);
nor U11485 (N_11485,N_4888,N_6461);
nor U11486 (N_11486,N_6788,N_7368);
or U11487 (N_11487,N_6292,N_7345);
and U11488 (N_11488,N_5135,N_7756);
or U11489 (N_11489,N_5633,N_6202);
and U11490 (N_11490,N_7454,N_7772);
nor U11491 (N_11491,N_6696,N_5509);
and U11492 (N_11492,N_5193,N_6779);
nor U11493 (N_11493,N_4909,N_5173);
or U11494 (N_11494,N_6711,N_7575);
and U11495 (N_11495,N_4285,N_4942);
and U11496 (N_11496,N_6319,N_4178);
and U11497 (N_11497,N_6491,N_7379);
nor U11498 (N_11498,N_6282,N_4998);
or U11499 (N_11499,N_6603,N_6126);
nand U11500 (N_11500,N_4004,N_5179);
and U11501 (N_11501,N_7667,N_7061);
or U11502 (N_11502,N_7491,N_4472);
and U11503 (N_11503,N_5960,N_7309);
nor U11504 (N_11504,N_6826,N_4258);
nor U11505 (N_11505,N_6212,N_4731);
nand U11506 (N_11506,N_4857,N_6087);
nor U11507 (N_11507,N_6521,N_4536);
or U11508 (N_11508,N_6025,N_6994);
and U11509 (N_11509,N_6813,N_6624);
nand U11510 (N_11510,N_7701,N_4786);
or U11511 (N_11511,N_5304,N_6220);
nor U11512 (N_11512,N_6852,N_4374);
nand U11513 (N_11513,N_7016,N_7098);
or U11514 (N_11514,N_5983,N_7028);
nand U11515 (N_11515,N_6934,N_6773);
or U11516 (N_11516,N_6785,N_4211);
or U11517 (N_11517,N_7557,N_7491);
nand U11518 (N_11518,N_6887,N_7620);
and U11519 (N_11519,N_4865,N_6097);
nand U11520 (N_11520,N_5609,N_7110);
or U11521 (N_11521,N_7750,N_7038);
nor U11522 (N_11522,N_5719,N_6757);
or U11523 (N_11523,N_6714,N_7438);
nor U11524 (N_11524,N_6196,N_7416);
nand U11525 (N_11525,N_4943,N_5040);
or U11526 (N_11526,N_4977,N_7201);
nor U11527 (N_11527,N_6991,N_6128);
nand U11528 (N_11528,N_7428,N_7999);
nand U11529 (N_11529,N_5790,N_4690);
nor U11530 (N_11530,N_7535,N_7839);
nor U11531 (N_11531,N_7644,N_7268);
or U11532 (N_11532,N_6610,N_5773);
or U11533 (N_11533,N_6508,N_7001);
or U11534 (N_11534,N_6051,N_7706);
nor U11535 (N_11535,N_5702,N_5217);
nor U11536 (N_11536,N_4366,N_5065);
or U11537 (N_11537,N_4979,N_6571);
and U11538 (N_11538,N_5337,N_6995);
and U11539 (N_11539,N_7782,N_6752);
nor U11540 (N_11540,N_5449,N_4669);
nor U11541 (N_11541,N_7885,N_7965);
and U11542 (N_11542,N_7929,N_5416);
or U11543 (N_11543,N_5223,N_4385);
nor U11544 (N_11544,N_5726,N_6393);
or U11545 (N_11545,N_7667,N_6091);
nor U11546 (N_11546,N_6491,N_5158);
and U11547 (N_11547,N_4022,N_7733);
and U11548 (N_11548,N_5100,N_4804);
xnor U11549 (N_11549,N_4739,N_6045);
nand U11550 (N_11550,N_7789,N_7467);
and U11551 (N_11551,N_4304,N_4002);
and U11552 (N_11552,N_4454,N_6293);
nand U11553 (N_11553,N_5006,N_7007);
nor U11554 (N_11554,N_4590,N_4429);
or U11555 (N_11555,N_6525,N_5008);
or U11556 (N_11556,N_6075,N_6354);
nor U11557 (N_11557,N_4843,N_6257);
nand U11558 (N_11558,N_6328,N_7142);
and U11559 (N_11559,N_7576,N_6656);
nand U11560 (N_11560,N_4693,N_6942);
and U11561 (N_11561,N_4443,N_5905);
nor U11562 (N_11562,N_5851,N_5792);
nand U11563 (N_11563,N_5197,N_4881);
and U11564 (N_11564,N_7732,N_7465);
or U11565 (N_11565,N_7384,N_4097);
or U11566 (N_11566,N_7266,N_4741);
nor U11567 (N_11567,N_5220,N_4677);
nor U11568 (N_11568,N_5642,N_5101);
or U11569 (N_11569,N_4859,N_4390);
nor U11570 (N_11570,N_7469,N_6370);
or U11571 (N_11571,N_5082,N_6959);
nor U11572 (N_11572,N_4137,N_7945);
nand U11573 (N_11573,N_7824,N_4444);
or U11574 (N_11574,N_5204,N_5386);
nor U11575 (N_11575,N_6233,N_6878);
or U11576 (N_11576,N_4826,N_7713);
and U11577 (N_11577,N_4458,N_7871);
or U11578 (N_11578,N_6237,N_6655);
and U11579 (N_11579,N_7597,N_7161);
or U11580 (N_11580,N_5198,N_6223);
and U11581 (N_11581,N_7299,N_7497);
nand U11582 (N_11582,N_6867,N_4666);
and U11583 (N_11583,N_5295,N_6262);
nand U11584 (N_11584,N_6104,N_4159);
and U11585 (N_11585,N_5495,N_7722);
nand U11586 (N_11586,N_5537,N_7840);
and U11587 (N_11587,N_5719,N_6150);
nor U11588 (N_11588,N_6333,N_4099);
nor U11589 (N_11589,N_4559,N_6561);
or U11590 (N_11590,N_6874,N_6822);
and U11591 (N_11591,N_4660,N_7519);
or U11592 (N_11592,N_4448,N_6683);
nor U11593 (N_11593,N_6910,N_7485);
or U11594 (N_11594,N_6700,N_7619);
and U11595 (N_11595,N_6106,N_4448);
nor U11596 (N_11596,N_7169,N_6904);
nor U11597 (N_11597,N_5920,N_5805);
or U11598 (N_11598,N_6282,N_4949);
nor U11599 (N_11599,N_4753,N_6153);
nor U11600 (N_11600,N_5829,N_6861);
nor U11601 (N_11601,N_4947,N_7421);
nand U11602 (N_11602,N_4239,N_7824);
nand U11603 (N_11603,N_6493,N_6905);
nor U11604 (N_11604,N_5911,N_5192);
nand U11605 (N_11605,N_4137,N_7510);
and U11606 (N_11606,N_4378,N_6771);
or U11607 (N_11607,N_6690,N_6812);
and U11608 (N_11608,N_5221,N_5850);
nand U11609 (N_11609,N_6436,N_6991);
and U11610 (N_11610,N_5865,N_4817);
nor U11611 (N_11611,N_5057,N_4345);
or U11612 (N_11612,N_4216,N_6981);
and U11613 (N_11613,N_4565,N_6313);
nor U11614 (N_11614,N_5080,N_6521);
and U11615 (N_11615,N_4513,N_6560);
or U11616 (N_11616,N_5230,N_4118);
nor U11617 (N_11617,N_6136,N_5088);
or U11618 (N_11618,N_6199,N_5206);
or U11619 (N_11619,N_7195,N_4646);
and U11620 (N_11620,N_5011,N_5691);
nor U11621 (N_11621,N_6606,N_7378);
nand U11622 (N_11622,N_7004,N_7698);
nor U11623 (N_11623,N_7762,N_5189);
nor U11624 (N_11624,N_7851,N_5360);
and U11625 (N_11625,N_6218,N_7906);
nand U11626 (N_11626,N_6970,N_6735);
nand U11627 (N_11627,N_7957,N_6826);
or U11628 (N_11628,N_5563,N_7997);
or U11629 (N_11629,N_5726,N_6096);
and U11630 (N_11630,N_5209,N_7571);
xor U11631 (N_11631,N_4179,N_5121);
and U11632 (N_11632,N_7813,N_4729);
and U11633 (N_11633,N_6688,N_4757);
or U11634 (N_11634,N_5946,N_5486);
and U11635 (N_11635,N_5864,N_7575);
nor U11636 (N_11636,N_6079,N_4621);
or U11637 (N_11637,N_6614,N_7349);
nor U11638 (N_11638,N_5224,N_7714);
nand U11639 (N_11639,N_7664,N_7409);
nand U11640 (N_11640,N_4618,N_4725);
or U11641 (N_11641,N_4301,N_5145);
nor U11642 (N_11642,N_6133,N_7936);
nand U11643 (N_11643,N_4470,N_7770);
and U11644 (N_11644,N_7465,N_4431);
nand U11645 (N_11645,N_7712,N_7781);
nor U11646 (N_11646,N_5909,N_5013);
and U11647 (N_11647,N_7938,N_7057);
nor U11648 (N_11648,N_6926,N_7329);
or U11649 (N_11649,N_4373,N_4258);
nand U11650 (N_11650,N_6814,N_6288);
or U11651 (N_11651,N_4172,N_6943);
and U11652 (N_11652,N_7368,N_6559);
and U11653 (N_11653,N_4107,N_5222);
nand U11654 (N_11654,N_5813,N_5082);
and U11655 (N_11655,N_6253,N_5130);
and U11656 (N_11656,N_6898,N_4592);
nor U11657 (N_11657,N_5698,N_7223);
nor U11658 (N_11658,N_7663,N_4905);
or U11659 (N_11659,N_6820,N_5208);
and U11660 (N_11660,N_7351,N_4891);
nor U11661 (N_11661,N_6031,N_4084);
and U11662 (N_11662,N_5047,N_4910);
and U11663 (N_11663,N_6632,N_4659);
or U11664 (N_11664,N_4594,N_4850);
and U11665 (N_11665,N_7986,N_6641);
nor U11666 (N_11666,N_5784,N_5193);
nand U11667 (N_11667,N_6511,N_7289);
or U11668 (N_11668,N_7419,N_4531);
and U11669 (N_11669,N_6573,N_5491);
nand U11670 (N_11670,N_7917,N_7648);
or U11671 (N_11671,N_5297,N_6672);
nor U11672 (N_11672,N_5115,N_5210);
or U11673 (N_11673,N_4459,N_7550);
nand U11674 (N_11674,N_5848,N_5050);
and U11675 (N_11675,N_6645,N_5206);
or U11676 (N_11676,N_4063,N_6385);
or U11677 (N_11677,N_7930,N_7722);
nor U11678 (N_11678,N_7156,N_6832);
or U11679 (N_11679,N_5169,N_4283);
nand U11680 (N_11680,N_5103,N_6516);
nor U11681 (N_11681,N_7011,N_5955);
and U11682 (N_11682,N_4200,N_5912);
nor U11683 (N_11683,N_6223,N_4652);
and U11684 (N_11684,N_7095,N_6483);
or U11685 (N_11685,N_5825,N_7802);
nand U11686 (N_11686,N_6284,N_7786);
nor U11687 (N_11687,N_5038,N_7518);
or U11688 (N_11688,N_4945,N_5332);
or U11689 (N_11689,N_4554,N_6806);
or U11690 (N_11690,N_5217,N_6719);
and U11691 (N_11691,N_5197,N_5334);
and U11692 (N_11692,N_7269,N_7668);
and U11693 (N_11693,N_5371,N_7703);
and U11694 (N_11694,N_5623,N_4586);
or U11695 (N_11695,N_5774,N_4201);
nand U11696 (N_11696,N_5626,N_7240);
nor U11697 (N_11697,N_5020,N_4082);
and U11698 (N_11698,N_4352,N_5268);
nand U11699 (N_11699,N_6502,N_5020);
or U11700 (N_11700,N_5759,N_4133);
nor U11701 (N_11701,N_6203,N_5300);
and U11702 (N_11702,N_4471,N_5313);
nor U11703 (N_11703,N_6203,N_5951);
nand U11704 (N_11704,N_4647,N_5762);
nand U11705 (N_11705,N_6414,N_7323);
and U11706 (N_11706,N_6530,N_4382);
or U11707 (N_11707,N_4369,N_7249);
and U11708 (N_11708,N_4681,N_7515);
xnor U11709 (N_11709,N_4965,N_5537);
and U11710 (N_11710,N_7900,N_7620);
or U11711 (N_11711,N_4659,N_5985);
nand U11712 (N_11712,N_6884,N_5725);
or U11713 (N_11713,N_5148,N_7444);
or U11714 (N_11714,N_7115,N_4691);
or U11715 (N_11715,N_4307,N_6459);
nand U11716 (N_11716,N_5775,N_7358);
nor U11717 (N_11717,N_5575,N_5715);
nor U11718 (N_11718,N_6410,N_7755);
xnor U11719 (N_11719,N_5304,N_7027);
and U11720 (N_11720,N_5088,N_6229);
nor U11721 (N_11721,N_7505,N_4233);
nor U11722 (N_11722,N_4336,N_4082);
and U11723 (N_11723,N_4070,N_4307);
and U11724 (N_11724,N_6784,N_7290);
and U11725 (N_11725,N_4464,N_6498);
nand U11726 (N_11726,N_5780,N_5251);
nor U11727 (N_11727,N_7415,N_5208);
and U11728 (N_11728,N_4323,N_5936);
or U11729 (N_11729,N_4511,N_7333);
nor U11730 (N_11730,N_5400,N_7201);
and U11731 (N_11731,N_6401,N_6658);
or U11732 (N_11732,N_5336,N_6792);
nor U11733 (N_11733,N_5826,N_5875);
or U11734 (N_11734,N_6406,N_5773);
nor U11735 (N_11735,N_6611,N_4901);
nor U11736 (N_11736,N_7623,N_6972);
and U11737 (N_11737,N_5392,N_5028);
nand U11738 (N_11738,N_5126,N_6457);
nand U11739 (N_11739,N_4104,N_7246);
or U11740 (N_11740,N_7815,N_6364);
or U11741 (N_11741,N_4642,N_5460);
and U11742 (N_11742,N_4102,N_6199);
or U11743 (N_11743,N_5507,N_7713);
nand U11744 (N_11744,N_5841,N_7045);
or U11745 (N_11745,N_6735,N_7302);
nand U11746 (N_11746,N_6921,N_4326);
nand U11747 (N_11747,N_4175,N_5456);
and U11748 (N_11748,N_6123,N_6757);
nor U11749 (N_11749,N_7745,N_7493);
nor U11750 (N_11750,N_7851,N_7918);
and U11751 (N_11751,N_6273,N_5868);
nand U11752 (N_11752,N_7023,N_4820);
or U11753 (N_11753,N_7573,N_5294);
or U11754 (N_11754,N_6302,N_5150);
nand U11755 (N_11755,N_4771,N_7018);
nand U11756 (N_11756,N_6376,N_4930);
nand U11757 (N_11757,N_7412,N_7215);
or U11758 (N_11758,N_4395,N_7185);
or U11759 (N_11759,N_4644,N_7821);
nor U11760 (N_11760,N_5419,N_5187);
or U11761 (N_11761,N_7408,N_5847);
and U11762 (N_11762,N_6399,N_7350);
nand U11763 (N_11763,N_7824,N_6448);
or U11764 (N_11764,N_7398,N_6904);
xor U11765 (N_11765,N_7684,N_7881);
and U11766 (N_11766,N_4614,N_7595);
or U11767 (N_11767,N_6649,N_4221);
or U11768 (N_11768,N_5738,N_4573);
and U11769 (N_11769,N_4411,N_4093);
or U11770 (N_11770,N_5804,N_5763);
nand U11771 (N_11771,N_7429,N_6286);
nor U11772 (N_11772,N_4566,N_4624);
nand U11773 (N_11773,N_6885,N_6559);
and U11774 (N_11774,N_5583,N_6824);
nor U11775 (N_11775,N_7870,N_7092);
and U11776 (N_11776,N_6413,N_4071);
nor U11777 (N_11777,N_7895,N_7134);
or U11778 (N_11778,N_7362,N_5742);
nand U11779 (N_11779,N_6425,N_6522);
nor U11780 (N_11780,N_7250,N_7477);
xor U11781 (N_11781,N_6668,N_4151);
or U11782 (N_11782,N_6835,N_4590);
nor U11783 (N_11783,N_5232,N_5021);
or U11784 (N_11784,N_6467,N_4042);
nor U11785 (N_11785,N_6766,N_5740);
xor U11786 (N_11786,N_5149,N_7502);
nor U11787 (N_11787,N_6439,N_7110);
nand U11788 (N_11788,N_4349,N_6488);
nor U11789 (N_11789,N_6135,N_4901);
nand U11790 (N_11790,N_4243,N_4421);
nor U11791 (N_11791,N_7413,N_6138);
nor U11792 (N_11792,N_6858,N_4533);
and U11793 (N_11793,N_7429,N_6908);
or U11794 (N_11794,N_7124,N_4154);
nor U11795 (N_11795,N_7136,N_7003);
and U11796 (N_11796,N_5185,N_7674);
or U11797 (N_11797,N_4554,N_7680);
or U11798 (N_11798,N_5601,N_5377);
and U11799 (N_11799,N_6292,N_7303);
or U11800 (N_11800,N_6750,N_4387);
or U11801 (N_11801,N_6269,N_5241);
nand U11802 (N_11802,N_5416,N_5669);
nor U11803 (N_11803,N_6232,N_6114);
nand U11804 (N_11804,N_5817,N_6376);
nor U11805 (N_11805,N_7819,N_7384);
and U11806 (N_11806,N_7760,N_6988);
nand U11807 (N_11807,N_7353,N_5297);
nand U11808 (N_11808,N_4088,N_4258);
nor U11809 (N_11809,N_7501,N_4126);
or U11810 (N_11810,N_6198,N_4538);
nor U11811 (N_11811,N_4743,N_7871);
or U11812 (N_11812,N_5018,N_6194);
nor U11813 (N_11813,N_7506,N_4623);
nand U11814 (N_11814,N_6128,N_4065);
or U11815 (N_11815,N_7284,N_6895);
nand U11816 (N_11816,N_5897,N_6225);
and U11817 (N_11817,N_7705,N_5887);
nand U11818 (N_11818,N_6296,N_6811);
nor U11819 (N_11819,N_4115,N_6801);
or U11820 (N_11820,N_4129,N_7069);
or U11821 (N_11821,N_5030,N_4884);
and U11822 (N_11822,N_6743,N_7757);
nor U11823 (N_11823,N_4512,N_4102);
nor U11824 (N_11824,N_6593,N_5220);
and U11825 (N_11825,N_7533,N_5669);
or U11826 (N_11826,N_6798,N_7603);
nor U11827 (N_11827,N_4346,N_6775);
or U11828 (N_11828,N_4217,N_4469);
and U11829 (N_11829,N_5351,N_7619);
nor U11830 (N_11830,N_5116,N_6467);
nor U11831 (N_11831,N_5063,N_6476);
nand U11832 (N_11832,N_6668,N_5287);
nand U11833 (N_11833,N_6287,N_7157);
nand U11834 (N_11834,N_4828,N_6075);
nor U11835 (N_11835,N_4365,N_5480);
nor U11836 (N_11836,N_5543,N_7315);
nand U11837 (N_11837,N_4738,N_5586);
and U11838 (N_11838,N_7734,N_7889);
and U11839 (N_11839,N_5474,N_7090);
and U11840 (N_11840,N_7493,N_6061);
nor U11841 (N_11841,N_6833,N_5834);
and U11842 (N_11842,N_6103,N_5053);
nand U11843 (N_11843,N_7622,N_7024);
and U11844 (N_11844,N_4184,N_5633);
and U11845 (N_11845,N_6068,N_4128);
nor U11846 (N_11846,N_6701,N_6184);
or U11847 (N_11847,N_5176,N_7764);
and U11848 (N_11848,N_7583,N_7200);
nand U11849 (N_11849,N_7961,N_6192);
nor U11850 (N_11850,N_7232,N_7659);
or U11851 (N_11851,N_4257,N_4069);
and U11852 (N_11852,N_5762,N_5541);
nor U11853 (N_11853,N_6130,N_6536);
and U11854 (N_11854,N_4061,N_5539);
nor U11855 (N_11855,N_7923,N_4279);
nor U11856 (N_11856,N_6306,N_4483);
nor U11857 (N_11857,N_6054,N_5330);
or U11858 (N_11858,N_6269,N_7824);
or U11859 (N_11859,N_7537,N_6344);
nor U11860 (N_11860,N_5201,N_5882);
and U11861 (N_11861,N_7472,N_4038);
and U11862 (N_11862,N_7346,N_7907);
nand U11863 (N_11863,N_4270,N_7898);
nand U11864 (N_11864,N_4671,N_5896);
and U11865 (N_11865,N_5924,N_4319);
and U11866 (N_11866,N_7562,N_6499);
or U11867 (N_11867,N_7675,N_4857);
and U11868 (N_11868,N_7623,N_4651);
nand U11869 (N_11869,N_4764,N_7631);
nor U11870 (N_11870,N_6923,N_4634);
and U11871 (N_11871,N_4084,N_6704);
or U11872 (N_11872,N_4912,N_5187);
or U11873 (N_11873,N_4302,N_6483);
nand U11874 (N_11874,N_7666,N_4897);
and U11875 (N_11875,N_4999,N_4488);
or U11876 (N_11876,N_6542,N_7344);
or U11877 (N_11877,N_6500,N_6901);
or U11878 (N_11878,N_5998,N_4991);
nand U11879 (N_11879,N_4239,N_7092);
nor U11880 (N_11880,N_5390,N_4873);
nand U11881 (N_11881,N_6979,N_4676);
nand U11882 (N_11882,N_6776,N_5566);
nand U11883 (N_11883,N_4723,N_7987);
nor U11884 (N_11884,N_7974,N_6229);
nor U11885 (N_11885,N_5101,N_6564);
and U11886 (N_11886,N_5253,N_4881);
and U11887 (N_11887,N_6745,N_6470);
nor U11888 (N_11888,N_6024,N_5723);
nor U11889 (N_11889,N_6798,N_5031);
or U11890 (N_11890,N_6993,N_7506);
or U11891 (N_11891,N_6033,N_5197);
nand U11892 (N_11892,N_6306,N_7313);
nor U11893 (N_11893,N_5347,N_6229);
or U11894 (N_11894,N_7981,N_4507);
nand U11895 (N_11895,N_6638,N_4229);
or U11896 (N_11896,N_4543,N_7451);
or U11897 (N_11897,N_7185,N_4150);
nand U11898 (N_11898,N_4222,N_4133);
or U11899 (N_11899,N_7558,N_6076);
and U11900 (N_11900,N_4591,N_4459);
nand U11901 (N_11901,N_5864,N_5145);
nor U11902 (N_11902,N_6862,N_4126);
or U11903 (N_11903,N_4787,N_5523);
or U11904 (N_11904,N_5335,N_4590);
xnor U11905 (N_11905,N_4464,N_7648);
nand U11906 (N_11906,N_7556,N_5546);
or U11907 (N_11907,N_5152,N_4729);
and U11908 (N_11908,N_5921,N_6726);
or U11909 (N_11909,N_6471,N_6543);
nor U11910 (N_11910,N_7393,N_5587);
and U11911 (N_11911,N_5458,N_5985);
nand U11912 (N_11912,N_5466,N_4454);
nand U11913 (N_11913,N_6170,N_4183);
and U11914 (N_11914,N_5107,N_6966);
nor U11915 (N_11915,N_6076,N_4138);
or U11916 (N_11916,N_6985,N_4231);
and U11917 (N_11917,N_7880,N_7875);
nand U11918 (N_11918,N_7681,N_4222);
nand U11919 (N_11919,N_5308,N_7273);
and U11920 (N_11920,N_4843,N_7284);
nand U11921 (N_11921,N_6979,N_6618);
and U11922 (N_11922,N_6948,N_4781);
nor U11923 (N_11923,N_5872,N_7599);
nand U11924 (N_11924,N_7646,N_7947);
and U11925 (N_11925,N_6812,N_7928);
nor U11926 (N_11926,N_7349,N_4162);
nand U11927 (N_11927,N_5363,N_5527);
nand U11928 (N_11928,N_5572,N_7220);
nor U11929 (N_11929,N_6149,N_4872);
or U11930 (N_11930,N_7752,N_5280);
or U11931 (N_11931,N_6317,N_6732);
and U11932 (N_11932,N_4894,N_7912);
nand U11933 (N_11933,N_4136,N_6037);
nand U11934 (N_11934,N_7710,N_7553);
or U11935 (N_11935,N_4780,N_7357);
nand U11936 (N_11936,N_6014,N_5092);
nor U11937 (N_11937,N_4237,N_6804);
nor U11938 (N_11938,N_4888,N_4293);
and U11939 (N_11939,N_5227,N_7058);
or U11940 (N_11940,N_5829,N_7315);
or U11941 (N_11941,N_7227,N_6668);
nand U11942 (N_11942,N_4220,N_6818);
nand U11943 (N_11943,N_5133,N_4759);
nand U11944 (N_11944,N_5809,N_4619);
nand U11945 (N_11945,N_5373,N_5331);
or U11946 (N_11946,N_7395,N_6062);
nor U11947 (N_11947,N_6654,N_5295);
or U11948 (N_11948,N_7199,N_5768);
nor U11949 (N_11949,N_7712,N_6252);
nand U11950 (N_11950,N_7822,N_5321);
and U11951 (N_11951,N_7814,N_5312);
and U11952 (N_11952,N_7858,N_4045);
nand U11953 (N_11953,N_5088,N_4895);
nor U11954 (N_11954,N_4368,N_6563);
or U11955 (N_11955,N_7454,N_7203);
nor U11956 (N_11956,N_5893,N_6966);
nand U11957 (N_11957,N_5921,N_7144);
nor U11958 (N_11958,N_5351,N_4209);
nand U11959 (N_11959,N_6990,N_6031);
or U11960 (N_11960,N_6051,N_4283);
and U11961 (N_11961,N_7053,N_7652);
nor U11962 (N_11962,N_5302,N_4956);
nor U11963 (N_11963,N_5700,N_7579);
nor U11964 (N_11964,N_7765,N_4803);
nor U11965 (N_11965,N_7082,N_6033);
or U11966 (N_11966,N_5451,N_6611);
or U11967 (N_11967,N_7690,N_4050);
nor U11968 (N_11968,N_5344,N_7540);
and U11969 (N_11969,N_5486,N_7940);
nand U11970 (N_11970,N_6683,N_7733);
or U11971 (N_11971,N_5959,N_7789);
nand U11972 (N_11972,N_5234,N_4047);
and U11973 (N_11973,N_4196,N_5717);
xnor U11974 (N_11974,N_5274,N_6445);
and U11975 (N_11975,N_4831,N_5221);
and U11976 (N_11976,N_6901,N_5253);
or U11977 (N_11977,N_5454,N_6415);
and U11978 (N_11978,N_7013,N_6597);
nand U11979 (N_11979,N_5336,N_4169);
nor U11980 (N_11980,N_5868,N_5209);
or U11981 (N_11981,N_5899,N_6241);
and U11982 (N_11982,N_4904,N_7282);
nand U11983 (N_11983,N_6946,N_6805);
or U11984 (N_11984,N_4260,N_6071);
or U11985 (N_11985,N_7402,N_5665);
or U11986 (N_11986,N_6496,N_4726);
and U11987 (N_11987,N_7441,N_6323);
or U11988 (N_11988,N_7661,N_7835);
nor U11989 (N_11989,N_7994,N_7644);
nor U11990 (N_11990,N_4407,N_4509);
nand U11991 (N_11991,N_7021,N_5039);
nand U11992 (N_11992,N_6288,N_7024);
nor U11993 (N_11993,N_6046,N_7948);
or U11994 (N_11994,N_6577,N_4405);
nand U11995 (N_11995,N_6960,N_4813);
nor U11996 (N_11996,N_6590,N_6378);
nor U11997 (N_11997,N_4430,N_4953);
nor U11998 (N_11998,N_6058,N_7565);
nand U11999 (N_11999,N_7363,N_7906);
nor U12000 (N_12000,N_11208,N_8001);
nor U12001 (N_12001,N_10083,N_9436);
nor U12002 (N_12002,N_11065,N_9565);
nand U12003 (N_12003,N_11491,N_11281);
and U12004 (N_12004,N_10242,N_9474);
and U12005 (N_12005,N_10969,N_8314);
or U12006 (N_12006,N_8974,N_9465);
nor U12007 (N_12007,N_11853,N_9888);
and U12008 (N_12008,N_8643,N_11324);
and U12009 (N_12009,N_10732,N_9812);
or U12010 (N_12010,N_10116,N_8109);
nand U12011 (N_12011,N_10217,N_9306);
and U12012 (N_12012,N_9419,N_11096);
and U12013 (N_12013,N_8791,N_8692);
nand U12014 (N_12014,N_8651,N_8443);
nor U12015 (N_12015,N_9544,N_9904);
nor U12016 (N_12016,N_9412,N_10689);
and U12017 (N_12017,N_11871,N_8341);
or U12018 (N_12018,N_11997,N_11604);
nand U12019 (N_12019,N_10647,N_10776);
nand U12020 (N_12020,N_8076,N_9284);
or U12021 (N_12021,N_9616,N_8259);
or U12022 (N_12022,N_9134,N_10832);
nand U12023 (N_12023,N_11717,N_11756);
and U12024 (N_12024,N_10782,N_9829);
or U12025 (N_12025,N_11473,N_11850);
and U12026 (N_12026,N_8544,N_8801);
nand U12027 (N_12027,N_10106,N_8729);
and U12028 (N_12028,N_9732,N_9550);
nor U12029 (N_12029,N_9190,N_8576);
and U12030 (N_12030,N_8002,N_10025);
and U12031 (N_12031,N_11643,N_9362);
or U12032 (N_12032,N_10265,N_8162);
nand U12033 (N_12033,N_10707,N_10167);
nor U12034 (N_12034,N_11674,N_11825);
nor U12035 (N_12035,N_10912,N_9032);
and U12036 (N_12036,N_11579,N_11092);
or U12037 (N_12037,N_8937,N_8273);
nand U12038 (N_12038,N_9258,N_9885);
nand U12039 (N_12039,N_11452,N_8807);
or U12040 (N_12040,N_11036,N_9212);
xnor U12041 (N_12041,N_9064,N_9648);
nor U12042 (N_12042,N_11721,N_9047);
xor U12043 (N_12043,N_9595,N_10411);
nand U12044 (N_12044,N_8225,N_8233);
or U12045 (N_12045,N_11988,N_8193);
or U12046 (N_12046,N_10501,N_8442);
nand U12047 (N_12047,N_11939,N_8448);
nor U12048 (N_12048,N_11622,N_9516);
and U12049 (N_12049,N_11125,N_9561);
and U12050 (N_12050,N_11738,N_10087);
or U12051 (N_12051,N_8534,N_10416);
nand U12052 (N_12052,N_10539,N_11907);
nor U12053 (N_12053,N_11083,N_11039);
nor U12054 (N_12054,N_10282,N_9122);
nor U12055 (N_12055,N_9752,N_10101);
or U12056 (N_12056,N_9129,N_11440);
nand U12057 (N_12057,N_8201,N_9663);
nand U12058 (N_12058,N_8552,N_8599);
and U12059 (N_12059,N_8247,N_11327);
nor U12060 (N_12060,N_11639,N_8423);
and U12061 (N_12061,N_10724,N_9209);
and U12062 (N_12062,N_10768,N_10955);
nor U12063 (N_12063,N_10481,N_10581);
nor U12064 (N_12064,N_10311,N_9059);
or U12065 (N_12065,N_11856,N_9476);
nand U12066 (N_12066,N_10475,N_10960);
and U12067 (N_12067,N_11681,N_10373);
and U12068 (N_12068,N_10261,N_11922);
and U12069 (N_12069,N_11463,N_10677);
and U12070 (N_12070,N_8391,N_11926);
nor U12071 (N_12071,N_9869,N_10531);
nor U12072 (N_12072,N_10424,N_9243);
and U12073 (N_12073,N_8690,N_11268);
nor U12074 (N_12074,N_10553,N_10409);
nand U12075 (N_12075,N_11492,N_10850);
nand U12076 (N_12076,N_10097,N_9042);
nand U12077 (N_12077,N_10165,N_10488);
and U12078 (N_12078,N_9584,N_11205);
or U12079 (N_12079,N_10734,N_9119);
or U12080 (N_12080,N_11786,N_10253);
or U12081 (N_12081,N_11669,N_11170);
nor U12082 (N_12082,N_9349,N_8802);
nand U12083 (N_12083,N_10438,N_11221);
nor U12084 (N_12084,N_11768,N_9586);
nor U12085 (N_12085,N_10169,N_8988);
and U12086 (N_12086,N_8194,N_8210);
and U12087 (N_12087,N_10917,N_9463);
nand U12088 (N_12088,N_10508,N_8333);
nand U12089 (N_12089,N_10548,N_9100);
nand U12090 (N_12090,N_11619,N_11508);
and U12091 (N_12091,N_10512,N_9001);
or U12092 (N_12092,N_11200,N_10061);
nand U12093 (N_12093,N_9088,N_10194);
nor U12094 (N_12094,N_8593,N_11302);
nand U12095 (N_12095,N_10182,N_9056);
or U12096 (N_12096,N_10991,N_10403);
nand U12097 (N_12097,N_8340,N_8033);
nand U12098 (N_12098,N_10137,N_8600);
nor U12099 (N_12099,N_10994,N_9210);
nand U12100 (N_12100,N_11115,N_8098);
or U12101 (N_12101,N_8517,N_9016);
and U12102 (N_12102,N_8355,N_9542);
or U12103 (N_12103,N_10051,N_10420);
or U12104 (N_12104,N_10399,N_10476);
and U12105 (N_12105,N_9222,N_11692);
nor U12106 (N_12106,N_10212,N_11951);
and U12107 (N_12107,N_8641,N_8778);
nand U12108 (N_12108,N_9720,N_9922);
and U12109 (N_12109,N_8976,N_8920);
nand U12110 (N_12110,N_9235,N_8714);
nand U12111 (N_12111,N_8388,N_9748);
nor U12112 (N_12112,N_9854,N_10546);
nor U12113 (N_12113,N_9859,N_9774);
nand U12114 (N_12114,N_9912,N_10172);
or U12115 (N_12115,N_11316,N_11098);
and U12116 (N_12116,N_9985,N_10159);
and U12117 (N_12117,N_8568,N_11240);
or U12118 (N_12118,N_10002,N_9138);
nor U12119 (N_12119,N_11409,N_10214);
or U12120 (N_12120,N_11539,N_8334);
nor U12121 (N_12121,N_10946,N_9173);
nand U12122 (N_12122,N_9699,N_11304);
or U12123 (N_12123,N_9787,N_8711);
nor U12124 (N_12124,N_9089,N_8515);
or U12125 (N_12125,N_11338,N_9631);
and U12126 (N_12126,N_11472,N_8467);
and U12127 (N_12127,N_9657,N_9624);
nor U12128 (N_12128,N_9940,N_8788);
and U12129 (N_12129,N_8879,N_11074);
nand U12130 (N_12130,N_11760,N_8359);
nand U12131 (N_12131,N_8218,N_10594);
nand U12132 (N_12132,N_10164,N_8881);
or U12133 (N_12133,N_11586,N_8007);
xnor U12134 (N_12134,N_8382,N_9563);
or U12135 (N_12135,N_11362,N_9333);
nand U12136 (N_12136,N_10477,N_11054);
or U12137 (N_12137,N_11553,N_9499);
and U12138 (N_12138,N_10048,N_11724);
or U12139 (N_12139,N_8780,N_11015);
or U12140 (N_12140,N_9283,N_10400);
nand U12141 (N_12141,N_9756,N_10140);
and U12142 (N_12142,N_8762,N_8712);
and U12143 (N_12143,N_10430,N_11565);
nand U12144 (N_12144,N_10341,N_8689);
or U12145 (N_12145,N_9354,N_10323);
and U12146 (N_12146,N_10078,N_10934);
and U12147 (N_12147,N_11912,N_11405);
and U12148 (N_12148,N_10622,N_10777);
or U12149 (N_12149,N_11819,N_10175);
nor U12150 (N_12150,N_8005,N_11053);
nor U12151 (N_12151,N_9831,N_8983);
nand U12152 (N_12152,N_9014,N_8938);
and U12153 (N_12153,N_11864,N_11805);
or U12154 (N_12154,N_9705,N_10979);
and U12155 (N_12155,N_10120,N_9847);
nand U12156 (N_12156,N_11679,N_8962);
or U12157 (N_12157,N_10764,N_8510);
nand U12158 (N_12158,N_9470,N_9842);
or U12159 (N_12159,N_10421,N_10254);
or U12160 (N_12160,N_11902,N_10761);
or U12161 (N_12161,N_11547,N_11718);
and U12162 (N_12162,N_10950,N_10545);
and U12163 (N_12163,N_11900,N_8754);
or U12164 (N_12164,N_10988,N_10263);
nand U12165 (N_12165,N_10088,N_8206);
and U12166 (N_12166,N_9227,N_9447);
nor U12167 (N_12167,N_10931,N_9329);
nand U12168 (N_12168,N_11217,N_10729);
or U12169 (N_12169,N_9039,N_9038);
and U12170 (N_12170,N_11481,N_11211);
nand U12171 (N_12171,N_9634,N_8840);
and U12172 (N_12172,N_11439,N_8349);
nand U12173 (N_12173,N_8494,N_10852);
or U12174 (N_12174,N_9061,N_9311);
and U12175 (N_12175,N_11215,N_8250);
nor U12176 (N_12176,N_11391,N_10580);
nand U12177 (N_12177,N_8065,N_8398);
nand U12178 (N_12178,N_9415,N_10906);
nand U12179 (N_12179,N_11935,N_11204);
xnor U12180 (N_12180,N_9570,N_10465);
or U12181 (N_12181,N_8681,N_8948);
and U12182 (N_12182,N_10679,N_11842);
and U12183 (N_12183,N_11270,N_11796);
nand U12184 (N_12184,N_10069,N_8269);
nand U12185 (N_12185,N_10023,N_8727);
xor U12186 (N_12186,N_11141,N_11872);
nor U12187 (N_12187,N_11859,N_11567);
nor U12188 (N_12188,N_10533,N_11273);
nor U12189 (N_12189,N_9094,N_9576);
or U12190 (N_12190,N_9968,N_8258);
nor U12191 (N_12191,N_11573,N_9074);
nand U12192 (N_12192,N_11342,N_11753);
and U12193 (N_12193,N_10295,N_11929);
nor U12194 (N_12194,N_10805,N_9686);
xor U12195 (N_12195,N_11614,N_10609);
nand U12196 (N_12196,N_8630,N_11169);
nand U12197 (N_12197,N_11851,N_9606);
nor U12198 (N_12198,N_9673,N_9101);
nand U12199 (N_12199,N_11910,N_10305);
and U12200 (N_12200,N_10862,N_10774);
nor U12201 (N_12201,N_10076,N_9133);
and U12202 (N_12202,N_9428,N_10970);
or U12203 (N_12203,N_9203,N_9587);
or U12204 (N_12204,N_11574,N_11442);
nor U12205 (N_12205,N_9972,N_11359);
nand U12206 (N_12206,N_10181,N_8239);
nor U12207 (N_12207,N_10661,N_9568);
nand U12208 (N_12208,N_9521,N_11485);
and U12209 (N_12209,N_11070,N_10247);
nor U12210 (N_12210,N_10506,N_11745);
nand U12211 (N_12211,N_11399,N_8985);
nand U12212 (N_12212,N_11427,N_10352);
or U12213 (N_12213,N_10909,N_8991);
and U12214 (N_12214,N_9057,N_10693);
nand U12215 (N_12215,N_10031,N_8595);
and U12216 (N_12216,N_10132,N_9481);
nor U12217 (N_12217,N_8014,N_9392);
and U12218 (N_12218,N_9638,N_11131);
or U12219 (N_12219,N_9409,N_10691);
nor U12220 (N_12220,N_8179,N_10085);
and U12221 (N_12221,N_10466,N_11400);
or U12222 (N_12222,N_9166,N_9342);
nand U12223 (N_12223,N_9588,N_8796);
and U12224 (N_12224,N_8306,N_9178);
nand U12225 (N_12225,N_10462,N_8091);
nor U12226 (N_12226,N_10745,N_10826);
or U12227 (N_12227,N_11223,N_10814);
or U12228 (N_12228,N_8417,N_8880);
nand U12229 (N_12229,N_10490,N_10220);
and U12230 (N_12230,N_10916,N_8286);
nor U12231 (N_12231,N_8764,N_9023);
or U12232 (N_12232,N_10456,N_8449);
nor U12233 (N_12233,N_9374,N_10904);
or U12234 (N_12234,N_9386,N_8310);
and U12235 (N_12235,N_10928,N_9857);
nor U12236 (N_12236,N_10836,N_9969);
nor U12237 (N_12237,N_9684,N_10747);
nor U12238 (N_12238,N_11934,N_11068);
nor U12239 (N_12239,N_9455,N_8153);
nor U12240 (N_12240,N_8297,N_8939);
and U12241 (N_12241,N_8665,N_9942);
and U12242 (N_12242,N_11725,N_11996);
or U12243 (N_12243,N_10520,N_9421);
nor U12244 (N_12244,N_11720,N_11112);
nand U12245 (N_12245,N_9438,N_9697);
nand U12246 (N_12246,N_9809,N_11960);
nor U12247 (N_12247,N_9537,N_8447);
nand U12248 (N_12248,N_8832,N_8864);
or U12249 (N_12249,N_8242,N_10932);
nand U12250 (N_12250,N_9497,N_11602);
nand U12251 (N_12251,N_8759,N_10933);
or U12252 (N_12252,N_8933,N_8049);
nor U12253 (N_12253,N_9109,N_11874);
nand U12254 (N_12254,N_9769,N_8220);
xnor U12255 (N_12255,N_8722,N_9086);
nand U12256 (N_12256,N_8886,N_9077);
nor U12257 (N_12257,N_11019,N_11801);
or U12258 (N_12258,N_10586,N_8337);
and U12259 (N_12259,N_10020,N_10010);
xnor U12260 (N_12260,N_11630,N_9185);
nand U12261 (N_12261,N_8965,N_8578);
nor U12262 (N_12262,N_9102,N_8543);
and U12263 (N_12263,N_8949,N_9482);
or U12264 (N_12264,N_9641,N_8458);
or U12265 (N_12265,N_8611,N_9739);
and U12266 (N_12266,N_8079,N_10358);
and U12267 (N_12267,N_8397,N_10435);
or U12268 (N_12268,N_9155,N_9211);
or U12269 (N_12269,N_10047,N_8640);
xnor U12270 (N_12270,N_8350,N_11052);
and U12271 (N_12271,N_8083,N_8416);
nor U12272 (N_12272,N_9270,N_10390);
nor U12273 (N_12273,N_10349,N_10627);
and U12274 (N_12274,N_11228,N_8961);
nand U12275 (N_12275,N_8527,N_9823);
nor U12276 (N_12276,N_9949,N_9866);
xor U12277 (N_12277,N_10748,N_8495);
nand U12278 (N_12278,N_9960,N_10381);
and U12279 (N_12279,N_8736,N_10855);
or U12280 (N_12280,N_8374,N_9858);
nor U12281 (N_12281,N_10860,N_8473);
and U12282 (N_12282,N_9139,N_8463);
and U12283 (N_12283,N_10080,N_11153);
or U12284 (N_12284,N_11255,N_11017);
and U12285 (N_12285,N_10587,N_9886);
or U12286 (N_12286,N_11938,N_9669);
and U12287 (N_12287,N_11507,N_9466);
and U12288 (N_12288,N_11562,N_10943);
xor U12289 (N_12289,N_8257,N_9682);
nor U12290 (N_12290,N_10996,N_9099);
and U12291 (N_12291,N_8177,N_11940);
nand U12292 (N_12292,N_8698,N_10013);
and U12293 (N_12293,N_9737,N_9322);
nand U12294 (N_12294,N_10754,N_11608);
and U12295 (N_12295,N_11549,N_9401);
nand U12296 (N_12296,N_10359,N_8503);
or U12297 (N_12297,N_8781,N_8195);
or U12298 (N_12298,N_8246,N_11836);
or U12299 (N_12299,N_9926,N_11116);
or U12300 (N_12300,N_11398,N_11341);
or U12301 (N_12301,N_9344,N_10272);
nor U12302 (N_12302,N_8150,N_9893);
nor U12303 (N_12303,N_9987,N_10337);
or U12304 (N_12304,N_8148,N_9234);
or U12305 (N_12305,N_8276,N_10039);
or U12306 (N_12306,N_9795,N_8241);
nand U12307 (N_12307,N_10460,N_10110);
nand U12308 (N_12308,N_10919,N_8539);
nor U12309 (N_12309,N_10278,N_11531);
or U12310 (N_12310,N_8457,N_8163);
or U12311 (N_12311,N_11194,N_11008);
or U12312 (N_12312,N_10173,N_8236);
and U12313 (N_12313,N_9797,N_8121);
nor U12314 (N_12314,N_11354,N_8512);
or U12315 (N_12315,N_11793,N_10716);
or U12316 (N_12316,N_10316,N_10876);
nand U12317 (N_12317,N_9967,N_8010);
and U12318 (N_12318,N_11297,N_11100);
nor U12319 (N_12319,N_9505,N_11530);
and U12320 (N_12320,N_8378,N_11881);
or U12321 (N_12321,N_9671,N_10090);
or U12322 (N_12322,N_11256,N_8987);
nand U12323 (N_12323,N_8244,N_8016);
and U12324 (N_12324,N_8481,N_11397);
or U12325 (N_12325,N_8929,N_9801);
nand U12326 (N_12326,N_10063,N_10766);
nand U12327 (N_12327,N_8525,N_11883);
or U12328 (N_12328,N_11526,N_10197);
nor U12329 (N_12329,N_10326,N_11954);
or U12330 (N_12330,N_8942,N_10952);
or U12331 (N_12331,N_9053,N_11195);
and U12332 (N_12332,N_8431,N_8070);
nor U12333 (N_12333,N_8363,N_11469);
nor U12334 (N_12334,N_8931,N_8452);
and U12335 (N_12335,N_10752,N_9302);
or U12336 (N_12336,N_9934,N_9667);
and U12337 (N_12337,N_8410,N_9073);
or U12338 (N_12338,N_10470,N_9262);
and U12339 (N_12339,N_9282,N_9772);
or U12340 (N_12340,N_8797,N_8590);
nand U12341 (N_12341,N_11374,N_11182);
or U12342 (N_12342,N_8313,N_8528);
or U12343 (N_12343,N_11072,N_8906);
or U12344 (N_12344,N_11882,N_8436);
nor U12345 (N_12345,N_8655,N_10393);
xnor U12346 (N_12346,N_10050,N_10444);
nor U12347 (N_12347,N_8513,N_8221);
or U12348 (N_12348,N_8584,N_10765);
xnor U12349 (N_12349,N_9848,N_9723);
nor U12350 (N_12350,N_8744,N_8040);
nand U12351 (N_12351,N_11084,N_11828);
nand U12352 (N_12352,N_10666,N_11790);
nor U12353 (N_12353,N_8228,N_8684);
and U12354 (N_12354,N_11321,N_8586);
nand U12355 (N_12355,N_11841,N_8975);
or U12356 (N_12356,N_10221,N_8716);
nand U12357 (N_12357,N_10342,N_10330);
and U12358 (N_12358,N_10593,N_8779);
or U12359 (N_12359,N_11090,N_10074);
and U12360 (N_12360,N_8737,N_10676);
nor U12361 (N_12361,N_9903,N_9397);
and U12362 (N_12362,N_9520,N_10302);
nor U12363 (N_12363,N_11616,N_10551);
nor U12364 (N_12364,N_10985,N_10643);
and U12365 (N_12365,N_8914,N_9698);
or U12366 (N_12366,N_8498,N_9009);
nand U12367 (N_12367,N_9128,N_11632);
nor U12368 (N_12368,N_11584,N_10922);
nand U12369 (N_12369,N_9219,N_9821);
nand U12370 (N_12370,N_9316,N_8717);
and U12371 (N_12371,N_11438,N_11457);
nand U12372 (N_12372,N_10309,N_11502);
nand U12373 (N_12373,N_11818,N_9979);
or U12374 (N_12374,N_10902,N_10821);
and U12375 (N_12375,N_11826,N_10467);
and U12376 (N_12376,N_8955,N_8508);
and U12377 (N_12377,N_10125,N_11612);
or U12378 (N_12378,N_11855,N_11983);
nand U12379 (N_12379,N_8686,N_8856);
and U12380 (N_12380,N_9714,N_10463);
nor U12381 (N_12381,N_8919,N_9670);
nor U12382 (N_12382,N_10603,N_11425);
nor U12383 (N_12383,N_10186,N_11980);
or U12384 (N_12384,N_11587,N_9398);
nand U12385 (N_12385,N_11698,N_11174);
nor U12386 (N_12386,N_8224,N_8414);
or U12387 (N_12387,N_8154,N_11250);
or U12388 (N_12388,N_10151,N_10483);
nand U12389 (N_12389,N_9471,N_9216);
and U12390 (N_12390,N_9148,N_11458);
or U12391 (N_12391,N_11709,N_11747);
and U12392 (N_12392,N_8903,N_10800);
and U12393 (N_12393,N_11928,N_9837);
nand U12394 (N_12394,N_9161,N_8894);
and U12395 (N_12395,N_9054,N_11185);
xor U12396 (N_12396,N_9500,N_11213);
nand U12397 (N_12397,N_10288,N_11060);
and U12398 (N_12398,N_10699,N_10084);
nor U12399 (N_12399,N_10951,N_10901);
nand U12400 (N_12400,N_10735,N_8912);
nand U12401 (N_12401,N_8649,N_10713);
or U12402 (N_12402,N_9553,N_10152);
and U12403 (N_12403,N_11467,N_10495);
nand U12404 (N_12404,N_11641,N_10042);
and U12405 (N_12405,N_11599,N_9592);
or U12406 (N_12406,N_10993,N_10591);
nand U12407 (N_12407,N_11061,N_9759);
or U12408 (N_12408,N_11680,N_9878);
and U12409 (N_12409,N_8637,N_10036);
or U12410 (N_12410,N_11541,N_11411);
nand U12411 (N_12411,N_9524,N_10510);
or U12412 (N_12412,N_9389,N_10290);
or U12413 (N_12413,N_11843,N_9448);
nor U12414 (N_12414,N_9773,N_9376);
nand U12415 (N_12415,N_11772,N_10003);
or U12416 (N_12416,N_10678,N_8361);
and U12417 (N_12417,N_10222,N_10428);
and U12418 (N_12418,N_9399,N_9828);
or U12419 (N_12419,N_10398,N_11689);
or U12420 (N_12420,N_9585,N_8522);
nor U12421 (N_12421,N_9092,N_11050);
nor U12422 (N_12422,N_10953,N_11049);
or U12423 (N_12423,N_11150,N_9323);
or U12424 (N_12424,N_9582,N_8720);
nand U12425 (N_12425,N_11807,N_10705);
nand U12426 (N_12426,N_11198,N_9452);
or U12427 (N_12427,N_9765,N_10480);
nand U12428 (N_12428,N_8260,N_8057);
nor U12429 (N_12429,N_10554,N_10560);
or U12430 (N_12430,N_8144,N_8181);
or U12431 (N_12431,N_9143,N_11333);
and U12432 (N_12432,N_11335,N_8509);
or U12433 (N_12433,N_9492,N_9861);
nand U12434 (N_12434,N_9079,N_9798);
and U12435 (N_12435,N_8324,N_8113);
nor U12436 (N_12436,N_8296,N_11705);
and U12437 (N_12437,N_10174,N_10103);
nand U12438 (N_12438,N_10871,N_8281);
nand U12439 (N_12439,N_11279,N_11287);
xnor U12440 (N_12440,N_8045,N_9704);
or U12441 (N_12441,N_10161,N_9058);
or U12442 (N_12442,N_10812,N_8750);
nand U12443 (N_12443,N_10927,N_8291);
nand U12444 (N_12444,N_8345,N_10778);
nor U12445 (N_12445,N_9902,N_11782);
nand U12446 (N_12446,N_10544,N_11308);
nor U12447 (N_12447,N_9274,N_10243);
or U12448 (N_12448,N_10925,N_10312);
or U12449 (N_12449,N_9220,N_9724);
nor U12450 (N_12450,N_8996,N_9522);
and U12451 (N_12451,N_8472,N_11420);
or U12452 (N_12452,N_9540,N_8116);
or U12453 (N_12453,N_9567,N_9402);
and U12454 (N_12454,N_11212,N_10680);
and U12455 (N_12455,N_8657,N_8678);
nor U12456 (N_12456,N_10503,N_8709);
nand U12457 (N_12457,N_9690,N_9334);
nand U12458 (N_12458,N_11571,N_10308);
and U12459 (N_12459,N_8027,N_8899);
nand U12460 (N_12460,N_10668,N_9215);
nand U12461 (N_12461,N_9931,N_10441);
nor U12462 (N_12462,N_11190,N_10758);
and U12463 (N_12463,N_9367,N_9867);
and U12464 (N_12464,N_8837,N_9764);
nand U12465 (N_12465,N_11637,N_10297);
and U12466 (N_12466,N_8782,N_8580);
nand U12467 (N_12467,N_8497,N_11799);
or U12468 (N_12468,N_10958,N_9110);
nand U12469 (N_12469,N_11184,N_8621);
nor U12470 (N_12470,N_9423,N_9085);
nand U12471 (N_12471,N_11291,N_9011);
nor U12472 (N_12472,N_10740,N_9273);
nor U12473 (N_12473,N_9303,N_9453);
and U12474 (N_12474,N_8031,N_9687);
nand U12475 (N_12475,N_8707,N_11893);
and U12476 (N_12476,N_9218,N_11066);
nor U12477 (N_12477,N_8735,N_11991);
and U12478 (N_12478,N_9836,N_10659);
nand U12479 (N_12479,N_11601,N_9564);
nor U12480 (N_12480,N_11620,N_9906);
nand U12481 (N_12481,N_11834,N_10597);
xor U12482 (N_12482,N_8309,N_9622);
nand U12483 (N_12483,N_10015,N_11513);
nand U12484 (N_12484,N_10339,N_8756);
and U12485 (N_12485,N_9069,N_9791);
nand U12486 (N_12486,N_9048,N_8772);
and U12487 (N_12487,N_8904,N_10634);
nand U12488 (N_12488,N_9223,N_11241);
or U12489 (N_12489,N_11026,N_9070);
nor U12490 (N_12490,N_11787,N_10472);
or U12491 (N_12491,N_11102,N_8390);
or U12492 (N_12492,N_11575,N_10356);
nor U12493 (N_12493,N_10602,N_9735);
nand U12494 (N_12494,N_8989,N_11490);
nor U12495 (N_12495,N_9135,N_9021);
and U12496 (N_12496,N_8574,N_8504);
and U12497 (N_12497,N_10471,N_9924);
or U12498 (N_12498,N_8514,N_9531);
nor U12499 (N_12499,N_9830,N_11424);
or U12500 (N_12500,N_8741,N_8099);
nand U12501 (N_12501,N_8024,N_8289);
nand U12502 (N_12502,N_10303,N_11591);
nor U12503 (N_12503,N_10185,N_11740);
and U12504 (N_12504,N_8900,N_10223);
nand U12505 (N_12505,N_11361,N_11126);
or U12506 (N_12506,N_10639,N_9628);
and U12507 (N_12507,N_9017,N_9287);
nor U12508 (N_12508,N_10853,N_11143);
or U12509 (N_12509,N_11173,N_9962);
or U12510 (N_12510,N_11600,N_8120);
nor U12511 (N_12511,N_8969,N_11367);
or U12512 (N_12512,N_10660,N_11430);
nor U12513 (N_12513,N_10150,N_9664);
nand U12514 (N_12514,N_8170,N_8255);
nor U12515 (N_12515,N_8629,N_10605);
nand U12516 (N_12516,N_9361,N_11501);
nand U12517 (N_12517,N_9062,N_9182);
nand U12518 (N_12518,N_9326,N_10898);
nand U12519 (N_12519,N_11710,N_10549);
nor U12520 (N_12520,N_11414,N_8934);
nand U12521 (N_12521,N_9611,N_8923);
or U12522 (N_12522,N_11564,N_8542);
nor U12523 (N_12523,N_11538,N_10730);
xnor U12524 (N_12524,N_10191,N_10726);
or U12525 (N_12525,N_11583,N_9771);
and U12526 (N_12526,N_9654,N_11258);
and U12527 (N_12527,N_10289,N_11339);
or U12528 (N_12528,N_8097,N_11484);
nor U12529 (N_12529,N_11603,N_8908);
nor U12530 (N_12530,N_8862,N_11334);
or U12531 (N_12531,N_11403,N_9393);
nand U12532 (N_12532,N_9461,N_11237);
nand U12533 (N_12533,N_10314,N_10250);
nor U12534 (N_12534,N_10404,N_11609);
and U12535 (N_12535,N_11965,N_10457);
or U12536 (N_12536,N_8402,N_11970);
and U12537 (N_12537,N_9468,N_8475);
and U12538 (N_12538,N_9029,N_10870);
or U12539 (N_12539,N_8328,N_8317);
or U12540 (N_12540,N_11977,N_8489);
and U12541 (N_12541,N_11272,N_8385);
and U12542 (N_12542,N_11844,N_10771);
nand U12543 (N_12543,N_10062,N_9214);
or U12544 (N_12544,N_11088,N_11719);
nand U12545 (N_12545,N_10474,N_11697);
nand U12546 (N_12546,N_11890,N_9896);
or U12547 (N_12547,N_8956,N_10664);
nor U12548 (N_12548,N_8638,N_9207);
nand U12549 (N_12549,N_11758,N_9041);
nand U12550 (N_12550,N_9272,N_9841);
nand U12551 (N_12551,N_11062,N_8663);
nand U12552 (N_12552,N_11192,N_11920);
or U12553 (N_12553,N_8626,N_8485);
and U12554 (N_12554,N_10102,N_9457);
and U12555 (N_12555,N_9549,N_8563);
and U12556 (N_12556,N_11465,N_8601);
nor U12557 (N_12557,N_10757,N_9117);
or U12558 (N_12558,N_10144,N_8700);
nor U12559 (N_12559,N_9864,N_10837);
or U12560 (N_12560,N_11421,N_11845);
nor U12561 (N_12561,N_10266,N_9145);
xor U12562 (N_12562,N_9418,N_10180);
and U12563 (N_12563,N_9065,N_11498);
and U12564 (N_12564,N_8800,N_10851);
or U12565 (N_12565,N_8981,N_8389);
nand U12566 (N_12566,N_11383,N_8895);
nor U12567 (N_12567,N_10759,N_8178);
and U12568 (N_12568,N_10361,N_9675);
and U12569 (N_12569,N_9484,N_11703);
or U12570 (N_12570,N_9366,N_11108);
nor U12571 (N_12571,N_9758,N_10795);
or U12572 (N_12572,N_9084,N_10787);
nand U12573 (N_12573,N_11822,N_10847);
and U12574 (N_12574,N_11891,N_11447);
nor U12575 (N_12575,N_8827,N_11275);
and U12576 (N_12576,N_8478,N_11524);
and U12577 (N_12577,N_11560,N_8550);
or U12578 (N_12578,N_10281,N_11914);
and U12579 (N_12579,N_8364,N_11838);
nor U12580 (N_12580,N_10355,N_11797);
or U12581 (N_12581,N_10433,N_9839);
and U12582 (N_12582,N_9002,N_10494);
and U12583 (N_12583,N_9424,N_9179);
or U12584 (N_12584,N_10158,N_9925);
nand U12585 (N_12585,N_9037,N_10067);
nand U12586 (N_12586,N_11569,N_11441);
nand U12587 (N_12587,N_8400,N_8810);
and U12588 (N_12588,N_9431,N_8874);
nor U12589 (N_12589,N_8928,N_9341);
or U12590 (N_12590,N_8499,N_8524);
nor U12591 (N_12591,N_10009,N_10880);
nand U12592 (N_12592,N_10442,N_10617);
nand U12593 (N_12593,N_8135,N_9140);
nand U12594 (N_12594,N_8451,N_11777);
nor U12595 (N_12595,N_8435,N_11518);
and U12596 (N_12596,N_8460,N_8476);
and U12597 (N_12597,N_10296,N_9515);
nor U12598 (N_12598,N_9767,N_10949);
nand U12599 (N_12599,N_8365,N_8624);
nor U12600 (N_12600,N_11045,N_9168);
or U12601 (N_12601,N_10057,N_9874);
nand U12602 (N_12602,N_8352,N_9604);
nor U12603 (N_12603,N_10517,N_10208);
or U12604 (N_12604,N_11840,N_9181);
or U12605 (N_12605,N_11369,N_8702);
and U12606 (N_12606,N_10389,N_8824);
nand U12607 (N_12607,N_10267,N_11963);
or U12608 (N_12608,N_8261,N_11732);
and U12609 (N_12609,N_8077,N_8511);
or U12610 (N_12610,N_8723,N_9693);
or U12611 (N_12611,N_10938,N_10802);
nor U12612 (N_12612,N_11109,N_10091);
and U12613 (N_12613,N_9301,N_9248);
and U12614 (N_12614,N_10756,N_10439);
and U12615 (N_12615,N_10986,N_8582);
and U12616 (N_12616,N_10007,N_9808);
nand U12617 (N_12617,N_9933,N_10819);
and U12618 (N_12618,N_11631,N_8264);
or U12619 (N_12619,N_8393,N_11456);
or U12620 (N_12620,N_8480,N_11118);
and U12621 (N_12621,N_10863,N_10882);
or U12622 (N_12622,N_10899,N_10040);
or U12623 (N_12623,N_9937,N_8370);
and U12624 (N_12624,N_11582,N_9034);
nand U12625 (N_12625,N_9835,N_10947);
and U12626 (N_12626,N_8847,N_11487);
and U12627 (N_12627,N_11025,N_9560);
and U12628 (N_12628,N_11043,N_11154);
or U12629 (N_12629,N_9384,N_10717);
nand U12630 (N_12630,N_8585,N_11022);
nor U12631 (N_12631,N_10948,N_8531);
or U12632 (N_12632,N_10577,N_11937);
and U12633 (N_12633,N_8980,N_10446);
or U12634 (N_12634,N_9359,N_10888);
or U12635 (N_12635,N_10537,N_10555);
and U12636 (N_12636,N_8706,N_11848);
or U12637 (N_12637,N_11343,N_9862);
or U12638 (N_12638,N_11982,N_10168);
nor U12639 (N_12639,N_9403,N_8763);
and U12640 (N_12640,N_10072,N_10293);
nor U12641 (N_12641,N_11789,N_10742);
and U12642 (N_12642,N_9992,N_9892);
or U12643 (N_12643,N_8863,N_11358);
or U12644 (N_12644,N_11001,N_8198);
nand U12645 (N_12645,N_11964,N_10064);
nor U12646 (N_12646,N_8811,N_8752);
nand U12647 (N_12647,N_8231,N_10640);
and U12648 (N_12648,N_11806,N_9788);
nand U12649 (N_12649,N_8217,N_8842);
nand U12650 (N_12650,N_9183,N_11536);
or U12651 (N_12651,N_8058,N_11847);
or U12652 (N_12652,N_8533,N_11624);
and U12653 (N_12653,N_10644,N_8598);
nor U12654 (N_12654,N_9512,N_11242);
nand U12655 (N_12655,N_11105,N_9257);
nor U12656 (N_12656,N_10291,N_9003);
and U12657 (N_12657,N_8620,N_11728);
nand U12658 (N_12658,N_11917,N_8693);
or U12659 (N_12659,N_11076,N_8843);
nand U12660 (N_12660,N_8836,N_11879);
xor U12661 (N_12661,N_10744,N_10614);
nand U12662 (N_12662,N_8331,N_11726);
nor U12663 (N_12663,N_8831,N_11685);
and U12664 (N_12664,N_11873,N_11445);
nand U12665 (N_12665,N_11151,N_11089);
or U12666 (N_12666,N_11588,N_11780);
or U12667 (N_12667,N_8013,N_10688);
or U12668 (N_12668,N_9613,N_8559);
and U12669 (N_12669,N_8219,N_8661);
or U12670 (N_12670,N_11464,N_9620);
nor U12671 (N_12671,N_10579,N_10283);
nand U12672 (N_12672,N_8187,N_10383);
nor U12673 (N_12673,N_10279,N_8430);
nor U12674 (N_12674,N_9762,N_8786);
nand U12675 (N_12675,N_10327,N_10975);
nand U12676 (N_12676,N_8612,N_9701);
nand U12677 (N_12677,N_8243,N_11699);
nand U12678 (N_12678,N_10371,N_10633);
nor U12679 (N_12679,N_9027,N_11800);
nor U12680 (N_12680,N_8051,N_11552);
and U12681 (N_12681,N_9727,N_11336);
nor U12682 (N_12682,N_8215,N_9373);
or U12683 (N_12683,N_8588,N_10131);
xor U12684 (N_12684,N_8270,N_10516);
and U12685 (N_12685,N_11157,N_8348);
and U12686 (N_12686,N_11905,N_9413);
or U12687 (N_12687,N_8316,N_8048);
or U12688 (N_12688,N_11433,N_8379);
nor U12689 (N_12689,N_9378,N_8675);
and U12690 (N_12690,N_10041,N_10737);
and U12691 (N_12691,N_9952,N_11875);
or U12692 (N_12692,N_9725,N_8212);
nor U12693 (N_12693,N_9915,N_8158);
nor U12694 (N_12694,N_11323,N_8751);
or U12695 (N_12695,N_10842,N_11128);
and U12696 (N_12696,N_11972,N_8104);
nand U12697 (N_12697,N_11387,N_10978);
nor U12698 (N_12698,N_11653,N_9870);
nor U12699 (N_12699,N_9115,N_10825);
nor U12700 (N_12700,N_11064,N_10017);
or U12701 (N_12701,N_11227,N_10155);
nor U12702 (N_12702,N_8461,N_8890);
nand U12703 (N_12703,N_9261,N_10992);
and U12704 (N_12704,N_10028,N_8086);
nand U12705 (N_12705,N_9558,N_10453);
nor U12706 (N_12706,N_11226,N_10541);
or U12707 (N_12707,N_9763,N_10331);
nand U12708 (N_12708,N_10436,N_10783);
or U12709 (N_12709,N_10822,N_11436);
and U12710 (N_12710,N_9609,N_11349);
and U12711 (N_12711,N_8277,N_11733);
nand U12712 (N_12712,N_10130,N_8562);
and U12713 (N_12713,N_8785,N_8160);
nor U12714 (N_12714,N_10484,N_9196);
nor U12715 (N_12715,N_10763,N_9381);
nor U12716 (N_12716,N_8633,N_9943);
nor U12717 (N_12717,N_9379,N_9899);
nand U12718 (N_12718,N_10332,N_10532);
nor U12719 (N_12719,N_10437,N_10987);
and U12720 (N_12720,N_11776,N_9176);
or U12721 (N_12721,N_11396,N_9615);
nand U12722 (N_12722,N_9260,N_9633);
and U12723 (N_12723,N_11611,N_8392);
or U12724 (N_12724,N_8848,N_11058);
nor U12725 (N_12725,N_10527,N_9443);
nor U12726 (N_12726,N_10892,N_10866);
or U12727 (N_12727,N_10997,N_11244);
nand U12728 (N_12728,N_9126,N_8916);
and U12729 (N_12729,N_8816,N_8570);
nor U12730 (N_12730,N_9517,N_9793);
or U12731 (N_12731,N_10410,N_11662);
or U12732 (N_12732,N_8055,N_11534);
nor U12733 (N_12733,N_11664,N_10630);
nor U12734 (N_12734,N_8950,N_9973);
nor U12735 (N_12735,N_11816,N_9487);
nand U12736 (N_12736,N_8875,N_10671);
or U12737 (N_12737,N_10054,N_11332);
or U12738 (N_12738,N_10388,N_11751);
or U12739 (N_12739,N_9158,N_11921);
nor U12740 (N_12740,N_11328,N_10507);
or U12741 (N_12741,N_9232,N_11379);
nand U12742 (N_12742,N_8743,N_10187);
nor U12743 (N_12743,N_10374,N_10478);
or U12744 (N_12744,N_9004,N_8203);
nor U12745 (N_12745,N_11031,N_10900);
and U12746 (N_12746,N_9060,N_8535);
nand U12747 (N_12747,N_11765,N_8540);
xnor U12748 (N_12748,N_10413,N_11543);
or U12749 (N_12749,N_9394,N_11408);
or U12750 (N_12750,N_10567,N_11781);
or U12751 (N_12751,N_8642,N_9824);
or U12752 (N_12752,N_8635,N_10665);
nor U12753 (N_12753,N_9944,N_11267);
nor U12754 (N_12754,N_9951,N_11953);
or U12755 (N_12755,N_11130,N_9665);
nor U12756 (N_12756,N_10112,N_9519);
nand U12757 (N_12757,N_9033,N_11499);
nor U12758 (N_12758,N_10427,N_9111);
nand U12759 (N_12759,N_10366,N_10698);
nor U12760 (N_12760,N_10372,N_8610);
and U12761 (N_12761,N_10535,N_10770);
and U12762 (N_12762,N_8733,N_10669);
nand U12763 (N_12763,N_9694,N_8304);
or U12764 (N_12764,N_9954,N_9127);
and U12765 (N_12765,N_11529,N_11916);
or U12766 (N_12766,N_9747,N_9891);
nor U12767 (N_12767,N_10963,N_9276);
nand U12768 (N_12768,N_8844,N_10370);
and U12769 (N_12769,N_9642,N_8268);
and U12770 (N_12770,N_9777,N_9480);
and U12771 (N_12771,N_9146,N_11201);
and U12772 (N_12772,N_10701,N_11999);
nand U12773 (N_12773,N_8819,N_10111);
nand U12774 (N_12774,N_10396,N_9177);
nand U12775 (N_12775,N_10251,N_9872);
and U12776 (N_12776,N_11210,N_8288);
nor U12777 (N_12777,N_9731,N_11149);
or U12778 (N_12778,N_8947,N_8335);
nor U12779 (N_12779,N_9445,N_9982);
nor U12780 (N_12780,N_8664,N_11136);
nor U12781 (N_12781,N_10817,N_9729);
and U12782 (N_12782,N_11589,N_8792);
nor U12783 (N_12783,N_11073,N_9796);
xor U12784 (N_12784,N_10872,N_9297);
nand U12785 (N_12785,N_8484,N_10769);
nand U12786 (N_12786,N_9525,N_11550);
or U12787 (N_12787,N_9538,N_9596);
or U12788 (N_12788,N_10710,N_11263);
nor U12789 (N_12789,N_8669,N_8793);
nor U12790 (N_12790,N_9923,N_8644);
nor U12791 (N_12791,N_10071,N_11309);
nand U12792 (N_12792,N_8136,N_10720);
nor U12793 (N_12793,N_11870,N_10809);
nand U12794 (N_12794,N_11628,N_11815);
nor U12795 (N_12795,N_9172,N_8506);
and U12796 (N_12796,N_11471,N_9013);
nor U12797 (N_12797,N_11081,N_8616);
and U12798 (N_12798,N_10686,N_9692);
and U12799 (N_12799,N_11642,N_11968);
nor U12800 (N_12800,N_8553,N_10511);
or U12801 (N_12801,N_9233,N_11007);
nor U12802 (N_12802,N_9348,N_10109);
or U12803 (N_12803,N_10957,N_9820);
nor U12804 (N_12804,N_8926,N_8877);
nand U12805 (N_12805,N_10493,N_8672);
or U12806 (N_12806,N_9330,N_8917);
nand U12807 (N_12807,N_10599,N_11798);
and U12808 (N_12808,N_9849,N_9938);
nor U12809 (N_12809,N_9681,N_10236);
or U12810 (N_12810,N_9430,N_11948);
or U12811 (N_12811,N_11961,N_10449);
or U12812 (N_12812,N_9305,N_10298);
nand U12813 (N_12813,N_11544,N_8992);
and U12814 (N_12814,N_10491,N_9813);
nor U12815 (N_12815,N_8551,N_11598);
and U12816 (N_12816,N_8523,N_8227);
and U12817 (N_12817,N_10199,N_8042);
and U12818 (N_12818,N_11663,N_9832);
nor U12819 (N_12819,N_8411,N_11372);
or U12820 (N_12820,N_9999,N_11752);
nand U12821 (N_12821,N_11650,N_10205);
nand U12822 (N_12822,N_9882,N_11876);
nor U12823 (N_12823,N_8653,N_10881);
and U12824 (N_12824,N_9818,N_9163);
nor U12825 (N_12825,N_9137,N_11122);
nor U12826 (N_12826,N_8953,N_11494);
nor U12827 (N_12827,N_10616,N_9159);
nor U12828 (N_12828,N_11357,N_11158);
or U12829 (N_12829,N_10492,N_9022);
and U12830 (N_12830,N_9990,N_8487);
nand U12831 (N_12831,N_11027,N_9589);
nand U12832 (N_12832,N_11545,N_9715);
and U12833 (N_12833,N_11231,N_8647);
and U12834 (N_12834,N_10108,N_10445);
nor U12835 (N_12835,N_8234,N_10683);
nand U12836 (N_12836,N_10195,N_8977);
xor U12837 (N_12837,N_11597,N_11981);
or U12838 (N_12838,N_8093,N_11278);
nand U12839 (N_12839,N_10415,N_11249);
nor U12840 (N_12840,N_11978,N_10104);
and U12841 (N_12841,N_9575,N_8123);
or U12842 (N_12842,N_8897,N_9000);
nand U12843 (N_12843,N_9467,N_10012);
nor U12844 (N_12844,N_10482,N_9509);
nor U12845 (N_12845,N_10649,N_9192);
and U12846 (N_12846,N_8325,N_8697);
or U12847 (N_12847,N_10380,N_10561);
and U12848 (N_12848,N_8419,N_9573);
or U12849 (N_12849,N_9327,N_11803);
or U12850 (N_12850,N_11312,N_11059);
nand U12851 (N_12851,N_10791,N_10275);
and U12852 (N_12852,N_8787,N_8691);
nor U12853 (N_12853,N_8256,N_8757);
or U12854 (N_12854,N_8927,N_10200);
nor U12855 (N_12855,N_11315,N_9237);
and U12856 (N_12856,N_11775,N_8375);
nand U12857 (N_12857,N_11693,N_11080);
nand U12858 (N_12858,N_8577,N_9939);
nand U12859 (N_12859,N_11269,N_11700);
nand U12860 (N_12860,N_8356,N_11225);
and U12861 (N_12861,N_10935,N_10582);
nor U12862 (N_12862,N_11230,N_10611);
or U12863 (N_12863,N_11171,N_11095);
nor U12864 (N_12864,N_9995,N_10696);
and U12865 (N_12865,N_8347,N_9208);
nand U12866 (N_12866,N_9066,N_10026);
or U12867 (N_12867,N_11915,N_9722);
and U12868 (N_12868,N_10455,N_10937);
or U12869 (N_12869,N_11561,N_9372);
and U12870 (N_12870,N_10391,N_10307);
nand U12871 (N_12871,N_8825,N_9905);
nand U12872 (N_12872,N_10153,N_11943);
nor U12873 (N_12873,N_11504,N_8015);
nand U12874 (N_12874,N_9655,N_10518);
and U12875 (N_12875,N_9559,N_8196);
and U12876 (N_12876,N_11593,N_9935);
or U12877 (N_12877,N_8823,N_11144);
and U12878 (N_12878,N_10498,N_9157);
or U12879 (N_12879,N_11313,N_9898);
and U12880 (N_12880,N_8437,N_11239);
nor U12881 (N_12881,N_8151,N_8701);
nand U12882 (N_12882,N_10121,N_10369);
nor U12883 (N_12883,N_9067,N_10335);
and U12884 (N_12884,N_9434,N_10395);
and U12885 (N_12885,N_9175,N_10971);
nand U12886 (N_12886,N_8742,N_8384);
and U12887 (N_12887,N_11993,N_9541);
or U12888 (N_12888,N_11030,N_9024);
nand U12889 (N_12889,N_9514,N_9097);
nor U12890 (N_12890,N_11288,N_9929);
and U12891 (N_12891,N_11989,N_10114);
and U12892 (N_12892,N_8765,N_11119);
or U12893 (N_12893,N_9807,N_9789);
nor U12894 (N_12894,N_10889,N_8229);
and U12895 (N_12895,N_8770,N_9426);
or U12896 (N_12896,N_8060,N_9251);
and U12897 (N_12897,N_8718,N_9167);
or U12898 (N_12898,N_9745,N_9721);
or U12899 (N_12899,N_11004,N_8902);
nor U12900 (N_12900,N_8748,N_10271);
nand U12901 (N_12901,N_9734,N_9320);
and U12902 (N_12902,N_11021,N_11187);
nand U12903 (N_12903,N_8915,N_9782);
nand U12904 (N_12904,N_8695,N_10458);
nor U12905 (N_12905,N_9608,N_10592);
nand U12906 (N_12906,N_8951,N_8935);
or U12907 (N_12907,N_11975,N_9554);
nand U12908 (N_12908,N_8280,N_9365);
and U12909 (N_12909,N_9685,N_9347);
and U12910 (N_12910,N_8175,N_11480);
or U12911 (N_12911,N_9810,N_9356);
or U12912 (N_12912,N_9130,N_8749);
or U12913 (N_12913,N_10684,N_9383);
or U12914 (N_12914,N_11933,N_8486);
nand U12915 (N_12915,N_8471,N_9229);
and U12916 (N_12916,N_10803,N_10913);
and U12917 (N_12917,N_10552,N_10405);
nand U12918 (N_12918,N_10099,N_10011);
nor U12919 (N_12919,N_10006,N_8833);
nor U12920 (N_12920,N_8518,N_9169);
or U12921 (N_12921,N_10999,N_10100);
nand U12922 (N_12922,N_9425,N_11363);
and U12923 (N_12923,N_11331,N_9932);
nand U12924 (N_12924,N_8739,N_11468);
nor U12925 (N_12925,N_11682,N_10653);
nand U12926 (N_12926,N_8982,N_10454);
or U12927 (N_12927,N_10499,N_8602);
nor U12928 (N_12928,N_11220,N_9275);
nand U12929 (N_12929,N_10721,N_10697);
nor U12930 (N_12930,N_11773,N_9513);
nor U12931 (N_12931,N_8084,N_8569);
nand U12932 (N_12932,N_11956,N_9231);
or U12933 (N_12933,N_11903,N_9191);
and U12934 (N_12934,N_10620,N_11355);
and U12935 (N_12935,N_9689,N_10514);
nand U12936 (N_12936,N_9860,N_10001);
nor U12937 (N_12937,N_10924,N_8368);
nor U12938 (N_12938,N_8004,N_8038);
nand U12939 (N_12939,N_8554,N_10918);
and U12940 (N_12940,N_10575,N_10824);
nand U12941 (N_12941,N_10038,N_10229);
or U12942 (N_12942,N_11412,N_8202);
nor U12943 (N_12943,N_10974,N_11476);
nor U12944 (N_12944,N_11138,N_10094);
or U12945 (N_12945,N_8536,N_11854);
nor U12946 (N_12946,N_8371,N_9385);
nand U12947 (N_12947,N_9785,N_8556);
and U12948 (N_12948,N_9927,N_11094);
or U12949 (N_12949,N_11887,N_9711);
xor U12950 (N_12950,N_9877,N_8166);
nor U12951 (N_12951,N_8829,N_10628);
nor U12952 (N_12952,N_10030,N_9803);
nand U12953 (N_12953,N_8846,N_11647);
nor U12954 (N_12954,N_11152,N_9324);
and U12955 (N_12955,N_9610,N_11423);
nor U12956 (N_12956,N_8000,N_8338);
and U12957 (N_12957,N_10662,N_10672);
nand U12958 (N_12958,N_11114,N_9096);
nor U12959 (N_12959,N_11303,N_8185);
and U12960 (N_12960,N_9153,N_9799);
or U12961 (N_12961,N_8216,N_9494);
nand U12962 (N_12962,N_8089,N_11431);
or U12963 (N_12963,N_10600,N_10722);
nor U12964 (N_12964,N_9307,N_8548);
or U12965 (N_12965,N_11044,N_11389);
and U12966 (N_12966,N_8139,N_8354);
nor U12967 (N_12967,N_10246,N_8687);
nand U12968 (N_12968,N_8835,N_8157);
nor U12969 (N_12969,N_10854,N_11568);
and U12970 (N_12970,N_10000,N_11103);
and U12971 (N_12971,N_11592,N_8235);
or U12972 (N_12972,N_11688,N_9277);
or U12973 (N_12973,N_9965,N_9242);
and U12974 (N_12974,N_11040,N_11318);
nor U12975 (N_12975,N_9802,N_10760);
nand U12976 (N_12976,N_10385,N_9331);
nand U12977 (N_12977,N_11766,N_10419);
nor U12978 (N_12978,N_9406,N_9213);
or U12979 (N_12979,N_10915,N_8403);
or U12980 (N_12980,N_8433,N_11701);
and U12981 (N_12981,N_11962,N_8604);
nand U12982 (N_12982,N_9977,N_8469);
nor U12983 (N_12983,N_8888,N_8190);
and U12984 (N_12984,N_11771,N_9581);
nor U12985 (N_12985,N_9264,N_9627);
and U12986 (N_12986,N_8191,N_8883);
or U12987 (N_12987,N_11657,N_10464);
or U12988 (N_12988,N_9195,N_11958);
or U12989 (N_12989,N_10785,N_10249);
or U12990 (N_12990,N_9293,N_8567);
or U12991 (N_12991,N_10024,N_9853);
nor U12992 (N_12992,N_8838,N_10869);
nor U12993 (N_12993,N_10954,N_10397);
nand U12994 (N_12994,N_8615,N_8973);
or U12995 (N_12995,N_8129,N_10681);
nor U12996 (N_12996,N_11837,N_9188);
and U12997 (N_12997,N_9296,N_8817);
and U12998 (N_12998,N_8117,N_10829);
nand U12999 (N_12999,N_10142,N_10700);
and U13000 (N_13000,N_9408,N_11636);
nand U13001 (N_13001,N_9652,N_11146);
nand U13002 (N_13002,N_10738,N_11265);
and U13003 (N_13003,N_10834,N_11949);
or U13004 (N_13004,N_11941,N_10650);
nand U13005 (N_13005,N_11784,N_8381);
nand U13006 (N_13006,N_9696,N_9717);
or U13007 (N_13007,N_8806,N_8418);
or U13008 (N_13008,N_10566,N_10929);
nand U13009 (N_13009,N_8747,N_11711);
nor U13010 (N_13010,N_8295,N_10032);
nand U13011 (N_13011,N_9919,N_8589);
nand U13012 (N_13012,N_10376,N_10068);
nand U13013 (N_13013,N_10967,N_8761);
nand U13014 (N_13014,N_11888,N_11572);
and U13015 (N_13015,N_8087,N_11140);
or U13016 (N_13016,N_9414,N_10425);
or U13017 (N_13017,N_8857,N_8872);
and U13018 (N_13018,N_11446,N_8294);
nor U13019 (N_13019,N_10285,N_8821);
and U13020 (N_13020,N_11254,N_8940);
nand U13021 (N_13021,N_8870,N_8127);
nor U13022 (N_13022,N_11957,N_9827);
nor U13023 (N_13023,N_11952,N_8979);
or U13024 (N_13024,N_8081,N_8783);
or U13025 (N_13025,N_8252,N_10879);
nor U13026 (N_13026,N_8869,N_11832);
nand U13027 (N_13027,N_11734,N_8538);
nand U13028 (N_13028,N_8432,N_9983);
and U13029 (N_13029,N_10942,N_9049);
nor U13030 (N_13030,N_11159,N_11566);
nand U13031 (N_13031,N_8878,N_11395);
nor U13032 (N_13032,N_8516,N_9617);
nor U13033 (N_13033,N_10619,N_10367);
nor U13034 (N_13034,N_11930,N_8491);
nor U13035 (N_13035,N_8984,N_10711);
and U13036 (N_13036,N_9246,N_9794);
or U13037 (N_13037,N_8775,N_10210);
or U13038 (N_13038,N_11450,N_10234);
or U13039 (N_13039,N_10422,N_11224);
or U13040 (N_13040,N_8892,N_8952);
and U13041 (N_13041,N_9035,N_8103);
nor U13042 (N_13042,N_8734,N_8245);
nor U13043 (N_13043,N_11010,N_10343);
or U13044 (N_13044,N_9974,N_9851);
and U13045 (N_13045,N_9051,N_8966);
and U13046 (N_13046,N_8625,N_11594);
nor U13047 (N_13047,N_8326,N_8813);
and U13048 (N_13048,N_11678,N_10328);
or U13049 (N_13049,N_8572,N_8884);
or U13050 (N_13050,N_9304,N_8130);
nor U13051 (N_13051,N_8998,N_10060);
and U13052 (N_13052,N_8685,N_10695);
or U13053 (N_13053,N_8446,N_9920);
nor U13054 (N_13054,N_9672,N_11390);
nand U13055 (N_13055,N_11521,N_10583);
or U13056 (N_13056,N_11051,N_9569);
nand U13057 (N_13057,N_9112,N_8278);
xor U13058 (N_13058,N_10907,N_9071);
and U13059 (N_13059,N_8732,N_8999);
nand U13060 (N_13060,N_8464,N_9695);
or U13061 (N_13061,N_8809,N_10772);
or U13062 (N_13062,N_11238,N_9946);
nand U13063 (N_13063,N_11849,N_10423);
nand U13064 (N_13064,N_8918,N_8803);
and U13065 (N_13065,N_8358,N_10709);
or U13066 (N_13066,N_8867,N_9632);
or U13067 (N_13067,N_11179,N_10939);
nand U13068 (N_13068,N_9318,N_10798);
nand U13069 (N_13069,N_10572,N_11880);
or U13070 (N_13070,N_11896,N_11134);
nand U13071 (N_13071,N_11908,N_11462);
xor U13072 (N_13072,N_9551,N_9052);
nor U13073 (N_13073,N_10176,N_8932);
nand U13074 (N_13074,N_8253,N_10564);
nand U13075 (N_13075,N_9574,N_11792);
or U13076 (N_13076,N_10417,N_9868);
nand U13077 (N_13077,N_8930,N_9055);
and U13078 (N_13078,N_9015,N_10648);
and U13079 (N_13079,N_8142,N_8332);
nand U13080 (N_13080,N_9957,N_10324);
or U13081 (N_13081,N_11402,N_10313);
nand U13082 (N_13082,N_8165,N_11177);
nand U13083 (N_13083,N_9647,N_8910);
or U13084 (N_13084,N_8575,N_8971);
nand U13085 (N_13085,N_9947,N_11163);
nand U13086 (N_13086,N_9046,N_8866);
and U13087 (N_13087,N_9887,N_11496);
nand U13088 (N_13088,N_11091,N_8406);
nor U13089 (N_13089,N_8924,N_10431);
nor U13090 (N_13090,N_8957,N_8526);
and U13091 (N_13091,N_9749,N_11416);
nand U13092 (N_13092,N_8376,N_11634);
nand U13093 (N_13093,N_8603,N_9335);
nand U13094 (N_13094,N_8439,N_11509);
nor U13095 (N_13095,N_9351,N_11282);
nor U13096 (N_13096,N_11407,N_9025);
nand U13097 (N_13097,N_9479,N_11863);
nor U13098 (N_13098,N_8174,N_11551);
nand U13099 (N_13099,N_10652,N_8581);
nor U13100 (N_13100,N_11444,N_11525);
nor U13101 (N_13101,N_11764,N_8954);
nor U13102 (N_13102,N_11802,N_11489);
or U13103 (N_13103,N_10479,N_9876);
nand U13104 (N_13104,N_8994,N_10828);
and U13105 (N_13105,N_10292,N_11063);
nor U13106 (N_13106,N_10258,N_11337);
and U13107 (N_13107,N_9879,N_8080);
or U13108 (N_13108,N_8850,N_8606);
nor U13109 (N_13109,N_8654,N_8440);
or U13110 (N_13110,N_10235,N_11661);
or U13111 (N_13111,N_11111,N_11835);
or U13112 (N_13112,N_8360,N_8483);
and U13113 (N_13113,N_11590,N_9459);
nand U13114 (N_13114,N_9856,N_9643);
nor U13115 (N_13115,N_8594,N_9761);
nor U13116 (N_13116,N_8232,N_9645);
and U13117 (N_13117,N_10703,N_9151);
nor U13118 (N_13118,N_11459,N_9556);
and U13119 (N_13119,N_9018,N_9478);
and U13120 (N_13120,N_9880,N_8459);
and U13121 (N_13121,N_8674,N_8596);
nand U13122 (N_13122,N_8351,N_10692);
and U13123 (N_13123,N_8020,N_11295);
nand U13124 (N_13124,N_9953,N_8614);
nand U13125 (N_13125,N_9844,N_10233);
nand U13126 (N_13126,N_8566,N_8383);
nor U13127 (N_13127,N_9225,N_10334);
nor U13128 (N_13128,N_11137,N_11483);
or U13129 (N_13129,N_8017,N_11020);
nor U13130 (N_13130,N_9733,N_10301);
xnor U13131 (N_13131,N_9562,N_11723);
and U13132 (N_13132,N_8039,N_9160);
and U13133 (N_13133,N_8342,N_8725);
nor U13134 (N_13134,N_10319,N_10983);
nand U13135 (N_13135,N_11706,N_8455);
nand U13136 (N_13136,N_10815,N_11460);
nor U13137 (N_13137,N_8545,N_10861);
nand U13138 (N_13138,N_10157,N_10117);
nand U13139 (N_13139,N_8003,N_8011);
and U13140 (N_13140,N_10280,N_9713);
nor U13141 (N_13141,N_11559,N_10226);
or U13142 (N_13142,N_8107,N_8683);
nor U13143 (N_13143,N_11535,N_9368);
nor U13144 (N_13144,N_10632,N_8450);
nand U13145 (N_13145,N_11714,N_10329);
and U13146 (N_13146,N_9189,N_9475);
or U13147 (N_13147,N_10521,N_10122);
or U13148 (N_13148,N_8680,N_9125);
nor U13149 (N_13149,N_9598,N_10941);
and U13150 (N_13150,N_8500,N_8226);
nand U13151 (N_13151,N_8794,N_8909);
nand U13152 (N_13152,N_9936,N_9928);
nor U13153 (N_13153,N_9469,N_9198);
nand U13154 (N_13154,N_8054,N_8650);
nor U13155 (N_13155,N_9490,N_8026);
nor U13156 (N_13156,N_9150,N_8262);
nand U13157 (N_13157,N_10751,N_11795);
or U13158 (N_13158,N_8565,N_10663);
or U13159 (N_13159,N_10218,N_10793);
and U13160 (N_13160,N_11329,N_11919);
and U13161 (N_13161,N_9433,N_8758);
and U13162 (N_13162,N_10345,N_9597);
nor U13163 (N_13163,N_9388,N_10304);
nand U13164 (N_13164,N_9072,N_10021);
or U13165 (N_13165,N_10193,N_11517);
nor U13166 (N_13166,N_11904,N_11071);
and U13167 (N_13167,N_8409,N_10375);
nor U13168 (N_13168,N_11186,N_10118);
nor U13169 (N_13169,N_8673,N_8623);
nor U13170 (N_13170,N_10461,N_9845);
nand U13171 (N_13171,N_8632,N_11394);
nor U13172 (N_13172,N_10270,N_11985);
and U13173 (N_13173,N_10723,N_11037);
nand U13174 (N_13174,N_10995,N_8143);
or U13175 (N_13175,N_11046,N_11932);
and U13176 (N_13176,N_8019,N_9131);
nand U13177 (N_13177,N_11527,N_11746);
nor U13178 (N_13178,N_10273,N_11969);
or U13179 (N_13179,N_10027,N_8936);
and U13180 (N_13180,N_8429,N_10202);
nand U13181 (N_13181,N_9291,N_9741);
nand U13182 (N_13182,N_9709,N_9477);
nand U13183 (N_13183,N_11615,N_10811);
nand U13184 (N_13184,N_8028,N_11546);
or U13185 (N_13185,N_10718,N_9660);
nand U13186 (N_13186,N_11715,N_9778);
and U13187 (N_13187,N_10382,N_11093);
nor U13188 (N_13188,N_11548,N_10613);
or U13189 (N_13189,N_8186,N_9429);
nor U13190 (N_13190,N_10841,N_10244);
and U13191 (N_13191,N_9290,N_10198);
or U13192 (N_13192,N_10618,N_8688);
nand U13193 (N_13193,N_10127,N_9464);
nor U13194 (N_13194,N_11892,N_11032);
nand U13195 (N_13195,N_11514,N_11175);
and U13196 (N_13196,N_10364,N_10767);
or U13197 (N_13197,N_11280,N_10801);
nor U13198 (N_13198,N_9825,N_11923);
or U13199 (N_13199,N_11754,N_9325);
nor U13200 (N_13200,N_9020,N_11757);
and U13201 (N_13201,N_10596,N_11635);
nor U13202 (N_13202,N_9486,N_8366);
and U13203 (N_13203,N_11648,N_10145);
nand U13204 (N_13204,N_10412,N_8052);
nand U13205 (N_13205,N_9114,N_10274);
nand U13206 (N_13206,N_8205,N_8986);
nor U13207 (N_13207,N_9751,N_9612);
nand U13208 (N_13208,N_11627,N_10418);
nand U13209 (N_13209,N_10287,N_8826);
nor U13210 (N_13210,N_10890,N_8815);
nor U13211 (N_13211,N_8468,N_8453);
nand U13212 (N_13212,N_8549,N_11376);
and U13213 (N_13213,N_11886,N_10598);
and U13214 (N_13214,N_9450,N_11352);
and U13215 (N_13215,N_11783,N_11884);
and U13216 (N_13216,N_8362,N_8428);
nand U13217 (N_13217,N_11386,N_8860);
nand U13218 (N_13218,N_10790,N_9204);
and U13219 (N_13219,N_8845,N_9712);
nand U13220 (N_13220,N_11077,N_11651);
or U13221 (N_13221,N_10610,N_10753);
or U13222 (N_13222,N_8605,N_11435);
nand U13223 (N_13223,N_9352,N_10190);
and U13224 (N_13224,N_9404,N_8085);
or U13225 (N_13225,N_10578,N_8882);
or U13226 (N_13226,N_9911,N_8426);
nor U13227 (N_13227,N_11713,N_8959);
and U13228 (N_13228,N_10123,N_10725);
and U13229 (N_13229,N_10333,N_11247);
nor U13230 (N_13230,N_9377,N_11668);
or U13231 (N_13231,N_9590,N_9783);
nor U13232 (N_13232,N_8583,N_9651);
nor U13233 (N_13233,N_9491,N_10284);
nor U13234 (N_13234,N_9572,N_10538);
nand U13235 (N_13235,N_11676,N_8789);
nor U13236 (N_13236,N_9528,N_9105);
nand U13237 (N_13237,N_10089,N_8479);
or U13238 (N_13238,N_9583,N_11808);
xnor U13239 (N_13239,N_9104,N_8199);
and U13240 (N_13240,N_8704,N_11704);
nand U13241 (N_13241,N_11942,N_11207);
nor U13242 (N_13242,N_9950,N_9579);
and U13243 (N_13243,N_10746,N_10049);
or U13244 (N_13244,N_9076,N_9976);
and U13245 (N_13245,N_8373,N_11821);
nand U13246 (N_13246,N_11317,N_8035);
nand U13247 (N_13247,N_10896,N_11511);
or U13248 (N_13248,N_10154,N_8275);
and U13249 (N_13249,N_8705,N_11984);
nand U13250 (N_13250,N_9141,N_8346);
nand U13251 (N_13251,N_11404,N_9193);
nor U13252 (N_13252,N_9786,N_11618);
or U13253 (N_13253,N_10874,N_10225);
or U13254 (N_13254,N_8339,N_8071);
and U13255 (N_13255,N_8272,N_9081);
nor U13256 (N_13256,N_9504,N_9005);
nor U13257 (N_13257,N_11846,N_8043);
and U13258 (N_13258,N_11129,N_10973);
and U13259 (N_13259,N_11563,N_9010);
nand U13260 (N_13260,N_10959,N_8132);
or U13261 (N_13261,N_11644,N_8456);
nand U13262 (N_13262,N_11448,N_8062);
and U13263 (N_13263,N_8183,N_10624);
or U13264 (N_13264,N_11665,N_9508);
nand U13265 (N_13265,N_11028,N_10056);
nor U13266 (N_13266,N_11301,N_10522);
nor U13267 (N_13267,N_9909,N_9980);
and U13268 (N_13268,N_10806,N_10886);
or U13269 (N_13269,N_9790,N_9439);
and U13270 (N_13270,N_11191,N_11722);
nand U13271 (N_13271,N_11348,N_10559);
or U13272 (N_13272,N_9811,N_9350);
xnor U13273 (N_13273,N_11012,N_11580);
or U13274 (N_13274,N_9552,N_11296);
and U13275 (N_13275,N_11833,N_8138);
or U13276 (N_13276,N_11690,N_9991);
and U13277 (N_13277,N_11523,N_10868);
or U13278 (N_13278,N_8876,N_11809);
nand U13279 (N_13279,N_9623,N_11606);
nor U13280 (N_13280,N_8871,N_11041);
and U13281 (N_13281,N_10394,N_8030);
or U13282 (N_13282,N_8521,N_11537);
nand U13283 (N_13283,N_10820,N_8126);
nor U13284 (N_13284,N_10447,N_9206);
nand U13285 (N_13285,N_10816,N_8887);
or U13286 (N_13286,N_9964,N_9165);
and U13287 (N_13287,N_9007,N_10576);
nand U13288 (N_13288,N_8591,N_10945);
nor U13289 (N_13289,N_11913,N_8474);
nor U13290 (N_13290,N_8715,N_11056);
nor U13291 (N_13291,N_11142,N_8865);
nor U13292 (N_13292,N_9371,N_11533);
or U13293 (N_13293,N_8021,N_10505);
nor U13294 (N_13294,N_11162,N_10093);
nand U13295 (N_13295,N_11283,N_8646);
or U13296 (N_13296,N_10623,N_8958);
nand U13297 (N_13297,N_8046,N_8301);
nand U13298 (N_13298,N_8141,N_11121);
nand U13299 (N_13299,N_8719,N_11432);
nand U13300 (N_13300,N_9288,N_9152);
or U13301 (N_13301,N_11585,N_9454);
nand U13302 (N_13302,N_11262,N_8405);
and U13303 (N_13303,N_8114,N_10259);
nor U13304 (N_13304,N_10773,N_11276);
and U13305 (N_13305,N_11311,N_11451);
or U13306 (N_13306,N_9440,N_9901);
nor U13307 (N_13307,N_10797,N_10547);
or U13308 (N_13308,N_8609,N_10584);
nand U13309 (N_13309,N_10524,N_11286);
nand U13310 (N_13310,N_11936,N_9106);
or U13311 (N_13311,N_9781,N_11625);
and U13312 (N_13312,N_8188,N_10989);
and U13313 (N_13313,N_11762,N_11749);
nand U13314 (N_13314,N_8266,N_9147);
nor U13315 (N_13315,N_8799,N_8176);
nor U13316 (N_13316,N_8659,N_9535);
and U13317 (N_13317,N_8462,N_10972);
or U13318 (N_13318,N_9435,N_11621);
and U13319 (N_13319,N_11737,N_11124);
nand U13320 (N_13320,N_9894,N_10574);
nand U13321 (N_13321,N_8907,N_10818);
and U13322 (N_13322,N_8771,N_10136);
nand U13323 (N_13323,N_10487,N_9895);
and U13324 (N_13324,N_11744,N_9963);
and U13325 (N_13325,N_10750,N_10231);
nand U13326 (N_13326,N_8111,N_10306);
or U13327 (N_13327,N_9742,N_11172);
or U13328 (N_13328,N_8855,N_9819);
or U13329 (N_13329,N_11878,N_11944);
or U13330 (N_13330,N_11417,N_10556);
and U13331 (N_13331,N_11673,N_10590);
and U13332 (N_13332,N_8204,N_9012);
or U13333 (N_13333,N_10035,N_11257);
nor U13334 (N_13334,N_9422,N_11113);
and U13335 (N_13335,N_9315,N_10256);
nand U13336 (N_13336,N_8161,N_9577);
nor U13337 (N_13337,N_10322,N_9473);
nand U13338 (N_13338,N_8315,N_9566);
and U13339 (N_13339,N_9044,N_8412);
or U13340 (N_13340,N_9666,N_8380);
nor U13341 (N_13341,N_9154,N_9996);
nor U13342 (N_13342,N_9599,N_9171);
or U13343 (N_13343,N_10893,N_9501);
nor U13344 (N_13344,N_8738,N_11428);
nand U13345 (N_13345,N_10702,N_9411);
and U13346 (N_13346,N_8438,N_10897);
nand U13347 (N_13347,N_10079,N_11222);
and U13348 (N_13348,N_10362,N_11419);
and U13349 (N_13349,N_10563,N_8282);
nor U13350 (N_13350,N_8149,N_10651);
or U13351 (N_13351,N_10529,N_11708);
or U13352 (N_13352,N_11406,N_10320);
and U13353 (N_13353,N_10053,N_10486);
nor U13354 (N_13354,N_10058,N_10146);
or U13355 (N_13355,N_11729,N_11474);
nor U13356 (N_13356,N_11346,N_9170);
nor U13357 (N_13357,N_9834,N_9988);
nand U13358 (N_13358,N_9780,N_11865);
and U13359 (N_13359,N_9545,N_11418);
or U13360 (N_13360,N_9328,N_8263);
and U13361 (N_13361,N_9241,N_8444);
nand U13362 (N_13362,N_11823,N_9346);
and U13363 (N_13363,N_9826,N_10965);
or U13364 (N_13364,N_11994,N_8564);
and U13365 (N_13365,N_10550,N_8125);
and U13366 (N_13366,N_11743,N_11788);
xor U13367 (N_13367,N_8645,N_10357);
and U13368 (N_13368,N_11770,N_11897);
nor U13369 (N_13369,N_11351,N_10911);
nand U13370 (N_13370,N_10621,N_11345);
or U13371 (N_13371,N_8617,N_11830);
or U13372 (N_13372,N_9555,N_8943);
nor U13373 (N_13373,N_9852,N_9239);
nand U13374 (N_13374,N_11512,N_8108);
and U13375 (N_13375,N_11079,N_10694);
and U13376 (N_13376,N_8767,N_11794);
and U13377 (N_13377,N_10903,N_10673);
and U13378 (N_13378,N_11901,N_8037);
and U13379 (N_13379,N_8898,N_11486);
or U13380 (N_13380,N_11646,N_9360);
nor U13381 (N_13381,N_8636,N_11804);
and U13382 (N_13382,N_10891,N_9493);
or U13383 (N_13383,N_11307,N_10607);
nor U13384 (N_13384,N_11219,N_11640);
nor U13385 (N_13385,N_10864,N_11364);
nand U13386 (N_13386,N_10865,N_8271);
nor U13387 (N_13387,N_8995,N_11482);
xnor U13388 (N_13388,N_11086,N_10914);
nand U13389 (N_13389,N_11139,N_11478);
nand U13390 (N_13390,N_9618,N_11147);
or U13391 (N_13391,N_11924,N_10264);
or U13392 (N_13392,N_9728,N_8618);
and U13393 (N_13393,N_11667,N_8798);
or U13394 (N_13394,N_11931,N_11686);
and U13395 (N_13395,N_10045,N_8300);
and U13396 (N_13396,N_11761,N_10318);
nor U13397 (N_13397,N_9653,N_10070);
and U13398 (N_13398,N_11097,N_8597);
nor U13399 (N_13399,N_9768,N_10496);
xor U13400 (N_13400,N_10908,N_8357);
and U13401 (N_13401,N_8941,N_9706);
nand U13402 (N_13402,N_9776,N_9917);
nand U13403 (N_13403,N_8329,N_10392);
and U13404 (N_13404,N_8507,N_11437);
and U13405 (N_13405,N_11857,N_9571);
nand U13406 (N_13406,N_8997,N_10241);
and U13407 (N_13407,N_9910,N_10469);
xor U13408 (N_13408,N_8639,N_11885);
or U13409 (N_13409,N_9530,N_11750);
and U13410 (N_13410,N_9873,N_10608);
nor U13411 (N_13411,N_8561,N_11694);
nand U13412 (N_13412,N_8396,N_10277);
nor U13413 (N_13413,N_8067,N_9815);
nor U13414 (N_13414,N_8214,N_10134);
nand U13415 (N_13415,N_11326,N_11898);
nand U13416 (N_13416,N_10601,N_11998);
or U13417 (N_13417,N_8292,N_11918);
nor U13418 (N_13418,N_9738,N_9770);
and U13419 (N_13419,N_10119,N_11895);
nor U13420 (N_13420,N_11375,N_9661);
or U13421 (N_13421,N_10065,N_9658);
nand U13422 (N_13422,N_10473,N_9364);
and U13423 (N_13423,N_8769,N_10252);
or U13424 (N_13424,N_10401,N_8424);
nand U13425 (N_13425,N_10804,N_11666);
nand U13426 (N_13426,N_8501,N_10792);
or U13427 (N_13427,N_9529,N_11677);
or U13428 (N_13428,N_8490,N_11990);
nor U13429 (N_13429,N_10310,N_9298);
or U13430 (N_13430,N_10018,N_10485);
nand U13431 (N_13431,N_8036,N_8859);
or U13432 (N_13432,N_10107,N_11947);
or U13433 (N_13433,N_11992,N_10354);
nand U13434 (N_13434,N_9164,N_11735);
nor U13435 (N_13435,N_9619,N_9006);
and U13436 (N_13436,N_8299,N_8658);
or U13437 (N_13437,N_10571,N_11009);
nor U13438 (N_13438,N_8182,N_11078);
and U13439 (N_13439,N_9908,N_9136);
and U13440 (N_13440,N_9255,N_10452);
nand U13441 (N_13441,N_10883,N_11160);
or U13442 (N_13442,N_8213,N_9792);
nor U13443 (N_13443,N_8237,N_11506);
nand U13444 (N_13444,N_9547,N_10325);
or U13445 (N_13445,N_8323,N_9390);
and U13446 (N_13446,N_10636,N_10799);
nor U13447 (N_13447,N_10685,N_10196);
nor U13448 (N_13448,N_11755,N_11684);
nand U13449 (N_13449,N_11607,N_10936);
and U13450 (N_13450,N_9662,N_9149);
or U13451 (N_13451,N_11360,N_11687);
nor U13452 (N_13452,N_9495,N_9420);
nor U13453 (N_13453,N_9269,N_8100);
nor U13454 (N_13454,N_10075,N_10655);
nor U13455 (N_13455,N_9236,N_9083);
and U13456 (N_13456,N_11812,N_9914);
nand U13457 (N_13457,N_8372,N_11271);
nor U13458 (N_13458,N_11974,N_10269);
nor U13459 (N_13459,N_9975,N_11373);
and U13460 (N_13460,N_8096,N_9503);
or U13461 (N_13461,N_8110,N_9649);
nand U13462 (N_13462,N_10082,N_9082);
nand U13463 (N_13463,N_9405,N_10232);
or U13464 (N_13464,N_8069,N_8679);
or U13465 (N_13465,N_8911,N_9483);
nand U13466 (N_13466,N_8106,N_11161);
or U13467 (N_13467,N_8238,N_8652);
or U13468 (N_13468,N_9496,N_8427);
nand U13469 (N_13469,N_10706,N_11862);
nor U13470 (N_13470,N_8171,N_9295);
nor U13471 (N_13471,N_11422,N_11774);
nand U13472 (N_13472,N_11202,N_8901);
nand U13473 (N_13473,N_8408,N_10631);
nor U13474 (N_13474,N_8386,N_9907);
nor U13475 (N_13475,N_8147,N_8724);
or U13476 (N_13476,N_8413,N_9108);
nand U13477 (N_13477,N_8537,N_11670);
or U13478 (N_13478,N_9629,N_10350);
nand U13479 (N_13479,N_9640,N_11867);
or U13480 (N_13480,N_11370,N_8682);
or U13481 (N_13481,N_8828,N_11655);
nor U13482 (N_13482,N_9313,N_10224);
and U13483 (N_13483,N_8094,N_10962);
nor U13484 (N_13484,N_10387,N_10429);
nor U13485 (N_13485,N_9833,N_11658);
nor U13486 (N_13486,N_10923,N_9441);
or U13487 (N_13487,N_11294,N_8726);
nor U13488 (N_13488,N_10384,N_9278);
nand U13489 (N_13489,N_11739,N_9916);
or U13490 (N_13490,N_10029,N_8970);
xor U13491 (N_13491,N_10340,N_10239);
and U13492 (N_13492,N_11216,N_9594);
nand U13493 (N_13493,N_10426,N_11477);
nand U13494 (N_13494,N_9031,N_8211);
or U13495 (N_13495,N_10675,N_10353);
nand U13496 (N_13496,N_11251,N_8189);
and U13497 (N_13497,N_11495,N_9614);
or U13498 (N_13498,N_10414,N_10743);
and U13499 (N_13499,N_9312,N_9626);
and U13500 (N_13500,N_11986,N_10588);
or U13501 (N_13501,N_11814,N_9656);
or U13502 (N_13502,N_10786,N_11214);
nand U13503 (N_13503,N_11528,N_9132);
or U13504 (N_13504,N_10562,N_8730);
nand U13505 (N_13505,N_8265,N_10823);
or U13506 (N_13506,N_10885,N_10344);
nor U13507 (N_13507,N_8441,N_8818);
and U13508 (N_13508,N_11347,N_10019);
and U13509 (N_13509,N_10497,N_8415);
and U13510 (N_13510,N_9263,N_9358);
and U13511 (N_13511,N_8804,N_8731);
nor U13512 (N_13512,N_8868,N_10595);
and U13513 (N_13513,N_11183,N_11542);
or U13514 (N_13514,N_11382,N_9708);
or U13515 (N_13515,N_9718,N_9268);
nand U13516 (N_13516,N_11290,N_9030);
or U13517 (N_13517,N_9279,N_11475);
and U13518 (N_13518,N_9319,N_8267);
and U13519 (N_13519,N_11252,N_11488);
and U13520 (N_13520,N_11246,N_8336);
nor U13521 (N_13521,N_10887,N_8555);
or U13522 (N_13522,N_10878,N_8972);
nor U13523 (N_13523,N_9913,N_8131);
or U13524 (N_13524,N_10379,N_11946);
nor U13525 (N_13525,N_9080,N_11652);
nand U13526 (N_13526,N_9703,N_9343);
nand U13527 (N_13527,N_11085,N_9314);
nand U13528 (N_13528,N_8032,N_8713);
or U13529 (N_13529,N_10844,N_10162);
and U13530 (N_13530,N_10201,N_9889);
and U13531 (N_13531,N_11736,N_11261);
and U13532 (N_13532,N_10877,N_9308);
nand U13533 (N_13533,N_9400,N_11284);
or U13534 (N_13534,N_9118,N_11516);
nor U13535 (N_13535,N_8851,N_11029);
nand U13536 (N_13536,N_11769,N_9040);
xnor U13537 (N_13537,N_9750,N_9201);
nand U13538 (N_13538,N_8008,N_9395);
and U13539 (N_13539,N_9945,N_10827);
or U13540 (N_13540,N_11945,N_9814);
nor U13541 (N_13541,N_11810,N_8834);
nor U13542 (N_13542,N_8128,N_8557);
nor U13543 (N_13543,N_8249,N_11515);
nor U13544 (N_13544,N_9416,N_10052);
and U13545 (N_13545,N_8377,N_11443);
and U13546 (N_13546,N_8422,N_8493);
nor U13547 (N_13547,N_8852,N_8579);
and U13548 (N_13548,N_10557,N_10645);
and U13549 (N_13549,N_8248,N_11378);
or U13550 (N_13550,N_9357,N_9956);
nor U13551 (N_13551,N_9716,N_9382);
nor U13552 (N_13552,N_9726,N_10407);
nand U13553 (N_13553,N_11274,N_9087);
or U13554 (N_13554,N_8327,N_9244);
or U13555 (N_13555,N_8353,N_9205);
nor U13556 (N_13556,N_11617,N_9187);
nor U13557 (N_13557,N_8619,N_10894);
or U13558 (N_13558,N_10095,N_10124);
and U13559 (N_13559,N_10004,N_10300);
nor U13560 (N_13560,N_9997,N_8230);
nand U13561 (N_13561,N_10450,N_9271);
and U13562 (N_13562,N_10589,N_10406);
nand U13563 (N_13563,N_10749,N_8668);
or U13564 (N_13564,N_9174,N_9636);
or U13565 (N_13565,N_10736,N_8861);
and U13566 (N_13566,N_8627,N_11966);
or U13567 (N_13567,N_11069,N_9387);
and U13568 (N_13568,N_10166,N_9507);
nor U13569 (N_13569,N_10755,N_11023);
or U13570 (N_13570,N_9659,N_9026);
or U13571 (N_13571,N_8822,N_10286);
nand U13572 (N_13572,N_10081,N_9285);
or U13573 (N_13573,N_11558,N_8063);
or U13574 (N_13574,N_8044,N_10833);
or U13575 (N_13575,N_11791,N_11626);
or U13576 (N_13576,N_9337,N_11659);
xnor U13577 (N_13577,N_10245,N_8466);
and U13578 (N_13578,N_10073,N_10096);
xor U13579 (N_13579,N_9294,N_8660);
nor U13580 (N_13580,N_11540,N_10338);
nor U13581 (N_13581,N_8746,N_10238);
nand U13582 (N_13582,N_10543,N_9224);
and U13583 (N_13583,N_8180,N_10530);
nor U13584 (N_13584,N_9321,N_11767);
and U13585 (N_13585,N_8571,N_9396);
nor U13586 (N_13586,N_8776,N_9986);
or U13587 (N_13587,N_11340,N_9280);
or U13588 (N_13588,N_9250,N_10378);
and U13589 (N_13589,N_8774,N_8922);
nor U13590 (N_13590,N_8387,N_11505);
nand U13591 (N_13591,N_11322,N_10143);
nor U13592 (N_13592,N_11013,N_11117);
nor U13593 (N_13593,N_10260,N_8529);
nor U13594 (N_13594,N_9238,N_9630);
xor U13595 (N_13595,N_8240,N_10982);
and U13596 (N_13596,N_10926,N_10113);
xor U13597 (N_13597,N_9506,N_11556);
nor U13598 (N_13598,N_10839,N_10848);
or U13599 (N_13599,N_8012,N_11218);
or U13600 (N_13600,N_9676,N_9098);
nand U13601 (N_13601,N_8041,N_8921);
or U13602 (N_13602,N_11748,N_11730);
nand U13603 (N_13603,N_10712,N_11319);
xor U13604 (N_13604,N_10204,N_8330);
or U13605 (N_13605,N_11048,N_9338);
and U13606 (N_13606,N_10542,N_8694);
nor U13607 (N_13607,N_8133,N_11955);
and U13608 (N_13608,N_11696,N_8112);
nand U13609 (N_13609,N_10178,N_9410);
nor U13610 (N_13610,N_9674,N_10604);
and U13611 (N_13611,N_9678,N_8343);
or U13612 (N_13612,N_9800,N_10775);
or U13613 (N_13613,N_11434,N_9370);
nor U13614 (N_13614,N_8293,N_11320);
nor U13615 (N_13615,N_10895,N_9650);
nand U13616 (N_13616,N_8092,N_9226);
nand U13617 (N_13617,N_10654,N_11206);
nand U13618 (N_13618,N_10921,N_11950);
nand U13619 (N_13619,N_8222,N_10219);
nor U13620 (N_13620,N_11155,N_8766);
and U13621 (N_13621,N_8197,N_10315);
nor U13622 (N_13622,N_11877,N_8303);
nor U13623 (N_13623,N_11299,N_9228);
nand U13624 (N_13624,N_9472,N_9755);
nor U13625 (N_13625,N_10184,N_8407);
nand U13626 (N_13626,N_8140,N_9121);
or U13627 (N_13627,N_10568,N_10739);
or U13628 (N_13628,N_11181,N_9532);
nand U13629 (N_13629,N_11236,N_11429);
and U13630 (N_13630,N_8849,N_11577);
nand U13631 (N_13631,N_10719,N_9502);
nand U13632 (N_13632,N_9966,N_11785);
and U13633 (N_13633,N_9677,N_10014);
and U13634 (N_13634,N_8134,N_11702);
nand U13635 (N_13635,N_9510,N_8145);
and U13636 (N_13636,N_8006,N_9806);
nor U13637 (N_13637,N_11285,N_11581);
and U13638 (N_13638,N_9310,N_8677);
nor U13639 (N_13639,N_10859,N_10526);
and U13640 (N_13640,N_10105,N_10704);
and U13641 (N_13641,N_9336,N_8082);
or U13642 (N_13642,N_8078,N_11166);
nor U13643 (N_13643,N_9989,N_11306);
or U13644 (N_13644,N_8755,N_9784);
nand U13645 (N_13645,N_8029,N_9897);
or U13646 (N_13646,N_11660,N_10569);
nand U13647 (N_13647,N_10443,N_8305);
or U13648 (N_13648,N_10794,N_10171);
nand U13649 (N_13649,N_9635,N_9900);
nand U13650 (N_13650,N_10346,N_11057);
or U13651 (N_13651,N_11454,N_10055);
nor U13652 (N_13652,N_10741,N_11519);
xnor U13653 (N_13653,N_9994,N_8283);
nand U13654 (N_13654,N_8896,N_11178);
or U13655 (N_13655,N_11497,N_8622);
nor U13656 (N_13656,N_10046,N_10149);
nor U13657 (N_13657,N_11987,N_11868);
or U13658 (N_13658,N_9602,N_11675);
nor U13659 (N_13659,N_10715,N_9518);
and U13660 (N_13660,N_10796,N_8968);
nand U13661 (N_13661,N_8945,N_9883);
and U13662 (N_13662,N_10188,N_8913);
nand U13663 (N_13663,N_10944,N_9462);
nor U13664 (N_13664,N_9197,N_8505);
nor U13665 (N_13665,N_10177,N_9489);
or U13666 (N_13666,N_10500,N_9539);
nor U13667 (N_13667,N_8925,N_8059);
nor U13668 (N_13668,N_8721,N_11820);
nor U13669 (N_13669,N_8401,N_8119);
or U13670 (N_13670,N_9918,N_9533);
and U13671 (N_13671,N_10468,N_11741);
nand U13672 (N_13672,N_8670,N_10163);
nand U13673 (N_13673,N_8990,N_8520);
nand U13674 (N_13674,N_8960,N_9417);
nor U13675 (N_13675,N_10515,N_8066);
nand U13676 (N_13676,N_11107,N_11035);
or U13677 (N_13677,N_9245,N_8631);
and U13678 (N_13678,N_11623,N_8369);
nand U13679 (N_13679,N_8477,N_11203);
nand U13680 (N_13680,N_10459,N_9816);
and U13681 (N_13681,N_9427,N_10856);
nor U13682 (N_13682,N_9523,N_10043);
nand U13683 (N_13683,N_11002,N_11148);
nor U13684 (N_13684,N_11695,N_9317);
or U13685 (N_13685,N_11520,N_10642);
nor U13686 (N_13686,N_9744,N_9683);
or U13687 (N_13687,N_10034,N_8560);
or U13688 (N_13688,N_10240,N_8841);
nand U13689 (N_13689,N_10840,N_9621);
and U13690 (N_13690,N_9380,N_8050);
and U13691 (N_13691,N_9332,N_10207);
nor U13692 (N_13692,N_8541,N_9753);
or U13693 (N_13693,N_8445,N_8073);
nand U13694 (N_13694,N_10674,N_10133);
nor U13695 (N_13695,N_9107,N_9442);
or U13696 (N_13696,N_10504,N_11645);
nor U13697 (N_13697,N_9194,N_10525);
nand U13698 (N_13698,N_9527,N_10115);
nand U13699 (N_13699,N_8284,N_11811);
nor U13700 (N_13700,N_9644,N_8312);
nor U13701 (N_13701,N_11300,N_10299);
or U13702 (N_13702,N_8167,N_11344);
and U13703 (N_13703,N_8784,N_10183);
nor U13704 (N_13704,N_8465,N_11759);
or U13705 (N_13705,N_9978,N_10956);
and U13706 (N_13706,N_11016,N_9090);
nand U13707 (N_13707,N_10682,N_9299);
or U13708 (N_13708,N_9247,N_10502);
and U13709 (N_13709,N_11380,N_10129);
nor U13710 (N_13710,N_8137,N_10781);
nand U13711 (N_13711,N_9688,N_11005);
nor U13712 (N_13712,N_9601,N_10022);
nand U13713 (N_13713,N_9981,N_8946);
nand U13714 (N_13714,N_9456,N_9971);
nand U13715 (N_13715,N_10432,N_9043);
nor U13716 (N_13716,N_9534,N_10884);
or U13717 (N_13717,N_10237,N_9369);
nor U13718 (N_13718,N_10727,N_11415);
and U13719 (N_13719,N_9355,N_10044);
or U13720 (N_13720,N_9881,N_9123);
nor U13721 (N_13721,N_8547,N_8208);
or U13722 (N_13722,N_11656,N_8699);
nor U13723 (N_13723,N_11248,N_11193);
nor U13724 (N_13724,N_9221,N_10363);
nand U13725 (N_13725,N_10016,N_10606);
or U13726 (N_13726,N_10976,N_11120);
or U13727 (N_13727,N_8773,N_8696);
nand U13728 (N_13728,N_10808,N_10626);
and U13729 (N_13729,N_10565,N_10635);
and U13730 (N_13730,N_8893,N_8399);
nand U13731 (N_13731,N_11145,N_10875);
nor U13732 (N_13732,N_10139,N_9668);
or U13733 (N_13733,N_11259,N_11727);
nor U13734 (N_13734,N_11038,N_10037);
nor U13735 (N_13735,N_8274,N_9162);
and U13736 (N_13736,N_10867,N_10509);
nand U13737 (N_13737,N_8530,N_10489);
or U13738 (N_13738,N_8061,N_11707);
nor U13739 (N_13739,N_11006,N_9267);
xor U13740 (N_13740,N_9536,N_8124);
nand U13741 (N_13741,N_10294,N_11817);
or U13742 (N_13742,N_9775,N_8156);
and U13743 (N_13743,N_8308,N_8287);
or U13744 (N_13744,N_10625,N_11293);
or U13745 (N_13745,N_11106,N_8710);
nor U13746 (N_13746,N_10348,N_8873);
nand U13747 (N_13747,N_9144,N_10807);
and U13748 (N_13748,N_10990,N_10262);
nand U13749 (N_13749,N_10846,N_9743);
and U13750 (N_13750,N_11979,N_10637);
or U13751 (N_13751,N_11330,N_9292);
and U13752 (N_13752,N_10708,N_10386);
nor U13753 (N_13753,N_9217,N_11716);
nor U13754 (N_13754,N_8964,N_11000);
and U13755 (N_13755,N_10940,N_8053);
nand U13756 (N_13756,N_9036,N_11671);
nor U13757 (N_13757,N_11779,N_11742);
and U13758 (N_13758,N_10209,N_11033);
or U13759 (N_13759,N_11385,N_8967);
nor U13760 (N_13760,N_9437,N_11289);
nor U13761 (N_13761,N_11453,N_10656);
or U13762 (N_13762,N_10211,N_8318);
and U13763 (N_13763,N_11595,N_10213);
and U13764 (N_13764,N_9345,N_11906);
or U13765 (N_13765,N_10255,N_8367);
and U13766 (N_13766,N_9746,N_10192);
and U13767 (N_13767,N_11087,N_9884);
and U13768 (N_13768,N_9200,N_11188);
nor U13769 (N_13769,N_11388,N_10534);
nor U13770 (N_13770,N_11605,N_9890);
nor U13771 (N_13771,N_10536,N_10141);
and U13772 (N_13772,N_8095,N_9984);
nor U13773 (N_13773,N_11180,N_11522);
or U13774 (N_13774,N_8394,N_10831);
nand U13775 (N_13775,N_8023,N_10966);
nand U13776 (N_13776,N_9578,N_10570);
or U13777 (N_13777,N_8285,N_9045);
nor U13778 (N_13778,N_11229,N_8192);
and U13779 (N_13779,N_11894,N_9008);
nor U13780 (N_13780,N_8047,N_10615);
and U13781 (N_13781,N_8056,N_9805);
nand U13782 (N_13782,N_11925,N_11298);
nand U13783 (N_13783,N_10910,N_10402);
and U13784 (N_13784,N_9485,N_11350);
and U13785 (N_13785,N_10789,N_9339);
and U13786 (N_13786,N_9707,N_10098);
and U13787 (N_13787,N_11691,N_9353);
nand U13788 (N_13788,N_8790,N_9871);
and U13789 (N_13789,N_11381,N_9446);
and U13790 (N_13790,N_10066,N_11869);
nor U13791 (N_13791,N_10408,N_9281);
nor U13792 (N_13792,N_8184,N_8805);
nand U13793 (N_13793,N_11712,N_10519);
and U13794 (N_13794,N_10228,N_9184);
nand U13795 (N_13795,N_8146,N_8676);
nor U13796 (N_13796,N_8978,N_10216);
nor U13797 (N_13797,N_10728,N_10268);
nand U13798 (N_13798,N_11654,N_10981);
or U13799 (N_13799,N_10317,N_10961);
and U13800 (N_13800,N_8320,N_11034);
nand U13801 (N_13801,N_8322,N_8298);
and U13802 (N_13802,N_11839,N_8666);
and U13803 (N_13803,N_10788,N_9679);
nand U13804 (N_13804,N_9580,N_9637);
nand U13805 (N_13805,N_8820,N_10365);
nand U13806 (N_13806,N_8022,N_11377);
nor U13807 (N_13807,N_11557,N_10179);
xor U13808 (N_13808,N_8502,N_11633);
or U13809 (N_13809,N_9961,N_8546);
nand U13810 (N_13810,N_11554,N_10528);
or U13811 (N_13811,N_10203,N_9309);
nor U13812 (N_13812,N_9498,N_9840);
or U13813 (N_13813,N_9930,N_11101);
or U13814 (N_13814,N_11233,N_9103);
nor U13815 (N_13815,N_8307,N_9702);
xnor U13816 (N_13816,N_10779,N_11683);
nand U13817 (N_13817,N_10059,N_8839);
nand U13818 (N_13818,N_8254,N_9230);
nand U13819 (N_13819,N_9591,N_11763);
and U13820 (N_13820,N_8891,N_9757);
nand U13821 (N_13821,N_9050,N_9254);
or U13822 (N_13822,N_9253,N_8159);
and U13823 (N_13823,N_11310,N_9921);
or U13824 (N_13824,N_8795,N_11860);
or U13825 (N_13825,N_9375,N_11082);
and U13826 (N_13826,N_11392,N_8587);
and U13827 (N_13827,N_10843,N_8088);
nor U13828 (N_13828,N_10905,N_9639);
or U13829 (N_13829,N_10612,N_10360);
or U13830 (N_13830,N_9407,N_11899);
nand U13831 (N_13831,N_11909,N_9186);
nand U13832 (N_13832,N_9091,N_8470);
and U13833 (N_13833,N_9600,N_8344);
and U13834 (N_13834,N_9843,N_11277);
nor U13835 (N_13835,N_10513,N_11133);
nand U13836 (N_13836,N_11055,N_9363);
nor U13837 (N_13837,N_10977,N_11813);
nand U13838 (N_13838,N_11384,N_11165);
xnor U13839 (N_13839,N_11168,N_11995);
or U13840 (N_13840,N_11413,N_9063);
nand U13841 (N_13841,N_8993,N_9958);
nand U13842 (N_13842,N_11610,N_9736);
or U13843 (N_13843,N_10573,N_9432);
nor U13844 (N_13844,N_11314,N_9252);
nand U13845 (N_13845,N_10033,N_9526);
nand U13846 (N_13846,N_8592,N_10845);
nand U13847 (N_13847,N_11067,N_9095);
nor U13848 (N_13848,N_10558,N_9838);
nor U13849 (N_13849,N_8115,N_9286);
or U13850 (N_13850,N_11356,N_8404);
and U13851 (N_13851,N_8656,N_10351);
nor U13852 (N_13852,N_8420,N_10126);
or U13853 (N_13853,N_8223,N_8090);
and U13854 (N_13854,N_8532,N_11470);
and U13855 (N_13855,N_11532,N_9028);
nor U13856 (N_13856,N_11449,N_11829);
and U13857 (N_13857,N_9075,N_10657);
nor U13858 (N_13858,N_8854,N_11911);
and U13859 (N_13859,N_9142,N_10998);
nor U13860 (N_13860,N_9593,N_11410);
or U13861 (N_13861,N_11366,N_8488);
or U13862 (N_13862,N_8662,N_9116);
nand U13863 (N_13863,N_8608,N_10005);
and U13864 (N_13864,N_8251,N_11959);
and U13865 (N_13865,N_11209,N_8152);
and U13866 (N_13866,N_10968,N_10227);
nor U13867 (N_13867,N_8944,N_8169);
or U13868 (N_13868,N_11253,N_9300);
and U13869 (N_13869,N_8519,N_9822);
nor U13870 (N_13870,N_11196,N_9804);
nor U13871 (N_13871,N_9180,N_11461);
and U13872 (N_13872,N_10813,N_10086);
and U13873 (N_13873,N_8395,N_9970);
nand U13874 (N_13874,N_8558,N_9120);
nand U13875 (N_13875,N_11365,N_10160);
nand U13876 (N_13876,N_11638,N_8102);
and U13877 (N_13877,N_11649,N_8173);
nor U13878 (N_13878,N_9124,N_9766);
and U13879 (N_13879,N_10835,N_10646);
and U13880 (N_13880,N_8613,N_9719);
nor U13881 (N_13881,N_9113,N_10448);
nor U13882 (N_13882,N_11305,N_9266);
and U13883 (N_13883,N_8753,N_8768);
or U13884 (N_13884,N_11371,N_8118);
or U13885 (N_13885,N_8068,N_9557);
and U13886 (N_13886,N_8209,N_8064);
nand U13887 (N_13887,N_11967,N_9548);
nor U13888 (N_13888,N_9740,N_8573);
or U13889 (N_13889,N_11672,N_11260);
and U13890 (N_13890,N_11858,N_11003);
nor U13891 (N_13891,N_8319,N_10762);
or U13892 (N_13892,N_10336,N_10276);
or U13893 (N_13893,N_10434,N_10731);
nor U13894 (N_13894,N_10440,N_9863);
and U13895 (N_13895,N_10321,N_11024);
nor U13896 (N_13896,N_10540,N_11510);
nor U13897 (N_13897,N_10138,N_9488);
nand U13898 (N_13898,N_11866,N_10687);
and U13899 (N_13899,N_11596,N_11011);
nor U13900 (N_13900,N_10670,N_10980);
nand U13901 (N_13901,N_8200,N_11014);
and U13902 (N_13902,N_11127,N_10451);
nor U13903 (N_13903,N_9846,N_9607);
nor U13904 (N_13904,N_10008,N_9993);
or U13905 (N_13905,N_11167,N_8889);
or U13906 (N_13906,N_8105,N_9156);
nand U13907 (N_13907,N_9959,N_9078);
nor U13908 (N_13908,N_11831,N_11353);
xnor U13909 (N_13909,N_9850,N_8667);
and U13910 (N_13910,N_10641,N_10667);
and U13911 (N_13911,N_8290,N_11500);
nor U13912 (N_13912,N_9199,N_9460);
nand U13913 (N_13913,N_11264,N_9543);
nand U13914 (N_13914,N_11075,N_10148);
nand U13915 (N_13915,N_11164,N_11861);
nand U13916 (N_13916,N_9068,N_8607);
nor U13917 (N_13917,N_11503,N_8777);
nor U13918 (N_13918,N_9451,N_8454);
or U13919 (N_13919,N_11393,N_8905);
nand U13920 (N_13920,N_8740,N_11466);
and U13921 (N_13921,N_10368,N_9955);
and U13922 (N_13922,N_11018,N_11455);
or U13923 (N_13923,N_8760,N_11243);
nor U13924 (N_13924,N_10830,N_11234);
nand U13925 (N_13925,N_10780,N_8814);
xnor U13926 (N_13926,N_10638,N_9779);
or U13927 (N_13927,N_11110,N_8482);
nor U13928 (N_13928,N_10092,N_8009);
nor U13929 (N_13929,N_9444,N_10206);
nand U13930 (N_13930,N_9511,N_10170);
nor U13931 (N_13931,N_11973,N_11570);
or U13932 (N_13932,N_11232,N_8808);
and U13933 (N_13933,N_11156,N_9240);
or U13934 (N_13934,N_10858,N_11629);
and U13935 (N_13935,N_8858,N_8628);
and U13936 (N_13936,N_11778,N_8101);
and U13937 (N_13937,N_11479,N_8634);
and U13938 (N_13938,N_9259,N_8434);
or U13939 (N_13939,N_11426,N_11189);
nor U13940 (N_13940,N_11197,N_11401);
and U13941 (N_13941,N_9948,N_9646);
and U13942 (N_13942,N_8302,N_10930);
nor U13943 (N_13943,N_10215,N_8745);
nand U13944 (N_13944,N_9093,N_9019);
nor U13945 (N_13945,N_10857,N_9875);
nor U13946 (N_13946,N_9700,N_8034);
nand U13947 (N_13947,N_8279,N_10873);
nor U13948 (N_13948,N_11555,N_10377);
and U13949 (N_13949,N_11199,N_8496);
and U13950 (N_13950,N_11047,N_10147);
or U13951 (N_13951,N_10733,N_10128);
and U13952 (N_13952,N_11852,N_10156);
nor U13953 (N_13953,N_11927,N_11578);
and U13954 (N_13954,N_8207,N_9998);
nand U13955 (N_13955,N_8321,N_10585);
or U13956 (N_13956,N_8671,N_11123);
nor U13957 (N_13957,N_11976,N_11889);
or U13958 (N_13958,N_11235,N_9249);
and U13959 (N_13959,N_8812,N_11292);
nand U13960 (N_13960,N_11325,N_9289);
or U13961 (N_13961,N_8172,N_8122);
or U13962 (N_13962,N_10523,N_11176);
and U13963 (N_13963,N_11266,N_11493);
and U13964 (N_13964,N_8164,N_11135);
nand U13965 (N_13965,N_8168,N_9855);
nor U13966 (N_13966,N_10248,N_10838);
and U13967 (N_13967,N_8885,N_8155);
or U13968 (N_13968,N_10849,N_9449);
nand U13969 (N_13969,N_8074,N_10189);
and U13970 (N_13970,N_9760,N_8728);
and U13971 (N_13971,N_9340,N_11099);
nand U13972 (N_13972,N_10784,N_9391);
or U13973 (N_13973,N_9603,N_11368);
and U13974 (N_13974,N_11245,N_11827);
and U13975 (N_13975,N_9680,N_10629);
nand U13976 (N_13976,N_9546,N_10984);
nor U13977 (N_13977,N_9817,N_9605);
nor U13978 (N_13978,N_10920,N_10964);
and U13979 (N_13979,N_11731,N_11104);
or U13980 (N_13980,N_8853,N_10347);
and U13981 (N_13981,N_10135,N_8703);
nor U13982 (N_13982,N_10690,N_9691);
nor U13983 (N_13983,N_9754,N_10810);
nor U13984 (N_13984,N_10077,N_11042);
and U13985 (N_13985,N_8421,N_11613);
or U13986 (N_13986,N_9256,N_11576);
nand U13987 (N_13987,N_9865,N_8018);
or U13988 (N_13988,N_8492,N_9265);
nor U13989 (N_13989,N_8075,N_9710);
nand U13990 (N_13990,N_9941,N_8425);
or U13991 (N_13991,N_10658,N_9730);
nand U13992 (N_13992,N_9202,N_8025);
nor U13993 (N_13993,N_8830,N_11824);
nand U13994 (N_13994,N_8708,N_9458);
and U13995 (N_13995,N_8311,N_11132);
nor U13996 (N_13996,N_8072,N_11971);
or U13997 (N_13997,N_10230,N_10257);
nand U13998 (N_13998,N_8648,N_10714);
or U13999 (N_13999,N_9625,N_8963);
nand U14000 (N_14000,N_11617,N_8489);
nand U14001 (N_14001,N_11076,N_11035);
nand U14002 (N_14002,N_9191,N_11602);
and U14003 (N_14003,N_10434,N_9995);
and U14004 (N_14004,N_11905,N_10617);
and U14005 (N_14005,N_8948,N_10226);
nand U14006 (N_14006,N_9197,N_9420);
or U14007 (N_14007,N_11378,N_8642);
nor U14008 (N_14008,N_11518,N_9627);
or U14009 (N_14009,N_8704,N_10828);
and U14010 (N_14010,N_10810,N_10163);
nand U14011 (N_14011,N_11505,N_10218);
nand U14012 (N_14012,N_9369,N_9585);
and U14013 (N_14013,N_11519,N_8763);
nor U14014 (N_14014,N_9156,N_10527);
nor U14015 (N_14015,N_9591,N_8463);
and U14016 (N_14016,N_9418,N_10352);
and U14017 (N_14017,N_10769,N_9417);
nor U14018 (N_14018,N_8600,N_9525);
nand U14019 (N_14019,N_11582,N_8608);
nand U14020 (N_14020,N_9279,N_9121);
nor U14021 (N_14021,N_10359,N_10159);
and U14022 (N_14022,N_8435,N_8859);
nor U14023 (N_14023,N_10437,N_10009);
nor U14024 (N_14024,N_10240,N_8390);
nand U14025 (N_14025,N_11648,N_9698);
nand U14026 (N_14026,N_8761,N_11167);
and U14027 (N_14027,N_8275,N_9835);
and U14028 (N_14028,N_10520,N_8269);
or U14029 (N_14029,N_9677,N_10055);
nor U14030 (N_14030,N_8501,N_10763);
nand U14031 (N_14031,N_9041,N_11218);
and U14032 (N_14032,N_11412,N_9803);
or U14033 (N_14033,N_11317,N_9468);
or U14034 (N_14034,N_9699,N_11810);
and U14035 (N_14035,N_8053,N_11867);
or U14036 (N_14036,N_8035,N_10887);
and U14037 (N_14037,N_8833,N_8497);
and U14038 (N_14038,N_11482,N_9489);
and U14039 (N_14039,N_8723,N_8507);
or U14040 (N_14040,N_10881,N_9145);
nand U14041 (N_14041,N_9335,N_8493);
nor U14042 (N_14042,N_8386,N_8502);
and U14043 (N_14043,N_8312,N_8372);
nand U14044 (N_14044,N_8044,N_11631);
and U14045 (N_14045,N_8083,N_8507);
nor U14046 (N_14046,N_9734,N_10485);
and U14047 (N_14047,N_11582,N_8077);
and U14048 (N_14048,N_9535,N_8046);
nor U14049 (N_14049,N_10880,N_8488);
and U14050 (N_14050,N_8571,N_8591);
and U14051 (N_14051,N_11458,N_10997);
nor U14052 (N_14052,N_10336,N_8487);
and U14053 (N_14053,N_11421,N_11115);
or U14054 (N_14054,N_9855,N_11006);
or U14055 (N_14055,N_11100,N_10475);
and U14056 (N_14056,N_10614,N_8608);
or U14057 (N_14057,N_11411,N_10749);
or U14058 (N_14058,N_8472,N_11876);
and U14059 (N_14059,N_10055,N_8602);
nand U14060 (N_14060,N_8391,N_11484);
or U14061 (N_14061,N_11044,N_11845);
and U14062 (N_14062,N_10433,N_8720);
and U14063 (N_14063,N_11862,N_8249);
and U14064 (N_14064,N_11371,N_9810);
nor U14065 (N_14065,N_9103,N_10115);
or U14066 (N_14066,N_9688,N_9105);
nor U14067 (N_14067,N_9875,N_10214);
nor U14068 (N_14068,N_8018,N_10079);
and U14069 (N_14069,N_10455,N_9773);
or U14070 (N_14070,N_11934,N_10033);
or U14071 (N_14071,N_8564,N_10373);
nand U14072 (N_14072,N_9355,N_10360);
nor U14073 (N_14073,N_9282,N_9080);
nor U14074 (N_14074,N_8628,N_9679);
and U14075 (N_14075,N_11533,N_11241);
nand U14076 (N_14076,N_8340,N_11554);
nor U14077 (N_14077,N_10335,N_8895);
or U14078 (N_14078,N_8190,N_10929);
and U14079 (N_14079,N_9937,N_10132);
or U14080 (N_14080,N_11654,N_9969);
or U14081 (N_14081,N_9677,N_8174);
and U14082 (N_14082,N_8186,N_8607);
nand U14083 (N_14083,N_11152,N_10952);
nand U14084 (N_14084,N_11118,N_10853);
nand U14085 (N_14085,N_8592,N_8363);
or U14086 (N_14086,N_11972,N_10642);
nand U14087 (N_14087,N_10779,N_11365);
and U14088 (N_14088,N_9135,N_11683);
nor U14089 (N_14089,N_8415,N_9494);
and U14090 (N_14090,N_9860,N_11030);
or U14091 (N_14091,N_11115,N_8352);
and U14092 (N_14092,N_9816,N_10594);
or U14093 (N_14093,N_9696,N_9992);
or U14094 (N_14094,N_9842,N_10494);
nor U14095 (N_14095,N_11133,N_11695);
nor U14096 (N_14096,N_10609,N_11221);
nor U14097 (N_14097,N_9966,N_10548);
or U14098 (N_14098,N_9132,N_9494);
nand U14099 (N_14099,N_10451,N_10858);
nand U14100 (N_14100,N_10303,N_8875);
and U14101 (N_14101,N_8837,N_9415);
nand U14102 (N_14102,N_10049,N_9249);
and U14103 (N_14103,N_9297,N_9171);
and U14104 (N_14104,N_11901,N_10602);
nand U14105 (N_14105,N_11087,N_10555);
or U14106 (N_14106,N_9067,N_10508);
nand U14107 (N_14107,N_10563,N_11169);
or U14108 (N_14108,N_10888,N_10644);
nand U14109 (N_14109,N_11711,N_11335);
nor U14110 (N_14110,N_8362,N_11833);
nand U14111 (N_14111,N_8363,N_9713);
nor U14112 (N_14112,N_9784,N_10873);
nor U14113 (N_14113,N_11019,N_10016);
or U14114 (N_14114,N_10717,N_9657);
nand U14115 (N_14115,N_11401,N_10578);
nand U14116 (N_14116,N_11751,N_9075);
or U14117 (N_14117,N_10238,N_11851);
nor U14118 (N_14118,N_8671,N_11132);
nand U14119 (N_14119,N_11265,N_11175);
or U14120 (N_14120,N_9811,N_10522);
or U14121 (N_14121,N_9258,N_8678);
nor U14122 (N_14122,N_8589,N_11868);
and U14123 (N_14123,N_11707,N_11192);
nor U14124 (N_14124,N_9591,N_11889);
nand U14125 (N_14125,N_8443,N_10567);
or U14126 (N_14126,N_10464,N_8126);
nor U14127 (N_14127,N_10493,N_8048);
nand U14128 (N_14128,N_11210,N_11931);
nand U14129 (N_14129,N_10425,N_10349);
nor U14130 (N_14130,N_11106,N_10420);
and U14131 (N_14131,N_8450,N_11604);
and U14132 (N_14132,N_11311,N_11780);
or U14133 (N_14133,N_8733,N_8159);
and U14134 (N_14134,N_11738,N_9896);
nor U14135 (N_14135,N_10632,N_11386);
or U14136 (N_14136,N_8544,N_8877);
nand U14137 (N_14137,N_9013,N_11513);
nand U14138 (N_14138,N_11444,N_9908);
and U14139 (N_14139,N_11944,N_11085);
and U14140 (N_14140,N_9607,N_11104);
nor U14141 (N_14141,N_8138,N_9022);
or U14142 (N_14142,N_9087,N_11569);
or U14143 (N_14143,N_11188,N_9215);
and U14144 (N_14144,N_11605,N_10148);
nand U14145 (N_14145,N_11484,N_10532);
or U14146 (N_14146,N_11965,N_9819);
nor U14147 (N_14147,N_10954,N_11491);
and U14148 (N_14148,N_10770,N_11676);
or U14149 (N_14149,N_9603,N_11003);
or U14150 (N_14150,N_11994,N_11728);
and U14151 (N_14151,N_9415,N_9417);
and U14152 (N_14152,N_11085,N_8640);
or U14153 (N_14153,N_10675,N_10945);
or U14154 (N_14154,N_11544,N_10723);
nor U14155 (N_14155,N_10304,N_8568);
nor U14156 (N_14156,N_10595,N_9241);
or U14157 (N_14157,N_8962,N_8036);
or U14158 (N_14158,N_11779,N_8242);
nor U14159 (N_14159,N_10770,N_10047);
nand U14160 (N_14160,N_11173,N_9767);
nor U14161 (N_14161,N_10842,N_9739);
nor U14162 (N_14162,N_10670,N_11256);
nand U14163 (N_14163,N_9455,N_10409);
or U14164 (N_14164,N_9028,N_9108);
or U14165 (N_14165,N_11020,N_10359);
nand U14166 (N_14166,N_9297,N_10063);
nor U14167 (N_14167,N_8325,N_8721);
or U14168 (N_14168,N_9866,N_9629);
and U14169 (N_14169,N_9218,N_9664);
and U14170 (N_14170,N_8851,N_10611);
and U14171 (N_14171,N_8511,N_8522);
and U14172 (N_14172,N_9137,N_9376);
nor U14173 (N_14173,N_8546,N_10583);
nor U14174 (N_14174,N_9628,N_9520);
or U14175 (N_14175,N_10632,N_9443);
and U14176 (N_14176,N_8030,N_10881);
or U14177 (N_14177,N_9127,N_10584);
and U14178 (N_14178,N_11919,N_8004);
nor U14179 (N_14179,N_11511,N_8089);
nor U14180 (N_14180,N_8257,N_9868);
nand U14181 (N_14181,N_8260,N_8099);
nand U14182 (N_14182,N_9594,N_8188);
or U14183 (N_14183,N_11716,N_8086);
and U14184 (N_14184,N_8696,N_9340);
nand U14185 (N_14185,N_11075,N_11088);
nand U14186 (N_14186,N_11976,N_11481);
nor U14187 (N_14187,N_11837,N_9476);
and U14188 (N_14188,N_9450,N_11889);
or U14189 (N_14189,N_9860,N_10898);
nor U14190 (N_14190,N_11411,N_11248);
or U14191 (N_14191,N_10294,N_11271);
or U14192 (N_14192,N_10603,N_10262);
nand U14193 (N_14193,N_8836,N_10558);
nor U14194 (N_14194,N_11371,N_11877);
or U14195 (N_14195,N_9678,N_8900);
or U14196 (N_14196,N_9679,N_10982);
and U14197 (N_14197,N_10484,N_10535);
or U14198 (N_14198,N_8595,N_11223);
or U14199 (N_14199,N_11669,N_9396);
nor U14200 (N_14200,N_10807,N_8273);
nor U14201 (N_14201,N_11337,N_11094);
nor U14202 (N_14202,N_9051,N_9726);
nand U14203 (N_14203,N_10133,N_9042);
nor U14204 (N_14204,N_11577,N_10696);
nor U14205 (N_14205,N_9057,N_9001);
nand U14206 (N_14206,N_11212,N_10028);
nor U14207 (N_14207,N_11619,N_10661);
nor U14208 (N_14208,N_9783,N_11517);
and U14209 (N_14209,N_10282,N_10483);
nor U14210 (N_14210,N_9030,N_10985);
or U14211 (N_14211,N_8849,N_9953);
nand U14212 (N_14212,N_9113,N_11395);
nand U14213 (N_14213,N_8613,N_9833);
and U14214 (N_14214,N_10773,N_10284);
or U14215 (N_14215,N_10266,N_11757);
or U14216 (N_14216,N_8417,N_11116);
nand U14217 (N_14217,N_8386,N_10561);
nand U14218 (N_14218,N_10185,N_9758);
or U14219 (N_14219,N_10326,N_11580);
and U14220 (N_14220,N_9966,N_11522);
nand U14221 (N_14221,N_10874,N_11257);
or U14222 (N_14222,N_8797,N_9269);
and U14223 (N_14223,N_9854,N_8426);
nor U14224 (N_14224,N_9321,N_10350);
or U14225 (N_14225,N_8615,N_10927);
and U14226 (N_14226,N_9393,N_8467);
nand U14227 (N_14227,N_8971,N_11296);
nor U14228 (N_14228,N_11966,N_10373);
or U14229 (N_14229,N_10447,N_10337);
nand U14230 (N_14230,N_10464,N_9886);
nor U14231 (N_14231,N_11495,N_9754);
and U14232 (N_14232,N_10723,N_9544);
and U14233 (N_14233,N_8336,N_9755);
and U14234 (N_14234,N_10077,N_8272);
or U14235 (N_14235,N_9053,N_8332);
nand U14236 (N_14236,N_9464,N_10994);
or U14237 (N_14237,N_9239,N_8894);
or U14238 (N_14238,N_8452,N_9282);
and U14239 (N_14239,N_10483,N_8840);
or U14240 (N_14240,N_9170,N_8924);
nand U14241 (N_14241,N_10683,N_11263);
or U14242 (N_14242,N_8017,N_10555);
nand U14243 (N_14243,N_9677,N_8501);
nand U14244 (N_14244,N_9947,N_9007);
nor U14245 (N_14245,N_8006,N_11324);
and U14246 (N_14246,N_9924,N_10671);
or U14247 (N_14247,N_10738,N_11797);
nand U14248 (N_14248,N_11337,N_10004);
nand U14249 (N_14249,N_8793,N_8152);
nand U14250 (N_14250,N_10279,N_9179);
nor U14251 (N_14251,N_8528,N_9694);
or U14252 (N_14252,N_10321,N_11845);
and U14253 (N_14253,N_9087,N_9640);
or U14254 (N_14254,N_8522,N_9903);
and U14255 (N_14255,N_10865,N_10871);
nand U14256 (N_14256,N_8897,N_10040);
nor U14257 (N_14257,N_8798,N_11597);
or U14258 (N_14258,N_11027,N_9915);
nand U14259 (N_14259,N_8447,N_11041);
and U14260 (N_14260,N_8296,N_11518);
nand U14261 (N_14261,N_9661,N_11032);
xnor U14262 (N_14262,N_8481,N_11020);
or U14263 (N_14263,N_10478,N_8315);
and U14264 (N_14264,N_8671,N_8465);
or U14265 (N_14265,N_10539,N_11047);
nor U14266 (N_14266,N_8963,N_11663);
nor U14267 (N_14267,N_11011,N_8341);
or U14268 (N_14268,N_10278,N_9681);
or U14269 (N_14269,N_10661,N_11494);
nand U14270 (N_14270,N_9160,N_10713);
or U14271 (N_14271,N_11709,N_8529);
nand U14272 (N_14272,N_10200,N_8704);
nand U14273 (N_14273,N_10759,N_11454);
nor U14274 (N_14274,N_10584,N_10550);
nand U14275 (N_14275,N_10882,N_8914);
or U14276 (N_14276,N_10920,N_10701);
or U14277 (N_14277,N_10597,N_11284);
and U14278 (N_14278,N_9770,N_10332);
or U14279 (N_14279,N_10444,N_8141);
nor U14280 (N_14280,N_9755,N_9720);
nand U14281 (N_14281,N_8276,N_11478);
nor U14282 (N_14282,N_11868,N_8910);
nor U14283 (N_14283,N_10498,N_9748);
nor U14284 (N_14284,N_10651,N_10266);
and U14285 (N_14285,N_9125,N_11491);
nor U14286 (N_14286,N_8373,N_11828);
nand U14287 (N_14287,N_9220,N_8245);
and U14288 (N_14288,N_8629,N_8214);
nand U14289 (N_14289,N_10425,N_10377);
or U14290 (N_14290,N_10285,N_10592);
or U14291 (N_14291,N_9757,N_10267);
nor U14292 (N_14292,N_11103,N_9908);
nand U14293 (N_14293,N_11558,N_9061);
nor U14294 (N_14294,N_11108,N_8087);
and U14295 (N_14295,N_10036,N_11315);
nand U14296 (N_14296,N_11934,N_8587);
and U14297 (N_14297,N_9761,N_10612);
or U14298 (N_14298,N_11564,N_11255);
and U14299 (N_14299,N_8877,N_9990);
nor U14300 (N_14300,N_10087,N_11669);
nor U14301 (N_14301,N_9002,N_10699);
and U14302 (N_14302,N_11275,N_11076);
nor U14303 (N_14303,N_10815,N_11296);
nor U14304 (N_14304,N_9377,N_8116);
nor U14305 (N_14305,N_11193,N_8291);
or U14306 (N_14306,N_8106,N_8834);
nor U14307 (N_14307,N_8428,N_9850);
or U14308 (N_14308,N_9599,N_11537);
or U14309 (N_14309,N_8147,N_10347);
or U14310 (N_14310,N_11046,N_9210);
nand U14311 (N_14311,N_9528,N_10071);
and U14312 (N_14312,N_10302,N_10726);
and U14313 (N_14313,N_10384,N_11564);
or U14314 (N_14314,N_8510,N_10955);
or U14315 (N_14315,N_9073,N_8111);
nand U14316 (N_14316,N_9439,N_10077);
nor U14317 (N_14317,N_11550,N_10093);
nand U14318 (N_14318,N_11170,N_9804);
nor U14319 (N_14319,N_11464,N_10501);
or U14320 (N_14320,N_9002,N_11135);
or U14321 (N_14321,N_8646,N_8490);
nor U14322 (N_14322,N_9858,N_9328);
or U14323 (N_14323,N_11208,N_11751);
or U14324 (N_14324,N_11527,N_10234);
and U14325 (N_14325,N_8423,N_9410);
and U14326 (N_14326,N_9714,N_10821);
or U14327 (N_14327,N_9246,N_10474);
and U14328 (N_14328,N_9681,N_9293);
or U14329 (N_14329,N_10886,N_10090);
and U14330 (N_14330,N_8164,N_11077);
nor U14331 (N_14331,N_9588,N_8059);
nand U14332 (N_14332,N_8993,N_10409);
nor U14333 (N_14333,N_8712,N_11700);
or U14334 (N_14334,N_8472,N_11947);
or U14335 (N_14335,N_10317,N_9795);
and U14336 (N_14336,N_8350,N_10213);
and U14337 (N_14337,N_8078,N_8311);
and U14338 (N_14338,N_10726,N_11661);
nand U14339 (N_14339,N_10582,N_10999);
or U14340 (N_14340,N_11983,N_9491);
nor U14341 (N_14341,N_8971,N_9098);
xor U14342 (N_14342,N_11654,N_10984);
nand U14343 (N_14343,N_8084,N_11543);
or U14344 (N_14344,N_11349,N_11138);
and U14345 (N_14345,N_11773,N_10181);
or U14346 (N_14346,N_9084,N_9509);
or U14347 (N_14347,N_9303,N_10780);
nand U14348 (N_14348,N_8643,N_9751);
and U14349 (N_14349,N_11088,N_10801);
or U14350 (N_14350,N_11227,N_9363);
and U14351 (N_14351,N_11995,N_9326);
nand U14352 (N_14352,N_11946,N_9379);
and U14353 (N_14353,N_10355,N_11435);
and U14354 (N_14354,N_11105,N_9790);
and U14355 (N_14355,N_8171,N_8112);
or U14356 (N_14356,N_8851,N_10896);
nand U14357 (N_14357,N_11641,N_10566);
nand U14358 (N_14358,N_9676,N_9759);
and U14359 (N_14359,N_11904,N_11484);
nand U14360 (N_14360,N_10148,N_11035);
nor U14361 (N_14361,N_10303,N_9291);
and U14362 (N_14362,N_8499,N_9212);
nor U14363 (N_14363,N_10848,N_8336);
or U14364 (N_14364,N_9640,N_11090);
or U14365 (N_14365,N_10793,N_8556);
and U14366 (N_14366,N_8174,N_11277);
and U14367 (N_14367,N_11218,N_11144);
nor U14368 (N_14368,N_9585,N_11519);
nand U14369 (N_14369,N_10892,N_10736);
nor U14370 (N_14370,N_10023,N_8785);
nand U14371 (N_14371,N_11051,N_11309);
nor U14372 (N_14372,N_9987,N_8107);
nor U14373 (N_14373,N_11437,N_9967);
nor U14374 (N_14374,N_9893,N_11374);
nand U14375 (N_14375,N_9255,N_8294);
and U14376 (N_14376,N_8190,N_10106);
and U14377 (N_14377,N_10273,N_9652);
nor U14378 (N_14378,N_8412,N_10986);
or U14379 (N_14379,N_10093,N_8148);
nor U14380 (N_14380,N_11508,N_9368);
and U14381 (N_14381,N_10101,N_8988);
nor U14382 (N_14382,N_11708,N_10565);
nand U14383 (N_14383,N_11383,N_11253);
nor U14384 (N_14384,N_8528,N_11569);
or U14385 (N_14385,N_8727,N_10172);
or U14386 (N_14386,N_9770,N_9010);
nor U14387 (N_14387,N_11216,N_9313);
nor U14388 (N_14388,N_10035,N_9411);
nand U14389 (N_14389,N_8710,N_9860);
nand U14390 (N_14390,N_11281,N_8137);
nand U14391 (N_14391,N_9912,N_11574);
or U14392 (N_14392,N_9430,N_11507);
nand U14393 (N_14393,N_10875,N_8979);
nor U14394 (N_14394,N_8288,N_10953);
and U14395 (N_14395,N_10665,N_8932);
nand U14396 (N_14396,N_10828,N_8809);
nor U14397 (N_14397,N_11028,N_10371);
nand U14398 (N_14398,N_10976,N_10451);
nand U14399 (N_14399,N_10010,N_8613);
and U14400 (N_14400,N_8211,N_8535);
nand U14401 (N_14401,N_10355,N_9317);
and U14402 (N_14402,N_11673,N_9420);
or U14403 (N_14403,N_11298,N_8908);
nand U14404 (N_14404,N_11797,N_8383);
and U14405 (N_14405,N_11416,N_9334);
nand U14406 (N_14406,N_10948,N_10616);
nand U14407 (N_14407,N_10084,N_11110);
and U14408 (N_14408,N_11845,N_11746);
nor U14409 (N_14409,N_9112,N_10289);
nand U14410 (N_14410,N_11414,N_9884);
nand U14411 (N_14411,N_11202,N_10272);
nor U14412 (N_14412,N_10747,N_11773);
or U14413 (N_14413,N_10723,N_9217);
nand U14414 (N_14414,N_8867,N_9537);
nor U14415 (N_14415,N_8662,N_9855);
nand U14416 (N_14416,N_11780,N_8971);
nor U14417 (N_14417,N_10769,N_10924);
or U14418 (N_14418,N_10493,N_10577);
nand U14419 (N_14419,N_10724,N_9794);
nand U14420 (N_14420,N_9978,N_8821);
or U14421 (N_14421,N_8479,N_11550);
and U14422 (N_14422,N_8422,N_11024);
nor U14423 (N_14423,N_10326,N_10180);
nand U14424 (N_14424,N_11933,N_9207);
nor U14425 (N_14425,N_11345,N_9561);
or U14426 (N_14426,N_11611,N_11590);
or U14427 (N_14427,N_9859,N_9051);
nor U14428 (N_14428,N_11457,N_11921);
and U14429 (N_14429,N_8646,N_11086);
and U14430 (N_14430,N_10444,N_8812);
and U14431 (N_14431,N_10918,N_10502);
nor U14432 (N_14432,N_8701,N_10915);
and U14433 (N_14433,N_11490,N_9633);
and U14434 (N_14434,N_10913,N_9247);
nor U14435 (N_14435,N_10207,N_11623);
or U14436 (N_14436,N_8119,N_9450);
or U14437 (N_14437,N_9678,N_8908);
and U14438 (N_14438,N_8799,N_10045);
nor U14439 (N_14439,N_8821,N_9145);
nor U14440 (N_14440,N_8400,N_8056);
and U14441 (N_14441,N_8826,N_9735);
and U14442 (N_14442,N_10623,N_11267);
or U14443 (N_14443,N_11506,N_10828);
nor U14444 (N_14444,N_9361,N_11231);
nor U14445 (N_14445,N_11181,N_9314);
or U14446 (N_14446,N_10111,N_11331);
nor U14447 (N_14447,N_9748,N_10090);
or U14448 (N_14448,N_8155,N_9190);
or U14449 (N_14449,N_10570,N_8436);
nor U14450 (N_14450,N_9807,N_11762);
and U14451 (N_14451,N_9235,N_9746);
and U14452 (N_14452,N_8770,N_8719);
nand U14453 (N_14453,N_10941,N_10546);
or U14454 (N_14454,N_9395,N_9057);
or U14455 (N_14455,N_8268,N_11659);
nand U14456 (N_14456,N_10268,N_10760);
nor U14457 (N_14457,N_11691,N_8009);
nor U14458 (N_14458,N_9710,N_11489);
nor U14459 (N_14459,N_8173,N_10951);
nor U14460 (N_14460,N_11521,N_9424);
nor U14461 (N_14461,N_11333,N_9947);
nand U14462 (N_14462,N_11256,N_11315);
and U14463 (N_14463,N_11164,N_11904);
and U14464 (N_14464,N_8931,N_10091);
or U14465 (N_14465,N_11809,N_11171);
or U14466 (N_14466,N_11626,N_11409);
and U14467 (N_14467,N_11322,N_8833);
nor U14468 (N_14468,N_11473,N_9315);
and U14469 (N_14469,N_8164,N_11268);
nand U14470 (N_14470,N_9024,N_10863);
or U14471 (N_14471,N_11485,N_9571);
and U14472 (N_14472,N_8720,N_9939);
nor U14473 (N_14473,N_11432,N_8135);
and U14474 (N_14474,N_8222,N_11332);
or U14475 (N_14475,N_8681,N_10762);
or U14476 (N_14476,N_9861,N_8092);
nor U14477 (N_14477,N_11435,N_8068);
or U14478 (N_14478,N_11607,N_9747);
xnor U14479 (N_14479,N_10676,N_11793);
nor U14480 (N_14480,N_10474,N_8706);
and U14481 (N_14481,N_9012,N_11572);
or U14482 (N_14482,N_8023,N_9844);
nor U14483 (N_14483,N_8866,N_8630);
or U14484 (N_14484,N_8825,N_8892);
nor U14485 (N_14485,N_8843,N_10222);
and U14486 (N_14486,N_11518,N_8126);
or U14487 (N_14487,N_11184,N_11211);
nand U14488 (N_14488,N_9165,N_10125);
and U14489 (N_14489,N_9568,N_9111);
xnor U14490 (N_14490,N_10740,N_8710);
nand U14491 (N_14491,N_8877,N_8490);
nand U14492 (N_14492,N_10758,N_10955);
and U14493 (N_14493,N_8981,N_11658);
or U14494 (N_14494,N_11251,N_10258);
nand U14495 (N_14495,N_8353,N_10951);
nand U14496 (N_14496,N_10556,N_11465);
or U14497 (N_14497,N_9274,N_9897);
nor U14498 (N_14498,N_8105,N_9421);
and U14499 (N_14499,N_9490,N_9362);
or U14500 (N_14500,N_11290,N_9807);
nor U14501 (N_14501,N_8338,N_10151);
nor U14502 (N_14502,N_8694,N_11251);
or U14503 (N_14503,N_8355,N_10912);
or U14504 (N_14504,N_8512,N_8677);
nor U14505 (N_14505,N_8164,N_11529);
xnor U14506 (N_14506,N_10855,N_8582);
or U14507 (N_14507,N_11413,N_10468);
and U14508 (N_14508,N_11729,N_8280);
and U14509 (N_14509,N_8679,N_9961);
or U14510 (N_14510,N_9436,N_11303);
nand U14511 (N_14511,N_9728,N_10104);
nand U14512 (N_14512,N_10554,N_8278);
nand U14513 (N_14513,N_11600,N_8963);
nand U14514 (N_14514,N_10853,N_11962);
nor U14515 (N_14515,N_9658,N_9751);
and U14516 (N_14516,N_9746,N_10111);
nor U14517 (N_14517,N_8747,N_8398);
nor U14518 (N_14518,N_11740,N_9419);
and U14519 (N_14519,N_10742,N_11457);
and U14520 (N_14520,N_8586,N_11703);
or U14521 (N_14521,N_8656,N_11457);
and U14522 (N_14522,N_9289,N_9740);
or U14523 (N_14523,N_11688,N_8633);
nand U14524 (N_14524,N_10714,N_9716);
or U14525 (N_14525,N_9385,N_8370);
and U14526 (N_14526,N_11840,N_9634);
and U14527 (N_14527,N_8422,N_8121);
or U14528 (N_14528,N_10747,N_10703);
xnor U14529 (N_14529,N_11617,N_10484);
or U14530 (N_14530,N_8196,N_8531);
nand U14531 (N_14531,N_10646,N_8070);
nor U14532 (N_14532,N_8654,N_9780);
or U14533 (N_14533,N_10721,N_8411);
nand U14534 (N_14534,N_11451,N_11207);
nor U14535 (N_14535,N_11021,N_8184);
nor U14536 (N_14536,N_10798,N_10213);
or U14537 (N_14537,N_8969,N_11877);
nor U14538 (N_14538,N_11075,N_11552);
nor U14539 (N_14539,N_11217,N_9152);
nor U14540 (N_14540,N_8123,N_9359);
or U14541 (N_14541,N_10234,N_10874);
nand U14542 (N_14542,N_10489,N_11764);
nor U14543 (N_14543,N_8472,N_8877);
or U14544 (N_14544,N_9027,N_11189);
and U14545 (N_14545,N_10335,N_10214);
nor U14546 (N_14546,N_11854,N_8022);
or U14547 (N_14547,N_9887,N_11019);
and U14548 (N_14548,N_10608,N_11989);
nor U14549 (N_14549,N_11313,N_10073);
nand U14550 (N_14550,N_11389,N_11983);
or U14551 (N_14551,N_11876,N_9513);
or U14552 (N_14552,N_10469,N_11745);
nor U14553 (N_14553,N_8543,N_9661);
or U14554 (N_14554,N_10557,N_9323);
or U14555 (N_14555,N_10797,N_11540);
and U14556 (N_14556,N_11719,N_10022);
and U14557 (N_14557,N_10193,N_10166);
and U14558 (N_14558,N_9576,N_9426);
nand U14559 (N_14559,N_11523,N_10924);
nand U14560 (N_14560,N_11026,N_10934);
and U14561 (N_14561,N_8067,N_11371);
and U14562 (N_14562,N_9961,N_8256);
and U14563 (N_14563,N_9632,N_10266);
or U14564 (N_14564,N_10611,N_11746);
or U14565 (N_14565,N_10804,N_11069);
nor U14566 (N_14566,N_11233,N_10741);
and U14567 (N_14567,N_11634,N_9425);
or U14568 (N_14568,N_8506,N_8746);
and U14569 (N_14569,N_8406,N_8725);
nor U14570 (N_14570,N_10109,N_11585);
and U14571 (N_14571,N_11198,N_11935);
nand U14572 (N_14572,N_8444,N_11949);
and U14573 (N_14573,N_9492,N_11629);
xor U14574 (N_14574,N_11589,N_8816);
nand U14575 (N_14575,N_10241,N_10439);
nand U14576 (N_14576,N_9291,N_10026);
and U14577 (N_14577,N_9690,N_10401);
or U14578 (N_14578,N_11807,N_8287);
nand U14579 (N_14579,N_10306,N_9472);
and U14580 (N_14580,N_8543,N_8439);
or U14581 (N_14581,N_11387,N_11910);
nand U14582 (N_14582,N_8206,N_8699);
nor U14583 (N_14583,N_10791,N_9387);
nand U14584 (N_14584,N_8927,N_9577);
or U14585 (N_14585,N_10461,N_9918);
or U14586 (N_14586,N_9693,N_11682);
and U14587 (N_14587,N_10565,N_10227);
nand U14588 (N_14588,N_10748,N_8875);
nand U14589 (N_14589,N_8700,N_9703);
and U14590 (N_14590,N_9056,N_10729);
and U14591 (N_14591,N_8637,N_10742);
nor U14592 (N_14592,N_9697,N_10230);
or U14593 (N_14593,N_11112,N_9498);
or U14594 (N_14594,N_9643,N_10641);
and U14595 (N_14595,N_11835,N_9495);
or U14596 (N_14596,N_10368,N_9556);
nor U14597 (N_14597,N_9793,N_9918);
or U14598 (N_14598,N_10385,N_11459);
nand U14599 (N_14599,N_10308,N_11745);
or U14600 (N_14600,N_8515,N_9845);
or U14601 (N_14601,N_8527,N_9621);
and U14602 (N_14602,N_11873,N_8416);
or U14603 (N_14603,N_10601,N_11406);
and U14604 (N_14604,N_9089,N_11561);
nand U14605 (N_14605,N_9377,N_10962);
and U14606 (N_14606,N_10399,N_11113);
and U14607 (N_14607,N_11725,N_9669);
nand U14608 (N_14608,N_11823,N_8029);
and U14609 (N_14609,N_8991,N_10556);
nand U14610 (N_14610,N_11868,N_10004);
and U14611 (N_14611,N_9724,N_10295);
or U14612 (N_14612,N_9196,N_9228);
nand U14613 (N_14613,N_9161,N_9401);
and U14614 (N_14614,N_10552,N_8384);
nand U14615 (N_14615,N_11222,N_10371);
or U14616 (N_14616,N_9071,N_9429);
and U14617 (N_14617,N_11784,N_11994);
and U14618 (N_14618,N_8894,N_11544);
nor U14619 (N_14619,N_10739,N_9906);
and U14620 (N_14620,N_11083,N_8765);
or U14621 (N_14621,N_9726,N_10491);
or U14622 (N_14622,N_9311,N_10470);
and U14623 (N_14623,N_8405,N_9184);
nor U14624 (N_14624,N_10472,N_10062);
nand U14625 (N_14625,N_8509,N_10763);
nor U14626 (N_14626,N_9167,N_9909);
and U14627 (N_14627,N_8131,N_10125);
nand U14628 (N_14628,N_9894,N_8230);
or U14629 (N_14629,N_11618,N_8583);
or U14630 (N_14630,N_10589,N_11708);
nor U14631 (N_14631,N_9032,N_9445);
nor U14632 (N_14632,N_11514,N_10338);
and U14633 (N_14633,N_9821,N_8960);
or U14634 (N_14634,N_10951,N_11722);
and U14635 (N_14635,N_9118,N_8480);
nor U14636 (N_14636,N_8808,N_9627);
nand U14637 (N_14637,N_11597,N_8182);
nand U14638 (N_14638,N_10483,N_10311);
and U14639 (N_14639,N_9038,N_8153);
and U14640 (N_14640,N_11872,N_8661);
or U14641 (N_14641,N_10513,N_8175);
and U14642 (N_14642,N_10581,N_10510);
nor U14643 (N_14643,N_10532,N_8433);
xor U14644 (N_14644,N_11776,N_10373);
nand U14645 (N_14645,N_8905,N_9142);
or U14646 (N_14646,N_9147,N_8881);
or U14647 (N_14647,N_8705,N_10335);
and U14648 (N_14648,N_10426,N_8683);
nor U14649 (N_14649,N_10672,N_10005);
xnor U14650 (N_14650,N_8373,N_9193);
and U14651 (N_14651,N_8604,N_11720);
nor U14652 (N_14652,N_8254,N_9745);
nand U14653 (N_14653,N_9958,N_9101);
nand U14654 (N_14654,N_11568,N_9533);
or U14655 (N_14655,N_11155,N_11413);
and U14656 (N_14656,N_11486,N_10589);
nand U14657 (N_14657,N_11839,N_11716);
nand U14658 (N_14658,N_10787,N_10616);
and U14659 (N_14659,N_11213,N_11978);
or U14660 (N_14660,N_8196,N_10404);
nand U14661 (N_14661,N_9389,N_11781);
nor U14662 (N_14662,N_9639,N_9770);
nor U14663 (N_14663,N_8125,N_11864);
or U14664 (N_14664,N_9977,N_8685);
and U14665 (N_14665,N_9519,N_11263);
and U14666 (N_14666,N_11773,N_10948);
or U14667 (N_14667,N_11339,N_9440);
or U14668 (N_14668,N_11513,N_11843);
nor U14669 (N_14669,N_8277,N_8865);
or U14670 (N_14670,N_10666,N_9411);
and U14671 (N_14671,N_10435,N_10308);
nand U14672 (N_14672,N_8982,N_11340);
nor U14673 (N_14673,N_11639,N_11339);
nand U14674 (N_14674,N_8997,N_9148);
nor U14675 (N_14675,N_9565,N_9017);
and U14676 (N_14676,N_8767,N_8921);
and U14677 (N_14677,N_11408,N_10865);
nor U14678 (N_14678,N_9429,N_9800);
and U14679 (N_14679,N_10763,N_9772);
and U14680 (N_14680,N_9351,N_11341);
nor U14681 (N_14681,N_8653,N_9060);
or U14682 (N_14682,N_9001,N_8258);
nor U14683 (N_14683,N_11022,N_8525);
nor U14684 (N_14684,N_11577,N_8989);
nor U14685 (N_14685,N_11274,N_8701);
or U14686 (N_14686,N_8693,N_8113);
nand U14687 (N_14687,N_8340,N_9885);
nand U14688 (N_14688,N_10383,N_9310);
and U14689 (N_14689,N_10171,N_8704);
or U14690 (N_14690,N_9552,N_11544);
and U14691 (N_14691,N_11961,N_10598);
nor U14692 (N_14692,N_8605,N_10309);
nand U14693 (N_14693,N_10675,N_9275);
nand U14694 (N_14694,N_10973,N_11307);
and U14695 (N_14695,N_10530,N_8548);
and U14696 (N_14696,N_8099,N_9298);
nand U14697 (N_14697,N_9563,N_9427);
nor U14698 (N_14698,N_9517,N_8994);
nand U14699 (N_14699,N_8237,N_8090);
or U14700 (N_14700,N_8134,N_8691);
and U14701 (N_14701,N_11096,N_10557);
and U14702 (N_14702,N_10538,N_11296);
nor U14703 (N_14703,N_10825,N_11136);
or U14704 (N_14704,N_8770,N_8666);
or U14705 (N_14705,N_10888,N_10370);
and U14706 (N_14706,N_10908,N_9820);
and U14707 (N_14707,N_11872,N_8543);
nand U14708 (N_14708,N_9200,N_8286);
and U14709 (N_14709,N_9539,N_9309);
nand U14710 (N_14710,N_10420,N_9783);
nor U14711 (N_14711,N_10769,N_8377);
nor U14712 (N_14712,N_10051,N_8490);
nor U14713 (N_14713,N_11367,N_8678);
nand U14714 (N_14714,N_8440,N_10351);
or U14715 (N_14715,N_11306,N_8705);
nor U14716 (N_14716,N_11737,N_11250);
or U14717 (N_14717,N_8589,N_11825);
or U14718 (N_14718,N_11420,N_8579);
nand U14719 (N_14719,N_11499,N_10396);
and U14720 (N_14720,N_11098,N_11575);
nand U14721 (N_14721,N_8508,N_10200);
or U14722 (N_14722,N_11125,N_10599);
nor U14723 (N_14723,N_10117,N_11676);
or U14724 (N_14724,N_11790,N_11533);
and U14725 (N_14725,N_9839,N_9638);
and U14726 (N_14726,N_10783,N_8174);
nand U14727 (N_14727,N_8970,N_11608);
xor U14728 (N_14728,N_8114,N_11961);
nor U14729 (N_14729,N_8280,N_11483);
or U14730 (N_14730,N_11606,N_8468);
nor U14731 (N_14731,N_10131,N_10878);
nor U14732 (N_14732,N_9704,N_8126);
nor U14733 (N_14733,N_11549,N_10433);
xnor U14734 (N_14734,N_9519,N_9256);
and U14735 (N_14735,N_8669,N_11761);
nor U14736 (N_14736,N_11633,N_8325);
and U14737 (N_14737,N_11662,N_8504);
nor U14738 (N_14738,N_9698,N_11313);
nand U14739 (N_14739,N_10568,N_11408);
nand U14740 (N_14740,N_10133,N_8033);
and U14741 (N_14741,N_9709,N_10702);
nor U14742 (N_14742,N_8832,N_8324);
nand U14743 (N_14743,N_9204,N_9838);
and U14744 (N_14744,N_10239,N_9296);
nand U14745 (N_14745,N_8553,N_10498);
nor U14746 (N_14746,N_10740,N_9211);
and U14747 (N_14747,N_8068,N_8928);
nand U14748 (N_14748,N_9000,N_9170);
and U14749 (N_14749,N_10993,N_11599);
or U14750 (N_14750,N_11414,N_11417);
or U14751 (N_14751,N_8992,N_11234);
nand U14752 (N_14752,N_8358,N_8391);
nand U14753 (N_14753,N_11361,N_11192);
nand U14754 (N_14754,N_10548,N_8847);
or U14755 (N_14755,N_8576,N_9755);
nor U14756 (N_14756,N_11762,N_8719);
nor U14757 (N_14757,N_10576,N_8854);
nand U14758 (N_14758,N_9629,N_9594);
or U14759 (N_14759,N_9190,N_10254);
or U14760 (N_14760,N_11304,N_11789);
nand U14761 (N_14761,N_11092,N_8606);
and U14762 (N_14762,N_10145,N_8881);
xnor U14763 (N_14763,N_8278,N_9255);
nand U14764 (N_14764,N_9257,N_9331);
or U14765 (N_14765,N_9160,N_9594);
and U14766 (N_14766,N_8157,N_11134);
and U14767 (N_14767,N_8758,N_11996);
or U14768 (N_14768,N_10783,N_8852);
or U14769 (N_14769,N_9749,N_11016);
or U14770 (N_14770,N_8019,N_10265);
xor U14771 (N_14771,N_9207,N_9812);
or U14772 (N_14772,N_10426,N_8492);
nand U14773 (N_14773,N_10549,N_11087);
or U14774 (N_14774,N_8806,N_10933);
and U14775 (N_14775,N_8314,N_9086);
nor U14776 (N_14776,N_9861,N_9898);
or U14777 (N_14777,N_11896,N_10073);
nand U14778 (N_14778,N_9561,N_8195);
nand U14779 (N_14779,N_9067,N_11870);
and U14780 (N_14780,N_11053,N_8779);
nor U14781 (N_14781,N_11058,N_10388);
nand U14782 (N_14782,N_11247,N_10646);
and U14783 (N_14783,N_11131,N_11824);
nor U14784 (N_14784,N_8240,N_11217);
or U14785 (N_14785,N_8452,N_9465);
and U14786 (N_14786,N_9526,N_10233);
or U14787 (N_14787,N_11016,N_10607);
nand U14788 (N_14788,N_10692,N_8237);
nand U14789 (N_14789,N_8819,N_11536);
and U14790 (N_14790,N_11601,N_8078);
nand U14791 (N_14791,N_10215,N_10353);
or U14792 (N_14792,N_10062,N_11651);
nand U14793 (N_14793,N_11725,N_9989);
nor U14794 (N_14794,N_9882,N_11186);
nand U14795 (N_14795,N_10411,N_11830);
nor U14796 (N_14796,N_10361,N_9765);
nor U14797 (N_14797,N_9159,N_11367);
and U14798 (N_14798,N_11876,N_10883);
and U14799 (N_14799,N_9608,N_10416);
xnor U14800 (N_14800,N_10461,N_11872);
and U14801 (N_14801,N_10221,N_11828);
nand U14802 (N_14802,N_8081,N_10979);
nor U14803 (N_14803,N_9113,N_10127);
nand U14804 (N_14804,N_11571,N_9942);
and U14805 (N_14805,N_9791,N_11028);
nor U14806 (N_14806,N_10587,N_9963);
nor U14807 (N_14807,N_10908,N_11310);
nor U14808 (N_14808,N_9225,N_10149);
nor U14809 (N_14809,N_9807,N_9374);
nor U14810 (N_14810,N_8610,N_11020);
nand U14811 (N_14811,N_11911,N_11174);
and U14812 (N_14812,N_9200,N_8055);
nand U14813 (N_14813,N_8970,N_10490);
and U14814 (N_14814,N_10254,N_8096);
nand U14815 (N_14815,N_8253,N_8857);
and U14816 (N_14816,N_10959,N_9837);
nand U14817 (N_14817,N_11767,N_10698);
and U14818 (N_14818,N_10614,N_10637);
and U14819 (N_14819,N_9292,N_8670);
or U14820 (N_14820,N_10728,N_10341);
or U14821 (N_14821,N_11721,N_10146);
and U14822 (N_14822,N_9934,N_10942);
nand U14823 (N_14823,N_8127,N_10634);
or U14824 (N_14824,N_11714,N_8631);
or U14825 (N_14825,N_10708,N_8733);
nor U14826 (N_14826,N_8224,N_10808);
nand U14827 (N_14827,N_8816,N_11572);
nand U14828 (N_14828,N_9604,N_9558);
or U14829 (N_14829,N_8885,N_10913);
nand U14830 (N_14830,N_8460,N_11803);
nor U14831 (N_14831,N_8851,N_8551);
nor U14832 (N_14832,N_8255,N_11936);
nor U14833 (N_14833,N_9199,N_8159);
nor U14834 (N_14834,N_9840,N_11799);
nand U14835 (N_14835,N_9383,N_10691);
nor U14836 (N_14836,N_10517,N_11104);
or U14837 (N_14837,N_9025,N_9506);
nand U14838 (N_14838,N_9981,N_11865);
or U14839 (N_14839,N_11518,N_8544);
nand U14840 (N_14840,N_9999,N_8810);
nor U14841 (N_14841,N_8532,N_8211);
and U14842 (N_14842,N_9332,N_8894);
and U14843 (N_14843,N_8892,N_9897);
and U14844 (N_14844,N_9673,N_10926);
or U14845 (N_14845,N_10187,N_11676);
and U14846 (N_14846,N_11070,N_10758);
nor U14847 (N_14847,N_10353,N_9906);
nor U14848 (N_14848,N_9654,N_9984);
and U14849 (N_14849,N_11224,N_9396);
nor U14850 (N_14850,N_9570,N_11818);
and U14851 (N_14851,N_11334,N_8457);
nand U14852 (N_14852,N_9434,N_11701);
and U14853 (N_14853,N_10364,N_11437);
nand U14854 (N_14854,N_8150,N_8680);
nor U14855 (N_14855,N_10428,N_9547);
or U14856 (N_14856,N_11944,N_8552);
or U14857 (N_14857,N_9405,N_10667);
or U14858 (N_14858,N_10898,N_9075);
or U14859 (N_14859,N_8209,N_11847);
xor U14860 (N_14860,N_8793,N_11814);
or U14861 (N_14861,N_9036,N_8456);
and U14862 (N_14862,N_8348,N_9236);
nand U14863 (N_14863,N_8879,N_8731);
or U14864 (N_14864,N_8306,N_8675);
and U14865 (N_14865,N_10961,N_8893);
nor U14866 (N_14866,N_8149,N_9573);
nor U14867 (N_14867,N_11136,N_10614);
nand U14868 (N_14868,N_8757,N_8162);
nand U14869 (N_14869,N_8412,N_8930);
or U14870 (N_14870,N_9918,N_8835);
and U14871 (N_14871,N_10499,N_11374);
nor U14872 (N_14872,N_9378,N_11364);
and U14873 (N_14873,N_10287,N_9642);
and U14874 (N_14874,N_8121,N_10199);
or U14875 (N_14875,N_10084,N_10929);
or U14876 (N_14876,N_11351,N_10368);
nand U14877 (N_14877,N_10853,N_11587);
and U14878 (N_14878,N_11655,N_8793);
nor U14879 (N_14879,N_10529,N_11931);
nand U14880 (N_14880,N_8125,N_9956);
nand U14881 (N_14881,N_10287,N_10715);
or U14882 (N_14882,N_10473,N_11010);
nor U14883 (N_14883,N_11442,N_9010);
or U14884 (N_14884,N_9399,N_10633);
xor U14885 (N_14885,N_10556,N_8134);
and U14886 (N_14886,N_8161,N_8733);
and U14887 (N_14887,N_10620,N_8769);
nand U14888 (N_14888,N_10310,N_8758);
and U14889 (N_14889,N_11678,N_10104);
nand U14890 (N_14890,N_8183,N_11467);
and U14891 (N_14891,N_9498,N_10595);
nor U14892 (N_14892,N_8782,N_8196);
nand U14893 (N_14893,N_8341,N_11098);
xor U14894 (N_14894,N_8818,N_8440);
nand U14895 (N_14895,N_9380,N_10679);
and U14896 (N_14896,N_10967,N_10133);
or U14897 (N_14897,N_9026,N_11911);
or U14898 (N_14898,N_9819,N_9528);
nor U14899 (N_14899,N_9760,N_8184);
or U14900 (N_14900,N_9611,N_11345);
nor U14901 (N_14901,N_11399,N_11960);
nor U14902 (N_14902,N_9615,N_9560);
nand U14903 (N_14903,N_9586,N_8349);
nor U14904 (N_14904,N_11764,N_11970);
nor U14905 (N_14905,N_9508,N_10567);
or U14906 (N_14906,N_8089,N_10197);
nand U14907 (N_14907,N_10499,N_9188);
or U14908 (N_14908,N_9098,N_11557);
nand U14909 (N_14909,N_10729,N_8561);
nor U14910 (N_14910,N_9839,N_9718);
and U14911 (N_14911,N_11244,N_9207);
or U14912 (N_14912,N_11903,N_11898);
nor U14913 (N_14913,N_11338,N_9968);
nand U14914 (N_14914,N_11708,N_11326);
or U14915 (N_14915,N_9041,N_11796);
nor U14916 (N_14916,N_8483,N_10366);
nor U14917 (N_14917,N_9568,N_8090);
or U14918 (N_14918,N_11975,N_10224);
or U14919 (N_14919,N_10354,N_10410);
and U14920 (N_14920,N_10327,N_9328);
nand U14921 (N_14921,N_9295,N_11074);
or U14922 (N_14922,N_10073,N_8765);
nor U14923 (N_14923,N_9376,N_11038);
xnor U14924 (N_14924,N_10601,N_8709);
or U14925 (N_14925,N_11552,N_11437);
nor U14926 (N_14926,N_11235,N_9764);
or U14927 (N_14927,N_11208,N_10989);
nand U14928 (N_14928,N_11456,N_9443);
or U14929 (N_14929,N_11885,N_11881);
and U14930 (N_14930,N_8724,N_9904);
nor U14931 (N_14931,N_10697,N_8129);
nand U14932 (N_14932,N_11412,N_9734);
nor U14933 (N_14933,N_11029,N_10504);
nor U14934 (N_14934,N_9028,N_9166);
or U14935 (N_14935,N_10222,N_9153);
and U14936 (N_14936,N_8774,N_11155);
or U14937 (N_14937,N_11139,N_10355);
nor U14938 (N_14938,N_8873,N_9348);
nand U14939 (N_14939,N_11290,N_10133);
nor U14940 (N_14940,N_8317,N_8877);
nor U14941 (N_14941,N_10325,N_8942);
and U14942 (N_14942,N_11484,N_10160);
nor U14943 (N_14943,N_11282,N_11299);
or U14944 (N_14944,N_11285,N_10042);
or U14945 (N_14945,N_10408,N_9897);
nor U14946 (N_14946,N_9825,N_9659);
nor U14947 (N_14947,N_11477,N_10477);
and U14948 (N_14948,N_11182,N_9881);
nor U14949 (N_14949,N_10206,N_8263);
nand U14950 (N_14950,N_10899,N_9157);
nand U14951 (N_14951,N_8832,N_10119);
and U14952 (N_14952,N_9350,N_8015);
nand U14953 (N_14953,N_10511,N_8267);
nor U14954 (N_14954,N_11554,N_8723);
nor U14955 (N_14955,N_11507,N_11620);
nand U14956 (N_14956,N_8691,N_10042);
and U14957 (N_14957,N_10292,N_9170);
nand U14958 (N_14958,N_8469,N_10203);
nand U14959 (N_14959,N_10468,N_11830);
nand U14960 (N_14960,N_9323,N_8736);
nor U14961 (N_14961,N_8501,N_8313);
nand U14962 (N_14962,N_11901,N_10352);
or U14963 (N_14963,N_10865,N_11475);
or U14964 (N_14964,N_10551,N_8447);
nand U14965 (N_14965,N_10849,N_10894);
nand U14966 (N_14966,N_9628,N_11484);
nand U14967 (N_14967,N_9709,N_10744);
and U14968 (N_14968,N_11842,N_8671);
nor U14969 (N_14969,N_10324,N_8898);
nor U14970 (N_14970,N_10759,N_11583);
nand U14971 (N_14971,N_9125,N_10476);
nand U14972 (N_14972,N_8429,N_11486);
nor U14973 (N_14973,N_8214,N_8229);
or U14974 (N_14974,N_9067,N_9251);
nand U14975 (N_14975,N_8817,N_10637);
and U14976 (N_14976,N_10801,N_9136);
and U14977 (N_14977,N_10524,N_11634);
nand U14978 (N_14978,N_10224,N_11166);
nand U14979 (N_14979,N_11495,N_10085);
and U14980 (N_14980,N_11199,N_9853);
nor U14981 (N_14981,N_9018,N_10987);
or U14982 (N_14982,N_9014,N_8120);
and U14983 (N_14983,N_10725,N_9590);
nor U14984 (N_14984,N_10899,N_9236);
or U14985 (N_14985,N_10384,N_10093);
and U14986 (N_14986,N_10760,N_11593);
or U14987 (N_14987,N_10496,N_8717);
nand U14988 (N_14988,N_11929,N_11743);
and U14989 (N_14989,N_11173,N_8057);
nand U14990 (N_14990,N_10299,N_9186);
nor U14991 (N_14991,N_8977,N_8342);
and U14992 (N_14992,N_10394,N_10633);
or U14993 (N_14993,N_10482,N_11449);
or U14994 (N_14994,N_10932,N_10325);
or U14995 (N_14995,N_9548,N_8835);
nand U14996 (N_14996,N_11425,N_9766);
or U14997 (N_14997,N_10699,N_11790);
nand U14998 (N_14998,N_11722,N_9789);
or U14999 (N_14999,N_10354,N_11321);
or U15000 (N_15000,N_10986,N_8887);
and U15001 (N_15001,N_8857,N_11406);
nor U15002 (N_15002,N_10425,N_11124);
or U15003 (N_15003,N_10693,N_10439);
and U15004 (N_15004,N_11185,N_11470);
nor U15005 (N_15005,N_11209,N_10554);
nand U15006 (N_15006,N_11238,N_8558);
nand U15007 (N_15007,N_10829,N_10181);
or U15008 (N_15008,N_8102,N_9870);
nand U15009 (N_15009,N_10593,N_9483);
and U15010 (N_15010,N_11809,N_10453);
nand U15011 (N_15011,N_11814,N_11027);
or U15012 (N_15012,N_10231,N_10689);
or U15013 (N_15013,N_10549,N_8055);
nand U15014 (N_15014,N_9953,N_11498);
nand U15015 (N_15015,N_9882,N_8673);
or U15016 (N_15016,N_9952,N_11127);
nand U15017 (N_15017,N_10041,N_8160);
nor U15018 (N_15018,N_11145,N_11621);
nor U15019 (N_15019,N_8875,N_10015);
and U15020 (N_15020,N_11717,N_10489);
nand U15021 (N_15021,N_10732,N_9648);
or U15022 (N_15022,N_11999,N_10661);
nand U15023 (N_15023,N_8878,N_8750);
or U15024 (N_15024,N_11226,N_11713);
or U15025 (N_15025,N_10500,N_10454);
nand U15026 (N_15026,N_11812,N_10309);
nor U15027 (N_15027,N_10827,N_11008);
nand U15028 (N_15028,N_9549,N_9513);
nand U15029 (N_15029,N_11350,N_8873);
and U15030 (N_15030,N_8280,N_9169);
nand U15031 (N_15031,N_10289,N_8554);
or U15032 (N_15032,N_8832,N_11968);
or U15033 (N_15033,N_10374,N_8760);
or U15034 (N_15034,N_10979,N_8330);
nor U15035 (N_15035,N_9155,N_10865);
and U15036 (N_15036,N_9905,N_8423);
and U15037 (N_15037,N_10163,N_9383);
xnor U15038 (N_15038,N_9462,N_8767);
or U15039 (N_15039,N_11890,N_10288);
and U15040 (N_15040,N_8392,N_11768);
nor U15041 (N_15041,N_9380,N_8372);
or U15042 (N_15042,N_11529,N_10699);
or U15043 (N_15043,N_10604,N_10311);
and U15044 (N_15044,N_11406,N_8633);
or U15045 (N_15045,N_9592,N_8342);
or U15046 (N_15046,N_8832,N_9779);
nand U15047 (N_15047,N_8749,N_11789);
nand U15048 (N_15048,N_9988,N_8590);
or U15049 (N_15049,N_11572,N_11474);
nor U15050 (N_15050,N_10167,N_11054);
nand U15051 (N_15051,N_10415,N_9476);
nand U15052 (N_15052,N_8185,N_10016);
and U15053 (N_15053,N_10929,N_10605);
or U15054 (N_15054,N_10705,N_9475);
nand U15055 (N_15055,N_9340,N_8924);
or U15056 (N_15056,N_10106,N_9522);
nor U15057 (N_15057,N_11098,N_8701);
or U15058 (N_15058,N_8971,N_8450);
nor U15059 (N_15059,N_8014,N_11134);
nor U15060 (N_15060,N_10652,N_11505);
nor U15061 (N_15061,N_9936,N_10561);
and U15062 (N_15062,N_11780,N_8717);
or U15063 (N_15063,N_10284,N_8062);
nand U15064 (N_15064,N_8861,N_10749);
and U15065 (N_15065,N_11439,N_10605);
or U15066 (N_15066,N_8601,N_11126);
nor U15067 (N_15067,N_9381,N_11772);
or U15068 (N_15068,N_9442,N_8590);
nor U15069 (N_15069,N_9395,N_8221);
and U15070 (N_15070,N_9611,N_8162);
and U15071 (N_15071,N_10942,N_11271);
nand U15072 (N_15072,N_8281,N_8192);
or U15073 (N_15073,N_11776,N_11855);
and U15074 (N_15074,N_11370,N_10618);
nor U15075 (N_15075,N_9173,N_9802);
or U15076 (N_15076,N_8097,N_11010);
nand U15077 (N_15077,N_10276,N_9143);
or U15078 (N_15078,N_10920,N_10318);
nor U15079 (N_15079,N_11711,N_8191);
or U15080 (N_15080,N_9802,N_8871);
and U15081 (N_15081,N_9263,N_8293);
and U15082 (N_15082,N_8053,N_8528);
nand U15083 (N_15083,N_9772,N_11559);
nor U15084 (N_15084,N_8105,N_9427);
or U15085 (N_15085,N_11168,N_9733);
and U15086 (N_15086,N_10504,N_11671);
or U15087 (N_15087,N_8438,N_10714);
nor U15088 (N_15088,N_11824,N_11287);
and U15089 (N_15089,N_11802,N_11219);
or U15090 (N_15090,N_10020,N_8640);
nand U15091 (N_15091,N_8410,N_9682);
or U15092 (N_15092,N_9029,N_8182);
nand U15093 (N_15093,N_9406,N_9216);
nand U15094 (N_15094,N_9710,N_9779);
nand U15095 (N_15095,N_9325,N_9335);
or U15096 (N_15096,N_10978,N_8172);
and U15097 (N_15097,N_9659,N_9057);
and U15098 (N_15098,N_10536,N_8120);
or U15099 (N_15099,N_10858,N_11581);
or U15100 (N_15100,N_9199,N_9524);
and U15101 (N_15101,N_9215,N_8716);
and U15102 (N_15102,N_8235,N_9539);
or U15103 (N_15103,N_8600,N_8879);
and U15104 (N_15104,N_8370,N_11994);
and U15105 (N_15105,N_10916,N_11796);
and U15106 (N_15106,N_8383,N_9775);
or U15107 (N_15107,N_9376,N_8894);
or U15108 (N_15108,N_8659,N_9919);
nor U15109 (N_15109,N_10538,N_11270);
or U15110 (N_15110,N_10089,N_11322);
and U15111 (N_15111,N_9317,N_11573);
and U15112 (N_15112,N_9723,N_9309);
or U15113 (N_15113,N_11998,N_11653);
and U15114 (N_15114,N_10429,N_11885);
nor U15115 (N_15115,N_8437,N_8875);
nand U15116 (N_15116,N_8232,N_9700);
nand U15117 (N_15117,N_9384,N_9161);
nor U15118 (N_15118,N_10788,N_9383);
nand U15119 (N_15119,N_8741,N_8493);
or U15120 (N_15120,N_8444,N_10252);
nor U15121 (N_15121,N_9867,N_9284);
nor U15122 (N_15122,N_8133,N_11731);
nand U15123 (N_15123,N_8783,N_11939);
and U15124 (N_15124,N_11052,N_8353);
and U15125 (N_15125,N_10847,N_9489);
and U15126 (N_15126,N_8971,N_10342);
and U15127 (N_15127,N_8827,N_8848);
and U15128 (N_15128,N_11800,N_9625);
nand U15129 (N_15129,N_9551,N_11732);
or U15130 (N_15130,N_8485,N_10196);
or U15131 (N_15131,N_9438,N_11284);
or U15132 (N_15132,N_10827,N_8016);
or U15133 (N_15133,N_11497,N_9660);
nand U15134 (N_15134,N_9456,N_8568);
nand U15135 (N_15135,N_10260,N_10032);
or U15136 (N_15136,N_10504,N_8863);
or U15137 (N_15137,N_9907,N_10695);
nor U15138 (N_15138,N_8739,N_11507);
nor U15139 (N_15139,N_11682,N_9272);
or U15140 (N_15140,N_9820,N_9655);
or U15141 (N_15141,N_9090,N_10522);
nand U15142 (N_15142,N_8608,N_10410);
and U15143 (N_15143,N_10197,N_8116);
nor U15144 (N_15144,N_10302,N_8865);
nor U15145 (N_15145,N_10171,N_9370);
nor U15146 (N_15146,N_8621,N_11651);
or U15147 (N_15147,N_9260,N_10795);
and U15148 (N_15148,N_10898,N_8036);
nand U15149 (N_15149,N_9746,N_8868);
nand U15150 (N_15150,N_8593,N_8459);
and U15151 (N_15151,N_11758,N_8816);
nand U15152 (N_15152,N_11025,N_11877);
or U15153 (N_15153,N_9337,N_10924);
nor U15154 (N_15154,N_8187,N_8296);
or U15155 (N_15155,N_8330,N_9142);
and U15156 (N_15156,N_9442,N_10915);
or U15157 (N_15157,N_8496,N_11828);
nor U15158 (N_15158,N_9886,N_11159);
or U15159 (N_15159,N_10059,N_11782);
nor U15160 (N_15160,N_11717,N_10568);
nand U15161 (N_15161,N_11653,N_9988);
or U15162 (N_15162,N_8186,N_10995);
and U15163 (N_15163,N_9167,N_10578);
and U15164 (N_15164,N_11509,N_10378);
or U15165 (N_15165,N_11195,N_8800);
and U15166 (N_15166,N_9371,N_8389);
nor U15167 (N_15167,N_8138,N_11860);
and U15168 (N_15168,N_11240,N_8377);
or U15169 (N_15169,N_10252,N_11499);
or U15170 (N_15170,N_8081,N_10713);
and U15171 (N_15171,N_9674,N_11527);
nor U15172 (N_15172,N_10376,N_8731);
or U15173 (N_15173,N_11017,N_8224);
and U15174 (N_15174,N_11886,N_10825);
or U15175 (N_15175,N_11698,N_10923);
and U15176 (N_15176,N_11708,N_11004);
nor U15177 (N_15177,N_10765,N_10635);
and U15178 (N_15178,N_8467,N_9196);
nand U15179 (N_15179,N_11653,N_10767);
nand U15180 (N_15180,N_10993,N_10648);
or U15181 (N_15181,N_10604,N_9598);
nand U15182 (N_15182,N_11712,N_10413);
or U15183 (N_15183,N_8354,N_10580);
and U15184 (N_15184,N_10898,N_9406);
or U15185 (N_15185,N_10698,N_8219);
or U15186 (N_15186,N_11065,N_11461);
and U15187 (N_15187,N_8894,N_10647);
nor U15188 (N_15188,N_8445,N_8496);
or U15189 (N_15189,N_9487,N_11497);
nand U15190 (N_15190,N_9701,N_8626);
nor U15191 (N_15191,N_10605,N_9461);
nand U15192 (N_15192,N_8900,N_9418);
nand U15193 (N_15193,N_9039,N_11970);
and U15194 (N_15194,N_8157,N_10784);
and U15195 (N_15195,N_10417,N_10511);
nor U15196 (N_15196,N_10890,N_10649);
nor U15197 (N_15197,N_11821,N_8395);
nand U15198 (N_15198,N_10211,N_8344);
and U15199 (N_15199,N_11957,N_11559);
nand U15200 (N_15200,N_11658,N_9767);
and U15201 (N_15201,N_8225,N_11677);
nand U15202 (N_15202,N_11235,N_10748);
nand U15203 (N_15203,N_8876,N_10953);
or U15204 (N_15204,N_11973,N_10794);
or U15205 (N_15205,N_10482,N_9512);
nor U15206 (N_15206,N_10504,N_9578);
nor U15207 (N_15207,N_8393,N_8599);
nand U15208 (N_15208,N_8491,N_11329);
nor U15209 (N_15209,N_8638,N_11177);
or U15210 (N_15210,N_10136,N_8331);
or U15211 (N_15211,N_11463,N_8750);
or U15212 (N_15212,N_9652,N_8997);
nand U15213 (N_15213,N_11710,N_9084);
nand U15214 (N_15214,N_8512,N_8807);
nand U15215 (N_15215,N_11745,N_10647);
nor U15216 (N_15216,N_8945,N_11321);
or U15217 (N_15217,N_10846,N_11003);
nand U15218 (N_15218,N_8001,N_8190);
nor U15219 (N_15219,N_9517,N_9786);
and U15220 (N_15220,N_11100,N_8117);
and U15221 (N_15221,N_10198,N_9087);
and U15222 (N_15222,N_9959,N_10959);
nor U15223 (N_15223,N_11516,N_8270);
nor U15224 (N_15224,N_9501,N_9640);
nor U15225 (N_15225,N_9844,N_10419);
nor U15226 (N_15226,N_11129,N_9532);
nor U15227 (N_15227,N_11217,N_8758);
nand U15228 (N_15228,N_9165,N_8172);
or U15229 (N_15229,N_11746,N_11859);
and U15230 (N_15230,N_8034,N_9831);
and U15231 (N_15231,N_9427,N_9637);
and U15232 (N_15232,N_8107,N_8334);
and U15233 (N_15233,N_10851,N_8879);
and U15234 (N_15234,N_8553,N_10472);
and U15235 (N_15235,N_11275,N_9716);
nor U15236 (N_15236,N_9286,N_9647);
or U15237 (N_15237,N_8450,N_10501);
nand U15238 (N_15238,N_11765,N_10974);
and U15239 (N_15239,N_9850,N_8404);
nor U15240 (N_15240,N_10863,N_9090);
or U15241 (N_15241,N_10223,N_8654);
nor U15242 (N_15242,N_11099,N_11113);
and U15243 (N_15243,N_10519,N_8674);
nor U15244 (N_15244,N_10061,N_10689);
and U15245 (N_15245,N_10776,N_11995);
nor U15246 (N_15246,N_11479,N_11093);
nor U15247 (N_15247,N_11012,N_10227);
and U15248 (N_15248,N_11578,N_10366);
nor U15249 (N_15249,N_8649,N_8647);
and U15250 (N_15250,N_11050,N_11697);
nand U15251 (N_15251,N_10783,N_11836);
and U15252 (N_15252,N_11045,N_10585);
nor U15253 (N_15253,N_10450,N_10042);
nor U15254 (N_15254,N_10970,N_10686);
nand U15255 (N_15255,N_10760,N_8452);
or U15256 (N_15256,N_10642,N_10416);
or U15257 (N_15257,N_9661,N_11272);
or U15258 (N_15258,N_8587,N_11785);
or U15259 (N_15259,N_11271,N_9865);
and U15260 (N_15260,N_9508,N_11560);
nor U15261 (N_15261,N_10029,N_10102);
and U15262 (N_15262,N_9729,N_11531);
nor U15263 (N_15263,N_9406,N_10599);
nor U15264 (N_15264,N_9476,N_11579);
nand U15265 (N_15265,N_11512,N_11572);
or U15266 (N_15266,N_8681,N_10873);
or U15267 (N_15267,N_9313,N_9090);
nand U15268 (N_15268,N_11451,N_8679);
nor U15269 (N_15269,N_10543,N_8932);
nand U15270 (N_15270,N_11907,N_9244);
nand U15271 (N_15271,N_9577,N_9666);
and U15272 (N_15272,N_9364,N_8613);
and U15273 (N_15273,N_8101,N_9315);
and U15274 (N_15274,N_9174,N_8965);
nor U15275 (N_15275,N_8750,N_8438);
nand U15276 (N_15276,N_8628,N_8188);
nor U15277 (N_15277,N_8198,N_8392);
or U15278 (N_15278,N_8393,N_11720);
or U15279 (N_15279,N_11083,N_8902);
or U15280 (N_15280,N_11083,N_8036);
nor U15281 (N_15281,N_9243,N_8872);
or U15282 (N_15282,N_10085,N_9799);
nor U15283 (N_15283,N_9104,N_8276);
nand U15284 (N_15284,N_8032,N_10310);
and U15285 (N_15285,N_8396,N_9823);
and U15286 (N_15286,N_11622,N_8732);
and U15287 (N_15287,N_10063,N_10152);
and U15288 (N_15288,N_11278,N_11243);
or U15289 (N_15289,N_10359,N_9390);
and U15290 (N_15290,N_8378,N_11955);
nor U15291 (N_15291,N_8512,N_8521);
nor U15292 (N_15292,N_10444,N_11401);
or U15293 (N_15293,N_8048,N_8976);
nor U15294 (N_15294,N_11558,N_10707);
nor U15295 (N_15295,N_10638,N_8789);
or U15296 (N_15296,N_11417,N_9416);
nand U15297 (N_15297,N_8661,N_8816);
nor U15298 (N_15298,N_8371,N_11890);
nand U15299 (N_15299,N_10016,N_9135);
nor U15300 (N_15300,N_9813,N_8044);
and U15301 (N_15301,N_11377,N_10034);
and U15302 (N_15302,N_10725,N_10377);
and U15303 (N_15303,N_10934,N_10079);
or U15304 (N_15304,N_9264,N_9144);
nor U15305 (N_15305,N_11032,N_8128);
or U15306 (N_15306,N_10494,N_10211);
nand U15307 (N_15307,N_10621,N_10913);
and U15308 (N_15308,N_11956,N_8930);
and U15309 (N_15309,N_10979,N_10453);
nand U15310 (N_15310,N_8458,N_11362);
nand U15311 (N_15311,N_10063,N_8212);
or U15312 (N_15312,N_10777,N_10679);
and U15313 (N_15313,N_10934,N_8463);
or U15314 (N_15314,N_11210,N_10381);
and U15315 (N_15315,N_11417,N_9972);
nand U15316 (N_15316,N_10894,N_10054);
or U15317 (N_15317,N_11734,N_8742);
nor U15318 (N_15318,N_8057,N_9250);
nor U15319 (N_15319,N_9098,N_11502);
or U15320 (N_15320,N_10549,N_9944);
and U15321 (N_15321,N_11211,N_8361);
or U15322 (N_15322,N_9397,N_10798);
or U15323 (N_15323,N_11599,N_9086);
nand U15324 (N_15324,N_8822,N_11685);
nand U15325 (N_15325,N_9609,N_8683);
or U15326 (N_15326,N_11525,N_8206);
nand U15327 (N_15327,N_10441,N_11054);
or U15328 (N_15328,N_9321,N_10972);
and U15329 (N_15329,N_11961,N_11714);
or U15330 (N_15330,N_8039,N_11624);
nand U15331 (N_15331,N_8085,N_10101);
nand U15332 (N_15332,N_11203,N_9644);
nand U15333 (N_15333,N_10148,N_11680);
or U15334 (N_15334,N_8865,N_11836);
or U15335 (N_15335,N_9169,N_10530);
nand U15336 (N_15336,N_9905,N_11980);
nor U15337 (N_15337,N_8559,N_8017);
nand U15338 (N_15338,N_10105,N_9748);
or U15339 (N_15339,N_10731,N_8607);
nor U15340 (N_15340,N_11962,N_8479);
and U15341 (N_15341,N_8969,N_11123);
and U15342 (N_15342,N_11028,N_11668);
nand U15343 (N_15343,N_8721,N_8636);
nor U15344 (N_15344,N_8954,N_11452);
and U15345 (N_15345,N_8104,N_8524);
nand U15346 (N_15346,N_10545,N_11175);
nand U15347 (N_15347,N_11482,N_9903);
or U15348 (N_15348,N_11426,N_9955);
and U15349 (N_15349,N_11115,N_8622);
and U15350 (N_15350,N_10309,N_10563);
nor U15351 (N_15351,N_11990,N_8702);
nor U15352 (N_15352,N_8881,N_11640);
xor U15353 (N_15353,N_8955,N_9926);
or U15354 (N_15354,N_8822,N_11745);
nand U15355 (N_15355,N_8544,N_10200);
and U15356 (N_15356,N_8168,N_8227);
or U15357 (N_15357,N_8793,N_11787);
and U15358 (N_15358,N_9642,N_8282);
and U15359 (N_15359,N_11399,N_10513);
or U15360 (N_15360,N_10676,N_9656);
or U15361 (N_15361,N_9152,N_9499);
nand U15362 (N_15362,N_10222,N_9156);
nand U15363 (N_15363,N_10020,N_9135);
and U15364 (N_15364,N_11668,N_10181);
or U15365 (N_15365,N_11018,N_9122);
and U15366 (N_15366,N_9507,N_10130);
nand U15367 (N_15367,N_11309,N_9821);
and U15368 (N_15368,N_10885,N_9433);
nor U15369 (N_15369,N_8854,N_10557);
nor U15370 (N_15370,N_11327,N_8772);
and U15371 (N_15371,N_8541,N_10747);
nor U15372 (N_15372,N_8495,N_10124);
nand U15373 (N_15373,N_9906,N_10407);
and U15374 (N_15374,N_11328,N_9940);
or U15375 (N_15375,N_11874,N_11410);
or U15376 (N_15376,N_8661,N_11919);
or U15377 (N_15377,N_8096,N_10436);
nand U15378 (N_15378,N_11666,N_9892);
and U15379 (N_15379,N_11161,N_11239);
or U15380 (N_15380,N_9188,N_8512);
nor U15381 (N_15381,N_10724,N_10388);
or U15382 (N_15382,N_11782,N_9188);
nand U15383 (N_15383,N_8162,N_10623);
or U15384 (N_15384,N_10640,N_8083);
and U15385 (N_15385,N_11300,N_8071);
nand U15386 (N_15386,N_11540,N_10473);
or U15387 (N_15387,N_10476,N_8137);
nand U15388 (N_15388,N_9669,N_10736);
or U15389 (N_15389,N_10848,N_9825);
xnor U15390 (N_15390,N_10023,N_8131);
or U15391 (N_15391,N_11863,N_10559);
nand U15392 (N_15392,N_11161,N_10664);
or U15393 (N_15393,N_11417,N_9328);
and U15394 (N_15394,N_10950,N_10501);
or U15395 (N_15395,N_8594,N_8206);
nand U15396 (N_15396,N_11451,N_10652);
and U15397 (N_15397,N_10666,N_10682);
or U15398 (N_15398,N_11063,N_8113);
and U15399 (N_15399,N_11152,N_10560);
nor U15400 (N_15400,N_11041,N_9879);
nor U15401 (N_15401,N_11337,N_10132);
nand U15402 (N_15402,N_10996,N_11171);
and U15403 (N_15403,N_10746,N_8838);
nand U15404 (N_15404,N_10910,N_11921);
nor U15405 (N_15405,N_10315,N_9121);
nor U15406 (N_15406,N_10480,N_9021);
nand U15407 (N_15407,N_8719,N_9194);
nor U15408 (N_15408,N_9681,N_8133);
or U15409 (N_15409,N_11492,N_8947);
or U15410 (N_15410,N_9248,N_10974);
and U15411 (N_15411,N_9686,N_9843);
or U15412 (N_15412,N_8535,N_9228);
and U15413 (N_15413,N_11668,N_10464);
or U15414 (N_15414,N_9059,N_11199);
xor U15415 (N_15415,N_10739,N_9646);
nand U15416 (N_15416,N_10843,N_8418);
or U15417 (N_15417,N_11941,N_11031);
xor U15418 (N_15418,N_11726,N_9892);
nand U15419 (N_15419,N_9609,N_9743);
and U15420 (N_15420,N_10713,N_8415);
nand U15421 (N_15421,N_10238,N_9469);
or U15422 (N_15422,N_8027,N_11660);
nand U15423 (N_15423,N_11505,N_10277);
or U15424 (N_15424,N_8792,N_11197);
nand U15425 (N_15425,N_10142,N_11706);
nor U15426 (N_15426,N_10694,N_11132);
nand U15427 (N_15427,N_10675,N_8944);
nand U15428 (N_15428,N_11241,N_8103);
nand U15429 (N_15429,N_11599,N_11048);
or U15430 (N_15430,N_9782,N_11315);
and U15431 (N_15431,N_11214,N_10514);
nand U15432 (N_15432,N_10231,N_10650);
nor U15433 (N_15433,N_10073,N_9638);
nor U15434 (N_15434,N_10018,N_11253);
nand U15435 (N_15435,N_10304,N_8511);
nor U15436 (N_15436,N_10923,N_11073);
and U15437 (N_15437,N_9843,N_9122);
and U15438 (N_15438,N_11740,N_10176);
nor U15439 (N_15439,N_10510,N_9008);
or U15440 (N_15440,N_9252,N_9618);
and U15441 (N_15441,N_10822,N_8453);
and U15442 (N_15442,N_8593,N_9859);
or U15443 (N_15443,N_11042,N_9629);
nand U15444 (N_15444,N_10377,N_11327);
or U15445 (N_15445,N_10719,N_11216);
xor U15446 (N_15446,N_11317,N_8321);
nand U15447 (N_15447,N_8257,N_11079);
xor U15448 (N_15448,N_11617,N_11857);
nor U15449 (N_15449,N_11115,N_9945);
or U15450 (N_15450,N_11340,N_8636);
nand U15451 (N_15451,N_10647,N_9250);
nand U15452 (N_15452,N_8920,N_10285);
nor U15453 (N_15453,N_9705,N_8240);
nor U15454 (N_15454,N_10769,N_11162);
or U15455 (N_15455,N_8119,N_8775);
or U15456 (N_15456,N_10573,N_11762);
nand U15457 (N_15457,N_11127,N_10427);
nand U15458 (N_15458,N_8533,N_9874);
or U15459 (N_15459,N_11907,N_10516);
or U15460 (N_15460,N_11636,N_9365);
or U15461 (N_15461,N_10172,N_9998);
or U15462 (N_15462,N_11970,N_8128);
or U15463 (N_15463,N_9795,N_8638);
nand U15464 (N_15464,N_10114,N_10889);
or U15465 (N_15465,N_8870,N_11003);
nor U15466 (N_15466,N_9111,N_10901);
nand U15467 (N_15467,N_8542,N_9759);
nand U15468 (N_15468,N_8166,N_9343);
and U15469 (N_15469,N_9128,N_10974);
nand U15470 (N_15470,N_11040,N_11221);
or U15471 (N_15471,N_11351,N_10995);
and U15472 (N_15472,N_8163,N_11302);
nor U15473 (N_15473,N_8284,N_10638);
nand U15474 (N_15474,N_10746,N_11127);
nor U15475 (N_15475,N_10524,N_10791);
nand U15476 (N_15476,N_9342,N_8203);
nor U15477 (N_15477,N_11057,N_8162);
and U15478 (N_15478,N_8064,N_9070);
and U15479 (N_15479,N_8529,N_8609);
nand U15480 (N_15480,N_9045,N_11976);
and U15481 (N_15481,N_9751,N_9417);
nand U15482 (N_15482,N_10614,N_11404);
nand U15483 (N_15483,N_9492,N_10801);
xor U15484 (N_15484,N_11695,N_9519);
and U15485 (N_15485,N_11199,N_9713);
nand U15486 (N_15486,N_9094,N_9030);
or U15487 (N_15487,N_11100,N_10737);
nor U15488 (N_15488,N_10680,N_11982);
nor U15489 (N_15489,N_8818,N_8213);
and U15490 (N_15490,N_10969,N_10871);
and U15491 (N_15491,N_9705,N_10117);
or U15492 (N_15492,N_11398,N_9153);
nor U15493 (N_15493,N_8960,N_11528);
nand U15494 (N_15494,N_10761,N_9953);
nand U15495 (N_15495,N_10540,N_9143);
nand U15496 (N_15496,N_8772,N_8802);
or U15497 (N_15497,N_9363,N_10194);
nand U15498 (N_15498,N_11368,N_9736);
nand U15499 (N_15499,N_10498,N_10215);
and U15500 (N_15500,N_9499,N_11210);
nor U15501 (N_15501,N_8312,N_9386);
and U15502 (N_15502,N_11809,N_8268);
and U15503 (N_15503,N_9529,N_11493);
nand U15504 (N_15504,N_9680,N_10427);
nand U15505 (N_15505,N_11363,N_9321);
and U15506 (N_15506,N_8444,N_11094);
or U15507 (N_15507,N_8802,N_10619);
and U15508 (N_15508,N_8631,N_11250);
and U15509 (N_15509,N_11859,N_9924);
and U15510 (N_15510,N_8883,N_9890);
or U15511 (N_15511,N_9508,N_9040);
nand U15512 (N_15512,N_8797,N_9689);
nand U15513 (N_15513,N_8178,N_10327);
and U15514 (N_15514,N_10141,N_9130);
nor U15515 (N_15515,N_11814,N_9416);
nor U15516 (N_15516,N_9522,N_10393);
and U15517 (N_15517,N_10160,N_9007);
nand U15518 (N_15518,N_11353,N_10826);
and U15519 (N_15519,N_8905,N_10746);
and U15520 (N_15520,N_10240,N_8810);
or U15521 (N_15521,N_11969,N_11260);
nor U15522 (N_15522,N_8726,N_9106);
or U15523 (N_15523,N_9578,N_8216);
nor U15524 (N_15524,N_8922,N_8342);
nand U15525 (N_15525,N_9173,N_8827);
nor U15526 (N_15526,N_10498,N_11270);
nand U15527 (N_15527,N_11485,N_11424);
nand U15528 (N_15528,N_8746,N_10793);
and U15529 (N_15529,N_8823,N_9139);
or U15530 (N_15530,N_9755,N_11847);
nand U15531 (N_15531,N_10381,N_10148);
or U15532 (N_15532,N_10330,N_9941);
xor U15533 (N_15533,N_10807,N_11658);
and U15534 (N_15534,N_8757,N_8371);
nand U15535 (N_15535,N_9053,N_11705);
or U15536 (N_15536,N_10372,N_9248);
nor U15537 (N_15537,N_9728,N_9532);
or U15538 (N_15538,N_8712,N_11379);
nand U15539 (N_15539,N_9464,N_10643);
nor U15540 (N_15540,N_8005,N_8139);
or U15541 (N_15541,N_11176,N_10334);
nand U15542 (N_15542,N_10323,N_11256);
nand U15543 (N_15543,N_10631,N_8386);
and U15544 (N_15544,N_11988,N_8487);
nand U15545 (N_15545,N_10505,N_8659);
nor U15546 (N_15546,N_9998,N_9091);
and U15547 (N_15547,N_8059,N_9990);
nand U15548 (N_15548,N_11842,N_11392);
nand U15549 (N_15549,N_9084,N_9895);
nand U15550 (N_15550,N_8405,N_8411);
and U15551 (N_15551,N_11920,N_9640);
and U15552 (N_15552,N_8167,N_11791);
or U15553 (N_15553,N_8820,N_11100);
and U15554 (N_15554,N_9258,N_11035);
nor U15555 (N_15555,N_10871,N_9429);
or U15556 (N_15556,N_9856,N_10560);
nand U15557 (N_15557,N_8351,N_10569);
or U15558 (N_15558,N_11001,N_10746);
nor U15559 (N_15559,N_11327,N_10401);
nand U15560 (N_15560,N_8562,N_8375);
nand U15561 (N_15561,N_11799,N_9837);
nand U15562 (N_15562,N_9747,N_11343);
nor U15563 (N_15563,N_9120,N_11307);
nor U15564 (N_15564,N_11245,N_9356);
or U15565 (N_15565,N_11883,N_10889);
and U15566 (N_15566,N_10071,N_11000);
nor U15567 (N_15567,N_10038,N_8782);
nor U15568 (N_15568,N_10571,N_9610);
or U15569 (N_15569,N_10286,N_8737);
nand U15570 (N_15570,N_8834,N_10289);
and U15571 (N_15571,N_9645,N_10495);
and U15572 (N_15572,N_11406,N_8585);
or U15573 (N_15573,N_8281,N_8630);
and U15574 (N_15574,N_10087,N_8986);
and U15575 (N_15575,N_11287,N_9243);
or U15576 (N_15576,N_8907,N_9825);
nor U15577 (N_15577,N_8529,N_9059);
or U15578 (N_15578,N_10829,N_10646);
and U15579 (N_15579,N_11357,N_10271);
nand U15580 (N_15580,N_9810,N_10844);
nor U15581 (N_15581,N_11738,N_10820);
and U15582 (N_15582,N_8414,N_10578);
or U15583 (N_15583,N_11282,N_10246);
nand U15584 (N_15584,N_9388,N_10537);
and U15585 (N_15585,N_9339,N_8065);
nor U15586 (N_15586,N_11973,N_11487);
nand U15587 (N_15587,N_8445,N_11626);
nand U15588 (N_15588,N_8874,N_10534);
nor U15589 (N_15589,N_8817,N_10361);
nand U15590 (N_15590,N_9200,N_9788);
and U15591 (N_15591,N_8674,N_11371);
or U15592 (N_15592,N_9690,N_8035);
nand U15593 (N_15593,N_11285,N_9953);
or U15594 (N_15594,N_10988,N_10301);
and U15595 (N_15595,N_10719,N_10007);
nor U15596 (N_15596,N_10328,N_8803);
or U15597 (N_15597,N_9903,N_8933);
and U15598 (N_15598,N_8055,N_9501);
nor U15599 (N_15599,N_10994,N_11510);
nor U15600 (N_15600,N_10891,N_11419);
and U15601 (N_15601,N_11232,N_9173);
and U15602 (N_15602,N_11827,N_11257);
or U15603 (N_15603,N_8618,N_9009);
nor U15604 (N_15604,N_11908,N_8797);
nand U15605 (N_15605,N_9682,N_11181);
and U15606 (N_15606,N_11653,N_11730);
nor U15607 (N_15607,N_8866,N_10828);
nor U15608 (N_15608,N_11239,N_8240);
nor U15609 (N_15609,N_10235,N_9777);
and U15610 (N_15610,N_8396,N_10856);
or U15611 (N_15611,N_10374,N_10989);
nand U15612 (N_15612,N_9827,N_11770);
nor U15613 (N_15613,N_9878,N_8260);
nor U15614 (N_15614,N_8254,N_8180);
nand U15615 (N_15615,N_11242,N_8866);
and U15616 (N_15616,N_8015,N_8018);
or U15617 (N_15617,N_11572,N_11972);
or U15618 (N_15618,N_8032,N_9057);
or U15619 (N_15619,N_10912,N_9569);
nor U15620 (N_15620,N_11725,N_9996);
and U15621 (N_15621,N_10401,N_11369);
nand U15622 (N_15622,N_9867,N_8602);
nor U15623 (N_15623,N_10766,N_9411);
nand U15624 (N_15624,N_10535,N_11219);
nand U15625 (N_15625,N_11479,N_11350);
nand U15626 (N_15626,N_8266,N_10968);
nor U15627 (N_15627,N_10007,N_11150);
nand U15628 (N_15628,N_8081,N_8768);
or U15629 (N_15629,N_9422,N_11794);
nand U15630 (N_15630,N_10973,N_9623);
nor U15631 (N_15631,N_8000,N_8190);
or U15632 (N_15632,N_10372,N_10189);
nor U15633 (N_15633,N_8113,N_8639);
or U15634 (N_15634,N_11267,N_11460);
or U15635 (N_15635,N_8244,N_10007);
or U15636 (N_15636,N_10625,N_9394);
or U15637 (N_15637,N_8838,N_11707);
or U15638 (N_15638,N_9096,N_10386);
nand U15639 (N_15639,N_9576,N_11019);
and U15640 (N_15640,N_8120,N_10300);
nand U15641 (N_15641,N_11179,N_8443);
or U15642 (N_15642,N_11715,N_9168);
nor U15643 (N_15643,N_11661,N_8128);
nand U15644 (N_15644,N_11343,N_11210);
or U15645 (N_15645,N_11384,N_9450);
nor U15646 (N_15646,N_8788,N_11077);
nand U15647 (N_15647,N_8562,N_10540);
or U15648 (N_15648,N_10978,N_8917);
nand U15649 (N_15649,N_10030,N_11680);
nand U15650 (N_15650,N_8269,N_10025);
nand U15651 (N_15651,N_9346,N_8345);
and U15652 (N_15652,N_10261,N_11970);
nor U15653 (N_15653,N_10244,N_10427);
or U15654 (N_15654,N_10432,N_8049);
or U15655 (N_15655,N_10108,N_9735);
and U15656 (N_15656,N_9886,N_11241);
or U15657 (N_15657,N_11684,N_8209);
or U15658 (N_15658,N_10503,N_11956);
nand U15659 (N_15659,N_8664,N_10786);
or U15660 (N_15660,N_11092,N_8148);
nor U15661 (N_15661,N_10883,N_10777);
or U15662 (N_15662,N_9404,N_8904);
or U15663 (N_15663,N_9464,N_8462);
and U15664 (N_15664,N_8655,N_8322);
or U15665 (N_15665,N_9610,N_10439);
nor U15666 (N_15666,N_10252,N_11785);
nor U15667 (N_15667,N_10767,N_10699);
or U15668 (N_15668,N_10156,N_10678);
nand U15669 (N_15669,N_9966,N_10399);
and U15670 (N_15670,N_9937,N_8145);
or U15671 (N_15671,N_10811,N_11066);
or U15672 (N_15672,N_9271,N_11318);
and U15673 (N_15673,N_11832,N_11745);
nor U15674 (N_15674,N_10079,N_9067);
and U15675 (N_15675,N_11329,N_9888);
or U15676 (N_15676,N_8405,N_11935);
or U15677 (N_15677,N_9854,N_10740);
nand U15678 (N_15678,N_8749,N_9115);
nor U15679 (N_15679,N_10789,N_11058);
or U15680 (N_15680,N_8792,N_9864);
nand U15681 (N_15681,N_10013,N_10673);
or U15682 (N_15682,N_8600,N_9290);
nand U15683 (N_15683,N_11808,N_9245);
nor U15684 (N_15684,N_10840,N_9090);
nor U15685 (N_15685,N_11239,N_9600);
nand U15686 (N_15686,N_9561,N_10042);
nor U15687 (N_15687,N_8071,N_9741);
nor U15688 (N_15688,N_10367,N_11156);
nor U15689 (N_15689,N_9408,N_8805);
or U15690 (N_15690,N_9841,N_10722);
or U15691 (N_15691,N_10930,N_10622);
nand U15692 (N_15692,N_10197,N_9689);
and U15693 (N_15693,N_9646,N_10190);
nand U15694 (N_15694,N_10940,N_11003);
or U15695 (N_15695,N_11886,N_9543);
and U15696 (N_15696,N_9056,N_9971);
xor U15697 (N_15697,N_11428,N_10637);
or U15698 (N_15698,N_11815,N_10155);
and U15699 (N_15699,N_8881,N_11992);
nand U15700 (N_15700,N_8102,N_8378);
or U15701 (N_15701,N_8756,N_9009);
nor U15702 (N_15702,N_10877,N_11468);
nand U15703 (N_15703,N_9726,N_11527);
or U15704 (N_15704,N_11409,N_9183);
nor U15705 (N_15705,N_11814,N_8234);
or U15706 (N_15706,N_10624,N_10144);
nor U15707 (N_15707,N_11909,N_8994);
and U15708 (N_15708,N_9018,N_8496);
and U15709 (N_15709,N_8064,N_9108);
nor U15710 (N_15710,N_11114,N_8319);
nor U15711 (N_15711,N_8034,N_10582);
or U15712 (N_15712,N_9749,N_8391);
nor U15713 (N_15713,N_9649,N_9152);
nand U15714 (N_15714,N_9948,N_9365);
xnor U15715 (N_15715,N_11851,N_11412);
or U15716 (N_15716,N_10766,N_9901);
or U15717 (N_15717,N_11180,N_9575);
nor U15718 (N_15718,N_10830,N_11036);
or U15719 (N_15719,N_11539,N_11222);
nand U15720 (N_15720,N_9826,N_9799);
and U15721 (N_15721,N_10542,N_9704);
nand U15722 (N_15722,N_11312,N_11555);
nor U15723 (N_15723,N_8475,N_9262);
nor U15724 (N_15724,N_11278,N_8956);
nand U15725 (N_15725,N_11817,N_10027);
and U15726 (N_15726,N_10567,N_8993);
nor U15727 (N_15727,N_11225,N_10284);
nand U15728 (N_15728,N_10276,N_10521);
nand U15729 (N_15729,N_11339,N_9687);
nand U15730 (N_15730,N_9799,N_9860);
nor U15731 (N_15731,N_9242,N_9485);
and U15732 (N_15732,N_9676,N_11525);
or U15733 (N_15733,N_10580,N_10231);
nand U15734 (N_15734,N_9673,N_11187);
nor U15735 (N_15735,N_8748,N_9896);
nor U15736 (N_15736,N_9011,N_11553);
or U15737 (N_15737,N_8825,N_11821);
or U15738 (N_15738,N_9643,N_8476);
nor U15739 (N_15739,N_8410,N_9789);
nand U15740 (N_15740,N_9735,N_9708);
or U15741 (N_15741,N_9202,N_8582);
or U15742 (N_15742,N_11287,N_11864);
nor U15743 (N_15743,N_11356,N_8042);
or U15744 (N_15744,N_10877,N_10330);
nor U15745 (N_15745,N_9919,N_9154);
or U15746 (N_15746,N_9862,N_11037);
nand U15747 (N_15747,N_11916,N_10803);
and U15748 (N_15748,N_8663,N_9497);
nand U15749 (N_15749,N_8612,N_8708);
nor U15750 (N_15750,N_11800,N_8534);
or U15751 (N_15751,N_9843,N_8946);
nand U15752 (N_15752,N_10182,N_11219);
or U15753 (N_15753,N_10991,N_8121);
nor U15754 (N_15754,N_10654,N_9590);
and U15755 (N_15755,N_8320,N_8373);
nor U15756 (N_15756,N_11782,N_10232);
nor U15757 (N_15757,N_10859,N_9731);
nand U15758 (N_15758,N_9803,N_8576);
nand U15759 (N_15759,N_10808,N_8988);
nor U15760 (N_15760,N_11089,N_10218);
or U15761 (N_15761,N_8848,N_9793);
nor U15762 (N_15762,N_8021,N_11406);
or U15763 (N_15763,N_9320,N_11137);
nand U15764 (N_15764,N_8557,N_9891);
or U15765 (N_15765,N_9116,N_9423);
and U15766 (N_15766,N_8630,N_9199);
and U15767 (N_15767,N_9186,N_9352);
or U15768 (N_15768,N_10953,N_11619);
or U15769 (N_15769,N_9469,N_11070);
nand U15770 (N_15770,N_11234,N_11383);
nand U15771 (N_15771,N_10279,N_10348);
nand U15772 (N_15772,N_9425,N_9091);
nand U15773 (N_15773,N_10400,N_8028);
nor U15774 (N_15774,N_11394,N_8702);
or U15775 (N_15775,N_8901,N_9300);
nand U15776 (N_15776,N_8435,N_10197);
nand U15777 (N_15777,N_8364,N_9549);
and U15778 (N_15778,N_10805,N_8654);
and U15779 (N_15779,N_10405,N_11730);
nand U15780 (N_15780,N_10559,N_9354);
or U15781 (N_15781,N_10880,N_11335);
and U15782 (N_15782,N_9395,N_8329);
and U15783 (N_15783,N_8848,N_11646);
and U15784 (N_15784,N_11876,N_9787);
nand U15785 (N_15785,N_9276,N_10521);
or U15786 (N_15786,N_10058,N_10203);
and U15787 (N_15787,N_10032,N_10063);
and U15788 (N_15788,N_10951,N_9658);
nor U15789 (N_15789,N_11095,N_10397);
and U15790 (N_15790,N_11845,N_11266);
nor U15791 (N_15791,N_11528,N_11084);
and U15792 (N_15792,N_8685,N_11596);
nand U15793 (N_15793,N_10231,N_9673);
nand U15794 (N_15794,N_11195,N_9720);
nor U15795 (N_15795,N_10732,N_11602);
or U15796 (N_15796,N_8766,N_8599);
or U15797 (N_15797,N_8231,N_8237);
and U15798 (N_15798,N_10362,N_11082);
nand U15799 (N_15799,N_8606,N_8656);
nand U15800 (N_15800,N_10956,N_8721);
nand U15801 (N_15801,N_10067,N_10441);
or U15802 (N_15802,N_8182,N_8654);
and U15803 (N_15803,N_8679,N_11576);
or U15804 (N_15804,N_9966,N_10184);
and U15805 (N_15805,N_10108,N_11963);
and U15806 (N_15806,N_11846,N_11325);
nor U15807 (N_15807,N_8877,N_9926);
nand U15808 (N_15808,N_8330,N_8241);
nand U15809 (N_15809,N_8698,N_9373);
nand U15810 (N_15810,N_9258,N_11583);
or U15811 (N_15811,N_10990,N_8825);
nor U15812 (N_15812,N_11837,N_11442);
nor U15813 (N_15813,N_9799,N_10249);
and U15814 (N_15814,N_11962,N_8017);
or U15815 (N_15815,N_10990,N_11882);
or U15816 (N_15816,N_9559,N_10839);
and U15817 (N_15817,N_8516,N_8282);
or U15818 (N_15818,N_11705,N_10713);
and U15819 (N_15819,N_9097,N_11057);
and U15820 (N_15820,N_9598,N_8637);
nor U15821 (N_15821,N_9927,N_11790);
nand U15822 (N_15822,N_8838,N_10661);
nand U15823 (N_15823,N_11222,N_8686);
nand U15824 (N_15824,N_11429,N_9912);
and U15825 (N_15825,N_10950,N_8417);
nand U15826 (N_15826,N_8223,N_10363);
and U15827 (N_15827,N_10445,N_11602);
nand U15828 (N_15828,N_9499,N_8246);
nand U15829 (N_15829,N_11370,N_9628);
nor U15830 (N_15830,N_9053,N_11944);
nand U15831 (N_15831,N_10392,N_10223);
nor U15832 (N_15832,N_8524,N_11362);
nand U15833 (N_15833,N_8449,N_10835);
and U15834 (N_15834,N_8361,N_10109);
xor U15835 (N_15835,N_11832,N_9604);
nand U15836 (N_15836,N_9449,N_8207);
and U15837 (N_15837,N_9848,N_11353);
or U15838 (N_15838,N_10321,N_9992);
nand U15839 (N_15839,N_9798,N_11651);
nand U15840 (N_15840,N_11639,N_9011);
nand U15841 (N_15841,N_9215,N_9820);
or U15842 (N_15842,N_8396,N_8141);
nor U15843 (N_15843,N_9992,N_9267);
and U15844 (N_15844,N_10297,N_9100);
and U15845 (N_15845,N_11465,N_10294);
and U15846 (N_15846,N_9951,N_10782);
and U15847 (N_15847,N_10826,N_8392);
nand U15848 (N_15848,N_11249,N_9603);
and U15849 (N_15849,N_9657,N_8080);
nand U15850 (N_15850,N_10551,N_8644);
nand U15851 (N_15851,N_8404,N_11326);
or U15852 (N_15852,N_9090,N_10589);
nand U15853 (N_15853,N_9409,N_10819);
nor U15854 (N_15854,N_10315,N_11960);
or U15855 (N_15855,N_10487,N_9081);
nor U15856 (N_15856,N_11075,N_9861);
and U15857 (N_15857,N_8025,N_8863);
nor U15858 (N_15858,N_11115,N_10254);
or U15859 (N_15859,N_9495,N_11971);
nand U15860 (N_15860,N_9902,N_9503);
nand U15861 (N_15861,N_11114,N_9513);
nor U15862 (N_15862,N_9069,N_10185);
nor U15863 (N_15863,N_11910,N_10851);
nor U15864 (N_15864,N_10210,N_11784);
nor U15865 (N_15865,N_9456,N_9477);
nor U15866 (N_15866,N_8423,N_11811);
nor U15867 (N_15867,N_8615,N_11490);
or U15868 (N_15868,N_10866,N_8572);
nor U15869 (N_15869,N_10105,N_8782);
or U15870 (N_15870,N_11093,N_10009);
nand U15871 (N_15871,N_8095,N_11682);
nor U15872 (N_15872,N_11687,N_8312);
nor U15873 (N_15873,N_10425,N_10830);
or U15874 (N_15874,N_11221,N_11274);
or U15875 (N_15875,N_11733,N_10792);
or U15876 (N_15876,N_9783,N_11400);
and U15877 (N_15877,N_11609,N_10862);
or U15878 (N_15878,N_8415,N_10172);
and U15879 (N_15879,N_9174,N_9300);
or U15880 (N_15880,N_8408,N_8370);
or U15881 (N_15881,N_11659,N_11700);
nand U15882 (N_15882,N_9550,N_8264);
nand U15883 (N_15883,N_10619,N_8583);
nand U15884 (N_15884,N_8018,N_10997);
and U15885 (N_15885,N_8051,N_8318);
or U15886 (N_15886,N_10981,N_11409);
nand U15887 (N_15887,N_9761,N_10237);
nor U15888 (N_15888,N_9425,N_8368);
nand U15889 (N_15889,N_10841,N_11182);
and U15890 (N_15890,N_11850,N_10134);
nand U15891 (N_15891,N_10872,N_9516);
and U15892 (N_15892,N_10258,N_11274);
or U15893 (N_15893,N_9773,N_8849);
and U15894 (N_15894,N_11102,N_8811);
or U15895 (N_15895,N_11271,N_8557);
and U15896 (N_15896,N_11314,N_11719);
and U15897 (N_15897,N_8531,N_8185);
nor U15898 (N_15898,N_10386,N_10734);
nand U15899 (N_15899,N_9444,N_10646);
nand U15900 (N_15900,N_9053,N_10504);
and U15901 (N_15901,N_10515,N_11005);
nand U15902 (N_15902,N_10940,N_9358);
nor U15903 (N_15903,N_10993,N_9002);
nand U15904 (N_15904,N_11835,N_8255);
and U15905 (N_15905,N_9565,N_11109);
or U15906 (N_15906,N_11912,N_11984);
and U15907 (N_15907,N_11145,N_10944);
or U15908 (N_15908,N_8865,N_8151);
or U15909 (N_15909,N_11045,N_8545);
nand U15910 (N_15910,N_10248,N_9484);
nor U15911 (N_15911,N_9149,N_9046);
and U15912 (N_15912,N_11384,N_11208);
nor U15913 (N_15913,N_9766,N_8746);
nor U15914 (N_15914,N_11376,N_11282);
nor U15915 (N_15915,N_8257,N_9747);
or U15916 (N_15916,N_8896,N_10729);
nor U15917 (N_15917,N_9570,N_11192);
nand U15918 (N_15918,N_8954,N_8540);
nand U15919 (N_15919,N_9469,N_8051);
nor U15920 (N_15920,N_11841,N_9201);
or U15921 (N_15921,N_8785,N_9621);
nor U15922 (N_15922,N_10239,N_11101);
and U15923 (N_15923,N_10018,N_10374);
or U15924 (N_15924,N_8826,N_9423);
nand U15925 (N_15925,N_8917,N_11489);
and U15926 (N_15926,N_9427,N_9726);
nor U15927 (N_15927,N_11476,N_9287);
nand U15928 (N_15928,N_8998,N_11301);
nand U15929 (N_15929,N_8552,N_9019);
nor U15930 (N_15930,N_10142,N_11819);
nand U15931 (N_15931,N_9789,N_8322);
nor U15932 (N_15932,N_10956,N_9401);
or U15933 (N_15933,N_9431,N_11259);
nor U15934 (N_15934,N_9278,N_8453);
and U15935 (N_15935,N_8723,N_9528);
nor U15936 (N_15936,N_10811,N_10915);
or U15937 (N_15937,N_11957,N_9673);
or U15938 (N_15938,N_8033,N_8985);
or U15939 (N_15939,N_11082,N_11940);
nor U15940 (N_15940,N_10915,N_11359);
or U15941 (N_15941,N_10984,N_8725);
nand U15942 (N_15942,N_9473,N_10813);
xnor U15943 (N_15943,N_9311,N_11791);
nor U15944 (N_15944,N_8361,N_8518);
and U15945 (N_15945,N_10829,N_8823);
xnor U15946 (N_15946,N_11658,N_8973);
nand U15947 (N_15947,N_8986,N_11480);
nor U15948 (N_15948,N_10345,N_9263);
and U15949 (N_15949,N_11742,N_9182);
nand U15950 (N_15950,N_10242,N_11861);
nand U15951 (N_15951,N_9238,N_8369);
and U15952 (N_15952,N_8894,N_9386);
or U15953 (N_15953,N_8952,N_9568);
and U15954 (N_15954,N_8294,N_9726);
and U15955 (N_15955,N_9645,N_9599);
or U15956 (N_15956,N_10107,N_10176);
nor U15957 (N_15957,N_8528,N_11927);
nand U15958 (N_15958,N_10625,N_10225);
nor U15959 (N_15959,N_8486,N_11865);
nand U15960 (N_15960,N_8208,N_8110);
nand U15961 (N_15961,N_9762,N_11598);
nand U15962 (N_15962,N_8140,N_11016);
and U15963 (N_15963,N_10502,N_9809);
nor U15964 (N_15964,N_10939,N_10212);
or U15965 (N_15965,N_10077,N_10394);
nor U15966 (N_15966,N_8393,N_11147);
or U15967 (N_15967,N_11203,N_11125);
nand U15968 (N_15968,N_10687,N_10385);
or U15969 (N_15969,N_11829,N_11903);
nand U15970 (N_15970,N_11830,N_10509);
and U15971 (N_15971,N_10469,N_8140);
and U15972 (N_15972,N_11149,N_8920);
or U15973 (N_15973,N_9458,N_9426);
nand U15974 (N_15974,N_9679,N_11872);
and U15975 (N_15975,N_8301,N_8224);
nand U15976 (N_15976,N_11218,N_10837);
nor U15977 (N_15977,N_11890,N_8133);
xnor U15978 (N_15978,N_9897,N_11560);
or U15979 (N_15979,N_10310,N_11723);
or U15980 (N_15980,N_11485,N_8473);
or U15981 (N_15981,N_10359,N_11000);
nand U15982 (N_15982,N_10103,N_10206);
or U15983 (N_15983,N_8069,N_9429);
and U15984 (N_15984,N_8671,N_10078);
and U15985 (N_15985,N_8409,N_9839);
nor U15986 (N_15986,N_9077,N_10295);
nand U15987 (N_15987,N_8777,N_8458);
and U15988 (N_15988,N_11443,N_11163);
nor U15989 (N_15989,N_10003,N_8687);
and U15990 (N_15990,N_8135,N_11849);
and U15991 (N_15991,N_11550,N_8814);
or U15992 (N_15992,N_8634,N_11856);
nor U15993 (N_15993,N_8730,N_9983);
nor U15994 (N_15994,N_11246,N_10580);
and U15995 (N_15995,N_10582,N_9441);
and U15996 (N_15996,N_8086,N_11608);
and U15997 (N_15997,N_8161,N_8185);
nor U15998 (N_15998,N_11514,N_11502);
nand U15999 (N_15999,N_11843,N_9450);
or U16000 (N_16000,N_14500,N_15009);
nand U16001 (N_16001,N_14064,N_15462);
or U16002 (N_16002,N_14712,N_12141);
nor U16003 (N_16003,N_15643,N_12800);
and U16004 (N_16004,N_14197,N_15568);
nand U16005 (N_16005,N_13676,N_12167);
nand U16006 (N_16006,N_13867,N_13420);
xor U16007 (N_16007,N_15631,N_14835);
nand U16008 (N_16008,N_15910,N_15639);
or U16009 (N_16009,N_13764,N_13616);
nand U16010 (N_16010,N_12654,N_13243);
and U16011 (N_16011,N_14677,N_12505);
nor U16012 (N_16012,N_12452,N_14971);
and U16013 (N_16013,N_12112,N_13060);
or U16014 (N_16014,N_15507,N_12570);
nand U16015 (N_16015,N_15021,N_14988);
nor U16016 (N_16016,N_14529,N_15946);
nor U16017 (N_16017,N_15618,N_15753);
or U16018 (N_16018,N_14515,N_12309);
or U16019 (N_16019,N_14323,N_15878);
nor U16020 (N_16020,N_13879,N_14125);
nand U16021 (N_16021,N_15525,N_15145);
xnor U16022 (N_16022,N_12757,N_14512);
or U16023 (N_16023,N_12753,N_14393);
and U16024 (N_16024,N_15258,N_14164);
or U16025 (N_16025,N_14796,N_14447);
nor U16026 (N_16026,N_15273,N_12731);
or U16027 (N_16027,N_13415,N_12154);
or U16028 (N_16028,N_12632,N_14918);
or U16029 (N_16029,N_12110,N_12701);
nand U16030 (N_16030,N_13461,N_15709);
and U16031 (N_16031,N_13891,N_15182);
or U16032 (N_16032,N_15126,N_14317);
or U16033 (N_16033,N_13050,N_14802);
or U16034 (N_16034,N_12558,N_12482);
or U16035 (N_16035,N_15896,N_14153);
and U16036 (N_16036,N_14487,N_13074);
and U16037 (N_16037,N_13794,N_14704);
or U16038 (N_16038,N_12267,N_12914);
nor U16039 (N_16039,N_13018,N_12774);
nor U16040 (N_16040,N_12605,N_12748);
nor U16041 (N_16041,N_12602,N_14110);
nand U16042 (N_16042,N_13257,N_13868);
xor U16043 (N_16043,N_13345,N_12087);
nor U16044 (N_16044,N_13985,N_14563);
nor U16045 (N_16045,N_14123,N_15841);
and U16046 (N_16046,N_14065,N_13184);
nor U16047 (N_16047,N_12035,N_15786);
nand U16048 (N_16048,N_12389,N_15201);
nor U16049 (N_16049,N_15606,N_13183);
nand U16050 (N_16050,N_13581,N_14538);
nor U16051 (N_16051,N_15204,N_13120);
nor U16052 (N_16052,N_15650,N_12916);
and U16053 (N_16053,N_14465,N_14265);
nor U16054 (N_16054,N_14302,N_13273);
and U16055 (N_16055,N_14630,N_14096);
or U16056 (N_16056,N_15808,N_13135);
nor U16057 (N_16057,N_14006,N_13466);
nor U16058 (N_16058,N_12079,N_12439);
and U16059 (N_16059,N_15607,N_15605);
nand U16060 (N_16060,N_15952,N_15647);
xor U16061 (N_16061,N_15084,N_15453);
nand U16062 (N_16062,N_13193,N_13195);
or U16063 (N_16063,N_12455,N_13075);
nand U16064 (N_16064,N_15397,N_15104);
nor U16065 (N_16065,N_15156,N_13815);
and U16066 (N_16066,N_14479,N_15064);
or U16067 (N_16067,N_15452,N_12320);
or U16068 (N_16068,N_12486,N_12226);
nand U16069 (N_16069,N_12624,N_15184);
or U16070 (N_16070,N_12064,N_15531);
nand U16071 (N_16071,N_13943,N_14685);
nand U16072 (N_16072,N_14762,N_15973);
nor U16073 (N_16073,N_12448,N_14594);
or U16074 (N_16074,N_15781,N_15333);
or U16075 (N_16075,N_15721,N_12495);
nor U16076 (N_16076,N_12750,N_14853);
nor U16077 (N_16077,N_13557,N_12433);
or U16078 (N_16078,N_12122,N_12722);
nand U16079 (N_16079,N_12123,N_14081);
nand U16080 (N_16080,N_15689,N_13423);
nor U16081 (N_16081,N_13539,N_12504);
nor U16082 (N_16082,N_12416,N_15746);
nand U16083 (N_16083,N_15839,N_15492);
nor U16084 (N_16084,N_14919,N_12712);
nor U16085 (N_16085,N_13725,N_15413);
nor U16086 (N_16086,N_13402,N_12521);
nand U16087 (N_16087,N_13928,N_13440);
and U16088 (N_16088,N_12596,N_15044);
and U16089 (N_16089,N_12865,N_13965);
or U16090 (N_16090,N_13459,N_14577);
and U16091 (N_16091,N_12590,N_12912);
nor U16092 (N_16092,N_13997,N_14368);
xnor U16093 (N_16093,N_12595,N_13613);
nand U16094 (N_16094,N_13651,N_13822);
and U16095 (N_16095,N_15293,N_13084);
nor U16096 (N_16096,N_14637,N_12686);
nor U16097 (N_16097,N_14751,N_12525);
nand U16098 (N_16098,N_15768,N_13190);
or U16099 (N_16099,N_15793,N_15642);
nor U16100 (N_16100,N_12084,N_12217);
or U16101 (N_16101,N_14388,N_13244);
nand U16102 (N_16102,N_12191,N_12446);
and U16103 (N_16103,N_13131,N_14733);
or U16104 (N_16104,N_15945,N_15949);
nand U16105 (N_16105,N_14203,N_14938);
nor U16106 (N_16106,N_14787,N_15058);
nor U16107 (N_16107,N_12833,N_15434);
nor U16108 (N_16108,N_14995,N_12435);
or U16109 (N_16109,N_13441,N_14216);
or U16110 (N_16110,N_14684,N_14230);
and U16111 (N_16111,N_15376,N_13372);
or U16112 (N_16112,N_15159,N_12434);
or U16113 (N_16113,N_13079,N_15911);
or U16114 (N_16114,N_13362,N_15623);
nor U16115 (N_16115,N_12432,N_12109);
nand U16116 (N_16116,N_13003,N_15033);
xnor U16117 (N_16117,N_15888,N_15707);
nand U16118 (N_16118,N_12113,N_15216);
or U16119 (N_16119,N_13721,N_13561);
nor U16120 (N_16120,N_12532,N_13984);
nor U16121 (N_16121,N_12585,N_14681);
or U16122 (N_16122,N_13795,N_14566);
nand U16123 (N_16123,N_12494,N_14463);
or U16124 (N_16124,N_15267,N_12421);
nand U16125 (N_16125,N_15343,N_14141);
and U16126 (N_16126,N_15890,N_13799);
and U16127 (N_16127,N_12149,N_13918);
nand U16128 (N_16128,N_13428,N_15597);
nand U16129 (N_16129,N_13233,N_12045);
and U16130 (N_16130,N_12888,N_13356);
and U16131 (N_16131,N_15116,N_14923);
nor U16132 (N_16132,N_15559,N_12732);
or U16133 (N_16133,N_12383,N_14861);
or U16134 (N_16134,N_14591,N_14799);
or U16135 (N_16135,N_13366,N_13546);
and U16136 (N_16136,N_14700,N_13365);
nand U16137 (N_16137,N_12048,N_14047);
and U16138 (N_16138,N_13645,N_12367);
or U16139 (N_16139,N_14968,N_13784);
or U16140 (N_16140,N_15139,N_15458);
and U16141 (N_16141,N_12204,N_15657);
nand U16142 (N_16142,N_15993,N_12337);
or U16143 (N_16143,N_14099,N_13885);
nor U16144 (N_16144,N_12622,N_13848);
and U16145 (N_16145,N_15918,N_12358);
or U16146 (N_16146,N_12101,N_15425);
nor U16147 (N_16147,N_14599,N_15970);
nor U16148 (N_16148,N_12874,N_13426);
and U16149 (N_16149,N_14622,N_13454);
and U16150 (N_16150,N_14370,N_15801);
nand U16151 (N_16151,N_12394,N_15899);
and U16152 (N_16152,N_13490,N_12864);
nor U16153 (N_16153,N_14905,N_12001);
nand U16154 (N_16154,N_13448,N_13198);
nor U16155 (N_16155,N_14127,N_13378);
and U16156 (N_16156,N_14911,N_14075);
and U16157 (N_16157,N_15416,N_12511);
and U16158 (N_16158,N_15706,N_12553);
and U16159 (N_16159,N_13560,N_14097);
and U16160 (N_16160,N_15769,N_14320);
and U16161 (N_16161,N_13104,N_13137);
or U16162 (N_16162,N_15645,N_12781);
or U16163 (N_16163,N_15554,N_15364);
nor U16164 (N_16164,N_14889,N_15003);
and U16165 (N_16165,N_14558,N_15621);
nand U16166 (N_16166,N_14629,N_13358);
or U16167 (N_16167,N_15188,N_14657);
nor U16168 (N_16168,N_14221,N_12291);
nor U16169 (N_16169,N_15763,N_14008);
or U16170 (N_16170,N_13293,N_14788);
and U16171 (N_16171,N_12951,N_13642);
or U16172 (N_16172,N_13703,N_15845);
and U16173 (N_16173,N_15468,N_15426);
nand U16174 (N_16174,N_13589,N_14495);
nand U16175 (N_16175,N_15260,N_12575);
nor U16176 (N_16176,N_13451,N_15245);
nand U16177 (N_16177,N_14419,N_12462);
nor U16178 (N_16178,N_15433,N_12148);
or U16179 (N_16179,N_15968,N_13923);
or U16180 (N_16180,N_15232,N_12906);
or U16181 (N_16181,N_14225,N_13988);
nor U16182 (N_16182,N_15542,N_12515);
and U16183 (N_16183,N_13032,N_14405);
or U16184 (N_16184,N_13882,N_14131);
nand U16185 (N_16185,N_13399,N_14150);
nor U16186 (N_16186,N_15697,N_12554);
or U16187 (N_16187,N_12893,N_14411);
nand U16188 (N_16188,N_13073,N_15826);
nand U16189 (N_16189,N_13773,N_14567);
or U16190 (N_16190,N_13383,N_14238);
or U16191 (N_16191,N_14448,N_14156);
nor U16192 (N_16192,N_12247,N_14138);
nand U16193 (N_16193,N_14244,N_14462);
nand U16194 (N_16194,N_12056,N_12033);
and U16195 (N_16195,N_13999,N_12051);
nand U16196 (N_16196,N_15236,N_15656);
nand U16197 (N_16197,N_15294,N_15956);
or U16198 (N_16198,N_13745,N_12310);
and U16199 (N_16199,N_14385,N_12603);
nor U16200 (N_16200,N_13013,N_15900);
and U16201 (N_16201,N_13898,N_13480);
nor U16202 (N_16202,N_13133,N_14459);
and U16203 (N_16203,N_12803,N_14754);
and U16204 (N_16204,N_14694,N_14732);
and U16205 (N_16205,N_12474,N_14533);
nand U16206 (N_16206,N_15338,N_13584);
or U16207 (N_16207,N_15868,N_12477);
nand U16208 (N_16208,N_14755,N_13256);
or U16209 (N_16209,N_12948,N_13986);
nand U16210 (N_16210,N_12060,N_12487);
and U16211 (N_16211,N_14426,N_15500);
or U16212 (N_16212,N_12094,N_12378);
nand U16213 (N_16213,N_13970,N_15894);
nand U16214 (N_16214,N_12301,N_14304);
and U16215 (N_16215,N_12422,N_12319);
or U16216 (N_16216,N_13841,N_15595);
nand U16217 (N_16217,N_13106,N_12355);
nor U16218 (N_16218,N_14017,N_13219);
nor U16219 (N_16219,N_12187,N_14683);
and U16220 (N_16220,N_14322,N_12871);
nand U16221 (N_16221,N_14642,N_14423);
or U16222 (N_16222,N_14055,N_13913);
nor U16223 (N_16223,N_15350,N_14996);
nand U16224 (N_16224,N_12576,N_13207);
or U16225 (N_16225,N_14336,N_14809);
and U16226 (N_16226,N_14434,N_15265);
and U16227 (N_16227,N_13349,N_13580);
or U16228 (N_16228,N_13171,N_15451);
nor U16229 (N_16229,N_12057,N_13200);
and U16230 (N_16230,N_14054,N_14387);
or U16231 (N_16231,N_14907,N_13511);
and U16232 (N_16232,N_13500,N_13886);
nand U16233 (N_16233,N_14417,N_15638);
and U16234 (N_16234,N_13523,N_12675);
and U16235 (N_16235,N_15566,N_15902);
xor U16236 (N_16236,N_14768,N_14281);
or U16237 (N_16237,N_12971,N_14070);
nor U16238 (N_16238,N_13883,N_12285);
or U16239 (N_16239,N_14767,N_14730);
nand U16240 (N_16240,N_12472,N_13628);
or U16241 (N_16241,N_14400,N_13031);
nand U16242 (N_16242,N_12138,N_15322);
nand U16243 (N_16243,N_12964,N_13012);
nand U16244 (N_16244,N_12074,N_13640);
or U16245 (N_16245,N_14836,N_12751);
nor U16246 (N_16246,N_13701,N_12046);
nand U16247 (N_16247,N_13481,N_13274);
nand U16248 (N_16248,N_15117,N_13929);
nand U16249 (N_16249,N_14789,N_13252);
or U16250 (N_16250,N_14314,N_15966);
nand U16251 (N_16251,N_12702,N_15023);
nor U16252 (N_16252,N_15648,N_15274);
nand U16253 (N_16253,N_14293,N_15812);
nor U16254 (N_16254,N_12844,N_15247);
nand U16255 (N_16255,N_15491,N_12198);
nand U16256 (N_16256,N_15423,N_14089);
nor U16257 (N_16257,N_14327,N_12920);
or U16258 (N_16258,N_13339,N_12336);
and U16259 (N_16259,N_13702,N_14993);
or U16260 (N_16260,N_15417,N_12506);
nand U16261 (N_16261,N_15177,N_14718);
or U16262 (N_16262,N_13896,N_12440);
nand U16263 (N_16263,N_13514,N_15115);
nand U16264 (N_16264,N_13384,N_12580);
or U16265 (N_16265,N_12929,N_14300);
or U16266 (N_16266,N_15742,N_13936);
or U16267 (N_16267,N_14872,N_12203);
nand U16268 (N_16268,N_15780,N_12837);
nor U16269 (N_16269,N_14309,N_13351);
nor U16270 (N_16270,N_13608,N_14009);
nand U16271 (N_16271,N_15620,N_14032);
or U16272 (N_16272,N_15050,N_15901);
or U16273 (N_16273,N_12497,N_12507);
nand U16274 (N_16274,N_12854,N_12918);
or U16275 (N_16275,N_14807,N_13638);
nand U16276 (N_16276,N_14210,N_15506);
nor U16277 (N_16277,N_14595,N_13101);
and U16278 (N_16278,N_13940,N_15479);
and U16279 (N_16279,N_12011,N_13809);
and U16280 (N_16280,N_13835,N_12130);
or U16281 (N_16281,N_13087,N_12542);
nor U16282 (N_16282,N_12273,N_15699);
or U16283 (N_16283,N_15985,N_14103);
or U16284 (N_16284,N_15442,N_15181);
nor U16285 (N_16285,N_13656,N_14093);
and U16286 (N_16286,N_15810,N_14416);
nor U16287 (N_16287,N_12526,N_15354);
nor U16288 (N_16288,N_15823,N_15516);
nor U16289 (N_16289,N_15220,N_14371);
nand U16290 (N_16290,N_14638,N_12681);
and U16291 (N_16291,N_15672,N_15591);
nor U16292 (N_16292,N_12409,N_12068);
nor U16293 (N_16293,N_12423,N_15436);
or U16294 (N_16294,N_13128,N_15019);
or U16295 (N_16295,N_12564,N_13317);
and U16296 (N_16296,N_15196,N_14610);
nor U16297 (N_16297,N_14570,N_12272);
and U16298 (N_16298,N_15961,N_13942);
and U16299 (N_16299,N_15983,N_13990);
and U16300 (N_16300,N_13673,N_15694);
or U16301 (N_16301,N_12952,N_15871);
and U16302 (N_16302,N_14428,N_15041);
and U16303 (N_16303,N_15846,N_12220);
or U16304 (N_16304,N_13832,N_14442);
and U16305 (N_16305,N_13141,N_13291);
xor U16306 (N_16306,N_13067,N_15406);
nand U16307 (N_16307,N_15308,N_14913);
or U16308 (N_16308,N_14697,N_12397);
nor U16309 (N_16309,N_14340,N_12129);
and U16310 (N_16310,N_12147,N_13321);
or U16311 (N_16311,N_13163,N_13532);
and U16312 (N_16312,N_13914,N_13768);
nor U16313 (N_16313,N_12746,N_15464);
nor U16314 (N_16314,N_14454,N_12509);
nand U16315 (N_16315,N_13464,N_13436);
or U16316 (N_16316,N_14198,N_13740);
nor U16317 (N_16317,N_15696,N_14239);
and U16318 (N_16318,N_13059,N_14876);
nand U16319 (N_16319,N_15277,N_14083);
nor U16320 (N_16320,N_12780,N_14643);
or U16321 (N_16321,N_15387,N_14022);
nor U16322 (N_16322,N_12533,N_15558);
nand U16323 (N_16323,N_12534,N_15884);
nor U16324 (N_16324,N_15392,N_12983);
and U16325 (N_16325,N_13718,N_12414);
or U16326 (N_16326,N_15482,N_14194);
nand U16327 (N_16327,N_12186,N_12881);
nand U16328 (N_16328,N_13911,N_12825);
or U16329 (N_16329,N_14987,N_12463);
or U16330 (N_16330,N_14379,N_13449);
and U16331 (N_16331,N_12841,N_15152);
nand U16332 (N_16332,N_12090,N_12838);
nand U16333 (N_16333,N_13267,N_12460);
or U16334 (N_16334,N_12073,N_15476);
nand U16335 (N_16335,N_12522,N_12279);
or U16336 (N_16336,N_14808,N_12680);
or U16337 (N_16337,N_13495,N_13294);
nor U16338 (N_16338,N_15284,N_12438);
and U16339 (N_16339,N_14845,N_13266);
nand U16340 (N_16340,N_13995,N_13176);
or U16341 (N_16341,N_12626,N_15711);
nor U16342 (N_16342,N_12721,N_12105);
and U16343 (N_16343,N_12255,N_14862);
and U16344 (N_16344,N_14575,N_12642);
nor U16345 (N_16345,N_13188,N_14355);
and U16346 (N_16346,N_15837,N_15800);
and U16347 (N_16347,N_13518,N_12822);
nand U16348 (N_16348,N_15632,N_13409);
and U16349 (N_16349,N_14217,N_15402);
or U16350 (N_16350,N_14908,N_15649);
nor U16351 (N_16351,N_12473,N_15712);
nand U16352 (N_16352,N_14646,N_12037);
nor U16353 (N_16353,N_15898,N_12411);
and U16354 (N_16354,N_12342,N_15092);
nand U16355 (N_16355,N_14435,N_15077);
or U16356 (N_16356,N_12608,N_14063);
nand U16357 (N_16357,N_15691,N_14250);
nor U16358 (N_16358,N_15324,N_14313);
nor U16359 (N_16359,N_15073,N_15378);
or U16360 (N_16360,N_15737,N_14849);
xnor U16361 (N_16361,N_15264,N_12262);
nand U16362 (N_16362,N_15553,N_12469);
nor U16363 (N_16363,N_15317,N_13042);
or U16364 (N_16364,N_14222,N_15303);
or U16365 (N_16365,N_15935,N_12671);
or U16366 (N_16366,N_14308,N_14820);
nand U16367 (N_16367,N_15081,N_14976);
nor U16368 (N_16368,N_15114,N_14170);
nor U16369 (N_16369,N_12259,N_13353);
or U16370 (N_16370,N_14852,N_13927);
nor U16371 (N_16371,N_14193,N_13865);
and U16372 (N_16372,N_13263,N_15678);
nor U16373 (N_16373,N_12341,N_13845);
and U16374 (N_16374,N_15856,N_14959);
nand U16375 (N_16375,N_12858,N_14476);
or U16376 (N_16376,N_14609,N_15330);
and U16377 (N_16377,N_12933,N_12012);
and U16378 (N_16378,N_15668,N_13234);
nor U16379 (N_16379,N_12972,N_15215);
or U16380 (N_16380,N_15046,N_13625);
or U16381 (N_16381,N_15562,N_14050);
and U16382 (N_16382,N_13978,N_14342);
or U16383 (N_16383,N_12795,N_15319);
nor U16384 (N_16384,N_15490,N_12708);
nand U16385 (N_16385,N_12565,N_15118);
or U16386 (N_16386,N_12799,N_15421);
xnor U16387 (N_16387,N_14506,N_12530);
nand U16388 (N_16388,N_12399,N_13738);
nand U16389 (N_16389,N_15610,N_14503);
or U16390 (N_16390,N_12095,N_14303);
or U16391 (N_16391,N_13802,N_15975);
and U16392 (N_16392,N_15596,N_12093);
nor U16393 (N_16393,N_13553,N_15222);
nand U16394 (N_16394,N_15738,N_14364);
xor U16395 (N_16395,N_14069,N_14255);
nand U16396 (N_16396,N_15399,N_14795);
nor U16397 (N_16397,N_13497,N_14786);
and U16398 (N_16398,N_15221,N_14329);
or U16399 (N_16399,N_14229,N_15589);
nor U16400 (N_16400,N_12878,N_15692);
nand U16401 (N_16401,N_12400,N_15863);
nand U16402 (N_16402,N_14235,N_12195);
or U16403 (N_16403,N_12980,N_15085);
or U16404 (N_16404,N_15893,N_15635);
nor U16405 (N_16405,N_13690,N_15055);
nor U16406 (N_16406,N_12713,N_15353);
nor U16407 (N_16407,N_14596,N_12975);
or U16408 (N_16408,N_12868,N_15172);
and U16409 (N_16409,N_12108,N_15448);
and U16410 (N_16410,N_14765,N_12763);
and U16411 (N_16411,N_13206,N_12922);
and U16412 (N_16412,N_13906,N_12213);
nand U16413 (N_16413,N_14029,N_12606);
nand U16414 (N_16414,N_12218,N_13429);
nand U16415 (N_16415,N_12027,N_14129);
nand U16416 (N_16416,N_15203,N_12207);
nand U16417 (N_16417,N_14678,N_14757);
nor U16418 (N_16418,N_12986,N_13756);
nor U16419 (N_16419,N_14548,N_14651);
or U16420 (N_16420,N_15428,N_12338);
and U16421 (N_16421,N_12995,N_13450);
or U16422 (N_16422,N_12492,N_15228);
nand U16423 (N_16423,N_15718,N_13653);
nand U16424 (N_16424,N_12339,N_12742);
and U16425 (N_16425,N_13685,N_13694);
nor U16426 (N_16426,N_13880,N_13958);
or U16427 (N_16427,N_13717,N_13471);
and U16428 (N_16428,N_12246,N_13543);
or U16429 (N_16429,N_14151,N_14626);
and U16430 (N_16430,N_12639,N_13873);
and U16431 (N_16431,N_15929,N_14812);
nand U16432 (N_16432,N_13818,N_12097);
nor U16433 (N_16433,N_14049,N_12866);
nand U16434 (N_16434,N_15716,N_13277);
or U16435 (N_16435,N_14251,N_12537);
or U16436 (N_16436,N_14747,N_14100);
nand U16437 (N_16437,N_14107,N_14201);
nand U16438 (N_16438,N_13682,N_14147);
nand U16439 (N_16439,N_12946,N_14177);
nor U16440 (N_16440,N_12555,N_13839);
and U16441 (N_16441,N_13318,N_15886);
nor U16442 (N_16442,N_12861,N_12164);
or U16443 (N_16443,N_15488,N_14016);
nor U16444 (N_16444,N_13082,N_12879);
and U16445 (N_16445,N_14869,N_12719);
and U16446 (N_16446,N_15733,N_12471);
nand U16447 (N_16447,N_15297,N_15660);
nor U16448 (N_16448,N_12323,N_14215);
and U16449 (N_16449,N_12594,N_14822);
and U16450 (N_16450,N_15539,N_13213);
nor U16451 (N_16451,N_12270,N_12444);
nand U16452 (N_16452,N_12171,N_14324);
nor U16453 (N_16453,N_13781,N_13493);
nor U16454 (N_16454,N_15480,N_12668);
nand U16455 (N_16455,N_15070,N_13649);
nor U16456 (N_16456,N_12165,N_13971);
or U16457 (N_16457,N_12417,N_13540);
nand U16458 (N_16458,N_12102,N_14924);
nand U16459 (N_16459,N_13966,N_14152);
nand U16460 (N_16460,N_12816,N_15210);
and U16461 (N_16461,N_13955,N_12156);
nand U16462 (N_16462,N_15235,N_12567);
nor U16463 (N_16463,N_13007,N_13636);
or U16464 (N_16464,N_14723,N_13586);
and U16465 (N_16465,N_12170,N_13117);
nor U16466 (N_16466,N_12278,N_12496);
nor U16467 (N_16467,N_13470,N_13693);
or U16468 (N_16468,N_14710,N_12340);
or U16469 (N_16469,N_15574,N_13438);
nand U16470 (N_16470,N_15914,N_14122);
nor U16471 (N_16471,N_13732,N_13535);
or U16472 (N_16472,N_14576,N_14051);
or U16473 (N_16473,N_13099,N_15741);
and U16474 (N_16474,N_13591,N_14585);
nand U16475 (N_16475,N_14199,N_14289);
nand U16476 (N_16476,N_14928,N_12300);
nor U16477 (N_16477,N_14021,N_12126);
or U16478 (N_16478,N_12321,N_14727);
nor U16479 (N_16479,N_13585,N_12481);
or U16480 (N_16480,N_13199,N_12911);
nand U16481 (N_16481,N_14436,N_12328);
nor U16482 (N_16482,N_13307,N_12257);
nand U16483 (N_16483,N_12225,N_13522);
and U16484 (N_16484,N_12254,N_12548);
or U16485 (N_16485,N_15953,N_13601);
or U16486 (N_16486,N_15435,N_13452);
nand U16487 (N_16487,N_13634,N_15807);
nor U16488 (N_16488,N_12313,N_12196);
or U16489 (N_16489,N_14593,N_15927);
or U16490 (N_16490,N_14895,N_15725);
nor U16491 (N_16491,N_15225,N_12233);
nand U16492 (N_16492,N_15499,N_13689);
and U16493 (N_16493,N_15103,N_15299);
and U16494 (N_16494,N_14382,N_12230);
nor U16495 (N_16495,N_14496,N_14984);
nand U16496 (N_16496,N_15804,N_12330);
nand U16497 (N_16497,N_15981,N_12183);
or U16498 (N_16498,N_15907,N_13215);
nand U16499 (N_16499,N_15300,N_15617);
and U16500 (N_16500,N_15527,N_15561);
nor U16501 (N_16501,N_13921,N_12846);
or U16502 (N_16502,N_15578,N_13157);
nand U16503 (N_16503,N_15359,N_15414);
and U16504 (N_16504,N_12633,N_13594);
and U16505 (N_16505,N_12821,N_12202);
and U16506 (N_16506,N_12677,N_12280);
or U16507 (N_16507,N_15459,N_13165);
or U16508 (N_16508,N_15349,N_12178);
nor U16509 (N_16509,N_15302,N_12107);
or U16510 (N_16510,N_13222,N_15677);
and U16511 (N_16511,N_15257,N_14776);
and U16512 (N_16512,N_12882,N_12769);
nor U16513 (N_16513,N_15987,N_12617);
and U16514 (N_16514,N_12706,N_13538);
nand U16515 (N_16515,N_12260,N_12849);
or U16516 (N_16516,N_13780,N_13335);
nor U16517 (N_16517,N_12917,N_13730);
nand U16518 (N_16518,N_14612,N_15105);
nand U16519 (N_16519,N_13377,N_14132);
and U16520 (N_16520,N_14187,N_12790);
or U16521 (N_16521,N_14276,N_14930);
or U16522 (N_16522,N_15504,N_14298);
nand U16523 (N_16523,N_15830,N_14450);
and U16524 (N_16524,N_15795,N_14475);
and U16525 (N_16525,N_12770,N_14983);
and U16526 (N_16526,N_12991,N_13404);
nand U16527 (N_16527,N_12249,N_13006);
nor U16528 (N_16528,N_14315,N_12696);
nor U16529 (N_16529,N_14145,N_15358);
nand U16530 (N_16530,N_14189,N_12306);
nor U16531 (N_16531,N_13786,N_14254);
or U16532 (N_16532,N_15796,N_15347);
and U16533 (N_16533,N_13741,N_15062);
nand U16534 (N_16534,N_15785,N_12752);
nand U16535 (N_16535,N_12904,N_14430);
and U16536 (N_16536,N_15205,N_12172);
nor U16537 (N_16537,N_15379,N_15076);
or U16538 (N_16538,N_13063,N_12019);
or U16539 (N_16539,N_15730,N_14915);
and U16540 (N_16540,N_12062,N_14580);
and U16541 (N_16541,N_13488,N_14902);
and U16542 (N_16542,N_15465,N_14743);
nor U16543 (N_16543,N_14188,N_14744);
nor U16544 (N_16544,N_12989,N_15093);
nor U16545 (N_16545,N_13325,N_14333);
nor U16546 (N_16546,N_14969,N_14856);
or U16547 (N_16547,N_15016,N_13797);
or U16548 (N_16548,N_15865,N_12711);
and U16549 (N_16549,N_15240,N_15143);
nand U16550 (N_16550,N_15519,N_15754);
or U16551 (N_16551,N_15685,N_14892);
or U16552 (N_16552,N_14242,N_13272);
or U16553 (N_16553,N_13662,N_13397);
nand U16554 (N_16554,N_12850,N_13919);
nor U16555 (N_16555,N_15870,N_14290);
or U16556 (N_16556,N_12245,N_13417);
nand U16557 (N_16557,N_13382,N_15000);
and U16558 (N_16558,N_12943,N_12356);
or U16559 (N_16559,N_15652,N_14654);
nor U16560 (N_16560,N_13981,N_12034);
and U16561 (N_16561,N_14890,N_12293);
nor U16562 (N_16562,N_12018,N_13536);
nor U16563 (N_16563,N_12010,N_14530);
nand U16564 (N_16564,N_15622,N_14542);
nand U16565 (N_16565,N_12992,N_12566);
nor U16566 (N_16566,N_13728,N_12930);
nor U16567 (N_16567,N_14130,N_12717);
nand U16568 (N_16568,N_15441,N_12450);
nor U16569 (N_16569,N_15748,N_13392);
or U16570 (N_16570,N_13465,N_12021);
nor U16571 (N_16571,N_13722,N_12857);
nand U16572 (N_16572,N_15681,N_14354);
or U16573 (N_16573,N_13765,N_13954);
nand U16574 (N_16574,N_13319,N_15306);
nor U16575 (N_16575,N_13129,N_12966);
nand U16576 (N_16576,N_15552,N_13161);
and U16577 (N_16577,N_12690,N_12392);
nand U16578 (N_16578,N_12197,N_14490);
nand U16579 (N_16579,N_13430,N_12891);
nor U16580 (N_16580,N_15341,N_15394);
nand U16581 (N_16581,N_15456,N_13907);
and U16582 (N_16582,N_15298,N_15025);
or U16583 (N_16583,N_13801,N_15400);
or U16584 (N_16584,N_13154,N_13805);
or U16585 (N_16585,N_12709,N_14884);
and U16586 (N_16586,N_12420,N_14172);
xnor U16587 (N_16587,N_14481,N_13427);
nand U16588 (N_16588,N_14603,N_15565);
nor U16589 (N_16589,N_12583,N_12977);
nand U16590 (N_16590,N_13785,N_13264);
or U16591 (N_16591,N_13599,N_13487);
nor U16592 (N_16592,N_12419,N_13287);
nand U16593 (N_16593,N_12551,N_15024);
and U16594 (N_16594,N_12664,N_15086);
nor U16595 (N_16595,N_13126,N_13631);
nand U16596 (N_16596,N_14071,N_13017);
and U16597 (N_16597,N_15474,N_13939);
or U16598 (N_16598,N_13665,N_14082);
xor U16599 (N_16599,N_15958,N_15332);
or U16600 (N_16600,N_14837,N_14554);
or U16601 (N_16601,N_12561,N_15749);
nor U16602 (N_16602,N_14875,N_15715);
or U16603 (N_16603,N_13113,N_12275);
nand U16604 (N_16604,N_12734,N_15089);
nor U16605 (N_16605,N_12653,N_12119);
or U16606 (N_16606,N_14607,N_13564);
nand U16607 (N_16607,N_13173,N_12634);
nand U16608 (N_16608,N_14384,N_15022);
nand U16609 (N_16609,N_15230,N_13664);
and U16610 (N_16610,N_14274,N_12256);
and U16611 (N_16611,N_15563,N_14278);
or U16612 (N_16612,N_15237,N_14154);
nor U16613 (N_16613,N_12998,N_12502);
or U16614 (N_16614,N_13422,N_15702);
and U16615 (N_16615,N_13160,N_13064);
nor U16616 (N_16616,N_15875,N_12683);
nand U16617 (N_16617,N_15765,N_12643);
or U16618 (N_16618,N_12022,N_14488);
nor U16619 (N_16619,N_13563,N_13014);
and U16620 (N_16620,N_15074,N_13076);
nand U16621 (N_16621,N_12386,N_15960);
nand U16622 (N_16622,N_14873,N_15690);
or U16623 (N_16623,N_13968,N_15615);
nand U16624 (N_16624,N_15582,N_13210);
nor U16625 (N_16625,N_13554,N_12649);
nand U16626 (N_16626,N_14719,N_12650);
nor U16627 (N_16627,N_14038,N_13419);
and U16628 (N_16628,N_12274,N_15431);
nor U16629 (N_16629,N_15029,N_12370);
and U16630 (N_16630,N_15905,N_15557);
or U16631 (N_16631,N_14963,N_13492);
or U16632 (N_16632,N_13072,N_14664);
nand U16633 (N_16633,N_15818,N_13504);
or U16634 (N_16634,N_12679,N_13840);
or U16635 (N_16635,N_14248,N_13225);
nor U16636 (N_16636,N_15897,N_13249);
and U16637 (N_16637,N_15129,N_12467);
or U16638 (N_16638,N_12479,N_13729);
and U16639 (N_16639,N_13941,N_13140);
and U16640 (N_16640,N_12276,N_15919);
or U16641 (N_16641,N_15250,N_14766);
nand U16642 (N_16642,N_13052,N_12809);
nand U16643 (N_16643,N_13295,N_13093);
nor U16644 (N_16644,N_13779,N_15751);
nor U16645 (N_16645,N_13519,N_12637);
or U16646 (N_16646,N_13559,N_15279);
and U16647 (N_16647,N_15992,N_14966);
nand U16648 (N_16648,N_12826,N_15057);
nor U16649 (N_16649,N_12261,N_14759);
and U16650 (N_16650,N_14665,N_14956);
nand U16651 (N_16651,N_14457,N_15495);
or U16652 (N_16652,N_15147,N_14404);
and U16653 (N_16653,N_12851,N_12015);
nor U16654 (N_16654,N_15457,N_13051);
nand U16655 (N_16655,N_12353,N_15174);
nand U16656 (N_16656,N_15040,N_14640);
and U16657 (N_16657,N_14738,N_12219);
nand U16658 (N_16658,N_12307,N_13905);
and U16659 (N_16659,N_14980,N_13747);
nand U16660 (N_16660,N_13211,N_15422);
nand U16661 (N_16661,N_15119,N_15560);
or U16662 (N_16662,N_14391,N_12513);
nor U16663 (N_16663,N_15533,N_13750);
and U16664 (N_16664,N_13590,N_14617);
nand U16665 (N_16665,N_13938,N_12308);
or U16666 (N_16666,N_15037,N_12557);
and U16667 (N_16667,N_12648,N_14589);
or U16668 (N_16668,N_14952,N_15923);
and U16669 (N_16669,N_14026,N_13713);
nor U16670 (N_16670,N_13127,N_13435);
or U16671 (N_16671,N_12937,N_15586);
or U16672 (N_16672,N_14334,N_12269);
nor U16673 (N_16673,N_15099,N_13770);
and U16674 (N_16674,N_13726,N_13895);
nor U16675 (N_16675,N_15278,N_12830);
and U16676 (N_16676,N_15471,N_14002);
nand U16677 (N_16677,N_12364,N_15515);
nor U16678 (N_16678,N_13328,N_15010);
nand U16679 (N_16679,N_12379,N_14429);
nand U16680 (N_16680,N_12252,N_15038);
or U16681 (N_16681,N_13315,N_12166);
or U16682 (N_16682,N_13655,N_12694);
nor U16683 (N_16683,N_14356,N_13387);
or U16684 (N_16684,N_12289,N_15628);
nor U16685 (N_16685,N_14741,N_14326);
or U16686 (N_16686,N_13220,N_12098);
nand U16687 (N_16687,N_15390,N_13010);
nand U16688 (N_16688,N_14810,N_14505);
nor U16689 (N_16689,N_14752,N_15339);
and U16690 (N_16690,N_14504,N_14414);
and U16691 (N_16691,N_15903,N_15053);
nor U16692 (N_16692,N_12630,N_15251);
or U16693 (N_16693,N_14105,N_13944);
or U16694 (N_16694,N_15301,N_13164);
and U16695 (N_16695,N_13537,N_15173);
nor U16696 (N_16696,N_14498,N_14024);
or U16697 (N_16697,N_14695,N_13248);
nor U16698 (N_16698,N_13499,N_15891);
nand U16699 (N_16699,N_14559,N_15192);
or U16700 (N_16700,N_13179,N_15307);
nand U16701 (N_16701,N_14590,N_14960);
nor U16702 (N_16702,N_14374,N_12014);
nand U16703 (N_16703,N_14121,N_13695);
nor U16704 (N_16704,N_12372,N_14906);
nor U16705 (N_16705,N_14109,N_12114);
or U16706 (N_16706,N_15083,N_15534);
or U16707 (N_16707,N_13374,N_13111);
or U16708 (N_16708,N_15776,N_12447);
nand U16709 (N_16709,N_15068,N_12823);
or U16710 (N_16710,N_15223,N_12127);
nor U16711 (N_16711,N_13897,N_13275);
nand U16712 (N_16712,N_15964,N_14510);
nor U16713 (N_16713,N_13652,N_15844);
xor U16714 (N_16714,N_15100,N_12973);
nand U16715 (N_16715,N_15090,N_13899);
and U16716 (N_16716,N_14839,N_14301);
nand U16717 (N_16717,N_15140,N_14307);
and U16718 (N_16718,N_15892,N_14756);
xnor U16719 (N_16719,N_15505,N_15101);
and U16720 (N_16720,N_12016,N_13731);
or U16721 (N_16721,N_13961,N_15132);
or U16722 (N_16722,N_13754,N_15430);
or U16723 (N_16723,N_13644,N_14933);
or U16724 (N_16724,N_12609,N_13411);
or U16725 (N_16725,N_15788,N_14040);
or U16726 (N_16726,N_13170,N_15489);
nand U16727 (N_16727,N_12066,N_13758);
or U16728 (N_16728,N_13527,N_13602);
nor U16729 (N_16729,N_15291,N_15701);
nor U16730 (N_16730,N_15005,N_12125);
nand U16731 (N_16731,N_12666,N_14218);
xnor U16732 (N_16732,N_15783,N_15373);
nor U16733 (N_16733,N_14631,N_13261);
and U16734 (N_16734,N_12005,N_13322);
nand U16735 (N_16735,N_13828,N_15375);
and U16736 (N_16736,N_13525,N_15381);
nand U16737 (N_16737,N_13798,N_13847);
or U16738 (N_16738,N_15687,N_13035);
and U16739 (N_16739,N_14805,N_13314);
nand U16740 (N_16740,N_12181,N_14532);
and U16741 (N_16741,N_14139,N_13265);
or U16742 (N_16742,N_14936,N_12700);
and U16743 (N_16743,N_15102,N_12806);
nand U16744 (N_16744,N_15385,N_12465);
nand U16745 (N_16745,N_12201,N_15082);
and U16746 (N_16746,N_14226,N_15758);
and U16747 (N_16747,N_12250,N_12128);
and U16748 (N_16748,N_12845,N_13716);
and U16749 (N_16749,N_14283,N_14232);
or U16750 (N_16750,N_13926,N_12627);
nor U16751 (N_16751,N_14556,N_15772);
and U16752 (N_16752,N_13720,N_14357);
or U16753 (N_16753,N_12374,N_15473);
nand U16754 (N_16754,N_14893,N_15997);
nor U16755 (N_16755,N_13236,N_12216);
and U16756 (N_16756,N_14920,N_14359);
xnor U16757 (N_16757,N_15493,N_15113);
or U16758 (N_16758,N_13789,N_15030);
nor U16759 (N_16759,N_14877,N_12877);
nor U16760 (N_16760,N_13963,N_12898);
and U16761 (N_16761,N_14363,N_12875);
nand U16762 (N_16762,N_12584,N_14826);
and U16763 (N_16763,N_12038,N_12574);
nor U16764 (N_16764,N_14466,N_13515);
or U16765 (N_16765,N_14039,N_13421);
and U16766 (N_16766,N_14433,N_13124);
nand U16767 (N_16767,N_12957,N_15972);
nor U16768 (N_16768,N_12023,N_15739);
nand U16769 (N_16769,N_12428,N_15693);
nor U16770 (N_16770,N_14739,N_12824);
or U16771 (N_16771,N_12902,N_12999);
nand U16772 (N_16772,N_12976,N_14746);
nand U16773 (N_16773,N_12070,N_13125);
nand U16774 (N_16774,N_15984,N_14880);
and U16775 (N_16775,N_12266,N_14000);
and U16776 (N_16776,N_12601,N_14823);
nand U16777 (N_16777,N_12402,N_12657);
and U16778 (N_16778,N_12510,N_13005);
or U16779 (N_16779,N_12464,N_15705);
or U16780 (N_16780,N_14292,N_13507);
and U16781 (N_16781,N_13544,N_14349);
nand U16782 (N_16782,N_13892,N_13846);
nor U16783 (N_16783,N_13829,N_12547);
and U16784 (N_16784,N_13416,N_12425);
xor U16785 (N_16785,N_12088,N_12485);
nand U16786 (N_16786,N_14380,N_14390);
and U16787 (N_16787,N_12945,N_12691);
and U16788 (N_16788,N_12331,N_14015);
and U16789 (N_16789,N_13932,N_15764);
nand U16790 (N_16790,N_12013,N_13463);
xor U16791 (N_16791,N_13587,N_12086);
nand U16792 (N_16792,N_12369,N_13168);
nand U16793 (N_16793,N_15806,N_13241);
nor U16794 (N_16794,N_15700,N_15467);
or U16795 (N_16795,N_13247,N_14833);
nand U16796 (N_16796,N_13837,N_12905);
nand U16797 (N_16797,N_12111,N_12085);
nor U16798 (N_16798,N_13453,N_13900);
or U16799 (N_16799,N_15179,N_13810);
nor U16800 (N_16800,N_14863,N_14376);
nor U16801 (N_16801,N_14478,N_15079);
nor U16802 (N_16802,N_14291,N_12235);
nor U16803 (N_16803,N_12938,N_14978);
or U16804 (N_16804,N_15481,N_15545);
and U16805 (N_16805,N_15937,N_13258);
and U16806 (N_16806,N_13737,N_15881);
nor U16807 (N_16807,N_15532,N_14418);
or U16808 (N_16808,N_13456,N_15853);
and U16809 (N_16809,N_12381,N_14137);
and U16810 (N_16810,N_13396,N_12672);
or U16811 (N_16811,N_12820,N_12593);
or U16812 (N_16812,N_12589,N_14142);
or U16813 (N_16813,N_15922,N_12699);
nor U16814 (N_16814,N_12518,N_13849);
nand U16815 (N_16815,N_14803,N_14581);
and U16816 (N_16816,N_13434,N_13477);
nor U16817 (N_16817,N_12560,N_13706);
nor U16818 (N_16818,N_12735,N_14702);
nor U16819 (N_16819,N_13245,N_15429);
nand U16820 (N_16820,N_14670,N_15828);
nand U16821 (N_16821,N_15537,N_15676);
nor U16822 (N_16822,N_14619,N_14828);
and U16823 (N_16823,N_14508,N_15614);
nor U16824 (N_16824,N_14181,N_12030);
or U16825 (N_16825,N_14970,N_13212);
and U16826 (N_16826,N_15180,N_14830);
or U16827 (N_16827,N_12059,N_14935);
or U16828 (N_16828,N_14650,N_13735);
or U16829 (N_16829,N_13308,N_15544);
nand U16830 (N_16830,N_14220,N_15189);
and U16831 (N_16831,N_12134,N_12028);
nand U16832 (N_16832,N_14867,N_12997);
nor U16833 (N_16833,N_14636,N_13341);
and U16834 (N_16834,N_15948,N_15990);
and U16835 (N_16835,N_15087,N_14394);
nand U16836 (N_16836,N_12333,N_15920);
and U16837 (N_16837,N_13903,N_13611);
or U16838 (N_16838,N_15455,N_13627);
or U16839 (N_16839,N_14275,N_15609);
nor U16840 (N_16840,N_14817,N_14480);
nor U16841 (N_16841,N_13289,N_12659);
or U16842 (N_16842,N_15405,N_15008);
or U16843 (N_16843,N_15728,N_14621);
or U16844 (N_16844,N_12544,N_12406);
nand U16845 (N_16845,N_15325,N_13512);
and U16846 (N_16846,N_13811,N_14740);
nand U16847 (N_16847,N_13619,N_13657);
nor U16848 (N_16848,N_13376,N_14335);
nand U16849 (N_16849,N_13547,N_15382);
nor U16850 (N_16850,N_12413,N_15162);
or U16851 (N_16851,N_15309,N_15026);
and U16852 (N_16852,N_13501,N_12921);
nor U16853 (N_16853,N_14742,N_15551);
or U16854 (N_16854,N_14310,N_14494);
and U16855 (N_16855,N_15288,N_12137);
nand U16856 (N_16856,N_12692,N_14815);
or U16857 (N_16857,N_13240,N_12185);
and U16858 (N_16858,N_14573,N_15636);
nor U16859 (N_16859,N_12040,N_14445);
nor U16860 (N_16860,N_15007,N_15659);
or U16861 (N_16861,N_15383,N_13517);
nor U16862 (N_16862,N_14144,N_13858);
nor U16863 (N_16863,N_15858,N_14518);
or U16864 (N_16864,N_14834,N_12158);
nand U16865 (N_16865,N_15536,N_13757);
nand U16866 (N_16866,N_12767,N_13684);
and U16867 (N_16867,N_13697,N_12880);
nand U16868 (N_16868,N_13095,N_14211);
nor U16869 (N_16869,N_12527,N_15164);
nor U16870 (N_16870,N_15014,N_14652);
or U16871 (N_16871,N_12036,N_12132);
or U16872 (N_16872,N_15779,N_15510);
nand U16873 (N_16873,N_14485,N_15243);
or U16874 (N_16874,N_15270,N_14432);
or U16875 (N_16875,N_14669,N_12959);
or U16876 (N_16876,N_12265,N_15882);
nand U16877 (N_16877,N_15031,N_15675);
or U16878 (N_16878,N_14422,N_15367);
or U16879 (N_16879,N_14444,N_15827);
nand U16880 (N_16880,N_13742,N_12177);
nor U16881 (N_16881,N_15368,N_13550);
or U16882 (N_16882,N_15619,N_15543);
nor U16883 (N_16883,N_13340,N_14456);
nor U16884 (N_16884,N_13395,N_15917);
and U16885 (N_16885,N_14555,N_13508);
nor U16886 (N_16886,N_12628,N_14989);
or U16887 (N_16887,N_15838,N_14072);
or U16888 (N_16888,N_14192,N_15054);
nor U16889 (N_16889,N_15494,N_13229);
and U16890 (N_16890,N_13071,N_15063);
and U16891 (N_16891,N_15318,N_12412);
or U16892 (N_16892,N_14114,N_12919);
nand U16893 (N_16893,N_14413,N_12978);
or U16894 (N_16894,N_14614,N_14060);
nor U16895 (N_16895,N_12160,N_12884);
or U16896 (N_16896,N_14062,N_14241);
nor U16897 (N_16897,N_15862,N_12818);
nand U16898 (N_16898,N_15750,N_13674);
and U16899 (N_16899,N_15463,N_12453);
nor U16900 (N_16900,N_12950,N_15778);
nand U16901 (N_16901,N_14330,N_14569);
nand U16902 (N_16902,N_15842,N_14399);
and U16903 (N_16903,N_13769,N_15971);
or U16904 (N_16904,N_14673,N_12348);
nand U16905 (N_16905,N_15111,N_13217);
or U16906 (N_16906,N_13282,N_15572);
nor U16907 (N_16907,N_14977,N_13610);
and U16908 (N_16908,N_13381,N_14057);
nand U16909 (N_16909,N_15241,N_14077);
nand U16910 (N_16910,N_14772,N_12611);
nand U16911 (N_16911,N_14373,N_12268);
and U16912 (N_16912,N_15310,N_13489);
nor U16913 (N_16913,N_14545,N_13792);
and U16914 (N_16914,N_15155,N_14325);
or U16915 (N_16915,N_12853,N_13576);
nand U16916 (N_16916,N_13989,N_14410);
or U16917 (N_16917,N_12443,N_14513);
nor U16918 (N_16918,N_12322,N_15167);
nand U16919 (N_16919,N_13259,N_13884);
nand U16920 (N_16920,N_15440,N_15175);
nand U16921 (N_16921,N_12150,N_15002);
nand U16922 (N_16922,N_15703,N_14899);
nor U16923 (N_16923,N_14184,N_13373);
nor U16924 (N_16924,N_15814,N_12248);
nor U16925 (N_16925,N_15889,N_14858);
nand U16926 (N_16926,N_15020,N_14842);
nand U16927 (N_16927,N_13705,N_12887);
or U16928 (N_16928,N_15450,N_12311);
or U16929 (N_16929,N_13842,N_14957);
nand U16930 (N_16930,N_14994,N_12025);
nand U16931 (N_16931,N_15091,N_14066);
nand U16932 (N_16932,N_13026,N_14331);
nand U16933 (N_16933,N_13311,N_14438);
nor U16934 (N_16934,N_14477,N_14471);
or U16935 (N_16935,N_15374,N_13231);
nand U16936 (N_16936,N_14169,N_15986);
or U16937 (N_16937,N_15686,N_14482);
nand U16938 (N_16938,N_12488,N_13203);
nand U16939 (N_16939,N_12054,N_14785);
and U16940 (N_16940,N_15477,N_13983);
nand U16941 (N_16941,N_13056,N_12749);
or U16942 (N_16942,N_14257,N_13091);
nor U16943 (N_16943,N_15994,N_14035);
nand U16944 (N_16944,N_15524,N_13001);
or U16945 (N_16945,N_14831,N_13881);
nand U16946 (N_16946,N_12418,N_14565);
nor U16947 (N_16947,N_13209,N_14102);
or U16948 (N_16948,N_13859,N_14543);
nand U16949 (N_16949,N_14903,N_13152);
and U16950 (N_16950,N_14846,N_14143);
and U16951 (N_16951,N_12136,N_15799);
or U16952 (N_16952,N_13573,N_12556);
nor U16953 (N_16953,N_12796,N_14910);
nor U16954 (N_16954,N_14098,N_12427);
nand U16955 (N_16955,N_14641,N_13987);
or U16956 (N_16956,N_12404,N_13040);
nand U16957 (N_16957,N_15773,N_12546);
nor U16958 (N_16958,N_12153,N_15296);
nor U16959 (N_16959,N_13654,N_15420);
and U16960 (N_16960,N_12552,N_13739);
or U16961 (N_16961,N_14605,N_12020);
and U16962 (N_16962,N_13808,N_13506);
and U16963 (N_16963,N_14223,N_15526);
nand U16964 (N_16964,N_12200,N_12963);
or U16965 (N_16965,N_12759,N_13775);
or U16966 (N_16966,N_13658,N_15883);
nor U16967 (N_16967,N_12512,N_12779);
or U16968 (N_16968,N_14339,N_14790);
or U16969 (N_16969,N_13876,N_15130);
nand U16970 (N_16970,N_12698,N_13850);
nor U16971 (N_16971,N_12135,N_13736);
nand U16972 (N_16972,N_15895,N_12133);
and U16973 (N_16973,N_14511,N_15511);
nor U16974 (N_16974,N_12359,N_15372);
nor U16975 (N_16975,N_13889,N_14461);
or U16976 (N_16976,N_15069,N_12354);
or U16977 (N_16977,N_14285,N_15938);
nor U16978 (N_16978,N_15158,N_12807);
and U16979 (N_16979,N_13869,N_14470);
and U16980 (N_16980,N_13278,N_12475);
and U16981 (N_16981,N_14119,N_13237);
or U16982 (N_16982,N_13197,N_15535);
and U16983 (N_16983,N_15336,N_12834);
and U16984 (N_16984,N_15266,N_12738);
nor U16985 (N_16985,N_15941,N_15497);
nand U16986 (N_16986,N_13853,N_14018);
or U16987 (N_16987,N_13394,N_12897);
and U16988 (N_16988,N_13595,N_12243);
and U16989 (N_16989,N_13753,N_14800);
or U16990 (N_16990,N_13872,N_14348);
or U16991 (N_16991,N_13098,N_13371);
nand U16992 (N_16992,N_14316,N_14541);
and U16993 (N_16993,N_15604,N_15066);
or U16994 (N_16994,N_14056,N_12939);
nor U16995 (N_16995,N_13201,N_14427);
or U16996 (N_16996,N_15564,N_14178);
and U16997 (N_16997,N_13692,N_15792);
nand U16998 (N_16998,N_12468,N_13223);
and U16999 (N_16999,N_15988,N_14031);
nor U17000 (N_17000,N_12489,N_14128);
nand U17001 (N_17001,N_13112,N_14207);
nor U17002 (N_17002,N_14243,N_15512);
or U17003 (N_17003,N_14632,N_14124);
or U17004 (N_17004,N_15954,N_12008);
or U17005 (N_17005,N_14458,N_14486);
nand U17006 (N_17006,N_12281,N_15612);
nor U17007 (N_17007,N_15855,N_13541);
nor U17008 (N_17008,N_15292,N_15186);
nor U17009 (N_17009,N_12332,N_14037);
xnor U17010 (N_17010,N_13185,N_12143);
nor U17011 (N_17011,N_12335,N_13251);
or U17012 (N_17012,N_13097,N_13503);
or U17013 (N_17013,N_14007,N_13524);
or U17014 (N_17014,N_13476,N_15784);
or U17015 (N_17015,N_14552,N_14492);
and U17016 (N_17016,N_13548,N_15695);
or U17017 (N_17017,N_15573,N_12856);
nand U17018 (N_17018,N_12343,N_13964);
and U17019 (N_17019,N_13232,N_12927);
or U17020 (N_17020,N_13457,N_13606);
nand U17021 (N_17021,N_14536,N_15439);
or U17022 (N_17022,N_12041,N_15819);
xor U17023 (N_17023,N_12629,N_13045);
and U17024 (N_17024,N_14167,N_13038);
nand U17025 (N_17025,N_14455,N_13182);
nand U17026 (N_17026,N_14706,N_13359);
nand U17027 (N_17027,N_14551,N_15833);
or U17028 (N_17028,N_14042,N_12592);
nor U17029 (N_17029,N_14701,N_14689);
and U17030 (N_17030,N_13817,N_12726);
or U17031 (N_17031,N_12403,N_12636);
or U17032 (N_17032,N_13260,N_14058);
nor U17033 (N_17033,N_12199,N_14014);
and U17034 (N_17034,N_13916,N_12067);
nand U17035 (N_17035,N_12491,N_15913);
nor U17036 (N_17036,N_13230,N_13156);
nor U17037 (N_17037,N_13583,N_13800);
and U17038 (N_17038,N_13582,N_13733);
or U17039 (N_17039,N_14550,N_12676);
or U17040 (N_17040,N_12723,N_15585);
nand U17041 (N_17041,N_13494,N_15226);
nand U17042 (N_17042,N_15601,N_15211);
or U17043 (N_17043,N_15342,N_13688);
nand U17044 (N_17044,N_12697,N_12890);
and U17045 (N_17045,N_13443,N_12009);
nand U17046 (N_17046,N_14403,N_15408);
nor U17047 (N_17047,N_14079,N_13116);
nor U17048 (N_17048,N_13136,N_15386);
nor U17049 (N_17049,N_13115,N_14753);
nand U17050 (N_17050,N_12077,N_12205);
and U17051 (N_17051,N_14113,N_13469);
nor U17052 (N_17052,N_12039,N_15944);
or U17053 (N_17053,N_13629,N_15682);
nor U17054 (N_17054,N_13034,N_13445);
or U17055 (N_17055,N_12120,N_13027);
and U17056 (N_17056,N_14527,N_14964);
nor U17057 (N_17057,N_14431,N_13575);
and U17058 (N_17058,N_12047,N_13609);
and U17059 (N_17059,N_14473,N_14501);
nand U17060 (N_17060,N_12739,N_13597);
or U17061 (N_17061,N_14048,N_14195);
nand U17062 (N_17062,N_14328,N_12892);
or U17063 (N_17063,N_12194,N_14437);
or U17064 (N_17064,N_13361,N_13479);
nor U17065 (N_17065,N_15683,N_13149);
or U17066 (N_17066,N_12913,N_14821);
nor U17067 (N_17067,N_12718,N_13065);
nor U17068 (N_17068,N_13812,N_12960);
or U17069 (N_17069,N_13836,N_13824);
xor U17070 (N_17070,N_13821,N_13439);
nor U17071 (N_17071,N_12519,N_13974);
nor U17072 (N_17072,N_14855,N_13724);
and U17073 (N_17073,N_12264,N_14864);
and U17074 (N_17074,N_14086,N_15835);
xnor U17075 (N_17075,N_12740,N_15885);
or U17076 (N_17076,N_15708,N_15569);
or U17077 (N_17077,N_12788,N_14745);
or U17078 (N_17078,N_12231,N_13138);
and U17079 (N_17079,N_15658,N_13979);
nand U17080 (N_17080,N_14491,N_12619);
and U17081 (N_17081,N_15362,N_15261);
and U17082 (N_17082,N_14166,N_12661);
and U17083 (N_17083,N_13596,N_15550);
and U17084 (N_17084,N_15822,N_12587);
nand U17085 (N_17085,N_15427,N_12819);
nor U17086 (N_17086,N_12829,N_15775);
and U17087 (N_17087,N_14731,N_14615);
or U17088 (N_17088,N_14816,N_14525);
or U17089 (N_17089,N_15925,N_12814);
xor U17090 (N_17090,N_15653,N_14940);
and U17091 (N_17091,N_13902,N_13593);
and U17092 (N_17092,N_12982,N_13778);
nor U17093 (N_17093,N_14791,N_14868);
nor U17094 (N_17094,N_13316,N_13969);
nand U17095 (N_17095,N_14011,N_12188);
nor U17096 (N_17096,N_14375,N_12304);
and U17097 (N_17097,N_12292,N_14883);
or U17098 (N_17098,N_12663,N_13189);
nand U17099 (N_17099,N_15148,N_13843);
nor U17100 (N_17100,N_12002,N_15015);
and U17101 (N_17101,N_12232,N_14992);
nor U17102 (N_17102,N_15234,N_12640);
and U17103 (N_17103,N_14117,N_14108);
nor U17104 (N_17104,N_14353,N_15168);
or U17105 (N_17105,N_15670,N_12935);
or U17106 (N_17106,N_12550,N_13530);
and U17107 (N_17107,N_12745,N_12258);
nor U17108 (N_17108,N_12539,N_13870);
and U17109 (N_17109,N_15662,N_15263);
and U17110 (N_17110,N_13337,N_12229);
nand U17111 (N_17111,N_13096,N_13679);
nand U17112 (N_17112,N_14841,N_13033);
and U17113 (N_17113,N_13570,N_13271);
and U17114 (N_17114,N_12180,N_15252);
nand U17115 (N_17115,N_13118,N_14392);
and U17116 (N_17116,N_15757,N_12176);
nor U17117 (N_17117,N_15224,N_14350);
or U17118 (N_17118,N_13187,N_15663);
or U17119 (N_17119,N_14696,N_14973);
nor U17120 (N_17120,N_13121,N_13413);
and U17121 (N_17121,N_12238,N_14682);
nand U17122 (N_17122,N_12901,N_13598);
nand U17123 (N_17123,N_15313,N_15253);
and U17124 (N_17124,N_14200,N_13178);
nand U17125 (N_17125,N_13482,N_14524);
or U17126 (N_17126,N_13838,N_14287);
or U17127 (N_17127,N_15503,N_12655);
xor U17128 (N_17128,N_13875,N_15840);
or U17129 (N_17129,N_13630,N_13061);
and U17130 (N_17130,N_14157,N_13648);
or U17131 (N_17131,N_15843,N_12096);
and U17132 (N_17132,N_13520,N_12813);
nand U17133 (N_17133,N_14415,N_15641);
nand U17134 (N_17134,N_12586,N_14955);
nand U17135 (N_17135,N_15153,N_14260);
nand U17136 (N_17136,N_14025,N_12212);
or U17137 (N_17137,N_13044,N_15877);
nand U17138 (N_17138,N_15600,N_13329);
and U17139 (N_17139,N_13364,N_12508);
and U17140 (N_17140,N_15962,N_14522);
nand U17141 (N_17141,N_12223,N_13367);
nand U17142 (N_17142,N_13177,N_13312);
nand U17143 (N_17143,N_15335,N_15160);
and U17144 (N_17144,N_13502,N_14717);
or U17145 (N_17145,N_15120,N_13528);
or U17146 (N_17146,N_14850,N_14279);
and U17147 (N_17147,N_13167,N_15384);
xor U17148 (N_17148,N_15575,N_13048);
and U17149 (N_17149,N_14975,N_12798);
nand U17150 (N_17150,N_15509,N_12499);
nor U17151 (N_17151,N_12984,N_15667);
and U17152 (N_17152,N_14499,N_15080);
or U17153 (N_17153,N_12872,N_15698);
or U17154 (N_17154,N_12562,N_13360);
and U17155 (N_17155,N_13216,N_15193);
nand U17156 (N_17156,N_15437,N_12688);
or U17157 (N_17157,N_15096,N_13572);
nor U17158 (N_17158,N_15233,N_12645);
nor U17159 (N_17159,N_15936,N_14777);
or U17160 (N_17160,N_14179,N_14460);
or U17161 (N_17161,N_14954,N_13343);
and U17162 (N_17162,N_13283,N_14361);
or U17163 (N_17163,N_13058,N_13306);
and U17164 (N_17164,N_13015,N_15932);
nand U17165 (N_17165,N_12942,N_15866);
and U17166 (N_17166,N_13447,N_13863);
and U17167 (N_17167,N_13460,N_14180);
and U17168 (N_17168,N_13296,N_15688);
or U17169 (N_17169,N_15323,N_13414);
and U17170 (N_17170,N_15634,N_14312);
nor U17171 (N_17171,N_15067,N_15039);
nor U17172 (N_17172,N_12693,N_14171);
nand U17173 (N_17173,N_13691,N_14483);
nand U17174 (N_17174,N_14667,N_12656);
nor U17175 (N_17175,N_13305,N_14362);
and U17176 (N_17176,N_12251,N_12876);
nand U17177 (N_17177,N_12388,N_14660);
nor U17178 (N_17178,N_15861,N_15829);
nor U17179 (N_17179,N_13947,N_12867);
or U17180 (N_17180,N_12408,N_14078);
and U17181 (N_17181,N_14750,N_12282);
nor U17182 (N_17182,N_13053,N_14711);
or U17183 (N_17183,N_12958,N_12061);
nand U17184 (N_17184,N_14775,N_12044);
nor U17185 (N_17185,N_12908,N_13683);
and U17186 (N_17186,N_13155,N_15713);
and U17187 (N_17187,N_13148,N_14981);
and U17188 (N_17188,N_14173,N_13304);
and U17189 (N_17189,N_14659,N_12965);
and U17190 (N_17190,N_15356,N_14860);
or U17191 (N_17191,N_14174,N_12786);
nor U17192 (N_17192,N_13744,N_13023);
nor U17193 (N_17193,N_14398,N_15249);
and U17194 (N_17194,N_13632,N_15395);
or U17195 (N_17195,N_15206,N_13196);
xnor U17196 (N_17196,N_13766,N_15847);
and U17197 (N_17197,N_13813,N_15315);
nand U17198 (N_17198,N_13994,N_15370);
nor U17199 (N_17199,N_15194,N_14946);
nand U17200 (N_17200,N_14080,N_15529);
nor U17201 (N_17201,N_12290,N_12026);
and U17202 (N_17202,N_14116,N_15248);
nor U17203 (N_17203,N_13313,N_14950);
and U17204 (N_17204,N_15346,N_13192);
or U17205 (N_17205,N_13285,N_13890);
and U17206 (N_17206,N_14087,N_14693);
nor U17207 (N_17207,N_12241,N_14389);
or U17208 (N_17208,N_14112,N_14043);
or U17209 (N_17209,N_13827,N_14770);
nand U17210 (N_17210,N_13672,N_13623);
nor U17211 (N_17211,N_13816,N_12437);
xnor U17212 (N_17212,N_15950,N_15873);
and U17213 (N_17213,N_14402,N_15637);
and U17214 (N_17214,N_15849,N_13162);
nand U17215 (N_17215,N_15345,N_14857);
or U17216 (N_17216,N_15816,N_15227);
nand U17217 (N_17217,N_12761,N_15142);
nor U17218 (N_17218,N_14655,N_13483);
nor U17219 (N_17219,N_13857,N_12764);
nand U17220 (N_17220,N_14297,N_12360);
or U17221 (N_17221,N_15859,N_12817);
or U17222 (N_17222,N_12470,N_14721);
and U17223 (N_17223,N_14467,N_15999);
nor U17224 (N_17224,N_14537,N_15443);
nor U17225 (N_17225,N_15042,N_14003);
nand U17226 (N_17226,N_15001,N_12604);
and U17227 (N_17227,N_13933,N_12317);
nor U17228 (N_17228,N_14749,N_13437);
nor U17229 (N_17229,N_15974,N_12843);
nor U17230 (N_17230,N_14780,N_14133);
nand U17231 (N_17231,N_14344,N_12297);
nor U17232 (N_17232,N_12886,N_13912);
nand U17233 (N_17233,N_12312,N_14231);
nand U17234 (N_17234,N_12674,N_13620);
or U17235 (N_17235,N_12863,N_12032);
and U17236 (N_17236,N_14282,N_12743);
or U17237 (N_17237,N_14149,N_15244);
or U17238 (N_17238,N_14574,N_15671);
nand U17239 (N_17239,N_14937,N_13462);
and U17240 (N_17240,N_13342,N_14874);
and U17241 (N_17241,N_12071,N_12545);
and U17242 (N_17242,N_13707,N_14921);
or U17243 (N_17243,N_14588,N_13830);
or U17244 (N_17244,N_14676,N_14793);
or U17245 (N_17245,N_14949,N_14763);
nand U17246 (N_17246,N_13107,N_13239);
nor U17247 (N_17247,N_13020,N_14859);
nor U17248 (N_17248,N_14267,N_12979);
nor U17249 (N_17249,N_15872,N_13407);
nor U17250 (N_17250,N_12667,N_14773);
nand U17251 (N_17251,N_12362,N_13957);
or U17252 (N_17252,N_12797,N_13030);
and U17253 (N_17253,N_12531,N_15219);
and U17254 (N_17254,N_14896,N_15912);
nor U17255 (N_17255,N_15255,N_13350);
and U17256 (N_17256,N_12121,N_15906);
or U17257 (N_17257,N_14885,N_13562);
and U17258 (N_17258,N_12915,N_14979);
nor U17259 (N_17259,N_13302,N_13975);
nor U17260 (N_17260,N_14088,N_15013);
or U17261 (N_17261,N_14546,N_12055);
nor U17262 (N_17262,N_15419,N_15289);
nor U17263 (N_17263,N_14233,N_15549);
nand U17264 (N_17264,N_12787,N_12944);
nor U17265 (N_17265,N_13100,N_14972);
or U17266 (N_17266,N_14005,N_14602);
nand U17267 (N_17267,N_15857,N_12801);
nand U17268 (N_17268,N_15579,N_15508);
nor U17269 (N_17269,N_12889,N_12043);
nor U17270 (N_17270,N_15242,N_15229);
nand U17271 (N_17271,N_14724,N_14961);
nor U17272 (N_17272,N_15454,N_14922);
nand U17273 (N_17273,N_14557,N_12326);
nor U17274 (N_17274,N_12615,N_14705);
and U17275 (N_17275,N_15825,N_15445);
and U17276 (N_17276,N_15502,N_13002);
and U17277 (N_17277,N_13521,N_13228);
nor U17278 (N_17278,N_14774,N_12614);
or U17279 (N_17279,N_13783,N_13670);
or U17280 (N_17280,N_15963,N_14758);
and U17281 (N_17281,N_15734,N_13934);
xnor U17282 (N_17282,N_12058,N_14866);
nor U17283 (N_17283,N_12514,N_15134);
nand U17284 (N_17284,N_15782,N_12625);
nor U17285 (N_17285,N_12685,N_14381);
and U17286 (N_17286,N_14713,N_13823);
nor U17287 (N_17287,N_14832,N_14115);
nor U17288 (N_17288,N_14947,N_15218);
and U17289 (N_17289,N_12695,N_15366);
or U17290 (N_17290,N_13208,N_13475);
nand U17291 (N_17291,N_14306,N_13004);
or U17292 (N_17292,N_15254,N_13825);
and U17293 (N_17293,N_14564,N_15664);
nor U17294 (N_17294,N_13777,N_14649);
nor U17295 (N_17295,N_13787,N_12996);
and U17296 (N_17296,N_14598,N_14094);
nand U17297 (N_17297,N_12961,N_14608);
nor U17298 (N_17298,N_13146,N_15329);
nor U17299 (N_17299,N_14341,N_13338);
or U17300 (N_17300,N_14299,N_12305);
or U17301 (N_17301,N_14813,N_14658);
nand U17302 (N_17302,N_12316,N_15802);
nor U17303 (N_17303,N_12325,N_15391);
or U17304 (N_17304,N_12658,N_15187);
nor U17305 (N_17305,N_15344,N_12240);
and U17306 (N_17306,N_13000,N_15043);
or U17307 (N_17307,N_12382,N_15626);
and U17308 (N_17308,N_13626,N_12184);
or U17309 (N_17309,N_15876,N_12083);
and U17310 (N_17310,N_14943,N_13235);
or U17311 (N_17311,N_15627,N_13066);
nor U17312 (N_17312,N_15625,N_12401);
xor U17313 (N_17313,N_13577,N_14722);
or U17314 (N_17314,N_12430,N_13615);
nand U17315 (N_17315,N_13993,N_13908);
or U17316 (N_17316,N_13566,N_13992);
nand U17317 (N_17317,N_13686,N_13893);
or U17318 (N_17318,N_14698,N_12363);
or U17319 (N_17319,N_12244,N_13668);
or U17320 (N_17320,N_12660,N_14582);
nor U17321 (N_17321,N_15124,N_12540);
nor U17322 (N_17322,N_14829,N_13569);
and U17323 (N_17323,N_14397,N_13355);
or U17324 (N_17324,N_15034,N_12744);
and U17325 (N_17325,N_13935,N_14578);
and U17326 (N_17326,N_12431,N_13804);
nor U17327 (N_17327,N_14571,N_12994);
and U17328 (N_17328,N_13571,N_12461);
nand U17329 (N_17329,N_14597,N_12396);
or U17330 (N_17330,N_12598,N_12284);
nor U17331 (N_17331,N_13604,N_14687);
and U17332 (N_17332,N_12687,N_15581);
nand U17333 (N_17333,N_15633,N_14604);
nor U17334 (N_17334,N_13380,N_14514);
nand U17335 (N_17335,N_12812,N_13700);
or U17336 (N_17336,N_15141,N_12451);
and U17337 (N_17337,N_12466,N_13910);
or U17338 (N_17338,N_12103,N_13851);
and U17339 (N_17339,N_12571,N_13348);
or U17340 (N_17340,N_13202,N_14118);
and U17341 (N_17341,N_14679,N_15166);
and U17342 (N_17342,N_13086,N_12903);
nor U17343 (N_17343,N_12516,N_14045);
nor U17344 (N_17344,N_13062,N_12214);
or U17345 (N_17345,N_13888,N_12762);
nand U17346 (N_17346,N_15271,N_12144);
or U17347 (N_17347,N_15854,N_13468);
nor U17348 (N_17348,N_12410,N_15472);
and U17349 (N_17349,N_15520,N_13389);
or U17350 (N_17350,N_13727,N_14268);
or U17351 (N_17351,N_12529,N_15444);
nor U17352 (N_17352,N_15732,N_12493);
and U17353 (N_17353,N_14369,N_15805);
and U17354 (N_17354,N_15200,N_15197);
or U17355 (N_17355,N_15710,N_14699);
or U17356 (N_17356,N_14716,N_12621);
nand U17357 (N_17357,N_14627,N_14161);
or U17358 (N_17358,N_13833,N_12391);
or U17359 (N_17359,N_14253,N_14600);
or U17360 (N_17360,N_12345,N_15570);
nand U17361 (N_17361,N_13806,N_13925);
nand U17362 (N_17362,N_12407,N_12387);
nand U17363 (N_17363,N_13950,N_12159);
nand U17364 (N_17364,N_13446,N_13977);
or U17365 (N_17365,N_15012,N_13854);
or U17366 (N_17366,N_13169,N_14635);
nand U17367 (N_17367,N_12155,N_14735);
nand U17368 (N_17368,N_13390,N_14120);
and U17369 (N_17369,N_15904,N_12081);
and U17370 (N_17370,N_14990,N_13288);
and U17371 (N_17371,N_13393,N_15035);
nor U17372 (N_17372,N_12597,N_15959);
nand U17373 (N_17373,N_15449,N_13647);
nor U17374 (N_17374,N_12277,N_12926);
and U17375 (N_17375,N_15409,N_15584);
xor U17376 (N_17376,N_14352,N_15337);
and U17377 (N_17377,N_12142,N_15061);
or U17378 (N_17378,N_13386,N_15665);
and U17379 (N_17379,N_13344,N_14004);
nor U17380 (N_17380,N_13262,N_15530);
nand U17381 (N_17381,N_12442,N_12705);
nor U17382 (N_17382,N_12384,N_14761);
or U17383 (N_17383,N_15629,N_13819);
or U17384 (N_17384,N_12480,N_13852);
or U17385 (N_17385,N_13280,N_15191);
or U17386 (N_17386,N_14778,N_13150);
nand U17387 (N_17387,N_12350,N_15214);
nor U17388 (N_17388,N_14965,N_13982);
nor U17389 (N_17389,N_12169,N_13549);
and U17390 (N_17390,N_15719,N_13887);
and U17391 (N_17391,N_15674,N_12222);
or U17392 (N_17392,N_13687,N_13368);
nor U17393 (N_17393,N_14421,N_14155);
or U17394 (N_17394,N_12578,N_12315);
and U17395 (N_17395,N_15613,N_13952);
nor U17396 (N_17396,N_12953,N_13172);
and U17397 (N_17397,N_14633,N_12896);
and U17398 (N_17398,N_12118,N_12146);
nand U17399 (N_17399,N_15136,N_15867);
nor U17400 (N_17400,N_15831,N_12993);
nand U17401 (N_17401,N_15521,N_13723);
or U17402 (N_17402,N_13861,N_12785);
nor U17403 (N_17403,N_15438,N_14358);
or U17404 (N_17404,N_12651,N_13763);
nand U17405 (N_17405,N_12715,N_14052);
or U17406 (N_17406,N_13621,N_15371);
nand U17407 (N_17407,N_15817,N_14932);
nor U17408 (N_17408,N_15815,N_12192);
nand U17409 (N_17409,N_15921,N_14343);
and U17410 (N_17410,N_13484,N_13948);
nand U17411 (N_17411,N_14041,N_15611);
nand U17412 (N_17412,N_12773,N_12140);
nor U17413 (N_17413,N_15198,N_14523);
nand U17414 (N_17414,N_12848,N_13269);
nand U17415 (N_17415,N_12828,N_13088);
and U17416 (N_17416,N_12283,N_12161);
and U17417 (N_17417,N_14662,N_12380);
nor U17418 (N_17418,N_12631,N_13931);
nand U17419 (N_17419,N_14378,N_13011);
and U17420 (N_17420,N_12728,N_13147);
and U17421 (N_17421,N_14728,N_13132);
nand U17422 (N_17422,N_12115,N_14134);
nand U17423 (N_17423,N_15576,N_14997);
and U17424 (N_17424,N_12116,N_15836);
or U17425 (N_17425,N_14395,N_13455);
or U17426 (N_17426,N_13391,N_14206);
or U17427 (N_17427,N_14092,N_12811);
nor U17428 (N_17428,N_12765,N_13529);
nor U17429 (N_17429,N_12644,N_13862);
or U17430 (N_17430,N_15011,N_12855);
and U17431 (N_17431,N_13643,N_13605);
and U17432 (N_17432,N_12669,N_12065);
nand U17433 (N_17433,N_15469,N_13255);
and U17434 (N_17434,N_13937,N_14824);
and U17435 (N_17435,N_13022,N_13122);
and U17436 (N_17436,N_14720,N_15144);
nand U17437 (N_17437,N_13089,N_12756);
and U17438 (N_17438,N_13545,N_13793);
nand U17439 (N_17439,N_13704,N_15165);
xnor U17440 (N_17440,N_15528,N_13070);
nand U17441 (N_17441,N_15195,N_15351);
and U17442 (N_17442,N_14587,N_12007);
and U17443 (N_17443,N_15072,N_15418);
nand U17444 (N_17444,N_15880,N_12673);
and U17445 (N_17445,N_12931,N_14453);
or U17446 (N_17446,N_13607,N_13103);
or U17447 (N_17447,N_12638,N_13991);
nor U17448 (N_17448,N_12288,N_15287);
nand U17449 (N_17449,N_15864,N_13019);
and U17450 (N_17450,N_13336,N_12616);
nand U17451 (N_17451,N_14967,N_15654);
or U17452 (N_17452,N_15874,N_13119);
or U17453 (N_17453,N_15517,N_13807);
nor U17454 (N_17454,N_15051,N_13996);
nor U17455 (N_17455,N_15555,N_14256);
and U17456 (N_17456,N_14023,N_14033);
nor U17457 (N_17457,N_15146,N_15290);
nand U17458 (N_17458,N_15735,N_13008);
or U17459 (N_17459,N_15887,N_12934);
xnor U17460 (N_17460,N_14236,N_15661);
or U17461 (N_17461,N_14346,N_13102);
nand U17462 (N_17462,N_12253,N_13036);
nand U17463 (N_17463,N_15316,N_15567);
nor U17464 (N_17464,N_14186,N_13734);
and U17465 (N_17465,N_14819,N_13403);
or U17466 (N_17466,N_14794,N_14059);
and U17467 (N_17467,N_12703,N_13946);
nand U17468 (N_17468,N_13617,N_12395);
nand U17469 (N_17469,N_15176,N_12361);
nor U17470 (N_17470,N_14263,N_13922);
and U17471 (N_17471,N_13834,N_15208);
nand U17472 (N_17472,N_13039,N_13144);
or U17473 (N_17473,N_13300,N_13151);
or U17474 (N_17474,N_13191,N_15834);
or U17475 (N_17475,N_14366,N_12541);
and U17476 (N_17476,N_13224,N_14783);
nand U17477 (N_17477,N_14912,N_12955);
and U17478 (N_17478,N_15571,N_13041);
nor U17479 (N_17479,N_14691,N_14998);
or U17480 (N_17480,N_13667,N_14882);
nor U17481 (N_17481,N_12859,N_12271);
and U17482 (N_17482,N_15787,N_15821);
or U17483 (N_17483,N_12974,N_14010);
or U17484 (N_17484,N_14840,N_15487);
and U17485 (N_17485,N_12478,N_12775);
nor U17486 (N_17486,N_14894,N_14944);
or U17487 (N_17487,N_15285,N_13826);
or U17488 (N_17488,N_13671,N_13105);
nand U17489 (N_17489,N_14715,N_14781);
xor U17490 (N_17490,N_14881,N_12724);
nand U17491 (N_17491,N_13114,N_12063);
nor U17492 (N_17492,N_14234,N_13864);
and U17493 (N_17493,N_15666,N_12802);
nand U17494 (N_17494,N_14601,N_14516);
or U17495 (N_17495,N_12707,N_15004);
and U17496 (N_17496,N_12907,N_12772);
nand U17497 (N_17497,N_13669,N_15744);
nand U17498 (N_17498,N_13949,N_15398);
nor U17499 (N_17499,N_15262,N_13661);
and U17500 (N_17500,N_13363,N_12373);
and U17501 (N_17501,N_13333,N_12607);
nand U17502 (N_17502,N_12839,N_15979);
nor U17503 (N_17503,N_13253,N_12050);
nor U17504 (N_17504,N_14748,N_12302);
nor U17505 (N_17505,N_13309,N_12768);
or U17506 (N_17506,N_14190,N_14916);
nor U17507 (N_17507,N_14917,N_14061);
nor U17508 (N_17508,N_13516,N_15655);
nand U17509 (N_17509,N_15989,N_15848);
or U17510 (N_17510,N_14273,N_13238);
nor U17511 (N_17511,N_15590,N_15726);
nand U17512 (N_17512,N_14579,N_15630);
nor U17513 (N_17513,N_13354,N_14703);
nor U17514 (N_17514,N_15352,N_15996);
nand U17515 (N_17515,N_14013,N_15170);
nand U17516 (N_17516,N_13796,N_15770);
nor U17517 (N_17517,N_15239,N_12234);
and U17518 (N_17518,N_15328,N_14028);
and U17519 (N_17519,N_12832,N_12069);
nor U17520 (N_17520,N_13759,N_12559);
xor U17521 (N_17521,N_13776,N_14671);
nand U17522 (N_17522,N_13425,N_12490);
nand U17523 (N_17523,N_14624,N_12885);
nand U17524 (N_17524,N_15108,N_14377);
nand U17525 (N_17525,N_14440,N_15978);
and U17526 (N_17526,N_14034,N_13659);
nor U17527 (N_17527,N_14526,N_14095);
or U17528 (N_17528,N_15717,N_12791);
or U17529 (N_17529,N_15798,N_13346);
nand U17530 (N_17530,N_15424,N_15389);
nor U17531 (N_17531,N_13485,N_13478);
nand U17532 (N_17532,N_14497,N_13057);
nor U17533 (N_17533,N_13298,N_13699);
nand U17534 (N_17534,N_13281,N_15131);
or U17535 (N_17535,N_12390,N_14259);
nor U17536 (N_17536,N_12899,N_15380);
or U17537 (N_17537,N_12941,N_14544);
and U17538 (N_17538,N_12157,N_14625);
and U17539 (N_17539,N_12612,N_12503);
nor U17540 (N_17540,N_12523,N_12457);
nor U17541 (N_17541,N_14811,N_14535);
or U17542 (N_17542,N_13600,N_13709);
or U17543 (N_17543,N_15075,N_14904);
nor U17544 (N_17544,N_13749,N_12208);
nand U17545 (N_17545,N_14044,N_12947);
nand U17546 (N_17546,N_15320,N_12793);
xnor U17547 (N_17547,N_14136,N_15275);
or U17548 (N_17548,N_13400,N_15256);
nand U17549 (N_17549,N_14214,N_14927);
and U17550 (N_17550,N_14798,N_15475);
or U17551 (N_17551,N_13771,N_14898);
or U17552 (N_17552,N_13083,N_13962);
nor U17553 (N_17553,N_15483,N_12295);
nand U17554 (N_17554,N_13790,N_12988);
nor U17555 (N_17555,N_13681,N_13650);
nand U17556 (N_17556,N_15212,N_15281);
and U17557 (N_17557,N_12577,N_12436);
and U17558 (N_17558,N_12329,N_13877);
nor U17559 (N_17559,N_14844,N_15624);
and U17560 (N_17560,N_14540,N_14284);
nand U17561 (N_17561,N_13719,N_15879);
and U17562 (N_17562,N_15977,N_15928);
or U17563 (N_17563,N_13592,N_12618);
and U17564 (N_17564,N_13567,N_12600);
nor U17565 (N_17565,N_15110,N_15006);
or U17566 (N_17566,N_12286,N_14986);
nand U17567 (N_17567,N_14865,N_15135);
and U17568 (N_17568,N_12080,N_12665);
nand U17569 (N_17569,N_12924,N_13431);
nand U17570 (N_17570,N_13552,N_12646);
nor U17571 (N_17571,N_15403,N_15125);
or U17572 (N_17572,N_12024,N_12227);
nor U17573 (N_17573,N_14204,N_14666);
nand U17574 (N_17574,N_14672,N_14209);
nor U17575 (N_17575,N_14396,N_13956);
nor U17576 (N_17576,N_15446,N_13379);
nand U17577 (N_17577,N_12969,N_15060);
or U17578 (N_17578,N_12730,N_15202);
nand U17579 (N_17579,N_14613,N_14053);
nor U17580 (N_17580,N_15790,N_14085);
or U17581 (N_17581,N_13513,N_15998);
or U17582 (N_17582,N_14104,N_12089);
nor U17583 (N_17583,N_13641,N_14318);
nor U17584 (N_17584,N_13024,N_12949);
and U17585 (N_17585,N_15355,N_12371);
nor U17586 (N_17586,N_14407,N_15272);
nor U17587 (N_17587,N_13761,N_12476);
nor U17588 (N_17588,N_15036,N_13748);
nand U17589 (N_17589,N_13505,N_12588);
xnor U17590 (N_17590,N_12296,N_12962);
nor U17591 (N_17591,N_12006,N_13442);
nand U17592 (N_17592,N_12720,N_14517);
and U17593 (N_17593,N_15789,N_15321);
and U17594 (N_17594,N_14237,N_14714);
or U17595 (N_17595,N_13633,N_13401);
or U17596 (N_17596,N_15760,N_13551);
and U17597 (N_17597,N_12352,N_15447);
or U17598 (N_17598,N_15282,N_13579);
and U17599 (N_17599,N_13860,N_13047);
nor U17600 (N_17600,N_13491,N_13139);
nand U17601 (N_17601,N_12365,N_14493);
or U17602 (N_17602,N_15348,N_12777);
nor U17603 (N_17603,N_15602,N_13531);
or U17604 (N_17604,N_15976,N_12754);
and U17605 (N_17605,N_13558,N_12104);
or U17606 (N_17606,N_14408,N_15593);
and U17607 (N_17607,N_14247,N_13284);
nand U17608 (N_17608,N_15183,N_15478);
and U17609 (N_17609,N_13108,N_15547);
nor U17610 (N_17610,N_12139,N_15723);
or U17611 (N_17611,N_13186,N_14616);
or U17612 (N_17612,N_15207,N_12635);
nand U17613 (N_17613,N_14801,N_13856);
or U17614 (N_17614,N_14311,N_12017);
nor U17615 (N_17615,N_15991,N_14468);
nor U17616 (N_17616,N_15727,N_14644);
and U17617 (N_17617,N_13612,N_14779);
nor U17618 (N_17618,N_14709,N_13675);
nand U17619 (N_17619,N_13054,N_12324);
nor U17620 (N_17620,N_12873,N_15369);
nand U17621 (N_17621,N_13526,N_12647);
nor U17622 (N_17622,N_14012,N_12808);
nor U17623 (N_17623,N_13622,N_14647);
nor U17624 (N_17624,N_15123,N_13326);
nor U17625 (N_17625,N_13831,N_14271);
and U17626 (N_17626,N_14507,N_15305);
or U17627 (N_17627,N_14205,N_15259);
nand U17628 (N_17628,N_12572,N_12100);
and U17629 (N_17629,N_14202,N_13398);
or U17630 (N_17630,N_15047,N_13473);
nor U17631 (N_17631,N_14528,N_13980);
nor U17632 (N_17632,N_15967,N_12910);
and U17633 (N_17633,N_15286,N_14760);
or U17634 (N_17634,N_12449,N_15933);
nand U17635 (N_17635,N_14321,N_12189);
nor U17636 (N_17636,N_13951,N_13578);
or U17637 (N_17637,N_13603,N_14240);
nor U17638 (N_17638,N_12582,N_12967);
and U17639 (N_17639,N_13204,N_13303);
nor U17640 (N_17640,N_15326,N_14305);
or U17641 (N_17641,N_15943,N_13166);
or U17642 (N_17642,N_12869,N_15238);
and U17643 (N_17643,N_15832,N_12909);
nor U17644 (N_17644,N_14771,N_15112);
and U17645 (N_17645,N_13762,N_12368);
nand U17646 (N_17646,N_13574,N_12441);
or U17647 (N_17647,N_12424,N_12925);
or U17648 (N_17648,N_14474,N_14272);
nand U17649 (N_17649,N_12163,N_13331);
nand U17650 (N_17650,N_14668,N_14764);
nor U17651 (N_17651,N_14951,N_13279);
and U17652 (N_17652,N_14347,N_15027);
and U17653 (N_17653,N_14606,N_12827);
and U17654 (N_17654,N_14680,N_12498);
or U17655 (N_17655,N_13174,N_14296);
nand U17656 (N_17656,N_15722,N_12075);
xor U17657 (N_17657,N_13043,N_12029);
nand U17658 (N_17658,N_15360,N_12162);
nor U17659 (N_17659,N_13915,N_13855);
nor U17660 (N_17660,N_12049,N_14219);
or U17661 (N_17661,N_13385,N_13375);
nor U17662 (N_17662,N_15217,N_14036);
nand U17663 (N_17663,N_15684,N_12426);
or U17664 (N_17664,N_13878,N_14165);
or U17665 (N_17665,N_15496,N_12840);
and U17666 (N_17666,N_15743,N_14639);
nand U17667 (N_17667,N_12182,N_15594);
nor U17668 (N_17668,N_13714,N_13357);
nand U17669 (N_17669,N_14074,N_12771);
and U17670 (N_17670,N_12623,N_13660);
and U17671 (N_17671,N_12620,N_13663);
and U17672 (N_17672,N_13820,N_15673);
nor U17673 (N_17673,N_15331,N_12990);
and U17674 (N_17674,N_14452,N_13945);
nor U17675 (N_17675,N_15766,N_12357);
nand U17676 (N_17676,N_15393,N_15231);
nor U17677 (N_17677,N_13568,N_12190);
or U17678 (N_17678,N_15334,N_13624);
or U17679 (N_17679,N_12000,N_15518);
nand U17680 (N_17680,N_14623,N_15940);
nand U17681 (N_17681,N_15127,N_13637);
nand U17682 (N_17682,N_15955,N_12454);
nor U17683 (N_17683,N_13081,N_13844);
or U17684 (N_17684,N_12042,N_14847);
and U17685 (N_17685,N_13276,N_12747);
and U17686 (N_17686,N_14424,N_15969);
nor U17687 (N_17687,N_12573,N_12299);
and U17688 (N_17688,N_15365,N_12215);
nor U17689 (N_17689,N_13710,N_14925);
nand U17690 (N_17690,N_13078,N_15106);
or U17691 (N_17691,N_12568,N_12591);
nand U17692 (N_17692,N_12725,N_15190);
or U17693 (N_17693,N_14091,N_12303);
or U17694 (N_17694,N_12429,N_14934);
nand U17695 (N_17695,N_13214,N_12298);
nor U17696 (N_17696,N_12168,N_14926);
and U17697 (N_17697,N_13130,N_12517);
nor U17698 (N_17698,N_13388,N_15939);
nor U17699 (N_17699,N_13712,N_14572);
nor U17700 (N_17700,N_13352,N_13250);
and U17701 (N_17701,N_12459,N_13324);
nor U17702 (N_17702,N_15669,N_12031);
and U17703 (N_17703,N_13080,N_14929);
and U17704 (N_17704,N_13646,N_14262);
xnor U17705 (N_17705,N_14870,N_14270);
or U17706 (N_17706,N_14827,N_15065);
nand U17707 (N_17707,N_13016,N_14953);
or U17708 (N_17708,N_13226,N_15327);
nor U17709 (N_17709,N_13334,N_15304);
nand U17710 (N_17710,N_14295,N_15363);
and U17711 (N_17711,N_12940,N_15178);
or U17712 (N_17712,N_12581,N_12987);
or U17713 (N_17713,N_12862,N_15128);
and U17714 (N_17714,N_14737,N_14412);
and U17715 (N_17715,N_14561,N_14420);
and U17716 (N_17716,N_12579,N_12610);
nor U17717 (N_17717,N_14090,N_12682);
nand U17718 (N_17718,N_12082,N_13901);
nand U17719 (N_17719,N_14126,N_15926);
and U17720 (N_17720,N_14208,N_14531);
nor U17721 (N_17721,N_12237,N_12641);
or U17722 (N_17722,N_13467,N_13774);
or U17723 (N_17723,N_15679,N_12174);
nor U17724 (N_17724,N_13297,N_12831);
or U17725 (N_17725,N_15056,N_14286);
and U17726 (N_17726,N_14962,N_13666);
and U17727 (N_17727,N_13444,N_14982);
xor U17728 (N_17728,N_12652,N_15813);
or U17729 (N_17729,N_14592,N_13092);
nand U17730 (N_17730,N_15942,N_14269);
nor U17731 (N_17731,N_13369,N_15388);
or U17732 (N_17732,N_14019,N_14212);
or U17733 (N_17733,N_15824,N_15777);
and U17734 (N_17734,N_13953,N_14001);
nand U17735 (N_17735,N_15185,N_15680);
nor U17736 (N_17736,N_14887,N_13077);
or U17737 (N_17737,N_12052,N_15276);
nor U17738 (N_17738,N_13301,N_15541);
nand U17739 (N_17739,N_13930,N_15157);
nor U17740 (N_17740,N_15934,N_13046);
and U17741 (N_17741,N_12366,N_14797);
xnor U17742 (N_17742,N_15088,N_13866);
nor U17743 (N_17743,N_12445,N_12741);
nand U17744 (N_17744,N_14446,N_15032);
nand U17745 (N_17745,N_14736,N_12458);
nand U17746 (N_17746,N_13110,N_13094);
and U17747 (N_17747,N_15485,N_12956);
or U17748 (N_17748,N_14784,N_14168);
and U17749 (N_17749,N_12760,N_15580);
nand U17750 (N_17750,N_13772,N_15484);
nand U17751 (N_17751,N_12932,N_12716);
or U17752 (N_17752,N_14224,N_12003);
nor U17753 (N_17753,N_14196,N_13037);
or U17754 (N_17754,N_13909,N_15094);
and U17755 (N_17755,N_14871,N_12092);
nor U17756 (N_17756,N_12078,N_13534);
nor U17757 (N_17757,N_12228,N_12327);
and U17758 (N_17758,N_14878,N_15411);
or U17759 (N_17759,N_14158,N_15461);
or U17760 (N_17760,N_15598,N_14425);
and U17761 (N_17761,N_14663,N_14675);
and U17762 (N_17762,N_15122,N_14620);
nor U17763 (N_17763,N_12524,N_13246);
nand U17764 (N_17764,N_15107,N_12099);
nand U17765 (N_17765,N_15982,N_15404);
and U17766 (N_17766,N_15295,N_13894);
or U17767 (N_17767,N_14266,N_14160);
nor U17768 (N_17768,N_15644,N_15470);
or U17769 (N_17769,N_14030,N_14084);
nand U17770 (N_17770,N_14804,N_13565);
nor U17771 (N_17771,N_14692,N_14135);
nand U17772 (N_17772,N_13678,N_12210);
nor U17773 (N_17773,N_13299,N_14319);
and U17774 (N_17774,N_14999,N_15869);
and U17775 (N_17775,N_15771,N_15410);
and U17776 (N_17776,N_12704,N_15209);
nand U17777 (N_17777,N_12870,N_15965);
xnor U17778 (N_17778,N_14067,N_15577);
and U17779 (N_17779,N_13408,N_13205);
nor U17780 (N_17780,N_15312,N_12737);
nand U17781 (N_17781,N_14246,N_13696);
and U17782 (N_17782,N_14261,N_15138);
or U17783 (N_17783,N_12484,N_14814);
and U17784 (N_17784,N_15947,N_12784);
or U17785 (N_17785,N_12179,N_14509);
nand U17786 (N_17786,N_15731,N_13009);
or U17787 (N_17787,N_14146,N_14562);
and U17788 (N_17788,N_14148,N_13330);
nand U17789 (N_17789,N_14674,N_14076);
nand U17790 (N_17790,N_15852,N_12804);
nand U17791 (N_17791,N_13788,N_12782);
nor U17792 (N_17792,N_13924,N_12710);
nor U17793 (N_17793,N_12895,N_12981);
nand U17794 (N_17794,N_14360,N_14227);
nor U17795 (N_17795,N_15587,N_14401);
and U17796 (N_17796,N_14176,N_14449);
nand U17797 (N_17797,N_14451,N_15980);
nor U17798 (N_17798,N_12836,N_15724);
nor U17799 (N_17799,N_15646,N_14469);
nor U17800 (N_17800,N_13332,N_12415);
nor U17801 (N_17801,N_13055,N_13618);
and U17802 (N_17802,N_14942,N_12789);
and U17803 (N_17803,N_13268,N_15154);
and U17804 (N_17804,N_13708,N_14534);
or U17805 (N_17805,N_12535,N_15803);
and U17806 (N_17806,N_13433,N_15311);
and U17807 (N_17807,N_15924,N_14252);
nand U17808 (N_17808,N_12783,N_15755);
nor U17809 (N_17809,N_12211,N_15246);
and U17810 (N_17810,N_12528,N_15850);
nand U17811 (N_17811,N_15028,N_15752);
or U17812 (N_17812,N_15361,N_12733);
nor U17813 (N_17813,N_15071,N_12852);
nand U17814 (N_17814,N_15150,N_14337);
and U17815 (N_17815,N_15756,N_15809);
or U17816 (N_17816,N_14521,N_14140);
or U17817 (N_17817,N_14661,N_14409);
or U17818 (N_17818,N_12405,N_14367);
nand U17819 (N_17819,N_12847,N_12193);
nor U17820 (N_17820,N_12842,N_13049);
or U17821 (N_17821,N_15109,N_15603);
and U17822 (N_17822,N_14945,N_14958);
nor U17823 (N_17823,N_15740,N_13472);
nand U17824 (N_17824,N_12778,N_12954);
or U17825 (N_17825,N_13069,N_14825);
nor U17826 (N_17826,N_12314,N_15909);
nor U17827 (N_17827,N_15931,N_14472);
nor U17828 (N_17828,N_15401,N_12670);
and U17829 (N_17829,N_15486,N_14769);
nand U17830 (N_17830,N_13181,N_12500);
nand U17831 (N_17831,N_14734,N_14851);
or U17832 (N_17832,N_14653,N_15995);
and U17833 (N_17833,N_15616,N_13767);
and U17834 (N_17834,N_12936,N_13677);
or U17835 (N_17835,N_12346,N_15407);
and U17836 (N_17836,N_14879,N_13458);
nor U17837 (N_17837,N_13242,N_14520);
nand U17838 (N_17838,N_12236,N_12287);
nor U17839 (N_17839,N_13498,N_13424);
nand U17840 (N_17840,N_14985,N_14729);
nand U17841 (N_17841,N_13090,N_14441);
nor U17842 (N_17842,N_13028,N_12106);
or U17843 (N_17843,N_15820,N_14688);
or U17844 (N_17844,N_12344,N_14185);
nand U17845 (N_17845,N_14891,N_13370);
nand U17846 (N_17846,N_15171,N_13405);
and U17847 (N_17847,N_12923,N_15860);
nand U17848 (N_17848,N_13752,N_15121);
and U17849 (N_17849,N_15736,N_14443);
or U17850 (N_17850,N_13153,N_12928);
nand U17851 (N_17851,N_14690,N_13021);
and U17852 (N_17852,N_13751,N_12776);
nor U17853 (N_17853,N_14843,N_12727);
nand U17854 (N_17854,N_12224,N_15767);
nor U17855 (N_17855,N_14586,N_12501);
or U17856 (N_17856,N_13142,N_15522);
nand U17857 (N_17857,N_15915,N_13323);
and U17858 (N_17858,N_15412,N_14560);
nor U17859 (N_17859,N_13134,N_14351);
nor U17860 (N_17860,N_13286,N_13533);
or U17861 (N_17861,N_13432,N_13347);
and U17862 (N_17862,N_14383,N_14900);
and U17863 (N_17863,N_15791,N_12968);
and U17864 (N_17864,N_13871,N_12209);
and U17865 (N_17865,N_12151,N_13639);
nor U17866 (N_17866,N_13614,N_13327);
and U17867 (N_17867,N_13782,N_12835);
xnor U17868 (N_17868,N_13158,N_14439);
nand U17869 (N_17869,N_15908,N_14726);
nor U17870 (N_17870,N_12173,N_14909);
and U17871 (N_17871,N_15774,N_14159);
nand U17872 (N_17872,N_12072,N_14806);
nand U17873 (N_17873,N_14645,N_13510);
nand U17874 (N_17874,N_14948,N_12076);
nand U17875 (N_17875,N_14294,N_12985);
or U17876 (N_17876,N_14792,N_15269);
or U17877 (N_17877,N_15163,N_14046);
or U17878 (N_17878,N_12131,N_12294);
nand U17879 (N_17879,N_12860,N_14464);
nor U17880 (N_17880,N_13410,N_14838);
or U17881 (N_17881,N_13418,N_14073);
or U17882 (N_17882,N_13068,N_13743);
and U17883 (N_17883,N_12393,N_14686);
nand U17884 (N_17884,N_12206,N_15761);
or U17885 (N_17885,N_13715,N_12883);
nand U17886 (N_17886,N_13109,N_14519);
nand U17887 (N_17887,N_13588,N_12456);
nand U17888 (N_17888,N_15811,N_13270);
and U17889 (N_17889,N_15762,N_14489);
nor U17890 (N_17890,N_15133,N_12569);
nor U17891 (N_17891,N_14611,N_15501);
nand U17892 (N_17892,N_12815,N_15608);
or U17893 (N_17893,N_12385,N_13556);
nor U17894 (N_17894,N_15415,N_12376);
or U17895 (N_17895,N_13194,N_14175);
nand U17896 (N_17896,N_12175,N_15583);
nor U17897 (N_17897,N_13803,N_15514);
nor U17898 (N_17898,N_15137,N_12520);
or U17899 (N_17899,N_15095,N_12242);
nor U17900 (N_17900,N_13290,N_13998);
or U17901 (N_17901,N_15049,N_12714);
nand U17902 (N_17902,N_15396,N_13486);
nor U17903 (N_17903,N_15556,N_15098);
nor U17904 (N_17904,N_15432,N_13254);
nor U17905 (N_17905,N_12091,N_15745);
or U17906 (N_17906,N_12678,N_14547);
or U17907 (N_17907,N_14549,N_15951);
nand U17908 (N_17908,N_13755,N_13874);
nor U17909 (N_17909,N_13159,N_12538);
and U17910 (N_17910,N_14264,N_15729);
nor U17911 (N_17911,N_13143,N_12810);
or U17912 (N_17912,N_13680,N_15357);
and U17913 (N_17913,N_14708,N_12689);
and U17914 (N_17914,N_14941,N_14213);
or U17915 (N_17915,N_14553,N_15714);
or U17916 (N_17916,N_15377,N_15498);
nor U17917 (N_17917,N_12117,N_13320);
nor U17918 (N_17918,N_14618,N_15599);
nor U17919 (N_17919,N_14182,N_13791);
or U17920 (N_17920,N_13025,N_14888);
nand U17921 (N_17921,N_14484,N_13145);
or U17922 (N_17922,N_14258,N_15540);
and U17923 (N_17923,N_15538,N_15213);
nor U17924 (N_17924,N_12152,N_14332);
nand U17925 (N_17925,N_14648,N_14162);
nor U17926 (N_17926,N_14245,N_13973);
or U17927 (N_17927,N_15169,N_15018);
and U17928 (N_17928,N_15759,N_14584);
nor U17929 (N_17929,N_15314,N_13904);
nand U17930 (N_17930,N_14707,N_12124);
nor U17931 (N_17931,N_13542,N_14277);
nand U17932 (N_17932,N_12004,N_15280);
nand U17933 (N_17933,N_15045,N_15199);
nor U17934 (N_17934,N_12684,N_13698);
nor U17935 (N_17935,N_14656,N_15957);
xor U17936 (N_17936,N_14939,N_15640);
or U17937 (N_17937,N_14974,N_15466);
nand U17938 (N_17938,N_14191,N_13412);
and U17939 (N_17939,N_15851,N_14848);
nor U17940 (N_17940,N_14228,N_14634);
nor U17941 (N_17941,N_14249,N_12334);
or U17942 (N_17942,N_14027,N_13917);
or U17943 (N_17943,N_13292,N_12736);
or U17944 (N_17944,N_14568,N_14020);
and U17945 (N_17945,N_14163,N_14931);
or U17946 (N_17946,N_14725,N_12347);
nand U17947 (N_17947,N_15059,N_12794);
and U17948 (N_17948,N_13972,N_14372);
nand U17949 (N_17949,N_15460,N_14280);
or U17950 (N_17950,N_12543,N_13920);
nor U17951 (N_17951,N_12536,N_15161);
or U17952 (N_17952,N_13635,N_12483);
nand U17953 (N_17953,N_12239,N_13406);
nand U17954 (N_17954,N_12349,N_15523);
nand U17955 (N_17955,N_14068,N_14854);
or U17956 (N_17956,N_12053,N_13123);
or U17957 (N_17957,N_14628,N_15704);
and U17958 (N_17958,N_12792,N_13960);
and U17959 (N_17959,N_12263,N_13180);
nor U17960 (N_17960,N_13175,N_13555);
or U17961 (N_17961,N_12613,N_12318);
nand U17962 (N_17962,N_14782,N_13967);
xor U17963 (N_17963,N_13711,N_15078);
and U17964 (N_17964,N_13746,N_15052);
or U17965 (N_17965,N_15151,N_12375);
xnor U17966 (N_17966,N_12351,N_12221);
nor U17967 (N_17967,N_13029,N_15548);
and U17968 (N_17968,N_14991,N_12805);
or U17969 (N_17969,N_14818,N_14106);
nand U17970 (N_17970,N_12563,N_14583);
or U17971 (N_17971,N_14539,N_13227);
and U17972 (N_17972,N_12900,N_13976);
nand U17973 (N_17973,N_13221,N_14365);
nor U17974 (N_17974,N_14886,N_15720);
and U17975 (N_17975,N_12766,N_15916);
nand U17976 (N_17976,N_15097,N_14111);
and U17977 (N_17977,N_12662,N_15747);
nand U17978 (N_17978,N_13218,N_13496);
nor U17979 (N_17979,N_13474,N_12377);
or U17980 (N_17980,N_15149,N_14183);
nor U17981 (N_17981,N_14502,N_15268);
or U17982 (N_17982,N_14288,N_15592);
nand U17983 (N_17983,N_15651,N_15797);
or U17984 (N_17984,N_12758,N_14897);
and U17985 (N_17985,N_15340,N_14345);
nand U17986 (N_17986,N_12599,N_14901);
nor U17987 (N_17987,N_15283,N_15588);
nand U17988 (N_17988,N_13760,N_15546);
or U17989 (N_17989,N_13509,N_12549);
or U17990 (N_17990,N_14386,N_14406);
and U17991 (N_17991,N_12398,N_13085);
nor U17992 (N_17992,N_15794,N_13814);
nand U17993 (N_17993,N_14914,N_12894);
and U17994 (N_17994,N_12970,N_15930);
or U17995 (N_17995,N_13310,N_15048);
nand U17996 (N_17996,N_12729,N_12755);
and U17997 (N_17997,N_15017,N_14101);
and U17998 (N_17998,N_15513,N_14338);
or U17999 (N_17999,N_13959,N_12145);
nand U18000 (N_18000,N_12332,N_15318);
nand U18001 (N_18001,N_12395,N_15542);
nand U18002 (N_18002,N_14240,N_12280);
and U18003 (N_18003,N_13864,N_13941);
and U18004 (N_18004,N_15314,N_14376);
or U18005 (N_18005,N_13648,N_14879);
nor U18006 (N_18006,N_12928,N_13857);
nor U18007 (N_18007,N_15396,N_12922);
and U18008 (N_18008,N_13316,N_13875);
or U18009 (N_18009,N_15121,N_13415);
nand U18010 (N_18010,N_15785,N_14533);
nand U18011 (N_18011,N_13093,N_14751);
or U18012 (N_18012,N_13780,N_14386);
nor U18013 (N_18013,N_15084,N_12978);
or U18014 (N_18014,N_15179,N_13138);
or U18015 (N_18015,N_14573,N_13572);
or U18016 (N_18016,N_12196,N_14038);
nor U18017 (N_18017,N_13521,N_13353);
and U18018 (N_18018,N_15185,N_12976);
nand U18019 (N_18019,N_14740,N_12008);
and U18020 (N_18020,N_13614,N_12596);
nand U18021 (N_18021,N_14893,N_14401);
nand U18022 (N_18022,N_14058,N_14396);
and U18023 (N_18023,N_15853,N_12064);
nor U18024 (N_18024,N_15325,N_12735);
nor U18025 (N_18025,N_14018,N_13181);
nor U18026 (N_18026,N_14696,N_12517);
and U18027 (N_18027,N_12563,N_12691);
or U18028 (N_18028,N_13147,N_12077);
nor U18029 (N_18029,N_12598,N_12285);
nor U18030 (N_18030,N_12466,N_12345);
and U18031 (N_18031,N_13565,N_14059);
or U18032 (N_18032,N_13924,N_15910);
nor U18033 (N_18033,N_12366,N_14119);
or U18034 (N_18034,N_12658,N_12800);
or U18035 (N_18035,N_14263,N_12984);
or U18036 (N_18036,N_13852,N_12682);
nor U18037 (N_18037,N_13217,N_14964);
and U18038 (N_18038,N_12482,N_14698);
or U18039 (N_18039,N_15347,N_13006);
or U18040 (N_18040,N_12132,N_12757);
or U18041 (N_18041,N_12794,N_14578);
nor U18042 (N_18042,N_14094,N_14091);
or U18043 (N_18043,N_14839,N_14247);
and U18044 (N_18044,N_13413,N_12332);
nor U18045 (N_18045,N_15520,N_14836);
or U18046 (N_18046,N_13829,N_13262);
nor U18047 (N_18047,N_13721,N_14101);
nand U18048 (N_18048,N_14109,N_14743);
or U18049 (N_18049,N_13116,N_14277);
nor U18050 (N_18050,N_15366,N_13629);
nand U18051 (N_18051,N_13325,N_12672);
or U18052 (N_18052,N_13139,N_13411);
and U18053 (N_18053,N_12811,N_13357);
or U18054 (N_18054,N_12267,N_12464);
nand U18055 (N_18055,N_12939,N_15033);
xor U18056 (N_18056,N_13518,N_14688);
or U18057 (N_18057,N_14866,N_12313);
nor U18058 (N_18058,N_12104,N_14183);
and U18059 (N_18059,N_15331,N_15343);
nor U18060 (N_18060,N_13621,N_15893);
and U18061 (N_18061,N_12620,N_14990);
and U18062 (N_18062,N_12351,N_12469);
or U18063 (N_18063,N_14399,N_12131);
or U18064 (N_18064,N_15584,N_12505);
and U18065 (N_18065,N_15267,N_14507);
and U18066 (N_18066,N_13173,N_14415);
and U18067 (N_18067,N_14355,N_15384);
nor U18068 (N_18068,N_15317,N_15878);
and U18069 (N_18069,N_13705,N_14151);
and U18070 (N_18070,N_15764,N_14681);
nor U18071 (N_18071,N_14452,N_15010);
or U18072 (N_18072,N_13331,N_13880);
nor U18073 (N_18073,N_15708,N_14923);
nor U18074 (N_18074,N_13901,N_13535);
nand U18075 (N_18075,N_12731,N_14277);
nor U18076 (N_18076,N_15065,N_13551);
nor U18077 (N_18077,N_15718,N_14562);
nand U18078 (N_18078,N_14825,N_15092);
and U18079 (N_18079,N_12341,N_15397);
and U18080 (N_18080,N_15760,N_14842);
nor U18081 (N_18081,N_14516,N_14401);
or U18082 (N_18082,N_15402,N_13680);
nor U18083 (N_18083,N_13047,N_12488);
or U18084 (N_18084,N_14010,N_14865);
nand U18085 (N_18085,N_15192,N_14380);
nand U18086 (N_18086,N_14195,N_13087);
nand U18087 (N_18087,N_13661,N_14708);
nor U18088 (N_18088,N_15969,N_13158);
nor U18089 (N_18089,N_13041,N_14600);
nor U18090 (N_18090,N_15679,N_13797);
nor U18091 (N_18091,N_15217,N_14217);
or U18092 (N_18092,N_12729,N_14454);
and U18093 (N_18093,N_13229,N_15051);
or U18094 (N_18094,N_14317,N_12579);
or U18095 (N_18095,N_13198,N_15792);
and U18096 (N_18096,N_14442,N_12468);
nor U18097 (N_18097,N_15779,N_14591);
nor U18098 (N_18098,N_14705,N_12854);
nor U18099 (N_18099,N_12618,N_13289);
nor U18100 (N_18100,N_15207,N_12208);
nand U18101 (N_18101,N_12934,N_13914);
nand U18102 (N_18102,N_12072,N_13319);
and U18103 (N_18103,N_15793,N_14372);
nor U18104 (N_18104,N_15846,N_15824);
and U18105 (N_18105,N_12298,N_12213);
nor U18106 (N_18106,N_12261,N_13533);
and U18107 (N_18107,N_14262,N_14813);
and U18108 (N_18108,N_15138,N_15816);
and U18109 (N_18109,N_13445,N_15002);
and U18110 (N_18110,N_13137,N_15662);
or U18111 (N_18111,N_12711,N_13746);
and U18112 (N_18112,N_13489,N_15004);
nand U18113 (N_18113,N_13974,N_15086);
or U18114 (N_18114,N_14359,N_14303);
and U18115 (N_18115,N_13865,N_14643);
or U18116 (N_18116,N_13937,N_14371);
nor U18117 (N_18117,N_13807,N_13693);
and U18118 (N_18118,N_14598,N_12370);
or U18119 (N_18119,N_14453,N_13772);
or U18120 (N_18120,N_14264,N_15063);
nand U18121 (N_18121,N_15807,N_12232);
and U18122 (N_18122,N_15042,N_12970);
nand U18123 (N_18123,N_14978,N_12187);
nor U18124 (N_18124,N_14251,N_13131);
or U18125 (N_18125,N_14226,N_15527);
and U18126 (N_18126,N_14925,N_14691);
or U18127 (N_18127,N_15964,N_13661);
and U18128 (N_18128,N_13156,N_12328);
nor U18129 (N_18129,N_12030,N_12267);
or U18130 (N_18130,N_13705,N_14002);
and U18131 (N_18131,N_15873,N_14177);
xnor U18132 (N_18132,N_13847,N_13632);
nand U18133 (N_18133,N_15821,N_14533);
or U18134 (N_18134,N_14166,N_14542);
or U18135 (N_18135,N_15358,N_12131);
nor U18136 (N_18136,N_14726,N_13416);
and U18137 (N_18137,N_13558,N_14600);
and U18138 (N_18138,N_15794,N_13981);
nor U18139 (N_18139,N_12727,N_12985);
nand U18140 (N_18140,N_15103,N_15561);
nand U18141 (N_18141,N_15395,N_14271);
nor U18142 (N_18142,N_15581,N_15729);
and U18143 (N_18143,N_15422,N_12324);
and U18144 (N_18144,N_13472,N_12113);
or U18145 (N_18145,N_14970,N_15068);
and U18146 (N_18146,N_15760,N_13043);
and U18147 (N_18147,N_12036,N_12386);
or U18148 (N_18148,N_12061,N_13049);
and U18149 (N_18149,N_12329,N_12583);
nand U18150 (N_18150,N_15884,N_14052);
or U18151 (N_18151,N_13771,N_14330);
and U18152 (N_18152,N_14675,N_13979);
nor U18153 (N_18153,N_13549,N_15899);
nor U18154 (N_18154,N_12785,N_14728);
or U18155 (N_18155,N_12194,N_12589);
nand U18156 (N_18156,N_13260,N_12154);
nand U18157 (N_18157,N_14185,N_14673);
nor U18158 (N_18158,N_12573,N_13145);
or U18159 (N_18159,N_12765,N_13233);
nor U18160 (N_18160,N_15109,N_13114);
or U18161 (N_18161,N_13137,N_14703);
nor U18162 (N_18162,N_15965,N_12419);
nor U18163 (N_18163,N_13177,N_15280);
or U18164 (N_18164,N_12622,N_12471);
nor U18165 (N_18165,N_14918,N_12380);
and U18166 (N_18166,N_12387,N_15289);
and U18167 (N_18167,N_13381,N_12624);
nand U18168 (N_18168,N_14888,N_12747);
xnor U18169 (N_18169,N_14938,N_14436);
nor U18170 (N_18170,N_15210,N_12176);
and U18171 (N_18171,N_13847,N_12163);
and U18172 (N_18172,N_15408,N_12861);
and U18173 (N_18173,N_14234,N_13636);
nor U18174 (N_18174,N_15737,N_14408);
or U18175 (N_18175,N_15293,N_15371);
nor U18176 (N_18176,N_15522,N_15638);
and U18177 (N_18177,N_14410,N_15504);
or U18178 (N_18178,N_15138,N_14042);
or U18179 (N_18179,N_13962,N_13847);
or U18180 (N_18180,N_14030,N_12800);
and U18181 (N_18181,N_12061,N_13152);
and U18182 (N_18182,N_15967,N_14830);
nand U18183 (N_18183,N_14752,N_14109);
nor U18184 (N_18184,N_14679,N_15262);
nor U18185 (N_18185,N_15209,N_14001);
or U18186 (N_18186,N_13571,N_14598);
or U18187 (N_18187,N_14217,N_12646);
or U18188 (N_18188,N_15129,N_14902);
nand U18189 (N_18189,N_14027,N_12341);
nor U18190 (N_18190,N_14913,N_14423);
nand U18191 (N_18191,N_12786,N_14654);
nor U18192 (N_18192,N_12227,N_12961);
and U18193 (N_18193,N_12303,N_13313);
and U18194 (N_18194,N_15565,N_12515);
nor U18195 (N_18195,N_15711,N_14059);
nand U18196 (N_18196,N_12956,N_13284);
and U18197 (N_18197,N_13005,N_13241);
nor U18198 (N_18198,N_13673,N_14031);
nand U18199 (N_18199,N_13432,N_12713);
nand U18200 (N_18200,N_12762,N_14347);
xor U18201 (N_18201,N_12058,N_13891);
and U18202 (N_18202,N_13093,N_14580);
nand U18203 (N_18203,N_15278,N_13328);
or U18204 (N_18204,N_14167,N_14658);
and U18205 (N_18205,N_14301,N_12557);
nand U18206 (N_18206,N_15462,N_15776);
nor U18207 (N_18207,N_15473,N_14188);
nand U18208 (N_18208,N_13918,N_15096);
nand U18209 (N_18209,N_13675,N_13919);
nand U18210 (N_18210,N_15376,N_13865);
nor U18211 (N_18211,N_14095,N_12978);
or U18212 (N_18212,N_14640,N_13400);
nand U18213 (N_18213,N_13682,N_14653);
and U18214 (N_18214,N_12581,N_14991);
and U18215 (N_18215,N_15261,N_15216);
or U18216 (N_18216,N_12061,N_15416);
and U18217 (N_18217,N_12028,N_12330);
or U18218 (N_18218,N_15917,N_13551);
nor U18219 (N_18219,N_15638,N_13685);
nand U18220 (N_18220,N_13266,N_13012);
nand U18221 (N_18221,N_13817,N_14788);
nand U18222 (N_18222,N_12574,N_13678);
nand U18223 (N_18223,N_13653,N_14640);
or U18224 (N_18224,N_12561,N_15607);
or U18225 (N_18225,N_12644,N_12620);
and U18226 (N_18226,N_15869,N_12267);
nand U18227 (N_18227,N_13563,N_15250);
and U18228 (N_18228,N_15077,N_13623);
or U18229 (N_18229,N_15528,N_13240);
or U18230 (N_18230,N_14868,N_12771);
and U18231 (N_18231,N_15778,N_15154);
and U18232 (N_18232,N_12580,N_12803);
nor U18233 (N_18233,N_12928,N_13616);
nand U18234 (N_18234,N_13816,N_15030);
nor U18235 (N_18235,N_13175,N_12653);
or U18236 (N_18236,N_14845,N_12338);
nand U18237 (N_18237,N_15113,N_12596);
nor U18238 (N_18238,N_15844,N_12185);
or U18239 (N_18239,N_13489,N_15336);
nand U18240 (N_18240,N_14033,N_13500);
or U18241 (N_18241,N_15389,N_15332);
and U18242 (N_18242,N_13483,N_13464);
or U18243 (N_18243,N_12915,N_15863);
or U18244 (N_18244,N_14029,N_15805);
nand U18245 (N_18245,N_15530,N_15151);
or U18246 (N_18246,N_12459,N_12821);
nor U18247 (N_18247,N_14148,N_12279);
and U18248 (N_18248,N_13826,N_12858);
nand U18249 (N_18249,N_14605,N_13702);
and U18250 (N_18250,N_14464,N_15636);
nand U18251 (N_18251,N_14555,N_13273);
nand U18252 (N_18252,N_14355,N_15008);
and U18253 (N_18253,N_15727,N_12364);
or U18254 (N_18254,N_15075,N_13945);
and U18255 (N_18255,N_15619,N_12411);
and U18256 (N_18256,N_14439,N_13849);
and U18257 (N_18257,N_12330,N_14138);
and U18258 (N_18258,N_13588,N_14172);
xnor U18259 (N_18259,N_13524,N_12872);
nor U18260 (N_18260,N_13894,N_12416);
or U18261 (N_18261,N_13413,N_12531);
nand U18262 (N_18262,N_15884,N_13779);
and U18263 (N_18263,N_13473,N_13825);
nor U18264 (N_18264,N_13031,N_15797);
or U18265 (N_18265,N_13964,N_12242);
or U18266 (N_18266,N_13631,N_13587);
or U18267 (N_18267,N_13349,N_12941);
and U18268 (N_18268,N_12565,N_15797);
xnor U18269 (N_18269,N_12842,N_12869);
nand U18270 (N_18270,N_13084,N_13090);
or U18271 (N_18271,N_15287,N_13926);
nor U18272 (N_18272,N_13693,N_14260);
or U18273 (N_18273,N_15573,N_14225);
nand U18274 (N_18274,N_15834,N_14601);
and U18275 (N_18275,N_15487,N_15729);
nand U18276 (N_18276,N_12776,N_12685);
nand U18277 (N_18277,N_15481,N_14183);
nand U18278 (N_18278,N_13609,N_15430);
and U18279 (N_18279,N_12456,N_15865);
nand U18280 (N_18280,N_15690,N_14418);
nand U18281 (N_18281,N_14675,N_14319);
and U18282 (N_18282,N_13493,N_12516);
and U18283 (N_18283,N_14243,N_15021);
nand U18284 (N_18284,N_14761,N_15673);
nor U18285 (N_18285,N_15879,N_14065);
nand U18286 (N_18286,N_12424,N_14754);
or U18287 (N_18287,N_15935,N_12363);
or U18288 (N_18288,N_15447,N_15702);
and U18289 (N_18289,N_15687,N_14829);
nor U18290 (N_18290,N_12352,N_13296);
nand U18291 (N_18291,N_14233,N_13678);
and U18292 (N_18292,N_14060,N_15327);
or U18293 (N_18293,N_13909,N_13717);
nor U18294 (N_18294,N_12726,N_13352);
nor U18295 (N_18295,N_13998,N_13180);
nand U18296 (N_18296,N_14729,N_14327);
and U18297 (N_18297,N_12185,N_15570);
xnor U18298 (N_18298,N_13583,N_13775);
nor U18299 (N_18299,N_13956,N_13556);
nand U18300 (N_18300,N_14198,N_12163);
or U18301 (N_18301,N_14251,N_14573);
nor U18302 (N_18302,N_13886,N_12777);
and U18303 (N_18303,N_13681,N_12115);
and U18304 (N_18304,N_13032,N_13649);
nand U18305 (N_18305,N_14442,N_13404);
nand U18306 (N_18306,N_14841,N_13816);
nor U18307 (N_18307,N_15467,N_14484);
and U18308 (N_18308,N_12695,N_13700);
and U18309 (N_18309,N_15171,N_12041);
or U18310 (N_18310,N_15949,N_14681);
or U18311 (N_18311,N_15896,N_14423);
nand U18312 (N_18312,N_12249,N_12501);
or U18313 (N_18313,N_14250,N_14903);
or U18314 (N_18314,N_14840,N_13600);
nand U18315 (N_18315,N_13446,N_13246);
or U18316 (N_18316,N_14832,N_15485);
nor U18317 (N_18317,N_12564,N_14681);
nor U18318 (N_18318,N_13631,N_14628);
or U18319 (N_18319,N_15674,N_13227);
nand U18320 (N_18320,N_15369,N_14600);
and U18321 (N_18321,N_14916,N_13907);
or U18322 (N_18322,N_14540,N_12053);
and U18323 (N_18323,N_15486,N_15073);
nand U18324 (N_18324,N_13941,N_12429);
nand U18325 (N_18325,N_13694,N_12639);
or U18326 (N_18326,N_14393,N_14553);
or U18327 (N_18327,N_13166,N_12829);
or U18328 (N_18328,N_15657,N_15984);
or U18329 (N_18329,N_14206,N_14995);
and U18330 (N_18330,N_14260,N_13937);
or U18331 (N_18331,N_12070,N_13865);
nand U18332 (N_18332,N_14310,N_15412);
or U18333 (N_18333,N_12369,N_15262);
nand U18334 (N_18334,N_14178,N_14303);
or U18335 (N_18335,N_12229,N_15320);
or U18336 (N_18336,N_15025,N_14952);
or U18337 (N_18337,N_15128,N_14555);
nand U18338 (N_18338,N_15545,N_14827);
nand U18339 (N_18339,N_12838,N_15548);
or U18340 (N_18340,N_13021,N_12924);
or U18341 (N_18341,N_14315,N_13422);
nand U18342 (N_18342,N_13343,N_13442);
or U18343 (N_18343,N_15127,N_13849);
nor U18344 (N_18344,N_15693,N_13894);
and U18345 (N_18345,N_12928,N_13087);
and U18346 (N_18346,N_14662,N_14442);
nand U18347 (N_18347,N_12096,N_12866);
and U18348 (N_18348,N_14973,N_14293);
or U18349 (N_18349,N_14203,N_14172);
nand U18350 (N_18350,N_12696,N_13361);
and U18351 (N_18351,N_12397,N_15917);
nor U18352 (N_18352,N_13248,N_13745);
nor U18353 (N_18353,N_15924,N_12881);
or U18354 (N_18354,N_13609,N_13202);
nor U18355 (N_18355,N_14994,N_15867);
and U18356 (N_18356,N_15926,N_14949);
nor U18357 (N_18357,N_12358,N_15163);
nand U18358 (N_18358,N_12360,N_14746);
and U18359 (N_18359,N_12758,N_14557);
or U18360 (N_18360,N_14204,N_13118);
and U18361 (N_18361,N_15878,N_14037);
nor U18362 (N_18362,N_12266,N_14527);
and U18363 (N_18363,N_12414,N_13083);
or U18364 (N_18364,N_13954,N_15410);
and U18365 (N_18365,N_13332,N_13601);
or U18366 (N_18366,N_12630,N_13064);
nand U18367 (N_18367,N_15997,N_15729);
and U18368 (N_18368,N_15975,N_14500);
nand U18369 (N_18369,N_12062,N_15046);
nand U18370 (N_18370,N_15896,N_14548);
nand U18371 (N_18371,N_14679,N_15513);
nor U18372 (N_18372,N_13594,N_13101);
and U18373 (N_18373,N_13853,N_15027);
nor U18374 (N_18374,N_12546,N_15332);
and U18375 (N_18375,N_15541,N_14798);
or U18376 (N_18376,N_14004,N_12345);
nand U18377 (N_18377,N_15348,N_13931);
and U18378 (N_18378,N_14541,N_13228);
nor U18379 (N_18379,N_14442,N_12128);
nand U18380 (N_18380,N_15367,N_13316);
nand U18381 (N_18381,N_14203,N_14476);
and U18382 (N_18382,N_12885,N_14400);
or U18383 (N_18383,N_12762,N_14231);
nor U18384 (N_18384,N_14176,N_13569);
nor U18385 (N_18385,N_12048,N_15182);
and U18386 (N_18386,N_12195,N_14776);
nand U18387 (N_18387,N_14088,N_14231);
and U18388 (N_18388,N_14299,N_13836);
nand U18389 (N_18389,N_14802,N_12444);
nand U18390 (N_18390,N_13591,N_14645);
and U18391 (N_18391,N_13563,N_12739);
or U18392 (N_18392,N_14369,N_12080);
nand U18393 (N_18393,N_14750,N_12709);
or U18394 (N_18394,N_15800,N_12260);
nor U18395 (N_18395,N_13718,N_12876);
or U18396 (N_18396,N_12545,N_13429);
or U18397 (N_18397,N_13609,N_12108);
and U18398 (N_18398,N_12265,N_14348);
nor U18399 (N_18399,N_12274,N_12886);
or U18400 (N_18400,N_15486,N_15435);
and U18401 (N_18401,N_15020,N_13046);
nand U18402 (N_18402,N_14815,N_13747);
and U18403 (N_18403,N_15487,N_14325);
or U18404 (N_18404,N_13046,N_12293);
nor U18405 (N_18405,N_13219,N_14518);
and U18406 (N_18406,N_13192,N_14250);
and U18407 (N_18407,N_15957,N_14645);
or U18408 (N_18408,N_15441,N_15743);
nor U18409 (N_18409,N_12680,N_12681);
nand U18410 (N_18410,N_12882,N_14297);
or U18411 (N_18411,N_13562,N_14288);
or U18412 (N_18412,N_15666,N_13255);
or U18413 (N_18413,N_13219,N_15314);
or U18414 (N_18414,N_12533,N_13849);
nand U18415 (N_18415,N_12012,N_12282);
nor U18416 (N_18416,N_15947,N_15289);
nor U18417 (N_18417,N_15567,N_15835);
nor U18418 (N_18418,N_12271,N_15970);
or U18419 (N_18419,N_12369,N_12697);
nand U18420 (N_18420,N_14642,N_13761);
nor U18421 (N_18421,N_14052,N_12961);
and U18422 (N_18422,N_15566,N_13363);
nor U18423 (N_18423,N_12319,N_12904);
nand U18424 (N_18424,N_12153,N_12344);
or U18425 (N_18425,N_12356,N_15250);
nand U18426 (N_18426,N_12219,N_15662);
and U18427 (N_18427,N_15926,N_15192);
nand U18428 (N_18428,N_12450,N_14583);
and U18429 (N_18429,N_13128,N_13501);
and U18430 (N_18430,N_15981,N_14115);
nand U18431 (N_18431,N_13673,N_15209);
or U18432 (N_18432,N_15751,N_14344);
nor U18433 (N_18433,N_12169,N_15539);
and U18434 (N_18434,N_13565,N_13231);
nand U18435 (N_18435,N_14985,N_14587);
or U18436 (N_18436,N_14266,N_15730);
nor U18437 (N_18437,N_12390,N_15032);
nor U18438 (N_18438,N_15387,N_15865);
or U18439 (N_18439,N_14438,N_15730);
and U18440 (N_18440,N_13935,N_15037);
xnor U18441 (N_18441,N_15142,N_12554);
and U18442 (N_18442,N_12292,N_12740);
or U18443 (N_18443,N_13636,N_13156);
nand U18444 (N_18444,N_12459,N_14124);
nand U18445 (N_18445,N_15461,N_14257);
nand U18446 (N_18446,N_14327,N_12930);
and U18447 (N_18447,N_14700,N_13920);
nor U18448 (N_18448,N_13154,N_15586);
nor U18449 (N_18449,N_14595,N_14224);
or U18450 (N_18450,N_12236,N_12822);
nor U18451 (N_18451,N_12026,N_13980);
or U18452 (N_18452,N_13067,N_13191);
nor U18453 (N_18453,N_14195,N_12364);
or U18454 (N_18454,N_15755,N_12464);
or U18455 (N_18455,N_12591,N_12761);
or U18456 (N_18456,N_12692,N_15474);
and U18457 (N_18457,N_15682,N_13984);
nor U18458 (N_18458,N_15745,N_14449);
nand U18459 (N_18459,N_13992,N_12228);
and U18460 (N_18460,N_14206,N_12984);
nor U18461 (N_18461,N_14791,N_13431);
nand U18462 (N_18462,N_14057,N_15304);
nand U18463 (N_18463,N_15468,N_14427);
and U18464 (N_18464,N_14606,N_13043);
nand U18465 (N_18465,N_15727,N_14776);
nor U18466 (N_18466,N_12851,N_12568);
or U18467 (N_18467,N_15662,N_12310);
nand U18468 (N_18468,N_14306,N_12908);
or U18469 (N_18469,N_14578,N_12701);
and U18470 (N_18470,N_14182,N_15826);
nand U18471 (N_18471,N_15379,N_14788);
nor U18472 (N_18472,N_12935,N_13727);
or U18473 (N_18473,N_12834,N_12304);
xnor U18474 (N_18474,N_14235,N_12966);
nor U18475 (N_18475,N_15257,N_13211);
nand U18476 (N_18476,N_13945,N_14673);
or U18477 (N_18477,N_12650,N_15938);
or U18478 (N_18478,N_13940,N_12393);
nand U18479 (N_18479,N_12718,N_14742);
nand U18480 (N_18480,N_15928,N_12779);
nor U18481 (N_18481,N_14891,N_12085);
nor U18482 (N_18482,N_13771,N_15810);
and U18483 (N_18483,N_14424,N_15846);
nor U18484 (N_18484,N_13536,N_13829);
and U18485 (N_18485,N_14983,N_15103);
nand U18486 (N_18486,N_13679,N_15907);
nor U18487 (N_18487,N_13112,N_15789);
and U18488 (N_18488,N_15670,N_15462);
nor U18489 (N_18489,N_15180,N_14532);
or U18490 (N_18490,N_14371,N_12555);
nor U18491 (N_18491,N_12141,N_15107);
and U18492 (N_18492,N_15612,N_12346);
or U18493 (N_18493,N_15657,N_15304);
or U18494 (N_18494,N_15523,N_14295);
and U18495 (N_18495,N_15191,N_13145);
and U18496 (N_18496,N_14402,N_14944);
nand U18497 (N_18497,N_12338,N_12628);
and U18498 (N_18498,N_13474,N_14522);
or U18499 (N_18499,N_15937,N_15092);
or U18500 (N_18500,N_13693,N_13326);
nor U18501 (N_18501,N_13698,N_12771);
or U18502 (N_18502,N_12237,N_14708);
or U18503 (N_18503,N_15188,N_12924);
and U18504 (N_18504,N_15081,N_12597);
and U18505 (N_18505,N_12051,N_13017);
and U18506 (N_18506,N_13725,N_15347);
nand U18507 (N_18507,N_15415,N_13200);
nand U18508 (N_18508,N_14698,N_14916);
and U18509 (N_18509,N_12062,N_14341);
and U18510 (N_18510,N_12487,N_12467);
or U18511 (N_18511,N_12526,N_14435);
nand U18512 (N_18512,N_13272,N_12028);
or U18513 (N_18513,N_13496,N_14205);
or U18514 (N_18514,N_13105,N_13919);
nand U18515 (N_18515,N_14822,N_12020);
and U18516 (N_18516,N_14187,N_13761);
nand U18517 (N_18517,N_13715,N_14216);
and U18518 (N_18518,N_14957,N_13711);
nor U18519 (N_18519,N_15908,N_12368);
and U18520 (N_18520,N_14159,N_12035);
or U18521 (N_18521,N_12412,N_12813);
nand U18522 (N_18522,N_15420,N_13635);
nor U18523 (N_18523,N_13685,N_13559);
or U18524 (N_18524,N_12206,N_15091);
xnor U18525 (N_18525,N_14212,N_14764);
and U18526 (N_18526,N_15512,N_14118);
or U18527 (N_18527,N_13074,N_12279);
nor U18528 (N_18528,N_13541,N_13738);
nand U18529 (N_18529,N_12189,N_13621);
nor U18530 (N_18530,N_14023,N_13727);
or U18531 (N_18531,N_15993,N_12859);
or U18532 (N_18532,N_13632,N_14026);
and U18533 (N_18533,N_14982,N_14401);
nor U18534 (N_18534,N_15588,N_15570);
nor U18535 (N_18535,N_13128,N_14477);
or U18536 (N_18536,N_14206,N_13708);
nor U18537 (N_18537,N_13724,N_12593);
and U18538 (N_18538,N_13895,N_14048);
or U18539 (N_18539,N_15896,N_14114);
and U18540 (N_18540,N_14057,N_14181);
and U18541 (N_18541,N_13299,N_12158);
or U18542 (N_18542,N_13106,N_14716);
nand U18543 (N_18543,N_14513,N_14236);
nor U18544 (N_18544,N_12011,N_13656);
nor U18545 (N_18545,N_12369,N_13695);
nor U18546 (N_18546,N_12671,N_15057);
and U18547 (N_18547,N_12261,N_12513);
nand U18548 (N_18548,N_15778,N_13177);
or U18549 (N_18549,N_12223,N_15168);
or U18550 (N_18550,N_15788,N_15400);
nand U18551 (N_18551,N_13675,N_13477);
and U18552 (N_18552,N_12428,N_12917);
nand U18553 (N_18553,N_15460,N_14495);
nand U18554 (N_18554,N_13807,N_12869);
or U18555 (N_18555,N_12357,N_15570);
or U18556 (N_18556,N_13924,N_12276);
nand U18557 (N_18557,N_14040,N_13503);
nand U18558 (N_18558,N_14010,N_13506);
and U18559 (N_18559,N_13144,N_15826);
and U18560 (N_18560,N_13120,N_12260);
nor U18561 (N_18561,N_15121,N_14445);
nor U18562 (N_18562,N_15091,N_12783);
or U18563 (N_18563,N_13499,N_14700);
nand U18564 (N_18564,N_14052,N_15431);
and U18565 (N_18565,N_12970,N_13259);
nor U18566 (N_18566,N_14490,N_14872);
nor U18567 (N_18567,N_15507,N_12179);
and U18568 (N_18568,N_13489,N_12311);
and U18569 (N_18569,N_13421,N_15918);
nor U18570 (N_18570,N_12595,N_14717);
or U18571 (N_18571,N_13101,N_13525);
nor U18572 (N_18572,N_14276,N_15179);
and U18573 (N_18573,N_12031,N_15503);
and U18574 (N_18574,N_14441,N_12930);
or U18575 (N_18575,N_13953,N_12175);
or U18576 (N_18576,N_12156,N_15018);
or U18577 (N_18577,N_13564,N_14850);
nor U18578 (N_18578,N_12450,N_12355);
nand U18579 (N_18579,N_15094,N_12871);
nand U18580 (N_18580,N_14462,N_12497);
or U18581 (N_18581,N_13003,N_13149);
nand U18582 (N_18582,N_15872,N_13428);
or U18583 (N_18583,N_13723,N_12025);
nand U18584 (N_18584,N_14338,N_15742);
nand U18585 (N_18585,N_14301,N_14684);
nand U18586 (N_18586,N_13199,N_12908);
nand U18587 (N_18587,N_15094,N_13453);
or U18588 (N_18588,N_12267,N_15758);
nand U18589 (N_18589,N_12542,N_14025);
nand U18590 (N_18590,N_15254,N_15963);
or U18591 (N_18591,N_12012,N_13132);
nor U18592 (N_18592,N_13876,N_14157);
and U18593 (N_18593,N_15684,N_13097);
nand U18594 (N_18594,N_15674,N_15934);
or U18595 (N_18595,N_14103,N_15599);
or U18596 (N_18596,N_12836,N_13599);
nor U18597 (N_18597,N_12147,N_12283);
nor U18598 (N_18598,N_14175,N_15853);
nor U18599 (N_18599,N_12367,N_12983);
or U18600 (N_18600,N_12857,N_13539);
and U18601 (N_18601,N_12019,N_13484);
nor U18602 (N_18602,N_12181,N_13324);
and U18603 (N_18603,N_13157,N_14918);
or U18604 (N_18604,N_12560,N_14132);
and U18605 (N_18605,N_15748,N_15043);
nor U18606 (N_18606,N_12671,N_14469);
nor U18607 (N_18607,N_15079,N_14245);
or U18608 (N_18608,N_15891,N_13909);
xor U18609 (N_18609,N_14872,N_15392);
and U18610 (N_18610,N_12193,N_15442);
or U18611 (N_18611,N_15523,N_13626);
and U18612 (N_18612,N_12274,N_14582);
nand U18613 (N_18613,N_12496,N_14560);
nand U18614 (N_18614,N_13166,N_14414);
nor U18615 (N_18615,N_14813,N_15590);
or U18616 (N_18616,N_14698,N_12818);
nor U18617 (N_18617,N_14194,N_15623);
or U18618 (N_18618,N_12287,N_14949);
or U18619 (N_18619,N_14439,N_12683);
nand U18620 (N_18620,N_12551,N_14371);
nand U18621 (N_18621,N_15819,N_15839);
or U18622 (N_18622,N_15642,N_15457);
or U18623 (N_18623,N_14374,N_13958);
and U18624 (N_18624,N_12056,N_12653);
nor U18625 (N_18625,N_12016,N_15613);
nor U18626 (N_18626,N_13457,N_14929);
and U18627 (N_18627,N_14211,N_14328);
nor U18628 (N_18628,N_12046,N_14582);
nor U18629 (N_18629,N_12541,N_14712);
and U18630 (N_18630,N_14419,N_12208);
and U18631 (N_18631,N_14530,N_12627);
or U18632 (N_18632,N_14717,N_14090);
nand U18633 (N_18633,N_12964,N_15674);
nand U18634 (N_18634,N_15157,N_14361);
and U18635 (N_18635,N_15025,N_15911);
nand U18636 (N_18636,N_12316,N_13275);
or U18637 (N_18637,N_13321,N_12527);
and U18638 (N_18638,N_15956,N_14061);
and U18639 (N_18639,N_12972,N_13480);
nor U18640 (N_18640,N_12403,N_12604);
nand U18641 (N_18641,N_14936,N_15169);
or U18642 (N_18642,N_15927,N_15644);
and U18643 (N_18643,N_15550,N_13112);
nor U18644 (N_18644,N_15932,N_14791);
or U18645 (N_18645,N_12040,N_15604);
or U18646 (N_18646,N_15052,N_13952);
nor U18647 (N_18647,N_15541,N_13113);
nor U18648 (N_18648,N_14850,N_15348);
nor U18649 (N_18649,N_15486,N_14066);
and U18650 (N_18650,N_13437,N_15314);
or U18651 (N_18651,N_14165,N_12062);
nor U18652 (N_18652,N_15342,N_14355);
nand U18653 (N_18653,N_15713,N_12346);
or U18654 (N_18654,N_13850,N_13564);
or U18655 (N_18655,N_12458,N_13461);
or U18656 (N_18656,N_13859,N_15153);
and U18657 (N_18657,N_14793,N_14918);
nand U18658 (N_18658,N_12210,N_14041);
nor U18659 (N_18659,N_15937,N_15044);
and U18660 (N_18660,N_12736,N_12552);
and U18661 (N_18661,N_13447,N_14786);
nand U18662 (N_18662,N_15677,N_12452);
xor U18663 (N_18663,N_13871,N_15077);
and U18664 (N_18664,N_13265,N_15323);
nand U18665 (N_18665,N_12328,N_14210);
nor U18666 (N_18666,N_13184,N_15847);
nand U18667 (N_18667,N_14036,N_13997);
nor U18668 (N_18668,N_13135,N_13103);
and U18669 (N_18669,N_12912,N_15948);
or U18670 (N_18670,N_14733,N_15823);
nand U18671 (N_18671,N_15704,N_15342);
or U18672 (N_18672,N_13700,N_14023);
and U18673 (N_18673,N_13198,N_15120);
xnor U18674 (N_18674,N_13456,N_13076);
or U18675 (N_18675,N_13115,N_13480);
and U18676 (N_18676,N_14555,N_15730);
or U18677 (N_18677,N_14346,N_14984);
nor U18678 (N_18678,N_15189,N_13782);
nand U18679 (N_18679,N_14431,N_15621);
nor U18680 (N_18680,N_15464,N_14973);
and U18681 (N_18681,N_12643,N_13976);
and U18682 (N_18682,N_13115,N_14218);
and U18683 (N_18683,N_13084,N_12800);
or U18684 (N_18684,N_13042,N_15744);
or U18685 (N_18685,N_14877,N_14554);
or U18686 (N_18686,N_12087,N_12118);
and U18687 (N_18687,N_15284,N_13589);
and U18688 (N_18688,N_15752,N_15446);
nand U18689 (N_18689,N_15320,N_14741);
nand U18690 (N_18690,N_12704,N_15450);
or U18691 (N_18691,N_12767,N_14951);
nor U18692 (N_18692,N_12373,N_13847);
xnor U18693 (N_18693,N_14346,N_15018);
nand U18694 (N_18694,N_15848,N_13673);
or U18695 (N_18695,N_14265,N_13773);
nand U18696 (N_18696,N_14219,N_14467);
nand U18697 (N_18697,N_13999,N_13630);
and U18698 (N_18698,N_15710,N_15796);
and U18699 (N_18699,N_14576,N_14498);
nor U18700 (N_18700,N_13528,N_13889);
or U18701 (N_18701,N_15677,N_14745);
and U18702 (N_18702,N_15866,N_12801);
nand U18703 (N_18703,N_12369,N_12074);
nand U18704 (N_18704,N_13325,N_12303);
nor U18705 (N_18705,N_12761,N_12061);
nor U18706 (N_18706,N_14744,N_12638);
or U18707 (N_18707,N_14655,N_14739);
or U18708 (N_18708,N_13740,N_13630);
or U18709 (N_18709,N_12847,N_15499);
and U18710 (N_18710,N_13763,N_12701);
nand U18711 (N_18711,N_15695,N_15434);
and U18712 (N_18712,N_14538,N_14595);
and U18713 (N_18713,N_14956,N_12574);
nor U18714 (N_18714,N_14215,N_15381);
or U18715 (N_18715,N_14568,N_13409);
and U18716 (N_18716,N_15428,N_15997);
and U18717 (N_18717,N_15138,N_14331);
nor U18718 (N_18718,N_12222,N_14861);
or U18719 (N_18719,N_15517,N_13316);
nand U18720 (N_18720,N_15027,N_15272);
and U18721 (N_18721,N_14182,N_13968);
and U18722 (N_18722,N_13645,N_12494);
and U18723 (N_18723,N_15639,N_12275);
nand U18724 (N_18724,N_15372,N_14815);
and U18725 (N_18725,N_13101,N_14081);
nand U18726 (N_18726,N_13129,N_12230);
nand U18727 (N_18727,N_14378,N_14726);
nand U18728 (N_18728,N_12591,N_13474);
nor U18729 (N_18729,N_13959,N_14331);
or U18730 (N_18730,N_13283,N_13865);
and U18731 (N_18731,N_14812,N_14520);
nand U18732 (N_18732,N_12410,N_12538);
and U18733 (N_18733,N_12613,N_13616);
nand U18734 (N_18734,N_14382,N_12063);
nand U18735 (N_18735,N_15933,N_12332);
and U18736 (N_18736,N_14620,N_15899);
nand U18737 (N_18737,N_13722,N_13444);
or U18738 (N_18738,N_14668,N_12672);
or U18739 (N_18739,N_15689,N_15900);
or U18740 (N_18740,N_15468,N_14839);
nor U18741 (N_18741,N_12107,N_15647);
or U18742 (N_18742,N_13710,N_12652);
nand U18743 (N_18743,N_15840,N_14279);
or U18744 (N_18744,N_15127,N_12668);
and U18745 (N_18745,N_15919,N_12715);
nand U18746 (N_18746,N_12924,N_13128);
nor U18747 (N_18747,N_13126,N_14526);
nor U18748 (N_18748,N_12876,N_15290);
and U18749 (N_18749,N_14218,N_13255);
nand U18750 (N_18750,N_15358,N_12313);
or U18751 (N_18751,N_12280,N_15036);
nor U18752 (N_18752,N_12043,N_15345);
and U18753 (N_18753,N_13735,N_15064);
or U18754 (N_18754,N_15389,N_13714);
nor U18755 (N_18755,N_13204,N_14970);
and U18756 (N_18756,N_13304,N_15810);
nand U18757 (N_18757,N_12519,N_14718);
or U18758 (N_18758,N_14221,N_13332);
nor U18759 (N_18759,N_13405,N_15432);
xor U18760 (N_18760,N_15275,N_12302);
and U18761 (N_18761,N_13630,N_14503);
nand U18762 (N_18762,N_12445,N_13303);
xnor U18763 (N_18763,N_13026,N_14085);
nand U18764 (N_18764,N_15174,N_14864);
nor U18765 (N_18765,N_12230,N_14481);
and U18766 (N_18766,N_13895,N_13470);
nand U18767 (N_18767,N_13912,N_15957);
nor U18768 (N_18768,N_12375,N_14087);
nor U18769 (N_18769,N_12107,N_12775);
nor U18770 (N_18770,N_14704,N_15833);
nand U18771 (N_18771,N_14240,N_14845);
nor U18772 (N_18772,N_15321,N_15837);
nand U18773 (N_18773,N_15498,N_12661);
xor U18774 (N_18774,N_12244,N_14292);
or U18775 (N_18775,N_13251,N_14926);
and U18776 (N_18776,N_15578,N_12408);
nor U18777 (N_18777,N_15228,N_15659);
nor U18778 (N_18778,N_15538,N_15178);
and U18779 (N_18779,N_12878,N_12197);
or U18780 (N_18780,N_12189,N_15779);
or U18781 (N_18781,N_12569,N_15203);
and U18782 (N_18782,N_15001,N_12930);
and U18783 (N_18783,N_13678,N_13785);
or U18784 (N_18784,N_14965,N_14893);
nor U18785 (N_18785,N_12632,N_13314);
or U18786 (N_18786,N_15648,N_15162);
nand U18787 (N_18787,N_12127,N_13994);
nand U18788 (N_18788,N_12996,N_12665);
nand U18789 (N_18789,N_13535,N_15459);
or U18790 (N_18790,N_12281,N_12178);
nand U18791 (N_18791,N_12388,N_13338);
nand U18792 (N_18792,N_12971,N_15114);
and U18793 (N_18793,N_14104,N_12426);
or U18794 (N_18794,N_15975,N_12910);
or U18795 (N_18795,N_14963,N_12751);
nor U18796 (N_18796,N_15995,N_12470);
or U18797 (N_18797,N_12067,N_13157);
nor U18798 (N_18798,N_15148,N_15431);
nor U18799 (N_18799,N_13356,N_12467);
or U18800 (N_18800,N_15763,N_14314);
nor U18801 (N_18801,N_12777,N_13607);
or U18802 (N_18802,N_12808,N_12812);
or U18803 (N_18803,N_12356,N_14408);
nor U18804 (N_18804,N_13245,N_15209);
xor U18805 (N_18805,N_14313,N_13006);
and U18806 (N_18806,N_13947,N_14065);
and U18807 (N_18807,N_15827,N_14611);
nor U18808 (N_18808,N_13836,N_12858);
and U18809 (N_18809,N_13804,N_12982);
nor U18810 (N_18810,N_14064,N_12635);
nor U18811 (N_18811,N_13708,N_15440);
nor U18812 (N_18812,N_12489,N_13154);
nor U18813 (N_18813,N_13235,N_13629);
or U18814 (N_18814,N_15336,N_13156);
or U18815 (N_18815,N_12079,N_12158);
nor U18816 (N_18816,N_13883,N_14326);
nand U18817 (N_18817,N_12433,N_14369);
nand U18818 (N_18818,N_13371,N_13463);
nand U18819 (N_18819,N_14184,N_14746);
or U18820 (N_18820,N_12980,N_12455);
nor U18821 (N_18821,N_15398,N_13575);
nor U18822 (N_18822,N_14776,N_15882);
nor U18823 (N_18823,N_15478,N_14570);
nor U18824 (N_18824,N_13267,N_14084);
nand U18825 (N_18825,N_15295,N_14174);
nand U18826 (N_18826,N_13229,N_14896);
nor U18827 (N_18827,N_13393,N_14360);
and U18828 (N_18828,N_12537,N_12018);
nand U18829 (N_18829,N_13141,N_12849);
xnor U18830 (N_18830,N_12788,N_14286);
and U18831 (N_18831,N_12137,N_14269);
or U18832 (N_18832,N_14423,N_12861);
nand U18833 (N_18833,N_15437,N_14366);
and U18834 (N_18834,N_14532,N_12304);
nor U18835 (N_18835,N_12041,N_12285);
nor U18836 (N_18836,N_14222,N_15832);
and U18837 (N_18837,N_14302,N_14775);
nand U18838 (N_18838,N_14768,N_12588);
and U18839 (N_18839,N_13122,N_12981);
or U18840 (N_18840,N_13642,N_13588);
nand U18841 (N_18841,N_13288,N_12974);
nand U18842 (N_18842,N_15435,N_14737);
and U18843 (N_18843,N_13968,N_13884);
nand U18844 (N_18844,N_15755,N_13007);
nand U18845 (N_18845,N_14325,N_13067);
and U18846 (N_18846,N_14830,N_12177);
nor U18847 (N_18847,N_12496,N_12262);
nand U18848 (N_18848,N_12179,N_13591);
nand U18849 (N_18849,N_14477,N_14525);
nand U18850 (N_18850,N_12587,N_12420);
or U18851 (N_18851,N_12681,N_15073);
and U18852 (N_18852,N_13992,N_13898);
nor U18853 (N_18853,N_14351,N_14807);
or U18854 (N_18854,N_15497,N_13258);
and U18855 (N_18855,N_13115,N_13642);
nand U18856 (N_18856,N_12007,N_12237);
or U18857 (N_18857,N_15617,N_13220);
or U18858 (N_18858,N_13637,N_14171);
nand U18859 (N_18859,N_13398,N_12724);
xor U18860 (N_18860,N_15425,N_15008);
nor U18861 (N_18861,N_15247,N_12676);
nand U18862 (N_18862,N_12792,N_12657);
nand U18863 (N_18863,N_13391,N_14422);
or U18864 (N_18864,N_14548,N_14098);
or U18865 (N_18865,N_13315,N_15441);
and U18866 (N_18866,N_13919,N_14638);
nand U18867 (N_18867,N_14055,N_12474);
nand U18868 (N_18868,N_14224,N_15271);
nand U18869 (N_18869,N_12364,N_14613);
or U18870 (N_18870,N_12035,N_14118);
nand U18871 (N_18871,N_15319,N_12386);
or U18872 (N_18872,N_15045,N_14135);
and U18873 (N_18873,N_13182,N_15463);
and U18874 (N_18874,N_13876,N_15514);
nor U18875 (N_18875,N_12802,N_14174);
or U18876 (N_18876,N_14219,N_14961);
nor U18877 (N_18877,N_13922,N_13037);
or U18878 (N_18878,N_13536,N_13631);
nor U18879 (N_18879,N_13881,N_15106);
nor U18880 (N_18880,N_13426,N_12721);
nand U18881 (N_18881,N_12993,N_15766);
or U18882 (N_18882,N_14823,N_12262);
or U18883 (N_18883,N_12729,N_13232);
and U18884 (N_18884,N_12005,N_12911);
or U18885 (N_18885,N_12602,N_15589);
nand U18886 (N_18886,N_14171,N_14686);
and U18887 (N_18887,N_15531,N_14631);
nand U18888 (N_18888,N_13681,N_12338);
or U18889 (N_18889,N_15456,N_13949);
or U18890 (N_18890,N_14759,N_14218);
nand U18891 (N_18891,N_13614,N_13127);
or U18892 (N_18892,N_12566,N_14549);
and U18893 (N_18893,N_12850,N_15603);
nand U18894 (N_18894,N_15812,N_13301);
nor U18895 (N_18895,N_15183,N_12367);
nor U18896 (N_18896,N_15279,N_14666);
or U18897 (N_18897,N_15647,N_14970);
or U18898 (N_18898,N_15908,N_13998);
nor U18899 (N_18899,N_15417,N_13438);
or U18900 (N_18900,N_15704,N_15021);
nand U18901 (N_18901,N_13307,N_12083);
nor U18902 (N_18902,N_12360,N_14605);
nand U18903 (N_18903,N_14188,N_14835);
nor U18904 (N_18904,N_12386,N_13983);
and U18905 (N_18905,N_15546,N_13248);
and U18906 (N_18906,N_12464,N_12423);
or U18907 (N_18907,N_14260,N_15969);
nand U18908 (N_18908,N_13285,N_15211);
and U18909 (N_18909,N_15133,N_12495);
nor U18910 (N_18910,N_13093,N_13278);
or U18911 (N_18911,N_12490,N_15099);
nand U18912 (N_18912,N_15917,N_15429);
nand U18913 (N_18913,N_15600,N_13299);
or U18914 (N_18914,N_14415,N_15464);
nand U18915 (N_18915,N_12650,N_14493);
nand U18916 (N_18916,N_13007,N_14575);
nor U18917 (N_18917,N_12335,N_14953);
or U18918 (N_18918,N_12715,N_15280);
or U18919 (N_18919,N_15081,N_15029);
nand U18920 (N_18920,N_15312,N_12558);
nor U18921 (N_18921,N_14479,N_13471);
and U18922 (N_18922,N_13093,N_14684);
or U18923 (N_18923,N_15283,N_15385);
or U18924 (N_18924,N_14216,N_12830);
nor U18925 (N_18925,N_14736,N_12168);
or U18926 (N_18926,N_15184,N_13211);
nand U18927 (N_18927,N_14567,N_15032);
or U18928 (N_18928,N_13523,N_12403);
or U18929 (N_18929,N_14275,N_13592);
nor U18930 (N_18930,N_12335,N_13100);
nor U18931 (N_18931,N_14071,N_12785);
nor U18932 (N_18932,N_12230,N_12749);
or U18933 (N_18933,N_12630,N_15687);
nor U18934 (N_18934,N_14114,N_14347);
and U18935 (N_18935,N_13539,N_15597);
nor U18936 (N_18936,N_14475,N_15774);
or U18937 (N_18937,N_13449,N_13790);
and U18938 (N_18938,N_15488,N_12428);
or U18939 (N_18939,N_13395,N_12198);
or U18940 (N_18940,N_12303,N_12625);
and U18941 (N_18941,N_14362,N_12636);
or U18942 (N_18942,N_14925,N_15630);
or U18943 (N_18943,N_13222,N_15725);
or U18944 (N_18944,N_12538,N_12967);
nor U18945 (N_18945,N_14482,N_14735);
and U18946 (N_18946,N_12302,N_12775);
nor U18947 (N_18947,N_12711,N_12624);
or U18948 (N_18948,N_14134,N_12237);
nand U18949 (N_18949,N_12130,N_13096);
nor U18950 (N_18950,N_15741,N_14350);
or U18951 (N_18951,N_13704,N_15085);
and U18952 (N_18952,N_15098,N_13357);
and U18953 (N_18953,N_14432,N_15589);
nand U18954 (N_18954,N_13093,N_13770);
and U18955 (N_18955,N_14637,N_13446);
and U18956 (N_18956,N_15402,N_13510);
nor U18957 (N_18957,N_12544,N_15201);
or U18958 (N_18958,N_13231,N_14285);
or U18959 (N_18959,N_13035,N_15019);
nor U18960 (N_18960,N_12595,N_15526);
or U18961 (N_18961,N_15859,N_15119);
nand U18962 (N_18962,N_12918,N_14095);
nor U18963 (N_18963,N_13732,N_15904);
nand U18964 (N_18964,N_15356,N_14320);
or U18965 (N_18965,N_13616,N_13176);
nand U18966 (N_18966,N_13676,N_15275);
and U18967 (N_18967,N_12237,N_14717);
nor U18968 (N_18968,N_15086,N_13040);
nand U18969 (N_18969,N_12723,N_12369);
nor U18970 (N_18970,N_12550,N_14223);
nand U18971 (N_18971,N_13006,N_12105);
nand U18972 (N_18972,N_13061,N_15607);
nor U18973 (N_18973,N_15002,N_15804);
nor U18974 (N_18974,N_12867,N_14991);
nand U18975 (N_18975,N_12703,N_14361);
and U18976 (N_18976,N_14168,N_13957);
and U18977 (N_18977,N_13742,N_15609);
nor U18978 (N_18978,N_13134,N_13298);
and U18979 (N_18979,N_12633,N_14076);
nor U18980 (N_18980,N_12128,N_15870);
and U18981 (N_18981,N_13317,N_15867);
nor U18982 (N_18982,N_15120,N_15097);
nor U18983 (N_18983,N_14219,N_13071);
or U18984 (N_18984,N_14203,N_12213);
and U18985 (N_18985,N_13302,N_12903);
and U18986 (N_18986,N_14602,N_15536);
nand U18987 (N_18987,N_13398,N_15251);
and U18988 (N_18988,N_13868,N_13270);
and U18989 (N_18989,N_15537,N_14670);
nand U18990 (N_18990,N_12103,N_14717);
xor U18991 (N_18991,N_12341,N_12532);
nor U18992 (N_18992,N_12029,N_15411);
nor U18993 (N_18993,N_15861,N_14427);
and U18994 (N_18994,N_13451,N_13004);
nand U18995 (N_18995,N_15918,N_12608);
or U18996 (N_18996,N_12317,N_13858);
and U18997 (N_18997,N_14174,N_14652);
nor U18998 (N_18998,N_15847,N_12261);
nor U18999 (N_18999,N_13232,N_13490);
and U19000 (N_19000,N_13731,N_13320);
or U19001 (N_19001,N_13344,N_15237);
and U19002 (N_19002,N_13340,N_14773);
nand U19003 (N_19003,N_15537,N_15515);
nand U19004 (N_19004,N_15083,N_13104);
nand U19005 (N_19005,N_13781,N_14128);
nand U19006 (N_19006,N_13658,N_12505);
nor U19007 (N_19007,N_14328,N_15167);
or U19008 (N_19008,N_14336,N_13592);
nand U19009 (N_19009,N_15307,N_15377);
and U19010 (N_19010,N_14859,N_13937);
nor U19011 (N_19011,N_15331,N_13963);
and U19012 (N_19012,N_12618,N_15118);
and U19013 (N_19013,N_15683,N_13839);
and U19014 (N_19014,N_12023,N_13639);
nand U19015 (N_19015,N_12100,N_13913);
or U19016 (N_19016,N_13129,N_13185);
and U19017 (N_19017,N_13442,N_12350);
nand U19018 (N_19018,N_12694,N_14849);
nor U19019 (N_19019,N_14094,N_15821);
nor U19020 (N_19020,N_13936,N_14063);
or U19021 (N_19021,N_12566,N_15632);
and U19022 (N_19022,N_13616,N_13056);
nand U19023 (N_19023,N_15413,N_15067);
nor U19024 (N_19024,N_15173,N_15510);
and U19025 (N_19025,N_15963,N_12605);
or U19026 (N_19026,N_14601,N_14621);
nand U19027 (N_19027,N_13557,N_15267);
or U19028 (N_19028,N_15127,N_14599);
nor U19029 (N_19029,N_12367,N_15777);
xnor U19030 (N_19030,N_13707,N_15046);
and U19031 (N_19031,N_12551,N_12304);
or U19032 (N_19032,N_12083,N_12526);
and U19033 (N_19033,N_15474,N_14159);
nor U19034 (N_19034,N_14672,N_14013);
and U19035 (N_19035,N_14136,N_13237);
or U19036 (N_19036,N_15015,N_15675);
and U19037 (N_19037,N_15956,N_15352);
nor U19038 (N_19038,N_12487,N_15543);
or U19039 (N_19039,N_12922,N_14441);
and U19040 (N_19040,N_14610,N_13220);
or U19041 (N_19041,N_12010,N_12343);
xor U19042 (N_19042,N_15361,N_15784);
nand U19043 (N_19043,N_14969,N_12117);
and U19044 (N_19044,N_15913,N_14062);
or U19045 (N_19045,N_13803,N_15720);
xor U19046 (N_19046,N_15470,N_12939);
and U19047 (N_19047,N_14767,N_12784);
or U19048 (N_19048,N_15787,N_15939);
or U19049 (N_19049,N_12699,N_15892);
nand U19050 (N_19050,N_14987,N_14736);
nand U19051 (N_19051,N_12572,N_15957);
nor U19052 (N_19052,N_12288,N_14397);
nor U19053 (N_19053,N_15944,N_12697);
and U19054 (N_19054,N_15039,N_14783);
or U19055 (N_19055,N_14933,N_15847);
or U19056 (N_19056,N_12701,N_12520);
nor U19057 (N_19057,N_12756,N_15380);
and U19058 (N_19058,N_13796,N_12632);
or U19059 (N_19059,N_13767,N_14829);
and U19060 (N_19060,N_14877,N_12433);
and U19061 (N_19061,N_12082,N_12073);
and U19062 (N_19062,N_12674,N_14390);
nand U19063 (N_19063,N_14791,N_12727);
nor U19064 (N_19064,N_12684,N_14101);
nand U19065 (N_19065,N_15197,N_13689);
or U19066 (N_19066,N_12626,N_15684);
and U19067 (N_19067,N_14684,N_13806);
or U19068 (N_19068,N_14122,N_15778);
or U19069 (N_19069,N_12226,N_13878);
nand U19070 (N_19070,N_13511,N_12918);
nand U19071 (N_19071,N_12310,N_15571);
and U19072 (N_19072,N_14161,N_12423);
nor U19073 (N_19073,N_13639,N_13969);
nor U19074 (N_19074,N_14777,N_15914);
nand U19075 (N_19075,N_15175,N_14448);
nor U19076 (N_19076,N_12176,N_15312);
and U19077 (N_19077,N_12348,N_13702);
or U19078 (N_19078,N_15437,N_14628);
nand U19079 (N_19079,N_15232,N_15913);
nand U19080 (N_19080,N_13177,N_13703);
nor U19081 (N_19081,N_13250,N_15594);
nand U19082 (N_19082,N_13556,N_14637);
nand U19083 (N_19083,N_15869,N_13095);
or U19084 (N_19084,N_13946,N_15248);
nor U19085 (N_19085,N_12080,N_14787);
or U19086 (N_19086,N_13201,N_12922);
nand U19087 (N_19087,N_14443,N_14751);
and U19088 (N_19088,N_14623,N_14399);
or U19089 (N_19089,N_14022,N_13334);
or U19090 (N_19090,N_14141,N_14921);
and U19091 (N_19091,N_15985,N_14498);
nand U19092 (N_19092,N_15983,N_12907);
nor U19093 (N_19093,N_13139,N_14144);
and U19094 (N_19094,N_12086,N_13564);
nor U19095 (N_19095,N_15846,N_12340);
nor U19096 (N_19096,N_14414,N_15919);
or U19097 (N_19097,N_13627,N_12105);
and U19098 (N_19098,N_14372,N_14035);
and U19099 (N_19099,N_12801,N_15051);
nor U19100 (N_19100,N_13763,N_15141);
or U19101 (N_19101,N_12539,N_12106);
or U19102 (N_19102,N_13768,N_14166);
or U19103 (N_19103,N_12361,N_12663);
nand U19104 (N_19104,N_12284,N_14068);
nand U19105 (N_19105,N_14812,N_14497);
nand U19106 (N_19106,N_14364,N_13801);
and U19107 (N_19107,N_13510,N_15743);
nand U19108 (N_19108,N_13134,N_13273);
nand U19109 (N_19109,N_12029,N_14980);
and U19110 (N_19110,N_15329,N_14649);
and U19111 (N_19111,N_13093,N_14827);
and U19112 (N_19112,N_15781,N_15806);
nor U19113 (N_19113,N_15593,N_12644);
or U19114 (N_19114,N_13690,N_12817);
nand U19115 (N_19115,N_12947,N_13990);
nor U19116 (N_19116,N_12451,N_13545);
or U19117 (N_19117,N_15932,N_14989);
and U19118 (N_19118,N_15457,N_12435);
nor U19119 (N_19119,N_15152,N_15736);
or U19120 (N_19120,N_15818,N_14044);
and U19121 (N_19121,N_15353,N_13940);
or U19122 (N_19122,N_12026,N_14543);
and U19123 (N_19123,N_12321,N_13721);
or U19124 (N_19124,N_15187,N_14178);
nand U19125 (N_19125,N_14770,N_14220);
xor U19126 (N_19126,N_12414,N_14537);
or U19127 (N_19127,N_14761,N_15241);
nor U19128 (N_19128,N_14951,N_12357);
nand U19129 (N_19129,N_13766,N_12692);
nand U19130 (N_19130,N_14422,N_12092);
nand U19131 (N_19131,N_15324,N_14511);
or U19132 (N_19132,N_13717,N_15102);
and U19133 (N_19133,N_12783,N_13402);
or U19134 (N_19134,N_15016,N_13607);
nand U19135 (N_19135,N_13659,N_15569);
or U19136 (N_19136,N_15933,N_15988);
and U19137 (N_19137,N_14432,N_14055);
nand U19138 (N_19138,N_15901,N_13281);
and U19139 (N_19139,N_12692,N_15957);
and U19140 (N_19140,N_15918,N_13268);
nand U19141 (N_19141,N_13963,N_15085);
nand U19142 (N_19142,N_15478,N_13706);
and U19143 (N_19143,N_15125,N_12040);
nor U19144 (N_19144,N_12406,N_15754);
and U19145 (N_19145,N_14379,N_13133);
nor U19146 (N_19146,N_12949,N_12332);
and U19147 (N_19147,N_14019,N_15044);
or U19148 (N_19148,N_12547,N_12309);
and U19149 (N_19149,N_15312,N_13086);
and U19150 (N_19150,N_15866,N_13243);
nand U19151 (N_19151,N_14928,N_14830);
and U19152 (N_19152,N_14178,N_15325);
nor U19153 (N_19153,N_12403,N_12066);
nor U19154 (N_19154,N_12784,N_12496);
nand U19155 (N_19155,N_15095,N_12876);
and U19156 (N_19156,N_14728,N_14157);
or U19157 (N_19157,N_14845,N_14495);
and U19158 (N_19158,N_15538,N_12354);
and U19159 (N_19159,N_14802,N_13260);
nor U19160 (N_19160,N_13344,N_13975);
nor U19161 (N_19161,N_13302,N_15509);
and U19162 (N_19162,N_15208,N_12940);
or U19163 (N_19163,N_12407,N_12483);
nor U19164 (N_19164,N_14779,N_14985);
or U19165 (N_19165,N_14453,N_15848);
or U19166 (N_19166,N_14219,N_14088);
and U19167 (N_19167,N_14330,N_12375);
nand U19168 (N_19168,N_15533,N_15226);
nor U19169 (N_19169,N_12526,N_15101);
or U19170 (N_19170,N_14444,N_12681);
nand U19171 (N_19171,N_13614,N_12111);
xnor U19172 (N_19172,N_15827,N_14281);
nor U19173 (N_19173,N_13215,N_14763);
xnor U19174 (N_19174,N_14856,N_15233);
nor U19175 (N_19175,N_15404,N_15298);
nor U19176 (N_19176,N_13249,N_13728);
nor U19177 (N_19177,N_13731,N_13125);
nor U19178 (N_19178,N_13810,N_13996);
and U19179 (N_19179,N_14537,N_15014);
nor U19180 (N_19180,N_13354,N_15619);
nor U19181 (N_19181,N_13232,N_14321);
nand U19182 (N_19182,N_14367,N_15402);
and U19183 (N_19183,N_15945,N_12286);
or U19184 (N_19184,N_12978,N_15940);
nand U19185 (N_19185,N_15371,N_14238);
nor U19186 (N_19186,N_12056,N_12937);
nor U19187 (N_19187,N_15728,N_15379);
or U19188 (N_19188,N_13007,N_15370);
nor U19189 (N_19189,N_14810,N_13406);
nor U19190 (N_19190,N_12930,N_12582);
nand U19191 (N_19191,N_12961,N_14035);
nand U19192 (N_19192,N_14684,N_13375);
nand U19193 (N_19193,N_12834,N_13190);
and U19194 (N_19194,N_13289,N_13573);
or U19195 (N_19195,N_15002,N_15016);
and U19196 (N_19196,N_12709,N_13039);
nand U19197 (N_19197,N_13199,N_14352);
and U19198 (N_19198,N_15487,N_14892);
nor U19199 (N_19199,N_12999,N_12203);
or U19200 (N_19200,N_15749,N_12899);
or U19201 (N_19201,N_13585,N_12874);
nor U19202 (N_19202,N_15354,N_14395);
nand U19203 (N_19203,N_14674,N_12320);
nor U19204 (N_19204,N_12644,N_14847);
nand U19205 (N_19205,N_13653,N_13533);
or U19206 (N_19206,N_15884,N_13953);
and U19207 (N_19207,N_12215,N_13352);
and U19208 (N_19208,N_12190,N_15628);
nor U19209 (N_19209,N_15693,N_12888);
nand U19210 (N_19210,N_12602,N_15405);
or U19211 (N_19211,N_13223,N_15224);
and U19212 (N_19212,N_13541,N_13617);
nand U19213 (N_19213,N_14699,N_15678);
or U19214 (N_19214,N_15545,N_13993);
xnor U19215 (N_19215,N_15934,N_14745);
xnor U19216 (N_19216,N_13113,N_13047);
nor U19217 (N_19217,N_14571,N_13349);
and U19218 (N_19218,N_12892,N_12973);
and U19219 (N_19219,N_14842,N_15715);
nor U19220 (N_19220,N_14608,N_14345);
nand U19221 (N_19221,N_13969,N_14210);
or U19222 (N_19222,N_15017,N_12484);
or U19223 (N_19223,N_13965,N_15080);
and U19224 (N_19224,N_13610,N_13207);
nor U19225 (N_19225,N_14193,N_12872);
nor U19226 (N_19226,N_13860,N_12464);
nor U19227 (N_19227,N_12015,N_13806);
and U19228 (N_19228,N_15964,N_15175);
nor U19229 (N_19229,N_14813,N_12251);
and U19230 (N_19230,N_13147,N_12608);
and U19231 (N_19231,N_12140,N_15391);
nor U19232 (N_19232,N_13698,N_15654);
nor U19233 (N_19233,N_13619,N_15290);
nand U19234 (N_19234,N_15413,N_15705);
and U19235 (N_19235,N_13356,N_14524);
and U19236 (N_19236,N_14289,N_14001);
nor U19237 (N_19237,N_15856,N_13534);
nand U19238 (N_19238,N_15152,N_15000);
and U19239 (N_19239,N_13321,N_12949);
and U19240 (N_19240,N_12596,N_14587);
nor U19241 (N_19241,N_14849,N_14735);
nand U19242 (N_19242,N_14053,N_15406);
or U19243 (N_19243,N_13411,N_15258);
and U19244 (N_19244,N_14445,N_13411);
or U19245 (N_19245,N_13888,N_12441);
nor U19246 (N_19246,N_14300,N_13549);
or U19247 (N_19247,N_14021,N_13640);
or U19248 (N_19248,N_12540,N_14065);
or U19249 (N_19249,N_14905,N_14506);
nor U19250 (N_19250,N_14016,N_15101);
or U19251 (N_19251,N_12842,N_12230);
and U19252 (N_19252,N_13483,N_15882);
and U19253 (N_19253,N_12504,N_15889);
nor U19254 (N_19254,N_14872,N_12907);
and U19255 (N_19255,N_14659,N_13788);
or U19256 (N_19256,N_15628,N_15164);
nor U19257 (N_19257,N_13199,N_12297);
or U19258 (N_19258,N_12879,N_13112);
or U19259 (N_19259,N_13534,N_12892);
nor U19260 (N_19260,N_14175,N_13927);
nor U19261 (N_19261,N_13316,N_12692);
or U19262 (N_19262,N_15513,N_12968);
nor U19263 (N_19263,N_12059,N_14379);
or U19264 (N_19264,N_13960,N_13929);
and U19265 (N_19265,N_15052,N_12074);
and U19266 (N_19266,N_14827,N_13962);
or U19267 (N_19267,N_13975,N_12964);
nor U19268 (N_19268,N_14978,N_13162);
nor U19269 (N_19269,N_12933,N_15284);
nor U19270 (N_19270,N_13659,N_14032);
and U19271 (N_19271,N_14199,N_12667);
and U19272 (N_19272,N_14929,N_14797);
nand U19273 (N_19273,N_15163,N_14093);
or U19274 (N_19274,N_14927,N_13164);
nand U19275 (N_19275,N_15176,N_15197);
and U19276 (N_19276,N_13739,N_14428);
or U19277 (N_19277,N_13059,N_12518);
or U19278 (N_19278,N_14563,N_13398);
or U19279 (N_19279,N_12764,N_12172);
nand U19280 (N_19280,N_15706,N_12576);
and U19281 (N_19281,N_13914,N_14031);
nand U19282 (N_19282,N_13780,N_14248);
nand U19283 (N_19283,N_12547,N_13187);
nor U19284 (N_19284,N_12701,N_14249);
or U19285 (N_19285,N_15919,N_13204);
nand U19286 (N_19286,N_13485,N_14574);
xnor U19287 (N_19287,N_13750,N_15061);
and U19288 (N_19288,N_14716,N_14658);
nand U19289 (N_19289,N_12347,N_12185);
and U19290 (N_19290,N_13761,N_13025);
nor U19291 (N_19291,N_12473,N_15602);
and U19292 (N_19292,N_15516,N_15919);
or U19293 (N_19293,N_14895,N_12405);
and U19294 (N_19294,N_13272,N_12710);
or U19295 (N_19295,N_13596,N_15701);
or U19296 (N_19296,N_13201,N_12453);
or U19297 (N_19297,N_15460,N_15729);
or U19298 (N_19298,N_15353,N_13125);
and U19299 (N_19299,N_13288,N_13089);
or U19300 (N_19300,N_12927,N_12459);
or U19301 (N_19301,N_15144,N_13603);
nor U19302 (N_19302,N_14392,N_12170);
and U19303 (N_19303,N_14014,N_13990);
nand U19304 (N_19304,N_13950,N_12996);
nand U19305 (N_19305,N_15974,N_13134);
nand U19306 (N_19306,N_12664,N_13472);
or U19307 (N_19307,N_14344,N_13903);
and U19308 (N_19308,N_14742,N_15996);
or U19309 (N_19309,N_14332,N_15592);
nand U19310 (N_19310,N_14212,N_12405);
nor U19311 (N_19311,N_12814,N_13293);
and U19312 (N_19312,N_14973,N_12546);
nand U19313 (N_19313,N_12179,N_12068);
and U19314 (N_19314,N_14505,N_13648);
and U19315 (N_19315,N_13677,N_14952);
nor U19316 (N_19316,N_13019,N_12809);
nor U19317 (N_19317,N_15474,N_12914);
nand U19318 (N_19318,N_15461,N_14114);
or U19319 (N_19319,N_15629,N_12275);
nand U19320 (N_19320,N_13426,N_12285);
or U19321 (N_19321,N_14795,N_13238);
nand U19322 (N_19322,N_13318,N_15224);
or U19323 (N_19323,N_14310,N_14487);
or U19324 (N_19324,N_14510,N_13180);
nor U19325 (N_19325,N_12423,N_13482);
nand U19326 (N_19326,N_14307,N_14777);
nor U19327 (N_19327,N_14784,N_15460);
nor U19328 (N_19328,N_14025,N_13579);
nand U19329 (N_19329,N_15830,N_14448);
nor U19330 (N_19330,N_15193,N_13984);
or U19331 (N_19331,N_14123,N_13406);
nand U19332 (N_19332,N_13494,N_14813);
nand U19333 (N_19333,N_12772,N_14573);
nand U19334 (N_19334,N_12605,N_15459);
nand U19335 (N_19335,N_15905,N_14352);
or U19336 (N_19336,N_14197,N_13547);
nor U19337 (N_19337,N_15369,N_13945);
or U19338 (N_19338,N_13212,N_13603);
nand U19339 (N_19339,N_12046,N_15978);
and U19340 (N_19340,N_14730,N_12296);
and U19341 (N_19341,N_14438,N_13647);
nand U19342 (N_19342,N_15693,N_12359);
nor U19343 (N_19343,N_13390,N_13029);
nor U19344 (N_19344,N_15616,N_12729);
and U19345 (N_19345,N_12903,N_12926);
nor U19346 (N_19346,N_13768,N_15350);
and U19347 (N_19347,N_15183,N_13947);
nand U19348 (N_19348,N_12394,N_12841);
nand U19349 (N_19349,N_13310,N_14248);
or U19350 (N_19350,N_13537,N_15049);
nor U19351 (N_19351,N_15939,N_12564);
nand U19352 (N_19352,N_14391,N_13190);
nand U19353 (N_19353,N_14813,N_13903);
and U19354 (N_19354,N_14159,N_12436);
and U19355 (N_19355,N_12601,N_15398);
or U19356 (N_19356,N_13068,N_12925);
or U19357 (N_19357,N_13664,N_12585);
or U19358 (N_19358,N_13095,N_14778);
nand U19359 (N_19359,N_12842,N_14312);
nor U19360 (N_19360,N_14815,N_15843);
nand U19361 (N_19361,N_15011,N_12407);
or U19362 (N_19362,N_12335,N_12010);
and U19363 (N_19363,N_13222,N_12264);
nor U19364 (N_19364,N_14001,N_14728);
nor U19365 (N_19365,N_13663,N_15246);
or U19366 (N_19366,N_12583,N_13612);
or U19367 (N_19367,N_12275,N_15876);
and U19368 (N_19368,N_12668,N_15914);
or U19369 (N_19369,N_14048,N_15737);
nor U19370 (N_19370,N_13543,N_13214);
nand U19371 (N_19371,N_15646,N_14213);
and U19372 (N_19372,N_12313,N_13185);
nand U19373 (N_19373,N_13993,N_14470);
nor U19374 (N_19374,N_13929,N_14378);
nand U19375 (N_19375,N_13756,N_14089);
nor U19376 (N_19376,N_14564,N_15439);
and U19377 (N_19377,N_12111,N_15101);
and U19378 (N_19378,N_13444,N_12500);
or U19379 (N_19379,N_12292,N_13362);
nand U19380 (N_19380,N_15274,N_12115);
or U19381 (N_19381,N_15484,N_13466);
or U19382 (N_19382,N_15098,N_13305);
nand U19383 (N_19383,N_15323,N_13295);
nand U19384 (N_19384,N_13773,N_13962);
or U19385 (N_19385,N_14786,N_14228);
nand U19386 (N_19386,N_15197,N_13911);
nor U19387 (N_19387,N_12180,N_15190);
nand U19388 (N_19388,N_12968,N_15566);
xor U19389 (N_19389,N_15551,N_14098);
nor U19390 (N_19390,N_14769,N_14840);
or U19391 (N_19391,N_15034,N_12023);
nor U19392 (N_19392,N_15983,N_13101);
or U19393 (N_19393,N_12598,N_13517);
nor U19394 (N_19394,N_13878,N_15497);
nor U19395 (N_19395,N_12923,N_12429);
nor U19396 (N_19396,N_13723,N_14157);
and U19397 (N_19397,N_12890,N_14401);
or U19398 (N_19398,N_15087,N_15785);
or U19399 (N_19399,N_15606,N_14627);
nand U19400 (N_19400,N_15747,N_15396);
nor U19401 (N_19401,N_14366,N_13524);
and U19402 (N_19402,N_13187,N_13732);
and U19403 (N_19403,N_15381,N_15489);
or U19404 (N_19404,N_15032,N_13389);
nor U19405 (N_19405,N_12918,N_14291);
nand U19406 (N_19406,N_14467,N_14146);
nand U19407 (N_19407,N_15795,N_12943);
and U19408 (N_19408,N_14021,N_12590);
nor U19409 (N_19409,N_15390,N_12484);
nand U19410 (N_19410,N_14918,N_15740);
and U19411 (N_19411,N_15943,N_13227);
or U19412 (N_19412,N_12601,N_12987);
and U19413 (N_19413,N_14416,N_15670);
nor U19414 (N_19414,N_15021,N_13066);
nor U19415 (N_19415,N_14502,N_15475);
and U19416 (N_19416,N_12477,N_13475);
and U19417 (N_19417,N_12325,N_13245);
nor U19418 (N_19418,N_12966,N_12109);
or U19419 (N_19419,N_14518,N_15860);
nor U19420 (N_19420,N_12270,N_12130);
nand U19421 (N_19421,N_13395,N_14841);
and U19422 (N_19422,N_15657,N_15663);
or U19423 (N_19423,N_14605,N_12211);
nand U19424 (N_19424,N_15231,N_13765);
nor U19425 (N_19425,N_15152,N_12727);
and U19426 (N_19426,N_15063,N_13672);
or U19427 (N_19427,N_12204,N_13469);
and U19428 (N_19428,N_12297,N_15803);
nor U19429 (N_19429,N_15527,N_12228);
nand U19430 (N_19430,N_14241,N_15757);
and U19431 (N_19431,N_12271,N_13504);
or U19432 (N_19432,N_15205,N_12587);
and U19433 (N_19433,N_14054,N_14280);
and U19434 (N_19434,N_15114,N_15137);
and U19435 (N_19435,N_12642,N_14868);
nor U19436 (N_19436,N_14803,N_14889);
and U19437 (N_19437,N_14056,N_13273);
or U19438 (N_19438,N_13751,N_15143);
nor U19439 (N_19439,N_15951,N_14128);
nor U19440 (N_19440,N_14616,N_13695);
nand U19441 (N_19441,N_15578,N_12057);
and U19442 (N_19442,N_15803,N_14626);
nor U19443 (N_19443,N_14930,N_14319);
nand U19444 (N_19444,N_13902,N_15038);
or U19445 (N_19445,N_14587,N_14107);
or U19446 (N_19446,N_13852,N_13523);
nor U19447 (N_19447,N_14587,N_12739);
and U19448 (N_19448,N_13212,N_12845);
or U19449 (N_19449,N_15566,N_12817);
or U19450 (N_19450,N_15265,N_12365);
nand U19451 (N_19451,N_15665,N_13185);
nand U19452 (N_19452,N_15389,N_13332);
nand U19453 (N_19453,N_12734,N_15749);
and U19454 (N_19454,N_12669,N_14556);
nor U19455 (N_19455,N_13453,N_13378);
and U19456 (N_19456,N_12613,N_12097);
or U19457 (N_19457,N_14456,N_15648);
nor U19458 (N_19458,N_15315,N_15554);
or U19459 (N_19459,N_15874,N_12800);
nor U19460 (N_19460,N_12076,N_13548);
nand U19461 (N_19461,N_12834,N_14107);
or U19462 (N_19462,N_14001,N_13476);
and U19463 (N_19463,N_15286,N_14999);
and U19464 (N_19464,N_14842,N_15221);
or U19465 (N_19465,N_15070,N_15641);
and U19466 (N_19466,N_12098,N_13018);
nand U19467 (N_19467,N_12207,N_14038);
nand U19468 (N_19468,N_13897,N_13279);
nor U19469 (N_19469,N_13101,N_15658);
and U19470 (N_19470,N_13855,N_15573);
or U19471 (N_19471,N_14404,N_15965);
or U19472 (N_19472,N_13946,N_15590);
and U19473 (N_19473,N_12347,N_13988);
nor U19474 (N_19474,N_13663,N_14587);
or U19475 (N_19475,N_15359,N_15271);
nand U19476 (N_19476,N_12076,N_15214);
and U19477 (N_19477,N_15862,N_13678);
or U19478 (N_19478,N_15059,N_13401);
and U19479 (N_19479,N_12661,N_12059);
and U19480 (N_19480,N_12201,N_15611);
or U19481 (N_19481,N_13966,N_13904);
and U19482 (N_19482,N_14062,N_12681);
nand U19483 (N_19483,N_15260,N_12085);
nor U19484 (N_19484,N_14170,N_14608);
nor U19485 (N_19485,N_15059,N_12241);
nor U19486 (N_19486,N_13451,N_12552);
and U19487 (N_19487,N_15935,N_14119);
nand U19488 (N_19488,N_15856,N_14879);
nand U19489 (N_19489,N_12202,N_13709);
and U19490 (N_19490,N_15595,N_14053);
nor U19491 (N_19491,N_12726,N_12316);
nor U19492 (N_19492,N_15469,N_15160);
nor U19493 (N_19493,N_15381,N_14298);
nor U19494 (N_19494,N_12294,N_13448);
and U19495 (N_19495,N_13279,N_14341);
nor U19496 (N_19496,N_12837,N_12995);
and U19497 (N_19497,N_13602,N_13707);
nor U19498 (N_19498,N_15996,N_12294);
or U19499 (N_19499,N_14951,N_15047);
or U19500 (N_19500,N_15200,N_12563);
nor U19501 (N_19501,N_14138,N_13815);
or U19502 (N_19502,N_13370,N_15307);
and U19503 (N_19503,N_14892,N_12428);
and U19504 (N_19504,N_13115,N_15869);
and U19505 (N_19505,N_13429,N_14762);
or U19506 (N_19506,N_15153,N_15326);
or U19507 (N_19507,N_13662,N_12950);
and U19508 (N_19508,N_15675,N_15710);
nand U19509 (N_19509,N_13560,N_12905);
nand U19510 (N_19510,N_14349,N_14571);
or U19511 (N_19511,N_13035,N_12132);
nand U19512 (N_19512,N_15257,N_15531);
nand U19513 (N_19513,N_13120,N_15987);
or U19514 (N_19514,N_13568,N_12297);
nand U19515 (N_19515,N_13876,N_15236);
nor U19516 (N_19516,N_15141,N_12533);
or U19517 (N_19517,N_12736,N_13259);
nand U19518 (N_19518,N_14855,N_12327);
nor U19519 (N_19519,N_15655,N_15959);
nand U19520 (N_19520,N_12520,N_14340);
nand U19521 (N_19521,N_15454,N_15304);
and U19522 (N_19522,N_14115,N_14308);
nor U19523 (N_19523,N_14986,N_14634);
nand U19524 (N_19524,N_12210,N_14653);
or U19525 (N_19525,N_14146,N_15079);
nor U19526 (N_19526,N_14578,N_12301);
xor U19527 (N_19527,N_15096,N_14203);
or U19528 (N_19528,N_15551,N_14120);
or U19529 (N_19529,N_15902,N_14584);
and U19530 (N_19530,N_14950,N_15739);
and U19531 (N_19531,N_14581,N_14447);
nor U19532 (N_19532,N_15938,N_13209);
and U19533 (N_19533,N_12095,N_13510);
nor U19534 (N_19534,N_14289,N_15478);
and U19535 (N_19535,N_14577,N_14532);
nand U19536 (N_19536,N_15436,N_12623);
and U19537 (N_19537,N_14326,N_13993);
nand U19538 (N_19538,N_15309,N_13564);
and U19539 (N_19539,N_13244,N_12941);
nand U19540 (N_19540,N_13800,N_12335);
nor U19541 (N_19541,N_14503,N_13745);
nor U19542 (N_19542,N_13594,N_15078);
and U19543 (N_19543,N_12940,N_15843);
nor U19544 (N_19544,N_14962,N_12627);
nand U19545 (N_19545,N_12163,N_13794);
or U19546 (N_19546,N_14049,N_12251);
nand U19547 (N_19547,N_12464,N_15418);
or U19548 (N_19548,N_15640,N_13996);
or U19549 (N_19549,N_14340,N_13925);
and U19550 (N_19550,N_14726,N_13644);
nand U19551 (N_19551,N_14297,N_12367);
nor U19552 (N_19552,N_14580,N_13225);
xor U19553 (N_19553,N_13937,N_14280);
and U19554 (N_19554,N_15304,N_15670);
and U19555 (N_19555,N_14663,N_12420);
and U19556 (N_19556,N_13316,N_15539);
and U19557 (N_19557,N_15158,N_13401);
or U19558 (N_19558,N_13305,N_13481);
nand U19559 (N_19559,N_14710,N_15744);
nor U19560 (N_19560,N_15805,N_15430);
nor U19561 (N_19561,N_13884,N_12699);
or U19562 (N_19562,N_12279,N_14545);
or U19563 (N_19563,N_15688,N_12942);
or U19564 (N_19564,N_12408,N_15887);
and U19565 (N_19565,N_15434,N_13012);
or U19566 (N_19566,N_12240,N_13109);
nand U19567 (N_19567,N_13812,N_12147);
nor U19568 (N_19568,N_14579,N_13126);
or U19569 (N_19569,N_12947,N_12995);
or U19570 (N_19570,N_15949,N_12009);
nand U19571 (N_19571,N_13789,N_13811);
and U19572 (N_19572,N_14025,N_12653);
and U19573 (N_19573,N_13037,N_13358);
and U19574 (N_19574,N_13741,N_13467);
or U19575 (N_19575,N_15351,N_12305);
and U19576 (N_19576,N_13493,N_15788);
nor U19577 (N_19577,N_13649,N_13530);
or U19578 (N_19578,N_12950,N_15990);
or U19579 (N_19579,N_12923,N_15701);
and U19580 (N_19580,N_14199,N_13891);
nor U19581 (N_19581,N_14390,N_14794);
or U19582 (N_19582,N_13534,N_13121);
nand U19583 (N_19583,N_13117,N_13077);
and U19584 (N_19584,N_15870,N_15731);
or U19585 (N_19585,N_12647,N_13748);
nor U19586 (N_19586,N_12016,N_15965);
nand U19587 (N_19587,N_14998,N_14032);
or U19588 (N_19588,N_14193,N_14181);
nand U19589 (N_19589,N_13317,N_15011);
nor U19590 (N_19590,N_15564,N_15287);
or U19591 (N_19591,N_14052,N_14988);
nand U19592 (N_19592,N_15827,N_13171);
nor U19593 (N_19593,N_15925,N_14030);
nand U19594 (N_19594,N_13257,N_13769);
nand U19595 (N_19595,N_14312,N_12296);
xnor U19596 (N_19596,N_14722,N_13152);
nand U19597 (N_19597,N_14412,N_13150);
nand U19598 (N_19598,N_12315,N_12839);
or U19599 (N_19599,N_15055,N_15960);
and U19600 (N_19600,N_12550,N_14195);
nor U19601 (N_19601,N_12325,N_15143);
nand U19602 (N_19602,N_15568,N_13650);
or U19603 (N_19603,N_14691,N_15796);
nor U19604 (N_19604,N_15323,N_15609);
nand U19605 (N_19605,N_12524,N_14469);
nor U19606 (N_19606,N_12698,N_13825);
nor U19607 (N_19607,N_12886,N_12473);
and U19608 (N_19608,N_14336,N_13291);
or U19609 (N_19609,N_15655,N_15104);
and U19610 (N_19610,N_14782,N_14427);
xnor U19611 (N_19611,N_14155,N_14468);
and U19612 (N_19612,N_15582,N_12414);
and U19613 (N_19613,N_14864,N_12047);
nor U19614 (N_19614,N_15667,N_14627);
or U19615 (N_19615,N_13743,N_14118);
and U19616 (N_19616,N_14917,N_15152);
or U19617 (N_19617,N_14371,N_13039);
xor U19618 (N_19618,N_13518,N_14214);
or U19619 (N_19619,N_12981,N_13718);
or U19620 (N_19620,N_12533,N_13080);
and U19621 (N_19621,N_12294,N_13070);
nand U19622 (N_19622,N_14247,N_12455);
nand U19623 (N_19623,N_14955,N_14714);
or U19624 (N_19624,N_12970,N_13425);
or U19625 (N_19625,N_13096,N_12795);
nor U19626 (N_19626,N_13127,N_14847);
nand U19627 (N_19627,N_14120,N_12047);
nor U19628 (N_19628,N_13819,N_12023);
and U19629 (N_19629,N_12043,N_12209);
and U19630 (N_19630,N_15750,N_13035);
nor U19631 (N_19631,N_13599,N_15449);
nor U19632 (N_19632,N_12172,N_14003);
and U19633 (N_19633,N_15658,N_12525);
and U19634 (N_19634,N_15792,N_12072);
and U19635 (N_19635,N_14538,N_12660);
or U19636 (N_19636,N_12572,N_14195);
and U19637 (N_19637,N_12727,N_15241);
and U19638 (N_19638,N_13591,N_15578);
or U19639 (N_19639,N_13254,N_14730);
nand U19640 (N_19640,N_13693,N_14181);
and U19641 (N_19641,N_15284,N_14693);
nor U19642 (N_19642,N_14884,N_12436);
nand U19643 (N_19643,N_14888,N_14347);
nand U19644 (N_19644,N_12015,N_15326);
or U19645 (N_19645,N_13999,N_12693);
and U19646 (N_19646,N_13538,N_13960);
nand U19647 (N_19647,N_14226,N_12982);
and U19648 (N_19648,N_14241,N_15567);
or U19649 (N_19649,N_13967,N_15304);
or U19650 (N_19650,N_12308,N_14155);
or U19651 (N_19651,N_12333,N_12830);
nand U19652 (N_19652,N_14637,N_14906);
and U19653 (N_19653,N_13611,N_13390);
nor U19654 (N_19654,N_15624,N_13453);
and U19655 (N_19655,N_14661,N_15573);
or U19656 (N_19656,N_14321,N_12820);
nor U19657 (N_19657,N_14737,N_14242);
nor U19658 (N_19658,N_15936,N_15960);
or U19659 (N_19659,N_15405,N_12344);
nand U19660 (N_19660,N_15066,N_12939);
or U19661 (N_19661,N_12292,N_14622);
nor U19662 (N_19662,N_13139,N_15505);
nand U19663 (N_19663,N_15461,N_15018);
xor U19664 (N_19664,N_12251,N_15348);
nand U19665 (N_19665,N_12404,N_12675);
nor U19666 (N_19666,N_15211,N_14336);
nand U19667 (N_19667,N_15575,N_15955);
or U19668 (N_19668,N_13626,N_12158);
nor U19669 (N_19669,N_15134,N_14502);
nand U19670 (N_19670,N_13924,N_13422);
or U19671 (N_19671,N_13460,N_14548);
nor U19672 (N_19672,N_15550,N_14750);
or U19673 (N_19673,N_13236,N_15059);
or U19674 (N_19674,N_15849,N_14047);
nand U19675 (N_19675,N_14009,N_12884);
and U19676 (N_19676,N_13095,N_14688);
and U19677 (N_19677,N_14813,N_15820);
and U19678 (N_19678,N_12995,N_13891);
and U19679 (N_19679,N_13287,N_13764);
nor U19680 (N_19680,N_12127,N_12545);
nand U19681 (N_19681,N_14111,N_12559);
nand U19682 (N_19682,N_12373,N_13720);
nand U19683 (N_19683,N_14116,N_14203);
and U19684 (N_19684,N_14276,N_14844);
or U19685 (N_19685,N_14628,N_13215);
nor U19686 (N_19686,N_12114,N_12073);
or U19687 (N_19687,N_14798,N_12246);
and U19688 (N_19688,N_12475,N_14616);
and U19689 (N_19689,N_14045,N_12386);
and U19690 (N_19690,N_13615,N_14021);
or U19691 (N_19691,N_14514,N_14919);
nand U19692 (N_19692,N_14452,N_14099);
and U19693 (N_19693,N_12922,N_13111);
nand U19694 (N_19694,N_12719,N_15044);
and U19695 (N_19695,N_12356,N_15093);
nand U19696 (N_19696,N_14440,N_14774);
nor U19697 (N_19697,N_12949,N_14518);
nor U19698 (N_19698,N_15318,N_12680);
or U19699 (N_19699,N_14005,N_15259);
and U19700 (N_19700,N_12345,N_13962);
and U19701 (N_19701,N_15030,N_12494);
nor U19702 (N_19702,N_13238,N_12732);
nor U19703 (N_19703,N_14814,N_14215);
and U19704 (N_19704,N_13950,N_14048);
nand U19705 (N_19705,N_12741,N_13429);
or U19706 (N_19706,N_14258,N_15589);
nand U19707 (N_19707,N_13818,N_13899);
or U19708 (N_19708,N_13698,N_13502);
or U19709 (N_19709,N_13030,N_14159);
nor U19710 (N_19710,N_15600,N_12126);
and U19711 (N_19711,N_14714,N_15602);
and U19712 (N_19712,N_12497,N_14110);
xor U19713 (N_19713,N_12093,N_13652);
nor U19714 (N_19714,N_12221,N_14711);
or U19715 (N_19715,N_14421,N_12150);
nand U19716 (N_19716,N_13993,N_15042);
nor U19717 (N_19717,N_14717,N_14171);
nor U19718 (N_19718,N_12384,N_13849);
nand U19719 (N_19719,N_12466,N_14816);
or U19720 (N_19720,N_13176,N_13960);
nor U19721 (N_19721,N_15505,N_15706);
nor U19722 (N_19722,N_15855,N_12707);
nor U19723 (N_19723,N_14664,N_12276);
nand U19724 (N_19724,N_13427,N_12221);
nand U19725 (N_19725,N_12222,N_12526);
or U19726 (N_19726,N_15410,N_13464);
nand U19727 (N_19727,N_13919,N_12640);
or U19728 (N_19728,N_12993,N_12620);
and U19729 (N_19729,N_14181,N_13133);
and U19730 (N_19730,N_14142,N_12695);
or U19731 (N_19731,N_13559,N_14504);
nor U19732 (N_19732,N_14250,N_15709);
and U19733 (N_19733,N_14066,N_15226);
nor U19734 (N_19734,N_13177,N_12347);
nor U19735 (N_19735,N_15938,N_13842);
nand U19736 (N_19736,N_13606,N_13941);
or U19737 (N_19737,N_14404,N_14092);
and U19738 (N_19738,N_13646,N_14876);
nor U19739 (N_19739,N_14464,N_14122);
or U19740 (N_19740,N_13432,N_13080);
nor U19741 (N_19741,N_13590,N_13689);
nor U19742 (N_19742,N_15736,N_12742);
nand U19743 (N_19743,N_13291,N_13617);
nand U19744 (N_19744,N_13718,N_12938);
or U19745 (N_19745,N_13748,N_13711);
or U19746 (N_19746,N_14912,N_14477);
nor U19747 (N_19747,N_14054,N_13090);
or U19748 (N_19748,N_15886,N_12289);
and U19749 (N_19749,N_13868,N_12334);
and U19750 (N_19750,N_12488,N_15116);
and U19751 (N_19751,N_15671,N_13660);
nor U19752 (N_19752,N_15763,N_15463);
nand U19753 (N_19753,N_14563,N_15915);
nand U19754 (N_19754,N_12462,N_15491);
nand U19755 (N_19755,N_12537,N_12725);
nor U19756 (N_19756,N_15502,N_15402);
and U19757 (N_19757,N_13671,N_15962);
or U19758 (N_19758,N_15114,N_15413);
and U19759 (N_19759,N_13641,N_14879);
and U19760 (N_19760,N_14569,N_13597);
and U19761 (N_19761,N_12968,N_13091);
and U19762 (N_19762,N_15458,N_13691);
nand U19763 (N_19763,N_14291,N_14469);
nor U19764 (N_19764,N_12986,N_12883);
and U19765 (N_19765,N_12820,N_13024);
and U19766 (N_19766,N_15590,N_12530);
nor U19767 (N_19767,N_14708,N_14974);
and U19768 (N_19768,N_13517,N_14587);
nand U19769 (N_19769,N_12031,N_12599);
and U19770 (N_19770,N_12659,N_14237);
nor U19771 (N_19771,N_14046,N_14753);
nor U19772 (N_19772,N_14615,N_15046);
or U19773 (N_19773,N_12342,N_12437);
or U19774 (N_19774,N_12764,N_15805);
nor U19775 (N_19775,N_13950,N_13770);
or U19776 (N_19776,N_12908,N_13196);
and U19777 (N_19777,N_12666,N_14656);
nand U19778 (N_19778,N_14939,N_14509);
or U19779 (N_19779,N_15115,N_14710);
and U19780 (N_19780,N_15628,N_15670);
nor U19781 (N_19781,N_13477,N_13211);
or U19782 (N_19782,N_14522,N_13657);
nand U19783 (N_19783,N_13788,N_15677);
nor U19784 (N_19784,N_15311,N_12832);
or U19785 (N_19785,N_13745,N_13264);
nor U19786 (N_19786,N_13424,N_13683);
nand U19787 (N_19787,N_13847,N_13753);
and U19788 (N_19788,N_15333,N_13375);
nand U19789 (N_19789,N_14429,N_14286);
and U19790 (N_19790,N_14442,N_12862);
nor U19791 (N_19791,N_15367,N_14938);
nor U19792 (N_19792,N_13664,N_15926);
nor U19793 (N_19793,N_13569,N_12780);
nor U19794 (N_19794,N_12169,N_14090);
nand U19795 (N_19795,N_12427,N_15061);
and U19796 (N_19796,N_14673,N_12979);
nand U19797 (N_19797,N_13824,N_14015);
nor U19798 (N_19798,N_15619,N_14963);
nand U19799 (N_19799,N_13312,N_14824);
and U19800 (N_19800,N_13634,N_13443);
nor U19801 (N_19801,N_14595,N_15853);
and U19802 (N_19802,N_15796,N_14664);
or U19803 (N_19803,N_12549,N_15964);
nor U19804 (N_19804,N_13598,N_13744);
or U19805 (N_19805,N_13473,N_15957);
nand U19806 (N_19806,N_13586,N_15618);
nand U19807 (N_19807,N_13531,N_14411);
or U19808 (N_19808,N_12657,N_13929);
nor U19809 (N_19809,N_14720,N_13438);
nor U19810 (N_19810,N_13389,N_14020);
xnor U19811 (N_19811,N_12827,N_12649);
nor U19812 (N_19812,N_15729,N_15565);
or U19813 (N_19813,N_12590,N_12626);
and U19814 (N_19814,N_13871,N_15779);
and U19815 (N_19815,N_14621,N_14523);
xnor U19816 (N_19816,N_14787,N_13727);
and U19817 (N_19817,N_12222,N_13012);
nand U19818 (N_19818,N_14504,N_12114);
and U19819 (N_19819,N_14365,N_15694);
and U19820 (N_19820,N_14016,N_12459);
or U19821 (N_19821,N_12751,N_13031);
nor U19822 (N_19822,N_14386,N_15321);
or U19823 (N_19823,N_12551,N_12807);
nor U19824 (N_19824,N_15896,N_14539);
and U19825 (N_19825,N_12988,N_12577);
and U19826 (N_19826,N_15413,N_12527);
nor U19827 (N_19827,N_14965,N_12568);
nor U19828 (N_19828,N_15576,N_14615);
nand U19829 (N_19829,N_14544,N_12186);
nand U19830 (N_19830,N_12085,N_12092);
or U19831 (N_19831,N_14024,N_13149);
nand U19832 (N_19832,N_15386,N_14801);
or U19833 (N_19833,N_13380,N_13226);
and U19834 (N_19834,N_12045,N_14654);
nor U19835 (N_19835,N_13303,N_14986);
or U19836 (N_19836,N_13723,N_14688);
nand U19837 (N_19837,N_13294,N_15791);
nor U19838 (N_19838,N_12717,N_15916);
and U19839 (N_19839,N_14661,N_12869);
and U19840 (N_19840,N_12504,N_14598);
and U19841 (N_19841,N_13354,N_15457);
nor U19842 (N_19842,N_15047,N_13510);
nand U19843 (N_19843,N_13605,N_14995);
nand U19844 (N_19844,N_15622,N_13070);
or U19845 (N_19845,N_13640,N_12340);
nand U19846 (N_19846,N_12498,N_13702);
and U19847 (N_19847,N_15614,N_13605);
and U19848 (N_19848,N_15754,N_14159);
and U19849 (N_19849,N_13645,N_14499);
nor U19850 (N_19850,N_13078,N_12386);
nor U19851 (N_19851,N_15773,N_12387);
nand U19852 (N_19852,N_13341,N_15864);
and U19853 (N_19853,N_13314,N_12383);
and U19854 (N_19854,N_15528,N_14771);
or U19855 (N_19855,N_13336,N_13039);
nor U19856 (N_19856,N_12191,N_15015);
or U19857 (N_19857,N_14414,N_12659);
or U19858 (N_19858,N_12086,N_12949);
or U19859 (N_19859,N_15038,N_12082);
or U19860 (N_19860,N_13018,N_15920);
and U19861 (N_19861,N_12575,N_15417);
nor U19862 (N_19862,N_13229,N_13670);
nand U19863 (N_19863,N_12630,N_15893);
nor U19864 (N_19864,N_12354,N_14564);
and U19865 (N_19865,N_15843,N_14192);
or U19866 (N_19866,N_12876,N_12561);
nand U19867 (N_19867,N_15651,N_13303);
or U19868 (N_19868,N_12256,N_12570);
and U19869 (N_19869,N_14341,N_14380);
nand U19870 (N_19870,N_12109,N_13907);
nor U19871 (N_19871,N_12407,N_12499);
nor U19872 (N_19872,N_12815,N_12954);
or U19873 (N_19873,N_14768,N_13675);
or U19874 (N_19874,N_14270,N_12448);
and U19875 (N_19875,N_12885,N_14957);
nand U19876 (N_19876,N_13231,N_14753);
and U19877 (N_19877,N_12736,N_13733);
and U19878 (N_19878,N_15016,N_15107);
nand U19879 (N_19879,N_12018,N_15969);
and U19880 (N_19880,N_13544,N_12732);
or U19881 (N_19881,N_15622,N_13821);
nand U19882 (N_19882,N_15768,N_15619);
xnor U19883 (N_19883,N_13838,N_12518);
nand U19884 (N_19884,N_14057,N_13121);
nand U19885 (N_19885,N_15194,N_13022);
nor U19886 (N_19886,N_14935,N_12355);
or U19887 (N_19887,N_14082,N_12018);
nand U19888 (N_19888,N_13861,N_12509);
nand U19889 (N_19889,N_12528,N_15884);
and U19890 (N_19890,N_12884,N_14621);
or U19891 (N_19891,N_15854,N_13215);
and U19892 (N_19892,N_14630,N_15064);
and U19893 (N_19893,N_12601,N_14949);
nand U19894 (N_19894,N_14190,N_14256);
or U19895 (N_19895,N_12379,N_14457);
nand U19896 (N_19896,N_13274,N_12075);
nor U19897 (N_19897,N_13011,N_12294);
nor U19898 (N_19898,N_14102,N_13766);
or U19899 (N_19899,N_13245,N_12422);
and U19900 (N_19900,N_14274,N_14366);
or U19901 (N_19901,N_12156,N_13407);
and U19902 (N_19902,N_14872,N_15048);
and U19903 (N_19903,N_12570,N_15743);
nor U19904 (N_19904,N_15164,N_12410);
nand U19905 (N_19905,N_12643,N_13543);
nand U19906 (N_19906,N_12499,N_14548);
nor U19907 (N_19907,N_12166,N_14414);
or U19908 (N_19908,N_12545,N_12362);
or U19909 (N_19909,N_15931,N_15188);
and U19910 (N_19910,N_12856,N_12943);
nor U19911 (N_19911,N_14891,N_15393);
or U19912 (N_19912,N_14095,N_13345);
and U19913 (N_19913,N_15227,N_14312);
nor U19914 (N_19914,N_15376,N_12761);
and U19915 (N_19915,N_15165,N_12088);
and U19916 (N_19916,N_12807,N_14903);
or U19917 (N_19917,N_15507,N_15142);
nand U19918 (N_19918,N_15468,N_15448);
or U19919 (N_19919,N_15236,N_14025);
or U19920 (N_19920,N_15059,N_15817);
xor U19921 (N_19921,N_15144,N_15439);
or U19922 (N_19922,N_15847,N_14927);
and U19923 (N_19923,N_12217,N_12517);
or U19924 (N_19924,N_15732,N_15883);
nor U19925 (N_19925,N_14123,N_12574);
nor U19926 (N_19926,N_13527,N_13036);
and U19927 (N_19927,N_12049,N_13152);
and U19928 (N_19928,N_15047,N_14886);
nor U19929 (N_19929,N_15949,N_13638);
and U19930 (N_19930,N_12377,N_14777);
nand U19931 (N_19931,N_15248,N_12705);
nor U19932 (N_19932,N_14005,N_15153);
or U19933 (N_19933,N_15379,N_13727);
nand U19934 (N_19934,N_13290,N_15754);
nor U19935 (N_19935,N_12970,N_13508);
and U19936 (N_19936,N_13400,N_14720);
nand U19937 (N_19937,N_14104,N_15062);
nor U19938 (N_19938,N_12990,N_13828);
or U19939 (N_19939,N_13759,N_14096);
and U19940 (N_19940,N_15791,N_14914);
nand U19941 (N_19941,N_15495,N_15796);
and U19942 (N_19942,N_15451,N_12688);
and U19943 (N_19943,N_12323,N_12914);
or U19944 (N_19944,N_12995,N_15144);
nand U19945 (N_19945,N_12973,N_15935);
and U19946 (N_19946,N_14425,N_12740);
and U19947 (N_19947,N_15426,N_14089);
nand U19948 (N_19948,N_13802,N_15498);
nor U19949 (N_19949,N_15622,N_12112);
and U19950 (N_19950,N_13500,N_14094);
nand U19951 (N_19951,N_12740,N_12789);
nor U19952 (N_19952,N_15383,N_13621);
or U19953 (N_19953,N_12790,N_12765);
nor U19954 (N_19954,N_14944,N_14743);
or U19955 (N_19955,N_14474,N_12958);
nor U19956 (N_19956,N_12832,N_12805);
nand U19957 (N_19957,N_15081,N_13141);
nand U19958 (N_19958,N_15493,N_14189);
nand U19959 (N_19959,N_15096,N_12246);
or U19960 (N_19960,N_15231,N_15204);
or U19961 (N_19961,N_13145,N_14734);
nor U19962 (N_19962,N_15293,N_13147);
or U19963 (N_19963,N_13564,N_14229);
nand U19964 (N_19964,N_15139,N_13904);
or U19965 (N_19965,N_15045,N_15804);
nand U19966 (N_19966,N_12699,N_15600);
or U19967 (N_19967,N_13841,N_12377);
nand U19968 (N_19968,N_14188,N_12947);
nand U19969 (N_19969,N_13025,N_12210);
nand U19970 (N_19970,N_15050,N_13099);
nor U19971 (N_19971,N_13681,N_13612);
or U19972 (N_19972,N_14722,N_14843);
nor U19973 (N_19973,N_14358,N_15776);
or U19974 (N_19974,N_12303,N_12587);
xor U19975 (N_19975,N_15860,N_13672);
nor U19976 (N_19976,N_12896,N_14084);
and U19977 (N_19977,N_14877,N_14114);
nand U19978 (N_19978,N_15337,N_13034);
nor U19979 (N_19979,N_15312,N_15717);
nand U19980 (N_19980,N_15605,N_12925);
or U19981 (N_19981,N_12536,N_15743);
or U19982 (N_19982,N_14652,N_15957);
or U19983 (N_19983,N_13408,N_15867);
and U19984 (N_19984,N_13285,N_15513);
nand U19985 (N_19985,N_12088,N_13810);
and U19986 (N_19986,N_13570,N_15915);
and U19987 (N_19987,N_15623,N_15192);
nand U19988 (N_19988,N_12030,N_13487);
nor U19989 (N_19989,N_15371,N_13918);
or U19990 (N_19990,N_12236,N_13223);
nor U19991 (N_19991,N_12634,N_14298);
and U19992 (N_19992,N_12272,N_15110);
nand U19993 (N_19993,N_13448,N_12162);
and U19994 (N_19994,N_13650,N_14142);
nor U19995 (N_19995,N_13543,N_14020);
nand U19996 (N_19996,N_12778,N_12851);
nand U19997 (N_19997,N_12729,N_14178);
or U19998 (N_19998,N_12867,N_15725);
nand U19999 (N_19999,N_14369,N_13290);
nor UO_0 (O_0,N_16672,N_18964);
and UO_1 (O_1,N_17790,N_19611);
nor UO_2 (O_2,N_17889,N_18685);
or UO_3 (O_3,N_16553,N_16358);
nand UO_4 (O_4,N_19779,N_19187);
nor UO_5 (O_5,N_16886,N_17041);
and UO_6 (O_6,N_17312,N_17179);
and UO_7 (O_7,N_17574,N_19952);
nand UO_8 (O_8,N_17820,N_19425);
and UO_9 (O_9,N_17252,N_17181);
nor UO_10 (O_10,N_19212,N_19572);
nor UO_11 (O_11,N_17188,N_19918);
or UO_12 (O_12,N_19290,N_17713);
or UO_13 (O_13,N_16381,N_16854);
nand UO_14 (O_14,N_18032,N_18106);
and UO_15 (O_15,N_16624,N_18804);
and UO_16 (O_16,N_16030,N_18723);
nor UO_17 (O_17,N_17388,N_18122);
and UO_18 (O_18,N_18761,N_16359);
nor UO_19 (O_19,N_17618,N_18515);
and UO_20 (O_20,N_19402,N_17765);
and UO_21 (O_21,N_16528,N_19055);
nand UO_22 (O_22,N_19692,N_18780);
nand UO_23 (O_23,N_19798,N_19942);
and UO_24 (O_24,N_16267,N_17381);
and UO_25 (O_25,N_17784,N_17907);
nand UO_26 (O_26,N_16939,N_16995);
or UO_27 (O_27,N_17610,N_16552);
and UO_28 (O_28,N_18824,N_16903);
nor UO_29 (O_29,N_17238,N_19241);
nor UO_30 (O_30,N_17888,N_16668);
nor UO_31 (O_31,N_16159,N_16439);
and UO_32 (O_32,N_19500,N_16154);
nor UO_33 (O_33,N_19658,N_19309);
and UO_34 (O_34,N_18437,N_18086);
and UO_35 (O_35,N_17552,N_18033);
nor UO_36 (O_36,N_18543,N_16520);
nand UO_37 (O_37,N_18477,N_17852);
and UO_38 (O_38,N_18468,N_17902);
nor UO_39 (O_39,N_17687,N_16702);
nand UO_40 (O_40,N_17952,N_17835);
nand UO_41 (O_41,N_19549,N_17014);
nand UO_42 (O_42,N_18221,N_16636);
or UO_43 (O_43,N_16867,N_19263);
and UO_44 (O_44,N_16996,N_19122);
or UO_45 (O_45,N_17350,N_16949);
nor UO_46 (O_46,N_19132,N_17498);
nand UO_47 (O_47,N_18598,N_19144);
and UO_48 (O_48,N_17331,N_19824);
nor UO_49 (O_49,N_18559,N_16402);
or UO_50 (O_50,N_17385,N_16410);
and UO_51 (O_51,N_16301,N_16776);
or UO_52 (O_52,N_17085,N_16306);
or UO_53 (O_53,N_17060,N_18966);
nand UO_54 (O_54,N_17021,N_17123);
and UO_55 (O_55,N_18999,N_17577);
nor UO_56 (O_56,N_18381,N_18548);
nand UO_57 (O_57,N_18314,N_16050);
nand UO_58 (O_58,N_17037,N_18014);
nand UO_59 (O_59,N_17148,N_17348);
and UO_60 (O_60,N_17472,N_17424);
and UO_61 (O_61,N_16872,N_19818);
or UO_62 (O_62,N_18442,N_19321);
nor UO_63 (O_63,N_19073,N_18390);
or UO_64 (O_64,N_16827,N_18718);
nand UO_65 (O_65,N_18427,N_16254);
and UO_66 (O_66,N_17196,N_19322);
nand UO_67 (O_67,N_16608,N_16370);
and UO_68 (O_68,N_16394,N_19537);
or UO_69 (O_69,N_19603,N_19415);
and UO_70 (O_70,N_16184,N_18710);
nor UO_71 (O_71,N_19388,N_19650);
nand UO_72 (O_72,N_19174,N_17370);
or UO_73 (O_73,N_16491,N_16025);
nor UO_74 (O_74,N_17058,N_16190);
or UO_75 (O_75,N_18197,N_17342);
nor UO_76 (O_76,N_18520,N_18443);
or UO_77 (O_77,N_19784,N_19334);
and UO_78 (O_78,N_17440,N_16384);
or UO_79 (O_79,N_19018,N_17065);
or UO_80 (O_80,N_16689,N_19738);
and UO_81 (O_81,N_18717,N_17579);
or UO_82 (O_82,N_17262,N_19510);
or UO_83 (O_83,N_18798,N_16281);
nor UO_84 (O_84,N_16659,N_18184);
nand UO_85 (O_85,N_18213,N_16131);
or UO_86 (O_86,N_16928,N_16779);
or UO_87 (O_87,N_16725,N_17475);
nand UO_88 (O_88,N_18792,N_19991);
and UO_89 (O_89,N_17554,N_19993);
nand UO_90 (O_90,N_18361,N_18943);
and UO_91 (O_91,N_17207,N_16514);
or UO_92 (O_92,N_18251,N_17647);
nor UO_93 (O_93,N_16695,N_18216);
nor UO_94 (O_94,N_19314,N_17711);
nand UO_95 (O_95,N_17946,N_18592);
xnor UO_96 (O_96,N_18340,N_18174);
and UO_97 (O_97,N_19027,N_17176);
nand UO_98 (O_98,N_16752,N_17575);
and UO_99 (O_99,N_19637,N_16183);
or UO_100 (O_100,N_19639,N_16517);
and UO_101 (O_101,N_17091,N_19473);
or UO_102 (O_102,N_19459,N_18590);
nor UO_103 (O_103,N_19028,N_17456);
nor UO_104 (O_104,N_16133,N_18228);
and UO_105 (O_105,N_17212,N_17221);
and UO_106 (O_106,N_19717,N_18787);
and UO_107 (O_107,N_16162,N_16821);
and UO_108 (O_108,N_17443,N_16878);
or UO_109 (O_109,N_18489,N_18281);
nor UO_110 (O_110,N_17879,N_18406);
and UO_111 (O_111,N_17555,N_19147);
or UO_112 (O_112,N_17706,N_18752);
and UO_113 (O_113,N_19305,N_18451);
or UO_114 (O_114,N_16242,N_18985);
and UO_115 (O_115,N_16972,N_18410);
nor UO_116 (O_116,N_19195,N_16238);
xor UO_117 (O_117,N_18732,N_17022);
nand UO_118 (O_118,N_18560,N_18807);
nand UO_119 (O_119,N_19463,N_16753);
nand UO_120 (O_120,N_17049,N_17024);
or UO_121 (O_121,N_19235,N_19119);
or UO_122 (O_122,N_17770,N_19990);
nand UO_123 (O_123,N_19412,N_17121);
or UO_124 (O_124,N_17264,N_19137);
nand UO_125 (O_125,N_16052,N_16096);
or UO_126 (O_126,N_19169,N_16942);
and UO_127 (O_127,N_19328,N_16834);
or UO_128 (O_128,N_19781,N_18909);
nand UO_129 (O_129,N_17629,N_19173);
and UO_130 (O_130,N_18055,N_19360);
and UO_131 (O_131,N_16625,N_19703);
and UO_132 (O_132,N_16182,N_16351);
nand UO_133 (O_133,N_16563,N_16701);
or UO_134 (O_134,N_19103,N_16033);
nand UO_135 (O_135,N_17066,N_18554);
nor UO_136 (O_136,N_16156,N_17408);
or UO_137 (O_137,N_18739,N_16271);
nor UO_138 (O_138,N_17634,N_17566);
nor UO_139 (O_139,N_16897,N_19563);
nor UO_140 (O_140,N_19876,N_19504);
and UO_141 (O_141,N_17046,N_19377);
nor UO_142 (O_142,N_17752,N_17254);
or UO_143 (O_143,N_19795,N_19281);
and UO_144 (O_144,N_16164,N_18687);
nor UO_145 (O_145,N_16791,N_18386);
or UO_146 (O_146,N_16168,N_16051);
or UO_147 (O_147,N_17457,N_16290);
nand UO_148 (O_148,N_18384,N_18104);
and UO_149 (O_149,N_18445,N_16270);
or UO_150 (O_150,N_17860,N_16613);
or UO_151 (O_151,N_18425,N_18902);
nand UO_152 (O_152,N_18929,N_18015);
nor UO_153 (O_153,N_16469,N_17116);
nand UO_154 (O_154,N_18848,N_17129);
nor UO_155 (O_155,N_16259,N_18250);
nor UO_156 (O_156,N_17728,N_18273);
or UO_157 (O_157,N_18796,N_19750);
and UO_158 (O_158,N_17904,N_16814);
nor UO_159 (O_159,N_19105,N_16365);
xor UO_160 (O_160,N_18846,N_16951);
nand UO_161 (O_161,N_16587,N_17195);
nand UO_162 (O_162,N_16602,N_19594);
and UO_163 (O_163,N_19614,N_18911);
nor UO_164 (O_164,N_17451,N_18479);
nand UO_165 (O_165,N_18118,N_19701);
nor UO_166 (O_166,N_19668,N_16774);
or UO_167 (O_167,N_19357,N_16294);
and UO_168 (O_168,N_17096,N_16097);
or UO_169 (O_169,N_18223,N_19323);
nand UO_170 (O_170,N_18376,N_17467);
or UO_171 (O_171,N_16577,N_18293);
and UO_172 (O_172,N_17093,N_18756);
and UO_173 (O_173,N_19864,N_19411);
nor UO_174 (O_174,N_18593,N_18639);
nand UO_175 (O_175,N_17736,N_19862);
and UO_176 (O_176,N_18860,N_17643);
or UO_177 (O_177,N_18450,N_19722);
and UO_178 (O_178,N_18359,N_17444);
and UO_179 (O_179,N_19871,N_16031);
nand UO_180 (O_180,N_19436,N_16667);
and UO_181 (O_181,N_19109,N_19673);
and UO_182 (O_182,N_16148,N_16020);
nand UO_183 (O_183,N_18716,N_17341);
and UO_184 (O_184,N_17168,N_16628);
nand UO_185 (O_185,N_16506,N_17507);
nand UO_186 (O_186,N_16008,N_18936);
nand UO_187 (O_187,N_16409,N_19176);
nor UO_188 (O_188,N_16649,N_19589);
or UO_189 (O_189,N_18364,N_19514);
nor UO_190 (O_190,N_18036,N_18636);
xnor UO_191 (O_191,N_16251,N_17246);
or UO_192 (O_192,N_19139,N_19118);
or UO_193 (O_193,N_18031,N_16495);
or UO_194 (O_194,N_18185,N_18960);
nand UO_195 (O_195,N_19769,N_19488);
nand UO_196 (O_196,N_18480,N_16149);
and UO_197 (O_197,N_17158,N_16129);
or UO_198 (O_198,N_18857,N_17773);
nand UO_199 (O_199,N_16805,N_17681);
or UO_200 (O_200,N_16245,N_16125);
nor UO_201 (O_201,N_17817,N_19928);
or UO_202 (O_202,N_18662,N_19215);
or UO_203 (O_203,N_18083,N_19479);
nor UO_204 (O_204,N_19586,N_18316);
nand UO_205 (O_205,N_16798,N_17340);
xnor UO_206 (O_206,N_16161,N_19878);
nand UO_207 (O_207,N_17361,N_19880);
or UO_208 (O_208,N_17882,N_18694);
nand UO_209 (O_209,N_18283,N_16795);
nand UO_210 (O_210,N_19896,N_17110);
nand UO_211 (O_211,N_19354,N_17418);
and UO_212 (O_212,N_17015,N_19995);
or UO_213 (O_213,N_17847,N_17992);
or UO_214 (O_214,N_16079,N_16457);
nor UO_215 (O_215,N_18574,N_18170);
or UO_216 (O_216,N_16176,N_18510);
xor UO_217 (O_217,N_19346,N_16645);
and UO_218 (O_218,N_17814,N_19006);
or UO_219 (O_219,N_17949,N_19529);
or UO_220 (O_220,N_18538,N_18166);
and UO_221 (O_221,N_16952,N_17901);
and UO_222 (O_222,N_16492,N_19050);
or UO_223 (O_223,N_16990,N_18195);
nor UO_224 (O_224,N_17004,N_18850);
and UO_225 (O_225,N_17193,N_19753);
nand UO_226 (O_226,N_19929,N_17442);
nand UO_227 (O_227,N_19295,N_16320);
and UO_228 (O_228,N_16015,N_18614);
nand UO_229 (O_229,N_16111,N_18342);
nand UO_230 (O_230,N_19216,N_18308);
nor UO_231 (O_231,N_19909,N_16089);
and UO_232 (O_232,N_16062,N_16465);
nand UO_233 (O_233,N_19816,N_16198);
nor UO_234 (O_234,N_19455,N_16444);
xnor UO_235 (O_235,N_19131,N_18757);
nand UO_236 (O_236,N_17293,N_16948);
or UO_237 (O_237,N_19407,N_19149);
nand UO_238 (O_238,N_16157,N_17649);
and UO_239 (O_239,N_18226,N_16765);
nor UO_240 (O_240,N_16706,N_17987);
nor UO_241 (O_241,N_17375,N_16797);
or UO_242 (O_242,N_17153,N_16071);
or UO_243 (O_243,N_19945,N_19924);
or UO_244 (O_244,N_17874,N_19934);
or UO_245 (O_245,N_18493,N_19868);
or UO_246 (O_246,N_19957,N_19861);
nor UO_247 (O_247,N_18144,N_17655);
or UO_248 (O_248,N_16113,N_18894);
nor UO_249 (O_249,N_19792,N_19442);
nand UO_250 (O_250,N_18358,N_18151);
or UO_251 (O_251,N_16905,N_18832);
and UO_252 (O_252,N_18157,N_16039);
or UO_253 (O_253,N_17255,N_18374);
nand UO_254 (O_254,N_16677,N_16155);
nand UO_255 (O_255,N_17347,N_18217);
nand UO_256 (O_256,N_18124,N_19256);
nand UO_257 (O_257,N_16865,N_18534);
or UO_258 (O_258,N_16200,N_18641);
or UO_259 (O_259,N_18891,N_16219);
or UO_260 (O_260,N_17934,N_18490);
nand UO_261 (O_261,N_16327,N_19731);
nor UO_262 (O_262,N_17415,N_18870);
and UO_263 (O_263,N_16312,N_18663);
nor UO_264 (O_264,N_19202,N_16311);
nor UO_265 (O_265,N_18986,N_17540);
nor UO_266 (O_266,N_19237,N_16021);
nor UO_267 (O_267,N_16060,N_16041);
and UO_268 (O_268,N_18677,N_16375);
nor UO_269 (O_269,N_16575,N_16167);
nand UO_270 (O_270,N_17591,N_16704);
nor UO_271 (O_271,N_17229,N_16570);
and UO_272 (O_272,N_16782,N_19844);
or UO_273 (O_273,N_16241,N_16237);
and UO_274 (O_274,N_17758,N_17446);
nor UO_275 (O_275,N_19483,N_16697);
or UO_276 (O_276,N_18577,N_17755);
nor UO_277 (O_277,N_18191,N_16106);
nor UO_278 (O_278,N_17799,N_16102);
nand UO_279 (O_279,N_16804,N_18294);
nor UO_280 (O_280,N_19218,N_19944);
and UO_281 (O_281,N_19183,N_19114);
or UO_282 (O_282,N_18193,N_19946);
and UO_283 (O_283,N_17912,N_17725);
nor UO_284 (O_284,N_17559,N_16336);
nand UO_285 (O_285,N_18017,N_17623);
nor UO_286 (O_286,N_17178,N_19214);
or UO_287 (O_287,N_19533,N_16501);
nand UO_288 (O_288,N_17957,N_18212);
xor UO_289 (O_289,N_18512,N_17163);
or UO_290 (O_290,N_17202,N_19715);
and UO_291 (O_291,N_18957,N_16547);
nor UO_292 (O_292,N_19582,N_16346);
and UO_293 (O_293,N_18454,N_17132);
and UO_294 (O_294,N_16158,N_17514);
nor UO_295 (O_295,N_19624,N_18621);
and UO_296 (O_296,N_17300,N_16775);
or UO_297 (O_297,N_18939,N_18146);
and UO_298 (O_298,N_19794,N_17420);
nor UO_299 (O_299,N_19056,N_19293);
nand UO_300 (O_300,N_16635,N_18934);
nand UO_301 (O_301,N_16787,N_16266);
or UO_302 (O_302,N_19919,N_17972);
and UO_303 (O_303,N_18127,N_17526);
or UO_304 (O_304,N_19505,N_16236);
nor UO_305 (O_305,N_16973,N_16944);
xor UO_306 (O_306,N_18051,N_19793);
nand UO_307 (O_307,N_19828,N_17208);
nand UO_308 (O_308,N_19168,N_17117);
xor UO_309 (O_309,N_18279,N_18601);
or UO_310 (O_310,N_19487,N_18516);
nand UO_311 (O_311,N_16512,N_16048);
or UO_312 (O_312,N_18402,N_16152);
or UO_313 (O_313,N_18186,N_16314);
xor UO_314 (O_314,N_19016,N_18502);
and UO_315 (O_315,N_17945,N_19696);
and UO_316 (O_316,N_17541,N_18789);
and UO_317 (O_317,N_19219,N_18942);
and UO_318 (O_318,N_17989,N_19048);
or UO_319 (O_319,N_17596,N_18916);
and UO_320 (O_320,N_18123,N_16656);
nand UO_321 (O_321,N_16144,N_19426);
nor UO_322 (O_322,N_16045,N_19822);
nand UO_323 (O_323,N_18299,N_17286);
or UO_324 (O_324,N_16476,N_16616);
nand UO_325 (O_325,N_17700,N_17712);
and UO_326 (O_326,N_17005,N_19983);
and UO_327 (O_327,N_16172,N_16601);
or UO_328 (O_328,N_19665,N_17678);
nor UO_329 (O_329,N_17894,N_17106);
or UO_330 (O_330,N_17997,N_16429);
or UO_331 (O_331,N_19675,N_16524);
and UO_332 (O_332,N_19242,N_16746);
nand UO_333 (O_333,N_18499,N_16844);
or UO_334 (O_334,N_19842,N_19920);
or UO_335 (O_335,N_17809,N_16186);
and UO_336 (O_336,N_18712,N_17669);
and UO_337 (O_337,N_17651,N_17829);
xor UO_338 (O_338,N_16348,N_16521);
nand UO_339 (O_339,N_16206,N_18434);
or UO_340 (O_340,N_17701,N_19813);
or UO_341 (O_341,N_17143,N_18484);
nand UO_342 (O_342,N_17473,N_18674);
nor UO_343 (O_343,N_16377,N_19152);
nor UO_344 (O_344,N_16840,N_16315);
nand UO_345 (O_345,N_16417,N_18001);
and UO_346 (O_346,N_18951,N_18878);
or UO_347 (O_347,N_18486,N_19954);
nor UO_348 (O_348,N_17886,N_19347);
nand UO_349 (O_349,N_17914,N_19181);
nor UO_350 (O_350,N_16945,N_16059);
nand UO_351 (O_351,N_19493,N_18682);
nand UO_352 (O_352,N_18062,N_19023);
nor UO_353 (O_353,N_17365,N_18422);
nor UO_354 (O_354,N_16177,N_16115);
nand UO_355 (O_355,N_17013,N_17253);
and UO_356 (O_356,N_17920,N_16964);
nand UO_357 (O_357,N_18054,N_17307);
and UO_358 (O_358,N_17434,N_16374);
and UO_359 (O_359,N_17357,N_19517);
or UO_360 (O_360,N_17944,N_18653);
and UO_361 (O_361,N_18115,N_17558);
and UO_362 (O_362,N_19200,N_18919);
nand UO_363 (O_363,N_18136,N_16808);
and UO_364 (O_364,N_17219,N_18533);
nor UO_365 (O_365,N_18139,N_18416);
nor UO_366 (O_366,N_18130,N_17052);
and UO_367 (O_367,N_17818,N_19106);
or UO_368 (O_368,N_17787,N_16451);
nand UO_369 (O_369,N_18762,N_16666);
nor UO_370 (O_370,N_18976,N_18814);
and UO_371 (O_371,N_18389,N_16953);
nand UO_372 (O_372,N_18050,N_18781);
nand UO_373 (O_373,N_16698,N_17384);
nand UO_374 (O_374,N_17810,N_17236);
xor UO_375 (O_375,N_19233,N_19496);
nand UO_376 (O_376,N_18926,N_17162);
nor UO_377 (O_377,N_16389,N_16406);
and UO_378 (O_378,N_18931,N_16591);
and UO_379 (O_379,N_17968,N_18194);
nor UO_380 (O_380,N_17637,N_17975);
nor UO_381 (O_381,N_19799,N_19905);
nand UO_382 (O_382,N_19339,N_16076);
or UO_383 (O_383,N_19422,N_18765);
xnor UO_384 (O_384,N_19390,N_18012);
or UO_385 (O_385,N_18688,N_19331);
nand UO_386 (O_386,N_16582,N_16818);
nand UO_387 (O_387,N_18096,N_18834);
nor UO_388 (O_388,N_16383,N_18180);
xnor UO_389 (O_389,N_17607,N_17595);
or UO_390 (O_390,N_18369,N_16299);
nand UO_391 (O_391,N_19060,N_16369);
nor UO_392 (O_392,N_19034,N_18037);
nand UO_393 (O_393,N_16195,N_19561);
and UO_394 (O_394,N_19026,N_19626);
nor UO_395 (O_395,N_16907,N_17263);
nor UO_396 (O_396,N_19689,N_17848);
nor UO_397 (O_397,N_18282,N_17156);
nand UO_398 (O_398,N_19881,N_16009);
and UO_399 (O_399,N_19270,N_16906);
and UO_400 (O_400,N_18269,N_16362);
or UO_401 (O_401,N_19497,N_17265);
and UO_402 (O_402,N_18994,N_17853);
nor UO_403 (O_403,N_19975,N_16934);
nand UO_404 (O_404,N_16550,N_19210);
and UO_405 (O_405,N_18624,N_19443);
nand UO_406 (O_406,N_19349,N_19869);
and UO_407 (O_407,N_18457,N_16622);
nor UO_408 (O_408,N_19058,N_16163);
xor UO_409 (O_409,N_19428,N_16678);
nor UO_410 (O_410,N_17985,N_17867);
or UO_411 (O_411,N_18084,N_18722);
and UO_412 (O_412,N_19959,N_16825);
nor UO_413 (O_413,N_17648,N_16594);
or UO_414 (O_414,N_18690,N_18801);
or UO_415 (O_415,N_19516,N_16817);
nand UO_416 (O_416,N_16839,N_17460);
nand UO_417 (O_417,N_17023,N_16966);
nor UO_418 (O_418,N_17259,N_17812);
nand UO_419 (O_419,N_19134,N_19068);
and UO_420 (O_420,N_17506,N_18081);
nor UO_421 (O_421,N_19171,N_17576);
nand UO_422 (O_422,N_16005,N_17239);
nand UO_423 (O_423,N_17329,N_16340);
and UO_424 (O_424,N_18530,N_17922);
nor UO_425 (O_425,N_16118,N_19145);
and UO_426 (O_426,N_18736,N_16700);
nand UO_427 (O_427,N_17161,N_16954);
or UO_428 (O_428,N_16070,N_17421);
and UO_429 (O_429,N_18280,N_19299);
and UO_430 (O_430,N_19469,N_16705);
nor UO_431 (O_431,N_16056,N_16785);
nand UO_432 (O_432,N_18959,N_19100);
or UO_433 (O_433,N_17210,N_18049);
and UO_434 (O_434,N_16876,N_19012);
or UO_435 (O_435,N_16018,N_16502);
and UO_436 (O_436,N_16720,N_19079);
nand UO_437 (O_437,N_19306,N_19904);
and UO_438 (O_438,N_16571,N_18309);
and UO_439 (O_439,N_18921,N_19344);
and UO_440 (O_440,N_17534,N_17371);
nor UO_441 (O_441,N_17599,N_16412);
or UO_442 (O_442,N_19985,N_16038);
nand UO_443 (O_443,N_18551,N_17288);
or UO_444 (O_444,N_19608,N_16826);
or UO_445 (O_445,N_18529,N_19951);
nor UO_446 (O_446,N_18702,N_16484);
and UO_447 (O_447,N_17291,N_16755);
or UO_448 (O_448,N_17877,N_19752);
nor UO_449 (O_449,N_18209,N_18259);
or UO_450 (O_450,N_19859,N_18793);
nor UO_451 (O_451,N_17744,N_16407);
or UO_452 (O_452,N_17645,N_18896);
nor UO_453 (O_453,N_17282,N_16603);
or UO_454 (O_454,N_19686,N_18844);
and UO_455 (O_455,N_18405,N_17646);
and UO_456 (O_456,N_17226,N_19156);
nand UO_457 (O_457,N_18108,N_17636);
and UO_458 (O_458,N_18067,N_19398);
nor UO_459 (O_459,N_16043,N_17602);
nor UO_460 (O_460,N_17796,N_19254);
nand UO_461 (O_461,N_17154,N_19432);
nor UO_462 (O_462,N_19318,N_16082);
and UO_463 (O_463,N_17380,N_18331);
and UO_464 (O_464,N_16077,N_17466);
or UO_465 (O_465,N_16404,N_19401);
nor UO_466 (O_466,N_19629,N_17167);
and UO_467 (O_467,N_18803,N_18160);
nor UO_468 (O_468,N_17503,N_17099);
nand UO_469 (O_469,N_19645,N_17974);
or UO_470 (O_470,N_16803,N_16380);
nor UO_471 (O_471,N_16555,N_18073);
nand UO_472 (O_472,N_19705,N_18383);
nor UO_473 (O_473,N_17292,N_17978);
or UO_474 (O_474,N_18275,N_16764);
and UO_475 (O_475,N_19036,N_18946);
nor UO_476 (O_476,N_18159,N_16819);
or UO_477 (O_477,N_18058,N_19565);
and UO_478 (O_478,N_17959,N_17830);
nand UO_479 (O_479,N_16307,N_17626);
nor UO_480 (O_480,N_17501,N_18557);
nor UO_481 (O_481,N_19568,N_17330);
and UO_482 (O_482,N_19341,N_19950);
and UO_483 (O_483,N_17831,N_18910);
nor UO_484 (O_484,N_18107,N_17727);
nand UO_485 (O_485,N_19039,N_17751);
xnor UO_486 (O_486,N_19627,N_19728);
or UO_487 (O_487,N_19564,N_19045);
or UO_488 (O_488,N_17125,N_19431);
and UO_489 (O_489,N_16621,N_18060);
nand UO_490 (O_490,N_16970,N_18693);
or UO_491 (O_491,N_19730,N_19421);
nand UO_492 (O_492,N_16109,N_19833);
nand UO_493 (O_493,N_16049,N_18776);
nor UO_494 (O_494,N_19054,N_18989);
and UO_495 (O_495,N_17598,N_18046);
nand UO_496 (O_496,N_17604,N_17395);
and UO_497 (O_497,N_18021,N_17857);
and UO_498 (O_498,N_16280,N_19783);
nand UO_499 (O_499,N_18928,N_17851);
or UO_500 (O_500,N_19345,N_18238);
and UO_501 (O_501,N_19269,N_16640);
xor UO_502 (O_502,N_17967,N_19638);
nand UO_503 (O_503,N_19316,N_19684);
or UO_504 (O_504,N_16499,N_16345);
or UO_505 (O_505,N_17759,N_18320);
and UO_506 (O_506,N_19811,N_17363);
or UO_507 (O_507,N_18119,N_18211);
xor UO_508 (O_508,N_17726,N_18513);
nand UO_509 (O_509,N_19462,N_18887);
nand UO_510 (O_510,N_16946,N_16846);
or UO_511 (O_511,N_17275,N_16470);
or UO_512 (O_512,N_19856,N_19203);
or UO_513 (O_513,N_19980,N_16122);
nor UO_514 (O_514,N_19695,N_19451);
nor UO_515 (O_515,N_19926,N_19372);
or UO_516 (O_516,N_18013,N_17801);
or UO_517 (O_517,N_17050,N_17224);
nor UO_518 (O_518,N_18272,N_16851);
and UO_519 (O_519,N_17280,N_18222);
nor UO_520 (O_520,N_16017,N_16910);
nand UO_521 (O_521,N_16904,N_19337);
and UO_522 (O_522,N_16661,N_17025);
nor UO_523 (O_523,N_18378,N_17101);
and UO_524 (O_524,N_17225,N_17892);
nor UO_525 (O_525,N_18905,N_18845);
nand UO_526 (O_526,N_17743,N_18968);
nor UO_527 (O_527,N_16343,N_17209);
nand UO_528 (O_528,N_16478,N_17754);
and UO_529 (O_529,N_19076,N_17969);
nand UO_530 (O_530,N_19146,N_19808);
nand UO_531 (O_531,N_17432,N_18821);
and UO_532 (O_532,N_19646,N_18676);
nand UO_533 (O_533,N_17142,N_18362);
or UO_534 (O_534,N_19143,N_19083);
or UO_535 (O_535,N_19445,N_17299);
or UO_536 (O_536,N_17438,N_19265);
nand UO_537 (O_537,N_19576,N_17074);
and UO_538 (O_538,N_18284,N_18366);
nor UO_539 (O_539,N_17337,N_18315);
and UO_540 (O_540,N_17990,N_16449);
or UO_541 (O_541,N_18063,N_19704);
or UO_542 (O_542,N_16274,N_17469);
nor UO_543 (O_543,N_16729,N_17359);
and UO_544 (O_544,N_17245,N_18915);
nor UO_545 (O_545,N_17827,N_16998);
or UO_546 (O_546,N_16807,N_17753);
nand UO_547 (O_547,N_18313,N_16835);
nand UO_548 (O_548,N_16372,N_18167);
or UO_549 (O_549,N_16806,N_18698);
or UO_550 (O_550,N_19330,N_17377);
and UO_551 (O_551,N_17397,N_19204);
nor UO_552 (O_552,N_16091,N_17913);
or UO_553 (O_553,N_19153,N_16813);
nor UO_554 (O_554,N_18290,N_16396);
nor UO_555 (O_555,N_16321,N_17563);
nor UO_556 (O_556,N_17398,N_16534);
or UO_557 (O_557,N_18511,N_16887);
and UO_558 (O_558,N_18330,N_17980);
and UO_559 (O_559,N_16626,N_19471);
and UO_560 (O_560,N_18317,N_18758);
or UO_561 (O_561,N_19759,N_17319);
nand UO_562 (O_562,N_17791,N_18982);
nand UO_563 (O_563,N_19763,N_17935);
nor UO_564 (O_564,N_16974,N_17568);
or UO_565 (O_565,N_18882,N_19770);
nand UO_566 (O_566,N_19826,N_19960);
and UO_567 (O_567,N_18148,N_17031);
and UO_568 (O_568,N_16318,N_19352);
and UO_569 (O_569,N_17258,N_18439);
or UO_570 (O_570,N_17211,N_19840);
nand UO_571 (O_571,N_19829,N_17030);
and UO_572 (O_572,N_19380,N_19656);
and UO_573 (O_573,N_17057,N_17413);
xor UO_574 (O_574,N_17216,N_17256);
or UO_575 (O_575,N_16249,N_18572);
or UO_576 (O_576,N_19727,N_19849);
nand UO_577 (O_577,N_16816,N_16715);
and UO_578 (O_578,N_18553,N_19700);
nor UO_579 (O_579,N_18679,N_19266);
and UO_580 (O_580,N_18231,N_17931);
nand UO_581 (O_581,N_16099,N_19378);
nand UO_582 (O_582,N_16273,N_17274);
and UO_583 (O_583,N_19417,N_17793);
or UO_584 (O_584,N_18669,N_19807);
nand UO_585 (O_585,N_17730,N_17399);
nor UO_586 (O_586,N_17390,N_16739);
nor UO_587 (O_587,N_16800,N_16713);
nand UO_588 (O_588,N_18885,N_16576);
and UO_589 (O_589,N_18204,N_19198);
nand UO_590 (O_590,N_19963,N_17538);
and UO_591 (O_591,N_17779,N_16812);
nand UO_592 (O_592,N_19581,N_17864);
xor UO_593 (O_593,N_17749,N_17905);
nand UO_594 (O_594,N_16975,N_16302);
and UO_595 (O_595,N_17441,N_16319);
and UO_596 (O_596,N_16291,N_16831);
or UO_597 (O_597,N_16726,N_17313);
and UO_598 (O_598,N_16455,N_16277);
nor UO_599 (O_599,N_19854,N_17105);
nor UO_600 (O_600,N_19518,N_17657);
or UO_601 (O_601,N_17002,N_16992);
nor UO_602 (O_602,N_17476,N_19662);
and UO_603 (O_603,N_19771,N_19512);
and UO_604 (O_604,N_18099,N_19782);
nor UO_605 (O_605,N_17953,N_18345);
nand UO_606 (O_606,N_18802,N_19806);
or UO_607 (O_607,N_19282,N_19447);
or UO_608 (O_608,N_19931,N_19754);
nand UO_609 (O_609,N_18729,N_18790);
or UO_610 (O_610,N_18699,N_18901);
xor UO_611 (O_611,N_16742,N_16386);
or UO_612 (O_612,N_16557,N_16744);
nand UO_613 (O_613,N_18088,N_18089);
nand UO_614 (O_614,N_16898,N_16895);
nor UO_615 (O_615,N_16395,N_16324);
nand UO_616 (O_616,N_18234,N_16920);
nand UO_617 (O_617,N_17463,N_18686);
nand UO_618 (O_618,N_16884,N_19786);
nand UO_619 (O_619,N_16650,N_19418);
and UO_620 (O_620,N_19165,N_19562);
or UO_621 (O_621,N_16860,N_17660);
or UO_622 (O_622,N_18353,N_19391);
nand UO_623 (O_623,N_19597,N_16823);
and UO_624 (O_624,N_16403,N_18813);
and UO_625 (O_625,N_19043,N_18025);
nand UO_626 (O_626,N_19223,N_16642);
nor UO_627 (O_627,N_16420,N_16847);
and UO_628 (O_628,N_19405,N_18628);
nand UO_629 (O_629,N_17296,N_19338);
and UO_630 (O_630,N_17133,N_16142);
nor UO_631 (O_631,N_16126,N_19908);
or UO_632 (O_632,N_16732,N_16793);
nand UO_633 (O_633,N_16643,N_18413);
and UO_634 (O_634,N_17718,N_17615);
nand UO_635 (O_635,N_18997,N_19217);
or UO_636 (O_636,N_17654,N_19101);
nor UO_637 (O_637,N_17994,N_19205);
and UO_638 (O_638,N_18620,N_16686);
and UO_639 (O_639,N_18235,N_19461);
nand UO_640 (O_640,N_17089,N_16257);
nor UO_641 (O_641,N_16072,N_19138);
nand UO_642 (O_642,N_16529,N_16606);
or UO_643 (O_643,N_17808,N_18105);
or UO_644 (O_644,N_18255,N_18726);
nor UO_645 (O_645,N_16376,N_18815);
and UO_646 (O_646,N_16371,N_19802);
nand UO_647 (O_647,N_17496,N_19729);
and UO_648 (O_648,N_16391,N_16234);
xor UO_649 (O_649,N_19852,N_19010);
and UO_650 (O_650,N_17811,N_17314);
nand UO_651 (O_651,N_16578,N_19382);
or UO_652 (O_652,N_16246,N_18707);
nor UO_653 (O_653,N_18473,N_16428);
nand UO_654 (O_654,N_18961,N_19521);
and UO_655 (O_655,N_19569,N_18334);
or UO_656 (O_656,N_17372,N_18365);
nand UO_657 (O_657,N_17854,N_17289);
nor UO_658 (O_658,N_19932,N_16002);
xnor UO_659 (O_659,N_16537,N_18527);
and UO_660 (O_660,N_17861,N_16767);
nor UO_661 (O_661,N_18519,N_18187);
nand UO_662 (O_662,N_16509,N_18524);
nand UO_663 (O_663,N_16673,N_19579);
or UO_664 (O_664,N_17487,N_18969);
and UO_665 (O_665,N_19094,N_17492);
nor UO_666 (O_666,N_18271,N_18652);
nor UO_667 (O_667,N_18373,N_19851);
and UO_668 (O_668,N_17771,N_17322);
nor UO_669 (O_669,N_16344,N_16985);
and UO_670 (O_670,N_19972,N_18208);
and UO_671 (O_671,N_17508,N_16511);
nand UO_672 (O_672,N_16199,N_18302);
nor UO_673 (O_673,N_16671,N_19619);
and UO_674 (O_674,N_17394,N_19029);
nand UO_675 (O_675,N_19977,N_18506);
and UO_676 (O_676,N_17522,N_19085);
or UO_677 (O_677,N_19207,N_18498);
nand UO_678 (O_678,N_16539,N_17073);
nor UO_679 (O_679,N_16890,N_16053);
or UO_680 (O_680,N_19180,N_19628);
or UO_681 (O_681,N_16714,N_18517);
and UO_682 (O_682,N_18307,N_19067);
or UO_683 (O_683,N_17838,N_18646);
nor UO_684 (O_684,N_16331,N_17891);
or UO_685 (O_685,N_17064,N_16284);
nand UO_686 (O_686,N_19674,N_17710);
or UO_687 (O_687,N_16464,N_17437);
or UO_688 (O_688,N_18714,N_17173);
nand UO_689 (O_689,N_17517,N_17998);
nor UO_690 (O_690,N_19302,N_19587);
nand UO_691 (O_691,N_16352,N_17053);
and UO_692 (O_692,N_17631,N_18429);
nand UO_693 (O_693,N_17824,N_16110);
nor UO_694 (O_694,N_19604,N_16462);
nor UO_695 (O_695,N_19175,N_17317);
nor UO_696 (O_696,N_16426,N_18169);
or UO_697 (O_697,N_16029,N_16222);
nor UO_698 (O_698,N_16016,N_19630);
nand UO_699 (O_699,N_16994,N_18265);
nand UO_700 (O_700,N_16003,N_16483);
or UO_701 (O_701,N_18349,N_17822);
nor UO_702 (O_702,N_17924,N_17627);
nand UO_703 (O_703,N_18933,N_18401);
or UO_704 (O_704,N_19996,N_16893);
nand UO_705 (O_705,N_17360,N_17113);
and UO_706 (O_706,N_18455,N_18262);
and UO_707 (O_707,N_17960,N_19170);
and UO_708 (O_708,N_18875,N_16140);
or UO_709 (O_709,N_16378,N_18658);
nand UO_710 (O_710,N_18237,N_16988);
or UO_711 (O_711,N_16295,N_17690);
nor UO_712 (O_712,N_16453,N_19541);
nand UO_713 (O_713,N_16448,N_18129);
or UO_714 (O_714,N_17358,N_17608);
nor UO_715 (O_715,N_17766,N_18418);
and UO_716 (O_716,N_16513,N_16883);
or UO_717 (O_717,N_19987,N_19111);
or UO_718 (O_718,N_18731,N_19275);
nor UO_719 (O_719,N_16790,N_18521);
or UO_720 (O_720,N_18453,N_19452);
and UO_721 (O_721,N_16416,N_16518);
and UO_722 (O_722,N_17333,N_19088);
nor UO_723 (O_723,N_16353,N_18786);
nand UO_724 (O_724,N_18023,N_19677);
nand UO_725 (O_725,N_18830,N_19548);
or UO_726 (O_726,N_19948,N_16042);
or UO_727 (O_727,N_17092,N_17593);
nor UO_728 (O_728,N_18579,N_18395);
nor UO_729 (O_729,N_16965,N_18839);
and UO_730 (O_730,N_19552,N_17659);
or UO_731 (O_731,N_18854,N_16574);
nor UO_732 (O_732,N_18868,N_18629);
or UO_733 (O_733,N_17036,N_16252);
or UO_734 (O_734,N_17339,N_17760);
or UO_735 (O_735,N_16588,N_18670);
and UO_736 (O_736,N_17628,N_19413);
nor UO_737 (O_737,N_18449,N_18744);
nand UO_738 (O_738,N_18324,N_18440);
nand UO_739 (O_739,N_16235,N_18022);
nor UO_740 (O_740,N_16368,N_19659);
and UO_741 (O_741,N_17737,N_18544);
or UO_742 (O_742,N_17816,N_19890);
nor UO_743 (O_743,N_19141,N_19774);
and UO_744 (O_744,N_17351,N_17937);
or UO_745 (O_745,N_19877,N_16933);
or UO_746 (O_746,N_19192,N_18540);
nor UO_747 (O_747,N_19809,N_19547);
nand UO_748 (O_748,N_17735,N_18009);
nand UO_749 (O_749,N_17515,N_16364);
nor UO_750 (O_750,N_19066,N_19615);
nor UO_751 (O_751,N_18588,N_17141);
and UO_752 (O_752,N_16859,N_19866);
nand UO_753 (O_753,N_18141,N_18038);
or UO_754 (O_754,N_19358,N_19035);
nor UO_755 (O_755,N_17454,N_17189);
nor UO_756 (O_756,N_16692,N_18938);
nor UO_757 (O_757,N_19340,N_18820);
nor UO_758 (O_758,N_17513,N_16663);
nor UO_759 (O_759,N_16339,N_17177);
or UO_760 (O_760,N_18836,N_19259);
or UO_761 (O_761,N_17653,N_18149);
nor UO_762 (O_762,N_18771,N_16580);
nand UO_763 (O_763,N_18249,N_17374);
and UO_764 (O_764,N_18161,N_16723);
and UO_765 (O_765,N_19743,N_19440);
nor UO_766 (O_766,N_19883,N_16980);
and UO_767 (O_767,N_17704,N_16435);
xor UO_768 (O_768,N_19797,N_16683);
or UO_769 (O_769,N_17086,N_18647);
nand UO_770 (O_770,N_17652,N_19902);
and UO_771 (O_771,N_17430,N_18312);
or UO_772 (O_772,N_17686,N_18491);
and UO_773 (O_773,N_18370,N_16203);
nand UO_774 (O_774,N_17335,N_17644);
nor UO_775 (O_775,N_18179,N_17184);
or UO_776 (O_776,N_19967,N_17203);
and UO_777 (O_777,N_16289,N_16170);
or UO_778 (O_778,N_19923,N_16564);
or UO_779 (O_779,N_18150,N_19719);
nand UO_780 (O_780,N_16554,N_18623);
and UO_781 (O_781,N_19159,N_18225);
and UO_782 (O_782,N_16620,N_18203);
and UO_783 (O_783,N_18893,N_16107);
nor UO_784 (O_784,N_17054,N_18876);
xor UO_785 (O_785,N_19772,N_16684);
and UO_786 (O_786,N_17279,N_18475);
or UO_787 (O_787,N_17689,N_17785);
xor UO_788 (O_788,N_17984,N_19958);
nand UO_789 (O_789,N_16421,N_17589);
and UO_790 (O_790,N_19693,N_19898);
nand UO_791 (O_791,N_16925,N_17930);
and UO_792 (O_792,N_16305,N_16092);
or UO_793 (O_793,N_18256,N_19227);
and UO_794 (O_794,N_16674,N_16445);
or UO_795 (O_795,N_19151,N_18827);
nand UO_796 (O_796,N_19120,N_18525);
or UO_797 (O_797,N_19234,N_19392);
nor UO_798 (O_798,N_19941,N_19206);
and UO_799 (O_799,N_17461,N_16093);
nand UO_800 (O_800,N_16627,N_19089);
nand UO_801 (O_801,N_16078,N_17996);
nand UO_802 (O_802,N_18257,N_17619);
nand UO_803 (O_803,N_18178,N_19468);
or UO_804 (O_804,N_19311,N_17866);
and UO_805 (O_805,N_17641,N_16188);
nor UO_806 (O_806,N_17039,N_17724);
nor UO_807 (O_807,N_19194,N_17872);
and UO_808 (O_808,N_16433,N_16584);
or UO_809 (O_809,N_17079,N_18035);
nand UO_810 (O_810,N_16171,N_17899);
and UO_811 (O_811,N_16882,N_18612);
nand UO_812 (O_812,N_17103,N_19911);
and UO_813 (O_813,N_16792,N_18303);
nor UO_814 (O_814,N_19591,N_16716);
nor UO_815 (O_815,N_17519,N_18162);
and UO_816 (O_816,N_17625,N_17733);
nand UO_817 (O_817,N_17523,N_18917);
or UO_818 (O_818,N_16877,N_18352);
or UO_819 (O_819,N_18247,N_16330);
nand UO_820 (O_820,N_17427,N_19814);
nor UO_821 (O_821,N_19566,N_18177);
or UO_822 (O_822,N_16976,N_16772);
nor UO_823 (O_823,N_18724,N_17986);
or UO_824 (O_824,N_16211,N_16615);
and UO_825 (O_825,N_18563,N_17383);
and UO_826 (O_826,N_18190,N_16363);
or UO_827 (O_827,N_17963,N_18379);
or UO_828 (O_828,N_19113,N_17297);
nand UO_829 (O_829,N_19978,N_16922);
or UO_830 (O_830,N_19244,N_17664);
and UO_831 (O_831,N_19777,N_18098);
and UO_832 (O_832,N_19970,N_18327);
nand UO_833 (O_833,N_18016,N_17898);
and UO_834 (O_834,N_17747,N_17630);
and UO_835 (O_835,N_18613,N_19600);
nand UO_836 (O_836,N_17243,N_16991);
and UO_837 (O_837,N_19899,N_19209);
or UO_838 (O_838,N_19164,N_18138);
and UO_839 (O_839,N_19261,N_18863);
nor UO_840 (O_840,N_16356,N_19885);
nand UO_841 (O_841,N_19005,N_18091);
and UO_842 (O_842,N_18285,N_16337);
or UO_843 (O_843,N_16243,N_17777);
and UO_844 (O_844,N_17338,N_16028);
or UO_845 (O_845,N_18200,N_17768);
and UO_846 (O_846,N_19404,N_17087);
and UO_847 (O_847,N_18018,N_17032);
nor UO_848 (O_848,N_19655,N_17775);
nor UO_849 (O_849,N_19664,N_19157);
and UO_850 (O_850,N_17205,N_19891);
nand UO_851 (O_851,N_19370,N_18795);
nand UO_852 (O_852,N_19453,N_19858);
nor UO_853 (O_853,N_18709,N_17927);
nor UO_854 (O_854,N_16282,N_17836);
and UO_855 (O_855,N_16278,N_16486);
or UO_856 (O_856,N_17621,N_19511);
and UO_857 (O_857,N_19355,N_16214);
xnor UO_858 (O_858,N_16768,N_18773);
or UO_859 (O_859,N_16784,N_17353);
nor UO_860 (O_860,N_17723,N_19385);
and UO_861 (O_861,N_16758,N_16955);
nand UO_862 (O_862,N_18608,N_17298);
and UO_863 (O_863,N_17876,N_19524);
and UO_864 (O_864,N_17815,N_16971);
nor UO_865 (O_865,N_17102,N_16023);
or UO_866 (O_866,N_17233,N_19616);
and UO_867 (O_867,N_16738,N_18419);
nor UO_868 (O_868,N_17976,N_18040);
and UO_869 (O_869,N_16657,N_17556);
nand UO_870 (O_870,N_16610,N_18354);
nor UO_871 (O_871,N_17107,N_19599);
and UO_872 (O_872,N_17249,N_19882);
nor UO_873 (O_873,N_16843,N_19460);
and UO_874 (O_874,N_17272,N_17873);
nor UO_875 (O_875,N_19785,N_19838);
nand UO_876 (O_876,N_19974,N_17663);
nor UO_877 (O_877,N_17151,N_18561);
nor UO_878 (O_878,N_18619,N_19938);
nor UO_879 (O_879,N_16736,N_19246);
nand UO_880 (O_880,N_17884,N_17692);
nand UO_881 (O_881,N_19835,N_18823);
xor UO_882 (O_882,N_19557,N_17499);
nor UO_883 (O_883,N_16204,N_19559);
or UO_884 (O_884,N_16981,N_16248);
nand UO_885 (O_885,N_18667,N_16081);
nand UO_886 (O_886,N_19515,N_19760);
nor UO_887 (O_887,N_18321,N_16011);
or UO_888 (O_888,N_18210,N_18027);
or UO_889 (O_889,N_17373,N_19049);
or UO_890 (O_890,N_16960,N_19420);
nor UO_891 (O_891,N_17611,N_19749);
nor UO_892 (O_892,N_17480,N_18163);
or UO_893 (O_893,N_19699,N_17756);
nand UO_894 (O_894,N_19756,N_17806);
nand UO_895 (O_895,N_18912,N_19004);
nand UO_896 (O_896,N_16727,N_18057);
and UO_897 (O_897,N_17895,N_19697);
nand UO_898 (O_898,N_17164,N_17266);
nand UO_899 (O_899,N_18093,N_16611);
nor UO_900 (O_900,N_17995,N_19734);
nor UO_901 (O_901,N_18898,N_16533);
and UO_902 (O_902,N_17720,N_16401);
nand UO_903 (O_903,N_19718,N_19663);
nand UO_904 (O_904,N_17159,N_19976);
or UO_905 (O_905,N_19544,N_18377);
nand UO_906 (O_906,N_16006,N_19013);
and UO_907 (O_907,N_17192,N_18638);
nand UO_908 (O_908,N_18562,N_16367);
nand UO_909 (O_909,N_18880,N_18292);
nand UO_910 (O_910,N_17722,N_16519);
and UO_911 (O_911,N_16064,N_19788);
and UO_912 (O_912,N_16419,N_16596);
or UO_913 (O_913,N_18660,N_19895);
nor UO_914 (O_914,N_19419,N_19307);
nor UO_915 (O_915,N_19264,N_17150);
nand UO_916 (O_916,N_18372,N_18300);
nor UO_917 (O_917,N_16493,N_17433);
and UO_918 (O_918,N_19260,N_16989);
nand UO_919 (O_919,N_19943,N_17417);
nor UO_920 (O_920,N_17530,N_16279);
or UO_921 (O_921,N_19288,N_18747);
nand UO_922 (O_922,N_19061,N_17919);
or UO_923 (O_923,N_19353,N_18274);
nor UO_924 (O_924,N_17294,N_17926);
nand UO_925 (O_925,N_18531,N_17000);
xnor UO_926 (O_926,N_17308,N_17100);
nand UO_927 (O_927,N_17354,N_18258);
nor UO_928 (O_928,N_18077,N_18232);
nor UO_929 (O_929,N_18085,N_19062);
or UO_930 (O_930,N_16393,N_17696);
and UO_931 (O_931,N_17423,N_18202);
or UO_932 (O_932,N_16230,N_18864);
nor UO_933 (O_933,N_16208,N_19283);
nand UO_934 (O_934,N_19925,N_16915);
nand UO_935 (O_935,N_16507,N_16293);
and UO_936 (O_936,N_16773,N_16285);
nand UO_937 (O_937,N_17802,N_16658);
nor UO_938 (O_938,N_17068,N_18977);
nor UO_939 (O_939,N_19670,N_16454);
or UO_940 (O_940,N_17045,N_19484);
or UO_941 (O_941,N_18518,N_19277);
nand UO_942 (O_942,N_19248,N_17605);
and UO_943 (O_943,N_18810,N_16869);
nor UO_944 (O_944,N_18143,N_19930);
nor UO_945 (O_945,N_18819,N_16957);
or UO_946 (O_946,N_18573,N_17197);
and UO_947 (O_947,N_19327,N_17590);
nor UO_948 (O_948,N_18549,N_19042);
xor UO_949 (O_949,N_19179,N_16560);
or UO_950 (O_950,N_17269,N_18835);
and UO_951 (O_951,N_16931,N_18672);
nor UO_952 (O_952,N_19078,N_19446);
and UO_953 (O_953,N_16929,N_17488);
nor UO_954 (O_954,N_16498,N_18763);
or UO_955 (O_955,N_19535,N_16392);
or UO_956 (O_956,N_19498,N_18990);
and UO_957 (O_957,N_17326,N_16987);
or UO_958 (O_958,N_17982,N_17250);
nand UO_959 (O_959,N_16436,N_18000);
nor UO_960 (O_960,N_16881,N_19177);
or UO_961 (O_961,N_19188,N_19017);
and UO_962 (O_962,N_17521,N_18002);
nor UO_963 (O_963,N_17788,N_19474);
and UO_964 (O_964,N_17020,N_16527);
and UO_965 (O_965,N_18908,N_17400);
and UO_966 (O_966,N_18856,N_18241);
and UO_967 (O_967,N_18261,N_18778);
nor UO_968 (O_968,N_19383,N_16757);
nand UO_969 (O_969,N_17464,N_19044);
and UO_970 (O_970,N_17136,N_16239);
or UO_971 (O_971,N_16221,N_18586);
nor UO_972 (O_972,N_19825,N_16581);
nand UO_973 (O_973,N_18304,N_16414);
nor UO_974 (O_974,N_17910,N_17550);
nor UO_975 (O_975,N_17878,N_16761);
and UO_976 (O_976,N_16335,N_19494);
or UO_977 (O_977,N_18983,N_17483);
nor UO_978 (O_978,N_18812,N_19466);
nor UO_979 (O_979,N_19403,N_17152);
or UO_980 (O_980,N_16918,N_16083);
nand UO_981 (O_981,N_16473,N_16459);
nor UO_982 (O_982,N_18456,N_17029);
or UO_983 (O_983,N_19464,N_19543);
and UO_984 (O_984,N_18749,N_18643);
nor UO_985 (O_985,N_17916,N_17807);
and UO_986 (O_986,N_16165,N_18788);
nor UO_987 (O_987,N_16542,N_18164);
nor UO_988 (O_988,N_18583,N_17368);
or UO_989 (O_989,N_18125,N_17428);
nand UO_990 (O_990,N_17470,N_16901);
nand UO_991 (O_991,N_17104,N_17436);
nand UO_992 (O_992,N_17617,N_19125);
and UO_993 (O_993,N_19889,N_18597);
nor UO_994 (O_994,N_19735,N_19167);
nor UO_995 (O_995,N_16935,N_17112);
and UO_996 (O_996,N_18630,N_19080);
nand UO_997 (O_997,N_18869,N_19075);
nand UO_998 (O_998,N_17883,N_18501);
and UO_999 (O_999,N_16598,N_18655);
or UO_1000 (O_1000,N_16801,N_18651);
nor UO_1001 (O_1001,N_17938,N_19163);
nand UO_1002 (O_1002,N_18030,N_16408);
and UO_1003 (O_1003,N_16489,N_19361);
nand UO_1004 (O_1004,N_17187,N_19008);
or UO_1005 (O_1005,N_18142,N_17012);
nand UO_1006 (O_1006,N_19298,N_19640);
nor UO_1007 (O_1007,N_19577,N_16399);
nand UO_1008 (O_1008,N_19315,N_16471);
nand UO_1009 (O_1009,N_17201,N_19688);
or UO_1010 (O_1010,N_18266,N_18656);
or UO_1011 (O_1011,N_19456,N_19084);
or UO_1012 (O_1012,N_17584,N_19966);
and UO_1013 (O_1013,N_16515,N_19506);
or UO_1014 (O_1014,N_16780,N_17090);
or UO_1015 (O_1015,N_18806,N_17524);
nor UO_1016 (O_1016,N_18276,N_16541);
and UO_1017 (O_1017,N_17001,N_18704);
nand UO_1018 (O_1018,N_17635,N_19099);
or UO_1019 (O_1019,N_16196,N_19458);
or UO_1020 (O_1020,N_18145,N_19800);
xor UO_1021 (O_1021,N_18387,N_18859);
and UO_1022 (O_1022,N_17705,N_18610);
nor UO_1023 (O_1023,N_16413,N_17051);
nor UO_1024 (O_1024,N_16207,N_17135);
nor UO_1025 (O_1025,N_16799,N_18356);
nand UO_1026 (O_1026,N_16862,N_19874);
nand UO_1027 (O_1027,N_16477,N_19342);
nor UO_1028 (O_1028,N_16820,N_18913);
nand UO_1029 (O_1029,N_18861,N_18132);
and UO_1030 (O_1030,N_19116,N_19454);
nand UO_1031 (O_1031,N_18102,N_18478);
and UO_1032 (O_1032,N_19090,N_17594);
nand UO_1033 (O_1033,N_19475,N_17761);
xnor UO_1034 (O_1034,N_17676,N_17082);
nor UO_1035 (O_1035,N_16558,N_19860);
and UO_1036 (O_1036,N_16688,N_18637);
nand UO_1037 (O_1037,N_19741,N_16187);
and UO_1038 (O_1038,N_17325,N_18542);
nand UO_1039 (O_1039,N_16193,N_19748);
and UO_1040 (O_1040,N_16811,N_17180);
nor UO_1041 (O_1041,N_19546,N_18339);
or UO_1042 (O_1042,N_17324,N_16332);
nor UO_1043 (O_1043,N_19096,N_16460);
nand UO_1044 (O_1044,N_18436,N_16094);
nor UO_1045 (O_1045,N_19136,N_19300);
or UO_1046 (O_1046,N_18618,N_16763);
and UO_1047 (O_1047,N_17028,N_18426);
and UO_1048 (O_1048,N_18587,N_16411);
nor UO_1049 (O_1049,N_19397,N_18851);
and UO_1050 (O_1050,N_17139,N_16205);
and UO_1051 (O_1051,N_17933,N_17573);
nor UO_1052 (O_1052,N_18409,N_18872);
or UO_1053 (O_1053,N_18571,N_19230);
nand UO_1054 (O_1054,N_17478,N_18224);
or UO_1055 (O_1055,N_17063,N_16244);
nand UO_1056 (O_1056,N_17439,N_16864);
nor UO_1057 (O_1057,N_16229,N_18289);
nand UO_1058 (O_1058,N_19757,N_18974);
nand UO_1059 (O_1059,N_19030,N_18363);
and UO_1060 (O_1060,N_17603,N_16508);
and UO_1061 (O_1061,N_18975,N_17406);
and UO_1062 (O_1062,N_17740,N_16735);
and UO_1063 (O_1063,N_17532,N_16482);
nand UO_1064 (O_1064,N_18719,N_18319);
and UO_1065 (O_1065,N_18288,N_17364);
and UO_1066 (O_1066,N_18849,N_16447);
nand UO_1067 (O_1067,N_17336,N_19387);
or UO_1068 (O_1068,N_17988,N_18689);
or UO_1069 (O_1069,N_19406,N_19531);
or UO_1070 (O_1070,N_16947,N_17449);
nor UO_1071 (O_1071,N_17638,N_16750);
nand UO_1072 (O_1072,N_17234,N_18460);
nand UO_1073 (O_1073,N_17070,N_19801);
or UO_1074 (O_1074,N_17056,N_16607);
or UO_1075 (O_1075,N_17379,N_19393);
or UO_1076 (O_1076,N_17950,N_19092);
nor UO_1077 (O_1077,N_16938,N_17494);
nor UO_1078 (O_1078,N_16631,N_19578);
and UO_1079 (O_1079,N_17616,N_18487);
nand UO_1080 (O_1080,N_18697,N_17076);
nor UO_1081 (O_1081,N_18568,N_19893);
or UO_1082 (O_1082,N_16240,N_16141);
or UO_1083 (O_1083,N_16007,N_19095);
nand UO_1084 (O_1084,N_18430,N_18536);
and UO_1085 (O_1085,N_16516,N_19389);
nand UO_1086 (O_1086,N_18746,N_16522);
or UO_1087 (O_1087,N_16937,N_19160);
nand UO_1088 (O_1088,N_19303,N_19583);
or UO_1089 (O_1089,N_17977,N_16468);
nand UO_1090 (O_1090,N_19350,N_16641);
and UO_1091 (O_1091,N_16617,N_16879);
nand UO_1092 (O_1092,N_17485,N_19486);
nor UO_1093 (O_1093,N_16531,N_17890);
or UO_1094 (O_1094,N_17581,N_18888);
and UO_1095 (O_1095,N_17999,N_18420);
or UO_1096 (O_1096,N_16494,N_17993);
or UO_1097 (O_1097,N_17951,N_18668);
nand UO_1098 (O_1098,N_19917,N_19875);
or UO_1099 (O_1099,N_18152,N_16496);
nand UO_1100 (O_1100,N_16913,N_17215);
or UO_1101 (O_1101,N_19820,N_16427);
xor UO_1102 (O_1102,N_16328,N_19220);
nand UO_1103 (O_1103,N_17947,N_18069);
nand UO_1104 (O_1104,N_19257,N_17235);
and UO_1105 (O_1105,N_16342,N_18774);
and UO_1106 (O_1106,N_18173,N_19024);
nand UO_1107 (O_1107,N_17311,N_18244);
and UO_1108 (O_1108,N_18305,N_19359);
or UO_1109 (O_1109,N_18198,N_16063);
nor UO_1110 (O_1110,N_16936,N_19491);
or UO_1111 (O_1111,N_16220,N_17240);
nor UO_1112 (O_1112,N_17734,N_19238);
nand UO_1113 (O_1113,N_16850,N_17281);
nor UO_1114 (O_1114,N_17387,N_18547);
and UO_1115 (O_1115,N_16569,N_17055);
nand UO_1116 (O_1116,N_16614,N_19585);
nand UO_1117 (O_1117,N_18346,N_18246);
and UO_1118 (O_1118,N_16572,N_18463);
nor UO_1119 (O_1119,N_18497,N_17422);
or UO_1120 (O_1120,N_17991,N_16646);
or UO_1121 (O_1121,N_19588,N_16434);
or UO_1122 (O_1122,N_18019,N_16595);
and UO_1123 (O_1123,N_17486,N_19441);
nand UO_1124 (O_1124,N_17310,N_17170);
nand UO_1125 (O_1125,N_19492,N_19236);
nor UO_1126 (O_1126,N_16010,N_19648);
nor UO_1127 (O_1127,N_19679,N_17671);
and UO_1128 (O_1128,N_18700,N_19376);
nor UO_1129 (O_1129,N_16169,N_16734);
or UO_1130 (O_1130,N_17719,N_16651);
nand UO_1131 (O_1131,N_19287,N_17075);
and UO_1132 (O_1132,N_17033,N_16191);
or UO_1133 (O_1133,N_16848,N_17858);
nand UO_1134 (O_1134,N_16055,N_17896);
nand UO_1135 (O_1135,N_16556,N_18029);
nand UO_1136 (O_1136,N_18270,N_18775);
or UO_1137 (O_1137,N_16639,N_17459);
or UO_1138 (O_1138,N_16424,N_18734);
and UO_1139 (O_1139,N_16373,N_16815);
nand UO_1140 (O_1140,N_17261,N_17094);
and UO_1141 (O_1141,N_18278,N_16415);
or UO_1142 (O_1142,N_19091,N_19324);
and UO_1143 (O_1143,N_17010,N_18423);
and UO_1144 (O_1144,N_17925,N_19633);
nor UO_1145 (O_1145,N_18042,N_16456);
nor UO_1146 (O_1146,N_18298,N_17213);
or UO_1147 (O_1147,N_19892,N_19255);
nor UO_1148 (O_1148,N_16004,N_17828);
nand UO_1149 (O_1149,N_17009,N_18828);
and UO_1150 (O_1150,N_18779,N_18783);
and UO_1151 (O_1151,N_17490,N_18459);
nor UO_1152 (O_1152,N_16899,N_17062);
nand UO_1153 (O_1153,N_19251,N_19308);
or UO_1154 (O_1154,N_18397,N_17697);
nor UO_1155 (O_1155,N_18469,N_17131);
or UO_1156 (O_1156,N_19817,N_17140);
nor UO_1157 (O_1157,N_18922,N_16535);
nor UO_1158 (O_1158,N_16422,N_16604);
and UO_1159 (O_1159,N_16999,N_18865);
nand UO_1160 (O_1160,N_18941,N_18852);
nand UO_1161 (O_1161,N_19618,N_19501);
and UO_1162 (O_1162,N_19716,N_19040);
nand UO_1163 (O_1163,N_19573,N_19522);
nand UO_1164 (O_1164,N_17069,N_17134);
nand UO_1165 (O_1165,N_17493,N_16719);
and UO_1166 (O_1166,N_18394,N_19709);
or UO_1167 (O_1167,N_17979,N_19607);
and UO_1168 (O_1168,N_18837,N_18822);
nor UO_1169 (O_1169,N_16228,N_18368);
nand UO_1170 (O_1170,N_19081,N_19444);
xnor UO_1171 (O_1171,N_19747,N_18245);
nand UO_1172 (O_1172,N_19009,N_17186);
nand UO_1173 (O_1173,N_16075,N_18514);
nand UO_1174 (O_1174,N_18095,N_19184);
or UO_1175 (O_1175,N_19819,N_18768);
and UO_1176 (O_1176,N_16300,N_19038);
xnor UO_1177 (O_1177,N_16590,N_17081);
nor UO_1178 (O_1178,N_19253,N_19053);
and UO_1179 (O_1179,N_16019,N_17471);
nand UO_1180 (O_1180,N_16095,N_16260);
or UO_1181 (O_1181,N_18742,N_18602);
or UO_1182 (O_1182,N_18117,N_17315);
nand UO_1183 (O_1183,N_19348,N_17543);
nand UO_1184 (O_1184,N_19979,N_16283);
or UO_1185 (O_1185,N_19310,N_18351);
nor UO_1186 (O_1186,N_16117,N_18743);
nor UO_1187 (O_1187,N_19897,N_18020);
nand UO_1188 (O_1188,N_17797,N_17414);
nand UO_1189 (O_1189,N_17849,N_19416);
or UO_1190 (O_1190,N_19761,N_18622);
and UO_1191 (O_1191,N_19685,N_16253);
nor UO_1192 (O_1192,N_17396,N_16833);
or UO_1193 (O_1193,N_19832,N_17859);
or UO_1194 (O_1194,N_16037,N_17964);
nor UO_1195 (O_1195,N_17856,N_17119);
or UO_1196 (O_1196,N_18287,N_18962);
nand UO_1197 (O_1197,N_17553,N_18034);
or UO_1198 (O_1198,N_17328,N_16262);
or UO_1199 (O_1199,N_19276,N_18236);
nor UO_1200 (O_1200,N_18767,N_16292);
nor UO_1201 (O_1201,N_18566,N_19865);
nand UO_1202 (O_1202,N_16932,N_18920);
or UO_1203 (O_1203,N_18873,N_19525);
nor UO_1204 (O_1204,N_17277,N_18482);
or UO_1205 (O_1205,N_16629,N_16721);
and UO_1206 (O_1206,N_18026,N_19724);
nand UO_1207 (O_1207,N_19680,N_16652);
or UO_1208 (O_1208,N_17780,N_18052);
or UO_1209 (O_1209,N_17640,N_19268);
xnor UO_1210 (O_1210,N_16490,N_16731);
and UO_1211 (O_1211,N_19758,N_16218);
or UO_1212 (O_1212,N_17840,N_19962);
or UO_1213 (O_1213,N_16308,N_18609);
and UO_1214 (O_1214,N_16388,N_19258);
or UO_1215 (O_1215,N_19592,N_18980);
nand UO_1216 (O_1216,N_19787,N_17691);
or UO_1217 (O_1217,N_19476,N_18065);
and UO_1218 (O_1218,N_18987,N_17932);
nand UO_1219 (O_1219,N_16551,N_18970);
and UO_1220 (O_1220,N_17942,N_18550);
nor UO_1221 (O_1221,N_17656,N_18189);
nor UO_1222 (O_1222,N_18584,N_16565);
or UO_1223 (O_1223,N_19766,N_17750);
nor UO_1224 (O_1224,N_19706,N_17248);
nand UO_1225 (O_1225,N_18380,N_19620);
or UO_1226 (O_1226,N_18165,N_16737);
and UO_1227 (O_1227,N_16310,N_19182);
or UO_1228 (O_1228,N_18935,N_19714);
nor UO_1229 (O_1229,N_17943,N_19989);
nor UO_1230 (O_1230,N_18664,N_18570);
nor UO_1231 (O_1231,N_17040,N_18594);
nor UO_1232 (O_1232,N_18219,N_17048);
and UO_1233 (O_1233,N_18877,N_19108);
nand UO_1234 (O_1234,N_18075,N_16676);
nor UO_1235 (O_1235,N_19128,N_19193);
nand UO_1236 (O_1236,N_16014,N_18606);
or UO_1237 (O_1237,N_16703,N_17392);
and UO_1238 (O_1238,N_18733,N_17624);
and UO_1239 (O_1239,N_17694,N_16861);
and UO_1240 (O_1240,N_16687,N_18318);
or UO_1241 (O_1241,N_17247,N_19723);
and UO_1242 (O_1242,N_16258,N_16058);
or UO_1243 (O_1243,N_19610,N_19935);
nor UO_1244 (O_1244,N_17043,N_19682);
nor UO_1245 (O_1245,N_19804,N_16475);
and UO_1246 (O_1246,N_18721,N_16609);
and UO_1247 (O_1247,N_16567,N_18654);
or UO_1248 (O_1248,N_19745,N_17614);
nand UO_1249 (O_1249,N_19280,N_16956);
or UO_1250 (O_1250,N_16810,N_18120);
and UO_1251 (O_1251,N_18666,N_19927);
nand UO_1252 (O_1252,N_17474,N_18116);
nor UO_1253 (O_1253,N_19115,N_19097);
and UO_1254 (O_1254,N_17601,N_19485);
and UO_1255 (O_1255,N_17580,N_17061);
or UO_1256 (O_1256,N_18053,N_16766);
and UO_1257 (O_1257,N_18414,N_19982);
or UO_1258 (O_1258,N_17708,N_19847);
and UO_1259 (O_1259,N_19780,N_17204);
nand UO_1260 (O_1260,N_18500,N_17839);
nor UO_1261 (O_1261,N_19019,N_16868);
nor UO_1262 (O_1262,N_16001,N_19937);
and UO_1263 (O_1263,N_17609,N_16983);
nor UO_1264 (O_1264,N_16709,N_17382);
nor UO_1265 (O_1265,N_17588,N_16418);
nor UO_1266 (O_1266,N_17230,N_19011);
nor UO_1267 (O_1267,N_16354,N_17973);
nand UO_1268 (O_1268,N_16855,N_18805);
and UO_1269 (O_1269,N_18556,N_19313);
nand UO_1270 (O_1270,N_18461,N_19325);
nand UO_1271 (O_1271,N_18388,N_18090);
nor UO_1272 (O_1272,N_18168,N_17782);
or UO_1273 (O_1273,N_18024,N_19129);
nand UO_1274 (O_1274,N_19580,N_16561);
or UO_1275 (O_1275,N_16044,N_19538);
nand UO_1276 (O_1276,N_19765,N_19762);
nand UO_1277 (O_1277,N_17813,N_19955);
nor UO_1278 (O_1278,N_18201,N_16858);
and UO_1279 (O_1279,N_16880,N_19022);
nor UO_1280 (O_1280,N_18998,N_19332);
nor UO_1281 (O_1281,N_17763,N_17122);
or UO_1282 (O_1282,N_19912,N_18010);
or UO_1283 (O_1283,N_18659,N_19190);
or UO_1284 (O_1284,N_17542,N_18981);
nor UO_1285 (O_1285,N_16036,N_17679);
nor UO_1286 (O_1286,N_16497,N_18528);
nor UO_1287 (O_1287,N_16638,N_18205);
nor UO_1288 (O_1288,N_16908,N_19710);
and UO_1289 (O_1289,N_19069,N_17231);
nand UO_1290 (O_1290,N_18071,N_19590);
and UO_1291 (O_1291,N_16930,N_19558);
or UO_1292 (O_1292,N_19968,N_17346);
xnor UO_1293 (O_1293,N_18171,N_17819);
or UO_1294 (O_1294,N_19291,N_17355);
and UO_1295 (O_1295,N_19921,N_18809);
and UO_1296 (O_1296,N_17327,N_18432);
or UO_1297 (O_1297,N_16151,N_19065);
nor UO_1298 (O_1298,N_18555,N_19478);
and UO_1299 (O_1299,N_16275,N_19810);
nor UO_1300 (O_1300,N_18947,N_18537);
nand UO_1301 (O_1301,N_17409,N_17367);
or UO_1302 (O_1302,N_19296,N_17194);
nor UO_1303 (O_1303,N_16717,N_18522);
or UO_1304 (O_1304,N_19507,N_16762);
nand UO_1305 (O_1305,N_16786,N_17302);
nor UO_1306 (O_1306,N_17084,N_19660);
and UO_1307 (O_1307,N_17411,N_19657);
and UO_1308 (O_1308,N_16090,N_19773);
or UO_1309 (O_1309,N_16323,N_17732);
or UO_1310 (O_1310,N_18175,N_16863);
nand UO_1311 (O_1311,N_18011,N_18080);
and UO_1312 (O_1312,N_17865,N_19560);
nand UO_1313 (O_1313,N_16189,N_16360);
or UO_1314 (O_1314,N_17738,N_18192);
or UO_1315 (O_1315,N_18039,N_19612);
or UO_1316 (O_1316,N_18772,N_19449);
or UO_1317 (O_1317,N_16124,N_18605);
and UO_1318 (O_1318,N_18900,N_19364);
or UO_1319 (O_1319,N_16202,N_19647);
nand UO_1320 (O_1320,N_17662,N_18738);
and UO_1321 (O_1321,N_17218,N_17565);
nor UO_1322 (O_1322,N_16227,N_17018);
or UO_1323 (O_1323,N_16385,N_16984);
nor UO_1324 (O_1324,N_19644,N_18671);
or UO_1325 (O_1325,N_17165,N_19384);
or UO_1326 (O_1326,N_18569,N_17600);
and UO_1327 (O_1327,N_19676,N_17862);
nor UO_1328 (O_1328,N_19225,N_16366);
and UO_1329 (O_1329,N_18711,N_18907);
and UO_1330 (O_1330,N_19285,N_19555);
nor UO_1331 (O_1331,N_16226,N_18825);
nor UO_1332 (O_1332,N_16481,N_16247);
or UO_1333 (O_1333,N_18740,N_16425);
or UO_1334 (O_1334,N_18759,N_18367);
nor UO_1335 (O_1335,N_19973,N_17199);
nand UO_1336 (O_1336,N_19161,N_18156);
and UO_1337 (O_1337,N_18924,N_19508);
or UO_1338 (O_1338,N_17745,N_17683);
and UO_1339 (O_1339,N_16885,N_19622);
or UO_1340 (O_1340,N_18565,N_18092);
nand UO_1341 (O_1341,N_19830,N_19158);
nand UO_1342 (O_1342,N_18635,N_17709);
or UO_1343 (O_1343,N_17863,N_19386);
nand UO_1344 (O_1344,N_18971,N_16338);
or UO_1345 (O_1345,N_17911,N_17825);
or UO_1346 (O_1346,N_17798,N_19643);
and UO_1347 (O_1347,N_18188,N_18829);
and UO_1348 (O_1348,N_18295,N_19121);
or UO_1349 (O_1349,N_18048,N_16223);
nor UO_1350 (O_1350,N_19304,N_17077);
and UO_1351 (O_1351,N_18393,N_17769);
and UO_1352 (O_1352,N_17244,N_19654);
nor UO_1353 (O_1353,N_19713,N_18607);
nor UO_1354 (O_1354,N_16397,N_16958);
nor UO_1355 (O_1355,N_19708,N_17223);
or UO_1356 (O_1356,N_19470,N_19284);
nor UO_1357 (O_1357,N_16201,N_18526);
or UO_1358 (O_1358,N_17067,N_16914);
nand UO_1359 (O_1359,N_16054,N_17955);
nand UO_1360 (O_1360,N_19964,N_17672);
or UO_1361 (O_1361,N_18421,N_17803);
or UO_1362 (O_1362,N_17881,N_19613);
nor UO_1363 (O_1363,N_19301,N_18532);
nor UO_1364 (O_1364,N_19642,N_19503);
and UO_1365 (O_1365,N_16441,N_17789);
or UO_1366 (O_1366,N_18458,N_16150);
or UO_1367 (O_1367,N_18403,N_17185);
or UO_1368 (O_1368,N_17349,N_18183);
nand UO_1369 (O_1369,N_17352,N_16101);
and UO_1370 (O_1370,N_19595,N_19222);
nand UO_1371 (O_1371,N_17035,N_16940);
and UO_1372 (O_1372,N_16532,N_19853);
nand UO_1373 (O_1373,N_19901,N_16000);
and UO_1374 (O_1374,N_18992,N_18260);
nor UO_1375 (O_1375,N_16696,N_18675);
or UO_1376 (O_1376,N_18045,N_17512);
or UO_1377 (O_1377,N_17674,N_16022);
nand UO_1378 (O_1378,N_18634,N_19886);
nor UO_1379 (O_1379,N_16104,N_18043);
nand UO_1380 (O_1380,N_16175,N_16852);
nor UO_1381 (O_1381,N_19540,N_19150);
or UO_1382 (O_1382,N_19596,N_16467);
nand UO_1383 (O_1383,N_19678,N_16503);
and UO_1384 (O_1384,N_16361,N_19438);
or UO_1385 (O_1385,N_19776,N_17742);
or UO_1386 (O_1386,N_17583,N_18730);
and UO_1387 (O_1387,N_19063,N_16452);
nor UO_1388 (O_1388,N_16662,N_18355);
or UO_1389 (O_1389,N_18585,N_19687);
or UO_1390 (O_1390,N_19130,N_17757);
nor UO_1391 (O_1391,N_18509,N_16047);
or UO_1392 (O_1392,N_18005,N_19243);
and UO_1393 (O_1393,N_17551,N_17504);
and UO_1394 (O_1394,N_17673,N_18600);
or UO_1395 (O_1395,N_18874,N_17698);
or UO_1396 (O_1396,N_19712,N_19437);
or UO_1397 (O_1397,N_17569,N_18424);
nand UO_1398 (O_1398,N_19526,N_16430);
nor UO_1399 (O_1399,N_18906,N_19467);
or UO_1400 (O_1400,N_16438,N_18713);
nand UO_1401 (O_1401,N_18431,N_18766);
nor UO_1402 (O_1402,N_18979,N_19271);
nand UO_1403 (O_1403,N_19939,N_16912);
nand UO_1404 (O_1404,N_19278,N_18047);
or UO_1405 (O_1405,N_18895,N_17260);
or UO_1406 (O_1406,N_17518,N_17871);
or UO_1407 (O_1407,N_17402,N_17220);
nor UO_1408 (O_1408,N_17011,N_17160);
and UO_1409 (O_1409,N_16830,N_19999);
nor UO_1410 (O_1410,N_16173,N_18066);
or UO_1411 (O_1411,N_16265,N_17126);
nor UO_1412 (O_1412,N_16583,N_16728);
or UO_1413 (O_1413,N_19636,N_19457);
nor UO_1414 (O_1414,N_18811,N_16544);
nand UO_1415 (O_1415,N_17301,N_16618);
nand UO_1416 (O_1416,N_16829,N_18741);
and UO_1417 (O_1417,N_16297,N_16035);
nand UO_1418 (O_1418,N_17642,N_17903);
and UO_1419 (O_1419,N_16579,N_19556);
nand UO_1420 (O_1420,N_17764,N_17677);
nand UO_1421 (O_1421,N_16288,N_19326);
or UO_1422 (O_1422,N_19368,N_16530);
and UO_1423 (O_1423,N_18603,N_17570);
or UO_1424 (O_1424,N_16067,N_19805);
nor UO_1425 (O_1425,N_19279,N_18708);
or UO_1426 (O_1426,N_18408,N_17844);
or UO_1427 (O_1427,N_18239,N_17495);
nand UO_1428 (O_1428,N_16136,N_17095);
nand UO_1429 (O_1429,N_19213,N_18625);
and UO_1430 (O_1430,N_18753,N_18253);
nor UO_1431 (O_1431,N_16794,N_16902);
or UO_1432 (O_1432,N_17731,N_18847);
and UO_1433 (O_1433,N_18466,N_19617);
nand UO_1434 (O_1434,N_18950,N_17680);
or UO_1435 (O_1435,N_18886,N_16474);
or UO_1436 (O_1436,N_18745,N_19409);
or UO_1437 (O_1437,N_19606,N_17632);
or UO_1438 (O_1438,N_19381,N_19077);
nand UO_1439 (O_1439,N_16130,N_18006);
nand UO_1440 (O_1440,N_16675,N_19333);
nor UO_1441 (O_1441,N_19126,N_16634);
and UO_1442 (O_1442,N_16287,N_17948);
nor UO_1443 (O_1443,N_17232,N_19481);
nand UO_1444 (O_1444,N_16350,N_17528);
or UO_1445 (O_1445,N_16540,N_16751);
or UO_1446 (O_1446,N_19867,N_16431);
or UO_1447 (O_1447,N_16505,N_16069);
or UO_1448 (O_1448,N_17721,N_19528);
nand UO_1449 (O_1449,N_17909,N_19915);
nand UO_1450 (O_1450,N_18348,N_18407);
nor UO_1451 (O_1451,N_16329,N_18930);
and UO_1452 (O_1452,N_17120,N_16916);
nor UO_1453 (O_1453,N_18665,N_17124);
or UO_1454 (O_1454,N_19837,N_17746);
nor UO_1455 (O_1455,N_16046,N_17699);
and UO_1456 (O_1456,N_18094,N_19186);
or UO_1457 (O_1457,N_16224,N_18337);
and UO_1458 (O_1458,N_19367,N_16690);
and UO_1459 (O_1459,N_19916,N_17271);
or UO_1460 (O_1460,N_18944,N_18103);
nand UO_1461 (O_1461,N_18843,N_19046);
or UO_1462 (O_1462,N_16123,N_19623);
nor UO_1463 (O_1463,N_16853,N_16139);
and UO_1464 (O_1464,N_18816,N_16147);
and UO_1465 (O_1465,N_16546,N_18777);
xor UO_1466 (O_1466,N_17257,N_17531);
nor UO_1467 (O_1467,N_17965,N_19490);
and UO_1468 (O_1468,N_19208,N_18764);
nor UO_1469 (O_1469,N_16707,N_19434);
nor UO_1470 (O_1470,N_17545,N_17633);
nand UO_1471 (O_1471,N_19037,N_18112);
nor UO_1472 (O_1472,N_17431,N_17016);
xor UO_1473 (O_1473,N_19725,N_16670);
and UO_1474 (O_1474,N_19196,N_16217);
nor UO_1475 (O_1475,N_18415,N_18889);
or UO_1476 (O_1476,N_16309,N_16857);
nand UO_1477 (O_1477,N_16837,N_18867);
and UO_1478 (O_1478,N_18341,N_18109);
nor UO_1479 (O_1479,N_17435,N_18504);
or UO_1480 (O_1480,N_16180,N_19414);
nor UO_1481 (O_1481,N_17970,N_19148);
nor UO_1482 (O_1482,N_19424,N_19740);
nand UO_1483 (O_1483,N_17855,N_18956);
nand UO_1484 (O_1484,N_19651,N_16962);
nand UO_1485 (O_1485,N_19362,N_17666);
or UO_1486 (O_1486,N_19873,N_18153);
nand UO_1487 (O_1487,N_17983,N_17562);
or UO_1488 (O_1488,N_17227,N_18492);
and UO_1489 (O_1489,N_19969,N_16304);
or UO_1490 (O_1490,N_16276,N_19154);
and UO_1491 (O_1491,N_18755,N_16741);
nand UO_1492 (O_1492,N_19093,N_16138);
nand UO_1493 (O_1493,N_17366,N_19913);
nor UO_1494 (O_1494,N_17906,N_18126);
and UO_1495 (O_1495,N_17344,N_17928);
nand UO_1496 (O_1496,N_18706,N_17017);
nand UO_1497 (O_1497,N_18883,N_18441);
nand UO_1498 (O_1498,N_17306,N_18343);
nor UO_1499 (O_1499,N_19472,N_17845);
nor UO_1500 (O_1500,N_18382,N_17290);
or UO_1501 (O_1501,N_16510,N_17500);
or UO_1502 (O_1502,N_16633,N_19394);
nand UO_1503 (O_1503,N_19609,N_16600);
or UO_1504 (O_1504,N_18967,N_17560);
nor UO_1505 (O_1505,N_16442,N_16298);
and UO_1506 (O_1506,N_17520,N_18041);
nand UO_1507 (O_1507,N_19098,N_19683);
nor UO_1508 (O_1508,N_16679,N_18640);
nor UO_1509 (O_1509,N_17429,N_17940);
or UO_1510 (O_1510,N_17407,N_16488);
or UO_1511 (O_1511,N_19625,N_18785);
or UO_1512 (O_1512,N_17228,N_19791);
or UO_1513 (O_1513,N_16632,N_19400);
and UO_1514 (O_1514,N_16192,N_16317);
or UO_1515 (O_1515,N_16194,N_17870);
or UO_1516 (O_1516,N_18988,N_16405);
or UO_1517 (O_1517,N_18649,N_18310);
nor UO_1518 (O_1518,N_19823,N_16845);
nor UO_1519 (O_1519,N_19064,N_18181);
nor UO_1520 (O_1520,N_17509,N_16680);
nor UO_1521 (O_1521,N_18853,N_18728);
or UO_1522 (O_1522,N_16654,N_18233);
or UO_1523 (O_1523,N_18417,N_18505);
nand UO_1524 (O_1524,N_19570,N_16694);
and UO_1525 (O_1525,N_16873,N_18952);
and UO_1526 (O_1526,N_19191,N_16796);
and UO_1527 (O_1527,N_16921,N_17285);
and UO_1528 (O_1528,N_18329,N_18240);
nand UO_1529 (O_1529,N_18838,N_17675);
nand UO_1530 (O_1530,N_18467,N_16653);
nand UO_1531 (O_1531,N_18858,N_18433);
and UO_1532 (O_1532,N_18831,N_17108);
or UO_1533 (O_1533,N_18678,N_18871);
or UO_1534 (O_1534,N_19988,N_19366);
nand UO_1535 (O_1535,N_18082,N_17484);
nand UO_1536 (O_1536,N_19272,N_16982);
nor UO_1537 (O_1537,N_17715,N_18800);
nor UO_1538 (O_1538,N_18642,N_16432);
and UO_1539 (O_1539,N_19329,N_16693);
and UO_1540 (O_1540,N_17169,N_17410);
nor UO_1541 (O_1541,N_19450,N_17826);
nor UO_1542 (O_1542,N_17137,N_19074);
nand UO_1543 (O_1543,N_16128,N_17875);
and UO_1544 (O_1544,N_18110,N_16655);
nand UO_1545 (O_1545,N_18137,N_19815);
and UO_1546 (O_1546,N_19872,N_19790);
xnor UO_1547 (O_1547,N_18953,N_19681);
or UO_1548 (O_1548,N_18452,N_17537);
nand UO_1549 (O_1549,N_16586,N_16463);
nand UO_1550 (O_1550,N_17823,N_19857);
nor UO_1551 (O_1551,N_18995,N_17268);
and UO_1552 (O_1552,N_18404,N_17157);
or UO_1553 (O_1553,N_16256,N_16941);
nor UO_1554 (O_1554,N_19363,N_17027);
and UO_1555 (O_1555,N_16986,N_19690);
nand UO_1556 (O_1556,N_17448,N_17072);
nor UO_1557 (O_1557,N_18611,N_18648);
nor UO_1558 (O_1558,N_17080,N_19189);
nor UO_1559 (O_1559,N_19635,N_18508);
nor UO_1560 (O_1560,N_16822,N_19127);
nor UO_1561 (O_1561,N_17578,N_18691);
or UO_1562 (O_1562,N_19631,N_16691);
or UO_1563 (O_1563,N_16623,N_19739);
nor UO_1564 (O_1564,N_18705,N_16592);
and UO_1565 (O_1565,N_19940,N_19162);
or UO_1566 (O_1566,N_16712,N_18581);
nor UO_1567 (O_1567,N_19002,N_18400);
and UO_1568 (O_1568,N_19124,N_19317);
nand UO_1569 (O_1569,N_16968,N_17707);
and UO_1570 (O_1570,N_17606,N_19429);
and UO_1571 (O_1571,N_17003,N_17682);
or UO_1572 (O_1572,N_19744,N_18113);
or UO_1573 (O_1573,N_17832,N_19051);
or UO_1574 (O_1574,N_18963,N_19598);
and UO_1575 (O_1575,N_16135,N_19821);
and UO_1576 (O_1576,N_17386,N_16919);
and UO_1577 (O_1577,N_17639,N_19379);
or UO_1578 (O_1578,N_17557,N_18306);
or UO_1579 (O_1579,N_17776,N_16538);
or UO_1580 (O_1580,N_16179,N_17356);
or UO_1581 (O_1581,N_17145,N_16074);
nand UO_1582 (O_1582,N_19554,N_16443);
or UO_1583 (O_1583,N_17962,N_19032);
nand UO_1584 (O_1584,N_19764,N_19003);
nor UO_1585 (O_1585,N_17800,N_17183);
and UO_1586 (O_1586,N_16210,N_16824);
nand UO_1587 (O_1587,N_19667,N_17511);
nor UO_1588 (O_1588,N_19997,N_16710);
nor UO_1589 (O_1589,N_19047,N_16026);
and UO_1590 (O_1590,N_17544,N_17529);
nand UO_1591 (O_1591,N_17332,N_16480);
or UO_1592 (O_1592,N_18727,N_18396);
and UO_1593 (O_1593,N_17006,N_18028);
nor UO_1594 (O_1594,N_16325,N_17921);
or UO_1595 (O_1595,N_16272,N_16745);
nor UO_1596 (O_1596,N_16027,N_19250);
nor UO_1597 (O_1597,N_18471,N_18196);
nand UO_1598 (O_1598,N_19107,N_18158);
or UO_1599 (O_1599,N_18333,N_16174);
and UO_1600 (O_1600,N_18958,N_18064);
nand UO_1601 (O_1601,N_19789,N_18068);
nand UO_1602 (O_1602,N_16724,N_18291);
nand UO_1603 (O_1603,N_16889,N_18242);
nor UO_1604 (O_1604,N_16061,N_18371);
and UO_1605 (O_1605,N_17778,N_17549);
nand UO_1606 (O_1606,N_19408,N_17251);
or UO_1607 (O_1607,N_18903,N_16121);
or UO_1608 (O_1608,N_16085,N_17109);
or UO_1609 (O_1609,N_18539,N_19267);
or UO_1610 (O_1610,N_16213,N_19775);
or UO_1611 (O_1611,N_16197,N_16963);
nand UO_1612 (O_1612,N_16842,N_18890);
nand UO_1613 (O_1613,N_17842,N_16978);
or UO_1614 (O_1614,N_19025,N_17214);
nand UO_1615 (O_1615,N_17527,N_16231);
nor UO_1616 (O_1616,N_16926,N_17462);
and UO_1617 (O_1617,N_18199,N_17702);
nor UO_1618 (O_1618,N_18545,N_18008);
nand UO_1619 (O_1619,N_16523,N_19903);
nand UO_1620 (O_1620,N_17539,N_16440);
nand UO_1621 (O_1621,N_18128,N_18059);
or UO_1622 (O_1622,N_17981,N_18496);
or UO_1623 (O_1623,N_18617,N_19845);
nand UO_1624 (O_1624,N_19947,N_19166);
nand UO_1625 (O_1625,N_18412,N_17191);
nand UO_1626 (O_1626,N_18616,N_19742);
nor UO_1627 (O_1627,N_17885,N_18703);
or UO_1628 (O_1628,N_17401,N_18448);
nand UO_1629 (O_1629,N_16993,N_18892);
nor UO_1630 (O_1630,N_17222,N_18791);
and UO_1631 (O_1631,N_18927,N_17273);
or UO_1632 (O_1632,N_17008,N_18268);
nor UO_1633 (O_1633,N_17369,N_16748);
nand UO_1634 (O_1634,N_17502,N_18748);
xor UO_1635 (O_1635,N_16619,N_19228);
nand UO_1636 (O_1636,N_18350,N_19021);
nor UO_1637 (O_1637,N_16209,N_17323);
and UO_1638 (O_1638,N_17869,N_17182);
nand UO_1639 (O_1639,N_17954,N_18932);
or UO_1640 (O_1640,N_19803,N_17284);
or UO_1641 (O_1641,N_18087,N_17455);
or UO_1642 (O_1642,N_16303,N_17334);
nor UO_1643 (O_1643,N_17505,N_19841);
nor UO_1644 (O_1644,N_19698,N_17585);
nor UO_1645 (O_1645,N_16917,N_17278);
nor UO_1646 (O_1646,N_18754,N_16718);
or UO_1647 (O_1647,N_18332,N_17665);
or UO_1648 (O_1648,N_17489,N_19007);
or UO_1649 (O_1649,N_19274,N_17283);
and UO_1650 (O_1650,N_18996,N_18301);
nor UO_1651 (O_1651,N_19433,N_16313);
nand UO_1652 (O_1652,N_18984,N_16479);
nor UO_1653 (O_1653,N_19292,N_16924);
and UO_1654 (O_1654,N_19465,N_19226);
nor UO_1655 (O_1655,N_19671,N_18325);
or UO_1656 (O_1656,N_18799,N_18474);
nand UO_1657 (O_1657,N_16648,N_19602);
and UO_1658 (O_1658,N_19133,N_16500);
nor UO_1659 (O_1659,N_18833,N_17586);
nor UO_1660 (O_1660,N_19513,N_18056);
nand UO_1661 (O_1661,N_17146,N_17567);
or UO_1662 (O_1662,N_16977,N_19836);
or UO_1663 (O_1663,N_17510,N_18782);
and UO_1664 (O_1664,N_17320,N_17190);
nand UO_1665 (O_1665,N_16664,N_16759);
and UO_1666 (O_1666,N_18826,N_18615);
or UO_1667 (O_1667,N_17661,N_19057);
and UO_1668 (O_1668,N_19641,N_18494);
nor UO_1669 (O_1669,N_16711,N_17939);
nand UO_1670 (O_1670,N_19984,N_17200);
nand UO_1671 (O_1671,N_17477,N_18925);
and UO_1672 (O_1672,N_16599,N_16568);
nor UO_1673 (O_1673,N_18154,N_19135);
nor UO_1674 (O_1674,N_19634,N_17548);
nor UO_1675 (O_1675,N_16132,N_18411);
and UO_1676 (O_1676,N_19502,N_17026);
nand UO_1677 (O_1677,N_16802,N_17908);
nor UO_1678 (O_1678,N_16160,N_16485);
nor UO_1679 (O_1679,N_19653,N_19221);
or UO_1680 (O_1680,N_17915,N_16585);
and UO_1681 (O_1681,N_19399,N_17128);
nand UO_1682 (O_1682,N_18818,N_16382);
and UO_1683 (O_1683,N_16644,N_16836);
nand UO_1684 (O_1684,N_18481,N_16722);
nor UO_1685 (O_1685,N_16923,N_18794);
and UO_1686 (O_1686,N_19155,N_17217);
nand UO_1687 (O_1687,N_19539,N_16874);
nor UO_1688 (O_1688,N_16504,N_18277);
or UO_1689 (O_1689,N_16927,N_19395);
nand UO_1690 (O_1690,N_18101,N_16215);
nor UO_1691 (O_1691,N_18862,N_18535);
nand UO_1692 (O_1692,N_16185,N_17309);
nand UO_1693 (O_1693,N_17900,N_18507);
nand UO_1694 (O_1694,N_19666,N_18899);
and UO_1695 (O_1695,N_17267,N_19335);
or UO_1696 (O_1696,N_18495,N_19751);
nor UO_1697 (O_1697,N_19104,N_18286);
nor UO_1698 (O_1698,N_17287,N_19072);
nor UO_1699 (O_1699,N_19312,N_19914);
nor UO_1700 (O_1700,N_18243,N_17404);
and UO_1701 (O_1701,N_16446,N_17772);
and UO_1702 (O_1702,N_18446,N_19371);
and UO_1703 (O_1703,N_17741,N_19536);
and UO_1704 (O_1704,N_17149,N_16341);
and UO_1705 (O_1705,N_18254,N_17781);
or UO_1706 (O_1706,N_18695,N_17098);
and UO_1707 (O_1707,N_17717,N_19249);
nand UO_1708 (O_1708,N_18631,N_16526);
and UO_1709 (O_1709,N_16086,N_18079);
nand UO_1710 (O_1710,N_16326,N_18003);
and UO_1711 (O_1711,N_18842,N_17044);
or UO_1712 (O_1712,N_19229,N_18133);
and UO_1713 (O_1713,N_17958,N_18476);
and UO_1714 (O_1714,N_16543,N_19894);
or UO_1715 (O_1715,N_18684,N_18428);
or UO_1716 (O_1716,N_18904,N_18100);
nand UO_1717 (O_1717,N_16849,N_17303);
nor UO_1718 (O_1718,N_19247,N_17425);
or UO_1719 (O_1719,N_18097,N_18263);
or UO_1720 (O_1720,N_18769,N_16012);
nand UO_1721 (O_1721,N_17714,N_16743);
or UO_1722 (O_1722,N_19956,N_18485);
and UO_1723 (O_1723,N_18444,N_16166);
and UO_1724 (O_1724,N_16548,N_16080);
nor UO_1725 (O_1725,N_19224,N_17130);
or UO_1726 (O_1726,N_16894,N_17491);
nor UO_1727 (O_1727,N_16559,N_16068);
nor UO_1728 (O_1728,N_17118,N_18464);
nor UO_1729 (O_1729,N_16891,N_17695);
and UO_1730 (O_1730,N_17295,N_18701);
and UO_1731 (O_1731,N_17918,N_17088);
nand UO_1732 (O_1732,N_16153,N_16379);
or UO_1733 (O_1733,N_16040,N_18336);
nand UO_1734 (O_1734,N_18633,N_17821);
and UO_1735 (O_1735,N_18541,N_18578);
or UO_1736 (O_1736,N_17147,N_17389);
nor UO_1737 (O_1737,N_18604,N_17426);
nand UO_1738 (O_1738,N_17042,N_18311);
xor UO_1739 (O_1739,N_19605,N_19574);
nand UO_1740 (O_1740,N_17111,N_19211);
nand UO_1741 (O_1741,N_17481,N_16573);
or UO_1742 (O_1742,N_18599,N_18044);
nand UO_1743 (O_1743,N_19059,N_19086);
xor UO_1744 (O_1744,N_17929,N_18375);
nor UO_1745 (O_1745,N_16788,N_19480);
or UO_1746 (O_1746,N_18004,N_17321);
nor UO_1747 (O_1747,N_19178,N_16900);
nand UO_1748 (O_1748,N_19796,N_18114);
nand UO_1749 (O_1749,N_18147,N_17114);
nor UO_1750 (O_1750,N_19410,N_19239);
nor UO_1751 (O_1751,N_16255,N_18558);
nand UO_1752 (O_1752,N_17345,N_18220);
and UO_1753 (O_1753,N_18488,N_17155);
nor UO_1754 (O_1754,N_16896,N_18978);
or UO_1755 (O_1755,N_16100,N_18582);
nor UO_1756 (O_1756,N_19850,N_17343);
or UO_1757 (O_1757,N_19720,N_16770);
and UO_1758 (O_1758,N_19523,N_17007);
or UO_1759 (O_1759,N_19601,N_16146);
and UO_1760 (O_1760,N_16525,N_19082);
xnor UO_1761 (O_1761,N_17536,N_16398);
nand UO_1762 (O_1762,N_19933,N_17412);
or UO_1763 (O_1763,N_16105,N_19906);
nor UO_1764 (O_1764,N_16979,N_17561);
and UO_1765 (O_1765,N_16216,N_19575);
nand UO_1766 (O_1766,N_17783,N_19015);
nor UO_1767 (O_1767,N_19994,N_19001);
or UO_1768 (O_1768,N_18725,N_17097);
or UO_1769 (O_1769,N_17688,N_17587);
nor UO_1770 (O_1770,N_16637,N_19907);
or UO_1771 (O_1771,N_16487,N_19112);
and UO_1772 (O_1772,N_18680,N_17786);
nand UO_1773 (O_1773,N_19887,N_18627);
nand UO_1774 (O_1774,N_18840,N_16870);
nand UO_1775 (O_1775,N_19584,N_16233);
or UO_1776 (O_1776,N_16997,N_16630);
or UO_1777 (O_1777,N_18645,N_16783);
xnor UO_1778 (O_1778,N_18007,N_16545);
xnor UO_1779 (O_1779,N_16685,N_16605);
or UO_1780 (O_1780,N_19863,N_18155);
nand UO_1781 (O_1781,N_16950,N_18264);
xor UO_1782 (O_1782,N_16114,N_19232);
nor UO_1783 (O_1783,N_18296,N_16832);
nor UO_1784 (O_1784,N_18121,N_16749);
xnor UO_1785 (O_1785,N_18076,N_19477);
and UO_1786 (O_1786,N_19669,N_18338);
and UO_1787 (O_1787,N_16322,N_18111);
nand UO_1788 (O_1788,N_19831,N_19286);
nand UO_1789 (O_1789,N_17622,N_17868);
and UO_1790 (O_1790,N_19550,N_17729);
or UO_1791 (O_1791,N_17941,N_19846);
nor UO_1792 (O_1792,N_16708,N_19707);
and UO_1793 (O_1793,N_16296,N_17450);
or UO_1794 (O_1794,N_16316,N_19320);
or UO_1795 (O_1795,N_17582,N_18252);
nor UO_1796 (O_1796,N_17206,N_19000);
nand UO_1797 (O_1797,N_19435,N_16892);
nand UO_1798 (O_1798,N_19374,N_19031);
nand UO_1799 (O_1799,N_16263,N_16789);
or UO_1800 (O_1800,N_19052,N_17458);
and UO_1801 (O_1801,N_16334,N_18918);
and UO_1802 (O_1802,N_17479,N_16181);
and UO_1803 (O_1803,N_18176,N_16760);
nor UO_1804 (O_1804,N_19199,N_18596);
and UO_1805 (O_1805,N_18841,N_16112);
or UO_1806 (O_1806,N_16145,N_16589);
nor UO_1807 (O_1807,N_16225,N_17670);
or UO_1808 (O_1808,N_17684,N_18072);
and UO_1809 (O_1809,N_19495,N_17482);
nand UO_1810 (O_1810,N_19396,N_19509);
or UO_1811 (O_1811,N_19672,N_18750);
nand UO_1812 (O_1812,N_17887,N_17391);
and UO_1813 (O_1813,N_18399,N_18576);
nand UO_1814 (O_1814,N_18135,N_16747);
nand UO_1815 (O_1815,N_18575,N_19834);
or UO_1816 (O_1816,N_18462,N_18470);
or UO_1817 (O_1817,N_19430,N_17047);
or UO_1818 (O_1818,N_17667,N_19185);
nor UO_1819 (O_1819,N_19965,N_16961);
nor UO_1820 (O_1820,N_19649,N_16838);
or UO_1821 (O_1821,N_16390,N_17658);
and UO_1822 (O_1822,N_16682,N_18770);
nand UO_1823 (O_1823,N_18078,N_19778);
and UO_1824 (O_1824,N_18229,N_17936);
and UO_1825 (O_1825,N_18267,N_17739);
and UO_1826 (O_1826,N_18991,N_16828);
nand UO_1827 (O_1827,N_17547,N_16777);
and UO_1828 (O_1828,N_19231,N_16264);
or UO_1829 (O_1829,N_18696,N_18879);
and UO_1830 (O_1830,N_18948,N_16866);
nand UO_1831 (O_1831,N_18897,N_19879);
nand UO_1832 (O_1832,N_17270,N_18503);
and UO_1833 (O_1833,N_16087,N_16681);
and UO_1834 (O_1834,N_17166,N_19123);
or UO_1835 (O_1835,N_17546,N_19936);
and UO_1836 (O_1836,N_19142,N_17419);
nor UO_1837 (O_1837,N_19726,N_16536);
and UO_1838 (O_1838,N_18673,N_19014);
nor UO_1839 (O_1839,N_16871,N_18206);
nand UO_1840 (O_1840,N_16437,N_19117);
nor UO_1841 (O_1841,N_17794,N_18817);
and UO_1842 (O_1842,N_18297,N_16612);
and UO_1843 (O_1843,N_18392,N_19971);
and UO_1844 (O_1844,N_16647,N_19746);
nor UO_1845 (O_1845,N_18564,N_19140);
or UO_1846 (O_1846,N_18215,N_19986);
or UO_1847 (O_1847,N_17716,N_16250);
nand UO_1848 (O_1848,N_17612,N_18644);
nor UO_1849 (O_1849,N_18134,N_16013);
nand UO_1850 (O_1850,N_16888,N_18182);
nand UO_1851 (O_1851,N_19262,N_19297);
nand UO_1852 (O_1852,N_19343,N_16756);
and UO_1853 (O_1853,N_19110,N_18218);
nor UO_1854 (O_1854,N_17613,N_19070);
and UO_1855 (O_1855,N_19499,N_18580);
nor UO_1856 (O_1856,N_18447,N_17668);
nor UO_1857 (O_1857,N_19519,N_16740);
or UO_1858 (O_1858,N_19571,N_18248);
and UO_1859 (O_1859,N_18914,N_17564);
nand UO_1860 (O_1860,N_18328,N_19812);
and UO_1861 (O_1861,N_17597,N_19252);
nand UO_1862 (O_1862,N_19245,N_17468);
or UO_1863 (O_1863,N_17792,N_19839);
nor UO_1864 (O_1864,N_17038,N_16119);
nand UO_1865 (O_1865,N_16116,N_18808);
and UO_1866 (O_1866,N_17850,N_16911);
or UO_1867 (O_1867,N_19375,N_17071);
nor UO_1868 (O_1868,N_19567,N_18751);
or UO_1869 (O_1869,N_16057,N_16809);
nor UO_1870 (O_1870,N_17748,N_19998);
nor UO_1871 (O_1871,N_17956,N_19884);
nand UO_1872 (O_1872,N_19527,N_19336);
and UO_1873 (O_1873,N_18360,N_16032);
and UO_1874 (O_1874,N_17971,N_18335);
nand UO_1875 (O_1875,N_19721,N_18993);
nand UO_1876 (O_1876,N_16875,N_18595);
or UO_1877 (O_1877,N_19733,N_19289);
nand UO_1878 (O_1878,N_18070,N_17304);
and UO_1879 (O_1879,N_17516,N_17362);
and UO_1880 (O_1880,N_16024,N_19102);
or UO_1881 (O_1881,N_17034,N_17198);
nand UO_1882 (O_1882,N_18230,N_18973);
nor UO_1883 (O_1883,N_17774,N_16073);
or UO_1884 (O_1884,N_16771,N_18735);
nor UO_1885 (O_1885,N_16669,N_17685);
and UO_1886 (O_1886,N_16967,N_17378);
or UO_1887 (O_1887,N_19992,N_17837);
nor UO_1888 (O_1888,N_19545,N_19532);
nor UO_1889 (O_1889,N_17242,N_19294);
nand UO_1890 (O_1890,N_16458,N_19448);
and UO_1891 (O_1891,N_16699,N_17453);
or UO_1892 (O_1892,N_17019,N_19900);
or UO_1893 (O_1893,N_19489,N_16347);
nand UO_1894 (O_1894,N_17961,N_16754);
and UO_1895 (O_1895,N_19961,N_16461);
nand UO_1896 (O_1896,N_19922,N_18760);
and UO_1897 (O_1897,N_18214,N_19652);
nand UO_1898 (O_1898,N_16212,N_17592);
or UO_1899 (O_1899,N_19351,N_17078);
xor UO_1900 (O_1900,N_17843,N_19732);
and UO_1901 (O_1901,N_19702,N_19981);
nand UO_1902 (O_1902,N_19240,N_16909);
nand UO_1903 (O_1903,N_17533,N_18207);
nor UO_1904 (O_1904,N_16730,N_16127);
nand UO_1905 (O_1905,N_19534,N_17762);
nand UO_1906 (O_1906,N_16769,N_16143);
and UO_1907 (O_1907,N_19041,N_16232);
or UO_1908 (O_1908,N_18357,N_19711);
nor UO_1909 (O_1909,N_18715,N_19356);
or UO_1910 (O_1910,N_17175,N_18435);
or UO_1911 (O_1911,N_17846,N_16566);
xor UO_1912 (O_1912,N_18632,N_19848);
or UO_1913 (O_1913,N_17083,N_16268);
or UO_1914 (O_1914,N_19661,N_18172);
nand UO_1915 (O_1915,N_18954,N_16120);
nand UO_1916 (O_1916,N_16660,N_17917);
nand UO_1917 (O_1917,N_16286,N_17893);
or UO_1918 (O_1918,N_18591,N_19319);
and UO_1919 (O_1919,N_19553,N_18650);
nand UO_1920 (O_1920,N_18940,N_16969);
nand UO_1921 (O_1921,N_18955,N_19197);
nand UO_1922 (O_1922,N_16088,N_18227);
nand UO_1923 (O_1923,N_19767,N_18683);
nor UO_1924 (O_1924,N_17966,N_19755);
and UO_1925 (O_1925,N_17171,N_19373);
nor UO_1926 (O_1926,N_18131,N_16355);
and UO_1927 (O_1927,N_18626,N_17795);
nand UO_1928 (O_1928,N_18972,N_19520);
nand UO_1929 (O_1929,N_17571,N_18855);
nor UO_1930 (O_1930,N_16065,N_16357);
and UO_1931 (O_1931,N_18326,N_19827);
and UO_1932 (O_1932,N_17897,N_19910);
or UO_1933 (O_1933,N_17376,N_18344);
nor UO_1934 (O_1934,N_19369,N_17405);
or UO_1935 (O_1935,N_19482,N_17833);
nand UO_1936 (O_1936,N_17767,N_18681);
and UO_1937 (O_1937,N_16549,N_17445);
nand UO_1938 (O_1938,N_18140,N_19855);
nor UO_1939 (O_1939,N_19542,N_17138);
and UO_1940 (O_1940,N_17318,N_19551);
nand UO_1941 (O_1941,N_16108,N_17416);
nor UO_1942 (O_1942,N_17403,N_17447);
nand UO_1943 (O_1943,N_19694,N_16778);
nor UO_1944 (O_1944,N_17525,N_19087);
or UO_1945 (O_1945,N_16137,N_16593);
xor UO_1946 (O_1946,N_17237,N_16269);
and UO_1947 (O_1947,N_18866,N_18347);
nand UO_1948 (O_1948,N_18720,N_18567);
nor UO_1949 (O_1949,N_17880,N_18323);
or UO_1950 (O_1950,N_18438,N_17693);
nand UO_1951 (O_1951,N_18965,N_16084);
nor UO_1952 (O_1952,N_17127,N_18483);
and UO_1953 (O_1953,N_17497,N_19439);
and UO_1954 (O_1954,N_16066,N_19768);
or UO_1955 (O_1955,N_17535,N_17465);
nor UO_1956 (O_1956,N_17115,N_19953);
and UO_1957 (O_1957,N_19427,N_17841);
nor UO_1958 (O_1958,N_18552,N_16387);
nand UO_1959 (O_1959,N_16856,N_18061);
and UO_1960 (O_1960,N_17572,N_19737);
or UO_1961 (O_1961,N_17834,N_16103);
nand UO_1962 (O_1962,N_16943,N_16034);
or UO_1963 (O_1963,N_17650,N_17620);
nor UO_1964 (O_1964,N_16665,N_17144);
or UO_1965 (O_1965,N_16450,N_19621);
and UO_1966 (O_1966,N_16562,N_16959);
nand UO_1967 (O_1967,N_19632,N_18881);
xor UO_1968 (O_1968,N_17276,N_16423);
or UO_1969 (O_1969,N_19273,N_16841);
nand UO_1970 (O_1970,N_17452,N_17393);
and UO_1971 (O_1971,N_19172,N_18737);
nand UO_1972 (O_1972,N_19071,N_19020);
or UO_1973 (O_1973,N_18797,N_17804);
or UO_1974 (O_1974,N_19530,N_16400);
nor UO_1975 (O_1975,N_16134,N_18692);
nor UO_1976 (O_1976,N_16333,N_16466);
and UO_1977 (O_1977,N_16098,N_18589);
nand UO_1978 (O_1978,N_19949,N_18385);
and UO_1979 (O_1979,N_19033,N_19888);
and UO_1980 (O_1980,N_16178,N_16597);
nand UO_1981 (O_1981,N_17316,N_19843);
nand UO_1982 (O_1982,N_19736,N_18937);
nor UO_1983 (O_1983,N_17305,N_19365);
xor UO_1984 (O_1984,N_17172,N_19691);
nand UO_1985 (O_1985,N_16261,N_18949);
nor UO_1986 (O_1986,N_18657,N_18923);
or UO_1987 (O_1987,N_18784,N_16472);
and UO_1988 (O_1988,N_18472,N_19201);
nor UO_1989 (O_1989,N_18945,N_17059);
nand UO_1990 (O_1990,N_19870,N_18398);
and UO_1991 (O_1991,N_16349,N_17174);
nor UO_1992 (O_1992,N_19593,N_18322);
or UO_1993 (O_1993,N_18884,N_17923);
xnor UO_1994 (O_1994,N_16781,N_18546);
and UO_1995 (O_1995,N_18391,N_17805);
and UO_1996 (O_1996,N_18523,N_17241);
nor UO_1997 (O_1997,N_18074,N_18465);
nand UO_1998 (O_1998,N_16733,N_18661);
nand UO_1999 (O_1999,N_17703,N_19423);
or UO_2000 (O_2000,N_16659,N_16847);
and UO_2001 (O_2001,N_17177,N_19288);
and UO_2002 (O_2002,N_16073,N_19553);
nand UO_2003 (O_2003,N_17536,N_16093);
or UO_2004 (O_2004,N_19970,N_17072);
nand UO_2005 (O_2005,N_17237,N_19327);
or UO_2006 (O_2006,N_19850,N_18939);
nor UO_2007 (O_2007,N_17187,N_18288);
nand UO_2008 (O_2008,N_16104,N_17856);
and UO_2009 (O_2009,N_18050,N_17169);
nor UO_2010 (O_2010,N_18322,N_16448);
and UO_2011 (O_2011,N_18709,N_17475);
nand UO_2012 (O_2012,N_16488,N_19470);
nor UO_2013 (O_2013,N_19083,N_18656);
or UO_2014 (O_2014,N_17861,N_16186);
or UO_2015 (O_2015,N_16732,N_16367);
nand UO_2016 (O_2016,N_18772,N_16728);
nand UO_2017 (O_2017,N_18681,N_18080);
or UO_2018 (O_2018,N_18858,N_19581);
nor UO_2019 (O_2019,N_18298,N_17973);
nand UO_2020 (O_2020,N_19445,N_16499);
xnor UO_2021 (O_2021,N_16093,N_17591);
and UO_2022 (O_2022,N_16762,N_17300);
or UO_2023 (O_2023,N_17940,N_17924);
and UO_2024 (O_2024,N_19919,N_17625);
and UO_2025 (O_2025,N_18292,N_16516);
nand UO_2026 (O_2026,N_16963,N_16269);
or UO_2027 (O_2027,N_19707,N_17957);
and UO_2028 (O_2028,N_19485,N_18579);
nand UO_2029 (O_2029,N_16881,N_19152);
nor UO_2030 (O_2030,N_17714,N_19641);
nor UO_2031 (O_2031,N_18561,N_18853);
nor UO_2032 (O_2032,N_17028,N_16714);
and UO_2033 (O_2033,N_16504,N_18921);
nor UO_2034 (O_2034,N_18051,N_17193);
nor UO_2035 (O_2035,N_17838,N_17828);
and UO_2036 (O_2036,N_17847,N_18349);
nand UO_2037 (O_2037,N_18604,N_18347);
and UO_2038 (O_2038,N_19688,N_19759);
nor UO_2039 (O_2039,N_17116,N_17931);
or UO_2040 (O_2040,N_17710,N_19896);
and UO_2041 (O_2041,N_19812,N_18232);
or UO_2042 (O_2042,N_16338,N_19762);
nor UO_2043 (O_2043,N_18767,N_17243);
nand UO_2044 (O_2044,N_18693,N_16674);
nor UO_2045 (O_2045,N_19498,N_16621);
nand UO_2046 (O_2046,N_18805,N_16521);
nor UO_2047 (O_2047,N_19643,N_19113);
nand UO_2048 (O_2048,N_19812,N_19801);
nand UO_2049 (O_2049,N_18177,N_18868);
or UO_2050 (O_2050,N_19229,N_18159);
and UO_2051 (O_2051,N_18390,N_17347);
nor UO_2052 (O_2052,N_18839,N_18763);
nor UO_2053 (O_2053,N_17099,N_19030);
nand UO_2054 (O_2054,N_19794,N_16961);
nand UO_2055 (O_2055,N_17806,N_17998);
or UO_2056 (O_2056,N_19408,N_17211);
or UO_2057 (O_2057,N_18763,N_17224);
nor UO_2058 (O_2058,N_16268,N_19449);
nor UO_2059 (O_2059,N_19314,N_16885);
nor UO_2060 (O_2060,N_18643,N_16799);
or UO_2061 (O_2061,N_16975,N_18886);
and UO_2062 (O_2062,N_18070,N_16612);
nor UO_2063 (O_2063,N_16056,N_19652);
or UO_2064 (O_2064,N_18783,N_18042);
or UO_2065 (O_2065,N_19408,N_19072);
nor UO_2066 (O_2066,N_17731,N_18046);
nor UO_2067 (O_2067,N_18695,N_16756);
and UO_2068 (O_2068,N_19068,N_18662);
or UO_2069 (O_2069,N_18589,N_19952);
nor UO_2070 (O_2070,N_17435,N_18208);
or UO_2071 (O_2071,N_16317,N_19008);
and UO_2072 (O_2072,N_18155,N_18957);
or UO_2073 (O_2073,N_18329,N_18316);
or UO_2074 (O_2074,N_16283,N_17292);
nor UO_2075 (O_2075,N_17958,N_17886);
or UO_2076 (O_2076,N_18802,N_16462);
or UO_2077 (O_2077,N_17885,N_19374);
nand UO_2078 (O_2078,N_17425,N_18084);
and UO_2079 (O_2079,N_16883,N_16143);
or UO_2080 (O_2080,N_19988,N_17333);
and UO_2081 (O_2081,N_16700,N_19246);
and UO_2082 (O_2082,N_16076,N_19713);
and UO_2083 (O_2083,N_16200,N_17840);
or UO_2084 (O_2084,N_19469,N_19406);
nor UO_2085 (O_2085,N_16808,N_18836);
nand UO_2086 (O_2086,N_16793,N_17081);
or UO_2087 (O_2087,N_17199,N_17598);
nor UO_2088 (O_2088,N_18892,N_17572);
nor UO_2089 (O_2089,N_17114,N_19844);
and UO_2090 (O_2090,N_17842,N_19238);
or UO_2091 (O_2091,N_17405,N_18968);
nand UO_2092 (O_2092,N_17835,N_18649);
or UO_2093 (O_2093,N_17811,N_17185);
nor UO_2094 (O_2094,N_18343,N_16051);
nor UO_2095 (O_2095,N_18338,N_18486);
nor UO_2096 (O_2096,N_19577,N_17985);
and UO_2097 (O_2097,N_19931,N_17750);
nand UO_2098 (O_2098,N_18008,N_16493);
nor UO_2099 (O_2099,N_16488,N_16718);
nand UO_2100 (O_2100,N_19024,N_16234);
nand UO_2101 (O_2101,N_16350,N_16970);
nand UO_2102 (O_2102,N_16848,N_16335);
or UO_2103 (O_2103,N_19916,N_19001);
and UO_2104 (O_2104,N_19321,N_17036);
or UO_2105 (O_2105,N_19839,N_18997);
nand UO_2106 (O_2106,N_17826,N_16764);
or UO_2107 (O_2107,N_19415,N_19364);
nor UO_2108 (O_2108,N_18325,N_18866);
nor UO_2109 (O_2109,N_17621,N_18222);
and UO_2110 (O_2110,N_16567,N_19108);
nor UO_2111 (O_2111,N_16714,N_17799);
or UO_2112 (O_2112,N_19981,N_17196);
nand UO_2113 (O_2113,N_19422,N_17543);
and UO_2114 (O_2114,N_19008,N_16200);
nor UO_2115 (O_2115,N_16795,N_16233);
or UO_2116 (O_2116,N_16899,N_19724);
or UO_2117 (O_2117,N_18506,N_16816);
nor UO_2118 (O_2118,N_18241,N_19754);
nor UO_2119 (O_2119,N_18220,N_16411);
or UO_2120 (O_2120,N_19197,N_16138);
and UO_2121 (O_2121,N_18720,N_18972);
and UO_2122 (O_2122,N_19121,N_18331);
nor UO_2123 (O_2123,N_19233,N_17871);
nor UO_2124 (O_2124,N_17254,N_18062);
or UO_2125 (O_2125,N_18271,N_18484);
nor UO_2126 (O_2126,N_17986,N_19061);
and UO_2127 (O_2127,N_18061,N_16948);
and UO_2128 (O_2128,N_16085,N_17776);
and UO_2129 (O_2129,N_18678,N_17247);
nor UO_2130 (O_2130,N_19672,N_18857);
nand UO_2131 (O_2131,N_18225,N_19588);
or UO_2132 (O_2132,N_17805,N_17758);
nor UO_2133 (O_2133,N_18603,N_16022);
nor UO_2134 (O_2134,N_18223,N_19714);
nand UO_2135 (O_2135,N_19048,N_16188);
nand UO_2136 (O_2136,N_16962,N_16821);
nand UO_2137 (O_2137,N_16044,N_16534);
and UO_2138 (O_2138,N_19482,N_19564);
and UO_2139 (O_2139,N_18697,N_17593);
nand UO_2140 (O_2140,N_19138,N_18547);
nand UO_2141 (O_2141,N_17239,N_16215);
and UO_2142 (O_2142,N_17357,N_19468);
or UO_2143 (O_2143,N_18881,N_19672);
nand UO_2144 (O_2144,N_16626,N_19824);
or UO_2145 (O_2145,N_18255,N_18448);
or UO_2146 (O_2146,N_17141,N_18423);
nand UO_2147 (O_2147,N_18064,N_16100);
and UO_2148 (O_2148,N_17680,N_19965);
nor UO_2149 (O_2149,N_17959,N_18634);
and UO_2150 (O_2150,N_19046,N_18494);
xor UO_2151 (O_2151,N_19751,N_18963);
or UO_2152 (O_2152,N_16048,N_18043);
and UO_2153 (O_2153,N_17429,N_18365);
nor UO_2154 (O_2154,N_17650,N_16694);
and UO_2155 (O_2155,N_19448,N_18462);
nand UO_2156 (O_2156,N_16687,N_17773);
and UO_2157 (O_2157,N_16043,N_17076);
or UO_2158 (O_2158,N_19437,N_19165);
nand UO_2159 (O_2159,N_16571,N_16498);
nand UO_2160 (O_2160,N_19788,N_18444);
nand UO_2161 (O_2161,N_16337,N_19041);
nor UO_2162 (O_2162,N_18041,N_19419);
xor UO_2163 (O_2163,N_17233,N_17987);
nand UO_2164 (O_2164,N_17394,N_18463);
nor UO_2165 (O_2165,N_18031,N_18559);
nand UO_2166 (O_2166,N_17575,N_17195);
and UO_2167 (O_2167,N_18765,N_17163);
nand UO_2168 (O_2168,N_19151,N_19972);
nand UO_2169 (O_2169,N_19611,N_19252);
and UO_2170 (O_2170,N_18348,N_16334);
and UO_2171 (O_2171,N_16093,N_19875);
and UO_2172 (O_2172,N_17974,N_18602);
nand UO_2173 (O_2173,N_16632,N_17496);
and UO_2174 (O_2174,N_18683,N_17862);
and UO_2175 (O_2175,N_18067,N_18519);
xor UO_2176 (O_2176,N_18667,N_18301);
and UO_2177 (O_2177,N_19512,N_17943);
nor UO_2178 (O_2178,N_19232,N_19382);
nor UO_2179 (O_2179,N_16521,N_19603);
or UO_2180 (O_2180,N_16351,N_17044);
nor UO_2181 (O_2181,N_19339,N_19285);
nand UO_2182 (O_2182,N_16202,N_19537);
nor UO_2183 (O_2183,N_16455,N_17950);
and UO_2184 (O_2184,N_16216,N_17004);
nor UO_2185 (O_2185,N_19915,N_16571);
nand UO_2186 (O_2186,N_19978,N_19174);
nand UO_2187 (O_2187,N_18334,N_16827);
nand UO_2188 (O_2188,N_16575,N_18203);
nor UO_2189 (O_2189,N_17784,N_17121);
nand UO_2190 (O_2190,N_17814,N_18870);
nor UO_2191 (O_2191,N_16047,N_16411);
or UO_2192 (O_2192,N_16417,N_18983);
and UO_2193 (O_2193,N_17239,N_19360);
or UO_2194 (O_2194,N_16322,N_17737);
nor UO_2195 (O_2195,N_17935,N_16711);
nor UO_2196 (O_2196,N_17058,N_18764);
nand UO_2197 (O_2197,N_16474,N_19416);
or UO_2198 (O_2198,N_19383,N_18942);
nand UO_2199 (O_2199,N_16557,N_18749);
nor UO_2200 (O_2200,N_17043,N_19015);
and UO_2201 (O_2201,N_17313,N_16357);
or UO_2202 (O_2202,N_18498,N_17296);
nor UO_2203 (O_2203,N_17336,N_18969);
or UO_2204 (O_2204,N_19936,N_19810);
nor UO_2205 (O_2205,N_19482,N_17163);
nand UO_2206 (O_2206,N_18734,N_19023);
nand UO_2207 (O_2207,N_17484,N_18565);
nand UO_2208 (O_2208,N_16890,N_16342);
and UO_2209 (O_2209,N_16207,N_16576);
nor UO_2210 (O_2210,N_16946,N_19638);
nor UO_2211 (O_2211,N_17300,N_18369);
nor UO_2212 (O_2212,N_16304,N_17034);
or UO_2213 (O_2213,N_16745,N_17868);
and UO_2214 (O_2214,N_18656,N_19347);
nand UO_2215 (O_2215,N_17990,N_18214);
and UO_2216 (O_2216,N_17896,N_18469);
or UO_2217 (O_2217,N_18426,N_18654);
nor UO_2218 (O_2218,N_17497,N_17469);
or UO_2219 (O_2219,N_16731,N_19312);
or UO_2220 (O_2220,N_19806,N_18424);
nor UO_2221 (O_2221,N_16473,N_19548);
nor UO_2222 (O_2222,N_17446,N_18429);
nand UO_2223 (O_2223,N_16469,N_18684);
nand UO_2224 (O_2224,N_18950,N_17587);
and UO_2225 (O_2225,N_19870,N_16135);
or UO_2226 (O_2226,N_18347,N_18858);
nand UO_2227 (O_2227,N_16038,N_16485);
and UO_2228 (O_2228,N_16312,N_18550);
and UO_2229 (O_2229,N_16047,N_17156);
nor UO_2230 (O_2230,N_17751,N_16029);
nand UO_2231 (O_2231,N_18479,N_17421);
nor UO_2232 (O_2232,N_18256,N_18131);
or UO_2233 (O_2233,N_18335,N_17111);
or UO_2234 (O_2234,N_17522,N_16616);
nor UO_2235 (O_2235,N_18039,N_19092);
and UO_2236 (O_2236,N_18442,N_18218);
nor UO_2237 (O_2237,N_18533,N_19328);
or UO_2238 (O_2238,N_17517,N_19011);
nand UO_2239 (O_2239,N_16395,N_19054);
nor UO_2240 (O_2240,N_17353,N_17060);
and UO_2241 (O_2241,N_18817,N_18124);
or UO_2242 (O_2242,N_17825,N_18077);
nor UO_2243 (O_2243,N_18324,N_18959);
and UO_2244 (O_2244,N_18872,N_19739);
and UO_2245 (O_2245,N_19155,N_19383);
and UO_2246 (O_2246,N_18144,N_17795);
nor UO_2247 (O_2247,N_18596,N_18487);
nand UO_2248 (O_2248,N_16566,N_19630);
and UO_2249 (O_2249,N_19805,N_17245);
nor UO_2250 (O_2250,N_19969,N_16541);
and UO_2251 (O_2251,N_16868,N_17622);
and UO_2252 (O_2252,N_18503,N_16382);
and UO_2253 (O_2253,N_17694,N_17334);
nand UO_2254 (O_2254,N_19812,N_19923);
nand UO_2255 (O_2255,N_16837,N_19966);
nor UO_2256 (O_2256,N_19984,N_17776);
and UO_2257 (O_2257,N_19321,N_16694);
and UO_2258 (O_2258,N_18794,N_16979);
nor UO_2259 (O_2259,N_18684,N_19645);
and UO_2260 (O_2260,N_17029,N_18645);
nand UO_2261 (O_2261,N_18205,N_16363);
nand UO_2262 (O_2262,N_18972,N_19061);
and UO_2263 (O_2263,N_19900,N_17450);
nand UO_2264 (O_2264,N_17815,N_19972);
or UO_2265 (O_2265,N_19483,N_17130);
or UO_2266 (O_2266,N_17772,N_16997);
xnor UO_2267 (O_2267,N_17938,N_18369);
or UO_2268 (O_2268,N_18071,N_18908);
nand UO_2269 (O_2269,N_19250,N_18235);
or UO_2270 (O_2270,N_16285,N_18669);
nand UO_2271 (O_2271,N_18455,N_19160);
nand UO_2272 (O_2272,N_17404,N_17829);
nand UO_2273 (O_2273,N_19125,N_16104);
or UO_2274 (O_2274,N_18488,N_17432);
nand UO_2275 (O_2275,N_16401,N_18895);
nand UO_2276 (O_2276,N_17816,N_16267);
and UO_2277 (O_2277,N_17288,N_18596);
and UO_2278 (O_2278,N_16574,N_19645);
or UO_2279 (O_2279,N_17102,N_19317);
nand UO_2280 (O_2280,N_19160,N_17286);
and UO_2281 (O_2281,N_16827,N_19669);
or UO_2282 (O_2282,N_17384,N_16353);
or UO_2283 (O_2283,N_18810,N_19743);
nor UO_2284 (O_2284,N_17946,N_18363);
nand UO_2285 (O_2285,N_18025,N_19158);
nor UO_2286 (O_2286,N_19490,N_18711);
or UO_2287 (O_2287,N_17446,N_16171);
nor UO_2288 (O_2288,N_16702,N_16818);
nor UO_2289 (O_2289,N_17234,N_18290);
or UO_2290 (O_2290,N_19929,N_17156);
or UO_2291 (O_2291,N_18358,N_18609);
nor UO_2292 (O_2292,N_18919,N_16815);
nor UO_2293 (O_2293,N_16834,N_17602);
and UO_2294 (O_2294,N_18028,N_19790);
nor UO_2295 (O_2295,N_17038,N_18217);
nand UO_2296 (O_2296,N_18017,N_18522);
or UO_2297 (O_2297,N_19666,N_17066);
or UO_2298 (O_2298,N_17436,N_18800);
or UO_2299 (O_2299,N_16401,N_17741);
and UO_2300 (O_2300,N_19270,N_16192);
and UO_2301 (O_2301,N_18091,N_18430);
xnor UO_2302 (O_2302,N_17530,N_18693);
xor UO_2303 (O_2303,N_19857,N_17452);
or UO_2304 (O_2304,N_18191,N_16304);
and UO_2305 (O_2305,N_19586,N_16168);
nor UO_2306 (O_2306,N_16245,N_18137);
nor UO_2307 (O_2307,N_16284,N_19585);
nand UO_2308 (O_2308,N_18148,N_18408);
nor UO_2309 (O_2309,N_19863,N_17907);
nor UO_2310 (O_2310,N_17227,N_19988);
or UO_2311 (O_2311,N_18024,N_16708);
xnor UO_2312 (O_2312,N_18731,N_18171);
and UO_2313 (O_2313,N_19517,N_17796);
or UO_2314 (O_2314,N_18287,N_17417);
nor UO_2315 (O_2315,N_17797,N_16175);
nor UO_2316 (O_2316,N_18315,N_17779);
nor UO_2317 (O_2317,N_17764,N_16129);
nand UO_2318 (O_2318,N_16468,N_17006);
nor UO_2319 (O_2319,N_16070,N_19139);
nor UO_2320 (O_2320,N_19479,N_18806);
or UO_2321 (O_2321,N_19049,N_19353);
and UO_2322 (O_2322,N_17417,N_16307);
nor UO_2323 (O_2323,N_16230,N_16799);
nand UO_2324 (O_2324,N_17999,N_16674);
or UO_2325 (O_2325,N_17480,N_18652);
nor UO_2326 (O_2326,N_19236,N_18416);
or UO_2327 (O_2327,N_18849,N_17880);
and UO_2328 (O_2328,N_18002,N_17484);
nand UO_2329 (O_2329,N_19904,N_19459);
or UO_2330 (O_2330,N_19478,N_17379);
or UO_2331 (O_2331,N_18115,N_18689);
nor UO_2332 (O_2332,N_17390,N_17527);
nor UO_2333 (O_2333,N_16064,N_18921);
nor UO_2334 (O_2334,N_16680,N_18537);
nor UO_2335 (O_2335,N_17782,N_19072);
and UO_2336 (O_2336,N_16105,N_17844);
nand UO_2337 (O_2337,N_17178,N_18736);
nor UO_2338 (O_2338,N_16932,N_16614);
and UO_2339 (O_2339,N_17971,N_16534);
nor UO_2340 (O_2340,N_17897,N_17434);
nor UO_2341 (O_2341,N_16079,N_16884);
or UO_2342 (O_2342,N_18771,N_17788);
nor UO_2343 (O_2343,N_19584,N_16190);
or UO_2344 (O_2344,N_16361,N_16592);
nand UO_2345 (O_2345,N_16649,N_18344);
or UO_2346 (O_2346,N_18009,N_17588);
or UO_2347 (O_2347,N_16141,N_19131);
or UO_2348 (O_2348,N_17343,N_16317);
nor UO_2349 (O_2349,N_16049,N_18960);
nor UO_2350 (O_2350,N_17623,N_17032);
and UO_2351 (O_2351,N_16009,N_17371);
or UO_2352 (O_2352,N_18482,N_18353);
nand UO_2353 (O_2353,N_16683,N_17931);
nand UO_2354 (O_2354,N_19309,N_17282);
nor UO_2355 (O_2355,N_17207,N_19309);
nand UO_2356 (O_2356,N_19211,N_16756);
or UO_2357 (O_2357,N_16287,N_17052);
nand UO_2358 (O_2358,N_18754,N_16708);
and UO_2359 (O_2359,N_17169,N_18176);
or UO_2360 (O_2360,N_19206,N_16964);
and UO_2361 (O_2361,N_18839,N_17048);
nand UO_2362 (O_2362,N_16667,N_19713);
nor UO_2363 (O_2363,N_19789,N_17131);
nand UO_2364 (O_2364,N_17630,N_17735);
and UO_2365 (O_2365,N_18209,N_17978);
nor UO_2366 (O_2366,N_18079,N_17827);
and UO_2367 (O_2367,N_17385,N_18027);
or UO_2368 (O_2368,N_18777,N_16599);
nand UO_2369 (O_2369,N_16036,N_18907);
or UO_2370 (O_2370,N_18869,N_18255);
or UO_2371 (O_2371,N_16947,N_16225);
nor UO_2372 (O_2372,N_16233,N_18771);
nand UO_2373 (O_2373,N_16886,N_18667);
and UO_2374 (O_2374,N_19727,N_18919);
and UO_2375 (O_2375,N_19560,N_16371);
and UO_2376 (O_2376,N_17288,N_17067);
xnor UO_2377 (O_2377,N_16552,N_17243);
or UO_2378 (O_2378,N_18518,N_17842);
or UO_2379 (O_2379,N_18709,N_16612);
and UO_2380 (O_2380,N_19906,N_17262);
or UO_2381 (O_2381,N_19023,N_17800);
nand UO_2382 (O_2382,N_19723,N_18766);
nand UO_2383 (O_2383,N_19973,N_16401);
and UO_2384 (O_2384,N_16296,N_16117);
nor UO_2385 (O_2385,N_16976,N_18236);
nor UO_2386 (O_2386,N_19530,N_16640);
and UO_2387 (O_2387,N_19116,N_16458);
or UO_2388 (O_2388,N_16681,N_18684);
nor UO_2389 (O_2389,N_19492,N_18545);
nand UO_2390 (O_2390,N_18450,N_17516);
and UO_2391 (O_2391,N_17001,N_18575);
nand UO_2392 (O_2392,N_16118,N_19375);
and UO_2393 (O_2393,N_17989,N_16932);
and UO_2394 (O_2394,N_17407,N_17478);
or UO_2395 (O_2395,N_16087,N_18659);
nand UO_2396 (O_2396,N_19344,N_16051);
and UO_2397 (O_2397,N_18040,N_18589);
or UO_2398 (O_2398,N_17237,N_16715);
nor UO_2399 (O_2399,N_16950,N_16941);
or UO_2400 (O_2400,N_17576,N_19685);
nor UO_2401 (O_2401,N_18430,N_18664);
and UO_2402 (O_2402,N_16942,N_19638);
and UO_2403 (O_2403,N_17413,N_19374);
nor UO_2404 (O_2404,N_17882,N_17733);
nand UO_2405 (O_2405,N_18932,N_19773);
and UO_2406 (O_2406,N_18340,N_19235);
nor UO_2407 (O_2407,N_16715,N_19695);
or UO_2408 (O_2408,N_17896,N_16245);
nor UO_2409 (O_2409,N_16474,N_16773);
nand UO_2410 (O_2410,N_17688,N_19329);
nor UO_2411 (O_2411,N_17515,N_17944);
or UO_2412 (O_2412,N_19721,N_19663);
nand UO_2413 (O_2413,N_17988,N_18362);
or UO_2414 (O_2414,N_17712,N_19947);
nand UO_2415 (O_2415,N_17093,N_18188);
nor UO_2416 (O_2416,N_18263,N_16907);
or UO_2417 (O_2417,N_19178,N_18346);
or UO_2418 (O_2418,N_16960,N_19844);
nor UO_2419 (O_2419,N_18101,N_18306);
and UO_2420 (O_2420,N_18651,N_17785);
or UO_2421 (O_2421,N_18469,N_17331);
nand UO_2422 (O_2422,N_17085,N_16367);
or UO_2423 (O_2423,N_19919,N_17820);
nor UO_2424 (O_2424,N_18895,N_19331);
nand UO_2425 (O_2425,N_19240,N_19788);
nor UO_2426 (O_2426,N_17896,N_19496);
and UO_2427 (O_2427,N_17111,N_17534);
or UO_2428 (O_2428,N_19705,N_17085);
or UO_2429 (O_2429,N_19416,N_19380);
or UO_2430 (O_2430,N_17877,N_16848);
or UO_2431 (O_2431,N_18986,N_18116);
xor UO_2432 (O_2432,N_19346,N_17593);
or UO_2433 (O_2433,N_18862,N_16323);
or UO_2434 (O_2434,N_16232,N_19924);
nor UO_2435 (O_2435,N_19238,N_18894);
nor UO_2436 (O_2436,N_17745,N_17346);
or UO_2437 (O_2437,N_18109,N_16503);
or UO_2438 (O_2438,N_17903,N_16864);
or UO_2439 (O_2439,N_16364,N_19993);
and UO_2440 (O_2440,N_17444,N_16981);
nor UO_2441 (O_2441,N_18763,N_16906);
nor UO_2442 (O_2442,N_18478,N_16541);
nor UO_2443 (O_2443,N_19268,N_19164);
xnor UO_2444 (O_2444,N_17679,N_18262);
nand UO_2445 (O_2445,N_19468,N_16918);
nand UO_2446 (O_2446,N_16532,N_19376);
or UO_2447 (O_2447,N_19025,N_19391);
xor UO_2448 (O_2448,N_16809,N_18275);
or UO_2449 (O_2449,N_17391,N_16895);
nor UO_2450 (O_2450,N_17370,N_17516);
or UO_2451 (O_2451,N_17873,N_19044);
and UO_2452 (O_2452,N_16556,N_16811);
and UO_2453 (O_2453,N_16793,N_19512);
nand UO_2454 (O_2454,N_16278,N_16570);
or UO_2455 (O_2455,N_18744,N_18886);
or UO_2456 (O_2456,N_17133,N_18926);
nor UO_2457 (O_2457,N_17120,N_16911);
nand UO_2458 (O_2458,N_19966,N_19329);
nor UO_2459 (O_2459,N_17733,N_17537);
or UO_2460 (O_2460,N_18447,N_18251);
and UO_2461 (O_2461,N_18108,N_17898);
nor UO_2462 (O_2462,N_16898,N_16077);
nand UO_2463 (O_2463,N_18141,N_16099);
and UO_2464 (O_2464,N_19464,N_16339);
and UO_2465 (O_2465,N_17200,N_16858);
nor UO_2466 (O_2466,N_16219,N_19905);
nor UO_2467 (O_2467,N_18537,N_18109);
or UO_2468 (O_2468,N_18303,N_19753);
and UO_2469 (O_2469,N_19409,N_19336);
nor UO_2470 (O_2470,N_16220,N_18925);
nor UO_2471 (O_2471,N_18291,N_19742);
nand UO_2472 (O_2472,N_18000,N_17795);
or UO_2473 (O_2473,N_19011,N_16588);
nor UO_2474 (O_2474,N_19417,N_18882);
nor UO_2475 (O_2475,N_17673,N_17549);
and UO_2476 (O_2476,N_16944,N_16502);
and UO_2477 (O_2477,N_16700,N_18572);
and UO_2478 (O_2478,N_19280,N_16876);
and UO_2479 (O_2479,N_17480,N_16825);
nor UO_2480 (O_2480,N_18121,N_19396);
nand UO_2481 (O_2481,N_17661,N_17266);
nor UO_2482 (O_2482,N_16720,N_16719);
or UO_2483 (O_2483,N_17596,N_18450);
or UO_2484 (O_2484,N_18013,N_16753);
and UO_2485 (O_2485,N_18673,N_17050);
and UO_2486 (O_2486,N_18243,N_16968);
nor UO_2487 (O_2487,N_18604,N_19471);
and UO_2488 (O_2488,N_16860,N_18223);
and UO_2489 (O_2489,N_19788,N_17457);
nand UO_2490 (O_2490,N_19494,N_18306);
nand UO_2491 (O_2491,N_16104,N_18472);
or UO_2492 (O_2492,N_19008,N_17418);
and UO_2493 (O_2493,N_18277,N_18551);
nand UO_2494 (O_2494,N_19822,N_17829);
and UO_2495 (O_2495,N_18482,N_18672);
nor UO_2496 (O_2496,N_17535,N_16284);
and UO_2497 (O_2497,N_17164,N_18357);
nand UO_2498 (O_2498,N_16790,N_19273);
or UO_2499 (O_2499,N_16169,N_18696);
endmodule