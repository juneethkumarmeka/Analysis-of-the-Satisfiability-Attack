module basic_1000_10000_1500_4_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_145,In_739);
nand U1 (N_1,In_7,In_210);
and U2 (N_2,In_472,In_955);
nand U3 (N_3,In_759,In_932);
nor U4 (N_4,In_698,In_872);
or U5 (N_5,In_552,In_610);
nand U6 (N_6,In_352,In_405);
nand U7 (N_7,In_276,In_599);
nand U8 (N_8,In_369,In_485);
or U9 (N_9,In_650,In_306);
nor U10 (N_10,In_709,In_956);
nand U11 (N_11,In_526,In_200);
and U12 (N_12,In_152,In_434);
nor U13 (N_13,In_738,In_917);
nand U14 (N_14,In_179,In_656);
nand U15 (N_15,In_962,In_520);
nor U16 (N_16,In_398,In_300);
or U17 (N_17,In_879,In_451);
nand U18 (N_18,In_227,In_784);
nand U19 (N_19,In_742,In_201);
or U20 (N_20,In_726,In_802);
and U21 (N_21,In_565,In_176);
nand U22 (N_22,In_418,In_333);
nand U23 (N_23,In_861,In_59);
nor U24 (N_24,In_589,In_634);
nor U25 (N_25,In_484,In_312);
nand U26 (N_26,In_743,In_517);
or U27 (N_27,In_142,In_875);
nor U28 (N_28,In_797,In_211);
or U29 (N_29,In_389,In_426);
nand U30 (N_30,In_416,In_617);
or U31 (N_31,In_919,In_551);
or U32 (N_32,In_880,In_354);
nor U33 (N_33,In_275,In_323);
or U34 (N_34,In_453,In_625);
or U35 (N_35,In_81,In_162);
nand U36 (N_36,In_186,In_423);
nand U37 (N_37,In_606,In_713);
nand U38 (N_38,In_869,In_342);
or U39 (N_39,In_672,In_721);
or U40 (N_40,In_615,In_512);
nor U41 (N_41,In_645,In_490);
and U42 (N_42,In_251,In_464);
nand U43 (N_43,In_776,In_307);
or U44 (N_44,In_791,In_263);
nor U45 (N_45,In_437,In_278);
nand U46 (N_46,In_222,In_786);
or U47 (N_47,In_335,In_429);
nor U48 (N_48,In_487,In_384);
nand U49 (N_49,In_224,In_848);
nand U50 (N_50,In_385,In_737);
and U51 (N_51,In_936,In_193);
nor U52 (N_52,In_885,In_97);
and U53 (N_53,In_403,In_62);
or U54 (N_54,In_581,In_387);
and U55 (N_55,In_24,In_580);
or U56 (N_56,In_202,In_190);
nor U57 (N_57,In_697,In_447);
and U58 (N_58,In_772,In_233);
nor U59 (N_59,In_121,In_213);
or U60 (N_60,In_229,In_769);
nand U61 (N_61,In_89,In_184);
and U62 (N_62,In_253,In_185);
nor U63 (N_63,In_724,In_994);
and U64 (N_64,In_728,In_740);
nor U65 (N_65,In_432,In_35);
nor U66 (N_66,In_545,In_42);
or U67 (N_67,In_970,In_468);
nor U68 (N_68,In_481,In_667);
nor U69 (N_69,In_456,In_865);
and U70 (N_70,In_11,In_668);
nor U71 (N_71,In_63,In_633);
and U72 (N_72,In_639,In_789);
or U73 (N_73,In_58,In_735);
or U74 (N_74,In_979,In_187);
nor U75 (N_75,In_706,In_958);
nor U76 (N_76,In_264,In_167);
nand U77 (N_77,In_191,In_685);
nor U78 (N_78,In_569,In_584);
nor U79 (N_79,In_341,In_290);
nand U80 (N_80,In_65,In_654);
or U81 (N_81,In_273,In_47);
or U82 (N_82,In_553,In_46);
or U83 (N_83,In_324,In_678);
nand U84 (N_84,In_614,In_216);
nor U85 (N_85,In_501,In_281);
nand U86 (N_86,In_326,In_431);
and U87 (N_87,In_86,In_414);
or U88 (N_88,In_840,In_923);
nor U89 (N_89,In_477,In_198);
nor U90 (N_90,In_659,In_799);
or U91 (N_91,In_987,In_670);
nor U92 (N_92,In_831,In_636);
nor U93 (N_93,In_531,In_887);
nor U94 (N_94,In_541,In_394);
nor U95 (N_95,In_22,In_635);
and U96 (N_96,In_949,In_538);
and U97 (N_97,In_792,In_514);
nor U98 (N_98,In_367,In_988);
or U99 (N_99,In_856,In_37);
or U100 (N_100,In_108,In_124);
or U101 (N_101,In_572,In_19);
nor U102 (N_102,In_741,In_542);
and U103 (N_103,In_683,In_401);
nand U104 (N_104,In_469,In_128);
nor U105 (N_105,In_295,In_171);
nor U106 (N_106,In_376,In_313);
nand U107 (N_107,In_417,In_149);
or U108 (N_108,In_82,In_924);
nand U109 (N_109,In_379,In_12);
and U110 (N_110,In_293,In_116);
or U111 (N_111,In_87,In_353);
and U112 (N_112,In_357,In_274);
and U113 (N_113,In_556,In_498);
and U114 (N_114,In_262,In_360);
nand U115 (N_115,In_812,In_348);
or U116 (N_116,In_876,In_653);
or U117 (N_117,In_460,In_444);
nand U118 (N_118,In_340,In_494);
nand U119 (N_119,In_246,In_72);
nor U120 (N_120,In_2,In_813);
and U121 (N_121,In_647,In_648);
nor U122 (N_122,In_180,In_199);
and U123 (N_123,In_240,In_985);
or U124 (N_124,In_359,In_903);
and U125 (N_125,In_252,In_934);
nand U126 (N_126,In_129,In_155);
nor U127 (N_127,In_952,In_302);
or U128 (N_128,In_286,In_623);
nor U129 (N_129,In_242,In_515);
and U130 (N_130,In_60,In_957);
and U131 (N_131,In_337,In_440);
or U132 (N_132,In_627,In_356);
and U133 (N_133,In_132,In_669);
or U134 (N_134,In_343,In_36);
nor U135 (N_135,In_753,In_810);
nor U136 (N_136,In_691,In_704);
nand U137 (N_137,In_806,In_297);
and U138 (N_138,In_871,In_798);
or U139 (N_139,In_752,In_311);
nand U140 (N_140,In_680,In_539);
or U141 (N_141,In_732,In_504);
and U142 (N_142,In_57,In_622);
or U143 (N_143,In_762,In_33);
and U144 (N_144,In_43,In_347);
and U145 (N_145,In_996,In_393);
nor U146 (N_146,In_349,In_800);
nand U147 (N_147,In_30,In_696);
nand U148 (N_148,In_820,In_513);
or U149 (N_149,In_154,In_906);
or U150 (N_150,In_649,In_819);
nor U151 (N_151,In_510,In_744);
and U152 (N_152,In_409,In_954);
or U153 (N_153,In_68,In_272);
nor U154 (N_154,In_466,In_334);
nand U155 (N_155,In_383,In_913);
and U156 (N_156,In_266,In_104);
nand U157 (N_157,In_172,In_603);
or U158 (N_158,In_974,In_587);
and U159 (N_159,In_549,In_849);
or U160 (N_160,In_9,In_712);
nand U161 (N_161,In_972,In_688);
and U162 (N_162,In_548,In_345);
nand U163 (N_163,In_236,In_953);
nor U164 (N_164,In_908,In_136);
nand U165 (N_165,In_321,In_567);
nor U166 (N_166,In_767,In_404);
and U167 (N_167,In_138,In_117);
nand U168 (N_168,In_506,In_938);
nor U169 (N_169,In_50,In_305);
and U170 (N_170,In_443,In_363);
or U171 (N_171,In_38,In_845);
nand U172 (N_172,In_768,In_226);
nand U173 (N_173,In_44,In_463);
nor U174 (N_174,In_14,In_568);
nor U175 (N_175,In_45,In_106);
nor U176 (N_176,In_257,In_571);
nand U177 (N_177,In_984,In_407);
nor U178 (N_178,In_771,In_935);
nor U179 (N_179,In_143,In_566);
nand U180 (N_180,In_937,In_716);
and U181 (N_181,In_13,In_616);
nand U182 (N_182,In_904,In_748);
or U183 (N_183,In_110,In_554);
nand U184 (N_184,In_694,In_787);
or U185 (N_185,In_632,In_818);
nor U186 (N_186,In_505,In_564);
nand U187 (N_187,In_245,In_521);
nor U188 (N_188,In_465,In_316);
and U189 (N_189,In_746,In_159);
and U190 (N_190,In_722,In_594);
nor U191 (N_191,In_339,In_918);
and U192 (N_192,In_399,In_239);
and U193 (N_193,In_61,In_663);
nor U194 (N_194,In_835,In_986);
nand U195 (N_195,In_682,In_84);
nor U196 (N_196,In_32,In_577);
nand U197 (N_197,In_146,In_674);
and U198 (N_198,In_518,In_930);
and U199 (N_199,In_194,In_854);
and U200 (N_200,In_248,In_543);
and U201 (N_201,In_26,In_288);
nand U202 (N_202,In_372,In_609);
and U203 (N_203,In_419,In_449);
nor U204 (N_204,In_225,In_509);
and U205 (N_205,In_249,In_1);
or U206 (N_206,In_950,In_891);
and U207 (N_207,In_782,In_575);
nand U208 (N_208,In_710,In_220);
nor U209 (N_209,In_626,In_476);
or U210 (N_210,In_424,In_592);
nand U211 (N_211,In_579,In_999);
and U212 (N_212,In_829,In_751);
nor U213 (N_213,In_79,In_303);
or U214 (N_214,In_330,In_600);
and U215 (N_215,In_530,In_174);
nand U216 (N_216,In_754,In_676);
or U217 (N_217,In_665,In_516);
or U218 (N_218,In_230,In_34);
nand U219 (N_219,In_692,In_749);
nand U220 (N_220,In_20,In_758);
nor U221 (N_221,In_408,In_486);
or U222 (N_222,In_18,In_804);
and U223 (N_223,In_382,In_99);
nand U224 (N_224,In_166,In_178);
xor U225 (N_225,In_452,In_964);
and U226 (N_226,In_168,In_315);
nor U227 (N_227,In_247,In_846);
nor U228 (N_228,In_939,In_107);
nand U229 (N_229,In_80,In_375);
or U230 (N_230,In_708,In_458);
nand U231 (N_231,In_147,In_719);
or U232 (N_232,In_783,In_977);
nand U233 (N_233,In_183,In_836);
or U234 (N_234,In_329,In_666);
nand U235 (N_235,In_889,In_470);
nor U236 (N_236,In_314,In_338);
xor U237 (N_237,In_827,In_137);
nor U238 (N_238,In_282,In_396);
nor U239 (N_239,In_662,In_319);
nor U240 (N_240,In_700,In_111);
nor U241 (N_241,In_40,In_661);
nand U242 (N_242,In_140,In_350);
and U243 (N_243,In_850,In_157);
and U244 (N_244,In_978,In_914);
or U245 (N_245,In_844,In_318);
nand U246 (N_246,In_277,In_816);
and U247 (N_247,In_997,In_292);
and U248 (N_248,In_215,In_714);
or U249 (N_249,In_660,In_637);
and U250 (N_250,In_862,In_777);
or U251 (N_251,In_85,In_294);
or U252 (N_252,In_995,In_53);
or U253 (N_253,In_165,In_943);
nand U254 (N_254,In_493,In_134);
or U255 (N_255,In_991,In_825);
nand U256 (N_256,In_638,In_896);
nand U257 (N_257,In_406,In_322);
or U258 (N_258,In_448,In_640);
or U259 (N_259,In_95,In_163);
and U260 (N_260,In_838,In_973);
nor U261 (N_261,In_90,In_528);
nand U262 (N_262,In_234,In_64);
and U263 (N_263,In_673,In_677);
nor U264 (N_264,In_809,In_852);
nor U265 (N_265,In_534,In_28);
or U266 (N_266,In_915,In_100);
nor U267 (N_267,In_781,In_595);
and U268 (N_268,In_540,In_940);
nand U269 (N_269,In_3,In_675);
or U270 (N_270,In_899,In_892);
and U271 (N_271,In_894,In_817);
nor U272 (N_272,In_750,In_808);
or U273 (N_273,In_878,In_495);
nor U274 (N_274,In_911,In_15);
nand U275 (N_275,In_31,In_392);
or U276 (N_276,In_355,In_438);
and U277 (N_277,In_830,In_241);
nand U278 (N_278,In_285,In_150);
and U279 (N_279,In_902,In_886);
nor U280 (N_280,In_88,In_83);
and U281 (N_281,In_944,In_982);
nand U282 (N_282,In_93,In_629);
nand U283 (N_283,In_55,In_371);
or U284 (N_284,In_169,In_259);
nand U285 (N_285,In_544,In_467);
and U286 (N_286,In_441,In_268);
or U287 (N_287,In_681,In_52);
nor U288 (N_288,In_841,In_400);
nor U289 (N_289,In_963,In_898);
and U290 (N_290,In_907,In_555);
or U291 (N_291,In_118,In_188);
and U292 (N_292,In_482,In_537);
and U293 (N_293,In_182,In_17);
nor U294 (N_294,In_821,In_427);
or U295 (N_295,In_664,In_496);
nor U296 (N_296,In_25,In_561);
and U297 (N_297,In_428,In_320);
nand U298 (N_298,In_612,In_267);
nand U299 (N_299,In_283,In_583);
or U300 (N_300,In_926,In_101);
nor U301 (N_301,In_959,In_679);
and U302 (N_302,In_796,In_27);
nand U303 (N_303,In_261,In_547);
nor U304 (N_304,In_402,In_655);
nand U305 (N_305,In_597,In_364);
or U306 (N_306,In_492,In_279);
and U307 (N_307,In_430,In_527);
nor U308 (N_308,In_446,In_232);
and U309 (N_309,In_833,In_843);
nor U310 (N_310,In_702,In_578);
or U311 (N_311,In_73,In_975);
or U312 (N_312,In_803,In_559);
nand U313 (N_313,In_192,In_299);
nand U314 (N_314,In_435,In_790);
and U315 (N_315,In_927,In_29);
or U316 (N_316,In_961,In_112);
nand U317 (N_317,In_671,In_524);
nand U318 (N_318,In_863,In_102);
and U319 (N_319,In_601,In_828);
nand U320 (N_320,In_951,In_920);
xnor U321 (N_321,In_207,In_851);
or U322 (N_322,In_703,In_223);
and U323 (N_323,In_832,In_814);
and U324 (N_324,In_49,In_374);
nand U325 (N_325,In_373,In_618);
and U326 (N_326,In_455,In_66);
nand U327 (N_327,In_76,In_195);
nor U328 (N_328,In_442,In_701);
and U329 (N_329,In_41,In_6);
nand U330 (N_330,In_270,In_642);
nand U331 (N_331,In_717,In_388);
nor U332 (N_332,In_380,In_491);
nand U333 (N_333,In_855,In_868);
and U334 (N_334,In_151,In_502);
nand U335 (N_335,In_361,In_945);
or U336 (N_336,In_362,In_218);
nand U337 (N_337,In_309,In_631);
or U338 (N_338,In_461,In_933);
nand U339 (N_339,In_582,In_127);
nor U340 (N_340,In_258,In_98);
or U341 (N_341,In_96,In_250);
nor U342 (N_342,In_822,In_105);
nand U343 (N_343,In_707,In_115);
and U344 (N_344,In_237,In_459);
nand U345 (N_345,In_882,In_901);
nor U346 (N_346,In_756,In_895);
nand U347 (N_347,In_328,In_280);
nor U348 (N_348,In_170,In_536);
nor U349 (N_349,In_607,In_588);
nand U350 (N_350,In_826,In_546);
nor U351 (N_351,In_770,In_815);
nand U352 (N_352,In_327,In_624);
nor U353 (N_353,In_238,In_523);
and U354 (N_354,In_734,In_308);
nand U355 (N_355,In_805,In_761);
or U356 (N_356,In_420,In_929);
or U357 (N_357,In_8,In_499);
and U358 (N_358,In_503,In_763);
and U359 (N_359,In_658,In_109);
or U360 (N_360,In_197,In_126);
or U361 (N_361,In_585,In_968);
nand U362 (N_362,In_228,In_471);
or U363 (N_363,In_344,In_120);
nor U364 (N_364,In_160,In_877);
or U365 (N_365,In_103,In_204);
nand U366 (N_366,In_508,In_765);
nor U367 (N_367,In_0,In_386);
nor U368 (N_368,In_941,In_39);
and U369 (N_369,In_346,In_764);
and U370 (N_370,In_593,In_71);
and U371 (N_371,In_890,In_947);
and U372 (N_372,In_203,In_693);
nor U373 (N_373,In_243,In_859);
or U374 (N_374,In_525,In_173);
nor U375 (N_375,In_867,In_175);
or U376 (N_376,In_590,In_10);
or U377 (N_377,In_395,In_883);
or U378 (N_378,In_760,In_628);
or U379 (N_379,In_421,In_834);
nand U380 (N_380,In_507,In_265);
or U381 (N_381,In_687,In_390);
nand U382 (N_382,In_370,In_874);
or U383 (N_383,In_221,In_269);
xor U384 (N_384,In_412,In_921);
nand U385 (N_385,In_591,In_522);
and U386 (N_386,In_774,In_310);
nor U387 (N_387,In_425,In_77);
nor U388 (N_388,In_870,In_156);
or U389 (N_389,In_92,In_766);
nor U390 (N_390,In_780,In_596);
nor U391 (N_391,In_793,In_158);
nand U392 (N_392,In_646,In_657);
nand U393 (N_393,In_535,In_897);
nor U394 (N_394,In_946,In_271);
nor U395 (N_395,In_317,In_980);
or U396 (N_396,In_839,In_332);
and U397 (N_397,In_928,In_21);
nor U398 (N_398,In_212,In_570);
nand U399 (N_399,In_489,In_550);
nand U400 (N_400,In_711,In_990);
nand U401 (N_401,In_720,In_873);
or U402 (N_402,In_148,In_778);
nor U403 (N_403,In_260,In_16);
nand U404 (N_404,In_368,In_235);
nand U405 (N_405,In_613,In_298);
or U406 (N_406,In_358,In_445);
or U407 (N_407,In_699,In_351);
nor U408 (N_408,In_966,In_775);
or U409 (N_409,In_70,In_289);
and U410 (N_410,In_847,In_860);
nor U411 (N_411,In_133,In_910);
nand U412 (N_412,In_557,In_244);
nor U413 (N_413,In_651,In_900);
nor U414 (N_414,In_325,In_256);
or U415 (N_415,In_478,In_377);
nand U416 (N_416,In_866,In_189);
and U417 (N_417,In_51,In_916);
nor U418 (N_418,In_336,In_969);
and U419 (N_419,In_153,In_113);
or U420 (N_420,In_532,In_811);
and U421 (N_421,In_391,In_718);
and U422 (N_422,In_415,In_139);
nor U423 (N_423,In_123,In_563);
or U424 (N_424,In_439,In_284);
and U425 (N_425,In_993,In_255);
nor U426 (N_426,In_287,In_208);
nand U427 (N_427,In_365,In_67);
nor U428 (N_428,In_652,In_745);
nor U429 (N_429,In_690,In_620);
nand U430 (N_430,In_948,In_586);
or U431 (N_431,In_795,In_981);
or U432 (N_432,In_196,In_644);
and U433 (N_433,In_942,In_598);
nor U434 (N_434,In_574,In_807);
nand U435 (N_435,In_511,In_976);
and U436 (N_436,In_122,In_558);
nor U437 (N_437,In_378,In_56);
or U438 (N_438,In_705,In_967);
nand U439 (N_439,In_462,In_733);
xnor U440 (N_440,In_960,In_621);
nand U441 (N_441,In_164,In_983);
nand U442 (N_442,In_864,In_209);
or U443 (N_443,In_130,In_480);
and U444 (N_444,In_643,In_608);
and U445 (N_445,In_450,In_433);
or U446 (N_446,In_161,In_881);
nor U447 (N_447,In_231,In_736);
nand U448 (N_448,In_695,In_965);
or U449 (N_449,In_78,In_135);
and U450 (N_450,In_757,In_747);
nor U451 (N_451,In_205,In_837);
and U452 (N_452,In_125,In_304);
nand U453 (N_453,In_641,In_729);
nor U454 (N_454,In_630,In_773);
nand U455 (N_455,In_366,In_54);
xor U456 (N_456,In_331,In_131);
nand U457 (N_457,In_119,In_560);
nand U458 (N_458,In_785,In_301);
nor U459 (N_459,In_893,In_611);
nor U460 (N_460,In_483,In_5);
nand U461 (N_461,In_931,In_602);
nor U462 (N_462,In_992,In_731);
nand U463 (N_463,In_686,In_413);
and U464 (N_464,In_214,In_619);
or U465 (N_465,In_144,In_562);
or U466 (N_466,In_605,In_23);
nor U467 (N_467,In_801,In_457);
nor U468 (N_468,In_989,In_475);
nor U469 (N_469,In_254,In_823);
or U470 (N_470,In_909,In_500);
or U471 (N_471,In_884,In_715);
and U472 (N_472,In_888,In_217);
and U473 (N_473,In_206,In_474);
nand U474 (N_474,In_779,In_689);
nor U475 (N_475,In_488,In_497);
and U476 (N_476,In_48,In_75);
nor U477 (N_477,In_177,In_912);
and U478 (N_478,In_454,In_411);
and U479 (N_479,In_94,In_181);
nor U480 (N_480,In_794,In_727);
and U481 (N_481,In_69,In_533);
or U482 (N_482,In_922,In_576);
or U483 (N_483,In_755,In_397);
or U484 (N_484,In_998,In_436);
or U485 (N_485,In_857,In_905);
nand U486 (N_486,In_853,In_141);
nand U487 (N_487,In_4,In_725);
and U488 (N_488,In_519,In_479);
and U489 (N_489,In_925,In_296);
nand U490 (N_490,In_422,In_573);
xor U491 (N_491,In_824,In_91);
or U492 (N_492,In_858,In_114);
or U493 (N_493,In_219,In_74);
nor U494 (N_494,In_604,In_971);
and U495 (N_495,In_788,In_529);
nand U496 (N_496,In_381,In_473);
or U497 (N_497,In_291,In_684);
nor U498 (N_498,In_842,In_730);
nor U499 (N_499,In_723,In_410);
and U500 (N_500,In_674,In_927);
or U501 (N_501,In_114,In_87);
and U502 (N_502,In_64,In_120);
nor U503 (N_503,In_413,In_305);
and U504 (N_504,In_473,In_58);
xor U505 (N_505,In_903,In_769);
or U506 (N_506,In_667,In_55);
nand U507 (N_507,In_752,In_278);
nor U508 (N_508,In_315,In_29);
nor U509 (N_509,In_440,In_533);
or U510 (N_510,In_785,In_52);
nand U511 (N_511,In_746,In_122);
nand U512 (N_512,In_736,In_669);
or U513 (N_513,In_10,In_929);
nand U514 (N_514,In_7,In_909);
nor U515 (N_515,In_588,In_53);
nor U516 (N_516,In_264,In_648);
nand U517 (N_517,In_762,In_527);
and U518 (N_518,In_113,In_280);
or U519 (N_519,In_416,In_379);
or U520 (N_520,In_456,In_931);
nand U521 (N_521,In_128,In_172);
or U522 (N_522,In_445,In_258);
nand U523 (N_523,In_272,In_1);
or U524 (N_524,In_543,In_101);
or U525 (N_525,In_365,In_305);
or U526 (N_526,In_183,In_661);
and U527 (N_527,In_831,In_551);
and U528 (N_528,In_539,In_237);
or U529 (N_529,In_964,In_85);
nand U530 (N_530,In_665,In_504);
or U531 (N_531,In_881,In_182);
or U532 (N_532,In_204,In_21);
and U533 (N_533,In_496,In_294);
or U534 (N_534,In_665,In_760);
nor U535 (N_535,In_186,In_721);
and U536 (N_536,In_322,In_207);
or U537 (N_537,In_80,In_59);
nor U538 (N_538,In_73,In_524);
xor U539 (N_539,In_650,In_557);
and U540 (N_540,In_811,In_788);
nand U541 (N_541,In_776,In_471);
nor U542 (N_542,In_596,In_169);
and U543 (N_543,In_429,In_651);
nand U544 (N_544,In_363,In_988);
nand U545 (N_545,In_904,In_722);
nand U546 (N_546,In_619,In_275);
and U547 (N_547,In_412,In_841);
or U548 (N_548,In_519,In_875);
xnor U549 (N_549,In_174,In_527);
nor U550 (N_550,In_505,In_770);
and U551 (N_551,In_183,In_513);
nor U552 (N_552,In_386,In_683);
and U553 (N_553,In_424,In_119);
or U554 (N_554,In_433,In_839);
and U555 (N_555,In_234,In_538);
nand U556 (N_556,In_829,In_144);
and U557 (N_557,In_731,In_476);
and U558 (N_558,In_781,In_226);
nand U559 (N_559,In_272,In_692);
nand U560 (N_560,In_6,In_0);
and U561 (N_561,In_244,In_370);
or U562 (N_562,In_912,In_784);
and U563 (N_563,In_30,In_430);
nor U564 (N_564,In_648,In_416);
nand U565 (N_565,In_904,In_808);
or U566 (N_566,In_688,In_298);
and U567 (N_567,In_447,In_540);
or U568 (N_568,In_803,In_673);
nor U569 (N_569,In_311,In_979);
or U570 (N_570,In_125,In_858);
nand U571 (N_571,In_873,In_17);
nand U572 (N_572,In_997,In_921);
or U573 (N_573,In_199,In_569);
nand U574 (N_574,In_17,In_998);
or U575 (N_575,In_881,In_912);
or U576 (N_576,In_244,In_610);
nand U577 (N_577,In_691,In_581);
nand U578 (N_578,In_718,In_709);
nand U579 (N_579,In_227,In_212);
or U580 (N_580,In_319,In_748);
and U581 (N_581,In_973,In_368);
and U582 (N_582,In_589,In_83);
or U583 (N_583,In_140,In_642);
and U584 (N_584,In_895,In_809);
nand U585 (N_585,In_705,In_143);
or U586 (N_586,In_182,In_430);
or U587 (N_587,In_737,In_946);
and U588 (N_588,In_465,In_497);
and U589 (N_589,In_737,In_468);
nor U590 (N_590,In_55,In_21);
nor U591 (N_591,In_661,In_806);
nor U592 (N_592,In_518,In_343);
nand U593 (N_593,In_848,In_762);
nand U594 (N_594,In_128,In_921);
nand U595 (N_595,In_477,In_916);
nor U596 (N_596,In_216,In_337);
or U597 (N_597,In_281,In_324);
or U598 (N_598,In_707,In_837);
nor U599 (N_599,In_855,In_311);
or U600 (N_600,In_580,In_283);
and U601 (N_601,In_895,In_536);
nor U602 (N_602,In_455,In_770);
nor U603 (N_603,In_779,In_838);
nand U604 (N_604,In_523,In_540);
and U605 (N_605,In_573,In_8);
and U606 (N_606,In_51,In_238);
or U607 (N_607,In_720,In_469);
nor U608 (N_608,In_928,In_27);
nor U609 (N_609,In_298,In_273);
nand U610 (N_610,In_655,In_909);
nor U611 (N_611,In_482,In_404);
nor U612 (N_612,In_40,In_802);
nand U613 (N_613,In_705,In_384);
nor U614 (N_614,In_877,In_7);
or U615 (N_615,In_143,In_35);
or U616 (N_616,In_192,In_992);
nand U617 (N_617,In_655,In_569);
or U618 (N_618,In_869,In_809);
and U619 (N_619,In_609,In_332);
and U620 (N_620,In_447,In_777);
and U621 (N_621,In_171,In_930);
nor U622 (N_622,In_396,In_10);
nand U623 (N_623,In_39,In_965);
or U624 (N_624,In_588,In_312);
and U625 (N_625,In_845,In_955);
nand U626 (N_626,In_509,In_920);
nor U627 (N_627,In_755,In_466);
and U628 (N_628,In_685,In_962);
nand U629 (N_629,In_461,In_3);
nor U630 (N_630,In_232,In_372);
and U631 (N_631,In_977,In_879);
and U632 (N_632,In_329,In_723);
nor U633 (N_633,In_657,In_279);
and U634 (N_634,In_723,In_144);
or U635 (N_635,In_750,In_787);
nor U636 (N_636,In_814,In_914);
nand U637 (N_637,In_547,In_263);
nand U638 (N_638,In_335,In_169);
nor U639 (N_639,In_863,In_226);
and U640 (N_640,In_271,In_466);
nand U641 (N_641,In_333,In_68);
or U642 (N_642,In_568,In_381);
nand U643 (N_643,In_267,In_627);
nor U644 (N_644,In_189,In_862);
nand U645 (N_645,In_998,In_755);
or U646 (N_646,In_326,In_985);
or U647 (N_647,In_683,In_277);
and U648 (N_648,In_866,In_677);
nor U649 (N_649,In_148,In_816);
nand U650 (N_650,In_591,In_248);
and U651 (N_651,In_797,In_625);
nand U652 (N_652,In_577,In_162);
or U653 (N_653,In_171,In_736);
or U654 (N_654,In_752,In_620);
and U655 (N_655,In_284,In_427);
nand U656 (N_656,In_953,In_892);
nand U657 (N_657,In_340,In_252);
or U658 (N_658,In_595,In_363);
nand U659 (N_659,In_392,In_455);
nand U660 (N_660,In_65,In_469);
and U661 (N_661,In_155,In_860);
or U662 (N_662,In_316,In_283);
nor U663 (N_663,In_843,In_46);
and U664 (N_664,In_991,In_197);
and U665 (N_665,In_921,In_956);
or U666 (N_666,In_450,In_4);
nand U667 (N_667,In_748,In_123);
nand U668 (N_668,In_44,In_411);
nor U669 (N_669,In_731,In_565);
nand U670 (N_670,In_839,In_365);
or U671 (N_671,In_395,In_811);
nand U672 (N_672,In_89,In_764);
or U673 (N_673,In_976,In_852);
and U674 (N_674,In_893,In_815);
nor U675 (N_675,In_639,In_302);
and U676 (N_676,In_426,In_342);
or U677 (N_677,In_799,In_594);
nor U678 (N_678,In_705,In_50);
nor U679 (N_679,In_933,In_193);
nor U680 (N_680,In_347,In_902);
nand U681 (N_681,In_848,In_203);
and U682 (N_682,In_372,In_333);
or U683 (N_683,In_174,In_25);
nor U684 (N_684,In_647,In_8);
xor U685 (N_685,In_958,In_818);
nand U686 (N_686,In_752,In_730);
and U687 (N_687,In_337,In_324);
nand U688 (N_688,In_221,In_44);
nor U689 (N_689,In_124,In_302);
nand U690 (N_690,In_854,In_85);
nor U691 (N_691,In_654,In_68);
nand U692 (N_692,In_884,In_159);
nand U693 (N_693,In_120,In_415);
and U694 (N_694,In_915,In_226);
and U695 (N_695,In_909,In_952);
nor U696 (N_696,In_331,In_254);
nor U697 (N_697,In_375,In_356);
nand U698 (N_698,In_232,In_919);
and U699 (N_699,In_797,In_824);
xnor U700 (N_700,In_735,In_245);
and U701 (N_701,In_194,In_506);
nand U702 (N_702,In_534,In_652);
nand U703 (N_703,In_217,In_626);
and U704 (N_704,In_903,In_338);
or U705 (N_705,In_629,In_293);
nand U706 (N_706,In_854,In_624);
or U707 (N_707,In_460,In_373);
nor U708 (N_708,In_698,In_264);
and U709 (N_709,In_828,In_495);
or U710 (N_710,In_414,In_840);
and U711 (N_711,In_156,In_563);
nand U712 (N_712,In_132,In_61);
or U713 (N_713,In_157,In_744);
nand U714 (N_714,In_832,In_663);
and U715 (N_715,In_720,In_172);
and U716 (N_716,In_885,In_368);
nand U717 (N_717,In_211,In_34);
nor U718 (N_718,In_100,In_884);
or U719 (N_719,In_615,In_238);
or U720 (N_720,In_341,In_622);
nand U721 (N_721,In_863,In_332);
nand U722 (N_722,In_372,In_998);
nand U723 (N_723,In_500,In_844);
nor U724 (N_724,In_552,In_444);
nor U725 (N_725,In_323,In_760);
or U726 (N_726,In_248,In_322);
nand U727 (N_727,In_734,In_652);
and U728 (N_728,In_857,In_829);
nand U729 (N_729,In_18,In_865);
nor U730 (N_730,In_895,In_664);
nand U731 (N_731,In_89,In_55);
nor U732 (N_732,In_258,In_221);
and U733 (N_733,In_9,In_658);
nand U734 (N_734,In_279,In_736);
nor U735 (N_735,In_414,In_309);
or U736 (N_736,In_777,In_608);
or U737 (N_737,In_940,In_646);
and U738 (N_738,In_642,In_221);
nor U739 (N_739,In_455,In_246);
nor U740 (N_740,In_39,In_204);
and U741 (N_741,In_484,In_50);
nor U742 (N_742,In_391,In_962);
and U743 (N_743,In_825,In_809);
and U744 (N_744,In_191,In_509);
or U745 (N_745,In_244,In_699);
and U746 (N_746,In_637,In_143);
or U747 (N_747,In_901,In_278);
or U748 (N_748,In_483,In_60);
or U749 (N_749,In_194,In_207);
nor U750 (N_750,In_140,In_105);
or U751 (N_751,In_95,In_981);
nand U752 (N_752,In_567,In_377);
and U753 (N_753,In_204,In_476);
nand U754 (N_754,In_158,In_157);
nand U755 (N_755,In_107,In_962);
nand U756 (N_756,In_872,In_152);
xnor U757 (N_757,In_539,In_899);
nand U758 (N_758,In_280,In_821);
and U759 (N_759,In_979,In_722);
and U760 (N_760,In_499,In_30);
nand U761 (N_761,In_887,In_685);
nand U762 (N_762,In_170,In_244);
nand U763 (N_763,In_975,In_361);
nand U764 (N_764,In_740,In_744);
and U765 (N_765,In_299,In_726);
nand U766 (N_766,In_475,In_215);
or U767 (N_767,In_828,In_364);
nand U768 (N_768,In_973,In_883);
or U769 (N_769,In_847,In_817);
nor U770 (N_770,In_359,In_693);
nand U771 (N_771,In_620,In_280);
nand U772 (N_772,In_930,In_427);
nor U773 (N_773,In_934,In_80);
or U774 (N_774,In_694,In_972);
or U775 (N_775,In_504,In_307);
or U776 (N_776,In_392,In_239);
or U777 (N_777,In_145,In_281);
and U778 (N_778,In_750,In_454);
or U779 (N_779,In_428,In_264);
or U780 (N_780,In_946,In_80);
nor U781 (N_781,In_202,In_480);
and U782 (N_782,In_641,In_590);
nand U783 (N_783,In_143,In_804);
or U784 (N_784,In_316,In_509);
nand U785 (N_785,In_47,In_732);
or U786 (N_786,In_864,In_980);
nor U787 (N_787,In_116,In_785);
nand U788 (N_788,In_265,In_819);
nand U789 (N_789,In_558,In_927);
nor U790 (N_790,In_616,In_73);
nor U791 (N_791,In_309,In_634);
and U792 (N_792,In_504,In_560);
nor U793 (N_793,In_859,In_254);
nand U794 (N_794,In_860,In_831);
nor U795 (N_795,In_253,In_329);
and U796 (N_796,In_466,In_919);
or U797 (N_797,In_814,In_781);
nor U798 (N_798,In_811,In_118);
nor U799 (N_799,In_286,In_228);
and U800 (N_800,In_679,In_43);
nor U801 (N_801,In_258,In_859);
nor U802 (N_802,In_718,In_886);
nand U803 (N_803,In_652,In_111);
or U804 (N_804,In_302,In_585);
nand U805 (N_805,In_137,In_276);
and U806 (N_806,In_505,In_753);
nand U807 (N_807,In_27,In_465);
or U808 (N_808,In_73,In_469);
nor U809 (N_809,In_273,In_128);
or U810 (N_810,In_14,In_803);
or U811 (N_811,In_2,In_137);
nor U812 (N_812,In_806,In_613);
nor U813 (N_813,In_136,In_977);
and U814 (N_814,In_271,In_213);
nand U815 (N_815,In_694,In_263);
or U816 (N_816,In_467,In_575);
or U817 (N_817,In_831,In_529);
nor U818 (N_818,In_319,In_629);
and U819 (N_819,In_59,In_437);
nand U820 (N_820,In_594,In_378);
or U821 (N_821,In_249,In_206);
nand U822 (N_822,In_924,In_118);
nand U823 (N_823,In_978,In_877);
nand U824 (N_824,In_365,In_633);
nor U825 (N_825,In_325,In_712);
and U826 (N_826,In_676,In_698);
nand U827 (N_827,In_649,In_697);
or U828 (N_828,In_994,In_48);
nor U829 (N_829,In_532,In_205);
or U830 (N_830,In_884,In_430);
nor U831 (N_831,In_201,In_738);
nand U832 (N_832,In_303,In_198);
nand U833 (N_833,In_372,In_380);
and U834 (N_834,In_239,In_352);
and U835 (N_835,In_690,In_689);
nor U836 (N_836,In_563,In_16);
nor U837 (N_837,In_956,In_157);
and U838 (N_838,In_998,In_900);
nor U839 (N_839,In_831,In_208);
nor U840 (N_840,In_34,In_792);
and U841 (N_841,In_74,In_890);
or U842 (N_842,In_958,In_971);
or U843 (N_843,In_488,In_173);
or U844 (N_844,In_911,In_594);
nand U845 (N_845,In_678,In_59);
nor U846 (N_846,In_221,In_877);
nor U847 (N_847,In_30,In_496);
and U848 (N_848,In_45,In_6);
and U849 (N_849,In_777,In_877);
and U850 (N_850,In_651,In_678);
nand U851 (N_851,In_485,In_446);
or U852 (N_852,In_305,In_830);
and U853 (N_853,In_388,In_647);
nand U854 (N_854,In_98,In_968);
or U855 (N_855,In_528,In_512);
nand U856 (N_856,In_139,In_82);
and U857 (N_857,In_971,In_279);
nand U858 (N_858,In_853,In_110);
xor U859 (N_859,In_252,In_633);
or U860 (N_860,In_729,In_346);
nor U861 (N_861,In_445,In_394);
or U862 (N_862,In_954,In_565);
and U863 (N_863,In_504,In_304);
nand U864 (N_864,In_583,In_19);
or U865 (N_865,In_918,In_889);
nor U866 (N_866,In_825,In_505);
nor U867 (N_867,In_341,In_881);
and U868 (N_868,In_810,In_637);
or U869 (N_869,In_453,In_34);
and U870 (N_870,In_255,In_311);
nor U871 (N_871,In_911,In_817);
nand U872 (N_872,In_135,In_839);
nand U873 (N_873,In_909,In_139);
xnor U874 (N_874,In_872,In_489);
and U875 (N_875,In_868,In_944);
and U876 (N_876,In_312,In_368);
nand U877 (N_877,In_217,In_218);
nand U878 (N_878,In_733,In_453);
and U879 (N_879,In_462,In_860);
nand U880 (N_880,In_643,In_688);
nand U881 (N_881,In_947,In_532);
and U882 (N_882,In_211,In_557);
and U883 (N_883,In_506,In_461);
or U884 (N_884,In_286,In_84);
or U885 (N_885,In_664,In_354);
nand U886 (N_886,In_481,In_236);
nor U887 (N_887,In_7,In_305);
and U888 (N_888,In_998,In_165);
or U889 (N_889,In_107,In_850);
nand U890 (N_890,In_828,In_366);
or U891 (N_891,In_979,In_371);
nand U892 (N_892,In_595,In_640);
nand U893 (N_893,In_425,In_247);
and U894 (N_894,In_164,In_399);
nand U895 (N_895,In_32,In_415);
nand U896 (N_896,In_122,In_639);
and U897 (N_897,In_677,In_622);
and U898 (N_898,In_628,In_637);
nor U899 (N_899,In_216,In_215);
nand U900 (N_900,In_509,In_452);
nand U901 (N_901,In_853,In_811);
nor U902 (N_902,In_713,In_94);
and U903 (N_903,In_542,In_652);
or U904 (N_904,In_297,In_877);
nor U905 (N_905,In_786,In_891);
and U906 (N_906,In_818,In_132);
and U907 (N_907,In_466,In_853);
or U908 (N_908,In_790,In_224);
or U909 (N_909,In_572,In_867);
or U910 (N_910,In_256,In_98);
nor U911 (N_911,In_424,In_275);
nand U912 (N_912,In_387,In_505);
nand U913 (N_913,In_955,In_728);
nor U914 (N_914,In_801,In_654);
nor U915 (N_915,In_842,In_193);
nor U916 (N_916,In_733,In_80);
or U917 (N_917,In_379,In_184);
and U918 (N_918,In_918,In_549);
and U919 (N_919,In_951,In_278);
and U920 (N_920,In_667,In_698);
nand U921 (N_921,In_381,In_179);
and U922 (N_922,In_576,In_452);
nand U923 (N_923,In_393,In_909);
and U924 (N_924,In_935,In_210);
and U925 (N_925,In_348,In_388);
nor U926 (N_926,In_853,In_403);
nand U927 (N_927,In_139,In_903);
or U928 (N_928,In_232,In_40);
nand U929 (N_929,In_790,In_729);
nand U930 (N_930,In_437,In_62);
and U931 (N_931,In_100,In_514);
or U932 (N_932,In_416,In_183);
or U933 (N_933,In_562,In_297);
and U934 (N_934,In_323,In_15);
nand U935 (N_935,In_474,In_885);
nand U936 (N_936,In_669,In_415);
nor U937 (N_937,In_705,In_336);
and U938 (N_938,In_968,In_904);
and U939 (N_939,In_272,In_250);
and U940 (N_940,In_92,In_18);
and U941 (N_941,In_163,In_428);
and U942 (N_942,In_66,In_371);
and U943 (N_943,In_333,In_395);
and U944 (N_944,In_627,In_414);
and U945 (N_945,In_429,In_753);
and U946 (N_946,In_103,In_682);
or U947 (N_947,In_784,In_735);
or U948 (N_948,In_924,In_244);
or U949 (N_949,In_798,In_334);
nand U950 (N_950,In_99,In_829);
nor U951 (N_951,In_647,In_1);
nor U952 (N_952,In_999,In_774);
nor U953 (N_953,In_932,In_91);
and U954 (N_954,In_852,In_477);
nand U955 (N_955,In_828,In_542);
nor U956 (N_956,In_931,In_652);
and U957 (N_957,In_452,In_835);
nand U958 (N_958,In_81,In_508);
or U959 (N_959,In_720,In_105);
nor U960 (N_960,In_623,In_555);
or U961 (N_961,In_508,In_458);
and U962 (N_962,In_428,In_653);
nor U963 (N_963,In_646,In_692);
nand U964 (N_964,In_363,In_625);
or U965 (N_965,In_272,In_649);
or U966 (N_966,In_226,In_993);
nor U967 (N_967,In_47,In_303);
or U968 (N_968,In_8,In_297);
nand U969 (N_969,In_787,In_519);
nand U970 (N_970,In_916,In_619);
and U971 (N_971,In_652,In_539);
and U972 (N_972,In_246,In_302);
nand U973 (N_973,In_783,In_520);
nor U974 (N_974,In_153,In_711);
nand U975 (N_975,In_11,In_266);
or U976 (N_976,In_236,In_111);
nand U977 (N_977,In_637,In_938);
nand U978 (N_978,In_693,In_1);
and U979 (N_979,In_338,In_367);
and U980 (N_980,In_755,In_421);
nor U981 (N_981,In_432,In_898);
nand U982 (N_982,In_202,In_477);
or U983 (N_983,In_816,In_362);
or U984 (N_984,In_233,In_550);
nor U985 (N_985,In_255,In_261);
nand U986 (N_986,In_582,In_549);
and U987 (N_987,In_749,In_270);
and U988 (N_988,In_71,In_572);
nor U989 (N_989,In_946,In_117);
nor U990 (N_990,In_203,In_780);
and U991 (N_991,In_229,In_972);
and U992 (N_992,In_822,In_589);
nand U993 (N_993,In_461,In_336);
and U994 (N_994,In_875,In_675);
nand U995 (N_995,In_863,In_763);
and U996 (N_996,In_224,In_634);
nor U997 (N_997,In_322,In_796);
nor U998 (N_998,In_854,In_596);
nand U999 (N_999,In_28,In_871);
nor U1000 (N_1000,In_740,In_581);
or U1001 (N_1001,In_489,In_105);
nand U1002 (N_1002,In_320,In_650);
nor U1003 (N_1003,In_871,In_688);
nor U1004 (N_1004,In_96,In_806);
nand U1005 (N_1005,In_577,In_884);
nor U1006 (N_1006,In_374,In_692);
nand U1007 (N_1007,In_76,In_893);
nand U1008 (N_1008,In_741,In_779);
or U1009 (N_1009,In_487,In_253);
or U1010 (N_1010,In_365,In_722);
nor U1011 (N_1011,In_645,In_296);
or U1012 (N_1012,In_227,In_498);
nand U1013 (N_1013,In_781,In_829);
or U1014 (N_1014,In_430,In_84);
and U1015 (N_1015,In_73,In_542);
and U1016 (N_1016,In_623,In_169);
or U1017 (N_1017,In_613,In_300);
nand U1018 (N_1018,In_578,In_845);
or U1019 (N_1019,In_221,In_718);
and U1020 (N_1020,In_143,In_915);
and U1021 (N_1021,In_639,In_15);
or U1022 (N_1022,In_349,In_112);
nor U1023 (N_1023,In_761,In_926);
and U1024 (N_1024,In_739,In_724);
nand U1025 (N_1025,In_541,In_478);
and U1026 (N_1026,In_998,In_963);
or U1027 (N_1027,In_274,In_303);
nand U1028 (N_1028,In_107,In_652);
or U1029 (N_1029,In_311,In_237);
or U1030 (N_1030,In_613,In_372);
or U1031 (N_1031,In_774,In_361);
nand U1032 (N_1032,In_400,In_294);
or U1033 (N_1033,In_60,In_843);
nor U1034 (N_1034,In_310,In_319);
or U1035 (N_1035,In_4,In_216);
or U1036 (N_1036,In_927,In_177);
xor U1037 (N_1037,In_970,In_511);
nand U1038 (N_1038,In_18,In_238);
or U1039 (N_1039,In_15,In_739);
and U1040 (N_1040,In_941,In_417);
or U1041 (N_1041,In_649,In_326);
nand U1042 (N_1042,In_86,In_298);
nor U1043 (N_1043,In_58,In_942);
nand U1044 (N_1044,In_305,In_618);
nand U1045 (N_1045,In_621,In_222);
and U1046 (N_1046,In_894,In_156);
and U1047 (N_1047,In_851,In_646);
or U1048 (N_1048,In_645,In_654);
nand U1049 (N_1049,In_515,In_450);
xnor U1050 (N_1050,In_888,In_496);
nor U1051 (N_1051,In_615,In_245);
xnor U1052 (N_1052,In_216,In_982);
nand U1053 (N_1053,In_402,In_730);
or U1054 (N_1054,In_482,In_575);
nand U1055 (N_1055,In_464,In_973);
and U1056 (N_1056,In_811,In_986);
and U1057 (N_1057,In_358,In_335);
and U1058 (N_1058,In_811,In_641);
xor U1059 (N_1059,In_335,In_596);
nand U1060 (N_1060,In_752,In_608);
or U1061 (N_1061,In_169,In_180);
nor U1062 (N_1062,In_896,In_837);
nor U1063 (N_1063,In_519,In_252);
or U1064 (N_1064,In_918,In_790);
nand U1065 (N_1065,In_635,In_404);
nor U1066 (N_1066,In_522,In_18);
nor U1067 (N_1067,In_728,In_499);
nand U1068 (N_1068,In_694,In_229);
and U1069 (N_1069,In_696,In_964);
and U1070 (N_1070,In_150,In_262);
or U1071 (N_1071,In_73,In_40);
nor U1072 (N_1072,In_537,In_961);
or U1073 (N_1073,In_160,In_126);
nor U1074 (N_1074,In_377,In_969);
or U1075 (N_1075,In_369,In_660);
nor U1076 (N_1076,In_496,In_150);
nand U1077 (N_1077,In_2,In_332);
nand U1078 (N_1078,In_628,In_463);
nor U1079 (N_1079,In_264,In_442);
and U1080 (N_1080,In_831,In_760);
or U1081 (N_1081,In_172,In_71);
and U1082 (N_1082,In_665,In_513);
nand U1083 (N_1083,In_189,In_693);
or U1084 (N_1084,In_367,In_209);
nand U1085 (N_1085,In_1,In_890);
nand U1086 (N_1086,In_182,In_397);
or U1087 (N_1087,In_626,In_606);
nand U1088 (N_1088,In_280,In_386);
and U1089 (N_1089,In_936,In_633);
nand U1090 (N_1090,In_727,In_624);
nand U1091 (N_1091,In_383,In_89);
or U1092 (N_1092,In_569,In_204);
or U1093 (N_1093,In_462,In_116);
and U1094 (N_1094,In_138,In_802);
nor U1095 (N_1095,In_17,In_959);
nand U1096 (N_1096,In_323,In_431);
nand U1097 (N_1097,In_5,In_577);
or U1098 (N_1098,In_492,In_958);
nor U1099 (N_1099,In_541,In_954);
and U1100 (N_1100,In_167,In_104);
nor U1101 (N_1101,In_272,In_982);
nor U1102 (N_1102,In_843,In_218);
nand U1103 (N_1103,In_690,In_220);
nand U1104 (N_1104,In_626,In_207);
or U1105 (N_1105,In_233,In_934);
nor U1106 (N_1106,In_794,In_231);
nand U1107 (N_1107,In_697,In_312);
or U1108 (N_1108,In_526,In_494);
nor U1109 (N_1109,In_111,In_288);
nand U1110 (N_1110,In_243,In_688);
nand U1111 (N_1111,In_979,In_959);
and U1112 (N_1112,In_653,In_822);
nand U1113 (N_1113,In_859,In_76);
nor U1114 (N_1114,In_57,In_197);
or U1115 (N_1115,In_72,In_627);
nand U1116 (N_1116,In_797,In_709);
nor U1117 (N_1117,In_810,In_293);
nor U1118 (N_1118,In_199,In_327);
nand U1119 (N_1119,In_98,In_163);
xor U1120 (N_1120,In_241,In_904);
nand U1121 (N_1121,In_748,In_576);
nor U1122 (N_1122,In_413,In_154);
and U1123 (N_1123,In_440,In_17);
and U1124 (N_1124,In_340,In_170);
nor U1125 (N_1125,In_979,In_872);
and U1126 (N_1126,In_415,In_950);
nand U1127 (N_1127,In_113,In_805);
and U1128 (N_1128,In_79,In_161);
or U1129 (N_1129,In_654,In_268);
or U1130 (N_1130,In_177,In_3);
and U1131 (N_1131,In_39,In_21);
or U1132 (N_1132,In_229,In_570);
or U1133 (N_1133,In_259,In_665);
nor U1134 (N_1134,In_902,In_469);
nor U1135 (N_1135,In_650,In_149);
and U1136 (N_1136,In_421,In_932);
nor U1137 (N_1137,In_338,In_671);
nor U1138 (N_1138,In_193,In_615);
nand U1139 (N_1139,In_868,In_217);
nor U1140 (N_1140,In_277,In_539);
and U1141 (N_1141,In_436,In_645);
nand U1142 (N_1142,In_960,In_753);
nor U1143 (N_1143,In_585,In_516);
or U1144 (N_1144,In_472,In_791);
and U1145 (N_1145,In_906,In_465);
and U1146 (N_1146,In_882,In_715);
nand U1147 (N_1147,In_868,In_390);
and U1148 (N_1148,In_19,In_793);
nand U1149 (N_1149,In_416,In_377);
nor U1150 (N_1150,In_738,In_866);
nor U1151 (N_1151,In_613,In_566);
or U1152 (N_1152,In_459,In_663);
nand U1153 (N_1153,In_235,In_765);
nand U1154 (N_1154,In_805,In_811);
and U1155 (N_1155,In_667,In_464);
or U1156 (N_1156,In_595,In_39);
and U1157 (N_1157,In_370,In_731);
nor U1158 (N_1158,In_297,In_440);
nor U1159 (N_1159,In_677,In_890);
and U1160 (N_1160,In_629,In_141);
and U1161 (N_1161,In_333,In_989);
or U1162 (N_1162,In_47,In_787);
nand U1163 (N_1163,In_922,In_241);
nor U1164 (N_1164,In_605,In_651);
nor U1165 (N_1165,In_286,In_705);
and U1166 (N_1166,In_595,In_676);
nor U1167 (N_1167,In_138,In_975);
nor U1168 (N_1168,In_347,In_642);
and U1169 (N_1169,In_195,In_650);
nand U1170 (N_1170,In_37,In_460);
and U1171 (N_1171,In_451,In_889);
or U1172 (N_1172,In_269,In_472);
and U1173 (N_1173,In_835,In_497);
nand U1174 (N_1174,In_481,In_498);
or U1175 (N_1175,In_20,In_614);
and U1176 (N_1176,In_918,In_70);
and U1177 (N_1177,In_968,In_152);
nor U1178 (N_1178,In_984,In_207);
nor U1179 (N_1179,In_1,In_574);
nor U1180 (N_1180,In_285,In_884);
nor U1181 (N_1181,In_238,In_558);
nor U1182 (N_1182,In_17,In_573);
nand U1183 (N_1183,In_84,In_505);
nand U1184 (N_1184,In_928,In_872);
nor U1185 (N_1185,In_556,In_620);
or U1186 (N_1186,In_15,In_889);
or U1187 (N_1187,In_71,In_409);
nand U1188 (N_1188,In_983,In_507);
and U1189 (N_1189,In_861,In_838);
or U1190 (N_1190,In_687,In_760);
nor U1191 (N_1191,In_228,In_654);
nand U1192 (N_1192,In_840,In_752);
and U1193 (N_1193,In_252,In_994);
and U1194 (N_1194,In_264,In_273);
nand U1195 (N_1195,In_270,In_926);
nor U1196 (N_1196,In_859,In_505);
and U1197 (N_1197,In_492,In_798);
nand U1198 (N_1198,In_119,In_653);
nor U1199 (N_1199,In_632,In_817);
nand U1200 (N_1200,In_56,In_635);
and U1201 (N_1201,In_122,In_46);
and U1202 (N_1202,In_926,In_734);
xor U1203 (N_1203,In_812,In_962);
or U1204 (N_1204,In_230,In_17);
and U1205 (N_1205,In_223,In_382);
nand U1206 (N_1206,In_482,In_736);
nor U1207 (N_1207,In_301,In_645);
and U1208 (N_1208,In_223,In_480);
and U1209 (N_1209,In_867,In_600);
nand U1210 (N_1210,In_705,In_976);
and U1211 (N_1211,In_764,In_236);
nor U1212 (N_1212,In_975,In_747);
nand U1213 (N_1213,In_297,In_358);
nor U1214 (N_1214,In_352,In_377);
nor U1215 (N_1215,In_773,In_146);
nor U1216 (N_1216,In_301,In_693);
or U1217 (N_1217,In_209,In_107);
nor U1218 (N_1218,In_75,In_228);
nor U1219 (N_1219,In_881,In_657);
and U1220 (N_1220,In_900,In_759);
nand U1221 (N_1221,In_70,In_779);
or U1222 (N_1222,In_835,In_984);
nor U1223 (N_1223,In_402,In_255);
and U1224 (N_1224,In_547,In_702);
and U1225 (N_1225,In_343,In_432);
nand U1226 (N_1226,In_269,In_325);
or U1227 (N_1227,In_842,In_240);
and U1228 (N_1228,In_401,In_255);
nand U1229 (N_1229,In_565,In_622);
or U1230 (N_1230,In_850,In_193);
or U1231 (N_1231,In_776,In_173);
nand U1232 (N_1232,In_178,In_522);
and U1233 (N_1233,In_156,In_373);
or U1234 (N_1234,In_46,In_954);
or U1235 (N_1235,In_759,In_714);
or U1236 (N_1236,In_34,In_891);
and U1237 (N_1237,In_835,In_369);
xnor U1238 (N_1238,In_595,In_500);
or U1239 (N_1239,In_880,In_796);
or U1240 (N_1240,In_638,In_567);
nor U1241 (N_1241,In_228,In_268);
or U1242 (N_1242,In_17,In_499);
nor U1243 (N_1243,In_738,In_779);
xor U1244 (N_1244,In_461,In_812);
and U1245 (N_1245,In_195,In_755);
or U1246 (N_1246,In_196,In_688);
or U1247 (N_1247,In_463,In_868);
nand U1248 (N_1248,In_395,In_769);
and U1249 (N_1249,In_472,In_83);
nand U1250 (N_1250,In_529,In_622);
or U1251 (N_1251,In_868,In_682);
nor U1252 (N_1252,In_87,In_577);
and U1253 (N_1253,In_320,In_167);
nor U1254 (N_1254,In_827,In_586);
nor U1255 (N_1255,In_167,In_781);
nand U1256 (N_1256,In_569,In_701);
nand U1257 (N_1257,In_692,In_22);
or U1258 (N_1258,In_817,In_156);
xor U1259 (N_1259,In_905,In_597);
nor U1260 (N_1260,In_857,In_254);
and U1261 (N_1261,In_540,In_832);
or U1262 (N_1262,In_745,In_746);
or U1263 (N_1263,In_205,In_682);
or U1264 (N_1264,In_623,In_599);
or U1265 (N_1265,In_800,In_592);
nand U1266 (N_1266,In_722,In_194);
nor U1267 (N_1267,In_652,In_296);
nand U1268 (N_1268,In_707,In_208);
or U1269 (N_1269,In_410,In_259);
nand U1270 (N_1270,In_705,In_867);
or U1271 (N_1271,In_319,In_524);
and U1272 (N_1272,In_534,In_479);
or U1273 (N_1273,In_29,In_791);
and U1274 (N_1274,In_472,In_843);
nand U1275 (N_1275,In_747,In_615);
nor U1276 (N_1276,In_746,In_457);
and U1277 (N_1277,In_612,In_64);
or U1278 (N_1278,In_285,In_14);
nand U1279 (N_1279,In_733,In_719);
or U1280 (N_1280,In_546,In_245);
nor U1281 (N_1281,In_58,In_488);
nand U1282 (N_1282,In_719,In_434);
and U1283 (N_1283,In_477,In_274);
nor U1284 (N_1284,In_698,In_891);
nand U1285 (N_1285,In_44,In_850);
nand U1286 (N_1286,In_379,In_317);
nor U1287 (N_1287,In_26,In_621);
and U1288 (N_1288,In_556,In_507);
and U1289 (N_1289,In_646,In_120);
nand U1290 (N_1290,In_109,In_594);
and U1291 (N_1291,In_483,In_437);
nor U1292 (N_1292,In_66,In_267);
nor U1293 (N_1293,In_948,In_118);
and U1294 (N_1294,In_146,In_699);
or U1295 (N_1295,In_535,In_292);
and U1296 (N_1296,In_688,In_920);
nor U1297 (N_1297,In_730,In_693);
nor U1298 (N_1298,In_3,In_612);
and U1299 (N_1299,In_846,In_514);
nor U1300 (N_1300,In_546,In_437);
xnor U1301 (N_1301,In_413,In_517);
nor U1302 (N_1302,In_585,In_286);
and U1303 (N_1303,In_308,In_724);
nor U1304 (N_1304,In_80,In_655);
and U1305 (N_1305,In_992,In_814);
nand U1306 (N_1306,In_474,In_549);
nor U1307 (N_1307,In_539,In_860);
and U1308 (N_1308,In_534,In_492);
or U1309 (N_1309,In_864,In_435);
or U1310 (N_1310,In_57,In_559);
nand U1311 (N_1311,In_424,In_108);
nor U1312 (N_1312,In_253,In_912);
nand U1313 (N_1313,In_854,In_358);
nor U1314 (N_1314,In_494,In_535);
or U1315 (N_1315,In_763,In_743);
nor U1316 (N_1316,In_206,In_667);
nand U1317 (N_1317,In_933,In_78);
nand U1318 (N_1318,In_600,In_456);
and U1319 (N_1319,In_355,In_742);
or U1320 (N_1320,In_52,In_811);
or U1321 (N_1321,In_748,In_456);
and U1322 (N_1322,In_362,In_280);
nor U1323 (N_1323,In_660,In_725);
and U1324 (N_1324,In_843,In_864);
or U1325 (N_1325,In_677,In_555);
nor U1326 (N_1326,In_390,In_352);
nor U1327 (N_1327,In_769,In_512);
nand U1328 (N_1328,In_787,In_121);
nor U1329 (N_1329,In_767,In_528);
nand U1330 (N_1330,In_788,In_309);
nand U1331 (N_1331,In_627,In_321);
and U1332 (N_1332,In_105,In_672);
and U1333 (N_1333,In_719,In_646);
nand U1334 (N_1334,In_371,In_118);
and U1335 (N_1335,In_702,In_173);
or U1336 (N_1336,In_238,In_25);
nand U1337 (N_1337,In_345,In_81);
nand U1338 (N_1338,In_590,In_764);
nand U1339 (N_1339,In_607,In_889);
or U1340 (N_1340,In_572,In_20);
nor U1341 (N_1341,In_588,In_367);
nor U1342 (N_1342,In_904,In_120);
nand U1343 (N_1343,In_432,In_942);
or U1344 (N_1344,In_614,In_778);
or U1345 (N_1345,In_280,In_248);
and U1346 (N_1346,In_836,In_81);
or U1347 (N_1347,In_471,In_568);
and U1348 (N_1348,In_286,In_877);
nor U1349 (N_1349,In_858,In_146);
nand U1350 (N_1350,In_345,In_348);
or U1351 (N_1351,In_136,In_941);
and U1352 (N_1352,In_770,In_535);
xor U1353 (N_1353,In_961,In_158);
nor U1354 (N_1354,In_578,In_423);
nor U1355 (N_1355,In_450,In_257);
and U1356 (N_1356,In_974,In_137);
nor U1357 (N_1357,In_478,In_330);
and U1358 (N_1358,In_154,In_174);
and U1359 (N_1359,In_149,In_933);
and U1360 (N_1360,In_431,In_321);
or U1361 (N_1361,In_591,In_663);
and U1362 (N_1362,In_231,In_431);
or U1363 (N_1363,In_49,In_191);
nor U1364 (N_1364,In_907,In_537);
nor U1365 (N_1365,In_624,In_62);
nor U1366 (N_1366,In_358,In_715);
nor U1367 (N_1367,In_793,In_528);
or U1368 (N_1368,In_272,In_436);
and U1369 (N_1369,In_356,In_58);
xnor U1370 (N_1370,In_3,In_443);
nor U1371 (N_1371,In_901,In_191);
nor U1372 (N_1372,In_993,In_295);
or U1373 (N_1373,In_986,In_168);
and U1374 (N_1374,In_949,In_666);
or U1375 (N_1375,In_5,In_109);
or U1376 (N_1376,In_5,In_311);
and U1377 (N_1377,In_952,In_793);
nand U1378 (N_1378,In_380,In_920);
or U1379 (N_1379,In_804,In_919);
nor U1380 (N_1380,In_765,In_270);
nand U1381 (N_1381,In_571,In_979);
and U1382 (N_1382,In_815,In_565);
nor U1383 (N_1383,In_947,In_802);
nand U1384 (N_1384,In_406,In_613);
nand U1385 (N_1385,In_917,In_694);
nand U1386 (N_1386,In_663,In_621);
and U1387 (N_1387,In_802,In_975);
and U1388 (N_1388,In_128,In_969);
or U1389 (N_1389,In_386,In_48);
and U1390 (N_1390,In_352,In_738);
and U1391 (N_1391,In_444,In_637);
and U1392 (N_1392,In_442,In_249);
nand U1393 (N_1393,In_925,In_812);
nor U1394 (N_1394,In_864,In_765);
nand U1395 (N_1395,In_140,In_35);
or U1396 (N_1396,In_257,In_547);
nand U1397 (N_1397,In_400,In_589);
nor U1398 (N_1398,In_27,In_30);
or U1399 (N_1399,In_678,In_578);
nand U1400 (N_1400,In_952,In_113);
nand U1401 (N_1401,In_914,In_66);
or U1402 (N_1402,In_688,In_33);
nor U1403 (N_1403,In_135,In_696);
nor U1404 (N_1404,In_146,In_289);
nand U1405 (N_1405,In_688,In_745);
and U1406 (N_1406,In_29,In_27);
nor U1407 (N_1407,In_672,In_993);
and U1408 (N_1408,In_287,In_556);
nand U1409 (N_1409,In_119,In_962);
nor U1410 (N_1410,In_33,In_749);
nor U1411 (N_1411,In_679,In_762);
nor U1412 (N_1412,In_192,In_180);
nor U1413 (N_1413,In_803,In_960);
or U1414 (N_1414,In_658,In_525);
nand U1415 (N_1415,In_324,In_262);
or U1416 (N_1416,In_877,In_236);
nor U1417 (N_1417,In_718,In_361);
and U1418 (N_1418,In_1,In_430);
and U1419 (N_1419,In_667,In_241);
nor U1420 (N_1420,In_520,In_223);
or U1421 (N_1421,In_405,In_969);
and U1422 (N_1422,In_100,In_40);
nand U1423 (N_1423,In_221,In_497);
and U1424 (N_1424,In_209,In_227);
and U1425 (N_1425,In_59,In_494);
or U1426 (N_1426,In_447,In_516);
and U1427 (N_1427,In_521,In_38);
or U1428 (N_1428,In_63,In_994);
nand U1429 (N_1429,In_638,In_73);
nor U1430 (N_1430,In_729,In_532);
nand U1431 (N_1431,In_63,In_532);
or U1432 (N_1432,In_428,In_6);
nand U1433 (N_1433,In_743,In_572);
and U1434 (N_1434,In_271,In_415);
nor U1435 (N_1435,In_820,In_338);
and U1436 (N_1436,In_769,In_870);
nand U1437 (N_1437,In_884,In_307);
or U1438 (N_1438,In_695,In_108);
or U1439 (N_1439,In_769,In_117);
or U1440 (N_1440,In_118,In_454);
or U1441 (N_1441,In_407,In_454);
nor U1442 (N_1442,In_920,In_370);
or U1443 (N_1443,In_770,In_958);
or U1444 (N_1444,In_216,In_780);
or U1445 (N_1445,In_960,In_974);
nor U1446 (N_1446,In_940,In_337);
and U1447 (N_1447,In_355,In_114);
or U1448 (N_1448,In_399,In_661);
nor U1449 (N_1449,In_675,In_734);
or U1450 (N_1450,In_998,In_277);
nor U1451 (N_1451,In_466,In_459);
xnor U1452 (N_1452,In_384,In_693);
nor U1453 (N_1453,In_382,In_422);
xnor U1454 (N_1454,In_5,In_65);
nor U1455 (N_1455,In_884,In_164);
nand U1456 (N_1456,In_804,In_29);
nor U1457 (N_1457,In_532,In_293);
and U1458 (N_1458,In_657,In_298);
nand U1459 (N_1459,In_884,In_318);
nor U1460 (N_1460,In_332,In_92);
or U1461 (N_1461,In_952,In_221);
nand U1462 (N_1462,In_580,In_150);
nand U1463 (N_1463,In_446,In_613);
and U1464 (N_1464,In_193,In_36);
nor U1465 (N_1465,In_619,In_450);
xnor U1466 (N_1466,In_729,In_737);
nor U1467 (N_1467,In_698,In_116);
nor U1468 (N_1468,In_976,In_165);
nor U1469 (N_1469,In_449,In_112);
nand U1470 (N_1470,In_307,In_196);
nor U1471 (N_1471,In_587,In_180);
nand U1472 (N_1472,In_304,In_781);
or U1473 (N_1473,In_97,In_368);
or U1474 (N_1474,In_485,In_162);
nor U1475 (N_1475,In_624,In_343);
nand U1476 (N_1476,In_719,In_743);
or U1477 (N_1477,In_898,In_604);
and U1478 (N_1478,In_849,In_672);
xor U1479 (N_1479,In_382,In_786);
nor U1480 (N_1480,In_863,In_970);
nand U1481 (N_1481,In_491,In_525);
nand U1482 (N_1482,In_163,In_197);
and U1483 (N_1483,In_256,In_748);
and U1484 (N_1484,In_723,In_755);
nand U1485 (N_1485,In_532,In_997);
nand U1486 (N_1486,In_954,In_771);
xor U1487 (N_1487,In_317,In_779);
or U1488 (N_1488,In_736,In_519);
or U1489 (N_1489,In_880,In_671);
nor U1490 (N_1490,In_626,In_990);
and U1491 (N_1491,In_652,In_928);
or U1492 (N_1492,In_175,In_202);
and U1493 (N_1493,In_578,In_267);
nor U1494 (N_1494,In_602,In_475);
nor U1495 (N_1495,In_408,In_345);
and U1496 (N_1496,In_493,In_66);
nand U1497 (N_1497,In_921,In_29);
and U1498 (N_1498,In_381,In_209);
or U1499 (N_1499,In_775,In_656);
and U1500 (N_1500,In_952,In_790);
nand U1501 (N_1501,In_833,In_664);
nand U1502 (N_1502,In_239,In_869);
and U1503 (N_1503,In_477,In_721);
and U1504 (N_1504,In_715,In_447);
nand U1505 (N_1505,In_541,In_313);
and U1506 (N_1506,In_977,In_5);
and U1507 (N_1507,In_727,In_655);
nor U1508 (N_1508,In_337,In_249);
nand U1509 (N_1509,In_257,In_264);
nand U1510 (N_1510,In_466,In_494);
and U1511 (N_1511,In_190,In_471);
or U1512 (N_1512,In_334,In_753);
or U1513 (N_1513,In_856,In_308);
or U1514 (N_1514,In_714,In_539);
nor U1515 (N_1515,In_351,In_49);
nor U1516 (N_1516,In_969,In_268);
nand U1517 (N_1517,In_79,In_289);
or U1518 (N_1518,In_645,In_232);
and U1519 (N_1519,In_872,In_697);
nor U1520 (N_1520,In_44,In_18);
nor U1521 (N_1521,In_584,In_321);
and U1522 (N_1522,In_588,In_123);
nand U1523 (N_1523,In_986,In_385);
and U1524 (N_1524,In_863,In_273);
and U1525 (N_1525,In_893,In_977);
nand U1526 (N_1526,In_740,In_677);
nor U1527 (N_1527,In_737,In_577);
nand U1528 (N_1528,In_659,In_504);
nand U1529 (N_1529,In_127,In_753);
and U1530 (N_1530,In_888,In_991);
or U1531 (N_1531,In_531,In_124);
nand U1532 (N_1532,In_413,In_629);
or U1533 (N_1533,In_681,In_903);
or U1534 (N_1534,In_825,In_146);
or U1535 (N_1535,In_488,In_831);
nor U1536 (N_1536,In_176,In_504);
and U1537 (N_1537,In_581,In_36);
and U1538 (N_1538,In_900,In_663);
nand U1539 (N_1539,In_938,In_667);
and U1540 (N_1540,In_504,In_239);
nand U1541 (N_1541,In_765,In_260);
nand U1542 (N_1542,In_173,In_161);
nor U1543 (N_1543,In_529,In_996);
xnor U1544 (N_1544,In_669,In_381);
nand U1545 (N_1545,In_689,In_574);
and U1546 (N_1546,In_89,In_646);
and U1547 (N_1547,In_13,In_745);
or U1548 (N_1548,In_728,In_517);
or U1549 (N_1549,In_244,In_177);
and U1550 (N_1550,In_606,In_466);
or U1551 (N_1551,In_490,In_292);
nand U1552 (N_1552,In_475,In_525);
nand U1553 (N_1553,In_138,In_108);
nor U1554 (N_1554,In_994,In_293);
and U1555 (N_1555,In_291,In_237);
and U1556 (N_1556,In_871,In_815);
or U1557 (N_1557,In_498,In_624);
nor U1558 (N_1558,In_152,In_385);
and U1559 (N_1559,In_57,In_143);
and U1560 (N_1560,In_138,In_340);
nor U1561 (N_1561,In_627,In_432);
xor U1562 (N_1562,In_620,In_902);
nand U1563 (N_1563,In_773,In_697);
nor U1564 (N_1564,In_184,In_176);
and U1565 (N_1565,In_324,In_92);
nand U1566 (N_1566,In_725,In_548);
or U1567 (N_1567,In_451,In_685);
nor U1568 (N_1568,In_873,In_622);
nand U1569 (N_1569,In_846,In_156);
or U1570 (N_1570,In_909,In_18);
nor U1571 (N_1571,In_950,In_681);
nor U1572 (N_1572,In_945,In_563);
nor U1573 (N_1573,In_341,In_187);
or U1574 (N_1574,In_914,In_6);
nor U1575 (N_1575,In_17,In_108);
nor U1576 (N_1576,In_668,In_83);
or U1577 (N_1577,In_618,In_454);
nand U1578 (N_1578,In_693,In_833);
and U1579 (N_1579,In_672,In_744);
nor U1580 (N_1580,In_723,In_689);
nand U1581 (N_1581,In_0,In_817);
nand U1582 (N_1582,In_364,In_601);
nor U1583 (N_1583,In_446,In_450);
nand U1584 (N_1584,In_993,In_249);
and U1585 (N_1585,In_466,In_660);
and U1586 (N_1586,In_162,In_773);
or U1587 (N_1587,In_617,In_161);
nor U1588 (N_1588,In_926,In_698);
nor U1589 (N_1589,In_466,In_417);
nand U1590 (N_1590,In_962,In_531);
and U1591 (N_1591,In_697,In_758);
nand U1592 (N_1592,In_191,In_918);
or U1593 (N_1593,In_525,In_439);
and U1594 (N_1594,In_187,In_980);
or U1595 (N_1595,In_769,In_982);
nand U1596 (N_1596,In_736,In_504);
or U1597 (N_1597,In_785,In_960);
nor U1598 (N_1598,In_814,In_591);
nand U1599 (N_1599,In_961,In_241);
nor U1600 (N_1600,In_198,In_844);
nor U1601 (N_1601,In_28,In_599);
nor U1602 (N_1602,In_888,In_460);
nor U1603 (N_1603,In_804,In_365);
nand U1604 (N_1604,In_51,In_240);
and U1605 (N_1605,In_626,In_655);
and U1606 (N_1606,In_723,In_157);
nor U1607 (N_1607,In_986,In_445);
or U1608 (N_1608,In_861,In_206);
and U1609 (N_1609,In_657,In_271);
and U1610 (N_1610,In_940,In_63);
nor U1611 (N_1611,In_502,In_737);
nand U1612 (N_1612,In_343,In_439);
nand U1613 (N_1613,In_36,In_598);
nor U1614 (N_1614,In_933,In_507);
and U1615 (N_1615,In_989,In_589);
nand U1616 (N_1616,In_226,In_18);
and U1617 (N_1617,In_201,In_368);
and U1618 (N_1618,In_125,In_179);
nand U1619 (N_1619,In_180,In_193);
nor U1620 (N_1620,In_470,In_329);
or U1621 (N_1621,In_566,In_393);
nand U1622 (N_1622,In_365,In_706);
or U1623 (N_1623,In_35,In_251);
nand U1624 (N_1624,In_802,In_581);
and U1625 (N_1625,In_550,In_147);
nor U1626 (N_1626,In_56,In_681);
and U1627 (N_1627,In_345,In_339);
nand U1628 (N_1628,In_908,In_600);
or U1629 (N_1629,In_771,In_145);
or U1630 (N_1630,In_219,In_440);
nand U1631 (N_1631,In_293,In_342);
nand U1632 (N_1632,In_952,In_6);
and U1633 (N_1633,In_846,In_682);
nor U1634 (N_1634,In_158,In_156);
or U1635 (N_1635,In_448,In_804);
nand U1636 (N_1636,In_657,In_306);
or U1637 (N_1637,In_929,In_643);
or U1638 (N_1638,In_493,In_635);
and U1639 (N_1639,In_661,In_836);
nand U1640 (N_1640,In_182,In_502);
nand U1641 (N_1641,In_661,In_796);
nand U1642 (N_1642,In_931,In_342);
nor U1643 (N_1643,In_745,In_637);
nand U1644 (N_1644,In_901,In_119);
or U1645 (N_1645,In_997,In_867);
and U1646 (N_1646,In_245,In_79);
or U1647 (N_1647,In_68,In_199);
nor U1648 (N_1648,In_834,In_267);
or U1649 (N_1649,In_683,In_587);
nor U1650 (N_1650,In_872,In_97);
nor U1651 (N_1651,In_352,In_815);
nand U1652 (N_1652,In_718,In_122);
nand U1653 (N_1653,In_427,In_226);
or U1654 (N_1654,In_112,In_497);
or U1655 (N_1655,In_746,In_256);
nand U1656 (N_1656,In_772,In_566);
nor U1657 (N_1657,In_733,In_129);
nor U1658 (N_1658,In_828,In_392);
nor U1659 (N_1659,In_373,In_767);
and U1660 (N_1660,In_67,In_261);
nand U1661 (N_1661,In_866,In_386);
or U1662 (N_1662,In_793,In_459);
nor U1663 (N_1663,In_350,In_559);
nand U1664 (N_1664,In_861,In_520);
nor U1665 (N_1665,In_706,In_490);
or U1666 (N_1666,In_423,In_897);
xor U1667 (N_1667,In_608,In_590);
or U1668 (N_1668,In_241,In_371);
and U1669 (N_1669,In_146,In_654);
nand U1670 (N_1670,In_466,In_560);
nor U1671 (N_1671,In_536,In_917);
nor U1672 (N_1672,In_66,In_645);
and U1673 (N_1673,In_763,In_566);
nand U1674 (N_1674,In_685,In_340);
nand U1675 (N_1675,In_474,In_56);
nor U1676 (N_1676,In_433,In_106);
nor U1677 (N_1677,In_528,In_634);
nand U1678 (N_1678,In_816,In_648);
or U1679 (N_1679,In_502,In_284);
nand U1680 (N_1680,In_980,In_375);
or U1681 (N_1681,In_315,In_297);
and U1682 (N_1682,In_591,In_450);
or U1683 (N_1683,In_267,In_686);
nand U1684 (N_1684,In_323,In_137);
and U1685 (N_1685,In_324,In_809);
nand U1686 (N_1686,In_13,In_599);
nor U1687 (N_1687,In_829,In_915);
and U1688 (N_1688,In_831,In_44);
nand U1689 (N_1689,In_811,In_752);
and U1690 (N_1690,In_345,In_413);
nor U1691 (N_1691,In_971,In_730);
or U1692 (N_1692,In_103,In_608);
or U1693 (N_1693,In_12,In_920);
nor U1694 (N_1694,In_553,In_673);
nand U1695 (N_1695,In_581,In_955);
and U1696 (N_1696,In_426,In_115);
or U1697 (N_1697,In_324,In_284);
nand U1698 (N_1698,In_208,In_604);
or U1699 (N_1699,In_720,In_623);
nor U1700 (N_1700,In_87,In_589);
nand U1701 (N_1701,In_567,In_496);
nand U1702 (N_1702,In_391,In_61);
nor U1703 (N_1703,In_3,In_969);
nor U1704 (N_1704,In_726,In_543);
nor U1705 (N_1705,In_498,In_232);
or U1706 (N_1706,In_533,In_204);
nand U1707 (N_1707,In_542,In_971);
or U1708 (N_1708,In_997,In_748);
nor U1709 (N_1709,In_938,In_858);
nand U1710 (N_1710,In_696,In_528);
and U1711 (N_1711,In_681,In_381);
nor U1712 (N_1712,In_252,In_121);
nor U1713 (N_1713,In_243,In_979);
nor U1714 (N_1714,In_804,In_730);
nor U1715 (N_1715,In_209,In_232);
nand U1716 (N_1716,In_809,In_751);
or U1717 (N_1717,In_576,In_534);
nor U1718 (N_1718,In_883,In_404);
or U1719 (N_1719,In_713,In_821);
nand U1720 (N_1720,In_577,In_985);
nand U1721 (N_1721,In_142,In_379);
nor U1722 (N_1722,In_323,In_295);
or U1723 (N_1723,In_605,In_391);
nor U1724 (N_1724,In_346,In_858);
nand U1725 (N_1725,In_272,In_61);
or U1726 (N_1726,In_292,In_914);
nand U1727 (N_1727,In_88,In_756);
and U1728 (N_1728,In_617,In_446);
or U1729 (N_1729,In_521,In_985);
or U1730 (N_1730,In_694,In_383);
or U1731 (N_1731,In_813,In_452);
nand U1732 (N_1732,In_405,In_83);
nor U1733 (N_1733,In_602,In_806);
nand U1734 (N_1734,In_388,In_765);
or U1735 (N_1735,In_968,In_674);
and U1736 (N_1736,In_126,In_288);
nor U1737 (N_1737,In_533,In_738);
nand U1738 (N_1738,In_593,In_386);
nor U1739 (N_1739,In_669,In_617);
or U1740 (N_1740,In_987,In_593);
and U1741 (N_1741,In_120,In_549);
or U1742 (N_1742,In_283,In_23);
and U1743 (N_1743,In_616,In_771);
nor U1744 (N_1744,In_635,In_23);
and U1745 (N_1745,In_280,In_927);
and U1746 (N_1746,In_357,In_522);
and U1747 (N_1747,In_977,In_194);
nor U1748 (N_1748,In_374,In_95);
and U1749 (N_1749,In_959,In_493);
or U1750 (N_1750,In_779,In_183);
and U1751 (N_1751,In_39,In_547);
nor U1752 (N_1752,In_885,In_427);
or U1753 (N_1753,In_22,In_512);
nor U1754 (N_1754,In_652,In_88);
and U1755 (N_1755,In_564,In_559);
nand U1756 (N_1756,In_340,In_350);
and U1757 (N_1757,In_294,In_587);
nor U1758 (N_1758,In_572,In_773);
nor U1759 (N_1759,In_62,In_363);
nor U1760 (N_1760,In_505,In_449);
and U1761 (N_1761,In_222,In_608);
and U1762 (N_1762,In_72,In_839);
nor U1763 (N_1763,In_607,In_995);
and U1764 (N_1764,In_623,In_343);
or U1765 (N_1765,In_579,In_165);
nor U1766 (N_1766,In_838,In_651);
nand U1767 (N_1767,In_934,In_984);
nor U1768 (N_1768,In_801,In_778);
nor U1769 (N_1769,In_153,In_694);
and U1770 (N_1770,In_19,In_976);
or U1771 (N_1771,In_633,In_350);
or U1772 (N_1772,In_638,In_475);
and U1773 (N_1773,In_32,In_470);
nand U1774 (N_1774,In_670,In_105);
nor U1775 (N_1775,In_990,In_605);
and U1776 (N_1776,In_246,In_117);
nor U1777 (N_1777,In_441,In_661);
nor U1778 (N_1778,In_13,In_258);
nor U1779 (N_1779,In_607,In_327);
nor U1780 (N_1780,In_912,In_3);
nor U1781 (N_1781,In_204,In_45);
nor U1782 (N_1782,In_481,In_640);
nor U1783 (N_1783,In_267,In_586);
nor U1784 (N_1784,In_632,In_102);
and U1785 (N_1785,In_493,In_17);
nor U1786 (N_1786,In_393,In_760);
and U1787 (N_1787,In_650,In_704);
nand U1788 (N_1788,In_435,In_510);
nor U1789 (N_1789,In_9,In_836);
nor U1790 (N_1790,In_758,In_112);
nand U1791 (N_1791,In_473,In_435);
and U1792 (N_1792,In_863,In_874);
nor U1793 (N_1793,In_787,In_414);
or U1794 (N_1794,In_510,In_125);
nor U1795 (N_1795,In_703,In_695);
and U1796 (N_1796,In_965,In_996);
or U1797 (N_1797,In_665,In_847);
and U1798 (N_1798,In_395,In_352);
nor U1799 (N_1799,In_187,In_67);
nand U1800 (N_1800,In_123,In_859);
nor U1801 (N_1801,In_613,In_951);
and U1802 (N_1802,In_719,In_406);
and U1803 (N_1803,In_207,In_680);
nor U1804 (N_1804,In_693,In_672);
nor U1805 (N_1805,In_757,In_651);
and U1806 (N_1806,In_890,In_898);
or U1807 (N_1807,In_568,In_840);
nand U1808 (N_1808,In_294,In_232);
or U1809 (N_1809,In_423,In_942);
xor U1810 (N_1810,In_664,In_821);
nor U1811 (N_1811,In_972,In_437);
or U1812 (N_1812,In_893,In_884);
or U1813 (N_1813,In_113,In_603);
nand U1814 (N_1814,In_265,In_227);
or U1815 (N_1815,In_465,In_398);
nand U1816 (N_1816,In_309,In_286);
nand U1817 (N_1817,In_715,In_232);
or U1818 (N_1818,In_880,In_56);
nand U1819 (N_1819,In_25,In_829);
nand U1820 (N_1820,In_649,In_316);
nor U1821 (N_1821,In_228,In_660);
or U1822 (N_1822,In_89,In_895);
nor U1823 (N_1823,In_954,In_731);
nor U1824 (N_1824,In_707,In_186);
nand U1825 (N_1825,In_905,In_701);
nor U1826 (N_1826,In_250,In_890);
nand U1827 (N_1827,In_335,In_480);
or U1828 (N_1828,In_582,In_627);
nand U1829 (N_1829,In_128,In_60);
nor U1830 (N_1830,In_699,In_530);
nand U1831 (N_1831,In_505,In_950);
or U1832 (N_1832,In_595,In_335);
and U1833 (N_1833,In_435,In_680);
nand U1834 (N_1834,In_894,In_274);
nor U1835 (N_1835,In_305,In_411);
and U1836 (N_1836,In_685,In_535);
or U1837 (N_1837,In_413,In_321);
nand U1838 (N_1838,In_947,In_54);
xor U1839 (N_1839,In_974,In_844);
nor U1840 (N_1840,In_977,In_106);
and U1841 (N_1841,In_135,In_111);
nor U1842 (N_1842,In_830,In_26);
nand U1843 (N_1843,In_301,In_360);
xnor U1844 (N_1844,In_674,In_904);
nor U1845 (N_1845,In_803,In_329);
or U1846 (N_1846,In_560,In_809);
or U1847 (N_1847,In_213,In_33);
or U1848 (N_1848,In_119,In_862);
nand U1849 (N_1849,In_266,In_237);
nand U1850 (N_1850,In_194,In_769);
or U1851 (N_1851,In_623,In_183);
nor U1852 (N_1852,In_461,In_436);
or U1853 (N_1853,In_318,In_866);
nor U1854 (N_1854,In_961,In_843);
and U1855 (N_1855,In_27,In_44);
nor U1856 (N_1856,In_16,In_642);
and U1857 (N_1857,In_597,In_918);
nand U1858 (N_1858,In_848,In_706);
and U1859 (N_1859,In_821,In_199);
or U1860 (N_1860,In_900,In_335);
or U1861 (N_1861,In_424,In_629);
nor U1862 (N_1862,In_8,In_9);
nand U1863 (N_1863,In_264,In_422);
or U1864 (N_1864,In_498,In_614);
nand U1865 (N_1865,In_195,In_607);
nor U1866 (N_1866,In_537,In_290);
and U1867 (N_1867,In_668,In_970);
or U1868 (N_1868,In_784,In_696);
nand U1869 (N_1869,In_427,In_991);
nor U1870 (N_1870,In_114,In_704);
nor U1871 (N_1871,In_382,In_812);
and U1872 (N_1872,In_767,In_119);
nand U1873 (N_1873,In_361,In_197);
and U1874 (N_1874,In_930,In_920);
or U1875 (N_1875,In_448,In_750);
or U1876 (N_1876,In_779,In_113);
nand U1877 (N_1877,In_140,In_502);
nor U1878 (N_1878,In_95,In_895);
nand U1879 (N_1879,In_316,In_288);
or U1880 (N_1880,In_24,In_384);
nand U1881 (N_1881,In_707,In_351);
nand U1882 (N_1882,In_579,In_183);
nand U1883 (N_1883,In_797,In_762);
xnor U1884 (N_1884,In_500,In_307);
and U1885 (N_1885,In_900,In_720);
nor U1886 (N_1886,In_900,In_979);
nor U1887 (N_1887,In_217,In_294);
nand U1888 (N_1888,In_937,In_204);
nand U1889 (N_1889,In_333,In_368);
nor U1890 (N_1890,In_224,In_484);
nor U1891 (N_1891,In_307,In_905);
and U1892 (N_1892,In_268,In_711);
and U1893 (N_1893,In_729,In_579);
nor U1894 (N_1894,In_398,In_487);
nand U1895 (N_1895,In_728,In_652);
or U1896 (N_1896,In_727,In_82);
nand U1897 (N_1897,In_439,In_75);
or U1898 (N_1898,In_695,In_901);
and U1899 (N_1899,In_302,In_78);
or U1900 (N_1900,In_462,In_613);
nand U1901 (N_1901,In_709,In_974);
and U1902 (N_1902,In_167,In_731);
nand U1903 (N_1903,In_277,In_186);
nand U1904 (N_1904,In_243,In_731);
and U1905 (N_1905,In_873,In_907);
and U1906 (N_1906,In_623,In_300);
and U1907 (N_1907,In_772,In_924);
or U1908 (N_1908,In_524,In_614);
nand U1909 (N_1909,In_849,In_364);
nor U1910 (N_1910,In_974,In_24);
nand U1911 (N_1911,In_927,In_198);
or U1912 (N_1912,In_340,In_919);
or U1913 (N_1913,In_805,In_35);
xnor U1914 (N_1914,In_359,In_438);
and U1915 (N_1915,In_923,In_260);
and U1916 (N_1916,In_564,In_145);
nor U1917 (N_1917,In_757,In_586);
nand U1918 (N_1918,In_618,In_56);
and U1919 (N_1919,In_865,In_344);
nor U1920 (N_1920,In_597,In_151);
nand U1921 (N_1921,In_194,In_403);
or U1922 (N_1922,In_223,In_245);
or U1923 (N_1923,In_610,In_132);
or U1924 (N_1924,In_34,In_202);
and U1925 (N_1925,In_433,In_677);
nand U1926 (N_1926,In_698,In_855);
nor U1927 (N_1927,In_569,In_48);
or U1928 (N_1928,In_51,In_793);
nand U1929 (N_1929,In_172,In_972);
nand U1930 (N_1930,In_805,In_40);
nor U1931 (N_1931,In_623,In_613);
nor U1932 (N_1932,In_939,In_680);
nand U1933 (N_1933,In_345,In_218);
or U1934 (N_1934,In_147,In_242);
nand U1935 (N_1935,In_562,In_265);
nor U1936 (N_1936,In_420,In_275);
nand U1937 (N_1937,In_559,In_260);
xnor U1938 (N_1938,In_136,In_540);
and U1939 (N_1939,In_629,In_233);
or U1940 (N_1940,In_16,In_852);
nor U1941 (N_1941,In_160,In_549);
and U1942 (N_1942,In_284,In_803);
and U1943 (N_1943,In_988,In_395);
or U1944 (N_1944,In_328,In_780);
nand U1945 (N_1945,In_138,In_770);
nand U1946 (N_1946,In_350,In_260);
nor U1947 (N_1947,In_678,In_137);
and U1948 (N_1948,In_208,In_898);
or U1949 (N_1949,In_217,In_347);
nor U1950 (N_1950,In_178,In_140);
xor U1951 (N_1951,In_806,In_221);
or U1952 (N_1952,In_382,In_600);
or U1953 (N_1953,In_124,In_190);
and U1954 (N_1954,In_970,In_394);
or U1955 (N_1955,In_498,In_103);
nand U1956 (N_1956,In_760,In_801);
and U1957 (N_1957,In_639,In_473);
and U1958 (N_1958,In_870,In_707);
nor U1959 (N_1959,In_389,In_197);
or U1960 (N_1960,In_716,In_562);
or U1961 (N_1961,In_835,In_803);
xnor U1962 (N_1962,In_839,In_701);
nor U1963 (N_1963,In_949,In_914);
nor U1964 (N_1964,In_817,In_725);
or U1965 (N_1965,In_628,In_521);
nand U1966 (N_1966,In_545,In_613);
or U1967 (N_1967,In_775,In_226);
and U1968 (N_1968,In_280,In_837);
or U1969 (N_1969,In_343,In_200);
nand U1970 (N_1970,In_902,In_725);
nand U1971 (N_1971,In_399,In_514);
nand U1972 (N_1972,In_339,In_489);
and U1973 (N_1973,In_513,In_286);
and U1974 (N_1974,In_546,In_96);
and U1975 (N_1975,In_765,In_858);
nor U1976 (N_1976,In_811,In_793);
nand U1977 (N_1977,In_713,In_546);
or U1978 (N_1978,In_122,In_371);
nand U1979 (N_1979,In_984,In_749);
or U1980 (N_1980,In_920,In_975);
and U1981 (N_1981,In_507,In_51);
and U1982 (N_1982,In_884,In_317);
and U1983 (N_1983,In_505,In_104);
and U1984 (N_1984,In_201,In_520);
or U1985 (N_1985,In_283,In_287);
and U1986 (N_1986,In_299,In_575);
nand U1987 (N_1987,In_760,In_696);
nor U1988 (N_1988,In_193,In_242);
nand U1989 (N_1989,In_6,In_567);
and U1990 (N_1990,In_118,In_571);
nand U1991 (N_1991,In_733,In_551);
or U1992 (N_1992,In_912,In_190);
and U1993 (N_1993,In_906,In_80);
and U1994 (N_1994,In_859,In_428);
or U1995 (N_1995,In_566,In_685);
nand U1996 (N_1996,In_842,In_450);
nor U1997 (N_1997,In_954,In_447);
nand U1998 (N_1998,In_796,In_558);
and U1999 (N_1999,In_916,In_903);
nor U2000 (N_2000,In_479,In_818);
nor U2001 (N_2001,In_810,In_743);
or U2002 (N_2002,In_471,In_707);
nor U2003 (N_2003,In_904,In_375);
and U2004 (N_2004,In_459,In_756);
or U2005 (N_2005,In_246,In_448);
or U2006 (N_2006,In_303,In_331);
nor U2007 (N_2007,In_1,In_728);
nand U2008 (N_2008,In_456,In_955);
nand U2009 (N_2009,In_869,In_749);
nor U2010 (N_2010,In_804,In_960);
nor U2011 (N_2011,In_967,In_21);
nand U2012 (N_2012,In_74,In_765);
nor U2013 (N_2013,In_262,In_170);
and U2014 (N_2014,In_295,In_259);
and U2015 (N_2015,In_269,In_656);
nor U2016 (N_2016,In_237,In_684);
and U2017 (N_2017,In_667,In_134);
and U2018 (N_2018,In_39,In_479);
nand U2019 (N_2019,In_606,In_208);
nor U2020 (N_2020,In_771,In_604);
nor U2021 (N_2021,In_5,In_278);
nand U2022 (N_2022,In_442,In_404);
nor U2023 (N_2023,In_598,In_987);
nor U2024 (N_2024,In_794,In_559);
nor U2025 (N_2025,In_611,In_174);
nor U2026 (N_2026,In_900,In_429);
or U2027 (N_2027,In_582,In_79);
nand U2028 (N_2028,In_965,In_746);
nand U2029 (N_2029,In_340,In_513);
or U2030 (N_2030,In_892,In_28);
or U2031 (N_2031,In_468,In_492);
nor U2032 (N_2032,In_410,In_447);
nand U2033 (N_2033,In_96,In_1);
or U2034 (N_2034,In_856,In_780);
nor U2035 (N_2035,In_301,In_840);
nor U2036 (N_2036,In_296,In_672);
and U2037 (N_2037,In_931,In_5);
or U2038 (N_2038,In_971,In_614);
nor U2039 (N_2039,In_437,In_497);
nand U2040 (N_2040,In_351,In_766);
and U2041 (N_2041,In_274,In_931);
or U2042 (N_2042,In_378,In_881);
and U2043 (N_2043,In_248,In_752);
nor U2044 (N_2044,In_164,In_882);
and U2045 (N_2045,In_965,In_751);
nor U2046 (N_2046,In_209,In_496);
and U2047 (N_2047,In_573,In_356);
nor U2048 (N_2048,In_432,In_977);
nand U2049 (N_2049,In_80,In_897);
nand U2050 (N_2050,In_980,In_312);
and U2051 (N_2051,In_210,In_400);
nand U2052 (N_2052,In_812,In_188);
nor U2053 (N_2053,In_687,In_144);
and U2054 (N_2054,In_801,In_786);
nand U2055 (N_2055,In_678,In_564);
and U2056 (N_2056,In_617,In_455);
nor U2057 (N_2057,In_434,In_269);
and U2058 (N_2058,In_501,In_659);
or U2059 (N_2059,In_516,In_858);
nand U2060 (N_2060,In_726,In_47);
nor U2061 (N_2061,In_275,In_639);
nor U2062 (N_2062,In_394,In_206);
and U2063 (N_2063,In_132,In_681);
nor U2064 (N_2064,In_440,In_305);
and U2065 (N_2065,In_886,In_602);
nor U2066 (N_2066,In_627,In_175);
nand U2067 (N_2067,In_370,In_511);
or U2068 (N_2068,In_278,In_589);
nand U2069 (N_2069,In_67,In_800);
and U2070 (N_2070,In_412,In_807);
nand U2071 (N_2071,In_923,In_434);
nor U2072 (N_2072,In_759,In_196);
nand U2073 (N_2073,In_987,In_105);
or U2074 (N_2074,In_579,In_617);
and U2075 (N_2075,In_944,In_862);
nor U2076 (N_2076,In_250,In_665);
and U2077 (N_2077,In_58,In_86);
and U2078 (N_2078,In_841,In_570);
and U2079 (N_2079,In_198,In_534);
nand U2080 (N_2080,In_945,In_597);
and U2081 (N_2081,In_22,In_655);
or U2082 (N_2082,In_1,In_819);
nand U2083 (N_2083,In_612,In_894);
and U2084 (N_2084,In_144,In_719);
nand U2085 (N_2085,In_197,In_755);
or U2086 (N_2086,In_318,In_170);
or U2087 (N_2087,In_669,In_196);
or U2088 (N_2088,In_925,In_14);
or U2089 (N_2089,In_151,In_777);
and U2090 (N_2090,In_508,In_292);
nor U2091 (N_2091,In_94,In_923);
nand U2092 (N_2092,In_760,In_804);
and U2093 (N_2093,In_645,In_124);
or U2094 (N_2094,In_569,In_688);
nor U2095 (N_2095,In_90,In_218);
nand U2096 (N_2096,In_234,In_347);
nor U2097 (N_2097,In_932,In_720);
or U2098 (N_2098,In_115,In_133);
and U2099 (N_2099,In_552,In_187);
and U2100 (N_2100,In_89,In_691);
or U2101 (N_2101,In_449,In_994);
nand U2102 (N_2102,In_812,In_246);
or U2103 (N_2103,In_444,In_306);
nand U2104 (N_2104,In_531,In_191);
nor U2105 (N_2105,In_478,In_754);
or U2106 (N_2106,In_662,In_663);
or U2107 (N_2107,In_84,In_419);
and U2108 (N_2108,In_287,In_735);
nand U2109 (N_2109,In_96,In_650);
and U2110 (N_2110,In_992,In_756);
and U2111 (N_2111,In_996,In_522);
nand U2112 (N_2112,In_259,In_299);
and U2113 (N_2113,In_612,In_517);
nand U2114 (N_2114,In_10,In_600);
nand U2115 (N_2115,In_639,In_493);
or U2116 (N_2116,In_368,In_293);
nor U2117 (N_2117,In_405,In_537);
nor U2118 (N_2118,In_749,In_687);
nand U2119 (N_2119,In_367,In_369);
and U2120 (N_2120,In_789,In_936);
nand U2121 (N_2121,In_35,In_846);
or U2122 (N_2122,In_345,In_846);
and U2123 (N_2123,In_546,In_181);
xor U2124 (N_2124,In_49,In_333);
or U2125 (N_2125,In_903,In_126);
and U2126 (N_2126,In_383,In_376);
and U2127 (N_2127,In_143,In_808);
or U2128 (N_2128,In_959,In_386);
nand U2129 (N_2129,In_429,In_891);
and U2130 (N_2130,In_569,In_604);
xnor U2131 (N_2131,In_809,In_98);
nor U2132 (N_2132,In_235,In_336);
and U2133 (N_2133,In_755,In_467);
or U2134 (N_2134,In_945,In_744);
and U2135 (N_2135,In_773,In_41);
nand U2136 (N_2136,In_429,In_733);
nor U2137 (N_2137,In_995,In_206);
and U2138 (N_2138,In_560,In_582);
nor U2139 (N_2139,In_401,In_283);
nor U2140 (N_2140,In_940,In_436);
nand U2141 (N_2141,In_516,In_437);
nor U2142 (N_2142,In_601,In_720);
nand U2143 (N_2143,In_516,In_478);
or U2144 (N_2144,In_807,In_444);
and U2145 (N_2145,In_554,In_225);
and U2146 (N_2146,In_239,In_155);
and U2147 (N_2147,In_91,In_613);
and U2148 (N_2148,In_122,In_304);
xor U2149 (N_2149,In_689,In_784);
nand U2150 (N_2150,In_199,In_882);
nor U2151 (N_2151,In_413,In_383);
nor U2152 (N_2152,In_508,In_564);
and U2153 (N_2153,In_305,In_260);
nor U2154 (N_2154,In_595,In_683);
nor U2155 (N_2155,In_468,In_83);
nand U2156 (N_2156,In_928,In_708);
nand U2157 (N_2157,In_638,In_432);
nand U2158 (N_2158,In_650,In_416);
and U2159 (N_2159,In_643,In_360);
nand U2160 (N_2160,In_729,In_981);
or U2161 (N_2161,In_710,In_995);
nand U2162 (N_2162,In_153,In_716);
and U2163 (N_2163,In_939,In_851);
nor U2164 (N_2164,In_700,In_651);
and U2165 (N_2165,In_586,In_558);
or U2166 (N_2166,In_403,In_407);
nor U2167 (N_2167,In_716,In_229);
nor U2168 (N_2168,In_798,In_254);
nand U2169 (N_2169,In_150,In_95);
and U2170 (N_2170,In_438,In_14);
nand U2171 (N_2171,In_886,In_567);
nor U2172 (N_2172,In_464,In_261);
nor U2173 (N_2173,In_269,In_185);
and U2174 (N_2174,In_195,In_629);
and U2175 (N_2175,In_768,In_595);
nand U2176 (N_2176,In_53,In_975);
nor U2177 (N_2177,In_533,In_148);
or U2178 (N_2178,In_465,In_833);
or U2179 (N_2179,In_874,In_72);
and U2180 (N_2180,In_100,In_79);
nor U2181 (N_2181,In_260,In_108);
and U2182 (N_2182,In_594,In_50);
and U2183 (N_2183,In_625,In_353);
nand U2184 (N_2184,In_698,In_552);
nand U2185 (N_2185,In_651,In_62);
nor U2186 (N_2186,In_884,In_573);
or U2187 (N_2187,In_463,In_966);
and U2188 (N_2188,In_372,In_581);
and U2189 (N_2189,In_156,In_832);
nand U2190 (N_2190,In_561,In_64);
nand U2191 (N_2191,In_161,In_463);
nand U2192 (N_2192,In_664,In_394);
nand U2193 (N_2193,In_709,In_543);
nand U2194 (N_2194,In_81,In_239);
nand U2195 (N_2195,In_839,In_935);
nand U2196 (N_2196,In_474,In_57);
and U2197 (N_2197,In_261,In_892);
or U2198 (N_2198,In_307,In_242);
or U2199 (N_2199,In_919,In_184);
nand U2200 (N_2200,In_320,In_673);
or U2201 (N_2201,In_770,In_439);
or U2202 (N_2202,In_597,In_113);
or U2203 (N_2203,In_118,In_907);
nand U2204 (N_2204,In_589,In_910);
and U2205 (N_2205,In_677,In_689);
or U2206 (N_2206,In_384,In_411);
or U2207 (N_2207,In_263,In_379);
or U2208 (N_2208,In_337,In_796);
nand U2209 (N_2209,In_271,In_253);
xnor U2210 (N_2210,In_305,In_683);
and U2211 (N_2211,In_236,In_721);
or U2212 (N_2212,In_239,In_845);
and U2213 (N_2213,In_264,In_939);
and U2214 (N_2214,In_140,In_632);
or U2215 (N_2215,In_749,In_529);
nand U2216 (N_2216,In_500,In_667);
nor U2217 (N_2217,In_183,In_424);
or U2218 (N_2218,In_20,In_421);
and U2219 (N_2219,In_689,In_592);
xor U2220 (N_2220,In_261,In_454);
nand U2221 (N_2221,In_761,In_522);
or U2222 (N_2222,In_548,In_40);
nor U2223 (N_2223,In_498,In_983);
and U2224 (N_2224,In_242,In_254);
nor U2225 (N_2225,In_462,In_389);
and U2226 (N_2226,In_16,In_55);
and U2227 (N_2227,In_505,In_469);
nor U2228 (N_2228,In_467,In_607);
or U2229 (N_2229,In_280,In_232);
or U2230 (N_2230,In_676,In_881);
and U2231 (N_2231,In_200,In_936);
or U2232 (N_2232,In_709,In_217);
nand U2233 (N_2233,In_751,In_897);
or U2234 (N_2234,In_927,In_287);
nand U2235 (N_2235,In_41,In_273);
nor U2236 (N_2236,In_68,In_219);
and U2237 (N_2237,In_198,In_948);
or U2238 (N_2238,In_96,In_14);
and U2239 (N_2239,In_174,In_256);
nand U2240 (N_2240,In_915,In_949);
or U2241 (N_2241,In_712,In_526);
xor U2242 (N_2242,In_730,In_653);
and U2243 (N_2243,In_50,In_345);
nand U2244 (N_2244,In_219,In_262);
nor U2245 (N_2245,In_534,In_769);
nor U2246 (N_2246,In_989,In_591);
nand U2247 (N_2247,In_73,In_239);
nand U2248 (N_2248,In_639,In_787);
or U2249 (N_2249,In_955,In_223);
nand U2250 (N_2250,In_719,In_643);
or U2251 (N_2251,In_678,In_249);
nand U2252 (N_2252,In_632,In_230);
and U2253 (N_2253,In_421,In_270);
nand U2254 (N_2254,In_742,In_894);
nand U2255 (N_2255,In_27,In_848);
or U2256 (N_2256,In_140,In_716);
nor U2257 (N_2257,In_618,In_41);
nor U2258 (N_2258,In_254,In_613);
nor U2259 (N_2259,In_51,In_283);
nand U2260 (N_2260,In_671,In_67);
or U2261 (N_2261,In_979,In_404);
or U2262 (N_2262,In_377,In_427);
nand U2263 (N_2263,In_21,In_712);
nor U2264 (N_2264,In_987,In_464);
nand U2265 (N_2265,In_57,In_338);
nand U2266 (N_2266,In_695,In_624);
or U2267 (N_2267,In_463,In_65);
nor U2268 (N_2268,In_135,In_472);
or U2269 (N_2269,In_76,In_921);
or U2270 (N_2270,In_352,In_177);
or U2271 (N_2271,In_456,In_172);
nor U2272 (N_2272,In_791,In_729);
or U2273 (N_2273,In_647,In_35);
nand U2274 (N_2274,In_432,In_919);
nand U2275 (N_2275,In_569,In_35);
nor U2276 (N_2276,In_515,In_727);
and U2277 (N_2277,In_915,In_702);
nand U2278 (N_2278,In_600,In_213);
nand U2279 (N_2279,In_892,In_362);
nor U2280 (N_2280,In_715,In_865);
nor U2281 (N_2281,In_504,In_323);
nor U2282 (N_2282,In_391,In_602);
nor U2283 (N_2283,In_890,In_813);
nand U2284 (N_2284,In_892,In_99);
nand U2285 (N_2285,In_283,In_424);
nand U2286 (N_2286,In_734,In_136);
and U2287 (N_2287,In_237,In_582);
and U2288 (N_2288,In_577,In_37);
or U2289 (N_2289,In_815,In_505);
nand U2290 (N_2290,In_594,In_933);
nor U2291 (N_2291,In_104,In_846);
or U2292 (N_2292,In_491,In_533);
nor U2293 (N_2293,In_504,In_946);
nor U2294 (N_2294,In_683,In_78);
or U2295 (N_2295,In_70,In_681);
and U2296 (N_2296,In_624,In_483);
nand U2297 (N_2297,In_790,In_244);
or U2298 (N_2298,In_117,In_914);
nand U2299 (N_2299,In_710,In_464);
and U2300 (N_2300,In_379,In_771);
nand U2301 (N_2301,In_684,In_953);
nor U2302 (N_2302,In_889,In_14);
and U2303 (N_2303,In_294,In_202);
and U2304 (N_2304,In_988,In_419);
and U2305 (N_2305,In_743,In_806);
and U2306 (N_2306,In_317,In_165);
or U2307 (N_2307,In_550,In_142);
or U2308 (N_2308,In_885,In_778);
nor U2309 (N_2309,In_58,In_981);
nor U2310 (N_2310,In_446,In_283);
and U2311 (N_2311,In_939,In_749);
and U2312 (N_2312,In_565,In_644);
nand U2313 (N_2313,In_394,In_930);
or U2314 (N_2314,In_834,In_296);
and U2315 (N_2315,In_224,In_113);
nor U2316 (N_2316,In_35,In_261);
nor U2317 (N_2317,In_240,In_475);
or U2318 (N_2318,In_909,In_601);
nor U2319 (N_2319,In_625,In_14);
and U2320 (N_2320,In_194,In_701);
or U2321 (N_2321,In_982,In_290);
and U2322 (N_2322,In_560,In_544);
nand U2323 (N_2323,In_615,In_687);
nand U2324 (N_2324,In_728,In_33);
nor U2325 (N_2325,In_654,In_819);
nand U2326 (N_2326,In_850,In_740);
nand U2327 (N_2327,In_916,In_24);
nand U2328 (N_2328,In_688,In_715);
and U2329 (N_2329,In_645,In_369);
or U2330 (N_2330,In_612,In_412);
nor U2331 (N_2331,In_396,In_300);
nor U2332 (N_2332,In_161,In_197);
and U2333 (N_2333,In_808,In_489);
nor U2334 (N_2334,In_240,In_216);
nor U2335 (N_2335,In_667,In_964);
nand U2336 (N_2336,In_635,In_377);
nand U2337 (N_2337,In_418,In_481);
nor U2338 (N_2338,In_185,In_779);
and U2339 (N_2339,In_918,In_212);
and U2340 (N_2340,In_786,In_836);
or U2341 (N_2341,In_693,In_688);
and U2342 (N_2342,In_1,In_291);
and U2343 (N_2343,In_472,In_494);
or U2344 (N_2344,In_937,In_407);
nand U2345 (N_2345,In_547,In_829);
nand U2346 (N_2346,In_533,In_234);
nand U2347 (N_2347,In_892,In_519);
nor U2348 (N_2348,In_226,In_340);
nor U2349 (N_2349,In_118,In_234);
or U2350 (N_2350,In_322,In_515);
or U2351 (N_2351,In_544,In_145);
nor U2352 (N_2352,In_213,In_407);
nor U2353 (N_2353,In_182,In_577);
and U2354 (N_2354,In_424,In_731);
or U2355 (N_2355,In_48,In_294);
nor U2356 (N_2356,In_853,In_263);
nor U2357 (N_2357,In_68,In_879);
nand U2358 (N_2358,In_54,In_207);
nor U2359 (N_2359,In_796,In_682);
and U2360 (N_2360,In_606,In_575);
or U2361 (N_2361,In_368,In_273);
nor U2362 (N_2362,In_510,In_287);
or U2363 (N_2363,In_603,In_362);
and U2364 (N_2364,In_178,In_421);
or U2365 (N_2365,In_441,In_363);
or U2366 (N_2366,In_854,In_521);
or U2367 (N_2367,In_387,In_162);
nor U2368 (N_2368,In_712,In_226);
nand U2369 (N_2369,In_564,In_347);
nor U2370 (N_2370,In_816,In_464);
nand U2371 (N_2371,In_103,In_688);
and U2372 (N_2372,In_996,In_290);
and U2373 (N_2373,In_165,In_284);
nand U2374 (N_2374,In_463,In_234);
or U2375 (N_2375,In_705,In_327);
xor U2376 (N_2376,In_772,In_922);
or U2377 (N_2377,In_613,In_608);
nand U2378 (N_2378,In_210,In_800);
nand U2379 (N_2379,In_908,In_944);
or U2380 (N_2380,In_83,In_571);
nor U2381 (N_2381,In_558,In_304);
nor U2382 (N_2382,In_558,In_869);
or U2383 (N_2383,In_417,In_175);
or U2384 (N_2384,In_224,In_68);
nor U2385 (N_2385,In_979,In_500);
and U2386 (N_2386,In_725,In_640);
nand U2387 (N_2387,In_661,In_149);
nand U2388 (N_2388,In_357,In_420);
nor U2389 (N_2389,In_135,In_639);
nor U2390 (N_2390,In_860,In_829);
nand U2391 (N_2391,In_536,In_597);
or U2392 (N_2392,In_262,In_767);
and U2393 (N_2393,In_598,In_352);
xnor U2394 (N_2394,In_636,In_491);
nand U2395 (N_2395,In_53,In_816);
nand U2396 (N_2396,In_980,In_90);
and U2397 (N_2397,In_362,In_70);
or U2398 (N_2398,In_743,In_579);
nor U2399 (N_2399,In_829,In_799);
nor U2400 (N_2400,In_580,In_767);
nand U2401 (N_2401,In_252,In_219);
and U2402 (N_2402,In_907,In_539);
or U2403 (N_2403,In_165,In_447);
nor U2404 (N_2404,In_658,In_743);
or U2405 (N_2405,In_929,In_934);
and U2406 (N_2406,In_808,In_613);
or U2407 (N_2407,In_518,In_117);
or U2408 (N_2408,In_703,In_950);
or U2409 (N_2409,In_15,In_242);
or U2410 (N_2410,In_105,In_945);
and U2411 (N_2411,In_402,In_317);
or U2412 (N_2412,In_347,In_199);
nor U2413 (N_2413,In_850,In_967);
or U2414 (N_2414,In_115,In_383);
nor U2415 (N_2415,In_623,In_962);
and U2416 (N_2416,In_383,In_297);
and U2417 (N_2417,In_718,In_599);
nand U2418 (N_2418,In_57,In_259);
or U2419 (N_2419,In_494,In_830);
and U2420 (N_2420,In_163,In_835);
xnor U2421 (N_2421,In_101,In_179);
or U2422 (N_2422,In_893,In_478);
and U2423 (N_2423,In_477,In_173);
xnor U2424 (N_2424,In_69,In_316);
nand U2425 (N_2425,In_86,In_615);
nand U2426 (N_2426,In_164,In_64);
nor U2427 (N_2427,In_848,In_507);
nand U2428 (N_2428,In_433,In_131);
or U2429 (N_2429,In_254,In_172);
or U2430 (N_2430,In_212,In_963);
and U2431 (N_2431,In_710,In_285);
nor U2432 (N_2432,In_584,In_871);
or U2433 (N_2433,In_910,In_395);
nor U2434 (N_2434,In_252,In_584);
or U2435 (N_2435,In_64,In_254);
nand U2436 (N_2436,In_356,In_637);
or U2437 (N_2437,In_455,In_345);
and U2438 (N_2438,In_191,In_286);
nor U2439 (N_2439,In_724,In_31);
or U2440 (N_2440,In_285,In_941);
or U2441 (N_2441,In_372,In_889);
nand U2442 (N_2442,In_220,In_576);
or U2443 (N_2443,In_116,In_52);
nand U2444 (N_2444,In_663,In_449);
nor U2445 (N_2445,In_902,In_985);
or U2446 (N_2446,In_536,In_192);
or U2447 (N_2447,In_880,In_185);
and U2448 (N_2448,In_937,In_744);
and U2449 (N_2449,In_781,In_169);
nor U2450 (N_2450,In_351,In_210);
and U2451 (N_2451,In_998,In_148);
nor U2452 (N_2452,In_559,In_128);
nand U2453 (N_2453,In_602,In_762);
or U2454 (N_2454,In_536,In_828);
and U2455 (N_2455,In_863,In_891);
or U2456 (N_2456,In_756,In_270);
nand U2457 (N_2457,In_187,In_91);
or U2458 (N_2458,In_200,In_56);
or U2459 (N_2459,In_730,In_358);
nand U2460 (N_2460,In_67,In_55);
nand U2461 (N_2461,In_59,In_563);
nor U2462 (N_2462,In_504,In_218);
and U2463 (N_2463,In_637,In_983);
nand U2464 (N_2464,In_480,In_530);
and U2465 (N_2465,In_248,In_100);
and U2466 (N_2466,In_621,In_692);
nand U2467 (N_2467,In_43,In_373);
nand U2468 (N_2468,In_503,In_692);
or U2469 (N_2469,In_403,In_313);
and U2470 (N_2470,In_267,In_266);
nor U2471 (N_2471,In_361,In_100);
nand U2472 (N_2472,In_319,In_532);
and U2473 (N_2473,In_247,In_547);
nand U2474 (N_2474,In_942,In_420);
nand U2475 (N_2475,In_244,In_119);
and U2476 (N_2476,In_357,In_3);
nand U2477 (N_2477,In_391,In_423);
nand U2478 (N_2478,In_441,In_707);
nor U2479 (N_2479,In_121,In_345);
or U2480 (N_2480,In_487,In_591);
and U2481 (N_2481,In_546,In_640);
and U2482 (N_2482,In_719,In_226);
nand U2483 (N_2483,In_640,In_207);
nor U2484 (N_2484,In_638,In_251);
or U2485 (N_2485,In_19,In_144);
and U2486 (N_2486,In_740,In_237);
and U2487 (N_2487,In_551,In_754);
and U2488 (N_2488,In_228,In_561);
and U2489 (N_2489,In_477,In_743);
nand U2490 (N_2490,In_945,In_49);
and U2491 (N_2491,In_197,In_236);
and U2492 (N_2492,In_911,In_245);
and U2493 (N_2493,In_133,In_549);
nand U2494 (N_2494,In_394,In_528);
nor U2495 (N_2495,In_46,In_909);
or U2496 (N_2496,In_627,In_308);
nor U2497 (N_2497,In_923,In_111);
and U2498 (N_2498,In_749,In_82);
nor U2499 (N_2499,In_345,In_192);
nor U2500 (N_2500,N_598,N_2454);
and U2501 (N_2501,N_2000,N_2141);
or U2502 (N_2502,N_500,N_619);
and U2503 (N_2503,N_1401,N_1637);
and U2504 (N_2504,N_239,N_632);
nor U2505 (N_2505,N_1222,N_1970);
and U2506 (N_2506,N_1751,N_1670);
and U2507 (N_2507,N_614,N_2069);
or U2508 (N_2508,N_1536,N_1785);
nor U2509 (N_2509,N_235,N_553);
nand U2510 (N_2510,N_1172,N_2497);
nor U2511 (N_2511,N_1890,N_939);
and U2512 (N_2512,N_813,N_1052);
or U2513 (N_2513,N_1036,N_208);
or U2514 (N_2514,N_55,N_707);
nand U2515 (N_2515,N_1618,N_847);
nand U2516 (N_2516,N_1100,N_930);
nor U2517 (N_2517,N_514,N_279);
nor U2518 (N_2518,N_1136,N_1723);
nand U2519 (N_2519,N_521,N_1214);
or U2520 (N_2520,N_2470,N_1910);
nand U2521 (N_2521,N_1821,N_430);
or U2522 (N_2522,N_2476,N_1623);
nor U2523 (N_2523,N_1523,N_482);
or U2524 (N_2524,N_1883,N_487);
and U2525 (N_2525,N_1125,N_1671);
or U2526 (N_2526,N_1397,N_1763);
and U2527 (N_2527,N_2293,N_1162);
or U2528 (N_2528,N_151,N_1496);
nand U2529 (N_2529,N_1105,N_330);
nand U2530 (N_2530,N_1825,N_400);
or U2531 (N_2531,N_856,N_1895);
or U2532 (N_2532,N_902,N_2332);
nand U2533 (N_2533,N_2243,N_862);
or U2534 (N_2534,N_2240,N_977);
nand U2535 (N_2535,N_1188,N_1983);
nor U2536 (N_2536,N_1555,N_1363);
nand U2537 (N_2537,N_244,N_748);
or U2538 (N_2538,N_2196,N_32);
or U2539 (N_2539,N_1792,N_1131);
nand U2540 (N_2540,N_409,N_1873);
and U2541 (N_2541,N_2194,N_1589);
nand U2542 (N_2542,N_1416,N_1005);
and U2543 (N_2543,N_982,N_2094);
nor U2544 (N_2544,N_2166,N_2354);
or U2545 (N_2545,N_507,N_999);
or U2546 (N_2546,N_451,N_2415);
or U2547 (N_2547,N_2359,N_2182);
nand U2548 (N_2548,N_1077,N_1722);
and U2549 (N_2549,N_668,N_323);
nand U2550 (N_2550,N_936,N_273);
nand U2551 (N_2551,N_1559,N_2384);
or U2552 (N_2552,N_25,N_370);
nand U2553 (N_2553,N_70,N_531);
nor U2554 (N_2554,N_1761,N_322);
nand U2555 (N_2555,N_876,N_2098);
nor U2556 (N_2556,N_1046,N_633);
nor U2557 (N_2557,N_1231,N_192);
and U2558 (N_2558,N_1694,N_528);
and U2559 (N_2559,N_2330,N_1211);
nor U2560 (N_2560,N_1215,N_561);
nor U2561 (N_2561,N_2260,N_1123);
nor U2562 (N_2562,N_1715,N_1612);
or U2563 (N_2563,N_2372,N_2483);
nand U2564 (N_2564,N_1812,N_1894);
nor U2565 (N_2565,N_935,N_1993);
nor U2566 (N_2566,N_263,N_1846);
nor U2567 (N_2567,N_1610,N_866);
and U2568 (N_2568,N_144,N_2192);
and U2569 (N_2569,N_1340,N_1750);
and U2570 (N_2570,N_2324,N_1278);
or U2571 (N_2571,N_334,N_2177);
nand U2572 (N_2572,N_2073,N_307);
and U2573 (N_2573,N_1614,N_694);
nand U2574 (N_2574,N_1755,N_1980);
nor U2575 (N_2575,N_275,N_643);
or U2576 (N_2576,N_824,N_351);
nor U2577 (N_2577,N_563,N_1547);
or U2578 (N_2578,N_1598,N_1663);
nor U2579 (N_2579,N_420,N_1431);
or U2580 (N_2580,N_1691,N_1988);
or U2581 (N_2581,N_1674,N_1745);
or U2582 (N_2582,N_1251,N_538);
nor U2583 (N_2583,N_234,N_2199);
and U2584 (N_2584,N_529,N_242);
nor U2585 (N_2585,N_1704,N_1420);
or U2586 (N_2586,N_166,N_685);
nor U2587 (N_2587,N_600,N_392);
nor U2588 (N_2588,N_2011,N_455);
nand U2589 (N_2589,N_2429,N_286);
nand U2590 (N_2590,N_1133,N_1306);
or U2591 (N_2591,N_1078,N_419);
nor U2592 (N_2592,N_893,N_59);
nand U2593 (N_2593,N_1774,N_1398);
nand U2594 (N_2594,N_365,N_426);
nand U2595 (N_2595,N_319,N_2132);
and U2596 (N_2596,N_1327,N_312);
nor U2597 (N_2597,N_186,N_2418);
and U2598 (N_2598,N_708,N_2436);
or U2599 (N_2599,N_1659,N_1857);
nor U2600 (N_2600,N_2452,N_1951);
or U2601 (N_2601,N_2446,N_1926);
or U2602 (N_2602,N_1545,N_288);
or U2603 (N_2603,N_794,N_990);
and U2604 (N_2604,N_1570,N_1878);
nand U2605 (N_2605,N_2118,N_2028);
nor U2606 (N_2606,N_280,N_1180);
or U2607 (N_2607,N_1140,N_179);
xor U2608 (N_2608,N_1365,N_1483);
and U2609 (N_2609,N_2112,N_397);
and U2610 (N_2610,N_1702,N_301);
nor U2611 (N_2611,N_2485,N_1320);
nand U2612 (N_2612,N_126,N_1409);
nor U2613 (N_2613,N_372,N_639);
and U2614 (N_2614,N_1002,N_2250);
nand U2615 (N_2615,N_1054,N_806);
nor U2616 (N_2616,N_369,N_1647);
or U2617 (N_2617,N_595,N_2152);
nor U2618 (N_2618,N_1060,N_1047);
and U2619 (N_2619,N_1274,N_247);
and U2620 (N_2620,N_2216,N_249);
nand U2621 (N_2621,N_1777,N_1317);
nor U2622 (N_2622,N_1,N_2238);
or U2623 (N_2623,N_2374,N_1972);
or U2624 (N_2624,N_756,N_406);
nand U2625 (N_2625,N_122,N_1515);
nor U2626 (N_2626,N_2426,N_2060);
or U2627 (N_2627,N_2265,N_2311);
nor U2628 (N_2628,N_590,N_1403);
nor U2629 (N_2629,N_1126,N_997);
and U2630 (N_2630,N_2255,N_1958);
and U2631 (N_2631,N_676,N_548);
and U2632 (N_2632,N_1906,N_2278);
nand U2633 (N_2633,N_1175,N_1801);
and U2634 (N_2634,N_664,N_1497);
and U2635 (N_2635,N_408,N_2190);
and U2636 (N_2636,N_779,N_1934);
and U2637 (N_2637,N_1087,N_470);
and U2638 (N_2638,N_1262,N_102);
nand U2639 (N_2639,N_735,N_2154);
nand U2640 (N_2640,N_2391,N_497);
nand U2641 (N_2641,N_1527,N_1923);
nor U2642 (N_2642,N_1139,N_2191);
and U2643 (N_2643,N_1645,N_724);
nor U2644 (N_2644,N_276,N_27);
nor U2645 (N_2645,N_1423,N_1479);
nand U2646 (N_2646,N_1649,N_942);
or U2647 (N_2647,N_172,N_360);
nand U2648 (N_2648,N_2025,N_30);
or U2649 (N_2649,N_377,N_1221);
nand U2650 (N_2650,N_1535,N_1082);
nor U2651 (N_2651,N_927,N_1061);
or U2652 (N_2652,N_270,N_1503);
and U2653 (N_2653,N_989,N_1151);
and U2654 (N_2654,N_814,N_1045);
nor U2655 (N_2655,N_700,N_185);
xor U2656 (N_2656,N_2172,N_2258);
or U2657 (N_2657,N_587,N_907);
or U2658 (N_2658,N_568,N_1466);
or U2659 (N_2659,N_1871,N_325);
or U2660 (N_2660,N_599,N_1177);
or U2661 (N_2661,N_1626,N_1942);
and U2662 (N_2662,N_1815,N_1817);
nor U2663 (N_2663,N_2399,N_2394);
or U2664 (N_2664,N_456,N_2246);
nand U2665 (N_2665,N_2296,N_1309);
nand U2666 (N_2666,N_1952,N_106);
nand U2667 (N_2667,N_560,N_543);
and U2668 (N_2668,N_1676,N_630);
nor U2669 (N_2669,N_1584,N_875);
nand U2670 (N_2670,N_373,N_679);
nor U2671 (N_2671,N_383,N_506);
and U2672 (N_2672,N_692,N_1673);
nor U2673 (N_2673,N_1516,N_250);
and U2674 (N_2674,N_463,N_1322);
and U2675 (N_2675,N_1587,N_1549);
nand U2676 (N_2676,N_719,N_946);
and U2677 (N_2677,N_1014,N_1351);
and U2678 (N_2678,N_1482,N_2186);
nor U2679 (N_2679,N_2353,N_1839);
or U2680 (N_2680,N_2252,N_1369);
or U2681 (N_2681,N_1950,N_608);
or U2682 (N_2682,N_398,N_318);
and U2683 (N_2683,N_1622,N_2085);
nand U2684 (N_2684,N_264,N_1362);
and U2685 (N_2685,N_2035,N_403);
nor U2686 (N_2686,N_892,N_2213);
nand U2687 (N_2687,N_1399,N_1458);
and U2688 (N_2688,N_142,N_304);
or U2689 (N_2689,N_1684,N_1240);
or U2690 (N_2690,N_1281,N_647);
nand U2691 (N_2691,N_603,N_1744);
nor U2692 (N_2692,N_1764,N_2390);
or U2693 (N_2693,N_138,N_113);
nor U2694 (N_2694,N_1513,N_282);
and U2695 (N_2695,N_1145,N_18);
or U2696 (N_2696,N_1156,N_364);
and U2697 (N_2697,N_859,N_63);
and U2698 (N_2698,N_363,N_874);
and U2699 (N_2699,N_1245,N_1590);
and U2700 (N_2700,N_2107,N_1625);
and U2701 (N_2701,N_484,N_417);
and U2702 (N_2702,N_1802,N_520);
nand U2703 (N_2703,N_1696,N_1708);
or U2704 (N_2704,N_136,N_2496);
or U2705 (N_2705,N_786,N_910);
or U2706 (N_2706,N_2010,N_648);
or U2707 (N_2707,N_976,N_99);
and U2708 (N_2708,N_1630,N_1820);
nor U2709 (N_2709,N_1266,N_423);
nor U2710 (N_2710,N_165,N_2041);
nor U2711 (N_2711,N_1378,N_2326);
nor U2712 (N_2712,N_453,N_2468);
nor U2713 (N_2713,N_652,N_2198);
nor U2714 (N_2714,N_958,N_1079);
and U2715 (N_2715,N_1657,N_2205);
nor U2716 (N_2716,N_2122,N_1834);
or U2717 (N_2717,N_1091,N_1025);
nor U2718 (N_2718,N_810,N_2364);
nand U2719 (N_2719,N_1330,N_1434);
nand U2720 (N_2720,N_2153,N_566);
nand U2721 (N_2721,N_624,N_160);
nand U2722 (N_2722,N_836,N_156);
or U2723 (N_2723,N_436,N_1471);
nor U2724 (N_2724,N_326,N_311);
and U2725 (N_2725,N_747,N_1387);
or U2726 (N_2726,N_517,N_1581);
or U2727 (N_2727,N_1160,N_2480);
nor U2728 (N_2728,N_467,N_772);
nor U2729 (N_2729,N_2059,N_1573);
or U2730 (N_2730,N_1400,N_1049);
or U2731 (N_2731,N_914,N_1752);
nor U2732 (N_2732,N_2239,N_2076);
or U2733 (N_2733,N_1903,N_1294);
nand U2734 (N_2734,N_97,N_2437);
and U2735 (N_2735,N_511,N_1171);
and U2736 (N_2736,N_1796,N_1701);
nor U2737 (N_2737,N_1411,N_868);
nand U2738 (N_2738,N_1747,N_580);
or U2739 (N_2739,N_2314,N_491);
or U2740 (N_2740,N_127,N_1769);
and U2741 (N_2741,N_1944,N_840);
xor U2742 (N_2742,N_955,N_1628);
nand U2743 (N_2743,N_1203,N_585);
nand U2744 (N_2744,N_2207,N_783);
and U2745 (N_2745,N_1212,N_1687);
and U2746 (N_2746,N_1604,N_1068);
or U2747 (N_2747,N_1481,N_2375);
nor U2748 (N_2748,N_2458,N_35);
or U2749 (N_2749,N_1868,N_1608);
nand U2750 (N_2750,N_1185,N_2037);
nor U2751 (N_2751,N_1427,N_316);
and U2752 (N_2752,N_1896,N_1553);
nand U2753 (N_2753,N_1838,N_662);
nand U2754 (N_2754,N_2195,N_80);
nand U2755 (N_2755,N_488,N_2348);
nand U2756 (N_2756,N_2086,N_1973);
nand U2757 (N_2757,N_2280,N_336);
or U2758 (N_2758,N_1524,N_203);
nor U2759 (N_2759,N_920,N_1564);
and U2760 (N_2760,N_386,N_428);
and U2761 (N_2761,N_65,N_2309);
nor U2762 (N_2762,N_757,N_486);
or U2763 (N_2763,N_848,N_2137);
nand U2764 (N_2764,N_1227,N_680);
nor U2765 (N_2765,N_1338,N_1765);
or U2766 (N_2766,N_1729,N_909);
nor U2767 (N_2767,N_2170,N_1753);
or U2768 (N_2768,N_672,N_901);
nor U2769 (N_2769,N_2082,N_2469);
or U2770 (N_2770,N_1682,N_2471);
or U2771 (N_2771,N_303,N_2263);
nor U2772 (N_2772,N_1293,N_900);
and U2773 (N_2773,N_1603,N_464);
or U2774 (N_2774,N_1108,N_489);
and U2775 (N_2775,N_737,N_3);
nand U2776 (N_2776,N_1933,N_1858);
nand U2777 (N_2777,N_2481,N_1992);
or U2778 (N_2778,N_2108,N_1578);
or U2779 (N_2779,N_2413,N_254);
nand U2780 (N_2780,N_1022,N_2002);
nor U2781 (N_2781,N_36,N_492);
or U2782 (N_2782,N_434,N_960);
xnor U2783 (N_2783,N_744,N_2345);
nor U2784 (N_2784,N_642,N_2462);
nor U2785 (N_2785,N_272,N_1892);
nand U2786 (N_2786,N_1721,N_1885);
nor U2787 (N_2787,N_709,N_1342);
and U2788 (N_2788,N_758,N_1899);
nor U2789 (N_2789,N_2008,N_0);
and U2790 (N_2790,N_629,N_2004);
nor U2791 (N_2791,N_1234,N_554);
and U2792 (N_2792,N_178,N_495);
nand U2793 (N_2793,N_1571,N_1739);
nor U2794 (N_2794,N_2129,N_2030);
and U2795 (N_2795,N_971,N_682);
or U2796 (N_2796,N_2227,N_2165);
nor U2797 (N_2797,N_2395,N_803);
or U2798 (N_2798,N_1771,N_2441);
and U2799 (N_2799,N_512,N_1283);
and U2800 (N_2800,N_2264,N_1498);
nor U2801 (N_2801,N_2211,N_105);
nand U2802 (N_2802,N_1358,N_2036);
nand U2803 (N_2803,N_2079,N_1593);
and U2804 (N_2804,N_1104,N_1572);
and U2805 (N_2805,N_427,N_1472);
nand U2806 (N_2806,N_324,N_2224);
and U2807 (N_2807,N_1019,N_229);
and U2808 (N_2808,N_461,N_1562);
nor U2809 (N_2809,N_2498,N_508);
and U2810 (N_2810,N_1742,N_2051);
or U2811 (N_2811,N_1732,N_1018);
and U2812 (N_2812,N_1597,N_1360);
nor U2813 (N_2813,N_1357,N_1161);
or U2814 (N_2814,N_1965,N_800);
or U2815 (N_2815,N_1383,N_833);
and U2816 (N_2816,N_2155,N_2241);
or U2817 (N_2817,N_2229,N_2105);
and U2818 (N_2818,N_1759,N_344);
or U2819 (N_2819,N_83,N_1909);
and U2820 (N_2820,N_147,N_1441);
or U2821 (N_2821,N_1877,N_1219);
or U2822 (N_2822,N_1272,N_1666);
nand U2823 (N_2823,N_1734,N_2245);
and U2824 (N_2824,N_1001,N_496);
nor U2825 (N_2825,N_2163,N_1864);
nand U2826 (N_2826,N_2464,N_195);
and U2827 (N_2827,N_2231,N_2236);
or U2828 (N_2828,N_261,N_1258);
and U2829 (N_2829,N_1633,N_1493);
or U2830 (N_2830,N_1316,N_2253);
nor U2831 (N_2831,N_1452,N_657);
nor U2832 (N_2832,N_1716,N_769);
and U2833 (N_2833,N_1335,N_277);
and U2834 (N_2834,N_2456,N_1490);
or U2835 (N_2835,N_2408,N_2493);
or U2836 (N_2836,N_983,N_2113);
nor U2837 (N_2837,N_2467,N_245);
and U2838 (N_2838,N_1287,N_1127);
or U2839 (N_2839,N_1263,N_1756);
or U2840 (N_2840,N_466,N_56);
nor U2841 (N_2841,N_1345,N_1476);
nor U2842 (N_2842,N_1920,N_252);
and U2843 (N_2843,N_119,N_212);
and U2844 (N_2844,N_966,N_1308);
and U2845 (N_2845,N_755,N_1170);
or U2846 (N_2846,N_1067,N_968);
and U2847 (N_2847,N_2406,N_2400);
nand U2848 (N_2848,N_1261,N_950);
or U2849 (N_2849,N_2428,N_940);
nor U2850 (N_2850,N_1979,N_253);
nand U2851 (N_2851,N_547,N_957);
or U2852 (N_2852,N_1085,N_116);
nand U2853 (N_2853,N_1455,N_391);
nand U2854 (N_2854,N_2410,N_459);
and U2855 (N_2855,N_1824,N_385);
or U2856 (N_2856,N_2157,N_1310);
nand U2857 (N_2857,N_1806,N_2210);
nand U2858 (N_2858,N_1520,N_1505);
or U2859 (N_2859,N_760,N_1499);
or U2860 (N_2860,N_1787,N_2262);
or U2861 (N_2861,N_1960,N_2338);
and U2862 (N_2862,N_2461,N_359);
or U2863 (N_2863,N_2062,N_1908);
or U2864 (N_2864,N_751,N_1773);
and U2865 (N_2865,N_24,N_2499);
or U2866 (N_2866,N_1665,N_1971);
nand U2867 (N_2867,N_139,N_2201);
or U2868 (N_2868,N_851,N_73);
nor U2869 (N_2869,N_884,N_2465);
nand U2870 (N_2870,N_1333,N_2417);
nand U2871 (N_2871,N_745,N_518);
nor U2872 (N_2872,N_12,N_1433);
nor U2873 (N_2873,N_2063,N_223);
or U2874 (N_2874,N_291,N_636);
nand U2875 (N_2875,N_1617,N_21);
nor U2876 (N_2876,N_2351,N_1065);
and U2877 (N_2877,N_1440,N_2208);
and U2878 (N_2878,N_2222,N_1650);
nor U2879 (N_2879,N_1703,N_1738);
or U2880 (N_2880,N_1176,N_1827);
nor U2881 (N_2881,N_1639,N_1615);
or U2882 (N_2882,N_1237,N_797);
nand U2883 (N_2883,N_82,N_1426);
nand U2884 (N_2884,N_98,N_1024);
nor U2885 (N_2885,N_45,N_23);
and U2886 (N_2886,N_1999,N_191);
or U2887 (N_2887,N_2319,N_29);
or U2888 (N_2888,N_2443,N_2303);
nand U2889 (N_2889,N_1254,N_1737);
or U2890 (N_2890,N_665,N_1301);
nand U2891 (N_2891,N_739,N_450);
and U2892 (N_2892,N_357,N_1748);
or U2893 (N_2893,N_1495,N_623);
nand U2894 (N_2894,N_174,N_1985);
and U2895 (N_2895,N_1681,N_725);
and U2896 (N_2896,N_1887,N_1003);
xor U2897 (N_2897,N_196,N_339);
or U2898 (N_2898,N_1521,N_801);
and U2899 (N_2899,N_970,N_1379);
or U2900 (N_2900,N_534,N_2169);
nand U2901 (N_2901,N_266,N_979);
nor U2902 (N_2902,N_1494,N_292);
nor U2903 (N_2903,N_1350,N_332);
nand U2904 (N_2904,N_1749,N_565);
or U2905 (N_2905,N_790,N_1836);
or U2906 (N_2906,N_306,N_317);
and U2907 (N_2907,N_2267,N_1368);
nor U2908 (N_2908,N_422,N_887);
and U2909 (N_2909,N_678,N_1299);
nand U2910 (N_2910,N_2156,N_842);
nor U2911 (N_2911,N_1478,N_1804);
nand U2912 (N_2912,N_581,N_34);
nor U2913 (N_2913,N_148,N_175);
nand U2914 (N_2914,N_852,N_1809);
nand U2915 (N_2915,N_2420,N_1941);
nand U2916 (N_2916,N_1179,N_618);
and U2917 (N_2917,N_1332,N_1638);
nor U2918 (N_2918,N_1144,N_1150);
nor U2919 (N_2919,N_2386,N_469);
nand U2920 (N_2920,N_527,N_1193);
nand U2921 (N_2921,N_1092,N_827);
nand U2922 (N_2922,N_237,N_1057);
nor U2923 (N_2923,N_443,N_57);
or U2924 (N_2924,N_986,N_41);
nand U2925 (N_2925,N_331,N_1344);
and U2926 (N_2926,N_1252,N_1874);
nand U2927 (N_2927,N_1842,N_962);
or U2928 (N_2928,N_1392,N_28);
nor U2929 (N_2929,N_1473,N_1480);
nor U2930 (N_2930,N_1835,N_1925);
and U2931 (N_2931,N_1823,N_1929);
xor U2932 (N_2932,N_1337,N_429);
and U2933 (N_2933,N_2377,N_780);
nor U2934 (N_2934,N_870,N_540);
nor U2935 (N_2935,N_640,N_2382);
and U2936 (N_2936,N_1326,N_2193);
or U2937 (N_2937,N_2256,N_2230);
nor U2938 (N_2938,N_1157,N_220);
nand U2939 (N_2939,N_2075,N_1978);
and U2940 (N_2940,N_832,N_103);
and U2941 (N_2941,N_898,N_878);
and U2942 (N_2942,N_2214,N_40);
xnor U2943 (N_2943,N_207,N_787);
or U2944 (N_2944,N_2023,N_513);
nand U2945 (N_2945,N_1181,N_524);
nand U2946 (N_2946,N_2232,N_539);
nand U2947 (N_2947,N_115,N_1679);
and U2948 (N_2948,N_1566,N_96);
or U2949 (N_2949,N_2366,N_995);
nand U2950 (N_2950,N_1026,N_1475);
nor U2951 (N_2951,N_1852,N_1149);
and U2952 (N_2952,N_1347,N_802);
nand U2953 (N_2953,N_246,N_1532);
or U2954 (N_2954,N_924,N_869);
nor U2955 (N_2955,N_865,N_502);
and U2956 (N_2956,N_1788,N_219);
or U2957 (N_2957,N_728,N_380);
or U2958 (N_2958,N_731,N_394);
or U2959 (N_2959,N_2247,N_1940);
or U2960 (N_2960,N_1096,N_2147);
or U2961 (N_2961,N_1031,N_2038);
xnor U2962 (N_2962,N_1727,N_673);
and U2963 (N_2963,N_1793,N_2221);
and U2964 (N_2964,N_2181,N_2388);
nand U2965 (N_2965,N_754,N_1195);
and U2966 (N_2966,N_1995,N_2026);
nand U2967 (N_2967,N_1651,N_1064);
and U2968 (N_2968,N_1713,N_1805);
nor U2969 (N_2969,N_1135,N_621);
nor U2970 (N_2970,N_667,N_1289);
and U2971 (N_2971,N_1504,N_1236);
nor U2972 (N_2972,N_1173,N_1946);
nor U2973 (N_2973,N_2432,N_2021);
nand U2974 (N_2974,N_905,N_2312);
or U2975 (N_2975,N_2015,N_2286);
or U2976 (N_2976,N_2357,N_1724);
and U2977 (N_2977,N_1900,N_1303);
or U2978 (N_2978,N_2092,N_67);
and U2979 (N_2979,N_1582,N_155);
and U2980 (N_2980,N_2453,N_1405);
nand U2981 (N_2981,N_1662,N_1837);
or U2982 (N_2982,N_1102,N_2043);
or U2983 (N_2983,N_677,N_1246);
nor U2984 (N_2984,N_199,N_2187);
nor U2985 (N_2985,N_792,N_1530);
or U2986 (N_2986,N_882,N_998);
nand U2987 (N_2987,N_327,N_297);
nor U2988 (N_2988,N_2411,N_811);
and U2989 (N_2989,N_259,N_2111);
nor U2990 (N_2990,N_1841,N_1235);
or U2991 (N_2991,N_972,N_1938);
or U2992 (N_2992,N_438,N_2270);
or U2993 (N_2993,N_387,N_1453);
nand U2994 (N_2994,N_1314,N_663);
or U2995 (N_2995,N_650,N_2318);
or U2996 (N_2996,N_2091,N_634);
nor U2997 (N_2997,N_1353,N_1109);
nor U2998 (N_2998,N_1607,N_1717);
and U2999 (N_2999,N_1089,N_1845);
nor U3000 (N_3000,N_778,N_1451);
or U3001 (N_3001,N_1190,N_308);
nor U3002 (N_3002,N_1319,N_260);
nand U3003 (N_3003,N_1230,N_2218);
nor U3004 (N_3004,N_938,N_1683);
or U3005 (N_3005,N_346,N_2027);
and U3006 (N_3006,N_490,N_1244);
and U3007 (N_3007,N_516,N_925);
nand U3008 (N_3008,N_2033,N_752);
and U3009 (N_3009,N_2042,N_703);
nand U3010 (N_3010,N_1974,N_416);
and U3011 (N_3011,N_674,N_1982);
and U3012 (N_3012,N_2448,N_1056);
nand U3013 (N_3013,N_1830,N_53);
and U3014 (N_3014,N_460,N_2313);
or U3015 (N_3015,N_820,N_1594);
or U3016 (N_3016,N_1438,N_1776);
or U3017 (N_3017,N_1653,N_1027);
or U3018 (N_3018,N_189,N_72);
or U3019 (N_3019,N_919,N_382);
xnor U3020 (N_3020,N_981,N_2289);
or U3021 (N_3021,N_536,N_452);
nor U3022 (N_3022,N_975,N_454);
nor U3023 (N_3023,N_1506,N_433);
nor U3024 (N_3024,N_2093,N_1998);
nand U3025 (N_3025,N_375,N_1781);
nor U3026 (N_3026,N_162,N_807);
nand U3027 (N_3027,N_1205,N_695);
and U3028 (N_3028,N_2110,N_2304);
nand U3029 (N_3029,N_75,N_2449);
or U3030 (N_3030,N_2298,N_5);
nand U3031 (N_3031,N_544,N_2007);
or U3032 (N_3032,N_2327,N_750);
nand U3033 (N_3033,N_638,N_1063);
nand U3034 (N_3034,N_698,N_1115);
and U3035 (N_3035,N_2305,N_671);
or U3036 (N_3036,N_173,N_1276);
and U3037 (N_3037,N_1891,N_1201);
and U3038 (N_3038,N_1850,N_1218);
nand U3039 (N_3039,N_378,N_1356);
nor U3040 (N_3040,N_505,N_2370);
and U3041 (N_3041,N_1937,N_2233);
nor U3042 (N_3042,N_1017,N_1602);
and U3043 (N_3043,N_1847,N_562);
xnor U3044 (N_3044,N_2276,N_537);
or U3045 (N_3045,N_2189,N_1928);
or U3046 (N_3046,N_240,N_2487);
nand U3047 (N_3047,N_1086,N_1331);
nor U3048 (N_3048,N_2095,N_733);
or U3049 (N_3049,N_1620,N_171);
or U3050 (N_3050,N_1968,N_2358);
and U3051 (N_3051,N_2378,N_2459);
or U3052 (N_3052,N_1121,N_1599);
nor U3053 (N_3053,N_2102,N_2368);
or U3054 (N_3054,N_2225,N_2295);
nand U3055 (N_3055,N_233,N_863);
and U3056 (N_3056,N_1917,N_1011);
nand U3057 (N_3057,N_2425,N_215);
or U3058 (N_3058,N_1913,N_2018);
or U3059 (N_3059,N_853,N_1648);
nand U3060 (N_3060,N_2257,N_916);
or U3061 (N_3061,N_2056,N_1927);
or U3062 (N_3062,N_2254,N_1977);
xnor U3063 (N_3063,N_1849,N_1870);
nor U3064 (N_3064,N_33,N_38);
nand U3065 (N_3065,N_1292,N_1956);
or U3066 (N_3066,N_2299,N_917);
nand U3067 (N_3067,N_1991,N_2185);
nand U3068 (N_3068,N_1568,N_941);
nand U3069 (N_3069,N_2131,N_404);
or U3070 (N_3070,N_1912,N_341);
and U3071 (N_3071,N_1735,N_1543);
nor U3072 (N_3072,N_2174,N_973);
or U3073 (N_3073,N_1634,N_1758);
and U3074 (N_3074,N_1531,N_612);
nand U3075 (N_3075,N_903,N_1714);
or U3076 (N_3076,N_721,N_448);
and U3077 (N_3077,N_2342,N_1277);
nand U3078 (N_3078,N_1743,N_656);
and U3079 (N_3079,N_474,N_371);
nor U3080 (N_3080,N_954,N_2482);
or U3081 (N_3081,N_1265,N_68);
nor U3082 (N_3082,N_1829,N_111);
nor U3083 (N_3083,N_1556,N_1059);
nand U3084 (N_3084,N_1872,N_2204);
and U3085 (N_3085,N_1794,N_1038);
nand U3086 (N_3086,N_69,N_686);
nor U3087 (N_3087,N_501,N_1518);
nand U3088 (N_3088,N_890,N_1264);
or U3089 (N_3089,N_64,N_2114);
and U3090 (N_3090,N_120,N_1044);
nor U3091 (N_3091,N_1323,N_776);
nand U3092 (N_3092,N_2455,N_2197);
nand U3093 (N_3093,N_704,N_584);
and U3094 (N_3094,N_2472,N_335);
nand U3095 (N_3095,N_1307,N_1655);
or U3096 (N_3096,N_1296,N_1658);
or U3097 (N_3097,N_2149,N_765);
xnor U3098 (N_3098,N_1786,N_1424);
or U3099 (N_3099,N_1448,N_1538);
or U3100 (N_3100,N_1866,N_895);
or U3101 (N_3101,N_108,N_6);
and U3102 (N_3102,N_2419,N_1371);
nand U3103 (N_3103,N_123,N_1935);
nor U3104 (N_3104,N_2136,N_1601);
nor U3105 (N_3105,N_1110,N_169);
or U3106 (N_3106,N_2414,N_2080);
or U3107 (N_3107,N_2474,N_221);
nand U3108 (N_3108,N_396,N_1370);
or U3109 (N_3109,N_1685,N_2101);
or U3110 (N_3110,N_2128,N_2491);
nor U3111 (N_3111,N_904,N_2355);
nand U3112 (N_3112,N_200,N_348);
or U3113 (N_3113,N_723,N_1430);
nand U3114 (N_3114,N_2473,N_1364);
or U3115 (N_3115,N_948,N_2158);
and U3116 (N_3116,N_1922,N_2495);
and U3117 (N_3117,N_684,N_1989);
or U3118 (N_3118,N_2180,N_1486);
and U3119 (N_3119,N_188,N_2266);
and U3120 (N_3120,N_2064,N_302);
and U3121 (N_3121,N_606,N_218);
or U3122 (N_3122,N_187,N_993);
or U3123 (N_3123,N_1402,N_1826);
nand U3124 (N_3124,N_211,N_533);
or U3125 (N_3125,N_2292,N_294);
nand U3126 (N_3126,N_985,N_399);
and U3127 (N_3127,N_2442,N_1361);
nand U3128 (N_3128,N_225,N_846);
or U3129 (N_3129,N_1425,N_1012);
and U3130 (N_3130,N_734,N_345);
nand U3131 (N_3131,N_2089,N_390);
or U3132 (N_3132,N_2271,N_1346);
nand U3133 (N_3133,N_1224,N_1772);
nor U3134 (N_3134,N_1693,N_2401);
xnor U3135 (N_3135,N_46,N_2017);
and U3136 (N_3136,N_864,N_1010);
or U3137 (N_3137,N_1107,N_736);
or U3138 (N_3138,N_1419,N_2435);
and U3139 (N_3139,N_1321,N_493);
or U3140 (N_3140,N_2003,N_194);
and U3141 (N_3141,N_424,N_1832);
and U3142 (N_3142,N_2159,N_2273);
and U3143 (N_3143,N_1962,N_1437);
nand U3144 (N_3144,N_1828,N_710);
nand U3145 (N_3145,N_718,N_352);
or U3146 (N_3146,N_1707,N_125);
and U3147 (N_3147,N_615,N_697);
or U3148 (N_3148,N_62,N_1810);
nor U3149 (N_3149,N_519,N_577);
nor U3150 (N_3150,N_1624,N_1882);
nand U3151 (N_3151,N_818,N_2220);
nand U3152 (N_3152,N_2014,N_393);
or U3153 (N_3153,N_549,N_844);
and U3154 (N_3154,N_2290,N_931);
or U3155 (N_3155,N_2130,N_1611);
nand U3156 (N_3156,N_891,N_1491);
nor U3157 (N_3157,N_1981,N_2135);
or U3158 (N_3158,N_722,N_1754);
and U3159 (N_3159,N_1226,N_1862);
and U3160 (N_3160,N_164,N_1517);
nand U3161 (N_3161,N_1865,N_20);
or U3162 (N_3162,N_50,N_361);
or U3163 (N_3163,N_477,N_819);
nor U3164 (N_3164,N_1273,N_314);
and U3165 (N_3165,N_2183,N_2226);
nand U3166 (N_3166,N_1395,N_26);
and U3167 (N_3167,N_826,N_651);
and U3168 (N_3168,N_2223,N_1856);
and U3169 (N_3169,N_1198,N_2176);
nand U3170 (N_3170,N_2235,N_2297);
nor U3171 (N_3171,N_130,N_462);
and U3172 (N_3172,N_2047,N_996);
nor U3173 (N_3173,N_1120,N_741);
or U3174 (N_3174,N_1435,N_1153);
nor U3175 (N_3175,N_1697,N_1029);
or U3176 (N_3176,N_1931,N_2440);
and U3177 (N_3177,N_2178,N_2119);
nand U3178 (N_3178,N_410,N_1112);
nor U3179 (N_3179,N_1385,N_1418);
and U3180 (N_3180,N_1191,N_2045);
nor U3181 (N_3181,N_2209,N_1106);
nand U3182 (N_3182,N_596,N_227);
and U3183 (N_3183,N_1585,N_48);
and U3184 (N_3184,N_1510,N_310);
or U3185 (N_3185,N_1579,N_1879);
nor U3186 (N_3186,N_1275,N_753);
nand U3187 (N_3187,N_161,N_715);
nor U3188 (N_3188,N_54,N_1039);
xor U3189 (N_3189,N_1994,N_296);
and U3190 (N_3190,N_1421,N_95);
nor U3191 (N_3191,N_978,N_1447);
and U3192 (N_3192,N_956,N_2022);
or U3193 (N_3193,N_1297,N_2484);
or U3194 (N_3194,N_2302,N_349);
or U3195 (N_3195,N_425,N_987);
or U3196 (N_3196,N_575,N_255);
nand U3197 (N_3197,N_2168,N_705);
and U3198 (N_3198,N_224,N_1103);
and U3199 (N_3199,N_653,N_137);
and U3200 (N_3200,N_1901,N_1808);
or U3201 (N_3201,N_1605,N_845);
or U3202 (N_3202,N_1840,N_934);
or U3203 (N_3203,N_498,N_1467);
and U3204 (N_3204,N_526,N_1770);
or U3205 (N_3205,N_2335,N_278);
nor U3206 (N_3206,N_771,N_468);
and U3207 (N_3207,N_2433,N_867);
and U3208 (N_3208,N_1073,N_1963);
nand U3209 (N_3209,N_951,N_828);
nor U3210 (N_3210,N_2460,N_1228);
nand U3211 (N_3211,N_163,N_1627);
nand U3212 (N_3212,N_228,N_2373);
or U3213 (N_3213,N_2463,N_1800);
and U3214 (N_3214,N_1220,N_1004);
and U3215 (N_3215,N_1779,N_1677);
or U3216 (N_3216,N_885,N_1949);
or U3217 (N_3217,N_2084,N_1184);
and U3218 (N_3218,N_1782,N_1511);
or U3219 (N_3219,N_1390,N_2117);
nand U3220 (N_3220,N_1137,N_829);
nor U3221 (N_3221,N_494,N_1863);
nand U3222 (N_3222,N_1643,N_689);
or U3223 (N_3223,N_1728,N_49);
or U3224 (N_3224,N_81,N_1051);
xor U3225 (N_3225,N_1557,N_2034);
nand U3226 (N_3226,N_838,N_770);
or U3227 (N_3227,N_1396,N_649);
and U3228 (N_3228,N_1436,N_401);
and U3229 (N_3229,N_405,N_2275);
nand U3230 (N_3230,N_1186,N_2052);
and U3231 (N_3231,N_112,N_923);
and U3232 (N_3232,N_1030,N_589);
nor U3233 (N_3233,N_696,N_1194);
nor U3234 (N_3234,N_315,N_945);
or U3235 (N_3235,N_509,N_729);
and U3236 (N_3236,N_1417,N_782);
nand U3237 (N_3237,N_1860,N_2124);
and U3238 (N_3238,N_1146,N_952);
nand U3239 (N_3239,N_2049,N_967);
nand U3240 (N_3240,N_129,N_2269);
nand U3241 (N_3241,N_447,N_1329);
nor U3242 (N_3242,N_2329,N_134);
nand U3243 (N_3243,N_411,N_226);
nand U3244 (N_3244,N_1355,N_1621);
or U3245 (N_3245,N_131,N_1163);
nor U3246 (N_3246,N_798,N_1094);
and U3247 (N_3247,N_210,N_661);
or U3248 (N_3248,N_1813,N_1859);
and U3249 (N_3249,N_241,N_1730);
nand U3250 (N_3250,N_121,N_953);
and U3251 (N_3251,N_1667,N_1412);
nand U3252 (N_3252,N_1736,N_1148);
or U3253 (N_3253,N_1267,N_206);
and U3254 (N_3254,N_607,N_1035);
or U3255 (N_3255,N_1200,N_413);
and U3256 (N_3256,N_1636,N_974);
and U3257 (N_3257,N_1561,N_475);
nand U3258 (N_3258,N_2070,N_2383);
and U3259 (N_3259,N_2404,N_2012);
and U3260 (N_3260,N_1546,N_1656);
nor U3261 (N_3261,N_458,N_1242);
or U3262 (N_3262,N_13,N_1138);
or U3263 (N_3263,N_2421,N_31);
and U3264 (N_3264,N_376,N_713);
nand U3265 (N_3265,N_992,N_2040);
nor U3266 (N_3266,N_631,N_2251);
nand U3267 (N_3267,N_1848,N_439);
or U3268 (N_3268,N_1122,N_1996);
nand U3269 (N_3269,N_1341,N_2096);
nand U3270 (N_3270,N_881,N_1540);
and U3271 (N_3271,N_2115,N_2237);
nand U3272 (N_3272,N_1050,N_1592);
or U3273 (N_3273,N_2044,N_1542);
and U3274 (N_3274,N_1710,N_2466);
and U3275 (N_3275,N_1967,N_328);
nor U3276 (N_3276,N_1854,N_732);
or U3277 (N_3277,N_749,N_1288);
nand U3278 (N_3278,N_2248,N_2081);
nand U3279 (N_3279,N_1574,N_583);
nor U3280 (N_3280,N_1902,N_2356);
nor U3281 (N_3281,N_2188,N_578);
nand U3282 (N_3282,N_2300,N_1305);
nor U3283 (N_3283,N_1075,N_871);
nor U3284 (N_3284,N_1718,N_2104);
and U3285 (N_3285,N_132,N_2294);
nand U3286 (N_3286,N_9,N_785);
or U3287 (N_3287,N_2146,N_1790);
or U3288 (N_3288,N_888,N_1700);
nand U3289 (N_3289,N_1074,N_1833);
nand U3290 (N_3290,N_267,N_906);
and U3291 (N_3291,N_2099,N_2349);
nor U3292 (N_3292,N_918,N_2405);
or U3293 (N_3293,N_2145,N_641);
or U3294 (N_3294,N_204,N_822);
or U3295 (N_3295,N_2402,N_17);
or U3296 (N_3296,N_2065,N_7);
and U3297 (N_3297,N_1948,N_1202);
nand U3298 (N_3298,N_1855,N_16);
nor U3299 (N_3299,N_124,N_1298);
nand U3300 (N_3300,N_1313,N_706);
nor U3301 (N_3301,N_1196,N_1255);
or U3302 (N_3302,N_2140,N_690);
or U3303 (N_3303,N_1875,N_1575);
nor U3304 (N_3304,N_683,N_1932);
and U3305 (N_3305,N_1239,N_1006);
or U3306 (N_3306,N_1861,N_295);
nor U3307 (N_3307,N_182,N_104);
nand U3308 (N_3308,N_256,N_14);
nor U3309 (N_3309,N_236,N_479);
or U3310 (N_3310,N_1248,N_854);
nor U3311 (N_3311,N_1055,N_1924);
nor U3312 (N_3312,N_1629,N_1279);
nor U3313 (N_3313,N_622,N_117);
and U3314 (N_3314,N_1167,N_1088);
or U3315 (N_3315,N_2363,N_2259);
or U3316 (N_3316,N_1280,N_2350);
and U3317 (N_3317,N_611,N_687);
or U3318 (N_3318,N_1099,N_1898);
or U3319 (N_3319,N_2477,N_1619);
nand U3320 (N_3320,N_1111,N_1445);
or U3321 (N_3321,N_2125,N_761);
nand U3322 (N_3322,N_949,N_2316);
and U3323 (N_3323,N_834,N_2057);
or U3324 (N_3324,N_1129,N_8);
or U3325 (N_3325,N_764,N_353);
nor U3326 (N_3326,N_1954,N_1182);
xnor U3327 (N_3327,N_552,N_480);
and U3328 (N_3328,N_243,N_1550);
nand U3329 (N_3329,N_1376,N_184);
and U3330 (N_3330,N_1328,N_1889);
and U3331 (N_3331,N_457,N_1803);
and U3332 (N_3332,N_1132,N_2323);
nor U3333 (N_3333,N_15,N_2422);
nand U3334 (N_3334,N_1462,N_177);
and U3335 (N_3335,N_10,N_1097);
nand U3336 (N_3336,N_1128,N_717);
or U3337 (N_3337,N_1915,N_746);
or U3338 (N_3338,N_1339,N_412);
or U3339 (N_3339,N_1881,N_1485);
or U3340 (N_3340,N_1037,N_2365);
nor U3341 (N_3341,N_84,N_1208);
or U3342 (N_3342,N_1197,N_1853);
nor U3343 (N_3343,N_381,N_1519);
nand U3344 (N_3344,N_1282,N_2001);
nor U3345 (N_3345,N_1286,N_784);
nor U3346 (N_3346,N_525,N_2444);
nand U3347 (N_3347,N_1474,N_2055);
or U3348 (N_3348,N_1961,N_309);
and U3349 (N_3349,N_2074,N_1886);
nor U3350 (N_3350,N_1414,N_616);
nand U3351 (N_3351,N_159,N_197);
or U3352 (N_3352,N_1783,N_2389);
or U3353 (N_3353,N_1907,N_395);
or U3354 (N_3354,N_1720,N_354);
and U3355 (N_3355,N_2450,N_816);
nor U3356 (N_3356,N_880,N_1119);
and U3357 (N_3357,N_66,N_1450);
and U3358 (N_3358,N_913,N_1492);
and U3359 (N_3359,N_1407,N_2142);
nor U3360 (N_3360,N_1959,N_1811);
or U3361 (N_3361,N_1502,N_1217);
or U3362 (N_3362,N_190,N_2376);
nand U3363 (N_3363,N_994,N_154);
and U3364 (N_3364,N_1740,N_2328);
nor U3365 (N_3365,N_688,N_1174);
or U3366 (N_3366,N_285,N_2103);
nand U3367 (N_3367,N_1799,N_293);
and U3368 (N_3368,N_1489,N_805);
nand U3369 (N_3369,N_1484,N_503);
xor U3370 (N_3370,N_91,N_775);
nor U3371 (N_3371,N_670,N_437);
or U3372 (N_3372,N_2054,N_1367);
nand U3373 (N_3373,N_94,N_2212);
or U3374 (N_3374,N_1311,N_726);
or U3375 (N_3375,N_1943,N_2430);
or U3376 (N_3376,N_1207,N_355);
and U3377 (N_3377,N_2283,N_1746);
and U3378 (N_3378,N_2024,N_71);
or U3379 (N_3379,N_588,N_299);
or U3380 (N_3380,N_2416,N_1394);
nor U3381 (N_3381,N_1009,N_1921);
and U3382 (N_3382,N_1093,N_1822);
or U3383 (N_3383,N_158,N_1930);
nand U3384 (N_3384,N_289,N_2379);
and U3385 (N_3385,N_804,N_1013);
nand U3386 (N_3386,N_1576,N_912);
nand U3387 (N_3387,N_483,N_817);
and U3388 (N_3388,N_87,N_564);
nor U3389 (N_3389,N_2392,N_499);
or U3390 (N_3390,N_535,N_947);
and U3391 (N_3391,N_557,N_2284);
nand U3392 (N_3392,N_1969,N_1449);
and U3393 (N_3393,N_929,N_107);
nand U3394 (N_3394,N_1964,N_368);
nand U3395 (N_3395,N_1028,N_2072);
or U3396 (N_3396,N_2175,N_762);
nor U3397 (N_3397,N_198,N_379);
or U3398 (N_3398,N_1844,N_1905);
or U3399 (N_3399,N_1500,N_74);
or U3400 (N_3400,N_2048,N_1528);
or U3401 (N_3401,N_1375,N_1124);
and U3402 (N_3402,N_602,N_586);
nand U3403 (N_3403,N_2320,N_1042);
or U3404 (N_3404,N_504,N_153);
nand U3405 (N_3405,N_569,N_1253);
or U3406 (N_3406,N_2071,N_1613);
and U3407 (N_3407,N_1939,N_1284);
nor U3408 (N_3408,N_1271,N_1336);
nand U3409 (N_3409,N_1918,N_675);
nor U3410 (N_3410,N_1439,N_435);
nor U3411 (N_3411,N_1386,N_76);
or U3412 (N_3412,N_1034,N_1359);
or U3413 (N_3413,N_1526,N_1349);
nand U3414 (N_3414,N_2167,N_1062);
nor U3415 (N_3415,N_831,N_1987);
nand U3416 (N_3416,N_402,N_86);
nor U3417 (N_3417,N_1814,N_1731);
nor U3418 (N_3418,N_1534,N_2046);
or U3419 (N_3419,N_388,N_1733);
nand U3420 (N_3420,N_2486,N_655);
and U3421 (N_3421,N_321,N_22);
and U3422 (N_3422,N_11,N_1408);
or U3423 (N_3423,N_78,N_1460);
and U3424 (N_3424,N_1606,N_51);
nor U3425 (N_3425,N_1041,N_2334);
nand U3426 (N_3426,N_143,N_1117);
or U3427 (N_3427,N_1766,N_248);
nand U3428 (N_3428,N_1380,N_1053);
or U3429 (N_3429,N_1867,N_659);
nor U3430 (N_3430,N_2398,N_2397);
or U3431 (N_3431,N_2173,N_2412);
and U3432 (N_3432,N_1210,N_2050);
and U3433 (N_3433,N_1241,N_88);
and U3434 (N_3434,N_421,N_1204);
nor U3435 (N_3435,N_1413,N_2121);
nor U3436 (N_3436,N_2337,N_2352);
nand U3437 (N_3437,N_1514,N_1690);
nand U3438 (N_3438,N_691,N_1554);
nor U3439 (N_3439,N_274,N_1083);
nor U3440 (N_3440,N_541,N_1541);
and U3441 (N_3441,N_222,N_2031);
nand U3442 (N_3442,N_2457,N_701);
nor U3443 (N_3443,N_1512,N_546);
or U3444 (N_3444,N_857,N_1233);
and U3445 (N_3445,N_1000,N_109);
nor U3446 (N_3446,N_2261,N_2346);
nand U3447 (N_3447,N_1560,N_961);
nand U3448 (N_3448,N_1295,N_1415);
nor U3449 (N_3449,N_1957,N_1143);
nand U3450 (N_3450,N_1257,N_1644);
or U3451 (N_3451,N_2109,N_626);
nand U3452 (N_3452,N_702,N_1291);
and U3453 (N_3453,N_90,N_767);
nand U3454 (N_3454,N_1966,N_1071);
and U3455 (N_3455,N_1354,N_287);
nor U3456 (N_3456,N_356,N_2308);
nor U3457 (N_3457,N_1023,N_1509);
nand U3458 (N_3458,N_522,N_627);
nor U3459 (N_3459,N_2274,N_789);
nor U3460 (N_3460,N_2164,N_342);
and U3461 (N_3461,N_1348,N_2344);
or U3462 (N_3462,N_1043,N_414);
or U3463 (N_3463,N_1015,N_2306);
nand U3464 (N_3464,N_114,N_523);
nand U3465 (N_3465,N_2203,N_1147);
and U3466 (N_3466,N_1947,N_213);
and U3467 (N_3467,N_1544,N_542);
nor U3468 (N_3468,N_777,N_2206);
or U3469 (N_3469,N_92,N_2244);
nand U3470 (N_3470,N_2479,N_1076);
or U3471 (N_3471,N_2150,N_1640);
nor U3472 (N_3472,N_1260,N_795);
or U3473 (N_3473,N_530,N_167);
or U3474 (N_3474,N_933,N_2380);
nand U3475 (N_3475,N_1725,N_85);
or U3476 (N_3476,N_1304,N_681);
nor U3477 (N_3477,N_858,N_2331);
and U3478 (N_3478,N_742,N_2279);
nand U3479 (N_3479,N_1315,N_879);
nand U3480 (N_3480,N_1021,N_1444);
and U3481 (N_3481,N_262,N_2242);
nand U3482 (N_3482,N_1080,N_2179);
or U3483 (N_3483,N_47,N_2202);
or U3484 (N_3484,N_2200,N_209);
nor U3485 (N_3485,N_1352,N_1270);
and U3486 (N_3486,N_830,N_658);
or U3487 (N_3487,N_1807,N_720);
nand U3488 (N_3488,N_2215,N_2083);
nand U3489 (N_3489,N_157,N_1072);
nand U3490 (N_3490,N_2325,N_1232);
nor U3491 (N_3491,N_44,N_926);
nor U3492 (N_3492,N_1784,N_2362);
nand U3493 (N_3493,N_58,N_872);
nand U3494 (N_3494,N_202,N_407);
and U3495 (N_3495,N_1429,N_617);
nand U3496 (N_3496,N_693,N_168);
nand U3497 (N_3497,N_1851,N_1070);
nand U3498 (N_3498,N_944,N_1465);
or U3499 (N_3499,N_257,N_101);
nand U3500 (N_3500,N_284,N_1789);
nand U3501 (N_3501,N_781,N_1007);
nand U3502 (N_3502,N_2339,N_1470);
and U3503 (N_3503,N_2492,N_2144);
nand U3504 (N_3504,N_1469,N_1699);
nand U3505 (N_3505,N_579,N_1118);
nand U3506 (N_3506,N_774,N_889);
or U3507 (N_3507,N_1130,N_1446);
nor U3508 (N_3508,N_555,N_959);
or U3509 (N_3509,N_1381,N_711);
nor U3510 (N_3510,N_135,N_963);
nand U3511 (N_3511,N_362,N_1325);
and U3512 (N_3512,N_1567,N_1223);
or U3513 (N_3513,N_79,N_921);
or U3514 (N_3514,N_1084,N_37);
nor U3515 (N_3515,N_2291,N_969);
nand U3516 (N_3516,N_431,N_1876);
or U3517 (N_3517,N_343,N_556);
and U3518 (N_3518,N_1616,N_340);
and U3519 (N_3519,N_911,N_601);
nor U3520 (N_3520,N_573,N_1285);
and U3521 (N_3521,N_152,N_1259);
nor U3522 (N_3522,N_2090,N_1678);
or U3523 (N_3523,N_338,N_620);
or U3524 (N_3524,N_1652,N_593);
or U3525 (N_3525,N_699,N_1762);
and U3526 (N_3526,N_1166,N_2321);
nor U3527 (N_3527,N_471,N_100);
or U3528 (N_3528,N_1775,N_1768);
nor U3529 (N_3529,N_2361,N_320);
nor U3530 (N_3530,N_2143,N_271);
and U3531 (N_3531,N_1668,N_532);
and U3532 (N_3532,N_2016,N_1897);
and U3533 (N_3533,N_2116,N_1116);
nor U3534 (N_3534,N_1580,N_39);
nor U3535 (N_3535,N_2431,N_1098);
nor U3536 (N_3536,N_799,N_1631);
nor U3537 (N_3537,N_2061,N_1533);
nor U3538 (N_3538,N_2123,N_2336);
nor U3539 (N_3539,N_313,N_333);
and U3540 (N_3540,N_77,N_2148);
or U3541 (N_3541,N_432,N_1393);
nand U3542 (N_3542,N_1664,N_928);
nand U3543 (N_3543,N_1955,N_2393);
and U3544 (N_3544,N_1695,N_1069);
or U3545 (N_3545,N_1507,N_358);
or U3546 (N_3546,N_1916,N_849);
and U3547 (N_3547,N_654,N_2171);
nand U3548 (N_3548,N_2127,N_2133);
and U3549 (N_3549,N_1986,N_374);
nand U3550 (N_3550,N_2005,N_2078);
nor U3551 (N_3551,N_93,N_1428);
or U3552 (N_3552,N_1689,N_2006);
or U3553 (N_3553,N_763,N_1997);
nand U3554 (N_3554,N_1635,N_1032);
nor U3555 (N_3555,N_1183,N_183);
and U3556 (N_3556,N_2013,N_1020);
nor U3557 (N_3557,N_1780,N_740);
nor U3558 (N_3558,N_2333,N_1048);
and U3559 (N_3559,N_476,N_1463);
nand U3560 (N_3560,N_2161,N_442);
or U3561 (N_3561,N_1187,N_1798);
nand U3562 (N_3562,N_2301,N_217);
nand U3563 (N_3563,N_2053,N_1454);
and U3564 (N_3564,N_714,N_605);
or U3565 (N_3565,N_808,N_937);
and U3566 (N_3566,N_877,N_2067);
nand U3567 (N_3567,N_2347,N_841);
and U3568 (N_3568,N_128,N_1238);
nor U3569 (N_3569,N_570,N_1791);
nand U3570 (N_3570,N_1795,N_1990);
and U3571 (N_3571,N_1256,N_2488);
and U3572 (N_3572,N_1843,N_932);
and U3573 (N_3573,N_897,N_1975);
or U3574 (N_3574,N_628,N_591);
or U3575 (N_3575,N_1033,N_1302);
or U3576 (N_3576,N_980,N_1646);
nand U3577 (N_3577,N_2310,N_2322);
and U3578 (N_3578,N_1192,N_1008);
and U3579 (N_3579,N_635,N_444);
nand U3580 (N_3580,N_1113,N_660);
nand U3581 (N_3581,N_2439,N_216);
or U3582 (N_3582,N_1169,N_1243);
nand U3583 (N_3583,N_2387,N_886);
nand U3584 (N_3584,N_551,N_2438);
nor U3585 (N_3585,N_1178,N_2120);
and U3586 (N_3586,N_571,N_991);
nor U3587 (N_3587,N_1391,N_1442);
or U3588 (N_3588,N_1141,N_899);
or U3589 (N_3589,N_1374,N_449);
or U3590 (N_3590,N_1698,N_2);
nor U3591 (N_3591,N_1767,N_1389);
and U3592 (N_3592,N_1609,N_1373);
nand U3593 (N_3593,N_1090,N_2434);
or U3594 (N_3594,N_2020,N_1888);
nor U3595 (N_3595,N_2343,N_1249);
nor U3596 (N_3596,N_743,N_835);
xnor U3597 (N_3597,N_231,N_1596);
and U3598 (N_3598,N_290,N_1101);
xnor U3599 (N_3599,N_843,N_510);
and U3600 (N_3600,N_441,N_1165);
or U3601 (N_3601,N_1953,N_2367);
nand U3602 (N_3602,N_269,N_193);
nand U3603 (N_3603,N_1548,N_1377);
and U3604 (N_3604,N_2100,N_1705);
or U3605 (N_3605,N_2032,N_1459);
or U3606 (N_3606,N_446,N_759);
nor U3607 (N_3607,N_1488,N_738);
nor U3608 (N_3608,N_258,N_1040);
and U3609 (N_3609,N_1884,N_1706);
or U3610 (N_3610,N_1468,N_2381);
nand U3611 (N_3611,N_2219,N_2281);
or U3612 (N_3612,N_1936,N_839);
nand U3613 (N_3613,N_1410,N_1537);
or U3614 (N_3614,N_860,N_1711);
nor U3615 (N_3615,N_1164,N_1577);
or U3616 (N_3616,N_2285,N_150);
and U3617 (N_3617,N_265,N_2039);
nand U3618 (N_3618,N_1945,N_796);
and U3619 (N_3619,N_582,N_1477);
or U3620 (N_3620,N_1660,N_1893);
nand U3621 (N_3621,N_821,N_1300);
nand U3622 (N_3622,N_1404,N_984);
nand U3623 (N_3623,N_268,N_2088);
nor U3624 (N_3624,N_1797,N_1525);
and U3625 (N_3625,N_730,N_1142);
xnor U3626 (N_3626,N_768,N_1831);
nand U3627 (N_3627,N_2249,N_347);
nor U3628 (N_3628,N_1760,N_1688);
and U3629 (N_3629,N_1583,N_2287);
or U3630 (N_3630,N_576,N_2371);
or U3631 (N_3631,N_1661,N_1976);
and U3632 (N_3632,N_2160,N_305);
or U3633 (N_3633,N_2423,N_1388);
or U3634 (N_3634,N_550,N_592);
or U3635 (N_3635,N_727,N_1456);
or U3636 (N_3636,N_2360,N_1290);
or U3637 (N_3637,N_251,N_2447);
or U3638 (N_3638,N_2282,N_2162);
xnor U3639 (N_3639,N_2451,N_1880);
nor U3640 (N_3640,N_478,N_1406);
or U3641 (N_3641,N_2077,N_2341);
nor U3642 (N_3642,N_837,N_1552);
and U3643 (N_3643,N_1757,N_873);
nand U3644 (N_3644,N_1199,N_2068);
and U3645 (N_3645,N_1269,N_61);
and U3646 (N_3646,N_1443,N_712);
or U3647 (N_3647,N_812,N_1819);
or U3648 (N_3648,N_791,N_1569);
nor U3649 (N_3649,N_964,N_4);
and U3650 (N_3650,N_894,N_2066);
and U3651 (N_3651,N_1680,N_1675);
or U3652 (N_3652,N_2307,N_283);
or U3653 (N_3653,N_922,N_1229);
or U3654 (N_3654,N_1686,N_825);
or U3655 (N_3655,N_645,N_1058);
nor U3656 (N_3656,N_896,N_1586);
and U3657 (N_3657,N_788,N_2409);
or U3658 (N_3658,N_625,N_1669);
nor U3659 (N_3659,N_2403,N_1016);
nor U3660 (N_3660,N_1213,N_42);
and U3661 (N_3661,N_1268,N_2489);
or U3662 (N_3662,N_855,N_1672);
nor U3663 (N_3663,N_2277,N_2396);
nor U3664 (N_3664,N_1709,N_850);
nand U3665 (N_3665,N_1565,N_1595);
nor U3666 (N_3666,N_793,N_574);
and U3667 (N_3667,N_559,N_485);
nor U3668 (N_3668,N_2019,N_2126);
and U3669 (N_3669,N_1919,N_201);
or U3670 (N_3670,N_1984,N_1600);
or U3671 (N_3671,N_1312,N_367);
nor U3672 (N_3672,N_515,N_1588);
nor U3673 (N_3673,N_1334,N_146);
nand U3674 (N_3674,N_1522,N_118);
nor U3675 (N_3675,N_943,N_604);
and U3676 (N_3676,N_594,N_1778);
nor U3677 (N_3677,N_2445,N_1209);
or U3678 (N_3678,N_609,N_823);
or U3679 (N_3679,N_1818,N_646);
nor U3680 (N_3680,N_1154,N_384);
nor U3681 (N_3681,N_1508,N_669);
and U3682 (N_3682,N_1152,N_1114);
and U3683 (N_3683,N_2478,N_666);
and U3684 (N_3684,N_2288,N_418);
or U3685 (N_3685,N_1134,N_637);
nor U3686 (N_3686,N_558,N_1168);
and U3687 (N_3687,N_1501,N_861);
and U3688 (N_3688,N_2475,N_133);
xor U3689 (N_3689,N_1529,N_1432);
or U3690 (N_3690,N_43,N_2139);
and U3691 (N_3691,N_89,N_141);
nor U3692 (N_3692,N_2317,N_1551);
nor U3693 (N_3693,N_572,N_337);
or U3694 (N_3694,N_389,N_1654);
or U3695 (N_3695,N_2134,N_1159);
or U3696 (N_3696,N_1692,N_230);
nor U3697 (N_3697,N_567,N_440);
or U3698 (N_3698,N_1216,N_1372);
or U3699 (N_3699,N_2087,N_149);
and U3700 (N_3700,N_300,N_915);
nor U3701 (N_3701,N_1914,N_19);
nor U3702 (N_3702,N_238,N_1591);
or U3703 (N_3703,N_2228,N_1461);
nor U3704 (N_3704,N_232,N_1318);
xnor U3705 (N_3705,N_170,N_1911);
or U3706 (N_3706,N_1563,N_1081);
or U3707 (N_3707,N_472,N_1464);
or U3708 (N_3708,N_766,N_1904);
or U3709 (N_3709,N_1155,N_545);
and U3710 (N_3710,N_2009,N_815);
nand U3711 (N_3711,N_644,N_1324);
and U3712 (N_3712,N_205,N_716);
nor U3713 (N_3713,N_145,N_1250);
or U3714 (N_3714,N_1206,N_1457);
or U3715 (N_3715,N_2315,N_366);
or U3716 (N_3716,N_1712,N_610);
nand U3717 (N_3717,N_613,N_2234);
and U3718 (N_3718,N_473,N_2407);
nor U3719 (N_3719,N_2029,N_1726);
or U3720 (N_3720,N_176,N_2268);
or U3721 (N_3721,N_1343,N_281);
and U3722 (N_3722,N_2494,N_1247);
and U3723 (N_3723,N_965,N_465);
or U3724 (N_3724,N_415,N_1641);
and U3725 (N_3725,N_1816,N_2490);
nor U3726 (N_3726,N_350,N_1642);
nor U3727 (N_3727,N_1366,N_60);
or U3728 (N_3728,N_1719,N_2369);
or U3729 (N_3729,N_2151,N_2217);
nand U3730 (N_3730,N_1225,N_1095);
nor U3731 (N_3731,N_988,N_1869);
or U3732 (N_3732,N_1487,N_2424);
nor U3733 (N_3733,N_1158,N_1422);
and U3734 (N_3734,N_445,N_1539);
nor U3735 (N_3735,N_1382,N_1066);
nand U3736 (N_3736,N_110,N_1741);
and U3737 (N_3737,N_180,N_2138);
or U3738 (N_3738,N_908,N_481);
and U3739 (N_3739,N_773,N_1558);
or U3740 (N_3740,N_2184,N_1632);
nor U3741 (N_3741,N_809,N_2272);
or U3742 (N_3742,N_298,N_2097);
and U3743 (N_3743,N_597,N_181);
or U3744 (N_3744,N_2427,N_1189);
nand U3745 (N_3745,N_140,N_2385);
and U3746 (N_3746,N_1384,N_52);
and U3747 (N_3747,N_2058,N_883);
nor U3748 (N_3748,N_214,N_329);
or U3749 (N_3749,N_2106,N_2340);
nor U3750 (N_3750,N_1238,N_981);
nor U3751 (N_3751,N_2168,N_1743);
nand U3752 (N_3752,N_424,N_535);
nand U3753 (N_3753,N_407,N_1174);
or U3754 (N_3754,N_1644,N_500);
or U3755 (N_3755,N_2385,N_223);
or U3756 (N_3756,N_2349,N_1307);
nor U3757 (N_3757,N_2481,N_124);
or U3758 (N_3758,N_1218,N_1982);
nor U3759 (N_3759,N_2388,N_2138);
or U3760 (N_3760,N_1060,N_932);
nor U3761 (N_3761,N_277,N_1980);
nor U3762 (N_3762,N_1697,N_1558);
or U3763 (N_3763,N_1585,N_1951);
nor U3764 (N_3764,N_659,N_1875);
or U3765 (N_3765,N_2351,N_1940);
and U3766 (N_3766,N_1437,N_2126);
and U3767 (N_3767,N_1396,N_1303);
nand U3768 (N_3768,N_1353,N_1177);
or U3769 (N_3769,N_773,N_340);
nand U3770 (N_3770,N_255,N_509);
nand U3771 (N_3771,N_844,N_2247);
nor U3772 (N_3772,N_2142,N_1503);
nor U3773 (N_3773,N_1332,N_1093);
nor U3774 (N_3774,N_1089,N_122);
nor U3775 (N_3775,N_726,N_2446);
nand U3776 (N_3776,N_1902,N_1031);
nand U3777 (N_3777,N_484,N_2313);
nand U3778 (N_3778,N_2031,N_1914);
nor U3779 (N_3779,N_607,N_1369);
nand U3780 (N_3780,N_1175,N_1687);
or U3781 (N_3781,N_1235,N_707);
nor U3782 (N_3782,N_1469,N_13);
and U3783 (N_3783,N_276,N_2476);
or U3784 (N_3784,N_746,N_2480);
nor U3785 (N_3785,N_1725,N_469);
nand U3786 (N_3786,N_733,N_512);
nand U3787 (N_3787,N_846,N_756);
nor U3788 (N_3788,N_366,N_218);
nand U3789 (N_3789,N_2210,N_874);
or U3790 (N_3790,N_1234,N_1110);
nor U3791 (N_3791,N_1081,N_2019);
or U3792 (N_3792,N_92,N_214);
or U3793 (N_3793,N_1714,N_1769);
nor U3794 (N_3794,N_1132,N_403);
nor U3795 (N_3795,N_1577,N_2341);
nand U3796 (N_3796,N_193,N_848);
or U3797 (N_3797,N_1074,N_2046);
or U3798 (N_3798,N_1617,N_1575);
or U3799 (N_3799,N_1638,N_2408);
or U3800 (N_3800,N_571,N_899);
nand U3801 (N_3801,N_1713,N_2423);
nor U3802 (N_3802,N_661,N_113);
and U3803 (N_3803,N_1129,N_1674);
nor U3804 (N_3804,N_1831,N_1462);
and U3805 (N_3805,N_240,N_1085);
or U3806 (N_3806,N_1268,N_2158);
and U3807 (N_3807,N_2330,N_596);
nor U3808 (N_3808,N_943,N_785);
and U3809 (N_3809,N_815,N_2062);
and U3810 (N_3810,N_484,N_2477);
or U3811 (N_3811,N_404,N_1226);
or U3812 (N_3812,N_36,N_708);
nand U3813 (N_3813,N_1630,N_990);
xor U3814 (N_3814,N_1920,N_966);
nand U3815 (N_3815,N_1565,N_40);
xor U3816 (N_3816,N_369,N_2475);
nor U3817 (N_3817,N_2310,N_2108);
nand U3818 (N_3818,N_24,N_2046);
nand U3819 (N_3819,N_936,N_1984);
nor U3820 (N_3820,N_465,N_733);
and U3821 (N_3821,N_2440,N_2077);
nor U3822 (N_3822,N_467,N_301);
nor U3823 (N_3823,N_2090,N_252);
nand U3824 (N_3824,N_1531,N_2124);
nand U3825 (N_3825,N_407,N_1736);
nor U3826 (N_3826,N_2084,N_2378);
nand U3827 (N_3827,N_1220,N_1853);
and U3828 (N_3828,N_1454,N_569);
and U3829 (N_3829,N_1506,N_1296);
and U3830 (N_3830,N_1261,N_1489);
and U3831 (N_3831,N_945,N_548);
nor U3832 (N_3832,N_1937,N_534);
and U3833 (N_3833,N_1673,N_790);
nor U3834 (N_3834,N_226,N_462);
nor U3835 (N_3835,N_1691,N_2218);
and U3836 (N_3836,N_2388,N_2187);
nand U3837 (N_3837,N_1469,N_933);
and U3838 (N_3838,N_1437,N_1279);
or U3839 (N_3839,N_1069,N_2402);
nor U3840 (N_3840,N_1676,N_2216);
or U3841 (N_3841,N_893,N_333);
xor U3842 (N_3842,N_1508,N_2452);
nor U3843 (N_3843,N_1642,N_906);
or U3844 (N_3844,N_2011,N_1405);
nor U3845 (N_3845,N_2002,N_2495);
nor U3846 (N_3846,N_523,N_1257);
or U3847 (N_3847,N_256,N_1554);
and U3848 (N_3848,N_1348,N_2413);
and U3849 (N_3849,N_2136,N_2206);
nor U3850 (N_3850,N_620,N_1626);
or U3851 (N_3851,N_1163,N_2025);
nand U3852 (N_3852,N_1801,N_2453);
or U3853 (N_3853,N_2484,N_993);
nor U3854 (N_3854,N_253,N_1026);
nand U3855 (N_3855,N_46,N_2455);
or U3856 (N_3856,N_403,N_210);
nand U3857 (N_3857,N_305,N_1135);
nor U3858 (N_3858,N_488,N_1041);
and U3859 (N_3859,N_409,N_263);
nor U3860 (N_3860,N_1583,N_487);
or U3861 (N_3861,N_329,N_2426);
or U3862 (N_3862,N_2010,N_2397);
and U3863 (N_3863,N_383,N_2000);
or U3864 (N_3864,N_791,N_381);
nand U3865 (N_3865,N_937,N_1869);
nor U3866 (N_3866,N_650,N_1810);
nor U3867 (N_3867,N_1845,N_370);
and U3868 (N_3868,N_675,N_1473);
or U3869 (N_3869,N_602,N_1693);
or U3870 (N_3870,N_630,N_1454);
or U3871 (N_3871,N_667,N_1691);
or U3872 (N_3872,N_1845,N_1920);
or U3873 (N_3873,N_1164,N_544);
and U3874 (N_3874,N_790,N_1118);
nand U3875 (N_3875,N_620,N_1598);
nor U3876 (N_3876,N_790,N_2221);
nand U3877 (N_3877,N_1786,N_353);
nand U3878 (N_3878,N_343,N_1317);
or U3879 (N_3879,N_1707,N_164);
nand U3880 (N_3880,N_735,N_70);
nand U3881 (N_3881,N_893,N_980);
and U3882 (N_3882,N_291,N_1054);
or U3883 (N_3883,N_1923,N_1499);
xor U3884 (N_3884,N_2021,N_98);
and U3885 (N_3885,N_311,N_2318);
and U3886 (N_3886,N_2076,N_1091);
or U3887 (N_3887,N_1718,N_2318);
or U3888 (N_3888,N_677,N_2368);
and U3889 (N_3889,N_1382,N_91);
nand U3890 (N_3890,N_1365,N_2106);
or U3891 (N_3891,N_352,N_1693);
nand U3892 (N_3892,N_1373,N_741);
or U3893 (N_3893,N_24,N_1985);
or U3894 (N_3894,N_2341,N_2173);
nor U3895 (N_3895,N_795,N_2035);
nand U3896 (N_3896,N_1422,N_99);
or U3897 (N_3897,N_1680,N_1721);
nand U3898 (N_3898,N_412,N_378);
or U3899 (N_3899,N_1389,N_131);
nand U3900 (N_3900,N_1309,N_2141);
and U3901 (N_3901,N_134,N_334);
and U3902 (N_3902,N_884,N_863);
nor U3903 (N_3903,N_1735,N_300);
nand U3904 (N_3904,N_1198,N_882);
nor U3905 (N_3905,N_1012,N_403);
nand U3906 (N_3906,N_1382,N_640);
nor U3907 (N_3907,N_1288,N_360);
or U3908 (N_3908,N_702,N_557);
nand U3909 (N_3909,N_2068,N_1726);
or U3910 (N_3910,N_1341,N_2260);
and U3911 (N_3911,N_1949,N_1863);
nand U3912 (N_3912,N_581,N_190);
nand U3913 (N_3913,N_306,N_60);
or U3914 (N_3914,N_155,N_2128);
nor U3915 (N_3915,N_1610,N_1636);
and U3916 (N_3916,N_242,N_927);
or U3917 (N_3917,N_1842,N_398);
or U3918 (N_3918,N_2016,N_1154);
or U3919 (N_3919,N_1695,N_2470);
or U3920 (N_3920,N_444,N_109);
nor U3921 (N_3921,N_1916,N_589);
or U3922 (N_3922,N_1681,N_93);
nor U3923 (N_3923,N_2489,N_2424);
or U3924 (N_3924,N_2466,N_1751);
nand U3925 (N_3925,N_956,N_1906);
nand U3926 (N_3926,N_1005,N_2414);
or U3927 (N_3927,N_1767,N_1689);
or U3928 (N_3928,N_11,N_189);
and U3929 (N_3929,N_1113,N_70);
and U3930 (N_3930,N_1123,N_318);
and U3931 (N_3931,N_21,N_337);
and U3932 (N_3932,N_356,N_2342);
nand U3933 (N_3933,N_1396,N_132);
and U3934 (N_3934,N_1295,N_368);
nand U3935 (N_3935,N_1104,N_233);
and U3936 (N_3936,N_1561,N_1552);
and U3937 (N_3937,N_1207,N_2035);
xnor U3938 (N_3938,N_2146,N_2067);
or U3939 (N_3939,N_171,N_386);
or U3940 (N_3940,N_163,N_1353);
nand U3941 (N_3941,N_1292,N_1316);
and U3942 (N_3942,N_296,N_1625);
and U3943 (N_3943,N_2412,N_1335);
or U3944 (N_3944,N_192,N_1030);
or U3945 (N_3945,N_2058,N_1452);
or U3946 (N_3946,N_1088,N_2374);
nor U3947 (N_3947,N_1124,N_1224);
or U3948 (N_3948,N_1873,N_1757);
nor U3949 (N_3949,N_1599,N_1165);
and U3950 (N_3950,N_1385,N_1867);
and U3951 (N_3951,N_1956,N_2314);
or U3952 (N_3952,N_158,N_138);
or U3953 (N_3953,N_206,N_445);
nand U3954 (N_3954,N_2069,N_1141);
nor U3955 (N_3955,N_448,N_1381);
nand U3956 (N_3956,N_1805,N_1101);
and U3957 (N_3957,N_19,N_845);
and U3958 (N_3958,N_495,N_394);
nor U3959 (N_3959,N_1899,N_395);
nand U3960 (N_3960,N_2214,N_1782);
nor U3961 (N_3961,N_847,N_1277);
and U3962 (N_3962,N_1588,N_1827);
or U3963 (N_3963,N_698,N_2014);
or U3964 (N_3964,N_1001,N_2425);
or U3965 (N_3965,N_2229,N_1638);
or U3966 (N_3966,N_1284,N_439);
and U3967 (N_3967,N_1800,N_2462);
nand U3968 (N_3968,N_1615,N_1796);
or U3969 (N_3969,N_222,N_1084);
nor U3970 (N_3970,N_1792,N_2247);
nand U3971 (N_3971,N_1948,N_1737);
nand U3972 (N_3972,N_740,N_160);
or U3973 (N_3973,N_11,N_1429);
or U3974 (N_3974,N_448,N_1454);
nor U3975 (N_3975,N_1287,N_1913);
nor U3976 (N_3976,N_2489,N_298);
and U3977 (N_3977,N_1709,N_574);
nand U3978 (N_3978,N_1343,N_70);
and U3979 (N_3979,N_68,N_1980);
nand U3980 (N_3980,N_339,N_603);
and U3981 (N_3981,N_1301,N_2270);
nand U3982 (N_3982,N_1763,N_2236);
nand U3983 (N_3983,N_1234,N_2260);
and U3984 (N_3984,N_1996,N_16);
nor U3985 (N_3985,N_1907,N_983);
nand U3986 (N_3986,N_907,N_906);
nand U3987 (N_3987,N_1534,N_265);
or U3988 (N_3988,N_1771,N_1444);
and U3989 (N_3989,N_2227,N_1185);
or U3990 (N_3990,N_555,N_590);
nor U3991 (N_3991,N_1102,N_2361);
or U3992 (N_3992,N_1719,N_1210);
nand U3993 (N_3993,N_1256,N_1086);
nor U3994 (N_3994,N_1761,N_2314);
nand U3995 (N_3995,N_1404,N_481);
nand U3996 (N_3996,N_2476,N_259);
or U3997 (N_3997,N_2462,N_433);
nor U3998 (N_3998,N_137,N_570);
or U3999 (N_3999,N_922,N_916);
or U4000 (N_4000,N_2181,N_136);
or U4001 (N_4001,N_2091,N_2324);
and U4002 (N_4002,N_2261,N_2214);
or U4003 (N_4003,N_942,N_2321);
nand U4004 (N_4004,N_1888,N_620);
or U4005 (N_4005,N_1798,N_2427);
or U4006 (N_4006,N_369,N_2264);
or U4007 (N_4007,N_1939,N_1524);
and U4008 (N_4008,N_779,N_1970);
nor U4009 (N_4009,N_97,N_575);
nor U4010 (N_4010,N_2156,N_947);
nand U4011 (N_4011,N_2019,N_2219);
nor U4012 (N_4012,N_491,N_1665);
or U4013 (N_4013,N_2328,N_1668);
nor U4014 (N_4014,N_608,N_803);
nand U4015 (N_4015,N_1824,N_2406);
nand U4016 (N_4016,N_999,N_2110);
and U4017 (N_4017,N_145,N_1121);
or U4018 (N_4018,N_530,N_2097);
nand U4019 (N_4019,N_2252,N_178);
or U4020 (N_4020,N_1272,N_285);
and U4021 (N_4021,N_153,N_92);
or U4022 (N_4022,N_634,N_1601);
and U4023 (N_4023,N_493,N_1954);
nand U4024 (N_4024,N_1416,N_2027);
nand U4025 (N_4025,N_1278,N_2039);
nand U4026 (N_4026,N_654,N_1412);
and U4027 (N_4027,N_1245,N_2491);
nand U4028 (N_4028,N_1983,N_1000);
nand U4029 (N_4029,N_2070,N_1765);
or U4030 (N_4030,N_187,N_421);
and U4031 (N_4031,N_2358,N_268);
or U4032 (N_4032,N_2302,N_792);
and U4033 (N_4033,N_2302,N_382);
nand U4034 (N_4034,N_2081,N_1329);
and U4035 (N_4035,N_1269,N_1051);
or U4036 (N_4036,N_1831,N_1814);
nor U4037 (N_4037,N_903,N_1684);
nor U4038 (N_4038,N_2254,N_990);
and U4039 (N_4039,N_719,N_2347);
and U4040 (N_4040,N_561,N_579);
nand U4041 (N_4041,N_2250,N_1897);
nor U4042 (N_4042,N_1250,N_1860);
or U4043 (N_4043,N_1065,N_936);
nand U4044 (N_4044,N_2282,N_752);
xnor U4045 (N_4045,N_1102,N_1940);
and U4046 (N_4046,N_504,N_1044);
and U4047 (N_4047,N_1419,N_704);
or U4048 (N_4048,N_1251,N_1520);
or U4049 (N_4049,N_1759,N_548);
nand U4050 (N_4050,N_872,N_1178);
nor U4051 (N_4051,N_2363,N_191);
nand U4052 (N_4052,N_1820,N_1716);
and U4053 (N_4053,N_1443,N_261);
nand U4054 (N_4054,N_143,N_756);
nor U4055 (N_4055,N_381,N_1236);
nor U4056 (N_4056,N_858,N_2058);
nor U4057 (N_4057,N_351,N_853);
and U4058 (N_4058,N_1191,N_1827);
or U4059 (N_4059,N_506,N_1862);
or U4060 (N_4060,N_619,N_963);
nand U4061 (N_4061,N_1601,N_1964);
nor U4062 (N_4062,N_1865,N_130);
nand U4063 (N_4063,N_294,N_502);
nand U4064 (N_4064,N_1574,N_1962);
and U4065 (N_4065,N_289,N_1760);
nand U4066 (N_4066,N_1675,N_1842);
nand U4067 (N_4067,N_2003,N_2471);
nand U4068 (N_4068,N_1082,N_329);
or U4069 (N_4069,N_2343,N_2045);
or U4070 (N_4070,N_2299,N_249);
or U4071 (N_4071,N_882,N_736);
nor U4072 (N_4072,N_2429,N_92);
nand U4073 (N_4073,N_412,N_517);
nor U4074 (N_4074,N_298,N_1030);
nand U4075 (N_4075,N_1108,N_2262);
nor U4076 (N_4076,N_386,N_108);
and U4077 (N_4077,N_519,N_2433);
nor U4078 (N_4078,N_2458,N_1974);
nand U4079 (N_4079,N_2134,N_739);
nor U4080 (N_4080,N_527,N_277);
or U4081 (N_4081,N_863,N_463);
and U4082 (N_4082,N_1018,N_1241);
nand U4083 (N_4083,N_552,N_1070);
nor U4084 (N_4084,N_176,N_1366);
nor U4085 (N_4085,N_421,N_1036);
or U4086 (N_4086,N_2113,N_961);
xor U4087 (N_4087,N_1491,N_1856);
nor U4088 (N_4088,N_557,N_573);
nor U4089 (N_4089,N_527,N_1);
or U4090 (N_4090,N_281,N_1670);
nor U4091 (N_4091,N_2418,N_580);
nor U4092 (N_4092,N_674,N_964);
nor U4093 (N_4093,N_1606,N_544);
nand U4094 (N_4094,N_2224,N_178);
or U4095 (N_4095,N_496,N_31);
nor U4096 (N_4096,N_973,N_1957);
nand U4097 (N_4097,N_797,N_1969);
nand U4098 (N_4098,N_964,N_873);
and U4099 (N_4099,N_1050,N_851);
xnor U4100 (N_4100,N_55,N_1219);
xor U4101 (N_4101,N_270,N_917);
nand U4102 (N_4102,N_2392,N_14);
and U4103 (N_4103,N_450,N_2246);
or U4104 (N_4104,N_1877,N_718);
nor U4105 (N_4105,N_130,N_1905);
or U4106 (N_4106,N_1198,N_395);
or U4107 (N_4107,N_1399,N_2110);
nand U4108 (N_4108,N_1274,N_873);
or U4109 (N_4109,N_1435,N_895);
nand U4110 (N_4110,N_285,N_1618);
nor U4111 (N_4111,N_2479,N_2209);
or U4112 (N_4112,N_1777,N_621);
nand U4113 (N_4113,N_90,N_2494);
or U4114 (N_4114,N_1048,N_285);
or U4115 (N_4115,N_2095,N_1256);
and U4116 (N_4116,N_1414,N_1226);
and U4117 (N_4117,N_2431,N_1980);
and U4118 (N_4118,N_100,N_2335);
and U4119 (N_4119,N_1031,N_461);
nand U4120 (N_4120,N_405,N_2227);
nor U4121 (N_4121,N_1369,N_76);
nand U4122 (N_4122,N_347,N_914);
and U4123 (N_4123,N_2037,N_1002);
nor U4124 (N_4124,N_1501,N_1230);
and U4125 (N_4125,N_2151,N_1570);
nor U4126 (N_4126,N_652,N_841);
nor U4127 (N_4127,N_1674,N_49);
and U4128 (N_4128,N_2249,N_835);
nand U4129 (N_4129,N_1269,N_2447);
and U4130 (N_4130,N_1308,N_142);
and U4131 (N_4131,N_670,N_2440);
nand U4132 (N_4132,N_2354,N_2060);
and U4133 (N_4133,N_2433,N_71);
nand U4134 (N_4134,N_1193,N_852);
nand U4135 (N_4135,N_2347,N_2098);
or U4136 (N_4136,N_503,N_771);
nor U4137 (N_4137,N_1698,N_248);
xor U4138 (N_4138,N_125,N_998);
and U4139 (N_4139,N_2291,N_1905);
or U4140 (N_4140,N_2262,N_2374);
nor U4141 (N_4141,N_19,N_795);
nor U4142 (N_4142,N_1203,N_2198);
nor U4143 (N_4143,N_92,N_1062);
or U4144 (N_4144,N_770,N_1762);
and U4145 (N_4145,N_1448,N_272);
nor U4146 (N_4146,N_2216,N_875);
nor U4147 (N_4147,N_1946,N_395);
nor U4148 (N_4148,N_1819,N_1997);
or U4149 (N_4149,N_1031,N_2336);
or U4150 (N_4150,N_345,N_1587);
nor U4151 (N_4151,N_2393,N_639);
nor U4152 (N_4152,N_438,N_878);
or U4153 (N_4153,N_2038,N_1612);
nor U4154 (N_4154,N_397,N_585);
and U4155 (N_4155,N_1693,N_573);
or U4156 (N_4156,N_1157,N_1255);
or U4157 (N_4157,N_2231,N_2243);
or U4158 (N_4158,N_2196,N_133);
or U4159 (N_4159,N_900,N_2333);
and U4160 (N_4160,N_886,N_772);
nand U4161 (N_4161,N_659,N_1862);
and U4162 (N_4162,N_2076,N_400);
or U4163 (N_4163,N_1773,N_962);
and U4164 (N_4164,N_1804,N_2447);
or U4165 (N_4165,N_1886,N_1351);
nand U4166 (N_4166,N_2178,N_1844);
or U4167 (N_4167,N_121,N_2068);
or U4168 (N_4168,N_388,N_1512);
nand U4169 (N_4169,N_250,N_1102);
nand U4170 (N_4170,N_1036,N_1203);
or U4171 (N_4171,N_812,N_598);
and U4172 (N_4172,N_1289,N_1768);
or U4173 (N_4173,N_67,N_267);
nor U4174 (N_4174,N_1439,N_2397);
nand U4175 (N_4175,N_229,N_2415);
or U4176 (N_4176,N_775,N_2327);
nand U4177 (N_4177,N_446,N_1185);
or U4178 (N_4178,N_971,N_579);
and U4179 (N_4179,N_2466,N_514);
nand U4180 (N_4180,N_2044,N_685);
nor U4181 (N_4181,N_725,N_1707);
nor U4182 (N_4182,N_2351,N_560);
nor U4183 (N_4183,N_1703,N_1442);
or U4184 (N_4184,N_118,N_630);
or U4185 (N_4185,N_1613,N_872);
and U4186 (N_4186,N_971,N_1239);
and U4187 (N_4187,N_943,N_1009);
nand U4188 (N_4188,N_1951,N_67);
nand U4189 (N_4189,N_1518,N_175);
and U4190 (N_4190,N_847,N_584);
nor U4191 (N_4191,N_40,N_990);
or U4192 (N_4192,N_2490,N_1143);
nand U4193 (N_4193,N_1141,N_2436);
or U4194 (N_4194,N_891,N_2484);
or U4195 (N_4195,N_2103,N_2443);
nand U4196 (N_4196,N_2359,N_1219);
and U4197 (N_4197,N_1335,N_84);
nor U4198 (N_4198,N_746,N_1571);
or U4199 (N_4199,N_2319,N_518);
or U4200 (N_4200,N_590,N_1161);
or U4201 (N_4201,N_961,N_1432);
or U4202 (N_4202,N_1469,N_976);
or U4203 (N_4203,N_1784,N_955);
nor U4204 (N_4204,N_2211,N_212);
nor U4205 (N_4205,N_1206,N_2060);
or U4206 (N_4206,N_1552,N_2197);
nand U4207 (N_4207,N_2381,N_2090);
nand U4208 (N_4208,N_2059,N_65);
nand U4209 (N_4209,N_2368,N_2331);
nand U4210 (N_4210,N_1422,N_1819);
or U4211 (N_4211,N_1402,N_480);
or U4212 (N_4212,N_2057,N_656);
and U4213 (N_4213,N_1842,N_2418);
and U4214 (N_4214,N_2333,N_1428);
and U4215 (N_4215,N_1887,N_2335);
and U4216 (N_4216,N_829,N_862);
nor U4217 (N_4217,N_2132,N_249);
and U4218 (N_4218,N_867,N_877);
and U4219 (N_4219,N_2264,N_2159);
and U4220 (N_4220,N_1096,N_1001);
or U4221 (N_4221,N_1068,N_1225);
or U4222 (N_4222,N_254,N_1633);
nand U4223 (N_4223,N_554,N_1233);
and U4224 (N_4224,N_1641,N_189);
nor U4225 (N_4225,N_2151,N_2027);
and U4226 (N_4226,N_2116,N_358);
nor U4227 (N_4227,N_1775,N_1853);
nand U4228 (N_4228,N_2475,N_1096);
xnor U4229 (N_4229,N_1178,N_1050);
nor U4230 (N_4230,N_1099,N_1844);
and U4231 (N_4231,N_1776,N_995);
and U4232 (N_4232,N_1140,N_2366);
and U4233 (N_4233,N_2387,N_2236);
nand U4234 (N_4234,N_621,N_1748);
nor U4235 (N_4235,N_2017,N_1903);
or U4236 (N_4236,N_66,N_1115);
and U4237 (N_4237,N_430,N_1710);
nor U4238 (N_4238,N_2042,N_2374);
and U4239 (N_4239,N_667,N_154);
and U4240 (N_4240,N_80,N_1764);
nor U4241 (N_4241,N_677,N_2034);
nor U4242 (N_4242,N_2459,N_125);
or U4243 (N_4243,N_1755,N_1362);
or U4244 (N_4244,N_1558,N_2091);
nor U4245 (N_4245,N_2020,N_1809);
nor U4246 (N_4246,N_109,N_4);
nor U4247 (N_4247,N_1331,N_1092);
and U4248 (N_4248,N_1743,N_2470);
nor U4249 (N_4249,N_721,N_2242);
xnor U4250 (N_4250,N_2449,N_294);
and U4251 (N_4251,N_402,N_2123);
or U4252 (N_4252,N_224,N_1981);
nor U4253 (N_4253,N_1979,N_1639);
or U4254 (N_4254,N_1843,N_2275);
or U4255 (N_4255,N_939,N_68);
xor U4256 (N_4256,N_1935,N_1475);
nor U4257 (N_4257,N_1316,N_482);
nand U4258 (N_4258,N_809,N_1195);
nand U4259 (N_4259,N_1992,N_2007);
or U4260 (N_4260,N_2107,N_825);
nor U4261 (N_4261,N_135,N_339);
or U4262 (N_4262,N_2155,N_2194);
or U4263 (N_4263,N_1149,N_2176);
and U4264 (N_4264,N_555,N_2397);
nor U4265 (N_4265,N_18,N_825);
nor U4266 (N_4266,N_798,N_2355);
nand U4267 (N_4267,N_551,N_1895);
and U4268 (N_4268,N_2323,N_122);
nor U4269 (N_4269,N_331,N_574);
nor U4270 (N_4270,N_1484,N_1090);
and U4271 (N_4271,N_1636,N_1832);
nand U4272 (N_4272,N_1666,N_2018);
nor U4273 (N_4273,N_314,N_626);
and U4274 (N_4274,N_2430,N_1739);
nor U4275 (N_4275,N_1734,N_825);
or U4276 (N_4276,N_916,N_1216);
nand U4277 (N_4277,N_1167,N_638);
nand U4278 (N_4278,N_758,N_2008);
nor U4279 (N_4279,N_2468,N_484);
and U4280 (N_4280,N_669,N_488);
nor U4281 (N_4281,N_783,N_2275);
nand U4282 (N_4282,N_2087,N_77);
or U4283 (N_4283,N_808,N_1745);
or U4284 (N_4284,N_1114,N_173);
nand U4285 (N_4285,N_1512,N_665);
nand U4286 (N_4286,N_685,N_2070);
nor U4287 (N_4287,N_1914,N_1016);
nor U4288 (N_4288,N_368,N_38);
or U4289 (N_4289,N_793,N_1693);
or U4290 (N_4290,N_2487,N_797);
nand U4291 (N_4291,N_166,N_334);
nor U4292 (N_4292,N_108,N_1882);
or U4293 (N_4293,N_1660,N_2342);
nor U4294 (N_4294,N_191,N_897);
nor U4295 (N_4295,N_2277,N_2307);
nor U4296 (N_4296,N_173,N_196);
nor U4297 (N_4297,N_1163,N_1095);
or U4298 (N_4298,N_1900,N_320);
nor U4299 (N_4299,N_2454,N_1500);
nor U4300 (N_4300,N_721,N_2150);
or U4301 (N_4301,N_560,N_1486);
nand U4302 (N_4302,N_265,N_1719);
nand U4303 (N_4303,N_1200,N_1911);
or U4304 (N_4304,N_754,N_1);
or U4305 (N_4305,N_2380,N_1608);
or U4306 (N_4306,N_1833,N_548);
and U4307 (N_4307,N_1506,N_1690);
or U4308 (N_4308,N_841,N_1211);
nand U4309 (N_4309,N_1654,N_1666);
nor U4310 (N_4310,N_1494,N_477);
nand U4311 (N_4311,N_422,N_758);
nand U4312 (N_4312,N_1905,N_1566);
and U4313 (N_4313,N_1332,N_301);
and U4314 (N_4314,N_2364,N_1609);
nor U4315 (N_4315,N_323,N_30);
nor U4316 (N_4316,N_741,N_472);
or U4317 (N_4317,N_406,N_1566);
or U4318 (N_4318,N_1320,N_1311);
or U4319 (N_4319,N_2045,N_1695);
and U4320 (N_4320,N_1087,N_331);
nand U4321 (N_4321,N_1140,N_1817);
nand U4322 (N_4322,N_1148,N_1407);
or U4323 (N_4323,N_1639,N_2364);
nor U4324 (N_4324,N_2255,N_43);
or U4325 (N_4325,N_1713,N_1087);
nor U4326 (N_4326,N_359,N_1619);
or U4327 (N_4327,N_2134,N_1590);
and U4328 (N_4328,N_2257,N_774);
and U4329 (N_4329,N_161,N_2447);
nand U4330 (N_4330,N_2002,N_10);
nand U4331 (N_4331,N_2427,N_1569);
and U4332 (N_4332,N_61,N_1591);
or U4333 (N_4333,N_1246,N_223);
and U4334 (N_4334,N_1611,N_2183);
nor U4335 (N_4335,N_520,N_1756);
or U4336 (N_4336,N_458,N_1495);
and U4337 (N_4337,N_266,N_1455);
nor U4338 (N_4338,N_1053,N_586);
or U4339 (N_4339,N_1298,N_1196);
nor U4340 (N_4340,N_1971,N_844);
and U4341 (N_4341,N_1053,N_734);
and U4342 (N_4342,N_1680,N_2152);
nor U4343 (N_4343,N_2272,N_348);
nand U4344 (N_4344,N_224,N_1616);
nor U4345 (N_4345,N_2404,N_1228);
and U4346 (N_4346,N_1387,N_1120);
nor U4347 (N_4347,N_351,N_2241);
and U4348 (N_4348,N_885,N_168);
nand U4349 (N_4349,N_1331,N_1619);
or U4350 (N_4350,N_866,N_2013);
nor U4351 (N_4351,N_966,N_452);
nor U4352 (N_4352,N_104,N_2201);
or U4353 (N_4353,N_1528,N_2037);
or U4354 (N_4354,N_427,N_1367);
or U4355 (N_4355,N_103,N_370);
nand U4356 (N_4356,N_2260,N_138);
nor U4357 (N_4357,N_568,N_1586);
nor U4358 (N_4358,N_1881,N_487);
or U4359 (N_4359,N_2135,N_462);
and U4360 (N_4360,N_1261,N_148);
nor U4361 (N_4361,N_1594,N_1636);
or U4362 (N_4362,N_1630,N_231);
nand U4363 (N_4363,N_1219,N_1584);
nand U4364 (N_4364,N_225,N_944);
nor U4365 (N_4365,N_2189,N_1173);
and U4366 (N_4366,N_2343,N_130);
nor U4367 (N_4367,N_1774,N_2253);
nand U4368 (N_4368,N_1767,N_1665);
or U4369 (N_4369,N_516,N_1401);
nor U4370 (N_4370,N_2237,N_1580);
or U4371 (N_4371,N_1223,N_1187);
nor U4372 (N_4372,N_206,N_633);
and U4373 (N_4373,N_532,N_1915);
or U4374 (N_4374,N_2184,N_1364);
or U4375 (N_4375,N_1353,N_2137);
and U4376 (N_4376,N_2113,N_2432);
nand U4377 (N_4377,N_978,N_1811);
nand U4378 (N_4378,N_2439,N_2258);
nor U4379 (N_4379,N_873,N_2176);
nand U4380 (N_4380,N_912,N_111);
or U4381 (N_4381,N_1616,N_1138);
nor U4382 (N_4382,N_2423,N_634);
or U4383 (N_4383,N_2324,N_784);
nand U4384 (N_4384,N_1599,N_2373);
nor U4385 (N_4385,N_1451,N_1784);
or U4386 (N_4386,N_1360,N_1412);
or U4387 (N_4387,N_1590,N_1795);
or U4388 (N_4388,N_832,N_2288);
and U4389 (N_4389,N_627,N_1671);
nand U4390 (N_4390,N_1242,N_1901);
and U4391 (N_4391,N_1985,N_2420);
and U4392 (N_4392,N_2120,N_577);
nand U4393 (N_4393,N_1088,N_423);
nor U4394 (N_4394,N_59,N_4);
and U4395 (N_4395,N_499,N_2133);
or U4396 (N_4396,N_2080,N_298);
and U4397 (N_4397,N_2476,N_356);
nor U4398 (N_4398,N_213,N_236);
nor U4399 (N_4399,N_580,N_1971);
nand U4400 (N_4400,N_2347,N_2160);
nand U4401 (N_4401,N_1178,N_1292);
or U4402 (N_4402,N_961,N_1520);
nand U4403 (N_4403,N_2158,N_2180);
nor U4404 (N_4404,N_1072,N_1938);
nor U4405 (N_4405,N_2249,N_1525);
and U4406 (N_4406,N_332,N_1767);
nor U4407 (N_4407,N_190,N_146);
nand U4408 (N_4408,N_539,N_333);
or U4409 (N_4409,N_2107,N_56);
or U4410 (N_4410,N_2304,N_1527);
and U4411 (N_4411,N_674,N_109);
and U4412 (N_4412,N_2208,N_2441);
nor U4413 (N_4413,N_129,N_791);
and U4414 (N_4414,N_1824,N_1073);
and U4415 (N_4415,N_1194,N_2400);
and U4416 (N_4416,N_1754,N_1494);
nand U4417 (N_4417,N_2383,N_712);
xor U4418 (N_4418,N_2309,N_1660);
and U4419 (N_4419,N_1501,N_1892);
or U4420 (N_4420,N_358,N_321);
nand U4421 (N_4421,N_1554,N_1480);
and U4422 (N_4422,N_992,N_2153);
and U4423 (N_4423,N_2021,N_219);
nor U4424 (N_4424,N_1162,N_400);
nor U4425 (N_4425,N_1725,N_2482);
and U4426 (N_4426,N_2449,N_265);
nand U4427 (N_4427,N_2212,N_757);
or U4428 (N_4428,N_1994,N_1622);
nand U4429 (N_4429,N_1759,N_1243);
and U4430 (N_4430,N_268,N_2373);
nand U4431 (N_4431,N_671,N_912);
nand U4432 (N_4432,N_2089,N_26);
xor U4433 (N_4433,N_1625,N_838);
nand U4434 (N_4434,N_491,N_688);
and U4435 (N_4435,N_1902,N_2467);
nor U4436 (N_4436,N_551,N_717);
and U4437 (N_4437,N_1337,N_2169);
nor U4438 (N_4438,N_2289,N_1270);
nor U4439 (N_4439,N_1368,N_619);
or U4440 (N_4440,N_406,N_645);
or U4441 (N_4441,N_595,N_1372);
or U4442 (N_4442,N_658,N_1836);
nor U4443 (N_4443,N_859,N_930);
nor U4444 (N_4444,N_2200,N_1780);
or U4445 (N_4445,N_782,N_304);
nor U4446 (N_4446,N_551,N_1212);
and U4447 (N_4447,N_1798,N_1764);
or U4448 (N_4448,N_93,N_1187);
and U4449 (N_4449,N_1507,N_86);
and U4450 (N_4450,N_1428,N_2060);
or U4451 (N_4451,N_1890,N_517);
nand U4452 (N_4452,N_1788,N_406);
nand U4453 (N_4453,N_456,N_445);
and U4454 (N_4454,N_839,N_1544);
nand U4455 (N_4455,N_1988,N_450);
or U4456 (N_4456,N_1624,N_1704);
or U4457 (N_4457,N_1275,N_2025);
and U4458 (N_4458,N_2224,N_423);
nor U4459 (N_4459,N_967,N_1129);
nand U4460 (N_4460,N_2394,N_786);
and U4461 (N_4461,N_882,N_248);
xnor U4462 (N_4462,N_355,N_517);
and U4463 (N_4463,N_1576,N_1449);
nor U4464 (N_4464,N_921,N_938);
and U4465 (N_4465,N_1388,N_118);
or U4466 (N_4466,N_1639,N_496);
and U4467 (N_4467,N_352,N_1550);
nand U4468 (N_4468,N_1390,N_1535);
nand U4469 (N_4469,N_331,N_949);
and U4470 (N_4470,N_1908,N_1194);
nor U4471 (N_4471,N_1116,N_2457);
nor U4472 (N_4472,N_534,N_708);
and U4473 (N_4473,N_1495,N_841);
nor U4474 (N_4474,N_231,N_2456);
nor U4475 (N_4475,N_585,N_549);
nor U4476 (N_4476,N_1031,N_2310);
and U4477 (N_4477,N_453,N_23);
or U4478 (N_4478,N_464,N_799);
nand U4479 (N_4479,N_1749,N_895);
or U4480 (N_4480,N_48,N_1357);
or U4481 (N_4481,N_1449,N_287);
or U4482 (N_4482,N_685,N_2361);
or U4483 (N_4483,N_1569,N_2414);
nor U4484 (N_4484,N_2140,N_2020);
nand U4485 (N_4485,N_838,N_747);
nand U4486 (N_4486,N_915,N_1021);
nor U4487 (N_4487,N_392,N_2244);
nor U4488 (N_4488,N_2400,N_2211);
nand U4489 (N_4489,N_924,N_2344);
and U4490 (N_4490,N_1058,N_1283);
and U4491 (N_4491,N_1019,N_2077);
nand U4492 (N_4492,N_475,N_1259);
and U4493 (N_4493,N_1046,N_518);
and U4494 (N_4494,N_1513,N_265);
or U4495 (N_4495,N_1273,N_792);
or U4496 (N_4496,N_2146,N_239);
or U4497 (N_4497,N_2433,N_1653);
nand U4498 (N_4498,N_2280,N_2424);
and U4499 (N_4499,N_151,N_2007);
and U4500 (N_4500,N_1881,N_2488);
nand U4501 (N_4501,N_1451,N_2270);
nor U4502 (N_4502,N_1213,N_12);
and U4503 (N_4503,N_2074,N_2338);
nor U4504 (N_4504,N_750,N_2005);
nand U4505 (N_4505,N_476,N_221);
or U4506 (N_4506,N_1327,N_2008);
or U4507 (N_4507,N_638,N_577);
and U4508 (N_4508,N_1609,N_1311);
nand U4509 (N_4509,N_1590,N_832);
and U4510 (N_4510,N_2265,N_792);
nor U4511 (N_4511,N_5,N_178);
nand U4512 (N_4512,N_2244,N_1015);
or U4513 (N_4513,N_697,N_2122);
nor U4514 (N_4514,N_867,N_2233);
or U4515 (N_4515,N_330,N_701);
and U4516 (N_4516,N_99,N_2066);
or U4517 (N_4517,N_1372,N_5);
nor U4518 (N_4518,N_1932,N_1360);
nor U4519 (N_4519,N_2109,N_1926);
nor U4520 (N_4520,N_934,N_966);
nor U4521 (N_4521,N_247,N_453);
and U4522 (N_4522,N_1721,N_2306);
nand U4523 (N_4523,N_1738,N_762);
nand U4524 (N_4524,N_1127,N_2447);
and U4525 (N_4525,N_2384,N_863);
and U4526 (N_4526,N_2423,N_143);
and U4527 (N_4527,N_2029,N_764);
or U4528 (N_4528,N_741,N_708);
nand U4529 (N_4529,N_68,N_2234);
or U4530 (N_4530,N_1393,N_130);
nand U4531 (N_4531,N_1829,N_1214);
and U4532 (N_4532,N_993,N_59);
and U4533 (N_4533,N_2441,N_1207);
and U4534 (N_4534,N_1446,N_655);
nand U4535 (N_4535,N_2488,N_2047);
nor U4536 (N_4536,N_1519,N_2252);
and U4537 (N_4537,N_1829,N_901);
nor U4538 (N_4538,N_2343,N_175);
and U4539 (N_4539,N_1446,N_1555);
nor U4540 (N_4540,N_45,N_460);
nor U4541 (N_4541,N_1496,N_584);
and U4542 (N_4542,N_2267,N_2338);
or U4543 (N_4543,N_202,N_128);
nor U4544 (N_4544,N_1241,N_1246);
nor U4545 (N_4545,N_1357,N_58);
and U4546 (N_4546,N_422,N_1176);
nor U4547 (N_4547,N_959,N_2408);
and U4548 (N_4548,N_1056,N_2128);
and U4549 (N_4549,N_1437,N_989);
nand U4550 (N_4550,N_752,N_1965);
nor U4551 (N_4551,N_1685,N_1413);
nand U4552 (N_4552,N_1329,N_1036);
nor U4553 (N_4553,N_1988,N_1623);
or U4554 (N_4554,N_2137,N_1939);
nor U4555 (N_4555,N_568,N_63);
nor U4556 (N_4556,N_2278,N_1927);
nand U4557 (N_4557,N_2333,N_1607);
nand U4558 (N_4558,N_1965,N_2423);
nor U4559 (N_4559,N_376,N_2129);
or U4560 (N_4560,N_949,N_1292);
or U4561 (N_4561,N_1301,N_1027);
or U4562 (N_4562,N_528,N_1032);
nand U4563 (N_4563,N_2250,N_1712);
nand U4564 (N_4564,N_29,N_1817);
or U4565 (N_4565,N_1702,N_1327);
or U4566 (N_4566,N_1770,N_158);
or U4567 (N_4567,N_2061,N_2071);
nand U4568 (N_4568,N_680,N_2440);
and U4569 (N_4569,N_1285,N_1342);
nand U4570 (N_4570,N_965,N_692);
and U4571 (N_4571,N_1050,N_1544);
and U4572 (N_4572,N_1040,N_2479);
nor U4573 (N_4573,N_669,N_1046);
and U4574 (N_4574,N_950,N_1587);
nand U4575 (N_4575,N_1643,N_974);
nand U4576 (N_4576,N_160,N_1677);
or U4577 (N_4577,N_1291,N_1107);
xnor U4578 (N_4578,N_1167,N_2071);
xnor U4579 (N_4579,N_376,N_419);
nor U4580 (N_4580,N_2400,N_2338);
and U4581 (N_4581,N_1831,N_786);
and U4582 (N_4582,N_1958,N_2125);
nand U4583 (N_4583,N_538,N_2203);
nand U4584 (N_4584,N_646,N_1787);
and U4585 (N_4585,N_1661,N_2329);
or U4586 (N_4586,N_127,N_554);
or U4587 (N_4587,N_188,N_1352);
and U4588 (N_4588,N_434,N_952);
or U4589 (N_4589,N_2251,N_1026);
or U4590 (N_4590,N_606,N_2426);
or U4591 (N_4591,N_1267,N_2090);
xor U4592 (N_4592,N_76,N_2142);
or U4593 (N_4593,N_2035,N_1109);
or U4594 (N_4594,N_946,N_51);
or U4595 (N_4595,N_445,N_1108);
or U4596 (N_4596,N_1118,N_2480);
nand U4597 (N_4597,N_1254,N_2224);
or U4598 (N_4598,N_2168,N_1740);
nor U4599 (N_4599,N_1848,N_1621);
nor U4600 (N_4600,N_484,N_1735);
nand U4601 (N_4601,N_2280,N_1747);
or U4602 (N_4602,N_999,N_691);
or U4603 (N_4603,N_1155,N_2157);
nand U4604 (N_4604,N_1926,N_1711);
and U4605 (N_4605,N_196,N_1747);
or U4606 (N_4606,N_2445,N_58);
or U4607 (N_4607,N_288,N_1378);
nand U4608 (N_4608,N_2466,N_2349);
or U4609 (N_4609,N_1139,N_1782);
nand U4610 (N_4610,N_623,N_536);
nand U4611 (N_4611,N_2316,N_461);
nand U4612 (N_4612,N_1016,N_2470);
nand U4613 (N_4613,N_553,N_1952);
or U4614 (N_4614,N_1649,N_1922);
nor U4615 (N_4615,N_507,N_553);
and U4616 (N_4616,N_1825,N_2194);
and U4617 (N_4617,N_1166,N_395);
nor U4618 (N_4618,N_123,N_827);
nand U4619 (N_4619,N_806,N_752);
nand U4620 (N_4620,N_620,N_408);
or U4621 (N_4621,N_2423,N_1112);
and U4622 (N_4622,N_1176,N_2484);
and U4623 (N_4623,N_2160,N_2124);
nand U4624 (N_4624,N_4,N_1026);
nor U4625 (N_4625,N_828,N_1686);
nand U4626 (N_4626,N_1211,N_355);
and U4627 (N_4627,N_626,N_163);
nand U4628 (N_4628,N_2019,N_1661);
nand U4629 (N_4629,N_1574,N_1845);
and U4630 (N_4630,N_672,N_1667);
and U4631 (N_4631,N_34,N_893);
and U4632 (N_4632,N_642,N_289);
and U4633 (N_4633,N_527,N_1131);
nor U4634 (N_4634,N_1368,N_881);
or U4635 (N_4635,N_773,N_1075);
nand U4636 (N_4636,N_1147,N_1164);
nor U4637 (N_4637,N_1334,N_355);
or U4638 (N_4638,N_2456,N_886);
nor U4639 (N_4639,N_2440,N_1654);
nand U4640 (N_4640,N_2084,N_1330);
nor U4641 (N_4641,N_802,N_1991);
or U4642 (N_4642,N_1932,N_706);
nor U4643 (N_4643,N_1888,N_2363);
and U4644 (N_4644,N_637,N_749);
and U4645 (N_4645,N_2380,N_956);
and U4646 (N_4646,N_1254,N_1046);
xnor U4647 (N_4647,N_2495,N_2192);
nor U4648 (N_4648,N_1717,N_2298);
or U4649 (N_4649,N_474,N_745);
and U4650 (N_4650,N_297,N_2354);
nor U4651 (N_4651,N_166,N_24);
nor U4652 (N_4652,N_881,N_1102);
and U4653 (N_4653,N_475,N_1468);
and U4654 (N_4654,N_795,N_1176);
nand U4655 (N_4655,N_1590,N_82);
nor U4656 (N_4656,N_71,N_355);
nand U4657 (N_4657,N_1019,N_2182);
and U4658 (N_4658,N_2022,N_150);
or U4659 (N_4659,N_1443,N_2008);
or U4660 (N_4660,N_2188,N_272);
nor U4661 (N_4661,N_1792,N_1624);
nand U4662 (N_4662,N_2025,N_1270);
and U4663 (N_4663,N_1087,N_830);
and U4664 (N_4664,N_1470,N_2092);
or U4665 (N_4665,N_314,N_1930);
and U4666 (N_4666,N_459,N_682);
nor U4667 (N_4667,N_2489,N_288);
nand U4668 (N_4668,N_910,N_252);
nor U4669 (N_4669,N_1029,N_277);
nand U4670 (N_4670,N_156,N_1447);
nand U4671 (N_4671,N_1197,N_925);
nor U4672 (N_4672,N_1827,N_1475);
nor U4673 (N_4673,N_2021,N_2465);
and U4674 (N_4674,N_31,N_1904);
or U4675 (N_4675,N_2021,N_81);
or U4676 (N_4676,N_226,N_28);
nor U4677 (N_4677,N_691,N_908);
and U4678 (N_4678,N_233,N_2198);
and U4679 (N_4679,N_491,N_542);
or U4680 (N_4680,N_2455,N_110);
xor U4681 (N_4681,N_2483,N_755);
or U4682 (N_4682,N_241,N_1110);
or U4683 (N_4683,N_1442,N_223);
nand U4684 (N_4684,N_1830,N_1898);
and U4685 (N_4685,N_692,N_1430);
nor U4686 (N_4686,N_2109,N_68);
or U4687 (N_4687,N_1309,N_2190);
and U4688 (N_4688,N_1773,N_515);
nand U4689 (N_4689,N_1606,N_2283);
and U4690 (N_4690,N_1244,N_311);
and U4691 (N_4691,N_260,N_2178);
and U4692 (N_4692,N_1656,N_2305);
and U4693 (N_4693,N_1763,N_608);
nand U4694 (N_4694,N_1347,N_646);
nor U4695 (N_4695,N_297,N_699);
and U4696 (N_4696,N_2123,N_2387);
nor U4697 (N_4697,N_241,N_419);
nand U4698 (N_4698,N_207,N_1537);
nor U4699 (N_4699,N_684,N_1407);
and U4700 (N_4700,N_1220,N_171);
or U4701 (N_4701,N_870,N_955);
and U4702 (N_4702,N_1710,N_2369);
and U4703 (N_4703,N_1315,N_2255);
and U4704 (N_4704,N_1868,N_1032);
and U4705 (N_4705,N_316,N_758);
nor U4706 (N_4706,N_818,N_1255);
nand U4707 (N_4707,N_2181,N_2419);
or U4708 (N_4708,N_527,N_977);
nor U4709 (N_4709,N_486,N_872);
and U4710 (N_4710,N_1879,N_614);
nor U4711 (N_4711,N_1668,N_281);
or U4712 (N_4712,N_574,N_97);
or U4713 (N_4713,N_128,N_1444);
or U4714 (N_4714,N_265,N_706);
nand U4715 (N_4715,N_2187,N_302);
or U4716 (N_4716,N_2108,N_643);
or U4717 (N_4717,N_725,N_509);
nor U4718 (N_4718,N_1758,N_2319);
and U4719 (N_4719,N_244,N_598);
or U4720 (N_4720,N_984,N_2355);
or U4721 (N_4721,N_1157,N_153);
and U4722 (N_4722,N_1897,N_1968);
or U4723 (N_4723,N_643,N_120);
nand U4724 (N_4724,N_2480,N_919);
and U4725 (N_4725,N_1240,N_1916);
nand U4726 (N_4726,N_2260,N_876);
nand U4727 (N_4727,N_1504,N_981);
or U4728 (N_4728,N_388,N_190);
nand U4729 (N_4729,N_506,N_887);
nand U4730 (N_4730,N_87,N_819);
or U4731 (N_4731,N_1049,N_2435);
nand U4732 (N_4732,N_342,N_984);
or U4733 (N_4733,N_806,N_166);
nand U4734 (N_4734,N_770,N_477);
nand U4735 (N_4735,N_1115,N_854);
or U4736 (N_4736,N_982,N_1470);
nand U4737 (N_4737,N_374,N_1274);
nand U4738 (N_4738,N_663,N_976);
or U4739 (N_4739,N_2259,N_1631);
and U4740 (N_4740,N_1066,N_601);
nor U4741 (N_4741,N_316,N_1194);
nand U4742 (N_4742,N_2368,N_93);
nor U4743 (N_4743,N_1177,N_155);
or U4744 (N_4744,N_2463,N_1561);
nand U4745 (N_4745,N_1993,N_2481);
nand U4746 (N_4746,N_1746,N_778);
or U4747 (N_4747,N_2420,N_1275);
nand U4748 (N_4748,N_1398,N_1837);
nor U4749 (N_4749,N_1234,N_838);
and U4750 (N_4750,N_758,N_1946);
or U4751 (N_4751,N_791,N_449);
nand U4752 (N_4752,N_114,N_18);
and U4753 (N_4753,N_1525,N_1562);
nor U4754 (N_4754,N_794,N_600);
nand U4755 (N_4755,N_2352,N_696);
and U4756 (N_4756,N_2138,N_253);
nand U4757 (N_4757,N_1883,N_1793);
or U4758 (N_4758,N_44,N_809);
or U4759 (N_4759,N_1703,N_1211);
nor U4760 (N_4760,N_958,N_1881);
and U4761 (N_4761,N_1560,N_1906);
and U4762 (N_4762,N_2038,N_1871);
nand U4763 (N_4763,N_1136,N_1912);
nor U4764 (N_4764,N_1836,N_45);
nor U4765 (N_4765,N_422,N_1129);
or U4766 (N_4766,N_2450,N_556);
nor U4767 (N_4767,N_717,N_1940);
nand U4768 (N_4768,N_1022,N_665);
and U4769 (N_4769,N_93,N_1194);
and U4770 (N_4770,N_520,N_80);
nand U4771 (N_4771,N_1694,N_1214);
and U4772 (N_4772,N_1749,N_952);
and U4773 (N_4773,N_1956,N_1552);
nand U4774 (N_4774,N_1281,N_1400);
or U4775 (N_4775,N_536,N_177);
nor U4776 (N_4776,N_1242,N_1662);
nand U4777 (N_4777,N_2127,N_1153);
or U4778 (N_4778,N_2234,N_854);
or U4779 (N_4779,N_2436,N_1901);
and U4780 (N_4780,N_903,N_2200);
nand U4781 (N_4781,N_1548,N_1573);
or U4782 (N_4782,N_1281,N_2286);
nor U4783 (N_4783,N_826,N_1746);
nand U4784 (N_4784,N_938,N_2495);
and U4785 (N_4785,N_1413,N_1465);
or U4786 (N_4786,N_2469,N_709);
nor U4787 (N_4787,N_1504,N_1283);
and U4788 (N_4788,N_154,N_1198);
and U4789 (N_4789,N_255,N_774);
and U4790 (N_4790,N_2104,N_107);
or U4791 (N_4791,N_1489,N_743);
and U4792 (N_4792,N_1078,N_2423);
or U4793 (N_4793,N_332,N_866);
or U4794 (N_4794,N_2322,N_1878);
or U4795 (N_4795,N_453,N_264);
and U4796 (N_4796,N_563,N_2227);
nand U4797 (N_4797,N_1067,N_1697);
nor U4798 (N_4798,N_603,N_621);
or U4799 (N_4799,N_1677,N_2408);
or U4800 (N_4800,N_1207,N_1066);
and U4801 (N_4801,N_1840,N_895);
nor U4802 (N_4802,N_1393,N_369);
nand U4803 (N_4803,N_925,N_104);
nor U4804 (N_4804,N_53,N_1401);
and U4805 (N_4805,N_1326,N_224);
or U4806 (N_4806,N_348,N_198);
or U4807 (N_4807,N_2417,N_1620);
or U4808 (N_4808,N_2034,N_397);
and U4809 (N_4809,N_1320,N_637);
and U4810 (N_4810,N_1597,N_1886);
and U4811 (N_4811,N_2157,N_187);
nand U4812 (N_4812,N_1152,N_177);
nand U4813 (N_4813,N_1864,N_1649);
nand U4814 (N_4814,N_1180,N_2128);
nand U4815 (N_4815,N_1496,N_1378);
and U4816 (N_4816,N_764,N_1383);
or U4817 (N_4817,N_1845,N_1239);
nor U4818 (N_4818,N_758,N_1622);
nor U4819 (N_4819,N_2375,N_1673);
nor U4820 (N_4820,N_2366,N_1925);
nor U4821 (N_4821,N_449,N_2042);
and U4822 (N_4822,N_1273,N_1899);
or U4823 (N_4823,N_1784,N_542);
or U4824 (N_4824,N_1956,N_422);
nand U4825 (N_4825,N_1795,N_153);
and U4826 (N_4826,N_2383,N_526);
nand U4827 (N_4827,N_325,N_1428);
nor U4828 (N_4828,N_2037,N_2082);
and U4829 (N_4829,N_1826,N_2131);
or U4830 (N_4830,N_1591,N_490);
nor U4831 (N_4831,N_1576,N_1605);
and U4832 (N_4832,N_177,N_1115);
nand U4833 (N_4833,N_324,N_664);
or U4834 (N_4834,N_911,N_2087);
and U4835 (N_4835,N_1823,N_1411);
and U4836 (N_4836,N_1015,N_414);
and U4837 (N_4837,N_1687,N_1856);
or U4838 (N_4838,N_934,N_1821);
and U4839 (N_4839,N_1683,N_2428);
nor U4840 (N_4840,N_2192,N_1090);
nand U4841 (N_4841,N_1996,N_1968);
and U4842 (N_4842,N_1031,N_2089);
and U4843 (N_4843,N_343,N_865);
or U4844 (N_4844,N_243,N_2138);
xnor U4845 (N_4845,N_2091,N_1449);
nor U4846 (N_4846,N_2378,N_2262);
nor U4847 (N_4847,N_1979,N_1955);
nor U4848 (N_4848,N_1535,N_1216);
or U4849 (N_4849,N_733,N_658);
nor U4850 (N_4850,N_429,N_1139);
or U4851 (N_4851,N_1234,N_1977);
or U4852 (N_4852,N_1394,N_1235);
and U4853 (N_4853,N_1725,N_2419);
and U4854 (N_4854,N_31,N_38);
and U4855 (N_4855,N_2207,N_92);
or U4856 (N_4856,N_2397,N_1547);
or U4857 (N_4857,N_115,N_1659);
and U4858 (N_4858,N_1660,N_1976);
nand U4859 (N_4859,N_2242,N_1299);
nand U4860 (N_4860,N_1978,N_2362);
or U4861 (N_4861,N_1335,N_1998);
or U4862 (N_4862,N_1483,N_579);
nor U4863 (N_4863,N_75,N_2354);
or U4864 (N_4864,N_1975,N_1617);
and U4865 (N_4865,N_1490,N_1294);
nand U4866 (N_4866,N_270,N_509);
and U4867 (N_4867,N_1881,N_2496);
or U4868 (N_4868,N_519,N_1689);
and U4869 (N_4869,N_867,N_405);
and U4870 (N_4870,N_917,N_1884);
nand U4871 (N_4871,N_886,N_749);
nand U4872 (N_4872,N_504,N_697);
or U4873 (N_4873,N_2035,N_2155);
and U4874 (N_4874,N_2083,N_276);
or U4875 (N_4875,N_2034,N_1437);
and U4876 (N_4876,N_1257,N_797);
nand U4877 (N_4877,N_1612,N_1006);
or U4878 (N_4878,N_932,N_1655);
or U4879 (N_4879,N_362,N_26);
nand U4880 (N_4880,N_2033,N_1579);
and U4881 (N_4881,N_1637,N_1210);
or U4882 (N_4882,N_2239,N_451);
nand U4883 (N_4883,N_1265,N_1610);
nor U4884 (N_4884,N_1597,N_329);
nand U4885 (N_4885,N_400,N_2414);
nand U4886 (N_4886,N_300,N_74);
nor U4887 (N_4887,N_1585,N_1089);
nor U4888 (N_4888,N_1239,N_865);
xnor U4889 (N_4889,N_2178,N_2084);
and U4890 (N_4890,N_263,N_1431);
nor U4891 (N_4891,N_2465,N_1632);
and U4892 (N_4892,N_833,N_1746);
nor U4893 (N_4893,N_1948,N_1685);
and U4894 (N_4894,N_1696,N_1564);
xnor U4895 (N_4895,N_189,N_153);
or U4896 (N_4896,N_352,N_542);
or U4897 (N_4897,N_2468,N_2);
nand U4898 (N_4898,N_2227,N_1160);
or U4899 (N_4899,N_866,N_1452);
nand U4900 (N_4900,N_1524,N_1807);
or U4901 (N_4901,N_652,N_1083);
nor U4902 (N_4902,N_1716,N_2205);
nor U4903 (N_4903,N_760,N_990);
or U4904 (N_4904,N_2420,N_390);
nand U4905 (N_4905,N_2439,N_921);
or U4906 (N_4906,N_823,N_1220);
or U4907 (N_4907,N_1649,N_2128);
nor U4908 (N_4908,N_15,N_1150);
or U4909 (N_4909,N_1214,N_511);
nor U4910 (N_4910,N_701,N_2232);
nor U4911 (N_4911,N_161,N_364);
nor U4912 (N_4912,N_2416,N_2424);
nor U4913 (N_4913,N_1735,N_1485);
nand U4914 (N_4914,N_2476,N_549);
nor U4915 (N_4915,N_1401,N_1557);
or U4916 (N_4916,N_971,N_1874);
and U4917 (N_4917,N_1299,N_1314);
nand U4918 (N_4918,N_2139,N_1144);
nand U4919 (N_4919,N_631,N_1911);
nand U4920 (N_4920,N_1695,N_203);
and U4921 (N_4921,N_1397,N_665);
nand U4922 (N_4922,N_1165,N_2130);
and U4923 (N_4923,N_933,N_1666);
and U4924 (N_4924,N_170,N_1957);
xnor U4925 (N_4925,N_1294,N_1582);
nand U4926 (N_4926,N_1560,N_1579);
and U4927 (N_4927,N_817,N_1796);
nor U4928 (N_4928,N_34,N_2178);
or U4929 (N_4929,N_811,N_906);
nand U4930 (N_4930,N_324,N_546);
nand U4931 (N_4931,N_190,N_477);
or U4932 (N_4932,N_1028,N_1661);
or U4933 (N_4933,N_1950,N_1338);
and U4934 (N_4934,N_1490,N_1266);
nor U4935 (N_4935,N_488,N_1490);
nor U4936 (N_4936,N_2202,N_336);
nor U4937 (N_4937,N_1633,N_30);
or U4938 (N_4938,N_2296,N_876);
and U4939 (N_4939,N_2063,N_222);
nor U4940 (N_4940,N_2196,N_1239);
nand U4941 (N_4941,N_2289,N_2089);
or U4942 (N_4942,N_2043,N_1630);
and U4943 (N_4943,N_2244,N_2394);
and U4944 (N_4944,N_1932,N_1523);
or U4945 (N_4945,N_1938,N_1980);
or U4946 (N_4946,N_2230,N_1354);
nand U4947 (N_4947,N_863,N_539);
and U4948 (N_4948,N_2023,N_475);
or U4949 (N_4949,N_886,N_209);
or U4950 (N_4950,N_254,N_2187);
or U4951 (N_4951,N_1928,N_410);
nor U4952 (N_4952,N_966,N_589);
and U4953 (N_4953,N_24,N_1623);
nand U4954 (N_4954,N_1264,N_1694);
nor U4955 (N_4955,N_2309,N_2389);
or U4956 (N_4956,N_2076,N_2);
and U4957 (N_4957,N_1084,N_391);
and U4958 (N_4958,N_2056,N_1907);
and U4959 (N_4959,N_890,N_127);
nor U4960 (N_4960,N_437,N_2027);
nor U4961 (N_4961,N_1079,N_1175);
nor U4962 (N_4962,N_1268,N_1335);
nor U4963 (N_4963,N_384,N_2434);
or U4964 (N_4964,N_1735,N_1293);
and U4965 (N_4965,N_2461,N_850);
nor U4966 (N_4966,N_1296,N_2372);
nor U4967 (N_4967,N_2327,N_563);
and U4968 (N_4968,N_515,N_260);
xor U4969 (N_4969,N_366,N_975);
and U4970 (N_4970,N_1038,N_1654);
nand U4971 (N_4971,N_256,N_712);
or U4972 (N_4972,N_1815,N_1146);
nor U4973 (N_4973,N_2365,N_246);
nand U4974 (N_4974,N_1434,N_2132);
or U4975 (N_4975,N_2301,N_1821);
or U4976 (N_4976,N_1254,N_106);
and U4977 (N_4977,N_1474,N_1358);
nand U4978 (N_4978,N_2459,N_1080);
nand U4979 (N_4979,N_1272,N_2099);
nand U4980 (N_4980,N_1341,N_904);
or U4981 (N_4981,N_412,N_1486);
nand U4982 (N_4982,N_326,N_2140);
and U4983 (N_4983,N_757,N_2178);
and U4984 (N_4984,N_1106,N_2206);
nor U4985 (N_4985,N_1680,N_1984);
and U4986 (N_4986,N_82,N_881);
and U4987 (N_4987,N_1383,N_121);
and U4988 (N_4988,N_1741,N_1712);
nand U4989 (N_4989,N_470,N_625);
nor U4990 (N_4990,N_2,N_1746);
or U4991 (N_4991,N_1206,N_2027);
or U4992 (N_4992,N_791,N_379);
nand U4993 (N_4993,N_1736,N_2485);
nor U4994 (N_4994,N_549,N_2458);
nor U4995 (N_4995,N_1100,N_2233);
and U4996 (N_4996,N_1842,N_143);
or U4997 (N_4997,N_2441,N_1268);
nor U4998 (N_4998,N_745,N_1612);
nor U4999 (N_4999,N_1879,N_1628);
nand U5000 (N_5000,N_4804,N_2877);
nor U5001 (N_5001,N_4707,N_2593);
or U5002 (N_5002,N_4339,N_3257);
and U5003 (N_5003,N_4004,N_4485);
and U5004 (N_5004,N_3059,N_2873);
or U5005 (N_5005,N_4686,N_3160);
nor U5006 (N_5006,N_3451,N_3134);
nor U5007 (N_5007,N_2733,N_4308);
or U5008 (N_5008,N_3899,N_3590);
or U5009 (N_5009,N_2532,N_4952);
nor U5010 (N_5010,N_4653,N_3910);
nand U5011 (N_5011,N_4948,N_3981);
nor U5012 (N_5012,N_4394,N_3487);
nor U5013 (N_5013,N_4608,N_4412);
and U5014 (N_5014,N_3378,N_4060);
and U5015 (N_5015,N_4774,N_3064);
nor U5016 (N_5016,N_3815,N_2756);
or U5017 (N_5017,N_3669,N_4328);
nor U5018 (N_5018,N_4275,N_2770);
nand U5019 (N_5019,N_4118,N_3017);
and U5020 (N_5020,N_4041,N_4187);
nand U5021 (N_5021,N_4139,N_4518);
or U5022 (N_5022,N_4365,N_4972);
or U5023 (N_5023,N_4334,N_2922);
or U5024 (N_5024,N_3356,N_2902);
and U5025 (N_5025,N_2856,N_4907);
nand U5026 (N_5026,N_4613,N_3866);
nor U5027 (N_5027,N_4129,N_4807);
and U5028 (N_5028,N_4197,N_2546);
nand U5029 (N_5029,N_3148,N_3438);
nand U5030 (N_5030,N_4536,N_3222);
or U5031 (N_5031,N_3801,N_4370);
or U5032 (N_5032,N_3284,N_3410);
and U5033 (N_5033,N_4045,N_4356);
or U5034 (N_5034,N_4325,N_3407);
or U5035 (N_5035,N_2618,N_4940);
nand U5036 (N_5036,N_4759,N_4199);
nand U5037 (N_5037,N_2614,N_4243);
and U5038 (N_5038,N_4017,N_3977);
and U5039 (N_5039,N_3693,N_4285);
nand U5040 (N_5040,N_4306,N_4319);
or U5041 (N_5041,N_4315,N_3103);
or U5042 (N_5042,N_3250,N_3730);
or U5043 (N_5043,N_4383,N_2883);
and U5044 (N_5044,N_4542,N_2526);
or U5045 (N_5045,N_3542,N_4450);
nor U5046 (N_5046,N_3515,N_4871);
nor U5047 (N_5047,N_4223,N_4161);
and U5048 (N_5048,N_3945,N_3979);
nand U5049 (N_5049,N_2505,N_2884);
and U5050 (N_5050,N_4027,N_3950);
and U5051 (N_5051,N_4254,N_4090);
nor U5052 (N_5052,N_4321,N_3599);
or U5053 (N_5053,N_4215,N_3420);
nor U5054 (N_5054,N_4028,N_4996);
nor U5055 (N_5055,N_4337,N_3985);
or U5056 (N_5056,N_3644,N_3167);
nand U5057 (N_5057,N_3227,N_4358);
nor U5058 (N_5058,N_2829,N_4494);
nand U5059 (N_5059,N_4368,N_3499);
nand U5060 (N_5060,N_4722,N_3359);
nand U5061 (N_5061,N_3226,N_2631);
or U5062 (N_5062,N_4258,N_4206);
and U5063 (N_5063,N_4249,N_3992);
and U5064 (N_5064,N_4549,N_3835);
or U5065 (N_5065,N_2609,N_3741);
nor U5066 (N_5066,N_3965,N_4892);
nor U5067 (N_5067,N_2938,N_3791);
nor U5068 (N_5068,N_3010,N_2875);
nand U5069 (N_5069,N_2857,N_3204);
and U5070 (N_5070,N_4371,N_4976);
and U5071 (N_5071,N_4760,N_3102);
and U5072 (N_5072,N_3675,N_3849);
and U5073 (N_5073,N_3154,N_3474);
and U5074 (N_5074,N_3129,N_2662);
or U5075 (N_5075,N_2723,N_3221);
nor U5076 (N_5076,N_4550,N_4880);
and U5077 (N_5077,N_2792,N_4135);
nor U5078 (N_5078,N_3933,N_3347);
xnor U5079 (N_5079,N_3296,N_4583);
nand U5080 (N_5080,N_2894,N_4569);
nor U5081 (N_5081,N_4640,N_4154);
nor U5082 (N_5082,N_4283,N_3539);
and U5083 (N_5083,N_4826,N_4253);
and U5084 (N_5084,N_3271,N_3900);
nor U5085 (N_5085,N_4828,N_3655);
or U5086 (N_5086,N_3829,N_4240);
and U5087 (N_5087,N_3367,N_2850);
nand U5088 (N_5088,N_3351,N_4934);
and U5089 (N_5089,N_4734,N_4675);
nor U5090 (N_5090,N_4629,N_3365);
nor U5091 (N_5091,N_3259,N_2879);
and U5092 (N_5092,N_4967,N_4464);
or U5093 (N_5093,N_4172,N_3810);
or U5094 (N_5094,N_4516,N_4474);
nor U5095 (N_5095,N_3468,N_4255);
and U5096 (N_5096,N_2678,N_4529);
or U5097 (N_5097,N_3418,N_4532);
nand U5098 (N_5098,N_2570,N_4226);
and U5099 (N_5099,N_3708,N_3022);
or U5100 (N_5100,N_3984,N_4299);
or U5101 (N_5101,N_4987,N_4059);
nand U5102 (N_5102,N_3080,N_3715);
and U5103 (N_5103,N_3220,N_3691);
and U5104 (N_5104,N_4415,N_2929);
nand U5105 (N_5105,N_3563,N_4559);
nand U5106 (N_5106,N_3447,N_4801);
nand U5107 (N_5107,N_3285,N_2550);
or U5108 (N_5108,N_2786,N_3098);
and U5109 (N_5109,N_4773,N_2651);
or U5110 (N_5110,N_4721,N_2739);
and U5111 (N_5111,N_3300,N_3752);
or U5112 (N_5112,N_4350,N_3847);
or U5113 (N_5113,N_4248,N_4106);
nor U5114 (N_5114,N_4084,N_2784);
or U5115 (N_5115,N_3350,N_3932);
nand U5116 (N_5116,N_3289,N_3797);
nor U5117 (N_5117,N_3189,N_3237);
nor U5118 (N_5118,N_2639,N_2748);
or U5119 (N_5119,N_3995,N_3200);
or U5120 (N_5120,N_2645,N_4503);
and U5121 (N_5121,N_3853,N_2666);
nand U5122 (N_5122,N_2996,N_2983);
or U5123 (N_5123,N_2975,N_4098);
nand U5124 (N_5124,N_3842,N_4194);
or U5125 (N_5125,N_4844,N_4979);
nand U5126 (N_5126,N_4074,N_4471);
nand U5127 (N_5127,N_4500,N_4469);
and U5128 (N_5128,N_3032,N_3583);
or U5129 (N_5129,N_3223,N_4805);
or U5130 (N_5130,N_2868,N_4719);
and U5131 (N_5131,N_4511,N_3182);
and U5132 (N_5132,N_4341,N_2659);
and U5133 (N_5133,N_3677,N_3666);
nand U5134 (N_5134,N_4577,N_4793);
nand U5135 (N_5135,N_3051,N_3753);
nor U5136 (N_5136,N_2831,N_3239);
nand U5137 (N_5137,N_4740,N_4507);
and U5138 (N_5138,N_2924,N_4641);
and U5139 (N_5139,N_4751,N_4600);
nor U5140 (N_5140,N_3555,N_3460);
or U5141 (N_5141,N_3571,N_3744);
or U5142 (N_5142,N_3942,N_2945);
and U5143 (N_5143,N_3138,N_3111);
nand U5144 (N_5144,N_3746,N_3526);
nand U5145 (N_5145,N_2910,N_4652);
or U5146 (N_5146,N_4056,N_4975);
or U5147 (N_5147,N_4539,N_4749);
or U5148 (N_5148,N_3884,N_2762);
nand U5149 (N_5149,N_3124,N_3660);
or U5150 (N_5150,N_2616,N_3967);
or U5151 (N_5151,N_3633,N_2995);
nor U5152 (N_5152,N_4472,N_4762);
or U5153 (N_5153,N_2521,N_3212);
nor U5154 (N_5154,N_3600,N_4543);
and U5155 (N_5155,N_3537,N_2554);
nor U5156 (N_5156,N_3868,N_3676);
nor U5157 (N_5157,N_2845,N_3662);
and U5158 (N_5158,N_2992,N_3814);
xnor U5159 (N_5159,N_3150,N_3572);
xnor U5160 (N_5160,N_4505,N_3890);
and U5161 (N_5161,N_4456,N_2657);
nand U5162 (N_5162,N_4043,N_4739);
or U5163 (N_5163,N_2860,N_3724);
nand U5164 (N_5164,N_2926,N_3395);
nand U5165 (N_5165,N_4913,N_4572);
or U5166 (N_5166,N_3619,N_3798);
nor U5167 (N_5167,N_3926,N_4391);
nor U5168 (N_5168,N_3562,N_3400);
and U5169 (N_5169,N_4158,N_3568);
or U5170 (N_5170,N_3188,N_4202);
nor U5171 (N_5171,N_3806,N_4782);
and U5172 (N_5172,N_4263,N_4949);
nand U5173 (N_5173,N_2525,N_3825);
and U5174 (N_5174,N_3426,N_2778);
nand U5175 (N_5175,N_3862,N_3025);
or U5176 (N_5176,N_2644,N_4720);
nand U5177 (N_5177,N_4857,N_3037);
and U5178 (N_5178,N_4649,N_3661);
nor U5179 (N_5179,N_3228,N_3316);
and U5180 (N_5180,N_2518,N_4022);
and U5181 (N_5181,N_3839,N_4673);
or U5182 (N_5182,N_4439,N_2968);
or U5183 (N_5183,N_2899,N_3789);
and U5184 (N_5184,N_3119,N_4755);
nand U5185 (N_5185,N_2587,N_2569);
nand U5186 (N_5186,N_4433,N_4519);
or U5187 (N_5187,N_2946,N_3264);
xor U5188 (N_5188,N_4180,N_3428);
and U5189 (N_5189,N_4748,N_3003);
and U5190 (N_5190,N_4483,N_3796);
nand U5191 (N_5191,N_3101,N_3107);
nor U5192 (N_5192,N_3770,N_3192);
nor U5193 (N_5193,N_4728,N_4313);
nor U5194 (N_5194,N_2653,N_2650);
or U5195 (N_5195,N_3626,N_4228);
or U5196 (N_5196,N_2713,N_3126);
nand U5197 (N_5197,N_3303,N_3780);
or U5198 (N_5198,N_4627,N_3540);
and U5199 (N_5199,N_4637,N_4786);
or U5200 (N_5200,N_2911,N_4698);
nand U5201 (N_5201,N_3552,N_4747);
nor U5202 (N_5202,N_4445,N_3427);
nor U5203 (N_5203,N_4294,N_3557);
nor U5204 (N_5204,N_3766,N_3245);
or U5205 (N_5205,N_3486,N_3243);
or U5206 (N_5206,N_3904,N_4693);
nor U5207 (N_5207,N_4512,N_2755);
or U5208 (N_5208,N_4133,N_3355);
or U5209 (N_5209,N_4108,N_2765);
nand U5210 (N_5210,N_3864,N_4615);
nor U5211 (N_5211,N_4276,N_3507);
nand U5212 (N_5212,N_4790,N_2746);
nor U5213 (N_5213,N_3083,N_4959);
or U5214 (N_5214,N_2542,N_2963);
and U5215 (N_5215,N_2984,N_3597);
nor U5216 (N_5216,N_2597,N_3953);
nor U5217 (N_5217,N_4816,N_2527);
and U5218 (N_5218,N_4409,N_4495);
and U5219 (N_5219,N_4964,N_3137);
nor U5220 (N_5220,N_4692,N_4620);
nor U5221 (N_5221,N_3595,N_2617);
and U5222 (N_5222,N_4909,N_4633);
or U5223 (N_5223,N_3727,N_3251);
or U5224 (N_5224,N_4109,N_4396);
or U5225 (N_5225,N_4648,N_4278);
or U5226 (N_5226,N_4437,N_3412);
and U5227 (N_5227,N_3143,N_3672);
or U5228 (N_5228,N_4134,N_3936);
or U5229 (N_5229,N_4866,N_3858);
and U5230 (N_5230,N_2794,N_4184);
or U5231 (N_5231,N_4451,N_3915);
and U5232 (N_5232,N_3762,N_4576);
nand U5233 (N_5233,N_3719,N_3242);
and U5234 (N_5234,N_2512,N_4822);
or U5235 (N_5235,N_2823,N_3115);
or U5236 (N_5236,N_3193,N_2511);
nor U5237 (N_5237,N_3880,N_4737);
nor U5238 (N_5238,N_4677,N_4860);
nor U5239 (N_5239,N_3558,N_4933);
or U5240 (N_5240,N_3332,N_4430);
or U5241 (N_5241,N_3659,N_4667);
or U5242 (N_5242,N_4630,N_2730);
nand U5243 (N_5243,N_3409,N_2668);
or U5244 (N_5244,N_4668,N_4746);
and U5245 (N_5245,N_3882,N_3642);
nor U5246 (N_5246,N_3740,N_3721);
and U5247 (N_5247,N_3869,N_4750);
and U5248 (N_5248,N_3261,N_3755);
and U5249 (N_5249,N_4305,N_4917);
or U5250 (N_5250,N_3846,N_3692);
or U5251 (N_5251,N_3589,N_4890);
nand U5252 (N_5252,N_3844,N_3877);
and U5253 (N_5253,N_3044,N_3382);
nor U5254 (N_5254,N_4556,N_2807);
nand U5255 (N_5255,N_3065,N_3463);
nand U5256 (N_5256,N_4210,N_4402);
nor U5257 (N_5257,N_4832,N_2571);
or U5258 (N_5258,N_4438,N_3905);
and U5259 (N_5259,N_3190,N_4568);
and U5260 (N_5260,N_3928,N_2613);
nor U5261 (N_5261,N_4855,N_4605);
nand U5262 (N_5262,N_2821,N_4757);
nor U5263 (N_5263,N_4928,N_4454);
and U5264 (N_5264,N_3068,N_4763);
nand U5265 (N_5265,N_2565,N_4024);
nand U5266 (N_5266,N_4850,N_3618);
nand U5267 (N_5267,N_2529,N_3828);
nand U5268 (N_5268,N_4968,N_4256);
or U5269 (N_5269,N_2660,N_4839);
nor U5270 (N_5270,N_2629,N_2661);
nor U5271 (N_5271,N_4209,N_2866);
nand U5272 (N_5272,N_3817,N_2835);
or U5273 (N_5273,N_2971,N_3371);
nand U5274 (N_5274,N_4422,N_3988);
and U5275 (N_5275,N_3452,N_3116);
nor U5276 (N_5276,N_4631,N_4477);
or U5277 (N_5277,N_4300,N_4318);
nor U5278 (N_5278,N_2632,N_4023);
nand U5279 (N_5279,N_4443,N_4099);
or U5280 (N_5280,N_3067,N_4522);
or U5281 (N_5281,N_3834,N_2890);
nand U5282 (N_5282,N_4390,N_3118);
nor U5283 (N_5283,N_3346,N_4944);
nor U5284 (N_5284,N_2698,N_4222);
and U5285 (N_5285,N_3874,N_2749);
nor U5286 (N_5286,N_3028,N_4271);
nand U5287 (N_5287,N_3229,N_3149);
nand U5288 (N_5288,N_4939,N_3450);
nor U5289 (N_5289,N_4514,N_4656);
or U5290 (N_5290,N_3650,N_4035);
nand U5291 (N_5291,N_3821,N_2669);
nand U5292 (N_5292,N_3501,N_2849);
and U5293 (N_5293,N_4352,N_2504);
and U5294 (N_5294,N_4843,N_4232);
nor U5295 (N_5295,N_2561,N_2791);
nor U5296 (N_5296,N_4725,N_4590);
or U5297 (N_5297,N_3016,N_3456);
nor U5298 (N_5298,N_4126,N_2772);
nor U5299 (N_5299,N_4973,N_3617);
or U5300 (N_5300,N_4128,N_4870);
and U5301 (N_5301,N_2767,N_4333);
or U5302 (N_5302,N_3972,N_4461);
or U5303 (N_5303,N_2751,N_4690);
nor U5304 (N_5304,N_4475,N_3402);
nand U5305 (N_5305,N_3586,N_3706);
nand U5306 (N_5306,N_3164,N_4761);
or U5307 (N_5307,N_4083,N_3807);
and U5308 (N_5308,N_3716,N_3053);
nor U5309 (N_5309,N_2851,N_3608);
nand U5310 (N_5310,N_3004,N_3924);
or U5311 (N_5311,N_3162,N_3913);
nor U5312 (N_5312,N_2841,N_4029);
nand U5313 (N_5313,N_4103,N_3034);
nor U5314 (N_5314,N_2834,N_4723);
or U5315 (N_5315,N_3231,N_4796);
or U5316 (N_5316,N_4513,N_3060);
nand U5317 (N_5317,N_4775,N_4825);
nand U5318 (N_5318,N_2626,N_3738);
nand U5319 (N_5319,N_3045,N_3286);
nand U5320 (N_5320,N_4718,N_4601);
and U5321 (N_5321,N_4480,N_3442);
nand U5322 (N_5322,N_4787,N_4487);
nor U5323 (N_5323,N_4538,N_3576);
and U5324 (N_5324,N_3343,N_3614);
and U5325 (N_5325,N_4324,N_2846);
and U5326 (N_5326,N_3443,N_3773);
or U5327 (N_5327,N_3041,N_4458);
or U5328 (N_5328,N_2538,N_3091);
nand U5329 (N_5329,N_4440,N_3811);
and U5330 (N_5330,N_4937,N_4320);
nand U5331 (N_5331,N_2878,N_3308);
nor U5332 (N_5332,N_4058,N_2827);
nand U5333 (N_5333,N_4326,N_3786);
nor U5334 (N_5334,N_2572,N_2918);
nand U5335 (N_5335,N_2993,N_3917);
nor U5336 (N_5336,N_3764,N_4366);
nand U5337 (N_5337,N_3968,N_4387);
nor U5338 (N_5338,N_4780,N_3704);
or U5339 (N_5339,N_3870,N_4791);
or U5340 (N_5340,N_3327,N_3449);
and U5341 (N_5341,N_4841,N_3497);
nor U5342 (N_5342,N_4727,N_3553);
nand U5343 (N_5343,N_4260,N_3769);
or U5344 (N_5344,N_2953,N_3405);
nor U5345 (N_5345,N_3374,N_4435);
nand U5346 (N_5346,N_3739,N_2900);
nand U5347 (N_5347,N_2582,N_4879);
nand U5348 (N_5348,N_3639,N_3511);
nor U5349 (N_5349,N_4811,N_3593);
nand U5350 (N_5350,N_3790,N_3029);
and U5351 (N_5351,N_3082,N_4163);
nand U5352 (N_5352,N_3702,N_4632);
nor U5353 (N_5353,N_2893,N_4237);
nor U5354 (N_5354,N_2921,N_3898);
and U5355 (N_5355,N_2633,N_3944);
and U5356 (N_5356,N_3725,N_4923);
nor U5357 (N_5357,N_2663,N_3912);
or U5358 (N_5358,N_3523,N_4696);
nor U5359 (N_5359,N_4063,N_3765);
and U5360 (N_5360,N_2981,N_3417);
or U5361 (N_5361,N_3320,N_4100);
and U5362 (N_5362,N_4457,N_3448);
nor U5363 (N_5363,N_3246,N_3973);
nor U5364 (N_5364,N_4654,N_4441);
nand U5365 (N_5365,N_3161,N_2998);
nand U5366 (N_5366,N_3681,N_3092);
nor U5367 (N_5367,N_3895,N_4882);
and U5368 (N_5368,N_2952,N_3437);
or U5369 (N_5369,N_2876,N_4754);
nor U5370 (N_5370,N_2658,N_2737);
and U5371 (N_5371,N_3483,N_3086);
nor U5372 (N_5372,N_2634,N_4587);
and U5373 (N_5373,N_4077,N_3006);
nand U5374 (N_5374,N_3396,N_4159);
nor U5375 (N_5375,N_3274,N_4466);
and U5376 (N_5376,N_3216,N_3278);
and U5377 (N_5377,N_4701,N_3411);
and U5378 (N_5378,N_3854,N_3310);
and U5379 (N_5379,N_4087,N_3133);
and U5380 (N_5380,N_3550,N_4898);
and U5381 (N_5381,N_3840,N_4927);
nand U5382 (N_5382,N_2578,N_4160);
and U5383 (N_5383,N_3761,N_3352);
nor U5384 (N_5384,N_3800,N_3827);
nor U5385 (N_5385,N_2567,N_2552);
or U5386 (N_5386,N_2764,N_3588);
nor U5387 (N_5387,N_2969,N_4779);
or U5388 (N_5388,N_3634,N_4508);
and U5389 (N_5389,N_4661,N_3033);
and U5390 (N_5390,N_4560,N_3156);
and U5391 (N_5391,N_3199,N_4638);
or U5392 (N_5392,N_4829,N_2721);
and U5393 (N_5393,N_4685,N_3206);
and U5394 (N_5394,N_4174,N_4069);
nor U5395 (N_5395,N_3577,N_2549);
or U5396 (N_5396,N_2826,N_3128);
nor U5397 (N_5397,N_3883,N_2560);
nor U5398 (N_5398,N_3643,N_3857);
and U5399 (N_5399,N_4875,N_3528);
or U5400 (N_5400,N_3808,N_4216);
nor U5401 (N_5401,N_3646,N_2568);
nor U5402 (N_5402,N_4684,N_3863);
or U5403 (N_5403,N_4858,N_3131);
or U5404 (N_5404,N_4465,N_4131);
nor U5405 (N_5405,N_3324,N_4355);
or U5406 (N_5406,N_3039,N_3982);
nor U5407 (N_5407,N_4296,N_4066);
nand U5408 (N_5408,N_2801,N_3071);
nor U5409 (N_5409,N_3094,N_3587);
nor U5410 (N_5410,N_3865,N_3978);
and U5411 (N_5411,N_2832,N_3309);
or U5412 (N_5412,N_2690,N_3360);
nor U5413 (N_5413,N_3485,N_3611);
and U5414 (N_5414,N_2734,N_4837);
nor U5415 (N_5415,N_4137,N_4419);
and U5416 (N_5416,N_4966,N_3479);
nor U5417 (N_5417,N_3969,N_3233);
or U5418 (N_5418,N_3641,N_3852);
nand U5419 (N_5419,N_2591,N_3415);
nand U5420 (N_5420,N_3194,N_4025);
or U5421 (N_5421,N_3891,N_4659);
xnor U5422 (N_5422,N_3224,N_3997);
nand U5423 (N_5423,N_4566,N_4189);
or U5424 (N_5424,N_3667,N_2558);
and U5425 (N_5425,N_2649,N_3722);
and U5426 (N_5426,N_4819,N_2592);
and U5427 (N_5427,N_4286,N_4778);
nand U5428 (N_5428,N_2501,N_4165);
nor U5429 (N_5429,N_4081,N_4030);
and U5430 (N_5430,N_2564,N_4935);
nand U5431 (N_5431,N_2908,N_3373);
and U5432 (N_5432,N_4195,N_2872);
nand U5433 (N_5433,N_3566,N_3657);
nor U5434 (N_5434,N_3023,N_2540);
nand U5435 (N_5435,N_4812,N_4117);
or U5436 (N_5436,N_3527,N_4428);
nor U5437 (N_5437,N_3737,N_3621);
and U5438 (N_5438,N_4288,N_4523);
or U5439 (N_5439,N_3348,N_3685);
nor U5440 (N_5440,N_4462,N_4104);
and U5441 (N_5441,N_4373,N_2769);
and U5442 (N_5442,N_2867,N_3787);
nand U5443 (N_5443,N_3873,N_4982);
nor U5444 (N_5444,N_2799,N_2881);
or U5445 (N_5445,N_4509,N_3850);
nor U5446 (N_5446,N_3901,N_3775);
nor U5447 (N_5447,N_3027,N_3191);
and U5448 (N_5448,N_3885,N_3598);
nor U5449 (N_5449,N_3845,N_4217);
and U5450 (N_5450,N_2886,N_4264);
and U5451 (N_5451,N_4783,N_4312);
nor U5452 (N_5452,N_3425,N_2604);
and U5453 (N_5453,N_2684,N_4006);
or U5454 (N_5454,N_3380,N_3108);
or U5455 (N_5455,N_4499,N_4894);
xor U5456 (N_5456,N_3057,N_3999);
and U5457 (N_5457,N_2500,N_2630);
or U5458 (N_5458,N_3836,N_4251);
and U5459 (N_5459,N_2759,N_4642);
nor U5460 (N_5460,N_3632,N_4119);
nor U5461 (N_5461,N_2514,N_2870);
or U5462 (N_5462,N_3419,N_4096);
nand U5463 (N_5463,N_4170,N_3441);
and U5464 (N_5464,N_4399,N_2588);
or U5465 (N_5465,N_3596,N_2729);
or U5466 (N_5466,N_3774,N_2806);
and U5467 (N_5467,N_2985,N_3078);
nand U5468 (N_5468,N_3794,N_4851);
or U5469 (N_5469,N_3688,N_3088);
nor U5470 (N_5470,N_4213,N_3085);
or U5471 (N_5471,N_3805,N_4002);
nor U5472 (N_5472,N_4921,N_4382);
nor U5473 (N_5473,N_3613,N_3957);
nor U5474 (N_5474,N_3482,N_3777);
nand U5475 (N_5475,N_4233,N_2701);
and U5476 (N_5476,N_4992,N_3818);
or U5477 (N_5477,N_3072,N_2903);
nor U5478 (N_5478,N_4279,N_3366);
nor U5479 (N_5479,N_4891,N_4658);
or U5480 (N_5480,N_4931,N_2859);
and U5481 (N_5481,N_2915,N_4845);
and U5482 (N_5482,N_4497,N_2607);
nand U5483 (N_5483,N_4622,N_2523);
nand U5484 (N_5484,N_3179,N_4246);
and U5485 (N_5485,N_3575,N_3640);
or U5486 (N_5486,N_4621,N_2744);
and U5487 (N_5487,N_3434,N_3491);
and U5488 (N_5488,N_2580,N_4799);
nor U5489 (N_5489,N_4088,N_2688);
nor U5490 (N_5490,N_4345,N_2958);
nor U5491 (N_5491,N_4930,N_4289);
or U5492 (N_5492,N_4595,N_2672);
and U5493 (N_5493,N_3021,N_4038);
or U5494 (N_5494,N_4986,N_3011);
and U5495 (N_5495,N_4182,N_2989);
or U5496 (N_5496,N_4484,N_4578);
nand U5497 (N_5497,N_2635,N_2809);
and U5498 (N_5498,N_3471,N_4191);
nand U5499 (N_5499,N_3684,N_4635);
nor U5500 (N_5500,N_4212,N_3931);
and U5501 (N_5501,N_3388,N_3887);
nor U5502 (N_5502,N_4795,N_4537);
and U5503 (N_5503,N_3622,N_2738);
or U5504 (N_5504,N_3291,N_4647);
or U5505 (N_5505,N_2931,N_3142);
nand U5506 (N_5506,N_3748,N_4421);
nor U5507 (N_5507,N_3455,N_3315);
or U5508 (N_5508,N_4478,N_4047);
and U5509 (N_5509,N_4257,N_2716);
or U5510 (N_5510,N_2820,N_2771);
or U5511 (N_5511,N_4245,N_4176);
nor U5512 (N_5512,N_3908,N_2677);
and U5513 (N_5513,N_4050,N_4157);
and U5514 (N_5514,N_3718,N_3710);
nand U5515 (N_5515,N_3998,N_3097);
and U5516 (N_5516,N_2731,N_2780);
and U5517 (N_5517,N_4708,N_4413);
and U5518 (N_5518,N_4124,N_2742);
and U5519 (N_5519,N_4385,N_3454);
nand U5520 (N_5520,N_4068,N_3837);
nand U5521 (N_5521,N_4567,N_2787);
nor U5522 (N_5522,N_4678,N_2961);
and U5523 (N_5523,N_3155,N_4776);
nor U5524 (N_5524,N_3276,N_3084);
and U5525 (N_5525,N_4846,N_3720);
and U5526 (N_5526,N_2986,N_4376);
nand U5527 (N_5527,N_2595,N_4910);
xor U5528 (N_5528,N_2954,N_2962);
or U5529 (N_5529,N_2934,N_3897);
or U5530 (N_5530,N_4151,N_3782);
nand U5531 (N_5531,N_3983,N_4551);
and U5532 (N_5532,N_3756,N_2863);
nand U5533 (N_5533,N_3270,N_4869);
or U5534 (N_5534,N_2988,N_4650);
and U5535 (N_5535,N_3430,N_4442);
and U5536 (N_5536,N_3819,N_2816);
nor U5537 (N_5537,N_4166,N_2732);
and U5538 (N_5538,N_2676,N_3255);
or U5539 (N_5539,N_3283,N_4336);
or U5540 (N_5540,N_3446,N_4342);
nor U5541 (N_5541,N_4584,N_3317);
xnor U5542 (N_5542,N_4717,N_4092);
or U5543 (N_5543,N_3364,N_2930);
nor U5544 (N_5544,N_3401,N_3337);
nand U5545 (N_5545,N_4219,N_2743);
and U5546 (N_5546,N_4893,N_3548);
nand U5547 (N_5547,N_4932,N_3990);
and U5548 (N_5548,N_3195,N_4889);
nor U5549 (N_5549,N_3263,N_2622);
or U5550 (N_5550,N_4814,N_4093);
or U5551 (N_5551,N_4453,N_3145);
xnor U5552 (N_5552,N_3993,N_4167);
nor U5553 (N_5553,N_2695,N_2696);
and U5554 (N_5554,N_3509,N_4624);
nor U5555 (N_5555,N_3605,N_2510);
nor U5556 (N_5556,N_4557,N_3493);
nand U5557 (N_5557,N_3620,N_2987);
or U5558 (N_5558,N_2798,N_3735);
or U5559 (N_5559,N_2818,N_3759);
nand U5560 (N_5560,N_2937,N_3288);
nand U5561 (N_5561,N_4227,N_3413);
and U5562 (N_5562,N_2611,N_2741);
nor U5563 (N_5563,N_3075,N_4302);
nand U5564 (N_5564,N_3181,N_4491);
nor U5565 (N_5565,N_3651,N_4169);
or U5566 (N_5566,N_3876,N_3647);
or U5567 (N_5567,N_4020,N_4459);
nand U5568 (N_5568,N_2556,N_3307);
and U5569 (N_5569,N_3795,N_4836);
nand U5570 (N_5570,N_4772,N_3604);
nand U5571 (N_5571,N_4317,N_3219);
nand U5572 (N_5572,N_3481,N_2577);
or U5573 (N_5573,N_2543,N_3368);
and U5574 (N_5574,N_3475,N_3656);
nor U5575 (N_5575,N_3260,N_4540);
and U5576 (N_5576,N_4899,N_2943);
xnor U5577 (N_5577,N_3267,N_4877);
nand U5578 (N_5578,N_3713,N_2722);
nand U5579 (N_5579,N_4574,N_3630);
nor U5580 (N_5580,N_4344,N_4962);
and U5581 (N_5581,N_4702,N_3989);
or U5582 (N_5582,N_3564,N_4639);
nor U5583 (N_5583,N_2916,N_4671);
and U5584 (N_5584,N_3824,N_3329);
nor U5585 (N_5585,N_3344,N_4848);
and U5586 (N_5586,N_3535,N_4925);
or U5587 (N_5587,N_4110,N_4669);
or U5588 (N_5588,N_2704,N_2977);
nor U5589 (N_5589,N_4603,N_2957);
and U5590 (N_5590,N_3211,N_2824);
nand U5591 (N_5591,N_3494,N_4406);
or U5592 (N_5592,N_3105,N_4021);
nand U5593 (N_5593,N_3937,N_3198);
or U5594 (N_5594,N_4838,N_4646);
nand U5595 (N_5595,N_3159,N_4918);
or U5596 (N_5596,N_4295,N_3240);
and U5597 (N_5597,N_4710,N_4183);
nor U5598 (N_5598,N_3545,N_4242);
nand U5599 (N_5599,N_3186,N_3768);
nand U5600 (N_5600,N_3763,N_4764);
and U5601 (N_5601,N_4410,N_2904);
nor U5602 (N_5602,N_2927,N_2819);
or U5603 (N_5603,N_4900,N_3066);
and U5604 (N_5604,N_4051,N_3648);
nand U5605 (N_5605,N_2608,N_3335);
nand U5606 (N_5606,N_2973,N_2935);
and U5607 (N_5607,N_3342,N_3757);
nand U5608 (N_5608,N_4951,N_4645);
and U5609 (N_5609,N_4061,N_4014);
or U5610 (N_5610,N_4831,N_4916);
and U5611 (N_5611,N_4823,N_4905);
nor U5612 (N_5612,N_4274,N_4552);
and U5613 (N_5613,N_4125,N_3214);
nand U5614 (N_5614,N_3743,N_4282);
or U5615 (N_5615,N_2773,N_3038);
and U5616 (N_5616,N_4388,N_3496);
nand U5617 (N_5617,N_3287,N_3040);
nor U5618 (N_5618,N_3421,N_4606);
nor U5619 (N_5619,N_4231,N_3394);
nand U5620 (N_5620,N_4052,N_2682);
or U5621 (N_5621,N_4745,N_3525);
and U5622 (N_5622,N_4113,N_4589);
and U5623 (N_5623,N_3152,N_3569);
and U5624 (N_5624,N_3238,N_2624);
and U5625 (N_5625,N_3831,N_4947);
nor U5626 (N_5626,N_4007,N_3247);
nor U5627 (N_5627,N_4741,N_3582);
nor U5628 (N_5628,N_3649,N_3964);
nand U5629 (N_5629,N_3484,N_4482);
nor U5630 (N_5630,N_4405,N_4963);
and U5631 (N_5631,N_2586,N_3971);
nor U5632 (N_5632,N_3026,N_3772);
and U5633 (N_5633,N_4447,N_3623);
and U5634 (N_5634,N_3398,N_4293);
and U5635 (N_5635,N_3703,N_4418);
nand U5636 (N_5636,N_4901,N_4140);
and U5637 (N_5637,N_3390,N_4040);
nor U5638 (N_5638,N_4374,N_4700);
nor U5639 (N_5639,N_3930,N_4817);
or U5640 (N_5640,N_3440,N_2956);
and U5641 (N_5641,N_4634,N_4236);
nand U5642 (N_5642,N_4476,N_2848);
or U5643 (N_5643,N_4150,N_3510);
nor U5644 (N_5644,N_3268,N_3168);
nand U5645 (N_5645,N_3218,N_3690);
or U5646 (N_5646,N_2974,N_3519);
and U5647 (N_5647,N_4348,N_2847);
or U5648 (N_5648,N_4926,N_3734);
nor U5649 (N_5649,N_2871,N_3054);
and U5650 (N_5650,N_4853,N_2966);
or U5651 (N_5651,N_3686,N_3860);
nand U5652 (N_5652,N_4013,N_2603);
and U5653 (N_5653,N_3363,N_3833);
or U5654 (N_5654,N_3391,N_2610);
nor U5655 (N_5655,N_4377,N_3745);
or U5656 (N_5656,N_4806,N_4821);
and U5657 (N_5657,N_2840,N_4353);
nand U5658 (N_5658,N_3472,N_4155);
nor U5659 (N_5659,N_3565,N_3573);
nor U5660 (N_5660,N_2895,N_3804);
nor U5661 (N_5661,N_4127,N_4380);
nor U5662 (N_5662,N_2686,N_4655);
xor U5663 (N_5663,N_4849,N_4874);
nand U5664 (N_5664,N_2906,N_2852);
xnor U5665 (N_5665,N_3784,N_4343);
nor U5666 (N_5666,N_3802,N_4207);
or U5667 (N_5667,N_3512,N_4046);
or U5668 (N_5668,N_3813,N_2726);
or U5669 (N_5669,N_2950,N_2796);
nor U5670 (N_5670,N_4897,N_4824);
nor U5671 (N_5671,N_3653,N_4582);
nor U5672 (N_5672,N_3861,N_4712);
nor U5673 (N_5673,N_4204,N_2955);
and U5674 (N_5674,N_3353,N_3146);
nor U5675 (N_5675,N_4460,N_2596);
and U5676 (N_5676,N_2530,N_3163);
nor U5677 (N_5677,N_4506,N_4859);
or U5678 (N_5678,N_2535,N_3615);
nor U5679 (N_5679,N_3697,N_2509);
xnor U5680 (N_5680,N_2531,N_4676);
or U5681 (N_5681,N_4965,N_4016);
nor U5682 (N_5682,N_3570,N_4896);
nor U5683 (N_5683,N_3878,N_4998);
nor U5684 (N_5684,N_3592,N_3478);
nor U5685 (N_5685,N_3424,N_3423);
nand U5686 (N_5686,N_4852,N_4280);
or U5687 (N_5687,N_4175,N_4034);
nor U5688 (N_5688,N_3609,N_2892);
nand U5689 (N_5689,N_3282,N_3297);
nand U5690 (N_5690,N_4919,N_2513);
or U5691 (N_5691,N_4417,N_3345);
or U5692 (N_5692,N_4501,N_2803);
nand U5693 (N_5693,N_2763,N_4868);
and U5694 (N_5694,N_3591,N_4062);
nand U5695 (N_5695,N_4147,N_4455);
nand U5696 (N_5696,N_3099,N_4980);
nand U5697 (N_5697,N_4680,N_4329);
or U5698 (N_5698,N_4895,N_3823);
and U5699 (N_5699,N_3379,N_4978);
or U5700 (N_5700,N_2896,N_3323);
nand U5701 (N_5701,N_3712,N_3336);
or U5702 (N_5702,N_3778,N_3546);
nor U5703 (N_5703,N_4771,N_3976);
nor U5704 (N_5704,N_4781,N_3520);
nand U5705 (N_5705,N_4834,N_3444);
or U5706 (N_5706,N_4815,N_2898);
or U5707 (N_5707,N_4942,N_3301);
nor U5708 (N_5708,N_4694,N_2563);
and U5709 (N_5709,N_4604,N_2654);
or U5710 (N_5710,N_3328,N_3435);
or U5711 (N_5711,N_3541,N_4904);
nand U5712 (N_5712,N_3422,N_2566);
nand U5713 (N_5713,N_3872,N_2623);
nand U5714 (N_5714,N_2728,N_4797);
nor U5715 (N_5715,N_2621,N_3173);
or U5716 (N_5716,N_3941,N_2967);
and U5717 (N_5717,N_4520,N_4623);
nor U5718 (N_5718,N_3464,N_3522);
nor U5719 (N_5719,N_4026,N_3732);
and U5720 (N_5720,N_2800,N_4908);
nand U5721 (N_5721,N_4414,N_4999);
or U5722 (N_5722,N_4713,N_2750);
or U5723 (N_5723,N_3996,N_4463);
nor U5724 (N_5724,N_2637,N_3416);
nor U5725 (N_5725,N_4072,N_4977);
nand U5726 (N_5726,N_2585,N_3241);
nor U5727 (N_5727,N_3911,N_4726);
or U5728 (N_5728,N_4179,N_3121);
xor U5729 (N_5729,N_4008,N_3326);
and U5730 (N_5730,N_3158,N_4609);
or U5731 (N_5731,N_4297,N_4149);
and U5732 (N_5732,N_3959,N_4434);
or U5733 (N_5733,N_4883,N_3729);
and U5734 (N_5734,N_3962,N_2711);
or U5735 (N_5735,N_4564,N_3952);
nand U5736 (N_5736,N_4071,N_3594);
nor U5737 (N_5737,N_4473,N_4752);
or U5738 (N_5738,N_4912,N_4527);
nand U5739 (N_5739,N_2844,N_3820);
nand U5740 (N_5740,N_2753,N_4162);
and U5741 (N_5741,N_3760,N_4314);
or U5742 (N_5742,N_2805,N_4524);
or U5743 (N_5743,N_4662,N_4357);
or U5744 (N_5744,N_3832,N_2865);
nand U5745 (N_5745,N_2508,N_4479);
nor U5746 (N_5746,N_2862,N_3073);
nand U5747 (N_5747,N_4444,N_3631);
and U5748 (N_5748,N_4012,N_3175);
or U5749 (N_5749,N_3292,N_3381);
and U5750 (N_5750,N_2717,N_4810);
nor U5751 (N_5751,N_3920,N_4292);
and U5752 (N_5752,N_4792,N_4349);
nor U5753 (N_5753,N_4015,N_2933);
nor U5754 (N_5754,N_2664,N_4515);
nand U5755 (N_5755,N_3549,N_3147);
or U5756 (N_5756,N_2813,N_2600);
or U5757 (N_5757,N_4830,N_4618);
or U5758 (N_5758,N_4252,N_2817);
and U5759 (N_5759,N_4316,N_2757);
or U5760 (N_5760,N_4247,N_2694);
nand U5761 (N_5761,N_3383,N_2740);
or U5762 (N_5762,N_4005,N_3906);
and U5763 (N_5763,N_3302,N_3130);
and U5764 (N_5764,N_4945,N_3689);
nand U5765 (N_5765,N_4758,N_4736);
and U5766 (N_5766,N_4259,N_4861);
nand U5767 (N_5767,N_2825,N_3986);
nand U5768 (N_5768,N_4181,N_4381);
or U5769 (N_5769,N_4818,N_3517);
nand U5770 (N_5770,N_4198,N_4186);
nor U5771 (N_5771,N_3458,N_4617);
nor U5772 (N_5772,N_3696,N_4188);
or U5773 (N_5773,N_4827,N_2708);
or U5774 (N_5774,N_3172,N_3665);
or U5775 (N_5775,N_4665,N_4340);
nor U5776 (N_5776,N_3892,N_3357);
nand U5777 (N_5777,N_4053,N_2541);
nor U5778 (N_5778,N_3473,N_3132);
nand U5779 (N_5779,N_4664,N_4599);
nand U5780 (N_5780,N_4924,N_2842);
and U5781 (N_5781,N_4610,N_3480);
nand U5782 (N_5782,N_3505,N_4886);
or U5783 (N_5783,N_4803,N_4842);
nand U5784 (N_5784,N_3749,N_3112);
and U5785 (N_5785,N_3171,N_3180);
or U5786 (N_5786,N_2897,N_3244);
or U5787 (N_5787,N_3728,N_3645);
nor U5788 (N_5788,N_4865,N_4971);
or U5789 (N_5789,N_4107,N_3500);
nor U5790 (N_5790,N_4200,N_4303);
and U5791 (N_5791,N_4802,N_3043);
nand U5792 (N_5792,N_4588,N_3354);
nand U5793 (N_5793,N_2812,N_4095);
and U5794 (N_5794,N_2628,N_2912);
nor U5795 (N_5795,N_2636,N_3369);
nor U5796 (N_5796,N_3377,N_4361);
nor U5797 (N_5797,N_4766,N_4273);
or U5798 (N_5798,N_3176,N_3530);
and U5799 (N_5799,N_3970,N_3980);
nor U5800 (N_5800,N_2656,N_4208);
nor U5801 (N_5801,N_3140,N_4398);
or U5802 (N_5802,N_2864,N_4153);
and U5803 (N_5803,N_4571,N_2795);
nand U5804 (N_5804,N_3894,N_3459);
and U5805 (N_5805,N_3638,N_4378);
or U5806 (N_5806,N_3579,N_3627);
nor U5807 (N_5807,N_3585,N_3318);
and U5808 (N_5808,N_4657,N_4663);
nor U5809 (N_5809,N_2793,N_2625);
nand U5810 (N_5810,N_4492,N_3498);
nor U5811 (N_5811,N_2942,N_3018);
nand U5812 (N_5812,N_4581,N_2640);
or U5813 (N_5813,N_3215,N_3758);
nand U5814 (N_5814,N_4744,N_3187);
nor U5815 (N_5815,N_4593,N_3855);
and U5816 (N_5816,N_4330,N_3465);
nor U5817 (N_5817,N_4395,N_2553);
and U5818 (N_5818,N_3298,N_4311);
nand U5819 (N_5819,N_4031,N_4545);
nor U5820 (N_5820,N_4903,N_2519);
and U5821 (N_5821,N_3536,N_2579);
or U5822 (N_5822,N_4086,N_2804);
and U5823 (N_5823,N_4432,N_4301);
nand U5824 (N_5824,N_3462,N_3612);
or U5825 (N_5825,N_3445,N_4094);
and U5826 (N_5826,N_3521,N_2783);
or U5827 (N_5827,N_3736,N_2854);
nand U5828 (N_5828,N_2972,N_3196);
and U5829 (N_5829,N_3886,N_2776);
nand U5830 (N_5830,N_3694,N_4716);
nor U5831 (N_5831,N_3678,N_3747);
nor U5832 (N_5832,N_3279,N_2941);
or U5833 (N_5833,N_4490,N_4784);
nor U5834 (N_5834,N_3939,N_2919);
nand U5835 (N_5835,N_4995,N_3321);
nor U5836 (N_5836,N_3280,N_2754);
or U5837 (N_5837,N_3208,N_4238);
nor U5838 (N_5838,N_3803,N_4528);
and U5839 (N_5839,N_3889,N_3076);
or U5840 (N_5840,N_4244,N_3466);
and U5841 (N_5841,N_3269,N_4510);
nor U5842 (N_5842,N_3556,N_3628);
and U5843 (N_5843,N_4468,N_3157);
or U5844 (N_5844,N_4619,N_3387);
and U5845 (N_5845,N_3063,N_2615);
nor U5846 (N_5846,N_2646,N_3049);
nand U5847 (N_5847,N_4936,N_4881);
and U5848 (N_5848,N_4863,N_3495);
xnor U5849 (N_5849,N_3429,N_4517);
nand U5850 (N_5850,N_4105,N_3012);
nor U5851 (N_5851,N_3095,N_2516);
and U5852 (N_5852,N_4310,N_2522);
nand U5853 (N_5853,N_3313,N_2843);
nand U5854 (N_5854,N_4102,N_4794);
and U5855 (N_5855,N_3751,N_4789);
or U5856 (N_5856,N_2788,N_3822);
nand U5857 (N_5857,N_2885,N_3122);
and U5858 (N_5858,N_2534,N_4544);
nor U5859 (N_5859,N_3331,N_4612);
or U5860 (N_5860,N_3927,N_2555);
nor U5861 (N_5861,N_4173,N_4682);
nor U5862 (N_5862,N_3120,N_4885);
nand U5863 (N_5863,N_4009,N_3046);
or U5864 (N_5864,N_2761,N_2714);
nand U5865 (N_5865,N_2736,N_3948);
nand U5866 (N_5866,N_4626,N_4057);
and U5867 (N_5867,N_4835,N_4145);
xnor U5868 (N_5868,N_2830,N_3397);
nand U5869 (N_5869,N_2675,N_4446);
and U5870 (N_5870,N_3404,N_3674);
nor U5871 (N_5871,N_3334,N_3074);
xnor U5872 (N_5872,N_3896,N_4876);
or U5873 (N_5873,N_3700,N_3918);
and U5874 (N_5874,N_4969,N_4674);
nand U5875 (N_5875,N_4970,N_4820);
or U5876 (N_5876,N_3177,N_4404);
and U5877 (N_5877,N_4032,N_3699);
nor U5878 (N_5878,N_2999,N_4190);
nand U5879 (N_5879,N_4400,N_3203);
nor U5880 (N_5880,N_4218,N_4290);
and U5881 (N_5881,N_4079,N_3372);
nand U5882 (N_5882,N_4547,N_3514);
nand U5883 (N_5883,N_2515,N_4055);
nor U5884 (N_5884,N_3089,N_4770);
or U5885 (N_5885,N_3603,N_2785);
nand U5886 (N_5886,N_4044,N_4367);
nand U5887 (N_5887,N_4943,N_3338);
nand U5888 (N_5888,N_3529,N_3534);
nand U5889 (N_5889,N_3561,N_3312);
or U5890 (N_5890,N_4489,N_2861);
and U5891 (N_5891,N_4493,N_4033);
nand U5892 (N_5892,N_3974,N_4347);
or U5893 (N_5893,N_4731,N_4116);
or U5894 (N_5894,N_2719,N_3090);
and U5895 (N_5895,N_2928,N_3826);
or U5896 (N_5896,N_4225,N_3625);
or U5897 (N_5897,N_2612,N_3030);
and U5898 (N_5898,N_4185,N_4408);
and U5899 (N_5899,N_3069,N_3955);
or U5900 (N_5900,N_4756,N_2601);
or U5901 (N_5901,N_4000,N_4873);
nor U5902 (N_5902,N_4706,N_3213);
or U5903 (N_5903,N_3714,N_3399);
nand U5904 (N_5904,N_3477,N_2725);
or U5905 (N_5905,N_3325,N_4467);
nor U5906 (N_5906,N_2774,N_2727);
and U5907 (N_5907,N_4130,N_4743);
nor U5908 (N_5908,N_3077,N_4003);
nor U5909 (N_5909,N_3954,N_3178);
nor U5910 (N_5910,N_2691,N_4065);
or U5911 (N_5911,N_4423,N_4262);
nor U5912 (N_5912,N_2917,N_4553);
nor U5913 (N_5913,N_2693,N_4555);
nand U5914 (N_5914,N_3717,N_2589);
nor U5915 (N_5915,N_2539,N_4192);
or U5916 (N_5916,N_3902,N_2828);
nand U5917 (N_5917,N_2606,N_4048);
or U5918 (N_5918,N_4878,N_4268);
or U5919 (N_5919,N_3436,N_2914);
nand U5920 (N_5920,N_2939,N_2758);
nor U5921 (N_5921,N_3461,N_2811);
and U5922 (N_5922,N_3453,N_2583);
or U5923 (N_5923,N_3184,N_3249);
or U5924 (N_5924,N_4867,N_2777);
nor U5925 (N_5925,N_4981,N_3058);
or U5926 (N_5926,N_3848,N_2562);
nor U5927 (N_5927,N_3518,N_3002);
nor U5928 (N_5928,N_4375,N_3559);
and U5929 (N_5929,N_2925,N_2960);
and U5930 (N_5930,N_3370,N_4309);
nor U5931 (N_5931,N_4148,N_4732);
and U5932 (N_5932,N_3492,N_2545);
and U5933 (N_5933,N_4602,N_2994);
or U5934 (N_5934,N_2940,N_3385);
nand U5935 (N_5935,N_4272,N_4813);
nor U5936 (N_5936,N_4298,N_4379);
nand U5937 (N_5937,N_2544,N_3602);
or U5938 (N_5938,N_2670,N_2970);
nand U5939 (N_5939,N_3601,N_2766);
nand U5940 (N_5940,N_2602,N_3209);
nor U5941 (N_5941,N_4327,N_2642);
or U5942 (N_5942,N_3938,N_3516);
nand U5943 (N_5943,N_2503,N_3024);
or U5944 (N_5944,N_3403,N_4809);
nor U5945 (N_5945,N_3290,N_3830);
and U5946 (N_5946,N_4112,N_4436);
and U5947 (N_5947,N_3683,N_4628);
nand U5948 (N_5948,N_3277,N_2718);
or U5949 (N_5949,N_4132,N_3109);
and U5950 (N_5950,N_4864,N_4136);
and U5951 (N_5951,N_3139,N_4416);
or U5952 (N_5952,N_2822,N_3754);
or U5953 (N_5953,N_2782,N_4580);
nor U5954 (N_5954,N_2980,N_3504);
nor U5955 (N_5955,N_2802,N_2598);
and U5956 (N_5956,N_3234,N_3532);
nor U5957 (N_5957,N_4644,N_3991);
or U5958 (N_5958,N_3015,N_3008);
nand U5959 (N_5959,N_3386,N_3711);
or U5960 (N_5960,N_4575,N_4234);
nand U5961 (N_5961,N_3392,N_4425);
or U5962 (N_5962,N_3907,N_3170);
and U5963 (N_5963,N_2683,N_2652);
nor U5964 (N_5964,N_4997,N_2702);
nor U5965 (N_5965,N_4541,N_2665);
and U5966 (N_5966,N_4954,N_2747);
and U5967 (N_5967,N_4168,N_4123);
and U5968 (N_5968,N_3508,N_3547);
nand U5969 (N_5969,N_4073,N_2699);
nand U5970 (N_5970,N_2976,N_3799);
and U5971 (N_5971,N_4429,N_4205);
or U5972 (N_5972,N_2936,N_3859);
or U5973 (N_5973,N_3951,N_3070);
or U5974 (N_5974,N_3333,N_4666);
or U5975 (N_5975,N_3169,N_2647);
nor U5976 (N_5976,N_4346,N_3680);
or U5977 (N_5977,N_3202,N_3106);
nand U5978 (N_5978,N_4950,N_3490);
nand U5979 (N_5979,N_3001,N_3909);
or U5980 (N_5980,N_2810,N_4765);
nor U5981 (N_5981,N_3629,N_3266);
and U5982 (N_5982,N_4498,N_3469);
nand U5983 (N_5983,N_4798,N_2680);
nor U5984 (N_5984,N_3687,N_2551);
or U5985 (N_5985,N_3750,N_3431);
or U5986 (N_5986,N_2888,N_3940);
or U5987 (N_5987,N_3197,N_2839);
nor U5988 (N_5988,N_3956,N_4496);
xor U5989 (N_5989,N_2605,N_4392);
or U5990 (N_5990,N_4424,N_3856);
nand U5991 (N_5991,N_2692,N_4990);
or U5992 (N_5992,N_3637,N_3538);
nor U5993 (N_5993,N_4941,N_2880);
nand U5994 (N_5994,N_3433,N_4579);
nand U5995 (N_5995,N_4573,N_2833);
and U5996 (N_5996,N_4241,N_4196);
or U5997 (N_5997,N_4957,N_3007);
nand U5998 (N_5998,N_3606,N_2760);
nand U5999 (N_5999,N_2891,N_4554);
nor U6000 (N_6000,N_4607,N_4070);
or U6001 (N_6001,N_4193,N_3809);
nand U6002 (N_6002,N_3079,N_3299);
or U6003 (N_6003,N_2991,N_4359);
or U6004 (N_6004,N_4938,N_3319);
nand U6005 (N_6005,N_4705,N_4558);
and U6006 (N_6006,N_4152,N_3947);
nor U6007 (N_6007,N_2706,N_3165);
nand U6008 (N_6008,N_4470,N_3994);
and U6009 (N_6009,N_4993,N_3934);
or U6010 (N_6010,N_2528,N_2978);
nor U6011 (N_6011,N_3635,N_3100);
and U6012 (N_6012,N_4526,N_2889);
or U6013 (N_6013,N_2641,N_4672);
nand U6014 (N_6014,N_4884,N_4201);
and U6015 (N_6015,N_4018,N_4742);
and U6016 (N_6016,N_3879,N_3658);
and U6017 (N_6017,N_4369,N_3975);
nand U6018 (N_6018,N_2685,N_4304);
nand U6019 (N_6019,N_4156,N_4397);
nor U6020 (N_6020,N_3531,N_3544);
nor U6021 (N_6021,N_3793,N_4709);
and U6022 (N_6022,N_4420,N_4010);
nor U6023 (N_6023,N_4291,N_4407);
and U6024 (N_6024,N_2537,N_4888);
and U6025 (N_6025,N_3254,N_3293);
and U6026 (N_6026,N_4920,N_3376);
or U6027 (N_6027,N_4178,N_2703);
or U6028 (N_6028,N_4714,N_3036);
nand U6029 (N_6029,N_2965,N_4856);
or U6030 (N_6030,N_4598,N_3061);
or U6031 (N_6031,N_4902,N_3723);
and U6032 (N_6032,N_2920,N_2932);
and U6033 (N_6033,N_4561,N_3235);
nand U6034 (N_6034,N_4037,N_3042);
and U6035 (N_6035,N_3987,N_3816);
or U6036 (N_6036,N_4101,N_4833);
and U6037 (N_6037,N_3093,N_2594);
nand U6038 (N_6038,N_3893,N_4946);
or U6039 (N_6039,N_4085,N_3843);
nor U6040 (N_6040,N_2533,N_3414);
or U6041 (N_6041,N_4660,N_2836);
xnor U6042 (N_6042,N_4067,N_3248);
or U6043 (N_6043,N_2735,N_4411);
or U6044 (N_6044,N_4591,N_4504);
nand U6045 (N_6045,N_4691,N_4144);
or U6046 (N_6046,N_3624,N_4534);
nor U6047 (N_6047,N_3673,N_3776);
and U6048 (N_6048,N_4586,N_3393);
or U6049 (N_6049,N_3183,N_3502);
nand U6050 (N_6050,N_4284,N_4753);
nand U6051 (N_6051,N_3707,N_3127);
or U6052 (N_6052,N_4697,N_2869);
or U6053 (N_6053,N_3670,N_2707);
nor U6054 (N_6054,N_3330,N_4914);
nor U6055 (N_6055,N_3258,N_4351);
nor U6056 (N_6056,N_4114,N_3921);
and U6057 (N_6057,N_2581,N_3087);
nand U6058 (N_6058,N_2720,N_3695);
or U6059 (N_6059,N_2506,N_4362);
nand U6060 (N_6060,N_3949,N_3432);
and U6061 (N_6061,N_3144,N_4211);
nor U6062 (N_6062,N_3488,N_4323);
or U6063 (N_6063,N_4958,N_4585);
nand U6064 (N_6064,N_3210,N_4788);
and U6065 (N_6065,N_3056,N_3439);
or U6066 (N_6066,N_4386,N_2674);
nand U6067 (N_6067,N_3574,N_3062);
nor U6068 (N_6068,N_2712,N_2700);
or U6069 (N_6069,N_3232,N_4929);
and U6070 (N_6070,N_3311,N_2671);
nor U6071 (N_6071,N_2964,N_3225);
nand U6072 (N_6072,N_2648,N_3581);
nand U6073 (N_6073,N_2507,N_2710);
nand U6074 (N_6074,N_3358,N_4338);
and U6075 (N_6075,N_4164,N_3306);
or U6076 (N_6076,N_3682,N_2547);
or U6077 (N_6077,N_2837,N_4389);
nand U6078 (N_6078,N_2638,N_4985);
nor U6079 (N_6079,N_3925,N_4974);
and U6080 (N_6080,N_2814,N_2959);
and U6081 (N_6081,N_2815,N_2909);
and U6082 (N_6082,N_2502,N_3668);
nor U6083 (N_6083,N_4679,N_3052);
or U6084 (N_6084,N_4360,N_2584);
nor U6085 (N_6085,N_3554,N_2982);
xor U6086 (N_6086,N_4177,N_4785);
nor U6087 (N_6087,N_4449,N_4393);
nand U6088 (N_6088,N_3929,N_4688);
nor U6089 (N_6089,N_2949,N_3867);
nor U6090 (N_6090,N_3914,N_4730);
and U6091 (N_6091,N_3314,N_4594);
or U6092 (N_6092,N_4922,N_3731);
and U6093 (N_6093,N_3174,N_3272);
or U6094 (N_6094,N_3304,N_4565);
nor U6095 (N_6095,N_4229,N_3035);
and U6096 (N_6096,N_3123,N_4531);
nand U6097 (N_6097,N_3467,N_4307);
nand U6098 (N_6098,N_3117,N_4562);
and U6099 (N_6099,N_3265,N_3871);
and U6100 (N_6100,N_3698,N_2948);
and U6101 (N_6101,N_3781,N_3943);
and U6102 (N_6102,N_3013,N_3785);
nor U6103 (N_6103,N_4141,N_3742);
nor U6104 (N_6104,N_2944,N_2905);
and U6105 (N_6105,N_3110,N_3339);
nand U6106 (N_6106,N_4111,N_2781);
nand U6107 (N_6107,N_3935,N_4220);
and U6108 (N_6108,N_3489,N_3812);
or U6109 (N_6109,N_4840,N_4082);
nor U6110 (N_6110,N_4138,N_3584);
nor U6111 (N_6111,N_4269,N_4769);
or U6112 (N_6112,N_3322,N_2990);
nand U6113 (N_6113,N_3767,N_4614);
or U6114 (N_6114,N_3771,N_4322);
and U6115 (N_6115,N_4777,N_4960);
nand U6116 (N_6116,N_4332,N_4078);
nor U6117 (N_6117,N_4115,N_2887);
or U6118 (N_6118,N_4800,N_2779);
nand U6119 (N_6119,N_3136,N_2858);
and U6120 (N_6120,N_2913,N_4372);
nand U6121 (N_6121,N_2574,N_3096);
or U6122 (N_6122,N_2667,N_4235);
nand U6123 (N_6123,N_4363,N_4143);
and U6124 (N_6124,N_3966,N_3230);
nor U6125 (N_6125,N_3705,N_2689);
nand U6126 (N_6126,N_4036,N_4287);
or U6127 (N_6127,N_3476,N_2681);
or U6128 (N_6128,N_4643,N_4267);
nor U6129 (N_6129,N_4735,N_4687);
and U6130 (N_6130,N_2643,N_3709);
or U6131 (N_6131,N_2709,N_3252);
or U6132 (N_6132,N_4887,N_4862);
or U6133 (N_6133,N_2673,N_4854);
and U6134 (N_6134,N_3253,N_2655);
nor U6135 (N_6135,N_3207,N_3788);
and U6136 (N_6136,N_3616,N_4042);
nand U6137 (N_6137,N_2715,N_3104);
or U6138 (N_6138,N_4906,N_3664);
and U6139 (N_6139,N_4611,N_3275);
or U6140 (N_6140,N_3663,N_4592);
nor U6141 (N_6141,N_4054,N_4265);
nand U6142 (N_6142,N_3679,N_4872);
nor U6143 (N_6143,N_3384,N_4354);
or U6144 (N_6144,N_3295,N_2874);
nor U6145 (N_6145,N_2979,N_2882);
nor U6146 (N_6146,N_3838,N_3217);
nand U6147 (N_6147,N_3881,N_4651);
nor U6148 (N_6148,N_4563,N_4488);
nor U6149 (N_6149,N_3733,N_3294);
and U6150 (N_6150,N_4715,N_3141);
or U6151 (N_6151,N_4767,N_3273);
nand U6152 (N_6152,N_4427,N_4221);
nor U6153 (N_6153,N_4699,N_4695);
and U6154 (N_6154,N_4121,N_3903);
and U6155 (N_6155,N_3201,N_2855);
and U6156 (N_6156,N_2853,N_2599);
nand U6157 (N_6157,N_3151,N_4689);
and U6158 (N_6158,N_4230,N_3888);
and U6159 (N_6159,N_3922,N_3055);
nand U6160 (N_6160,N_4546,N_4401);
or U6161 (N_6161,N_2997,N_3875);
or U6162 (N_6162,N_3349,N_3503);
and U6163 (N_6163,N_4670,N_4239);
or U6164 (N_6164,N_4724,N_2775);
nand U6165 (N_6165,N_3567,N_4075);
nor U6166 (N_6166,N_4953,N_3113);
xor U6167 (N_6167,N_3779,N_3457);
nand U6168 (N_6168,N_4142,N_4448);
nand U6169 (N_6169,N_4533,N_3923);
nor U6170 (N_6170,N_4426,N_3375);
or U6171 (N_6171,N_4039,N_2548);
nand U6172 (N_6172,N_4261,N_3783);
or U6173 (N_6173,N_4530,N_3919);
nor U6174 (N_6174,N_3135,N_4080);
or U6175 (N_6175,N_3341,N_4847);
nor U6176 (N_6176,N_3256,N_3305);
or U6177 (N_6177,N_4625,N_2687);
or U6178 (N_6178,N_3000,N_4994);
nand U6179 (N_6179,N_4431,N_2789);
or U6180 (N_6180,N_4011,N_3340);
nand U6181 (N_6181,N_3961,N_4983);
and U6182 (N_6182,N_4681,N_2576);
and U6183 (N_6183,N_4486,N_3636);
nand U6184 (N_6184,N_3408,N_4570);
nor U6185 (N_6185,N_4091,N_3362);
nor U6186 (N_6186,N_3009,N_3560);
nand U6187 (N_6187,N_2575,N_4266);
or U6188 (N_6188,N_4502,N_3652);
or U6189 (N_6189,N_2808,N_3047);
or U6190 (N_6190,N_3533,N_4738);
nand U6191 (N_6191,N_4403,N_3726);
nand U6192 (N_6192,N_2559,N_4704);
nor U6193 (N_6193,N_3513,N_3361);
nand U6194 (N_6194,N_3946,N_3671);
nor U6195 (N_6195,N_4956,N_3406);
nor U6196 (N_6196,N_3389,N_3543);
nand U6197 (N_6197,N_2620,N_3551);
nor U6198 (N_6198,N_3020,N_4596);
or U6199 (N_6199,N_4768,N_4076);
nor U6200 (N_6200,N_4991,N_2524);
nor U6201 (N_6201,N_3610,N_2947);
or U6202 (N_6202,N_4171,N_4911);
or U6203 (N_6203,N_3578,N_4331);
or U6204 (N_6204,N_4214,N_2557);
or U6205 (N_6205,N_3701,N_3236);
or U6206 (N_6206,N_4364,N_2838);
or U6207 (N_6207,N_4733,N_4120);
nor U6208 (N_6208,N_2752,N_3792);
or U6209 (N_6209,N_3185,N_3125);
or U6210 (N_6210,N_4988,N_4019);
nand U6211 (N_6211,N_4915,N_2517);
or U6212 (N_6212,N_4616,N_3019);
or U6213 (N_6213,N_4452,N_4281);
or U6214 (N_6214,N_2907,N_4729);
or U6215 (N_6215,N_3262,N_3050);
nand U6216 (N_6216,N_4224,N_2697);
or U6217 (N_6217,N_4521,N_4955);
or U6218 (N_6218,N_3960,N_3506);
nor U6219 (N_6219,N_4481,N_3081);
or U6220 (N_6220,N_3963,N_4146);
or U6221 (N_6221,N_2951,N_4270);
nor U6222 (N_6222,N_2679,N_4001);
and U6223 (N_6223,N_2619,N_4597);
nor U6224 (N_6224,N_4097,N_3916);
or U6225 (N_6225,N_2724,N_3958);
or U6226 (N_6226,N_3841,N_4703);
nand U6227 (N_6227,N_3281,N_4277);
nand U6228 (N_6228,N_4064,N_2705);
nor U6229 (N_6229,N_3851,N_3607);
or U6230 (N_6230,N_3524,N_4961);
nand U6231 (N_6231,N_4548,N_4808);
nor U6232 (N_6232,N_4525,N_3166);
nand U6233 (N_6233,N_4636,N_3654);
nor U6234 (N_6234,N_4203,N_3048);
nor U6235 (N_6235,N_4984,N_3114);
and U6236 (N_6236,N_4335,N_2590);
nor U6237 (N_6237,N_2573,N_2520);
nor U6238 (N_6238,N_2901,N_2536);
and U6239 (N_6239,N_4989,N_2745);
or U6240 (N_6240,N_3470,N_3153);
and U6241 (N_6241,N_3031,N_2790);
nand U6242 (N_6242,N_4384,N_3580);
nand U6243 (N_6243,N_4683,N_3205);
or U6244 (N_6244,N_2627,N_4250);
nand U6245 (N_6245,N_2768,N_2923);
and U6246 (N_6246,N_4535,N_4122);
and U6247 (N_6247,N_3005,N_4049);
and U6248 (N_6248,N_4089,N_2797);
and U6249 (N_6249,N_4711,N_3014);
or U6250 (N_6250,N_2555,N_3733);
or U6251 (N_6251,N_4602,N_2578);
and U6252 (N_6252,N_3307,N_2678);
and U6253 (N_6253,N_3451,N_4154);
nor U6254 (N_6254,N_3382,N_4064);
nor U6255 (N_6255,N_2778,N_3352);
and U6256 (N_6256,N_4873,N_4701);
nor U6257 (N_6257,N_2764,N_3773);
nand U6258 (N_6258,N_3488,N_3106);
and U6259 (N_6259,N_4290,N_3168);
or U6260 (N_6260,N_4502,N_3885);
nand U6261 (N_6261,N_2702,N_3868);
and U6262 (N_6262,N_4138,N_2879);
nand U6263 (N_6263,N_3103,N_4591);
or U6264 (N_6264,N_4849,N_2543);
nand U6265 (N_6265,N_4829,N_4711);
xnor U6266 (N_6266,N_4437,N_3459);
and U6267 (N_6267,N_4487,N_3586);
and U6268 (N_6268,N_4234,N_3086);
nor U6269 (N_6269,N_3130,N_3281);
nand U6270 (N_6270,N_2849,N_4521);
or U6271 (N_6271,N_3870,N_3534);
and U6272 (N_6272,N_4463,N_3932);
or U6273 (N_6273,N_3500,N_4674);
or U6274 (N_6274,N_3204,N_2889);
nor U6275 (N_6275,N_4467,N_4187);
nand U6276 (N_6276,N_4243,N_3680);
nor U6277 (N_6277,N_3219,N_3463);
or U6278 (N_6278,N_3216,N_2880);
nand U6279 (N_6279,N_4795,N_4580);
nor U6280 (N_6280,N_2636,N_2993);
nand U6281 (N_6281,N_4475,N_3350);
or U6282 (N_6282,N_3791,N_4440);
or U6283 (N_6283,N_4700,N_4872);
nand U6284 (N_6284,N_4214,N_4305);
or U6285 (N_6285,N_4011,N_3636);
nor U6286 (N_6286,N_3543,N_2839);
nand U6287 (N_6287,N_4090,N_4252);
xor U6288 (N_6288,N_3316,N_4959);
nor U6289 (N_6289,N_4562,N_3223);
nor U6290 (N_6290,N_3648,N_4932);
and U6291 (N_6291,N_3260,N_3003);
nand U6292 (N_6292,N_4222,N_3673);
and U6293 (N_6293,N_3883,N_3272);
and U6294 (N_6294,N_4819,N_3173);
and U6295 (N_6295,N_4360,N_3836);
nand U6296 (N_6296,N_4768,N_2827);
or U6297 (N_6297,N_3472,N_4107);
or U6298 (N_6298,N_3479,N_4338);
or U6299 (N_6299,N_2763,N_4840);
and U6300 (N_6300,N_2663,N_4444);
and U6301 (N_6301,N_3686,N_3765);
or U6302 (N_6302,N_3652,N_2517);
and U6303 (N_6303,N_4043,N_3748);
or U6304 (N_6304,N_3963,N_2920);
or U6305 (N_6305,N_4273,N_4151);
or U6306 (N_6306,N_3432,N_4058);
nor U6307 (N_6307,N_4909,N_4310);
nor U6308 (N_6308,N_3792,N_2870);
or U6309 (N_6309,N_4573,N_3709);
and U6310 (N_6310,N_4590,N_3538);
nor U6311 (N_6311,N_4457,N_3214);
or U6312 (N_6312,N_3806,N_3223);
or U6313 (N_6313,N_2534,N_3848);
or U6314 (N_6314,N_4968,N_4400);
nand U6315 (N_6315,N_3907,N_3238);
nor U6316 (N_6316,N_4473,N_2786);
nor U6317 (N_6317,N_4603,N_3941);
nor U6318 (N_6318,N_4582,N_3955);
nor U6319 (N_6319,N_2767,N_3133);
nand U6320 (N_6320,N_3133,N_2723);
nand U6321 (N_6321,N_4783,N_3194);
or U6322 (N_6322,N_3263,N_4591);
and U6323 (N_6323,N_2890,N_3262);
or U6324 (N_6324,N_4146,N_2542);
nor U6325 (N_6325,N_3672,N_3388);
nor U6326 (N_6326,N_2659,N_3325);
or U6327 (N_6327,N_3396,N_2873);
and U6328 (N_6328,N_3319,N_4840);
or U6329 (N_6329,N_2508,N_3932);
nand U6330 (N_6330,N_4889,N_3477);
nor U6331 (N_6331,N_4541,N_4766);
nand U6332 (N_6332,N_2887,N_2890);
nor U6333 (N_6333,N_4605,N_3253);
nand U6334 (N_6334,N_3794,N_3306);
or U6335 (N_6335,N_3398,N_2779);
nor U6336 (N_6336,N_3063,N_4225);
and U6337 (N_6337,N_4550,N_4457);
nand U6338 (N_6338,N_3204,N_4096);
nor U6339 (N_6339,N_3541,N_4187);
or U6340 (N_6340,N_4359,N_4184);
and U6341 (N_6341,N_4660,N_4727);
or U6342 (N_6342,N_4719,N_3073);
and U6343 (N_6343,N_2531,N_3068);
nand U6344 (N_6344,N_3187,N_4253);
nand U6345 (N_6345,N_3251,N_4680);
or U6346 (N_6346,N_2530,N_3918);
nor U6347 (N_6347,N_3824,N_3315);
or U6348 (N_6348,N_3355,N_3912);
and U6349 (N_6349,N_4228,N_3069);
or U6350 (N_6350,N_3731,N_2771);
or U6351 (N_6351,N_3458,N_2921);
and U6352 (N_6352,N_3472,N_3624);
or U6353 (N_6353,N_4122,N_4149);
or U6354 (N_6354,N_3575,N_3062);
nand U6355 (N_6355,N_3716,N_4416);
nand U6356 (N_6356,N_2695,N_2890);
or U6357 (N_6357,N_4668,N_2953);
or U6358 (N_6358,N_3597,N_3310);
nor U6359 (N_6359,N_2903,N_2765);
nand U6360 (N_6360,N_2942,N_3748);
and U6361 (N_6361,N_3645,N_3627);
nor U6362 (N_6362,N_2715,N_3368);
or U6363 (N_6363,N_3907,N_3491);
nand U6364 (N_6364,N_4328,N_3615);
or U6365 (N_6365,N_3656,N_4508);
nand U6366 (N_6366,N_2984,N_2584);
nand U6367 (N_6367,N_3514,N_3223);
nor U6368 (N_6368,N_3417,N_4843);
nor U6369 (N_6369,N_4967,N_3559);
nand U6370 (N_6370,N_4295,N_3364);
nor U6371 (N_6371,N_3619,N_3893);
and U6372 (N_6372,N_4295,N_4498);
or U6373 (N_6373,N_2982,N_2930);
or U6374 (N_6374,N_4988,N_4707);
or U6375 (N_6375,N_4021,N_2847);
nand U6376 (N_6376,N_3486,N_3795);
nand U6377 (N_6377,N_3642,N_4106);
nand U6378 (N_6378,N_3006,N_4315);
or U6379 (N_6379,N_3230,N_4795);
nor U6380 (N_6380,N_2697,N_3804);
nand U6381 (N_6381,N_2682,N_4866);
nor U6382 (N_6382,N_4934,N_3535);
or U6383 (N_6383,N_2968,N_3556);
and U6384 (N_6384,N_3750,N_4678);
nor U6385 (N_6385,N_4446,N_4095);
nor U6386 (N_6386,N_3346,N_2768);
nand U6387 (N_6387,N_3726,N_4715);
and U6388 (N_6388,N_3288,N_3470);
and U6389 (N_6389,N_4837,N_2781);
nor U6390 (N_6390,N_3861,N_3431);
or U6391 (N_6391,N_3434,N_4399);
nand U6392 (N_6392,N_2543,N_3687);
nand U6393 (N_6393,N_3795,N_3294);
and U6394 (N_6394,N_2903,N_3706);
or U6395 (N_6395,N_3701,N_4047);
nand U6396 (N_6396,N_3935,N_2592);
nor U6397 (N_6397,N_2813,N_3350);
or U6398 (N_6398,N_2837,N_4125);
and U6399 (N_6399,N_3340,N_2720);
or U6400 (N_6400,N_4147,N_3980);
or U6401 (N_6401,N_4065,N_3859);
and U6402 (N_6402,N_3167,N_4560);
nor U6403 (N_6403,N_3202,N_2628);
nand U6404 (N_6404,N_3986,N_4568);
and U6405 (N_6405,N_3299,N_4835);
xnor U6406 (N_6406,N_3995,N_3215);
xor U6407 (N_6407,N_3709,N_2599);
nor U6408 (N_6408,N_2882,N_3336);
or U6409 (N_6409,N_3853,N_4000);
nand U6410 (N_6410,N_4314,N_3495);
and U6411 (N_6411,N_3302,N_3288);
and U6412 (N_6412,N_3698,N_3484);
nor U6413 (N_6413,N_4589,N_4718);
or U6414 (N_6414,N_2594,N_4986);
nand U6415 (N_6415,N_4832,N_4899);
and U6416 (N_6416,N_3306,N_2625);
nand U6417 (N_6417,N_4213,N_4424);
or U6418 (N_6418,N_3570,N_3196);
nor U6419 (N_6419,N_2902,N_4007);
or U6420 (N_6420,N_3006,N_4819);
nand U6421 (N_6421,N_4526,N_4415);
and U6422 (N_6422,N_3170,N_2639);
or U6423 (N_6423,N_3470,N_3106);
nor U6424 (N_6424,N_2543,N_4222);
or U6425 (N_6425,N_4372,N_3887);
and U6426 (N_6426,N_3692,N_3310);
nor U6427 (N_6427,N_4420,N_4697);
and U6428 (N_6428,N_3507,N_4472);
nor U6429 (N_6429,N_3595,N_4639);
and U6430 (N_6430,N_2577,N_3301);
or U6431 (N_6431,N_2544,N_3705);
nand U6432 (N_6432,N_2561,N_3039);
nand U6433 (N_6433,N_2872,N_4259);
and U6434 (N_6434,N_3927,N_2572);
or U6435 (N_6435,N_4144,N_4491);
nand U6436 (N_6436,N_3814,N_4522);
and U6437 (N_6437,N_3154,N_4198);
or U6438 (N_6438,N_4590,N_4484);
and U6439 (N_6439,N_4123,N_3846);
and U6440 (N_6440,N_3829,N_4638);
nand U6441 (N_6441,N_4084,N_3921);
or U6442 (N_6442,N_2655,N_4467);
nor U6443 (N_6443,N_3714,N_4215);
and U6444 (N_6444,N_4153,N_2865);
or U6445 (N_6445,N_2877,N_4330);
and U6446 (N_6446,N_4600,N_4086);
and U6447 (N_6447,N_4617,N_3649);
xor U6448 (N_6448,N_3612,N_4224);
nand U6449 (N_6449,N_2847,N_3821);
and U6450 (N_6450,N_3199,N_3239);
and U6451 (N_6451,N_4350,N_4624);
nand U6452 (N_6452,N_4046,N_3693);
xor U6453 (N_6453,N_4628,N_3101);
nor U6454 (N_6454,N_3404,N_2844);
or U6455 (N_6455,N_4747,N_3898);
and U6456 (N_6456,N_4162,N_2526);
and U6457 (N_6457,N_3825,N_3815);
and U6458 (N_6458,N_4888,N_3854);
or U6459 (N_6459,N_4120,N_4530);
and U6460 (N_6460,N_4341,N_4605);
or U6461 (N_6461,N_2636,N_3561);
and U6462 (N_6462,N_2669,N_3549);
nor U6463 (N_6463,N_4075,N_3080);
nor U6464 (N_6464,N_4404,N_3902);
nand U6465 (N_6465,N_4346,N_4753);
nand U6466 (N_6466,N_4705,N_4348);
nor U6467 (N_6467,N_4907,N_4208);
nand U6468 (N_6468,N_4842,N_2983);
nor U6469 (N_6469,N_2836,N_3325);
nor U6470 (N_6470,N_4930,N_4772);
or U6471 (N_6471,N_4323,N_4526);
or U6472 (N_6472,N_3201,N_3812);
or U6473 (N_6473,N_2797,N_2634);
and U6474 (N_6474,N_3633,N_3064);
or U6475 (N_6475,N_4885,N_3552);
nor U6476 (N_6476,N_4720,N_4318);
nand U6477 (N_6477,N_3866,N_3982);
nor U6478 (N_6478,N_4172,N_4762);
nand U6479 (N_6479,N_3977,N_3190);
and U6480 (N_6480,N_3342,N_3282);
or U6481 (N_6481,N_4473,N_2744);
nor U6482 (N_6482,N_3858,N_3789);
or U6483 (N_6483,N_3997,N_3058);
nor U6484 (N_6484,N_4625,N_3818);
or U6485 (N_6485,N_3386,N_3063);
or U6486 (N_6486,N_3344,N_3197);
nand U6487 (N_6487,N_2517,N_4351);
nor U6488 (N_6488,N_3672,N_3997);
or U6489 (N_6489,N_4942,N_3245);
and U6490 (N_6490,N_3609,N_4362);
nor U6491 (N_6491,N_2950,N_4477);
or U6492 (N_6492,N_3519,N_2595);
and U6493 (N_6493,N_3700,N_3524);
nand U6494 (N_6494,N_2638,N_3930);
nand U6495 (N_6495,N_2550,N_4952);
nand U6496 (N_6496,N_4765,N_4526);
nor U6497 (N_6497,N_4339,N_3400);
and U6498 (N_6498,N_3107,N_2666);
nand U6499 (N_6499,N_4205,N_4242);
nand U6500 (N_6500,N_3695,N_3766);
nor U6501 (N_6501,N_4411,N_3211);
nor U6502 (N_6502,N_2923,N_3489);
nand U6503 (N_6503,N_4855,N_4716);
or U6504 (N_6504,N_2792,N_4633);
nor U6505 (N_6505,N_2941,N_3084);
nor U6506 (N_6506,N_4848,N_4337);
nor U6507 (N_6507,N_2572,N_3007);
nor U6508 (N_6508,N_3586,N_4647);
nand U6509 (N_6509,N_4518,N_4829);
nor U6510 (N_6510,N_3274,N_2847);
nor U6511 (N_6511,N_4974,N_3172);
or U6512 (N_6512,N_4049,N_3095);
nand U6513 (N_6513,N_3795,N_3411);
or U6514 (N_6514,N_3810,N_2917);
and U6515 (N_6515,N_4062,N_3564);
nand U6516 (N_6516,N_4515,N_4428);
or U6517 (N_6517,N_3491,N_4958);
and U6518 (N_6518,N_4534,N_3538);
or U6519 (N_6519,N_4890,N_2904);
nor U6520 (N_6520,N_2948,N_2770);
nor U6521 (N_6521,N_4976,N_3184);
nor U6522 (N_6522,N_3740,N_3417);
and U6523 (N_6523,N_4287,N_4989);
and U6524 (N_6524,N_4030,N_3352);
nor U6525 (N_6525,N_4201,N_3849);
nand U6526 (N_6526,N_2570,N_4273);
nand U6527 (N_6527,N_3787,N_2835);
or U6528 (N_6528,N_2852,N_4204);
nor U6529 (N_6529,N_3219,N_2583);
or U6530 (N_6530,N_2711,N_4843);
or U6531 (N_6531,N_2900,N_4030);
nand U6532 (N_6532,N_3966,N_4988);
and U6533 (N_6533,N_4842,N_4615);
nor U6534 (N_6534,N_3345,N_4531);
nand U6535 (N_6535,N_2558,N_3032);
nand U6536 (N_6536,N_3363,N_4968);
or U6537 (N_6537,N_4277,N_2555);
nand U6538 (N_6538,N_3576,N_2668);
or U6539 (N_6539,N_2634,N_3561);
nor U6540 (N_6540,N_3517,N_3046);
or U6541 (N_6541,N_2973,N_4974);
nand U6542 (N_6542,N_2915,N_3143);
or U6543 (N_6543,N_4168,N_3235);
nor U6544 (N_6544,N_2608,N_4379);
nor U6545 (N_6545,N_2824,N_4266);
or U6546 (N_6546,N_3498,N_3417);
or U6547 (N_6547,N_3477,N_4244);
or U6548 (N_6548,N_2725,N_2600);
nand U6549 (N_6549,N_3310,N_2971);
nand U6550 (N_6550,N_4813,N_3984);
nor U6551 (N_6551,N_3193,N_4586);
and U6552 (N_6552,N_4914,N_4260);
nor U6553 (N_6553,N_4020,N_4623);
or U6554 (N_6554,N_3595,N_3320);
nand U6555 (N_6555,N_3674,N_3420);
and U6556 (N_6556,N_4287,N_4240);
nand U6557 (N_6557,N_3673,N_4636);
or U6558 (N_6558,N_3949,N_3104);
or U6559 (N_6559,N_4873,N_3263);
xor U6560 (N_6560,N_3793,N_2966);
nand U6561 (N_6561,N_4561,N_4308);
nor U6562 (N_6562,N_4965,N_3389);
and U6563 (N_6563,N_3003,N_3420);
nor U6564 (N_6564,N_3577,N_3095);
nand U6565 (N_6565,N_3869,N_3188);
nand U6566 (N_6566,N_3809,N_3835);
and U6567 (N_6567,N_3600,N_3747);
and U6568 (N_6568,N_3903,N_2525);
and U6569 (N_6569,N_4531,N_2737);
nand U6570 (N_6570,N_3380,N_4212);
or U6571 (N_6571,N_4856,N_4586);
nand U6572 (N_6572,N_4532,N_2645);
nor U6573 (N_6573,N_3792,N_3361);
or U6574 (N_6574,N_3221,N_2749);
and U6575 (N_6575,N_3303,N_3240);
nor U6576 (N_6576,N_4492,N_3305);
nand U6577 (N_6577,N_3582,N_2748);
and U6578 (N_6578,N_4214,N_4331);
nand U6579 (N_6579,N_2658,N_3926);
or U6580 (N_6580,N_4861,N_3165);
and U6581 (N_6581,N_3061,N_4852);
nor U6582 (N_6582,N_4334,N_2762);
nor U6583 (N_6583,N_4371,N_3568);
and U6584 (N_6584,N_4271,N_4248);
nor U6585 (N_6585,N_4520,N_3505);
or U6586 (N_6586,N_2521,N_3486);
and U6587 (N_6587,N_4488,N_4545);
nor U6588 (N_6588,N_4218,N_4437);
nor U6589 (N_6589,N_3721,N_3487);
and U6590 (N_6590,N_4172,N_2619);
nor U6591 (N_6591,N_3969,N_2680);
nand U6592 (N_6592,N_3877,N_3926);
nor U6593 (N_6593,N_4637,N_2700);
or U6594 (N_6594,N_3397,N_2591);
or U6595 (N_6595,N_3302,N_2850);
nor U6596 (N_6596,N_4203,N_3013);
and U6597 (N_6597,N_4496,N_4615);
nand U6598 (N_6598,N_4154,N_4325);
and U6599 (N_6599,N_4776,N_2803);
or U6600 (N_6600,N_3985,N_3325);
nor U6601 (N_6601,N_2735,N_3547);
nor U6602 (N_6602,N_2894,N_3565);
nor U6603 (N_6603,N_2629,N_4127);
nand U6604 (N_6604,N_4311,N_4899);
nor U6605 (N_6605,N_2897,N_3756);
nor U6606 (N_6606,N_2607,N_3481);
nor U6607 (N_6607,N_3790,N_4701);
nand U6608 (N_6608,N_3292,N_4562);
xor U6609 (N_6609,N_4391,N_4319);
or U6610 (N_6610,N_4494,N_4880);
or U6611 (N_6611,N_2804,N_2715);
or U6612 (N_6612,N_2548,N_3723);
or U6613 (N_6613,N_4890,N_3267);
and U6614 (N_6614,N_4186,N_4712);
or U6615 (N_6615,N_3907,N_2783);
nor U6616 (N_6616,N_3367,N_3117);
nor U6617 (N_6617,N_2651,N_3677);
nand U6618 (N_6618,N_2645,N_2953);
nand U6619 (N_6619,N_4448,N_3170);
or U6620 (N_6620,N_4028,N_4997);
nand U6621 (N_6621,N_4578,N_2941);
and U6622 (N_6622,N_4806,N_2793);
or U6623 (N_6623,N_3873,N_3339);
nor U6624 (N_6624,N_2610,N_3520);
nor U6625 (N_6625,N_4788,N_4036);
nand U6626 (N_6626,N_4749,N_3657);
and U6627 (N_6627,N_3589,N_2708);
nand U6628 (N_6628,N_3348,N_4583);
nand U6629 (N_6629,N_3487,N_3802);
or U6630 (N_6630,N_3481,N_4311);
and U6631 (N_6631,N_3548,N_3995);
nand U6632 (N_6632,N_4415,N_3539);
nor U6633 (N_6633,N_3134,N_4142);
nor U6634 (N_6634,N_2812,N_2972);
nand U6635 (N_6635,N_3754,N_4721);
or U6636 (N_6636,N_4442,N_4623);
nor U6637 (N_6637,N_3105,N_3801);
and U6638 (N_6638,N_3960,N_3768);
and U6639 (N_6639,N_2900,N_2873);
or U6640 (N_6640,N_3722,N_4802);
and U6641 (N_6641,N_2634,N_3747);
and U6642 (N_6642,N_4600,N_4585);
nand U6643 (N_6643,N_2618,N_2677);
and U6644 (N_6644,N_4615,N_3233);
or U6645 (N_6645,N_4591,N_3309);
nand U6646 (N_6646,N_3868,N_2726);
nand U6647 (N_6647,N_2725,N_3410);
nand U6648 (N_6648,N_3512,N_2677);
nor U6649 (N_6649,N_3731,N_3968);
nor U6650 (N_6650,N_3609,N_3507);
and U6651 (N_6651,N_4016,N_4037);
and U6652 (N_6652,N_4563,N_3393);
nand U6653 (N_6653,N_4937,N_3081);
and U6654 (N_6654,N_4168,N_3019);
or U6655 (N_6655,N_3853,N_4324);
and U6656 (N_6656,N_3680,N_2932);
nor U6657 (N_6657,N_4012,N_4889);
and U6658 (N_6658,N_3216,N_2943);
nand U6659 (N_6659,N_2684,N_4602);
and U6660 (N_6660,N_3475,N_4622);
nand U6661 (N_6661,N_4903,N_4948);
nor U6662 (N_6662,N_4766,N_4333);
nor U6663 (N_6663,N_4994,N_4363);
nor U6664 (N_6664,N_4668,N_3861);
and U6665 (N_6665,N_3559,N_3082);
and U6666 (N_6666,N_4290,N_2810);
or U6667 (N_6667,N_4825,N_4659);
or U6668 (N_6668,N_3484,N_4602);
and U6669 (N_6669,N_3685,N_3687);
or U6670 (N_6670,N_4449,N_3844);
and U6671 (N_6671,N_4424,N_3327);
nand U6672 (N_6672,N_4881,N_4406);
and U6673 (N_6673,N_4676,N_4438);
nand U6674 (N_6674,N_4643,N_4405);
and U6675 (N_6675,N_3893,N_3794);
nand U6676 (N_6676,N_3002,N_4237);
and U6677 (N_6677,N_3559,N_2901);
or U6678 (N_6678,N_4885,N_3468);
nand U6679 (N_6679,N_4146,N_4635);
nand U6680 (N_6680,N_4894,N_4059);
nand U6681 (N_6681,N_2757,N_2603);
nor U6682 (N_6682,N_4181,N_3413);
or U6683 (N_6683,N_4888,N_2557);
or U6684 (N_6684,N_4833,N_4818);
or U6685 (N_6685,N_3653,N_3811);
or U6686 (N_6686,N_2677,N_4599);
nor U6687 (N_6687,N_4130,N_4949);
and U6688 (N_6688,N_2617,N_4847);
or U6689 (N_6689,N_4565,N_4488);
xor U6690 (N_6690,N_4180,N_4708);
and U6691 (N_6691,N_4762,N_4565);
and U6692 (N_6692,N_4668,N_2711);
or U6693 (N_6693,N_3848,N_3799);
and U6694 (N_6694,N_2846,N_2976);
nand U6695 (N_6695,N_4428,N_4395);
or U6696 (N_6696,N_3493,N_4116);
nor U6697 (N_6697,N_3504,N_4482);
nor U6698 (N_6698,N_4959,N_4128);
or U6699 (N_6699,N_4434,N_4917);
nand U6700 (N_6700,N_4052,N_3771);
and U6701 (N_6701,N_2865,N_4096);
nor U6702 (N_6702,N_4788,N_4911);
nand U6703 (N_6703,N_2518,N_3252);
nand U6704 (N_6704,N_4759,N_4639);
and U6705 (N_6705,N_4478,N_3567);
or U6706 (N_6706,N_3226,N_4968);
nand U6707 (N_6707,N_3589,N_4585);
nand U6708 (N_6708,N_3300,N_4702);
nor U6709 (N_6709,N_4895,N_4088);
or U6710 (N_6710,N_4039,N_4453);
and U6711 (N_6711,N_3502,N_4688);
or U6712 (N_6712,N_3526,N_3272);
and U6713 (N_6713,N_3589,N_4464);
or U6714 (N_6714,N_4208,N_3347);
nor U6715 (N_6715,N_2845,N_3198);
nor U6716 (N_6716,N_2935,N_4119);
nor U6717 (N_6717,N_4163,N_2786);
nand U6718 (N_6718,N_4551,N_4005);
or U6719 (N_6719,N_4923,N_2518);
nand U6720 (N_6720,N_3737,N_4585);
nand U6721 (N_6721,N_3526,N_4595);
or U6722 (N_6722,N_3672,N_2539);
nor U6723 (N_6723,N_2933,N_4450);
and U6724 (N_6724,N_3760,N_2852);
nor U6725 (N_6725,N_3619,N_3435);
nand U6726 (N_6726,N_4570,N_4711);
and U6727 (N_6727,N_3916,N_4045);
and U6728 (N_6728,N_3289,N_3458);
nand U6729 (N_6729,N_4035,N_2530);
nor U6730 (N_6730,N_4549,N_2924);
and U6731 (N_6731,N_2798,N_4439);
and U6732 (N_6732,N_3774,N_2614);
and U6733 (N_6733,N_3453,N_4343);
nor U6734 (N_6734,N_2744,N_4527);
and U6735 (N_6735,N_4932,N_4315);
nand U6736 (N_6736,N_3389,N_4145);
nand U6737 (N_6737,N_4747,N_2733);
nand U6738 (N_6738,N_4698,N_3438);
nand U6739 (N_6739,N_3699,N_4027);
nor U6740 (N_6740,N_4074,N_4737);
or U6741 (N_6741,N_3897,N_4493);
nand U6742 (N_6742,N_2765,N_4547);
nand U6743 (N_6743,N_3779,N_3599);
nand U6744 (N_6744,N_4744,N_2526);
or U6745 (N_6745,N_4048,N_4074);
nor U6746 (N_6746,N_3458,N_3102);
nand U6747 (N_6747,N_4414,N_4654);
nand U6748 (N_6748,N_4807,N_4875);
nand U6749 (N_6749,N_2830,N_4426);
nand U6750 (N_6750,N_3780,N_4561);
nor U6751 (N_6751,N_4890,N_4007);
nand U6752 (N_6752,N_3176,N_3097);
and U6753 (N_6753,N_3277,N_4705);
or U6754 (N_6754,N_3193,N_2892);
and U6755 (N_6755,N_3460,N_2655);
or U6756 (N_6756,N_2997,N_2981);
or U6757 (N_6757,N_4313,N_4166);
or U6758 (N_6758,N_3665,N_3857);
or U6759 (N_6759,N_4056,N_3697);
nor U6760 (N_6760,N_2529,N_2823);
nor U6761 (N_6761,N_4609,N_4197);
nor U6762 (N_6762,N_2761,N_3488);
and U6763 (N_6763,N_3611,N_3756);
and U6764 (N_6764,N_3629,N_4940);
or U6765 (N_6765,N_3304,N_4119);
nand U6766 (N_6766,N_4160,N_4020);
nand U6767 (N_6767,N_4344,N_3153);
nand U6768 (N_6768,N_3701,N_3243);
or U6769 (N_6769,N_3516,N_2950);
or U6770 (N_6770,N_3367,N_4153);
or U6771 (N_6771,N_4440,N_3902);
nand U6772 (N_6772,N_3231,N_4940);
or U6773 (N_6773,N_4011,N_2615);
and U6774 (N_6774,N_4954,N_3141);
and U6775 (N_6775,N_3945,N_4473);
and U6776 (N_6776,N_4318,N_4358);
or U6777 (N_6777,N_3851,N_3505);
and U6778 (N_6778,N_4229,N_4468);
or U6779 (N_6779,N_3185,N_4018);
or U6780 (N_6780,N_2566,N_3241);
and U6781 (N_6781,N_3221,N_4826);
nand U6782 (N_6782,N_4120,N_4503);
nor U6783 (N_6783,N_4274,N_3281);
nand U6784 (N_6784,N_3006,N_3444);
and U6785 (N_6785,N_2886,N_4585);
and U6786 (N_6786,N_4938,N_4882);
and U6787 (N_6787,N_3340,N_4267);
nor U6788 (N_6788,N_4834,N_3801);
nor U6789 (N_6789,N_4467,N_4689);
nand U6790 (N_6790,N_4889,N_4978);
nand U6791 (N_6791,N_3950,N_2779);
nand U6792 (N_6792,N_4287,N_3797);
and U6793 (N_6793,N_4690,N_4678);
nor U6794 (N_6794,N_3117,N_4780);
nor U6795 (N_6795,N_2973,N_4138);
nand U6796 (N_6796,N_3342,N_3201);
or U6797 (N_6797,N_4317,N_3349);
nand U6798 (N_6798,N_4550,N_3088);
and U6799 (N_6799,N_4210,N_3811);
nor U6800 (N_6800,N_3969,N_2549);
nand U6801 (N_6801,N_4286,N_3828);
nand U6802 (N_6802,N_4569,N_4199);
nor U6803 (N_6803,N_3451,N_2964);
nand U6804 (N_6804,N_4782,N_3508);
nor U6805 (N_6805,N_2660,N_4644);
nand U6806 (N_6806,N_3797,N_4931);
or U6807 (N_6807,N_4109,N_3176);
nor U6808 (N_6808,N_4812,N_4307);
or U6809 (N_6809,N_2929,N_2595);
or U6810 (N_6810,N_4147,N_3116);
and U6811 (N_6811,N_3438,N_4226);
or U6812 (N_6812,N_2894,N_2833);
nand U6813 (N_6813,N_3877,N_4131);
nand U6814 (N_6814,N_3150,N_4057);
nand U6815 (N_6815,N_4915,N_4491);
or U6816 (N_6816,N_4948,N_4681);
or U6817 (N_6817,N_3090,N_4210);
nand U6818 (N_6818,N_3884,N_4046);
nor U6819 (N_6819,N_3117,N_3133);
and U6820 (N_6820,N_4837,N_4298);
nand U6821 (N_6821,N_3998,N_4778);
nand U6822 (N_6822,N_3690,N_4197);
nand U6823 (N_6823,N_3528,N_4919);
nor U6824 (N_6824,N_4078,N_3932);
nor U6825 (N_6825,N_3137,N_2773);
or U6826 (N_6826,N_4719,N_2671);
nand U6827 (N_6827,N_3719,N_4279);
or U6828 (N_6828,N_3169,N_4966);
nor U6829 (N_6829,N_2674,N_4845);
or U6830 (N_6830,N_4753,N_3854);
nor U6831 (N_6831,N_3390,N_4763);
and U6832 (N_6832,N_3898,N_3748);
and U6833 (N_6833,N_4811,N_3877);
nand U6834 (N_6834,N_3847,N_2512);
and U6835 (N_6835,N_4356,N_3248);
nor U6836 (N_6836,N_4822,N_2564);
and U6837 (N_6837,N_4493,N_2976);
nand U6838 (N_6838,N_3541,N_4743);
or U6839 (N_6839,N_3476,N_4108);
and U6840 (N_6840,N_3336,N_3801);
nand U6841 (N_6841,N_2991,N_3098);
or U6842 (N_6842,N_2789,N_2719);
and U6843 (N_6843,N_3535,N_4073);
or U6844 (N_6844,N_3484,N_4403);
and U6845 (N_6845,N_3869,N_3868);
xor U6846 (N_6846,N_3523,N_4187);
nand U6847 (N_6847,N_4336,N_2973);
or U6848 (N_6848,N_2987,N_4787);
nand U6849 (N_6849,N_3563,N_3694);
and U6850 (N_6850,N_4968,N_3279);
nand U6851 (N_6851,N_4464,N_2588);
nor U6852 (N_6852,N_2573,N_3736);
or U6853 (N_6853,N_2903,N_4640);
nand U6854 (N_6854,N_3233,N_3042);
and U6855 (N_6855,N_3299,N_4621);
or U6856 (N_6856,N_3198,N_3354);
nand U6857 (N_6857,N_2836,N_3479);
nor U6858 (N_6858,N_4722,N_3700);
or U6859 (N_6859,N_4449,N_4122);
or U6860 (N_6860,N_3338,N_4404);
and U6861 (N_6861,N_2793,N_3492);
nor U6862 (N_6862,N_3493,N_3286);
nand U6863 (N_6863,N_4206,N_3031);
and U6864 (N_6864,N_2984,N_3651);
nand U6865 (N_6865,N_2936,N_3720);
nor U6866 (N_6866,N_3603,N_3666);
or U6867 (N_6867,N_4192,N_2518);
and U6868 (N_6868,N_4920,N_4057);
or U6869 (N_6869,N_2535,N_4862);
or U6870 (N_6870,N_4270,N_2576);
or U6871 (N_6871,N_4887,N_4589);
and U6872 (N_6872,N_3065,N_3835);
or U6873 (N_6873,N_3076,N_3786);
and U6874 (N_6874,N_3876,N_3047);
or U6875 (N_6875,N_3094,N_3596);
and U6876 (N_6876,N_4090,N_3489);
and U6877 (N_6877,N_3026,N_4947);
nor U6878 (N_6878,N_4154,N_4608);
nor U6879 (N_6879,N_3902,N_4279);
nand U6880 (N_6880,N_4585,N_4832);
nor U6881 (N_6881,N_3465,N_3396);
nor U6882 (N_6882,N_4574,N_3233);
and U6883 (N_6883,N_4681,N_4361);
nand U6884 (N_6884,N_4195,N_4834);
nand U6885 (N_6885,N_4988,N_4182);
nand U6886 (N_6886,N_2761,N_3474);
nor U6887 (N_6887,N_2867,N_3439);
and U6888 (N_6888,N_4346,N_3437);
and U6889 (N_6889,N_4938,N_3117);
or U6890 (N_6890,N_3586,N_4911);
nor U6891 (N_6891,N_4135,N_3405);
nand U6892 (N_6892,N_4553,N_4017);
nor U6893 (N_6893,N_3435,N_3873);
and U6894 (N_6894,N_3792,N_4683);
nand U6895 (N_6895,N_3233,N_4128);
nand U6896 (N_6896,N_2871,N_2619);
xor U6897 (N_6897,N_2917,N_4406);
nor U6898 (N_6898,N_2897,N_3458);
xnor U6899 (N_6899,N_4679,N_2796);
or U6900 (N_6900,N_4254,N_4361);
or U6901 (N_6901,N_3232,N_4642);
or U6902 (N_6902,N_4061,N_4710);
or U6903 (N_6903,N_4183,N_3230);
and U6904 (N_6904,N_2977,N_3773);
nor U6905 (N_6905,N_3564,N_2932);
nor U6906 (N_6906,N_3939,N_4473);
nor U6907 (N_6907,N_4104,N_4998);
or U6908 (N_6908,N_4453,N_3194);
nand U6909 (N_6909,N_4524,N_3584);
or U6910 (N_6910,N_4754,N_4203);
nand U6911 (N_6911,N_4601,N_4841);
nor U6912 (N_6912,N_4135,N_2768);
nand U6913 (N_6913,N_4944,N_2856);
and U6914 (N_6914,N_4528,N_2855);
nand U6915 (N_6915,N_4283,N_2747);
and U6916 (N_6916,N_4057,N_2931);
nor U6917 (N_6917,N_3509,N_4251);
nor U6918 (N_6918,N_2938,N_4125);
or U6919 (N_6919,N_4182,N_3692);
and U6920 (N_6920,N_3453,N_2893);
and U6921 (N_6921,N_2691,N_4634);
nand U6922 (N_6922,N_2805,N_3763);
and U6923 (N_6923,N_2546,N_4699);
nor U6924 (N_6924,N_4249,N_2972);
nor U6925 (N_6925,N_4139,N_3963);
nand U6926 (N_6926,N_3811,N_3634);
nor U6927 (N_6927,N_2549,N_3228);
and U6928 (N_6928,N_3561,N_3983);
nand U6929 (N_6929,N_4759,N_3419);
nand U6930 (N_6930,N_3336,N_3474);
nor U6931 (N_6931,N_4733,N_3551);
nand U6932 (N_6932,N_2616,N_2930);
or U6933 (N_6933,N_2894,N_2846);
and U6934 (N_6934,N_4616,N_3508);
nor U6935 (N_6935,N_3380,N_2605);
nor U6936 (N_6936,N_4835,N_3082);
nand U6937 (N_6937,N_4835,N_3929);
and U6938 (N_6938,N_4754,N_3549);
nor U6939 (N_6939,N_4457,N_3364);
and U6940 (N_6940,N_4279,N_3234);
nand U6941 (N_6941,N_4735,N_2637);
nand U6942 (N_6942,N_3687,N_4623);
nand U6943 (N_6943,N_3526,N_4602);
or U6944 (N_6944,N_4572,N_3425);
nor U6945 (N_6945,N_3105,N_2923);
or U6946 (N_6946,N_4000,N_4265);
or U6947 (N_6947,N_3603,N_3854);
nand U6948 (N_6948,N_4563,N_2531);
or U6949 (N_6949,N_3041,N_4761);
and U6950 (N_6950,N_4569,N_3839);
nand U6951 (N_6951,N_3264,N_3361);
xor U6952 (N_6952,N_4367,N_3465);
nor U6953 (N_6953,N_2502,N_3958);
nand U6954 (N_6954,N_3444,N_3849);
or U6955 (N_6955,N_4357,N_3754);
nand U6956 (N_6956,N_3899,N_3136);
nand U6957 (N_6957,N_2919,N_3590);
or U6958 (N_6958,N_2836,N_3068);
nor U6959 (N_6959,N_4096,N_2903);
nor U6960 (N_6960,N_4777,N_2886);
nor U6961 (N_6961,N_4664,N_3055);
or U6962 (N_6962,N_4136,N_3184);
nor U6963 (N_6963,N_3093,N_4845);
or U6964 (N_6964,N_3015,N_4791);
nor U6965 (N_6965,N_2809,N_4065);
nor U6966 (N_6966,N_3736,N_4127);
or U6967 (N_6967,N_3295,N_4907);
and U6968 (N_6968,N_3731,N_2995);
nand U6969 (N_6969,N_3672,N_3736);
and U6970 (N_6970,N_3939,N_4593);
or U6971 (N_6971,N_4756,N_3119);
nand U6972 (N_6972,N_4842,N_4201);
nand U6973 (N_6973,N_3830,N_4977);
or U6974 (N_6974,N_3656,N_3179);
or U6975 (N_6975,N_3022,N_2880);
nor U6976 (N_6976,N_4667,N_3925);
and U6977 (N_6977,N_3716,N_3875);
nand U6978 (N_6978,N_3550,N_3608);
nand U6979 (N_6979,N_4185,N_2503);
nor U6980 (N_6980,N_4578,N_3836);
nor U6981 (N_6981,N_4667,N_2839);
nor U6982 (N_6982,N_2509,N_3332);
nor U6983 (N_6983,N_2875,N_2742);
and U6984 (N_6984,N_2653,N_3758);
nand U6985 (N_6985,N_2880,N_2900);
nand U6986 (N_6986,N_3125,N_3074);
and U6987 (N_6987,N_4544,N_4769);
or U6988 (N_6988,N_4658,N_3540);
nor U6989 (N_6989,N_4814,N_2636);
nor U6990 (N_6990,N_3730,N_4516);
or U6991 (N_6991,N_4216,N_4336);
nand U6992 (N_6992,N_2727,N_2909);
nor U6993 (N_6993,N_2829,N_2577);
and U6994 (N_6994,N_2655,N_3280);
nand U6995 (N_6995,N_4113,N_2584);
nand U6996 (N_6996,N_4203,N_3706);
nand U6997 (N_6997,N_3816,N_3641);
nor U6998 (N_6998,N_4553,N_2901);
or U6999 (N_6999,N_3296,N_4138);
nor U7000 (N_7000,N_2520,N_3358);
nor U7001 (N_7001,N_4359,N_3553);
and U7002 (N_7002,N_4210,N_2536);
nand U7003 (N_7003,N_4653,N_4064);
or U7004 (N_7004,N_3436,N_2643);
or U7005 (N_7005,N_3763,N_4558);
or U7006 (N_7006,N_4364,N_4754);
nor U7007 (N_7007,N_2863,N_2689);
or U7008 (N_7008,N_4838,N_3851);
nand U7009 (N_7009,N_2993,N_4752);
and U7010 (N_7010,N_2658,N_2513);
nor U7011 (N_7011,N_2711,N_2570);
or U7012 (N_7012,N_4579,N_4332);
and U7013 (N_7013,N_3076,N_3938);
nor U7014 (N_7014,N_4577,N_3822);
nor U7015 (N_7015,N_2664,N_3390);
nor U7016 (N_7016,N_4486,N_3203);
xor U7017 (N_7017,N_4552,N_2828);
nand U7018 (N_7018,N_4648,N_4237);
nor U7019 (N_7019,N_3859,N_3456);
nor U7020 (N_7020,N_4087,N_3342);
nor U7021 (N_7021,N_4096,N_2651);
or U7022 (N_7022,N_4514,N_3030);
and U7023 (N_7023,N_4850,N_2637);
and U7024 (N_7024,N_4675,N_3057);
nor U7025 (N_7025,N_2987,N_4434);
nand U7026 (N_7026,N_4433,N_4246);
nand U7027 (N_7027,N_3561,N_4088);
nand U7028 (N_7028,N_2974,N_3520);
and U7029 (N_7029,N_4360,N_3112);
nand U7030 (N_7030,N_4154,N_4331);
nand U7031 (N_7031,N_4008,N_4100);
nor U7032 (N_7032,N_2614,N_3827);
or U7033 (N_7033,N_2847,N_4484);
and U7034 (N_7034,N_4196,N_2684);
nand U7035 (N_7035,N_4022,N_4323);
nor U7036 (N_7036,N_4410,N_3468);
nand U7037 (N_7037,N_4234,N_4323);
and U7038 (N_7038,N_4669,N_4333);
or U7039 (N_7039,N_3184,N_4205);
nand U7040 (N_7040,N_3003,N_3221);
nor U7041 (N_7041,N_3758,N_3379);
and U7042 (N_7042,N_4758,N_3100);
nor U7043 (N_7043,N_4617,N_4332);
nand U7044 (N_7044,N_3441,N_4996);
or U7045 (N_7045,N_4329,N_2740);
and U7046 (N_7046,N_4105,N_3180);
nor U7047 (N_7047,N_3350,N_3602);
nand U7048 (N_7048,N_4934,N_3884);
xnor U7049 (N_7049,N_4644,N_2540);
or U7050 (N_7050,N_4300,N_4851);
or U7051 (N_7051,N_4494,N_2859);
or U7052 (N_7052,N_3293,N_3195);
or U7053 (N_7053,N_3090,N_4341);
nand U7054 (N_7054,N_3649,N_2636);
or U7055 (N_7055,N_2502,N_4425);
or U7056 (N_7056,N_3014,N_4553);
or U7057 (N_7057,N_3034,N_4499);
and U7058 (N_7058,N_3763,N_3225);
nand U7059 (N_7059,N_4839,N_4166);
nand U7060 (N_7060,N_2989,N_2751);
or U7061 (N_7061,N_4348,N_2836);
nor U7062 (N_7062,N_4565,N_4080);
or U7063 (N_7063,N_4998,N_4382);
nor U7064 (N_7064,N_3241,N_3646);
and U7065 (N_7065,N_2794,N_2627);
nand U7066 (N_7066,N_3507,N_4245);
nand U7067 (N_7067,N_3003,N_3099);
and U7068 (N_7068,N_3352,N_3567);
or U7069 (N_7069,N_3890,N_4643);
and U7070 (N_7070,N_3668,N_2921);
or U7071 (N_7071,N_2653,N_3676);
or U7072 (N_7072,N_3167,N_4710);
nor U7073 (N_7073,N_4531,N_4194);
nand U7074 (N_7074,N_3556,N_3591);
nor U7075 (N_7075,N_3450,N_3006);
and U7076 (N_7076,N_2933,N_3775);
nor U7077 (N_7077,N_4102,N_4764);
nand U7078 (N_7078,N_3860,N_4770);
or U7079 (N_7079,N_3409,N_4060);
nor U7080 (N_7080,N_4075,N_4226);
nor U7081 (N_7081,N_3056,N_3264);
nand U7082 (N_7082,N_4908,N_4893);
and U7083 (N_7083,N_4268,N_3039);
nor U7084 (N_7084,N_3294,N_4944);
or U7085 (N_7085,N_3242,N_4323);
or U7086 (N_7086,N_3448,N_4377);
or U7087 (N_7087,N_4725,N_3772);
or U7088 (N_7088,N_3581,N_4849);
nor U7089 (N_7089,N_4284,N_4511);
and U7090 (N_7090,N_2905,N_3420);
nor U7091 (N_7091,N_3437,N_3703);
and U7092 (N_7092,N_3216,N_2700);
and U7093 (N_7093,N_4513,N_4882);
or U7094 (N_7094,N_4530,N_2522);
nor U7095 (N_7095,N_4479,N_3610);
nand U7096 (N_7096,N_4449,N_4458);
or U7097 (N_7097,N_2941,N_4439);
and U7098 (N_7098,N_3638,N_4415);
nor U7099 (N_7099,N_3204,N_2733);
or U7100 (N_7100,N_3164,N_4103);
nand U7101 (N_7101,N_3357,N_4109);
nand U7102 (N_7102,N_3380,N_2861);
or U7103 (N_7103,N_4157,N_2754);
xnor U7104 (N_7104,N_3424,N_3391);
nand U7105 (N_7105,N_2844,N_2573);
nand U7106 (N_7106,N_3400,N_4701);
nand U7107 (N_7107,N_3806,N_4958);
nand U7108 (N_7108,N_3759,N_3230);
nand U7109 (N_7109,N_3604,N_3640);
and U7110 (N_7110,N_4149,N_4946);
and U7111 (N_7111,N_2979,N_4668);
nor U7112 (N_7112,N_4186,N_3347);
nand U7113 (N_7113,N_3110,N_4701);
and U7114 (N_7114,N_4233,N_2538);
or U7115 (N_7115,N_3423,N_3978);
or U7116 (N_7116,N_2658,N_4380);
nor U7117 (N_7117,N_3918,N_2968);
nor U7118 (N_7118,N_3934,N_4260);
or U7119 (N_7119,N_4247,N_4265);
nor U7120 (N_7120,N_3510,N_4189);
or U7121 (N_7121,N_3869,N_2999);
nor U7122 (N_7122,N_2655,N_4543);
nand U7123 (N_7123,N_3885,N_4628);
nand U7124 (N_7124,N_3773,N_3206);
or U7125 (N_7125,N_4315,N_3214);
or U7126 (N_7126,N_3159,N_3050);
and U7127 (N_7127,N_2550,N_3413);
nand U7128 (N_7128,N_4443,N_3123);
or U7129 (N_7129,N_4900,N_3878);
or U7130 (N_7130,N_3219,N_4238);
nor U7131 (N_7131,N_3767,N_3704);
nand U7132 (N_7132,N_3768,N_3302);
nor U7133 (N_7133,N_2924,N_4136);
nand U7134 (N_7134,N_3730,N_4816);
nand U7135 (N_7135,N_3572,N_3502);
or U7136 (N_7136,N_4609,N_3354);
and U7137 (N_7137,N_2810,N_3833);
or U7138 (N_7138,N_3467,N_4884);
nand U7139 (N_7139,N_3779,N_4207);
or U7140 (N_7140,N_3402,N_4490);
and U7141 (N_7141,N_2834,N_4882);
and U7142 (N_7142,N_3343,N_3198);
nand U7143 (N_7143,N_4603,N_3339);
or U7144 (N_7144,N_3804,N_4876);
or U7145 (N_7145,N_4111,N_3359);
or U7146 (N_7146,N_4348,N_4638);
or U7147 (N_7147,N_4348,N_4720);
nand U7148 (N_7148,N_3663,N_4041);
and U7149 (N_7149,N_3228,N_2706);
nand U7150 (N_7150,N_3834,N_4039);
nor U7151 (N_7151,N_3382,N_3558);
nand U7152 (N_7152,N_4590,N_3557);
nor U7153 (N_7153,N_3120,N_2767);
nand U7154 (N_7154,N_4771,N_4405);
and U7155 (N_7155,N_4269,N_2765);
or U7156 (N_7156,N_3328,N_3546);
nor U7157 (N_7157,N_3856,N_2979);
nor U7158 (N_7158,N_3538,N_3133);
nor U7159 (N_7159,N_3258,N_4870);
or U7160 (N_7160,N_3592,N_3461);
and U7161 (N_7161,N_4365,N_2534);
nand U7162 (N_7162,N_3196,N_3961);
nor U7163 (N_7163,N_4292,N_3293);
or U7164 (N_7164,N_3253,N_4292);
nor U7165 (N_7165,N_2667,N_2754);
nand U7166 (N_7166,N_2869,N_4935);
or U7167 (N_7167,N_4530,N_4345);
nor U7168 (N_7168,N_2750,N_3629);
nor U7169 (N_7169,N_4390,N_4349);
nor U7170 (N_7170,N_4842,N_4893);
or U7171 (N_7171,N_4054,N_3774);
nand U7172 (N_7172,N_4298,N_2636);
nor U7173 (N_7173,N_4516,N_3098);
nand U7174 (N_7174,N_2696,N_3764);
nor U7175 (N_7175,N_3472,N_2572);
or U7176 (N_7176,N_4736,N_3861);
nor U7177 (N_7177,N_4907,N_4998);
and U7178 (N_7178,N_3843,N_3465);
nor U7179 (N_7179,N_2705,N_3411);
nand U7180 (N_7180,N_3937,N_4561);
nor U7181 (N_7181,N_4619,N_2732);
nand U7182 (N_7182,N_4681,N_4223);
and U7183 (N_7183,N_4775,N_4782);
and U7184 (N_7184,N_3319,N_3380);
nor U7185 (N_7185,N_3266,N_3419);
nor U7186 (N_7186,N_3002,N_3586);
and U7187 (N_7187,N_4857,N_3121);
and U7188 (N_7188,N_2589,N_3735);
xor U7189 (N_7189,N_4360,N_4647);
nor U7190 (N_7190,N_2771,N_2596);
nand U7191 (N_7191,N_3726,N_3705);
nand U7192 (N_7192,N_4265,N_3809);
nor U7193 (N_7193,N_4892,N_4968);
nor U7194 (N_7194,N_4376,N_4590);
nand U7195 (N_7195,N_4500,N_2904);
or U7196 (N_7196,N_3735,N_3646);
or U7197 (N_7197,N_3064,N_4707);
nor U7198 (N_7198,N_2874,N_4187);
or U7199 (N_7199,N_4983,N_3635);
nand U7200 (N_7200,N_2624,N_4613);
nor U7201 (N_7201,N_4730,N_4270);
and U7202 (N_7202,N_4902,N_4669);
and U7203 (N_7203,N_3618,N_3087);
nor U7204 (N_7204,N_2548,N_3503);
nand U7205 (N_7205,N_4486,N_4922);
xor U7206 (N_7206,N_3432,N_3220);
nor U7207 (N_7207,N_2740,N_3807);
nor U7208 (N_7208,N_4886,N_2639);
nand U7209 (N_7209,N_3642,N_4037);
nor U7210 (N_7210,N_4651,N_3463);
or U7211 (N_7211,N_4036,N_2627);
and U7212 (N_7212,N_4860,N_3709);
nor U7213 (N_7213,N_4186,N_3722);
and U7214 (N_7214,N_3774,N_4201);
nor U7215 (N_7215,N_2643,N_3558);
and U7216 (N_7216,N_4443,N_3963);
and U7217 (N_7217,N_4831,N_4371);
or U7218 (N_7218,N_4749,N_3559);
nand U7219 (N_7219,N_2602,N_4745);
and U7220 (N_7220,N_3270,N_2812);
nor U7221 (N_7221,N_4199,N_3616);
and U7222 (N_7222,N_4668,N_4191);
nand U7223 (N_7223,N_4184,N_2702);
or U7224 (N_7224,N_4316,N_3796);
or U7225 (N_7225,N_4467,N_2899);
nor U7226 (N_7226,N_3935,N_2628);
and U7227 (N_7227,N_4787,N_4187);
nand U7228 (N_7228,N_4939,N_4054);
or U7229 (N_7229,N_3346,N_2673);
or U7230 (N_7230,N_4906,N_4949);
nor U7231 (N_7231,N_3127,N_4808);
nand U7232 (N_7232,N_3839,N_4033);
or U7233 (N_7233,N_4084,N_2798);
nor U7234 (N_7234,N_2648,N_4368);
nand U7235 (N_7235,N_3178,N_4718);
nor U7236 (N_7236,N_2734,N_4062);
nor U7237 (N_7237,N_2596,N_3243);
nor U7238 (N_7238,N_3296,N_4946);
or U7239 (N_7239,N_3051,N_4536);
or U7240 (N_7240,N_3520,N_3758);
nor U7241 (N_7241,N_4393,N_4076);
nor U7242 (N_7242,N_3773,N_2972);
or U7243 (N_7243,N_4857,N_4435);
or U7244 (N_7244,N_3693,N_3989);
or U7245 (N_7245,N_3297,N_3795);
or U7246 (N_7246,N_4808,N_3004);
nand U7247 (N_7247,N_3206,N_4523);
or U7248 (N_7248,N_2721,N_4415);
and U7249 (N_7249,N_2729,N_4010);
nand U7250 (N_7250,N_3137,N_4820);
or U7251 (N_7251,N_3404,N_4945);
and U7252 (N_7252,N_4890,N_2660);
and U7253 (N_7253,N_2853,N_2975);
nand U7254 (N_7254,N_3085,N_4318);
and U7255 (N_7255,N_3732,N_4888);
nor U7256 (N_7256,N_3531,N_3046);
xnor U7257 (N_7257,N_4198,N_3533);
nand U7258 (N_7258,N_4715,N_3880);
or U7259 (N_7259,N_3389,N_2980);
or U7260 (N_7260,N_4588,N_3451);
and U7261 (N_7261,N_3722,N_3314);
nand U7262 (N_7262,N_3986,N_4657);
and U7263 (N_7263,N_3746,N_3302);
and U7264 (N_7264,N_2923,N_3293);
nor U7265 (N_7265,N_4422,N_2920);
and U7266 (N_7266,N_3053,N_3911);
nand U7267 (N_7267,N_2899,N_2950);
nand U7268 (N_7268,N_3242,N_2550);
nor U7269 (N_7269,N_4063,N_3240);
nor U7270 (N_7270,N_3581,N_4090);
nor U7271 (N_7271,N_3709,N_4445);
and U7272 (N_7272,N_3621,N_3216);
or U7273 (N_7273,N_4201,N_3681);
nor U7274 (N_7274,N_3812,N_3814);
nor U7275 (N_7275,N_4630,N_4866);
nand U7276 (N_7276,N_4093,N_3141);
nor U7277 (N_7277,N_4562,N_4843);
nand U7278 (N_7278,N_2962,N_3941);
and U7279 (N_7279,N_3812,N_2567);
nor U7280 (N_7280,N_3347,N_3734);
nand U7281 (N_7281,N_2789,N_4056);
nand U7282 (N_7282,N_4887,N_3050);
nand U7283 (N_7283,N_4805,N_4271);
nand U7284 (N_7284,N_2659,N_4610);
or U7285 (N_7285,N_3611,N_4313);
nor U7286 (N_7286,N_3569,N_4995);
nand U7287 (N_7287,N_4730,N_2755);
or U7288 (N_7288,N_3360,N_3587);
and U7289 (N_7289,N_3876,N_3560);
nor U7290 (N_7290,N_2935,N_4136);
or U7291 (N_7291,N_3468,N_2688);
or U7292 (N_7292,N_3038,N_4706);
nor U7293 (N_7293,N_2651,N_3991);
or U7294 (N_7294,N_2719,N_4265);
nor U7295 (N_7295,N_4209,N_3812);
and U7296 (N_7296,N_3791,N_3488);
nor U7297 (N_7297,N_4838,N_4085);
nand U7298 (N_7298,N_2797,N_3612);
nand U7299 (N_7299,N_2957,N_3085);
nand U7300 (N_7300,N_2759,N_4697);
nand U7301 (N_7301,N_3415,N_3859);
or U7302 (N_7302,N_3992,N_3043);
and U7303 (N_7303,N_3589,N_3704);
nor U7304 (N_7304,N_3381,N_4917);
and U7305 (N_7305,N_3777,N_2609);
or U7306 (N_7306,N_4367,N_4931);
or U7307 (N_7307,N_4400,N_3377);
nor U7308 (N_7308,N_3883,N_3191);
nor U7309 (N_7309,N_2947,N_4462);
nor U7310 (N_7310,N_2855,N_4985);
nand U7311 (N_7311,N_2630,N_4396);
nand U7312 (N_7312,N_2946,N_3705);
or U7313 (N_7313,N_3119,N_4280);
or U7314 (N_7314,N_3044,N_3979);
nand U7315 (N_7315,N_4809,N_4106);
nor U7316 (N_7316,N_3175,N_4825);
xor U7317 (N_7317,N_4826,N_3879);
nand U7318 (N_7318,N_4596,N_4740);
nand U7319 (N_7319,N_3003,N_4407);
or U7320 (N_7320,N_3749,N_4978);
and U7321 (N_7321,N_4902,N_3256);
nand U7322 (N_7322,N_3900,N_4568);
or U7323 (N_7323,N_3929,N_3785);
and U7324 (N_7324,N_4939,N_4353);
nor U7325 (N_7325,N_3851,N_3171);
nor U7326 (N_7326,N_3295,N_4489);
nand U7327 (N_7327,N_2717,N_4727);
nor U7328 (N_7328,N_4201,N_3295);
nor U7329 (N_7329,N_4010,N_3824);
nor U7330 (N_7330,N_4190,N_3744);
nor U7331 (N_7331,N_3841,N_2717);
or U7332 (N_7332,N_4436,N_2941);
and U7333 (N_7333,N_3746,N_3883);
nand U7334 (N_7334,N_3067,N_4957);
and U7335 (N_7335,N_2628,N_2751);
nor U7336 (N_7336,N_3577,N_2872);
nand U7337 (N_7337,N_3409,N_4271);
and U7338 (N_7338,N_3093,N_3800);
or U7339 (N_7339,N_3842,N_4374);
nor U7340 (N_7340,N_3886,N_2651);
nand U7341 (N_7341,N_4264,N_3332);
nand U7342 (N_7342,N_4285,N_3793);
nand U7343 (N_7343,N_4716,N_2745);
or U7344 (N_7344,N_3607,N_2798);
nor U7345 (N_7345,N_2971,N_3692);
and U7346 (N_7346,N_3265,N_4033);
nand U7347 (N_7347,N_4112,N_4640);
or U7348 (N_7348,N_4274,N_2940);
and U7349 (N_7349,N_4194,N_2697);
and U7350 (N_7350,N_3824,N_2949);
and U7351 (N_7351,N_3142,N_4044);
nor U7352 (N_7352,N_3643,N_3071);
nor U7353 (N_7353,N_4308,N_2831);
or U7354 (N_7354,N_4162,N_4228);
and U7355 (N_7355,N_3523,N_3257);
nor U7356 (N_7356,N_4877,N_2886);
nor U7357 (N_7357,N_4982,N_3587);
and U7358 (N_7358,N_3390,N_3220);
or U7359 (N_7359,N_4777,N_3959);
and U7360 (N_7360,N_4671,N_3980);
nand U7361 (N_7361,N_2582,N_2760);
or U7362 (N_7362,N_2866,N_4379);
nand U7363 (N_7363,N_3594,N_4062);
nor U7364 (N_7364,N_3772,N_4342);
and U7365 (N_7365,N_3338,N_4605);
and U7366 (N_7366,N_4588,N_2725);
and U7367 (N_7367,N_3528,N_3448);
and U7368 (N_7368,N_2535,N_4787);
nor U7369 (N_7369,N_4670,N_4244);
nand U7370 (N_7370,N_4844,N_2654);
nand U7371 (N_7371,N_4318,N_2923);
and U7372 (N_7372,N_4309,N_3547);
nor U7373 (N_7373,N_3748,N_2595);
nor U7374 (N_7374,N_2585,N_3987);
and U7375 (N_7375,N_2528,N_4699);
or U7376 (N_7376,N_3220,N_4675);
nand U7377 (N_7377,N_4511,N_3638);
nand U7378 (N_7378,N_3600,N_3468);
nand U7379 (N_7379,N_4125,N_3302);
nor U7380 (N_7380,N_3077,N_3286);
nand U7381 (N_7381,N_3583,N_4456);
and U7382 (N_7382,N_3430,N_3611);
nand U7383 (N_7383,N_3088,N_3703);
nor U7384 (N_7384,N_4671,N_4528);
or U7385 (N_7385,N_2603,N_3857);
or U7386 (N_7386,N_4225,N_2500);
and U7387 (N_7387,N_2734,N_3358);
nand U7388 (N_7388,N_3831,N_3134);
and U7389 (N_7389,N_3855,N_3614);
nand U7390 (N_7390,N_3640,N_4851);
or U7391 (N_7391,N_3597,N_4141);
or U7392 (N_7392,N_3883,N_4240);
nand U7393 (N_7393,N_4070,N_3582);
nand U7394 (N_7394,N_4183,N_3615);
and U7395 (N_7395,N_4214,N_4855);
or U7396 (N_7396,N_4841,N_4992);
nor U7397 (N_7397,N_2825,N_4377);
nand U7398 (N_7398,N_3672,N_4456);
nor U7399 (N_7399,N_4009,N_2761);
and U7400 (N_7400,N_2578,N_4644);
and U7401 (N_7401,N_3404,N_2941);
nor U7402 (N_7402,N_4131,N_4528);
or U7403 (N_7403,N_2892,N_4174);
nand U7404 (N_7404,N_4103,N_2889);
nor U7405 (N_7405,N_2519,N_3444);
nand U7406 (N_7406,N_2731,N_2842);
nand U7407 (N_7407,N_3864,N_4525);
or U7408 (N_7408,N_2899,N_3897);
nand U7409 (N_7409,N_4360,N_4082);
and U7410 (N_7410,N_4284,N_4543);
nor U7411 (N_7411,N_3484,N_4931);
nor U7412 (N_7412,N_3933,N_2694);
nand U7413 (N_7413,N_3478,N_3913);
and U7414 (N_7414,N_2509,N_2644);
and U7415 (N_7415,N_3444,N_4635);
and U7416 (N_7416,N_4409,N_3111);
nor U7417 (N_7417,N_3624,N_4768);
nand U7418 (N_7418,N_4457,N_2617);
nor U7419 (N_7419,N_4058,N_2555);
or U7420 (N_7420,N_4877,N_3505);
nand U7421 (N_7421,N_3077,N_4753);
xor U7422 (N_7422,N_4871,N_2715);
or U7423 (N_7423,N_4883,N_4324);
nand U7424 (N_7424,N_2626,N_4641);
nor U7425 (N_7425,N_3443,N_4586);
and U7426 (N_7426,N_4288,N_4468);
nand U7427 (N_7427,N_4718,N_3423);
nor U7428 (N_7428,N_2992,N_3964);
and U7429 (N_7429,N_4876,N_4699);
nor U7430 (N_7430,N_3193,N_4195);
nor U7431 (N_7431,N_3922,N_3263);
nor U7432 (N_7432,N_3474,N_3921);
and U7433 (N_7433,N_2511,N_3387);
and U7434 (N_7434,N_4966,N_3813);
or U7435 (N_7435,N_3169,N_4254);
nand U7436 (N_7436,N_4114,N_3959);
and U7437 (N_7437,N_2983,N_3405);
and U7438 (N_7438,N_3225,N_3570);
and U7439 (N_7439,N_3810,N_3784);
nand U7440 (N_7440,N_2820,N_4618);
or U7441 (N_7441,N_3853,N_3855);
or U7442 (N_7442,N_2677,N_3446);
or U7443 (N_7443,N_4678,N_4424);
xor U7444 (N_7444,N_2728,N_4005);
nor U7445 (N_7445,N_2513,N_3218);
nor U7446 (N_7446,N_2675,N_2910);
and U7447 (N_7447,N_2928,N_4684);
nand U7448 (N_7448,N_4973,N_3329);
or U7449 (N_7449,N_2932,N_2706);
and U7450 (N_7450,N_3465,N_3889);
nand U7451 (N_7451,N_3074,N_3738);
nand U7452 (N_7452,N_3004,N_4144);
and U7453 (N_7453,N_2707,N_2869);
and U7454 (N_7454,N_3853,N_4508);
nand U7455 (N_7455,N_2999,N_4533);
or U7456 (N_7456,N_2697,N_4518);
nand U7457 (N_7457,N_3499,N_2562);
nor U7458 (N_7458,N_2720,N_3292);
nor U7459 (N_7459,N_3216,N_4312);
nand U7460 (N_7460,N_3270,N_3129);
nor U7461 (N_7461,N_4723,N_4972);
nor U7462 (N_7462,N_3491,N_3808);
nand U7463 (N_7463,N_2623,N_4380);
nor U7464 (N_7464,N_4156,N_2699);
nor U7465 (N_7465,N_4787,N_2976);
or U7466 (N_7466,N_3388,N_2895);
nor U7467 (N_7467,N_2673,N_3639);
and U7468 (N_7468,N_3279,N_4877);
and U7469 (N_7469,N_4607,N_3266);
nor U7470 (N_7470,N_4320,N_4639);
nand U7471 (N_7471,N_4718,N_4709);
or U7472 (N_7472,N_4205,N_3723);
nand U7473 (N_7473,N_2561,N_3050);
and U7474 (N_7474,N_3367,N_3985);
nand U7475 (N_7475,N_4719,N_4987);
nor U7476 (N_7476,N_2942,N_4004);
nor U7477 (N_7477,N_2537,N_3104);
or U7478 (N_7478,N_4545,N_3126);
nand U7479 (N_7479,N_3489,N_4366);
or U7480 (N_7480,N_4171,N_4478);
or U7481 (N_7481,N_4398,N_4381);
or U7482 (N_7482,N_3920,N_4538);
and U7483 (N_7483,N_4854,N_3257);
nor U7484 (N_7484,N_3883,N_4047);
nor U7485 (N_7485,N_3663,N_4672);
or U7486 (N_7486,N_3524,N_3711);
nand U7487 (N_7487,N_4372,N_2681);
nand U7488 (N_7488,N_4779,N_3122);
nand U7489 (N_7489,N_2979,N_4855);
and U7490 (N_7490,N_2678,N_2807);
and U7491 (N_7491,N_4715,N_4346);
or U7492 (N_7492,N_3879,N_2885);
nand U7493 (N_7493,N_3673,N_3417);
or U7494 (N_7494,N_3564,N_2750);
or U7495 (N_7495,N_3279,N_3267);
nor U7496 (N_7496,N_3764,N_4660);
and U7497 (N_7497,N_4150,N_4424);
nand U7498 (N_7498,N_4601,N_4387);
xnor U7499 (N_7499,N_4271,N_3904);
or U7500 (N_7500,N_6048,N_7012);
nand U7501 (N_7501,N_5102,N_5658);
nand U7502 (N_7502,N_5744,N_5407);
and U7503 (N_7503,N_7194,N_5435);
and U7504 (N_7504,N_5157,N_6888);
nand U7505 (N_7505,N_7297,N_5362);
and U7506 (N_7506,N_5560,N_6553);
or U7507 (N_7507,N_5418,N_5936);
nor U7508 (N_7508,N_6793,N_6255);
nor U7509 (N_7509,N_7287,N_5307);
nor U7510 (N_7510,N_7461,N_6096);
nand U7511 (N_7511,N_6786,N_6966);
nor U7512 (N_7512,N_5574,N_7002);
nand U7513 (N_7513,N_5991,N_5176);
nand U7514 (N_7514,N_7064,N_5737);
nor U7515 (N_7515,N_5538,N_6527);
or U7516 (N_7516,N_7184,N_6879);
and U7517 (N_7517,N_6004,N_5276);
and U7518 (N_7518,N_6635,N_6331);
nor U7519 (N_7519,N_5400,N_5845);
nand U7520 (N_7520,N_5838,N_5814);
or U7521 (N_7521,N_5897,N_5172);
and U7522 (N_7522,N_6273,N_5243);
nand U7523 (N_7523,N_6083,N_6479);
and U7524 (N_7524,N_5969,N_5074);
nand U7525 (N_7525,N_5644,N_7120);
nor U7526 (N_7526,N_6902,N_5395);
nor U7527 (N_7527,N_6768,N_7102);
nor U7528 (N_7528,N_5662,N_5588);
nand U7529 (N_7529,N_5776,N_5431);
nand U7530 (N_7530,N_5651,N_5563);
and U7531 (N_7531,N_6026,N_5391);
or U7532 (N_7532,N_6107,N_5187);
or U7533 (N_7533,N_7425,N_5620);
and U7534 (N_7534,N_5487,N_5808);
nand U7535 (N_7535,N_5014,N_6093);
nand U7536 (N_7536,N_6311,N_5708);
and U7537 (N_7537,N_5840,N_6952);
nor U7538 (N_7538,N_5943,N_5528);
nand U7539 (N_7539,N_6817,N_6954);
and U7540 (N_7540,N_7027,N_5861);
and U7541 (N_7541,N_6000,N_5165);
or U7542 (N_7542,N_6856,N_5634);
and U7543 (N_7543,N_5210,N_5993);
or U7544 (N_7544,N_6468,N_6665);
or U7545 (N_7545,N_6304,N_5095);
nand U7546 (N_7546,N_5041,N_5606);
or U7547 (N_7547,N_5581,N_6851);
nor U7548 (N_7548,N_6429,N_6741);
and U7549 (N_7549,N_5515,N_7398);
and U7550 (N_7550,N_7079,N_7411);
nor U7551 (N_7551,N_5971,N_6079);
or U7552 (N_7552,N_6764,N_6327);
nor U7553 (N_7553,N_6217,N_6341);
nor U7554 (N_7554,N_6846,N_6784);
or U7555 (N_7555,N_7443,N_5793);
or U7556 (N_7556,N_7445,N_5850);
or U7557 (N_7557,N_6470,N_6416);
nor U7558 (N_7558,N_7291,N_5393);
and U7559 (N_7559,N_5447,N_5485);
nor U7560 (N_7560,N_5050,N_5541);
and U7561 (N_7561,N_5119,N_7199);
or U7562 (N_7562,N_5822,N_5690);
and U7563 (N_7563,N_7213,N_6742);
or U7564 (N_7564,N_5779,N_5898);
and U7565 (N_7565,N_6514,N_6729);
nand U7566 (N_7566,N_5137,N_5445);
nand U7567 (N_7567,N_6143,N_6707);
and U7568 (N_7568,N_6644,N_6338);
nand U7569 (N_7569,N_5423,N_6020);
nor U7570 (N_7570,N_6296,N_5605);
and U7571 (N_7571,N_5408,N_7065);
nand U7572 (N_7572,N_5373,N_7178);
nor U7573 (N_7573,N_5016,N_5412);
nand U7574 (N_7574,N_6188,N_5295);
or U7575 (N_7575,N_7166,N_5381);
or U7576 (N_7576,N_6750,N_5275);
and U7577 (N_7577,N_5592,N_7243);
nand U7578 (N_7578,N_6886,N_6989);
and U7579 (N_7579,N_7438,N_7327);
nand U7580 (N_7580,N_6818,N_5156);
or U7581 (N_7581,N_6447,N_5181);
and U7582 (N_7582,N_6908,N_5555);
or U7583 (N_7583,N_6552,N_6946);
nor U7584 (N_7584,N_5013,N_5313);
nor U7585 (N_7585,N_7201,N_7402);
or U7586 (N_7586,N_6618,N_6100);
and U7587 (N_7587,N_5584,N_5207);
nand U7588 (N_7588,N_7433,N_6874);
and U7589 (N_7589,N_6598,N_7227);
nand U7590 (N_7590,N_5748,N_6628);
nand U7591 (N_7591,N_5753,N_5451);
or U7592 (N_7592,N_7476,N_5027);
nand U7593 (N_7593,N_7003,N_6633);
nand U7594 (N_7594,N_6207,N_7488);
nor U7595 (N_7595,N_6686,N_5490);
or U7596 (N_7596,N_5614,N_7190);
xor U7597 (N_7597,N_6382,N_5399);
or U7598 (N_7598,N_6190,N_7099);
nor U7599 (N_7599,N_6920,N_6463);
nor U7600 (N_7600,N_7109,N_5472);
nor U7601 (N_7601,N_6254,N_6008);
and U7602 (N_7602,N_6828,N_6054);
xnor U7603 (N_7603,N_5323,N_6816);
nor U7604 (N_7604,N_7377,N_5937);
and U7605 (N_7605,N_5880,N_5402);
nor U7606 (N_7606,N_5926,N_5632);
nand U7607 (N_7607,N_6277,N_6513);
nand U7608 (N_7608,N_7464,N_5561);
nor U7609 (N_7609,N_6825,N_6007);
nor U7610 (N_7610,N_5450,N_5772);
and U7611 (N_7611,N_6924,N_5785);
and U7612 (N_7612,N_7192,N_5653);
nand U7613 (N_7613,N_6839,N_5828);
and U7614 (N_7614,N_5031,N_5734);
or U7615 (N_7615,N_5401,N_6643);
nor U7616 (N_7616,N_7395,N_5815);
nor U7617 (N_7617,N_5092,N_6047);
xnor U7618 (N_7618,N_5234,N_6791);
nor U7619 (N_7619,N_7352,N_6883);
and U7620 (N_7620,N_5083,N_6948);
and U7621 (N_7621,N_6744,N_7479);
nand U7622 (N_7622,N_7207,N_7378);
or U7623 (N_7623,N_5512,N_5694);
nor U7624 (N_7624,N_5405,N_5446);
and U7625 (N_7625,N_5069,N_6101);
nand U7626 (N_7626,N_7058,N_6522);
and U7627 (N_7627,N_6295,N_5202);
or U7628 (N_7628,N_5842,N_6415);
nand U7629 (N_7629,N_5059,N_6484);
nand U7630 (N_7630,N_6657,N_5624);
nand U7631 (N_7631,N_7333,N_5701);
nand U7632 (N_7632,N_6350,N_7100);
nor U7633 (N_7633,N_5433,N_5497);
nand U7634 (N_7634,N_6528,N_6547);
nand U7635 (N_7635,N_5827,N_5676);
nand U7636 (N_7636,N_6170,N_7034);
nor U7637 (N_7637,N_6861,N_5343);
and U7638 (N_7638,N_5328,N_6570);
and U7639 (N_7639,N_5826,N_7257);
nand U7640 (N_7640,N_6291,N_7339);
and U7641 (N_7641,N_6352,N_5292);
nor U7642 (N_7642,N_6494,N_6044);
nand U7643 (N_7643,N_5319,N_5854);
nand U7644 (N_7644,N_5832,N_7359);
or U7645 (N_7645,N_7215,N_6746);
and U7646 (N_7646,N_5000,N_6132);
nand U7647 (N_7647,N_5824,N_5650);
and U7648 (N_7648,N_6042,N_5612);
or U7649 (N_7649,N_6560,N_7161);
nor U7650 (N_7650,N_7165,N_5018);
and U7651 (N_7651,N_6660,N_5720);
and U7652 (N_7652,N_5930,N_7038);
or U7653 (N_7653,N_5914,N_6235);
nand U7654 (N_7654,N_6421,N_7442);
nand U7655 (N_7655,N_6252,N_6388);
nor U7656 (N_7656,N_5968,N_5966);
and U7657 (N_7657,N_5342,N_6670);
or U7658 (N_7658,N_7258,N_7299);
nand U7659 (N_7659,N_5962,N_6664);
or U7660 (N_7660,N_5033,N_5678);
nor U7661 (N_7661,N_7407,N_5590);
or U7662 (N_7662,N_7022,N_6781);
or U7663 (N_7663,N_5061,N_5378);
and U7664 (N_7664,N_5766,N_6442);
nor U7665 (N_7665,N_6226,N_5194);
or U7666 (N_7666,N_5078,N_5049);
or U7667 (N_7667,N_6033,N_5552);
or U7668 (N_7668,N_6676,N_5046);
or U7669 (N_7669,N_7073,N_6929);
nor U7670 (N_7670,N_5934,N_5261);
nor U7671 (N_7671,N_5454,N_5311);
and U7672 (N_7672,N_5422,N_5645);
and U7673 (N_7673,N_6540,N_6530);
nand U7674 (N_7674,N_6059,N_5274);
nor U7675 (N_7675,N_5992,N_6790);
nand U7676 (N_7676,N_6474,N_5289);
nand U7677 (N_7677,N_6538,N_5834);
and U7678 (N_7678,N_7310,N_7366);
or U7679 (N_7679,N_6003,N_5995);
or U7680 (N_7680,N_7233,N_6408);
nand U7681 (N_7681,N_7264,N_6144);
nor U7682 (N_7682,N_5548,N_7342);
nand U7683 (N_7683,N_7228,N_6844);
or U7684 (N_7684,N_6994,N_5988);
nand U7685 (N_7685,N_6820,N_7152);
or U7686 (N_7686,N_6916,N_6848);
or U7687 (N_7687,N_5558,N_5038);
and U7688 (N_7688,N_5750,N_7029);
nand U7689 (N_7689,N_5367,N_5794);
or U7690 (N_7690,N_6890,N_6605);
and U7691 (N_7691,N_6455,N_5689);
nor U7692 (N_7692,N_5478,N_7195);
nor U7693 (N_7693,N_5536,N_5216);
nor U7694 (N_7694,N_6775,N_6885);
nand U7695 (N_7695,N_5121,N_6477);
or U7696 (N_7696,N_5388,N_7451);
nand U7697 (N_7697,N_5514,N_6977);
nand U7698 (N_7698,N_7295,N_7103);
nand U7699 (N_7699,N_7094,N_5191);
and U7700 (N_7700,N_5819,N_7119);
nand U7701 (N_7701,N_6165,N_6765);
and U7702 (N_7702,N_7343,N_5666);
and U7703 (N_7703,N_5652,N_6968);
nor U7704 (N_7704,N_6336,N_5831);
or U7705 (N_7705,N_6580,N_6070);
nor U7706 (N_7706,N_7289,N_6257);
or U7707 (N_7707,N_7429,N_5231);
or U7708 (N_7708,N_6533,N_7322);
nor U7709 (N_7709,N_5709,N_5304);
or U7710 (N_7710,N_5603,N_6053);
nor U7711 (N_7711,N_5477,N_6519);
or U7712 (N_7712,N_7332,N_6131);
nor U7713 (N_7713,N_5359,N_7140);
and U7714 (N_7714,N_5707,N_6164);
and U7715 (N_7715,N_6064,N_6082);
nand U7716 (N_7716,N_5628,N_7096);
and U7717 (N_7717,N_7414,N_6094);
nand U7718 (N_7718,N_5580,N_5519);
nand U7719 (N_7719,N_6616,N_6127);
or U7720 (N_7720,N_6162,N_7121);
or U7721 (N_7721,N_6115,N_5120);
or U7722 (N_7722,N_6783,N_7284);
and U7723 (N_7723,N_7173,N_6403);
nand U7724 (N_7724,N_6495,N_7259);
or U7725 (N_7725,N_6205,N_6762);
and U7726 (N_7726,N_6667,N_6544);
nand U7727 (N_7727,N_7468,N_6089);
nor U7728 (N_7728,N_5017,N_5111);
nor U7729 (N_7729,N_6011,N_7315);
nor U7730 (N_7730,N_5566,N_5736);
or U7731 (N_7731,N_7293,N_6090);
nor U7732 (N_7732,N_6505,N_7338);
and U7733 (N_7733,N_6045,N_6326);
or U7734 (N_7734,N_5532,N_7495);
and U7735 (N_7735,N_6542,N_5055);
nor U7736 (N_7736,N_5812,N_5193);
nor U7737 (N_7737,N_6088,N_6725);
nand U7738 (N_7738,N_7350,N_7057);
nor U7739 (N_7739,N_5250,N_5019);
nor U7740 (N_7740,N_7018,N_5467);
or U7741 (N_7741,N_5476,N_5201);
nand U7742 (N_7742,N_6689,N_7313);
nand U7743 (N_7743,N_6923,N_7145);
nor U7744 (N_7744,N_5264,N_6963);
or U7745 (N_7745,N_7242,N_6136);
and U7746 (N_7746,N_6747,N_5646);
nor U7747 (N_7747,N_5168,N_6991);
nand U7748 (N_7748,N_7128,N_7281);
nor U7749 (N_7749,N_6401,N_5981);
and U7750 (N_7750,N_5414,N_6347);
nor U7751 (N_7751,N_6197,N_7000);
and U7752 (N_7752,N_6978,N_5260);
or U7753 (N_7753,N_6102,N_5475);
nand U7754 (N_7754,N_6106,N_6850);
or U7755 (N_7755,N_6843,N_5064);
and U7756 (N_7756,N_5858,N_5718);
nand U7757 (N_7757,N_6371,N_6752);
nand U7758 (N_7758,N_5463,N_7255);
or U7759 (N_7759,N_5335,N_6773);
or U7760 (N_7760,N_7172,N_7361);
nand U7761 (N_7761,N_5244,N_5852);
and U7762 (N_7762,N_5329,N_6551);
or U7763 (N_7763,N_5573,N_5839);
nor U7764 (N_7764,N_7372,N_6831);
nor U7765 (N_7765,N_6085,N_7216);
nand U7766 (N_7766,N_7142,N_6334);
nand U7767 (N_7767,N_7188,N_6889);
nand U7768 (N_7768,N_6105,N_5654);
nand U7769 (N_7769,N_6456,N_7447);
nand U7770 (N_7770,N_6322,N_6492);
and U7771 (N_7771,N_7204,N_5496);
nor U7772 (N_7772,N_7460,N_7063);
or U7773 (N_7773,N_7308,N_5615);
or U7774 (N_7774,N_5188,N_5642);
nand U7775 (N_7775,N_5398,N_6469);
nand U7776 (N_7776,N_7336,N_5686);
nor U7777 (N_7777,N_5209,N_7469);
or U7778 (N_7778,N_5136,N_5687);
and U7779 (N_7779,N_5762,N_5722);
nor U7780 (N_7780,N_5340,N_6737);
and U7781 (N_7781,N_7251,N_6405);
and U7782 (N_7782,N_6056,N_5942);
or U7783 (N_7783,N_5390,N_6880);
or U7784 (N_7784,N_6575,N_5910);
and U7785 (N_7785,N_5586,N_7351);
nand U7786 (N_7786,N_6976,N_6596);
nand U7787 (N_7787,N_7225,N_6537);
or U7788 (N_7788,N_5290,N_6699);
or U7789 (N_7789,N_5228,N_7101);
nor U7790 (N_7790,N_6718,N_7397);
or U7791 (N_7791,N_5413,N_6811);
nor U7792 (N_7792,N_7205,N_6599);
and U7793 (N_7793,N_7435,N_6263);
nor U7794 (N_7794,N_5011,N_5738);
nor U7795 (N_7795,N_5145,N_5219);
or U7796 (N_7796,N_7450,N_6005);
and U7797 (N_7797,N_6055,N_6753);
nand U7798 (N_7798,N_7448,N_5551);
nor U7799 (N_7799,N_5818,N_6185);
nor U7800 (N_7800,N_6545,N_7486);
or U7801 (N_7801,N_6182,N_6898);
nand U7802 (N_7802,N_5980,N_6803);
nand U7803 (N_7803,N_7422,N_6283);
nor U7804 (N_7804,N_5263,N_5425);
or U7805 (N_7805,N_5530,N_5987);
nor U7806 (N_7806,N_6970,N_6041);
nor U7807 (N_7807,N_7106,N_6097);
nand U7808 (N_7808,N_5203,N_5746);
nor U7809 (N_7809,N_6668,N_6719);
nand U7810 (N_7810,N_5177,N_7390);
nor U7811 (N_7811,N_7421,N_6275);
or U7812 (N_7812,N_5949,N_5090);
or U7813 (N_7813,N_6732,N_6853);
nor U7814 (N_7814,N_6662,N_6965);
nor U7815 (N_7815,N_5480,N_5301);
or U7816 (N_7816,N_5318,N_7298);
and U7817 (N_7817,N_6335,N_6493);
or U7818 (N_7818,N_6800,N_7371);
and U7819 (N_7819,N_6496,N_7091);
or U7820 (N_7820,N_6915,N_7381);
nand U7821 (N_7821,N_5035,N_6919);
nand U7822 (N_7822,N_6148,N_7485);
nand U7823 (N_7823,N_7380,N_6754);
and U7824 (N_7824,N_6647,N_7382);
or U7825 (N_7825,N_5449,N_6308);
or U7826 (N_7826,N_6434,N_5513);
and U7827 (N_7827,N_5043,N_5577);
or U7828 (N_7828,N_6807,N_5696);
nand U7829 (N_7829,N_5556,N_5841);
nor U7830 (N_7830,N_5559,N_7236);
or U7831 (N_7831,N_7023,N_6031);
and U7832 (N_7832,N_5887,N_5797);
nand U7833 (N_7833,N_7368,N_5075);
nand U7834 (N_7834,N_7048,N_5356);
and U7835 (N_7835,N_5982,N_6441);
nor U7836 (N_7836,N_5255,N_6156);
nand U7837 (N_7837,N_7246,N_5639);
and U7838 (N_7838,N_7417,N_6964);
or U7839 (N_7839,N_5892,N_5800);
and U7840 (N_7840,N_6397,N_7457);
or U7841 (N_7841,N_7412,N_5747);
or U7842 (N_7842,N_5594,N_6795);
or U7843 (N_7843,N_7498,N_5616);
nand U7844 (N_7844,N_7082,N_5110);
nor U7845 (N_7845,N_6183,N_5860);
and U7846 (N_7846,N_6481,N_5796);
and U7847 (N_7847,N_7051,N_6926);
nor U7848 (N_7848,N_5144,N_5032);
and U7849 (N_7849,N_6445,N_6634);
or U7850 (N_7850,N_7491,N_5941);
nand U7851 (N_7851,N_5855,N_5739);
nand U7852 (N_7852,N_7384,N_5166);
nand U7853 (N_7853,N_7266,N_7169);
or U7854 (N_7854,N_5811,N_7388);
or U7855 (N_7855,N_5932,N_5961);
nand U7856 (N_7856,N_5100,N_5715);
nand U7857 (N_7857,N_6412,N_6332);
and U7858 (N_7858,N_7115,N_6201);
nand U7859 (N_7859,N_5751,N_6906);
or U7860 (N_7860,N_6319,N_5656);
nand U7861 (N_7861,N_6681,N_7474);
or U7862 (N_7862,N_7108,N_5904);
xnor U7863 (N_7863,N_6424,N_7226);
or U7864 (N_7864,N_5847,N_6797);
and U7865 (N_7865,N_7047,N_6238);
nand U7866 (N_7866,N_6515,N_5979);
xor U7867 (N_7867,N_5890,N_6103);
nand U7868 (N_7868,N_5140,N_7276);
or U7869 (N_7869,N_6222,N_5062);
or U7870 (N_7870,N_5859,N_7092);
or U7871 (N_7871,N_6339,N_5186);
and U7872 (N_7872,N_5920,N_6563);
or U7873 (N_7873,N_5682,N_5358);
or U7874 (N_7874,N_6529,N_6849);
nor U7875 (N_7875,N_5221,N_5571);
and U7876 (N_7876,N_7473,N_6062);
or U7877 (N_7877,N_6711,N_5649);
nor U7878 (N_7878,N_6171,N_5023);
or U7879 (N_7879,N_6709,N_5491);
or U7880 (N_7880,N_7306,N_7348);
nor U7881 (N_7881,N_7329,N_5287);
or U7882 (N_7882,N_6697,N_5805);
and U7883 (N_7883,N_6050,N_5330);
nand U7884 (N_7884,N_5954,N_5147);
or U7885 (N_7885,N_7458,N_7168);
nor U7886 (N_7886,N_6632,N_5240);
or U7887 (N_7887,N_6900,N_5913);
nand U7888 (N_7888,N_7330,N_5444);
or U7889 (N_7889,N_5426,N_7084);
nor U7890 (N_7890,N_5317,N_6396);
nor U7891 (N_7891,N_5312,N_6242);
nor U7892 (N_7892,N_6858,N_5459);
or U7893 (N_7893,N_7186,N_5045);
or U7894 (N_7894,N_6159,N_5306);
or U7895 (N_7895,N_5565,N_5679);
or U7896 (N_7896,N_6907,N_6860);
and U7897 (N_7897,N_5099,N_7344);
nand U7898 (N_7898,N_5438,N_6569);
or U7899 (N_7899,N_5382,N_5956);
nand U7900 (N_7900,N_5909,N_7031);
and U7901 (N_7901,N_6812,N_6593);
nor U7902 (N_7902,N_7477,N_6438);
nand U7903 (N_7903,N_6595,N_7162);
and U7904 (N_7904,N_5777,N_5939);
nor U7905 (N_7905,N_5124,N_6859);
nand U7906 (N_7906,N_6389,N_7452);
nand U7907 (N_7907,N_5486,N_6951);
nand U7908 (N_7908,N_5989,N_7001);
and U7909 (N_7909,N_6895,N_7046);
nand U7910 (N_7910,N_7126,N_6611);
and U7911 (N_7911,N_6323,N_6546);
nor U7912 (N_7912,N_5249,N_6774);
nand U7913 (N_7913,N_5745,N_6169);
nor U7914 (N_7914,N_5637,N_5325);
nor U7915 (N_7915,N_6863,N_6225);
nand U7916 (N_7916,N_6381,N_6779);
nor U7917 (N_7917,N_6333,N_5460);
nor U7918 (N_7918,N_5123,N_6787);
or U7919 (N_7919,N_6678,N_5198);
nor U7920 (N_7920,N_7304,N_5305);
nand U7921 (N_7921,N_6717,N_6631);
and U7922 (N_7922,N_5053,N_6973);
nor U7923 (N_7923,N_6202,N_5661);
nor U7924 (N_7924,N_6700,N_5792);
nor U7925 (N_7925,N_6579,N_6240);
nor U7926 (N_7926,N_6276,N_6035);
or U7927 (N_7927,N_7033,N_6749);
nor U7928 (N_7928,N_6684,N_5667);
nor U7929 (N_7929,N_5504,N_7496);
nor U7930 (N_7930,N_5901,N_7363);
or U7931 (N_7931,N_6567,N_6637);
and U7932 (N_7932,N_7396,N_6629);
nor U7933 (N_7933,N_5948,N_6435);
or U7934 (N_7934,N_6357,N_5479);
nand U7935 (N_7935,N_6203,N_6586);
or U7936 (N_7936,N_5266,N_7326);
and U7937 (N_7937,N_7376,N_5820);
and U7938 (N_7938,N_6927,N_6426);
or U7939 (N_7939,N_6280,N_6785);
nor U7940 (N_7940,N_6654,N_7321);
or U7941 (N_7941,N_6258,N_7017);
and U7942 (N_7942,N_5967,N_6834);
or U7943 (N_7943,N_5782,N_5429);
and U7944 (N_7944,N_5308,N_6253);
and U7945 (N_7945,N_7229,N_7191);
or U7946 (N_7946,N_6359,N_6137);
nand U7947 (N_7947,N_7423,N_5494);
nor U7948 (N_7948,N_6153,N_7097);
or U7949 (N_7949,N_6782,N_7081);
nor U7950 (N_7950,N_5891,N_5204);
nand U7951 (N_7951,N_6982,N_5699);
nor U7952 (N_7952,N_6488,N_5761);
and U7953 (N_7953,N_6525,N_6271);
and U7954 (N_7954,N_7271,N_6723);
and U7955 (N_7955,N_7301,N_5303);
and U7956 (N_7956,N_7198,N_6361);
or U7957 (N_7957,N_6022,N_5173);
or U7958 (N_7958,N_5610,N_5767);
xnor U7959 (N_7959,N_5688,N_7116);
xor U7960 (N_7960,N_5112,N_6427);
nor U7961 (N_7961,N_5789,N_6413);
and U7962 (N_7962,N_6651,N_7095);
nor U7963 (N_7963,N_7056,N_5042);
nand U7964 (N_7964,N_5540,N_5741);
or U7965 (N_7965,N_5214,N_7497);
or U7966 (N_7966,N_7303,N_7285);
or U7967 (N_7967,N_5947,N_6471);
or U7968 (N_7968,N_5755,N_7171);
nor U7969 (N_7969,N_5543,N_7482);
or U7970 (N_7970,N_5732,N_6065);
nor U7971 (N_7971,N_6724,N_6069);
or U7972 (N_7972,N_5907,N_6030);
nor U7973 (N_7973,N_5279,N_5229);
and U7974 (N_7974,N_7130,N_6642);
nor U7975 (N_7975,N_6913,N_7394);
or U7976 (N_7976,N_5660,N_5621);
nand U7977 (N_7977,N_5576,N_5280);
nor U7978 (N_7978,N_7449,N_6340);
nor U7979 (N_7979,N_5754,N_5817);
nand U7980 (N_7980,N_5089,N_6037);
or U7981 (N_7981,N_7218,N_5833);
nor U7982 (N_7982,N_6953,N_6521);
and U7983 (N_7983,N_5622,N_6422);
or U7984 (N_7984,N_6076,N_5764);
nor U7985 (N_7985,N_6154,N_7203);
nor U7986 (N_7986,N_6652,N_6009);
and U7987 (N_7987,N_6236,N_5072);
and U7988 (N_7988,N_5786,N_5192);
nor U7989 (N_7989,N_6117,N_5081);
nor U7990 (N_7990,N_5242,N_5903);
and U7991 (N_7991,N_6983,N_7137);
nor U7992 (N_7992,N_6006,N_6769);
and U7993 (N_7993,N_6673,N_5285);
or U7994 (N_7994,N_5830,N_7153);
and U7995 (N_7995,N_6057,N_7456);
nor U7996 (N_7996,N_6049,N_5218);
and U7997 (N_7997,N_6206,N_6443);
nand U7998 (N_7998,N_5595,N_6324);
nand U7999 (N_7999,N_5468,N_6436);
or U8000 (N_8000,N_6852,N_7104);
and U8001 (N_8001,N_6186,N_5179);
nand U8002 (N_8002,N_6822,N_5795);
nand U8003 (N_8003,N_7222,N_6287);
or U8004 (N_8004,N_5728,N_6375);
nor U8005 (N_8005,N_7098,N_6534);
nand U8006 (N_8006,N_5269,N_5421);
or U8007 (N_8007,N_5184,N_5374);
nand U8008 (N_8008,N_5759,N_7061);
or U8009 (N_8009,N_6893,N_6536);
nor U8010 (N_8010,N_5355,N_5453);
and U8011 (N_8011,N_5195,N_6325);
and U8012 (N_8012,N_7405,N_5283);
or U8013 (N_8013,N_5148,N_6892);
nor U8014 (N_8014,N_7176,N_5030);
or U8015 (N_8015,N_6173,N_5868);
nand U8016 (N_8016,N_7280,N_6191);
nor U8017 (N_8017,N_7111,N_6104);
nor U8018 (N_8018,N_6690,N_5821);
nand U8019 (N_8019,N_5627,N_5685);
or U8020 (N_8020,N_6461,N_6655);
nor U8021 (N_8021,N_5091,N_5625);
nand U8022 (N_8022,N_6370,N_6451);
nand U8023 (N_8023,N_7231,N_7478);
nor U8024 (N_8024,N_6449,N_6979);
and U8025 (N_8025,N_7206,N_6387);
nand U8026 (N_8026,N_5237,N_5928);
and U8027 (N_8027,N_7312,N_6130);
or U8028 (N_8028,N_7267,N_5944);
nand U8029 (N_8029,N_7319,N_5619);
and U8030 (N_8030,N_6346,N_6420);
or U8031 (N_8031,N_5526,N_6077);
and U8032 (N_8032,N_6193,N_6910);
nor U8033 (N_8033,N_6824,N_5570);
nor U8034 (N_8034,N_5883,N_6761);
nand U8035 (N_8035,N_5005,N_6526);
nand U8036 (N_8036,N_7163,N_6229);
and U8037 (N_8037,N_6539,N_5309);
nand U8038 (N_8038,N_5587,N_6990);
and U8039 (N_8039,N_7235,N_5273);
and U8040 (N_8040,N_6423,N_6905);
nor U8041 (N_8041,N_6823,N_7252);
or U8042 (N_8042,N_7345,N_5152);
or U8043 (N_8043,N_5098,N_5958);
and U8044 (N_8044,N_7210,N_5001);
nand U8045 (N_8045,N_6981,N_7463);
nor U8046 (N_8046,N_7347,N_7354);
nor U8047 (N_8047,N_5684,N_6740);
nor U8048 (N_8048,N_7143,N_5710);
or U8049 (N_8049,N_6607,N_6310);
and U8050 (N_8050,N_7418,N_5375);
and U8051 (N_8051,N_7135,N_5057);
and U8052 (N_8052,N_5288,N_7328);
nor U8053 (N_8053,N_6486,N_5927);
nand U8054 (N_8054,N_7434,N_5579);
nor U8055 (N_8055,N_7230,N_6482);
and U8056 (N_8056,N_6448,N_5369);
nor U8057 (N_8057,N_6224,N_7290);
nor U8058 (N_8058,N_6814,N_7275);
nand U8059 (N_8059,N_7148,N_5134);
nand U8060 (N_8060,N_6692,N_7392);
nor U8061 (N_8061,N_6286,N_5068);
and U8062 (N_8062,N_7364,N_5863);
nand U8063 (N_8063,N_6425,N_6393);
or U8064 (N_8064,N_5681,N_7085);
and U8065 (N_8065,N_6584,N_7221);
or U8066 (N_8066,N_5670,N_7037);
or U8067 (N_8067,N_6602,N_5291);
nand U8068 (N_8068,N_7373,N_7060);
and U8069 (N_8069,N_5087,N_5417);
nand U8070 (N_8070,N_7237,N_5386);
and U8071 (N_8071,N_6141,N_6836);
and U8072 (N_8072,N_6944,N_5714);
or U8073 (N_8073,N_5963,N_7141);
and U8074 (N_8074,N_5293,N_6988);
nand U8075 (N_8075,N_6640,N_6517);
nand U8076 (N_8076,N_6653,N_5952);
nand U8077 (N_8077,N_5051,N_6181);
or U8078 (N_8078,N_5270,N_5131);
and U8079 (N_8079,N_6409,N_5321);
nor U8080 (N_8080,N_6815,N_5865);
nand U8081 (N_8081,N_5804,N_6878);
and U8082 (N_8082,N_5020,N_5474);
or U8083 (N_8083,N_5310,N_5006);
nand U8084 (N_8084,N_5582,N_6805);
nand U8085 (N_8085,N_6307,N_5550);
and U8086 (N_8086,N_6081,N_6021);
or U8087 (N_8087,N_6266,N_5048);
and U8088 (N_8088,N_6312,N_6184);
and U8089 (N_8089,N_7374,N_5315);
nand U8090 (N_8090,N_7197,N_5915);
nor U8091 (N_8091,N_6731,N_6282);
nor U8092 (N_8092,N_7150,N_7090);
or U8093 (N_8093,N_5919,N_7416);
and U8094 (N_8094,N_6572,N_6999);
or U8095 (N_8095,N_6316,N_7369);
or U8096 (N_8096,N_5097,N_5065);
or U8097 (N_8097,N_6221,N_6735);
and U8098 (N_8098,N_6087,N_5377);
xor U8099 (N_8099,N_6013,N_6394);
nor U8100 (N_8100,N_6264,N_5516);
and U8101 (N_8101,N_7202,N_6406);
or U8102 (N_8102,N_5239,N_7074);
nand U8103 (N_8103,N_5787,N_6400);
and U8104 (N_8104,N_5106,N_6918);
nand U8105 (N_8105,N_6223,N_7105);
nor U8106 (N_8106,N_6996,N_5326);
nand U8107 (N_8107,N_6245,N_7404);
nand U8108 (N_8108,N_6682,N_6380);
and U8109 (N_8109,N_6440,N_7386);
and U8110 (N_8110,N_6658,N_6122);
nand U8111 (N_8111,N_5502,N_5721);
nor U8112 (N_8112,N_6594,N_6896);
nor U8113 (N_8113,N_5257,N_6829);
or U8114 (N_8114,N_6483,N_6502);
nor U8115 (N_8115,N_5608,N_6279);
or U8116 (N_8116,N_5985,N_6597);
and U8117 (N_8117,N_6841,N_5034);
nor U8118 (N_8118,N_6523,N_6073);
or U8119 (N_8119,N_6986,N_6460);
and U8120 (N_8120,N_7436,N_5806);
nor U8121 (N_8121,N_7346,N_6950);
nand U8122 (N_8122,N_6454,N_7015);
nor U8123 (N_8123,N_5518,N_6876);
or U8124 (N_8124,N_6039,N_7177);
or U8125 (N_8125,N_5366,N_7494);
and U8126 (N_8126,N_6739,N_6962);
nand U8127 (N_8127,N_6024,N_5142);
nand U8128 (N_8128,N_6498,N_7005);
or U8129 (N_8129,N_6930,N_7415);
nor U8130 (N_8130,N_5547,N_5372);
or U8131 (N_8131,N_6758,N_5596);
and U8132 (N_8132,N_6095,N_5389);
and U8133 (N_8133,N_6114,N_6801);
nor U8134 (N_8134,N_6078,N_5212);
nand U8135 (N_8135,N_5531,N_6621);
nor U8136 (N_8136,N_6993,N_5916);
and U8137 (N_8137,N_7273,N_6733);
nor U8138 (N_8138,N_5442,N_5364);
and U8139 (N_8139,N_6998,N_6497);
and U8140 (N_8140,N_5430,N_6265);
nand U8141 (N_8141,N_6147,N_7013);
nand U8142 (N_8142,N_6175,N_6751);
or U8143 (N_8143,N_5211,N_5499);
and U8144 (N_8144,N_6002,N_7282);
nand U8145 (N_8145,N_6957,N_6507);
nor U8146 (N_8146,N_5357,N_5877);
nor U8147 (N_8147,N_6038,N_5671);
nand U8148 (N_8148,N_7160,N_5404);
nand U8149 (N_8149,N_5299,N_5052);
and U8150 (N_8150,N_5296,N_6196);
nor U8151 (N_8151,N_6365,N_5542);
nor U8152 (N_8152,N_5088,N_6485);
nand U8153 (N_8153,N_5895,N_7262);
and U8154 (N_8154,N_5509,N_5281);
and U8155 (N_8155,N_7341,N_5870);
or U8156 (N_8156,N_6583,N_5385);
and U8157 (N_8157,N_5252,N_7040);
and U8158 (N_8158,N_5470,N_6940);
nor U8159 (N_8159,N_7127,N_5054);
nor U8160 (N_8160,N_5823,N_5862);
and U8161 (N_8161,N_5416,N_5996);
nor U8162 (N_8162,N_6063,N_6955);
or U8163 (N_8163,N_6672,N_5545);
and U8164 (N_8164,N_7110,N_6656);
nor U8165 (N_8165,N_5039,N_7472);
nor U8166 (N_8166,N_6931,N_6166);
nor U8167 (N_8167,N_6591,N_5881);
or U8168 (N_8168,N_5025,N_7320);
and U8169 (N_8169,N_7083,N_6194);
or U8170 (N_8170,N_6172,N_6200);
nand U8171 (N_8171,N_5521,N_5851);
nor U8172 (N_8172,N_5672,N_5557);
or U8173 (N_8173,N_6418,N_6466);
and U8174 (N_8174,N_6428,N_7391);
nand U8175 (N_8175,N_5241,N_6472);
nand U8176 (N_8176,N_5864,N_7180);
and U8177 (N_8177,N_7028,N_6309);
nand U8178 (N_8178,N_5471,N_7200);
and U8179 (N_8179,N_5139,N_6620);
nor U8180 (N_8180,N_5770,N_5599);
or U8181 (N_8181,N_6972,N_6118);
nor U8182 (N_8182,N_7069,N_5638);
nand U8183 (N_8183,N_5683,N_6721);
or U8184 (N_8184,N_7410,N_7286);
nand U8185 (N_8185,N_5569,N_6367);
nand U8186 (N_8186,N_5973,N_5802);
nor U8187 (N_8187,N_6887,N_5529);
and U8188 (N_8188,N_6767,N_5659);
nand U8189 (N_8189,N_7400,N_6351);
and U8190 (N_8190,N_5505,N_5631);
and U8191 (N_8191,N_6080,N_6914);
nand U8192 (N_8192,N_6559,N_6138);
nor U8193 (N_8193,N_6262,N_6108);
nand U8194 (N_8194,N_7408,N_6541);
or U8195 (N_8195,N_6870,N_7470);
nor U8196 (N_8196,N_6376,N_6036);
or U8197 (N_8197,N_5103,N_5294);
nand U8198 (N_8198,N_6581,N_7401);
and U8199 (N_8199,N_7009,N_7189);
nor U8200 (N_8200,N_6120,N_5674);
nand U8201 (N_8201,N_6052,N_6873);
nor U8202 (N_8202,N_6487,N_6615);
and U8203 (N_8203,N_5409,N_7367);
nand U8204 (N_8204,N_5994,N_5829);
or U8205 (N_8205,N_6971,N_5809);
nor U8206 (N_8206,N_7307,N_5073);
or U8207 (N_8207,N_6504,N_5955);
nor U8208 (N_8208,N_5597,N_5783);
and U8209 (N_8209,N_5871,N_5905);
or U8210 (N_8210,N_6289,N_6608);
nand U8211 (N_8211,N_6124,N_5208);
nand U8212 (N_8212,N_6636,N_6407);
nor U8213 (N_8213,N_5259,N_5044);
and U8214 (N_8214,N_6789,N_5424);
nand U8215 (N_8215,N_6139,N_5983);
nand U8216 (N_8216,N_5302,N_5101);
and U8217 (N_8217,N_5116,N_5533);
and U8218 (N_8218,N_6759,N_6756);
nor U8219 (N_8219,N_5757,N_6437);
nor U8220 (N_8220,N_6027,N_6669);
nand U8221 (N_8221,N_7311,N_6809);
or U8222 (N_8222,N_5640,N_7164);
and U8223 (N_8223,N_6379,N_6489);
nand U8224 (N_8224,N_6297,N_7431);
nand U8225 (N_8225,N_5908,N_5591);
xnor U8226 (N_8226,N_6588,N_5197);
nor U8227 (N_8227,N_6301,N_6328);
nand U8228 (N_8228,N_7043,N_5893);
or U8229 (N_8229,N_5648,N_6722);
nor U8230 (N_8230,N_7212,N_5175);
or U8231 (N_8231,N_5466,N_5885);
and U8232 (N_8232,N_6404,N_7080);
and U8233 (N_8233,N_5115,N_5345);
or U8234 (N_8234,N_5807,N_5130);
nand U8235 (N_8235,N_5498,N_6392);
and U8236 (N_8236,N_7427,N_5912);
nor U8237 (N_8237,N_7409,N_6564);
nand U8238 (N_8238,N_6868,N_6562);
nand U8239 (N_8239,N_6720,N_6092);
or U8240 (N_8240,N_6086,N_6921);
and U8241 (N_8241,N_6119,N_6671);
and U8242 (N_8242,N_5262,N_6051);
nor U8243 (N_8243,N_7035,N_6627);
and U8244 (N_8244,N_5258,N_5886);
nor U8245 (N_8245,N_6619,N_5464);
nor U8246 (N_8246,N_5537,N_5008);
nor U8247 (N_8247,N_5428,N_5047);
and U8248 (N_8248,N_7365,N_5284);
or U8249 (N_8249,N_6126,N_5607);
nor U8250 (N_8250,N_7406,N_5609);
nor U8251 (N_8251,N_6974,N_6810);
and U8252 (N_8252,N_7337,N_5669);
and U8253 (N_8253,N_5507,N_5436);
and U8254 (N_8254,N_6476,N_7389);
or U8255 (N_8255,N_7151,N_6128);
or U8256 (N_8256,N_6373,N_5598);
or U8257 (N_8257,N_5007,N_7075);
or U8258 (N_8258,N_5848,N_6363);
or U8259 (N_8259,N_5951,N_5882);
or U8260 (N_8260,N_6374,N_6272);
and U8261 (N_8261,N_7093,N_5692);
nor U8262 (N_8262,N_6639,N_5735);
or U8263 (N_8263,N_5384,N_5161);
and U8264 (N_8264,N_7249,N_6992);
xor U8265 (N_8265,N_6155,N_5523);
or U8266 (N_8266,N_6244,N_7483);
nor U8267 (N_8267,N_6293,N_6587);
or U8268 (N_8268,N_6556,N_5432);
nor U8269 (N_8269,N_5931,N_6028);
and U8270 (N_8270,N_5675,N_6867);
nand U8271 (N_8271,N_5668,N_6945);
nor U8272 (N_8272,N_5836,N_5803);
or U8273 (N_8273,N_7147,N_6661);
and U8274 (N_8274,N_6622,N_6160);
nor U8275 (N_8275,N_6267,N_6685);
and U8276 (N_8276,N_5066,N_6904);
nand U8277 (N_8277,N_7453,N_5618);
and U8278 (N_8278,N_5127,N_5082);
nand U8279 (N_8279,N_6531,N_5940);
and U8280 (N_8280,N_5713,N_6663);
or U8281 (N_8281,N_5341,N_6135);
or U8282 (N_8282,N_5003,N_5233);
nor U8283 (N_8283,N_7314,N_7323);
nand U8284 (N_8284,N_5665,N_6516);
xor U8285 (N_8285,N_6446,N_6342);
or U8286 (N_8286,N_6248,N_5778);
and U8287 (N_8287,N_7379,N_7263);
nand U8288 (N_8288,N_7124,N_6804);
nor U8289 (N_8289,N_6075,N_6480);
or U8290 (N_8290,N_7010,N_6112);
or U8291 (N_8291,N_5365,N_6491);
or U8292 (N_8292,N_5071,N_5253);
nand U8293 (N_8293,N_5009,N_6799);
nand U8294 (N_8294,N_7349,N_6260);
nor U8295 (N_8295,N_7055,N_6702);
nand U8296 (N_8296,N_6189,N_5070);
nand U8297 (N_8297,N_5629,N_7265);
or U8298 (N_8298,N_5719,N_6023);
nand U8299 (N_8299,N_5420,N_6259);
nor U8300 (N_8300,N_5522,N_6696);
or U8301 (N_8301,N_5888,N_6865);
nand U8302 (N_8302,N_6099,N_5322);
or U8303 (N_8303,N_6019,N_5743);
and U8304 (N_8304,N_5448,N_6032);
nor U8305 (N_8305,N_7042,N_6734);
and U8306 (N_8306,N_6060,N_6688);
and U8307 (N_8307,N_5185,N_7136);
nand U8308 (N_8308,N_6214,N_5874);
nand U8309 (N_8309,N_5921,N_6984);
nand U8310 (N_8310,N_7484,N_5986);
or U8311 (N_8311,N_7238,N_5752);
nor U8312 (N_8312,N_5922,N_5427);
or U8313 (N_8313,N_6343,N_6305);
or U8314 (N_8314,N_5457,N_5037);
or U8315 (N_8315,N_7492,N_6453);
nand U8316 (N_8316,N_6705,N_5965);
nor U8317 (N_8317,N_5380,N_5403);
nand U8318 (N_8318,N_7370,N_6366);
nor U8319 (N_8319,N_6949,N_5578);
and U8320 (N_8320,N_7087,N_5562);
nand U8321 (N_8321,N_5217,N_5957);
nand U8322 (N_8322,N_5225,N_5664);
nand U8323 (N_8323,N_7292,N_5297);
or U8324 (N_8324,N_6362,N_6975);
nor U8325 (N_8325,N_5731,N_6808);
nand U8326 (N_8326,N_5534,N_7481);
and U8327 (N_8327,N_7245,N_6842);
and U8328 (N_8328,N_5925,N_5331);
or U8329 (N_8329,N_5138,N_6306);
nand U8330 (N_8330,N_5397,N_6777);
nor U8331 (N_8331,N_6158,N_5473);
nand U8332 (N_8332,N_7260,N_5702);
or U8333 (N_8333,N_6237,N_6576);
nor U8334 (N_8334,N_6875,N_6614);
nor U8335 (N_8335,N_5080,N_5500);
nand U8336 (N_8336,N_5554,N_5245);
and U8337 (N_8337,N_5984,N_6261);
nand U8338 (N_8338,N_6912,N_5114);
and U8339 (N_8339,N_6872,N_5079);
nand U8340 (N_8340,N_5853,N_5387);
and U8341 (N_8341,N_6178,N_6313);
or U8342 (N_8342,N_6645,N_5063);
nand U8343 (N_8343,N_5125,N_5857);
nor U8344 (N_8344,N_6167,N_6290);
nand U8345 (N_8345,N_5349,N_6941);
and U8346 (N_8346,N_7302,N_5278);
or U8347 (N_8347,N_5525,N_5492);
nor U8348 (N_8348,N_6691,N_6592);
and U8349 (N_8349,N_7139,N_5923);
or U8350 (N_8350,N_6706,N_5524);
nand U8351 (N_8351,N_5154,N_6317);
and U8352 (N_8352,N_7123,N_7430);
and U8353 (N_8353,N_6561,N_7420);
or U8354 (N_8354,N_5135,N_6368);
nor U8355 (N_8355,N_6302,N_5415);
nand U8356 (N_8356,N_6903,N_6891);
nand U8357 (N_8357,N_5462,N_5781);
and U8358 (N_8358,N_7441,N_6687);
and U8359 (N_8359,N_5029,N_6939);
nand U8360 (N_8360,N_5170,N_7475);
nand U8361 (N_8361,N_5232,N_6250);
nor U8362 (N_8362,N_6410,N_7144);
nand U8363 (N_8363,N_6467,N_5196);
and U8364 (N_8364,N_5844,N_5236);
and U8365 (N_8365,N_7305,N_5867);
nor U8366 (N_8366,N_5469,N_7357);
or U8367 (N_8367,N_6736,N_7253);
and U8368 (N_8368,N_6285,N_5724);
and U8369 (N_8369,N_5564,N_7244);
and U8370 (N_8370,N_5394,N_5604);
nor U8371 (N_8371,N_6802,N_5647);
nor U8372 (N_8372,N_7125,N_5978);
nand U8373 (N_8373,N_5151,N_5248);
and U8374 (N_8374,N_7489,N_6508);
nand U8375 (N_8375,N_6123,N_6922);
nand U8376 (N_8376,N_6384,N_7131);
nor U8377 (N_8377,N_5780,N_6819);
and U8378 (N_8378,N_6210,N_6246);
or U8379 (N_8379,N_7185,N_6219);
and U8380 (N_8380,N_7254,N_5383);
nor U8381 (N_8381,N_6641,N_7466);
and U8382 (N_8382,N_7133,N_5769);
or U8383 (N_8383,N_5643,N_6847);
nand U8384 (N_8384,N_5439,N_7072);
nor U8385 (N_8385,N_7465,N_7413);
or U8386 (N_8386,N_5268,N_5265);
and U8387 (N_8387,N_6046,N_5774);
or U8388 (N_8388,N_6772,N_7214);
nand U8389 (N_8389,N_6577,N_6358);
nor U8390 (N_8390,N_5076,N_5946);
nand U8391 (N_8391,N_6216,N_7032);
and U8392 (N_8392,N_7316,N_5902);
and U8393 (N_8393,N_5510,N_6649);
or U8394 (N_8394,N_6589,N_5879);
nand U8395 (N_8395,N_5972,N_5878);
and U8396 (N_8396,N_7113,N_6234);
and U8397 (N_8397,N_6585,N_7467);
and U8398 (N_8398,N_7487,N_5617);
nor U8399 (N_8399,N_6233,N_6712);
and U8400 (N_8400,N_5314,N_5641);
and U8401 (N_8401,N_5727,N_5481);
nand U8402 (N_8402,N_7455,N_6987);
and U8403 (N_8403,N_7353,N_6228);
and U8404 (N_8404,N_6798,N_5900);
nand U8405 (N_8405,N_5286,N_6071);
nand U8406 (N_8406,N_6535,N_7076);
and U8407 (N_8407,N_7138,N_5636);
or U8408 (N_8408,N_6256,N_5021);
nor U8409 (N_8409,N_6320,N_7088);
nand U8410 (N_8410,N_6199,N_6630);
and U8411 (N_8411,N_5945,N_5856);
nand U8412 (N_8412,N_6098,N_6715);
nor U8413 (N_8413,N_5222,N_6714);
nor U8414 (N_8414,N_6748,N_6826);
and U8415 (N_8415,N_7219,N_5169);
and U8416 (N_8416,N_5105,N_7211);
nor U8417 (N_8417,N_5730,N_5159);
nand U8418 (N_8418,N_7077,N_7066);
and U8419 (N_8419,N_5756,N_5368);
nor U8420 (N_8420,N_5697,N_6315);
nand U8421 (N_8421,N_7024,N_6001);
or U8422 (N_8422,N_7118,N_5929);
nor U8423 (N_8423,N_6281,N_5695);
or U8424 (N_8424,N_5869,N_6959);
nand U8425 (N_8425,N_5976,N_5443);
nand U8426 (N_8426,N_6145,N_6377);
or U8427 (N_8427,N_5760,N_6625);
or U8428 (N_8428,N_6303,N_5813);
nor U8429 (N_8429,N_6372,N_7239);
and U8430 (N_8430,N_5938,N_6624);
and U8431 (N_8431,N_5906,N_5899);
nor U8432 (N_8432,N_7317,N_5104);
nand U8433 (N_8433,N_6174,N_5816);
and U8434 (N_8434,N_6209,N_5601);
nor U8435 (N_8435,N_7175,N_5004);
and U8436 (N_8436,N_7157,N_6574);
nor U8437 (N_8437,N_7078,N_6213);
and U8438 (N_8438,N_6337,N_6911);
nor U8439 (N_8439,N_6152,N_6942);
nor U8440 (N_8440,N_5164,N_7499);
or U8441 (N_8441,N_5337,N_6603);
nand U8442 (N_8442,N_5527,N_6928);
and U8443 (N_8443,N_5691,N_5129);
or U8444 (N_8444,N_6149,N_5583);
nand U8445 (N_8445,N_5108,N_5441);
and U8446 (N_8446,N_6015,N_6398);
and U8447 (N_8447,N_6857,N_7025);
or U8448 (N_8448,N_6459,N_6518);
nor U8449 (N_8449,N_5517,N_7089);
xnor U8450 (N_8450,N_6960,N_5246);
nand U8451 (N_8451,N_6478,N_7008);
and U8452 (N_8452,N_6348,N_6694);
and U8453 (N_8453,N_7146,N_5143);
nand U8454 (N_8454,N_5825,N_5623);
nor U8455 (N_8455,N_6356,N_6877);
and U8456 (N_8456,N_5630,N_6195);
or U8457 (N_8457,N_6503,N_5235);
and U8458 (N_8458,N_5122,N_5028);
or U8459 (N_8459,N_5775,N_5224);
and U8460 (N_8460,N_5990,N_7196);
nand U8461 (N_8461,N_5199,N_5835);
or U8462 (N_8462,N_6116,N_7114);
nand U8463 (N_8463,N_5096,N_6909);
or U8464 (N_8464,N_6832,N_5086);
nand U8465 (N_8465,N_6344,N_7045);
nand U8466 (N_8466,N_7283,N_6299);
nor U8467 (N_8467,N_6755,N_7149);
nor U8468 (N_8468,N_5347,N_6058);
nor U8469 (N_8469,N_5153,N_6163);
nor U8470 (N_8470,N_7240,N_6626);
and U8471 (N_8471,N_6674,N_5729);
nand U8472 (N_8472,N_5396,N_7261);
and U8473 (N_8473,N_5094,N_6450);
or U8474 (N_8474,N_6730,N_5970);
xnor U8475 (N_8475,N_6284,N_7296);
and U8476 (N_8476,N_7155,N_7393);
nand U8477 (N_8477,N_5876,N_7232);
and U8478 (N_8478,N_7016,N_5488);
and U8479 (N_8479,N_5917,N_5677);
nand U8480 (N_8480,N_5238,N_5520);
nor U8481 (N_8481,N_6268,N_6766);
and U8482 (N_8482,N_6932,N_7335);
and U8483 (N_8483,N_7134,N_5215);
and U8484 (N_8484,N_7193,N_6509);
or U8485 (N_8485,N_6845,N_5350);
nand U8486 (N_8486,N_6208,N_6018);
nand U8487 (N_8487,N_5465,N_6967);
or U8488 (N_8488,N_5810,N_5740);
nand U8489 (N_8489,N_6142,N_6288);
xor U8490 (N_8490,N_6129,N_5704);
or U8491 (N_8491,N_7053,N_5613);
and U8492 (N_8492,N_7274,N_6943);
xor U8493 (N_8493,N_5655,N_5875);
and U8494 (N_8494,N_6871,N_5298);
nor U8495 (N_8495,N_5455,N_6395);
nor U8496 (N_8496,N_6110,N_7050);
or U8497 (N_8497,N_5205,N_6125);
and U8498 (N_8498,N_5370,N_5348);
nand U8499 (N_8499,N_6813,N_7041);
and U8500 (N_8500,N_7132,N_5109);
and U8501 (N_8501,N_6969,N_5959);
and U8502 (N_8502,N_5077,N_7325);
or U8503 (N_8503,N_5703,N_5392);
or U8504 (N_8504,N_7112,N_6270);
nand U8505 (N_8505,N_7318,N_6716);
nand U8506 (N_8506,N_6402,N_6566);
or U8507 (N_8507,N_7383,N_7270);
nand U8508 (N_8508,N_5711,N_5673);
and U8509 (N_8509,N_5107,N_5223);
and U8510 (N_8510,N_6464,N_7181);
or U8511 (N_8511,N_5339,N_6713);
or U8512 (N_8512,N_6947,N_7279);
and U8513 (N_8513,N_6590,N_5067);
nand U8514 (N_8514,N_5801,N_5163);
and U8515 (N_8515,N_5918,N_6355);
nor U8516 (N_8516,N_6227,N_6161);
or U8517 (N_8517,N_5911,N_6543);
nor U8518 (N_8518,N_5506,N_7067);
nand U8519 (N_8519,N_6770,N_5277);
or U8520 (N_8520,N_5118,N_7020);
and U8521 (N_8521,N_6369,N_6230);
nand U8522 (N_8522,N_5568,N_5773);
and U8523 (N_8523,N_6091,N_6010);
nor U8524 (N_8524,N_7462,N_5015);
nor U8525 (N_8525,N_6894,N_6980);
or U8526 (N_8526,N_6680,N_6935);
or U8527 (N_8527,N_6550,N_5351);
nand U8528 (N_8528,N_6606,N_5600);
nor U8529 (N_8529,N_6532,N_7014);
or U8530 (N_8530,N_6745,N_6330);
nor U8531 (N_8531,N_5213,N_5180);
nand U8532 (N_8532,N_7006,N_5126);
or U8533 (N_8533,N_6399,N_5132);
or U8534 (N_8534,N_5960,N_6251);
or U8535 (N_8535,N_7269,N_6623);
and U8536 (N_8536,N_6232,N_5742);
nor U8537 (N_8537,N_7459,N_5799);
and U8538 (N_8538,N_7241,N_7444);
nand U8539 (N_8539,N_7358,N_6294);
nand U8540 (N_8540,N_5508,N_5758);
and U8541 (N_8541,N_6617,N_6792);
and U8542 (N_8542,N_6349,N_6029);
nor U8543 (N_8543,N_7068,N_6433);
nand U8544 (N_8544,N_6157,N_7268);
and U8545 (N_8545,N_6524,N_6314);
nand U8546 (N_8546,N_5549,N_7256);
or U8547 (N_8547,N_5346,N_5056);
or U8548 (N_8548,N_6693,N_5036);
nand U8549 (N_8549,N_6961,N_7052);
and U8550 (N_8550,N_5160,N_6646);
nand U8551 (N_8551,N_7154,N_5493);
and U8552 (N_8552,N_6473,N_5589);
nand U8553 (N_8553,N_6648,N_5272);
and U8554 (N_8554,N_7209,N_5461);
and U8555 (N_8555,N_5999,N_7419);
and U8556 (N_8556,N_5002,N_6917);
nand U8557 (N_8557,N_5316,N_5178);
nand U8558 (N_8558,N_6329,N_7044);
nand U8559 (N_8559,N_6821,N_6833);
or U8560 (N_8560,N_5791,N_6757);
and U8561 (N_8561,N_6936,N_6134);
or U8562 (N_8562,N_7490,N_7432);
or U8563 (N_8563,N_6043,N_6806);
and U8564 (N_8564,N_5998,N_5133);
nor U8565 (N_8565,N_5974,N_5553);
nand U8566 (N_8566,N_6582,N_5146);
and U8567 (N_8567,N_6215,N_5484);
nand U8568 (N_8568,N_5371,N_6698);
or U8569 (N_8569,N_7159,N_5267);
or U8570 (N_8570,N_5022,N_7036);
nor U8571 (N_8571,N_5026,N_5010);
and U8572 (N_8572,N_5975,N_5771);
or U8573 (N_8573,N_7471,N_5894);
nand U8574 (N_8574,N_7446,N_6417);
nand U8575 (N_8575,N_6066,N_6788);
nor U8576 (N_8576,N_6708,N_6109);
nor U8577 (N_8577,N_5483,N_5733);
nor U8578 (N_8578,N_7117,N_6364);
or U8579 (N_8579,N_6411,N_5680);
and U8580 (N_8580,N_5873,N_6760);
nand U8581 (N_8581,N_7182,N_5440);
or U8582 (N_8582,N_6151,N_7122);
or U8583 (N_8583,N_6901,N_5141);
nand U8584 (N_8584,N_6506,N_5167);
nor U8585 (N_8585,N_5749,N_5226);
nand U8586 (N_8586,N_6192,N_7385);
and U8587 (N_8587,N_7426,N_6679);
and U8588 (N_8588,N_6869,N_6465);
or U8589 (N_8589,N_6168,N_5230);
nand U8590 (N_8590,N_6666,N_6613);
nor U8591 (N_8591,N_7220,N_5950);
nor U8592 (N_8592,N_7004,N_6726);
and U8593 (N_8593,N_5933,N_5501);
or U8594 (N_8594,N_7224,N_5768);
nor U8595 (N_8595,N_5220,N_6780);
nand U8596 (N_8596,N_7387,N_6933);
nand U8597 (N_8597,N_5320,N_6439);
and U8598 (N_8598,N_6360,N_7277);
or U8599 (N_8599,N_6074,N_5324);
and U8600 (N_8600,N_5410,N_7070);
nor U8601 (N_8601,N_6177,N_7480);
and U8602 (N_8602,N_7107,N_6016);
nand U8603 (N_8603,N_6899,N_5837);
and U8604 (N_8604,N_6659,N_5155);
or U8605 (N_8605,N_6600,N_5846);
nand U8606 (N_8606,N_5585,N_6995);
and U8607 (N_8607,N_7272,N_6180);
or U8608 (N_8608,N_7223,N_6830);
nor U8609 (N_8609,N_6241,N_6025);
and U8610 (N_8610,N_5150,N_5535);
nor U8611 (N_8611,N_5300,N_6012);
and U8612 (N_8612,N_5171,N_6609);
or U8613 (N_8613,N_6710,N_5189);
or U8614 (N_8614,N_7403,N_7030);
or U8615 (N_8615,N_6321,N_5866);
nand U8616 (N_8616,N_7039,N_6292);
and U8617 (N_8617,N_6827,N_6353);
nor U8618 (N_8618,N_6925,N_5693);
or U8619 (N_8619,N_6638,N_5872);
nor U8620 (N_8620,N_5332,N_7309);
nand U8621 (N_8621,N_5503,N_6610);
nand U8622 (N_8622,N_5798,N_6683);
or U8623 (N_8623,N_5251,N_6703);
and U8624 (N_8624,N_6430,N_6864);
and U8625 (N_8625,N_6837,N_6414);
and U8626 (N_8626,N_6796,N_6778);
or U8627 (N_8627,N_6958,N_6675);
nor U8628 (N_8628,N_6985,N_6499);
nand U8629 (N_8629,N_5572,N_6391);
nor U8630 (N_8630,N_6084,N_6354);
nand U8631 (N_8631,N_5128,N_6300);
nor U8632 (N_8632,N_6345,N_7026);
and U8633 (N_8633,N_6571,N_6204);
and U8634 (N_8634,N_5379,N_7454);
or U8635 (N_8635,N_6677,N_5790);
and U8636 (N_8636,N_7049,N_5567);
nor U8637 (N_8637,N_5997,N_5723);
nand U8638 (N_8638,N_5575,N_5896);
and U8639 (N_8639,N_6650,N_6239);
and U8640 (N_8640,N_5040,N_6390);
and U8641 (N_8641,N_5360,N_7375);
nand U8642 (N_8642,N_7187,N_5344);
or U8643 (N_8643,N_6520,N_5190);
nand U8644 (N_8644,N_5084,N_6763);
nor U8645 (N_8645,N_5352,N_7158);
nand U8646 (N_8646,N_5113,N_6510);
and U8647 (N_8647,N_6794,N_5602);
nand U8648 (N_8648,N_6247,N_5458);
and U8649 (N_8649,N_5363,N_5626);
and U8650 (N_8650,N_5593,N_6511);
nor U8651 (N_8651,N_6274,N_6862);
or U8652 (N_8652,N_7179,N_6462);
nand U8653 (N_8653,N_5200,N_5495);
nor U8654 (N_8654,N_6549,N_5705);
nor U8655 (N_8655,N_5546,N_7021);
and U8656 (N_8656,N_5706,N_6866);
nand U8657 (N_8657,N_5482,N_6512);
xnor U8658 (N_8658,N_5635,N_5784);
or U8659 (N_8659,N_6432,N_7250);
and U8660 (N_8660,N_7062,N_5327);
nor U8661 (N_8661,N_6854,N_5158);
or U8662 (N_8662,N_5162,N_6067);
and U8663 (N_8663,N_5282,N_6573);
or U8664 (N_8664,N_7300,N_5149);
or U8665 (N_8665,N_5716,N_7278);
and U8666 (N_8666,N_6218,N_6017);
or U8667 (N_8667,N_5663,N_7019);
nand U8668 (N_8668,N_6146,N_5633);
and U8669 (N_8669,N_5334,N_5452);
or U8670 (N_8670,N_5849,N_6121);
and U8671 (N_8671,N_6458,N_5271);
nand U8672 (N_8672,N_6187,N_5717);
and U8673 (N_8673,N_5712,N_5024);
or U8674 (N_8674,N_6937,N_5726);
and U8675 (N_8675,N_5419,N_6701);
or U8676 (N_8676,N_7174,N_6140);
nand U8677 (N_8677,N_5763,N_7248);
and U8678 (N_8678,N_6881,N_5884);
nand U8679 (N_8679,N_6771,N_5977);
nand U8680 (N_8680,N_5935,N_7071);
nor U8681 (N_8681,N_5511,N_6198);
and U8682 (N_8682,N_5765,N_6249);
nor U8683 (N_8683,N_7183,N_6211);
nand U8684 (N_8684,N_6150,N_5434);
nand U8685 (N_8685,N_5788,N_6385);
or U8686 (N_8686,N_6838,N_5411);
nand U8687 (N_8687,N_6897,N_6956);
and U8688 (N_8688,N_5206,N_5247);
nor U8689 (N_8689,N_6554,N_6457);
or U8690 (N_8690,N_7439,N_6938);
nand U8691 (N_8691,N_6034,N_5489);
or U8692 (N_8692,N_5657,N_7170);
nand U8693 (N_8693,N_6704,N_7334);
nor U8694 (N_8694,N_6386,N_5539);
or U8695 (N_8695,N_6934,N_5333);
or U8696 (N_8696,N_7493,N_5698);
xor U8697 (N_8697,N_6220,N_6243);
nor U8698 (N_8698,N_7440,N_7288);
nor U8699 (N_8699,N_6578,N_5338);
and U8700 (N_8700,N_6072,N_5183);
and U8701 (N_8701,N_6548,N_6111);
nand U8702 (N_8702,N_6068,N_5093);
xnor U8703 (N_8703,N_6231,N_5117);
nand U8704 (N_8704,N_6378,N_7217);
nor U8705 (N_8705,N_7340,N_7424);
and U8706 (N_8706,N_6601,N_5012);
nand U8707 (N_8707,N_5725,N_7129);
nand U8708 (N_8708,N_6298,N_6884);
nor U8709 (N_8709,N_6278,N_5060);
nor U8710 (N_8710,N_7294,N_6176);
nand U8711 (N_8711,N_7428,N_7437);
and U8712 (N_8712,N_6604,N_6501);
and U8713 (N_8713,N_5336,N_6728);
nor U8714 (N_8714,N_6179,N_7355);
nor U8715 (N_8715,N_6383,N_6014);
nand U8716 (N_8716,N_5353,N_7331);
nor U8717 (N_8717,N_5924,N_6040);
or U8718 (N_8718,N_6743,N_5256);
nor U8719 (N_8719,N_7399,N_7208);
nor U8720 (N_8720,N_6490,N_6738);
or U8721 (N_8721,N_6113,N_6565);
and U8722 (N_8722,N_5085,N_5611);
nor U8723 (N_8723,N_6840,N_7234);
nand U8724 (N_8724,N_6997,N_6568);
nand U8725 (N_8725,N_6695,N_7086);
and U8726 (N_8726,N_6612,N_6133);
nand U8727 (N_8727,N_6444,N_5254);
or U8728 (N_8728,N_5174,N_7324);
and U8729 (N_8729,N_6776,N_5889);
nand U8730 (N_8730,N_6431,N_6557);
nand U8731 (N_8731,N_5843,N_7167);
nand U8732 (N_8732,N_5544,N_6212);
nand U8733 (N_8733,N_6452,N_6555);
xor U8734 (N_8734,N_5456,N_5354);
and U8735 (N_8735,N_7356,N_7059);
or U8736 (N_8736,N_6475,N_6500);
or U8737 (N_8737,N_5406,N_6882);
and U8738 (N_8738,N_6835,N_5058);
and U8739 (N_8739,N_7362,N_7247);
nor U8740 (N_8740,N_6061,N_6269);
nand U8741 (N_8741,N_7360,N_6855);
or U8742 (N_8742,N_5227,N_5953);
or U8743 (N_8743,N_5964,N_7011);
nor U8744 (N_8744,N_7007,N_5700);
and U8745 (N_8745,N_7156,N_6318);
and U8746 (N_8746,N_6558,N_6419);
nand U8747 (N_8747,N_7054,N_5437);
and U8748 (N_8748,N_5361,N_5376);
and U8749 (N_8749,N_5182,N_6727);
nand U8750 (N_8750,N_5248,N_6424);
nor U8751 (N_8751,N_6375,N_6722);
nor U8752 (N_8752,N_5338,N_5447);
nand U8753 (N_8753,N_7118,N_5428);
nor U8754 (N_8754,N_5068,N_5768);
or U8755 (N_8755,N_5479,N_6391);
and U8756 (N_8756,N_5010,N_5529);
nand U8757 (N_8757,N_7114,N_7300);
or U8758 (N_8758,N_6533,N_7379);
and U8759 (N_8759,N_5646,N_5245);
or U8760 (N_8760,N_7254,N_6494);
and U8761 (N_8761,N_5999,N_5091);
and U8762 (N_8762,N_7085,N_5173);
or U8763 (N_8763,N_6301,N_7358);
nand U8764 (N_8764,N_6342,N_6444);
nor U8765 (N_8765,N_5980,N_6844);
nor U8766 (N_8766,N_6295,N_5859);
or U8767 (N_8767,N_7437,N_5164);
and U8768 (N_8768,N_5361,N_5760);
nand U8769 (N_8769,N_5531,N_5259);
nand U8770 (N_8770,N_6134,N_7233);
or U8771 (N_8771,N_5105,N_6111);
and U8772 (N_8772,N_6898,N_5312);
nand U8773 (N_8773,N_6454,N_6731);
nand U8774 (N_8774,N_6740,N_5812);
or U8775 (N_8775,N_6700,N_5729);
or U8776 (N_8776,N_6322,N_7033);
and U8777 (N_8777,N_7448,N_7072);
nor U8778 (N_8778,N_7470,N_6259);
or U8779 (N_8779,N_6790,N_5708);
nand U8780 (N_8780,N_5956,N_6268);
nor U8781 (N_8781,N_7235,N_5655);
nor U8782 (N_8782,N_6504,N_6003);
nor U8783 (N_8783,N_7031,N_6916);
or U8784 (N_8784,N_7057,N_7412);
and U8785 (N_8785,N_5474,N_5218);
or U8786 (N_8786,N_5164,N_7404);
nor U8787 (N_8787,N_6332,N_6995);
nor U8788 (N_8788,N_6806,N_6661);
nand U8789 (N_8789,N_5715,N_6233);
nor U8790 (N_8790,N_5108,N_5150);
or U8791 (N_8791,N_5574,N_6374);
and U8792 (N_8792,N_6195,N_5637);
nand U8793 (N_8793,N_5385,N_6253);
nand U8794 (N_8794,N_5324,N_7159);
and U8795 (N_8795,N_7054,N_6012);
or U8796 (N_8796,N_5219,N_6829);
and U8797 (N_8797,N_7153,N_6405);
and U8798 (N_8798,N_6117,N_6137);
and U8799 (N_8799,N_5553,N_6222);
nor U8800 (N_8800,N_6013,N_5612);
nand U8801 (N_8801,N_5699,N_7106);
nor U8802 (N_8802,N_5801,N_6066);
or U8803 (N_8803,N_7241,N_7034);
nand U8804 (N_8804,N_6763,N_6812);
or U8805 (N_8805,N_7406,N_7026);
nor U8806 (N_8806,N_5005,N_5008);
nor U8807 (N_8807,N_5479,N_7349);
nor U8808 (N_8808,N_7114,N_5134);
nand U8809 (N_8809,N_5753,N_5732);
and U8810 (N_8810,N_6002,N_7210);
or U8811 (N_8811,N_5862,N_5626);
or U8812 (N_8812,N_5744,N_6480);
nor U8813 (N_8813,N_5980,N_7113);
nor U8814 (N_8814,N_7024,N_7410);
nand U8815 (N_8815,N_5387,N_5678);
nand U8816 (N_8816,N_6186,N_7333);
and U8817 (N_8817,N_5208,N_5326);
or U8818 (N_8818,N_7325,N_7458);
and U8819 (N_8819,N_6304,N_6698);
or U8820 (N_8820,N_6323,N_6246);
nor U8821 (N_8821,N_7119,N_7264);
and U8822 (N_8822,N_5082,N_6790);
or U8823 (N_8823,N_5454,N_6040);
nand U8824 (N_8824,N_6104,N_7449);
or U8825 (N_8825,N_6710,N_5422);
nor U8826 (N_8826,N_5411,N_7258);
or U8827 (N_8827,N_6237,N_6001);
or U8828 (N_8828,N_6213,N_6472);
nand U8829 (N_8829,N_7293,N_6106);
nand U8830 (N_8830,N_6319,N_6021);
nor U8831 (N_8831,N_5741,N_5045);
and U8832 (N_8832,N_7380,N_6016);
or U8833 (N_8833,N_6056,N_5216);
or U8834 (N_8834,N_6367,N_6224);
and U8835 (N_8835,N_5931,N_6190);
and U8836 (N_8836,N_6759,N_6728);
nand U8837 (N_8837,N_5449,N_5897);
nand U8838 (N_8838,N_6115,N_5289);
nand U8839 (N_8839,N_6214,N_5659);
nand U8840 (N_8840,N_6838,N_5933);
nand U8841 (N_8841,N_5971,N_6409);
and U8842 (N_8842,N_6849,N_6949);
nor U8843 (N_8843,N_6189,N_5812);
nor U8844 (N_8844,N_5579,N_7320);
or U8845 (N_8845,N_6226,N_7092);
nand U8846 (N_8846,N_5540,N_6629);
or U8847 (N_8847,N_5488,N_6970);
or U8848 (N_8848,N_7367,N_6171);
xnor U8849 (N_8849,N_7040,N_6300);
or U8850 (N_8850,N_5319,N_6488);
nand U8851 (N_8851,N_7102,N_5387);
nor U8852 (N_8852,N_5821,N_6753);
or U8853 (N_8853,N_7306,N_5153);
nor U8854 (N_8854,N_6087,N_5991);
nor U8855 (N_8855,N_5377,N_5952);
nor U8856 (N_8856,N_5937,N_6449);
or U8857 (N_8857,N_6411,N_5716);
and U8858 (N_8858,N_6323,N_6178);
nor U8859 (N_8859,N_5301,N_5074);
and U8860 (N_8860,N_7018,N_5449);
nor U8861 (N_8861,N_7162,N_5663);
nor U8862 (N_8862,N_7050,N_6877);
and U8863 (N_8863,N_5703,N_5630);
nand U8864 (N_8864,N_6396,N_6617);
nand U8865 (N_8865,N_5805,N_7205);
and U8866 (N_8866,N_5104,N_7053);
nand U8867 (N_8867,N_5134,N_5627);
and U8868 (N_8868,N_6307,N_7460);
nor U8869 (N_8869,N_5455,N_5992);
and U8870 (N_8870,N_5509,N_6971);
nand U8871 (N_8871,N_5913,N_5730);
nor U8872 (N_8872,N_6301,N_7086);
nand U8873 (N_8873,N_5992,N_6034);
or U8874 (N_8874,N_6906,N_6661);
or U8875 (N_8875,N_5562,N_5526);
nand U8876 (N_8876,N_5739,N_5467);
nand U8877 (N_8877,N_7078,N_5234);
nor U8878 (N_8878,N_6662,N_5505);
nand U8879 (N_8879,N_5725,N_5716);
nor U8880 (N_8880,N_6506,N_5576);
nor U8881 (N_8881,N_5452,N_6222);
nand U8882 (N_8882,N_5381,N_5585);
and U8883 (N_8883,N_7172,N_5987);
nor U8884 (N_8884,N_5455,N_5395);
nand U8885 (N_8885,N_7175,N_6488);
or U8886 (N_8886,N_5000,N_6301);
nor U8887 (N_8887,N_6323,N_5790);
nor U8888 (N_8888,N_5430,N_5898);
or U8889 (N_8889,N_6862,N_7380);
and U8890 (N_8890,N_6892,N_5122);
or U8891 (N_8891,N_6765,N_5499);
and U8892 (N_8892,N_5191,N_5838);
nor U8893 (N_8893,N_5886,N_7322);
nor U8894 (N_8894,N_6455,N_6960);
nand U8895 (N_8895,N_5257,N_7206);
or U8896 (N_8896,N_7109,N_6461);
or U8897 (N_8897,N_5861,N_5634);
or U8898 (N_8898,N_5925,N_6300);
or U8899 (N_8899,N_5347,N_7173);
nand U8900 (N_8900,N_7251,N_7041);
nor U8901 (N_8901,N_6275,N_7339);
nand U8902 (N_8902,N_5276,N_5459);
nor U8903 (N_8903,N_5607,N_6961);
or U8904 (N_8904,N_7224,N_6669);
and U8905 (N_8905,N_6015,N_5147);
nand U8906 (N_8906,N_6465,N_6834);
and U8907 (N_8907,N_5712,N_6747);
or U8908 (N_8908,N_5279,N_7422);
or U8909 (N_8909,N_5760,N_7180);
or U8910 (N_8910,N_6065,N_6416);
and U8911 (N_8911,N_7034,N_6318);
or U8912 (N_8912,N_5968,N_5361);
and U8913 (N_8913,N_6424,N_5833);
nand U8914 (N_8914,N_5454,N_7271);
nand U8915 (N_8915,N_5477,N_6720);
or U8916 (N_8916,N_5722,N_6252);
or U8917 (N_8917,N_5624,N_5260);
nand U8918 (N_8918,N_6320,N_5591);
nor U8919 (N_8919,N_6073,N_5670);
or U8920 (N_8920,N_7339,N_5794);
and U8921 (N_8921,N_5083,N_7012);
nand U8922 (N_8922,N_7034,N_5215);
nor U8923 (N_8923,N_7333,N_6285);
or U8924 (N_8924,N_6023,N_6639);
or U8925 (N_8925,N_7265,N_6078);
and U8926 (N_8926,N_5707,N_7374);
and U8927 (N_8927,N_5836,N_6244);
nor U8928 (N_8928,N_6017,N_5066);
or U8929 (N_8929,N_6020,N_5039);
nor U8930 (N_8930,N_6623,N_6106);
nor U8931 (N_8931,N_7417,N_5006);
and U8932 (N_8932,N_5724,N_5441);
nand U8933 (N_8933,N_7023,N_5485);
xor U8934 (N_8934,N_6609,N_7423);
and U8935 (N_8935,N_7033,N_7106);
nand U8936 (N_8936,N_5359,N_5354);
nand U8937 (N_8937,N_5984,N_7135);
nand U8938 (N_8938,N_7390,N_5555);
or U8939 (N_8939,N_6320,N_6635);
or U8940 (N_8940,N_7239,N_6368);
or U8941 (N_8941,N_5667,N_5528);
or U8942 (N_8942,N_7158,N_7153);
and U8943 (N_8943,N_6057,N_5827);
nand U8944 (N_8944,N_6590,N_5805);
and U8945 (N_8945,N_6306,N_6788);
and U8946 (N_8946,N_7137,N_5751);
nand U8947 (N_8947,N_6638,N_5171);
nor U8948 (N_8948,N_6854,N_6559);
and U8949 (N_8949,N_6721,N_7121);
nor U8950 (N_8950,N_6015,N_5389);
nand U8951 (N_8951,N_7158,N_5699);
and U8952 (N_8952,N_6612,N_6293);
or U8953 (N_8953,N_6343,N_7100);
or U8954 (N_8954,N_6016,N_5109);
nor U8955 (N_8955,N_6245,N_7265);
or U8956 (N_8956,N_6652,N_5586);
nor U8957 (N_8957,N_5859,N_5522);
xor U8958 (N_8958,N_7413,N_6189);
or U8959 (N_8959,N_6782,N_5670);
nor U8960 (N_8960,N_5508,N_5292);
or U8961 (N_8961,N_5732,N_5543);
or U8962 (N_8962,N_7490,N_6222);
and U8963 (N_8963,N_7196,N_6561);
nor U8964 (N_8964,N_5929,N_7345);
nor U8965 (N_8965,N_7371,N_6058);
nor U8966 (N_8966,N_6811,N_7140);
or U8967 (N_8967,N_6834,N_6668);
or U8968 (N_8968,N_5848,N_6579);
and U8969 (N_8969,N_5737,N_6850);
and U8970 (N_8970,N_5473,N_5064);
nor U8971 (N_8971,N_7329,N_6914);
and U8972 (N_8972,N_5512,N_7172);
nor U8973 (N_8973,N_5890,N_5810);
nand U8974 (N_8974,N_6562,N_7259);
nor U8975 (N_8975,N_5549,N_5225);
nand U8976 (N_8976,N_7476,N_5720);
nand U8977 (N_8977,N_7091,N_7380);
and U8978 (N_8978,N_5042,N_5656);
nor U8979 (N_8979,N_5592,N_6120);
and U8980 (N_8980,N_5143,N_5437);
nand U8981 (N_8981,N_7293,N_5997);
and U8982 (N_8982,N_6230,N_5321);
or U8983 (N_8983,N_5837,N_6480);
nor U8984 (N_8984,N_6385,N_5317);
and U8985 (N_8985,N_5103,N_7046);
nor U8986 (N_8986,N_6824,N_5308);
or U8987 (N_8987,N_6883,N_6494);
nand U8988 (N_8988,N_7024,N_7084);
xnor U8989 (N_8989,N_5562,N_5550);
and U8990 (N_8990,N_6028,N_6517);
nand U8991 (N_8991,N_6210,N_6283);
and U8992 (N_8992,N_7061,N_7408);
nor U8993 (N_8993,N_6806,N_6847);
nor U8994 (N_8994,N_6746,N_5997);
nor U8995 (N_8995,N_5374,N_5334);
or U8996 (N_8996,N_5134,N_6177);
nand U8997 (N_8997,N_7082,N_6131);
nand U8998 (N_8998,N_6269,N_6980);
nor U8999 (N_8999,N_6466,N_7238);
or U9000 (N_9000,N_5259,N_6106);
and U9001 (N_9001,N_6377,N_6676);
or U9002 (N_9002,N_6397,N_5103);
and U9003 (N_9003,N_6045,N_6645);
and U9004 (N_9004,N_5928,N_5833);
nor U9005 (N_9005,N_6881,N_5284);
and U9006 (N_9006,N_7486,N_5521);
nor U9007 (N_9007,N_6238,N_5011);
and U9008 (N_9008,N_5120,N_5806);
nand U9009 (N_9009,N_5640,N_6525);
and U9010 (N_9010,N_6528,N_6632);
nor U9011 (N_9011,N_5053,N_5486);
and U9012 (N_9012,N_7286,N_5916);
nor U9013 (N_9013,N_6850,N_5841);
nor U9014 (N_9014,N_6108,N_6503);
xor U9015 (N_9015,N_6364,N_6757);
or U9016 (N_9016,N_6382,N_5950);
nand U9017 (N_9017,N_7402,N_6851);
or U9018 (N_9018,N_6414,N_7388);
or U9019 (N_9019,N_6858,N_5987);
nor U9020 (N_9020,N_5864,N_6901);
nand U9021 (N_9021,N_6924,N_5514);
nor U9022 (N_9022,N_7242,N_7259);
nand U9023 (N_9023,N_6312,N_5390);
nor U9024 (N_9024,N_6388,N_6958);
nand U9025 (N_9025,N_6450,N_7389);
or U9026 (N_9026,N_6113,N_5273);
or U9027 (N_9027,N_6653,N_6341);
nor U9028 (N_9028,N_7205,N_6774);
nor U9029 (N_9029,N_5707,N_5859);
and U9030 (N_9030,N_7064,N_6758);
nand U9031 (N_9031,N_6586,N_6333);
nand U9032 (N_9032,N_6924,N_5007);
nor U9033 (N_9033,N_6572,N_5370);
nand U9034 (N_9034,N_6619,N_7038);
xor U9035 (N_9035,N_6242,N_5086);
nor U9036 (N_9036,N_6384,N_5812);
or U9037 (N_9037,N_5473,N_5264);
nand U9038 (N_9038,N_6595,N_6610);
or U9039 (N_9039,N_6758,N_5811);
nor U9040 (N_9040,N_5668,N_6726);
nand U9041 (N_9041,N_6914,N_5030);
and U9042 (N_9042,N_6226,N_5840);
or U9043 (N_9043,N_5113,N_5261);
and U9044 (N_9044,N_7399,N_5672);
or U9045 (N_9045,N_6443,N_5480);
nor U9046 (N_9046,N_6878,N_7012);
and U9047 (N_9047,N_5348,N_6749);
nor U9048 (N_9048,N_7028,N_7199);
nor U9049 (N_9049,N_5890,N_7155);
and U9050 (N_9050,N_7485,N_6164);
and U9051 (N_9051,N_5271,N_7097);
or U9052 (N_9052,N_6817,N_7435);
and U9053 (N_9053,N_5324,N_6080);
nor U9054 (N_9054,N_5241,N_5756);
nand U9055 (N_9055,N_7122,N_7293);
nand U9056 (N_9056,N_5637,N_6061);
or U9057 (N_9057,N_7118,N_5878);
nor U9058 (N_9058,N_5327,N_5020);
nor U9059 (N_9059,N_6771,N_6601);
and U9060 (N_9060,N_6728,N_5713);
xnor U9061 (N_9061,N_5843,N_5522);
and U9062 (N_9062,N_6524,N_5081);
nand U9063 (N_9063,N_5156,N_5527);
nand U9064 (N_9064,N_5530,N_5249);
or U9065 (N_9065,N_5628,N_6328);
and U9066 (N_9066,N_6584,N_5433);
or U9067 (N_9067,N_5725,N_7294);
nand U9068 (N_9068,N_7094,N_5482);
nand U9069 (N_9069,N_5728,N_7110);
or U9070 (N_9070,N_5197,N_6489);
nor U9071 (N_9071,N_7414,N_6527);
nor U9072 (N_9072,N_6158,N_7468);
nand U9073 (N_9073,N_6810,N_7298);
and U9074 (N_9074,N_7224,N_6812);
nor U9075 (N_9075,N_7062,N_6096);
or U9076 (N_9076,N_5913,N_6820);
nand U9077 (N_9077,N_6882,N_6597);
and U9078 (N_9078,N_7245,N_5927);
nor U9079 (N_9079,N_6080,N_7105);
or U9080 (N_9080,N_6019,N_6708);
or U9081 (N_9081,N_5895,N_6941);
nand U9082 (N_9082,N_6994,N_5941);
or U9083 (N_9083,N_5002,N_6030);
and U9084 (N_9084,N_5196,N_6889);
nor U9085 (N_9085,N_5522,N_5744);
or U9086 (N_9086,N_6514,N_5337);
and U9087 (N_9087,N_7107,N_5937);
or U9088 (N_9088,N_6255,N_6319);
nand U9089 (N_9089,N_7087,N_6094);
and U9090 (N_9090,N_7345,N_7448);
nor U9091 (N_9091,N_6677,N_6579);
nand U9092 (N_9092,N_5357,N_5584);
and U9093 (N_9093,N_5424,N_6068);
xor U9094 (N_9094,N_6697,N_5576);
nand U9095 (N_9095,N_6593,N_6611);
nand U9096 (N_9096,N_6403,N_7014);
nand U9097 (N_9097,N_6409,N_5855);
or U9098 (N_9098,N_7376,N_5426);
nand U9099 (N_9099,N_7203,N_6534);
xor U9100 (N_9100,N_6868,N_6089);
and U9101 (N_9101,N_7000,N_7412);
and U9102 (N_9102,N_5365,N_6161);
or U9103 (N_9103,N_5215,N_5592);
nor U9104 (N_9104,N_5703,N_5490);
nand U9105 (N_9105,N_6310,N_7226);
nor U9106 (N_9106,N_6713,N_5852);
or U9107 (N_9107,N_5888,N_6368);
nor U9108 (N_9108,N_6641,N_5616);
or U9109 (N_9109,N_5126,N_5860);
nand U9110 (N_9110,N_5537,N_6420);
or U9111 (N_9111,N_6368,N_6320);
or U9112 (N_9112,N_7331,N_7409);
nor U9113 (N_9113,N_6324,N_6380);
and U9114 (N_9114,N_6205,N_7072);
and U9115 (N_9115,N_6662,N_5420);
nor U9116 (N_9116,N_5863,N_5614);
nor U9117 (N_9117,N_6193,N_5572);
nand U9118 (N_9118,N_5634,N_7344);
nor U9119 (N_9119,N_6047,N_6962);
or U9120 (N_9120,N_7272,N_6324);
nor U9121 (N_9121,N_6143,N_6477);
or U9122 (N_9122,N_5327,N_5964);
or U9123 (N_9123,N_5865,N_5015);
nand U9124 (N_9124,N_5802,N_6713);
or U9125 (N_9125,N_6652,N_6225);
nand U9126 (N_9126,N_5982,N_7204);
and U9127 (N_9127,N_5758,N_7059);
nor U9128 (N_9128,N_7182,N_6875);
or U9129 (N_9129,N_6881,N_6927);
or U9130 (N_9130,N_6402,N_5861);
nor U9131 (N_9131,N_7204,N_5926);
and U9132 (N_9132,N_5946,N_6332);
and U9133 (N_9133,N_5549,N_6368);
nor U9134 (N_9134,N_6307,N_6213);
nor U9135 (N_9135,N_6451,N_5890);
and U9136 (N_9136,N_5881,N_5115);
nand U9137 (N_9137,N_5931,N_7235);
and U9138 (N_9138,N_5189,N_6124);
nand U9139 (N_9139,N_6601,N_5811);
nand U9140 (N_9140,N_6969,N_6675);
or U9141 (N_9141,N_6081,N_5203);
or U9142 (N_9142,N_5451,N_7343);
nor U9143 (N_9143,N_5956,N_6239);
or U9144 (N_9144,N_6414,N_6601);
nor U9145 (N_9145,N_5960,N_7093);
nand U9146 (N_9146,N_7337,N_5031);
or U9147 (N_9147,N_5456,N_5804);
or U9148 (N_9148,N_6077,N_6224);
nand U9149 (N_9149,N_6438,N_5537);
nand U9150 (N_9150,N_6162,N_5764);
nand U9151 (N_9151,N_7388,N_7116);
nand U9152 (N_9152,N_6208,N_5124);
or U9153 (N_9153,N_5562,N_5796);
and U9154 (N_9154,N_5373,N_6622);
and U9155 (N_9155,N_6001,N_5203);
nor U9156 (N_9156,N_6443,N_6428);
and U9157 (N_9157,N_7027,N_5945);
nor U9158 (N_9158,N_6247,N_5376);
nand U9159 (N_9159,N_7392,N_6138);
nand U9160 (N_9160,N_6922,N_6103);
and U9161 (N_9161,N_7172,N_6531);
nand U9162 (N_9162,N_5548,N_6350);
nor U9163 (N_9163,N_5544,N_6214);
nor U9164 (N_9164,N_7414,N_5618);
nand U9165 (N_9165,N_6877,N_6526);
or U9166 (N_9166,N_7067,N_5650);
and U9167 (N_9167,N_5466,N_5893);
or U9168 (N_9168,N_6288,N_5348);
or U9169 (N_9169,N_5395,N_5564);
or U9170 (N_9170,N_5841,N_6050);
and U9171 (N_9171,N_6193,N_7394);
nor U9172 (N_9172,N_7063,N_6764);
or U9173 (N_9173,N_6763,N_6801);
nand U9174 (N_9174,N_5471,N_5947);
nor U9175 (N_9175,N_7476,N_7157);
or U9176 (N_9176,N_6665,N_5617);
and U9177 (N_9177,N_5922,N_7218);
nand U9178 (N_9178,N_6838,N_7419);
and U9179 (N_9179,N_6355,N_6019);
nor U9180 (N_9180,N_7002,N_6710);
nand U9181 (N_9181,N_7286,N_5046);
or U9182 (N_9182,N_6617,N_6057);
or U9183 (N_9183,N_6582,N_6114);
nor U9184 (N_9184,N_7292,N_7378);
or U9185 (N_9185,N_7411,N_5061);
or U9186 (N_9186,N_6939,N_5972);
and U9187 (N_9187,N_5838,N_5664);
nor U9188 (N_9188,N_6893,N_7150);
nand U9189 (N_9189,N_5656,N_6978);
nor U9190 (N_9190,N_5789,N_5417);
nor U9191 (N_9191,N_6369,N_5501);
or U9192 (N_9192,N_7499,N_7123);
nand U9193 (N_9193,N_6951,N_7069);
and U9194 (N_9194,N_6109,N_6992);
or U9195 (N_9195,N_7031,N_6911);
and U9196 (N_9196,N_7055,N_6970);
nor U9197 (N_9197,N_5496,N_5294);
nor U9198 (N_9198,N_6099,N_5849);
nor U9199 (N_9199,N_5634,N_6183);
nor U9200 (N_9200,N_5906,N_5819);
and U9201 (N_9201,N_6731,N_7409);
nand U9202 (N_9202,N_6242,N_7186);
and U9203 (N_9203,N_6599,N_6341);
or U9204 (N_9204,N_7308,N_7140);
nand U9205 (N_9205,N_6253,N_5955);
and U9206 (N_9206,N_5519,N_5932);
and U9207 (N_9207,N_5118,N_6609);
nor U9208 (N_9208,N_5071,N_5984);
xnor U9209 (N_9209,N_6679,N_7191);
and U9210 (N_9210,N_5343,N_6064);
nand U9211 (N_9211,N_6104,N_7455);
or U9212 (N_9212,N_6813,N_6827);
or U9213 (N_9213,N_6349,N_6286);
or U9214 (N_9214,N_6990,N_6809);
nor U9215 (N_9215,N_6950,N_6187);
nand U9216 (N_9216,N_5691,N_6993);
and U9217 (N_9217,N_6981,N_7325);
nor U9218 (N_9218,N_5991,N_5854);
nor U9219 (N_9219,N_6867,N_5480);
nor U9220 (N_9220,N_7256,N_5085);
or U9221 (N_9221,N_7470,N_7220);
or U9222 (N_9222,N_5010,N_6151);
nand U9223 (N_9223,N_7051,N_6601);
nand U9224 (N_9224,N_5695,N_6231);
nand U9225 (N_9225,N_5379,N_6492);
and U9226 (N_9226,N_6062,N_6273);
and U9227 (N_9227,N_7410,N_5448);
nor U9228 (N_9228,N_6373,N_5367);
nand U9229 (N_9229,N_5253,N_5421);
or U9230 (N_9230,N_5163,N_6907);
nor U9231 (N_9231,N_6392,N_6972);
nor U9232 (N_9232,N_6778,N_5562);
nor U9233 (N_9233,N_6012,N_6112);
nand U9234 (N_9234,N_6157,N_6278);
nand U9235 (N_9235,N_6322,N_7250);
nor U9236 (N_9236,N_5870,N_6507);
nor U9237 (N_9237,N_7128,N_5685);
and U9238 (N_9238,N_7206,N_6573);
and U9239 (N_9239,N_6326,N_6444);
nand U9240 (N_9240,N_6875,N_6613);
nand U9241 (N_9241,N_7013,N_5808);
nor U9242 (N_9242,N_5560,N_6614);
and U9243 (N_9243,N_7059,N_7280);
nand U9244 (N_9244,N_6531,N_6581);
nand U9245 (N_9245,N_7202,N_5207);
nand U9246 (N_9246,N_6976,N_7428);
nor U9247 (N_9247,N_7240,N_7113);
nand U9248 (N_9248,N_5409,N_5008);
nand U9249 (N_9249,N_6638,N_6244);
or U9250 (N_9250,N_6855,N_7067);
nand U9251 (N_9251,N_5694,N_5531);
nor U9252 (N_9252,N_5156,N_6336);
and U9253 (N_9253,N_6130,N_7395);
nor U9254 (N_9254,N_5487,N_5125);
nor U9255 (N_9255,N_6350,N_5879);
and U9256 (N_9256,N_5054,N_7285);
and U9257 (N_9257,N_5982,N_7245);
nand U9258 (N_9258,N_5269,N_5313);
nand U9259 (N_9259,N_6296,N_5884);
and U9260 (N_9260,N_7316,N_7088);
and U9261 (N_9261,N_6457,N_5912);
or U9262 (N_9262,N_6171,N_6324);
nand U9263 (N_9263,N_5024,N_6842);
nor U9264 (N_9264,N_5769,N_6972);
and U9265 (N_9265,N_6691,N_5860);
and U9266 (N_9266,N_5276,N_5785);
or U9267 (N_9267,N_5062,N_5246);
or U9268 (N_9268,N_6957,N_6940);
nand U9269 (N_9269,N_7360,N_5313);
and U9270 (N_9270,N_7455,N_7410);
nor U9271 (N_9271,N_5553,N_5673);
nor U9272 (N_9272,N_5094,N_5882);
nand U9273 (N_9273,N_5193,N_5496);
nor U9274 (N_9274,N_6325,N_6127);
or U9275 (N_9275,N_5078,N_5463);
or U9276 (N_9276,N_6886,N_7161);
and U9277 (N_9277,N_6215,N_7149);
nor U9278 (N_9278,N_5563,N_5587);
nand U9279 (N_9279,N_6565,N_5121);
nand U9280 (N_9280,N_5459,N_5311);
nor U9281 (N_9281,N_5206,N_7281);
and U9282 (N_9282,N_6112,N_5809);
nor U9283 (N_9283,N_5013,N_6644);
nand U9284 (N_9284,N_5901,N_6608);
nand U9285 (N_9285,N_5547,N_5391);
nor U9286 (N_9286,N_7237,N_6174);
or U9287 (N_9287,N_6568,N_5831);
nor U9288 (N_9288,N_5001,N_6286);
or U9289 (N_9289,N_5339,N_6942);
nand U9290 (N_9290,N_6612,N_5317);
nand U9291 (N_9291,N_7319,N_5628);
and U9292 (N_9292,N_5427,N_7063);
nand U9293 (N_9293,N_7260,N_5242);
or U9294 (N_9294,N_7481,N_5260);
nand U9295 (N_9295,N_7278,N_5237);
nand U9296 (N_9296,N_6493,N_6729);
and U9297 (N_9297,N_6628,N_5045);
and U9298 (N_9298,N_6652,N_5178);
nor U9299 (N_9299,N_6949,N_6595);
nand U9300 (N_9300,N_5295,N_5000);
or U9301 (N_9301,N_6962,N_6504);
nand U9302 (N_9302,N_5039,N_5179);
or U9303 (N_9303,N_6532,N_7247);
nor U9304 (N_9304,N_7087,N_6819);
and U9305 (N_9305,N_7038,N_5572);
nor U9306 (N_9306,N_6756,N_6000);
or U9307 (N_9307,N_5540,N_5366);
or U9308 (N_9308,N_7209,N_7206);
nor U9309 (N_9309,N_6086,N_5594);
nand U9310 (N_9310,N_6821,N_5720);
and U9311 (N_9311,N_5294,N_5269);
nand U9312 (N_9312,N_6502,N_5360);
and U9313 (N_9313,N_6745,N_6914);
nor U9314 (N_9314,N_6454,N_5935);
nor U9315 (N_9315,N_5628,N_5589);
xnor U9316 (N_9316,N_5991,N_7097);
and U9317 (N_9317,N_7253,N_5826);
nor U9318 (N_9318,N_5593,N_6740);
or U9319 (N_9319,N_5635,N_5174);
and U9320 (N_9320,N_5009,N_6795);
nand U9321 (N_9321,N_7353,N_6019);
nand U9322 (N_9322,N_5874,N_5406);
or U9323 (N_9323,N_5768,N_7472);
nand U9324 (N_9324,N_6343,N_5822);
or U9325 (N_9325,N_6616,N_6038);
nand U9326 (N_9326,N_5996,N_5706);
nor U9327 (N_9327,N_6768,N_5267);
or U9328 (N_9328,N_6733,N_6109);
nor U9329 (N_9329,N_6858,N_5866);
nor U9330 (N_9330,N_7275,N_6237);
nor U9331 (N_9331,N_7188,N_6944);
nor U9332 (N_9332,N_6569,N_5032);
nand U9333 (N_9333,N_7414,N_5485);
nor U9334 (N_9334,N_5417,N_5416);
and U9335 (N_9335,N_5201,N_5718);
nor U9336 (N_9336,N_6884,N_6125);
and U9337 (N_9337,N_7431,N_6977);
nand U9338 (N_9338,N_6022,N_6824);
nor U9339 (N_9339,N_7086,N_5248);
nand U9340 (N_9340,N_6234,N_6144);
nor U9341 (N_9341,N_6942,N_6487);
or U9342 (N_9342,N_5113,N_6995);
nor U9343 (N_9343,N_7020,N_5864);
nand U9344 (N_9344,N_7296,N_5040);
nor U9345 (N_9345,N_5035,N_5521);
nor U9346 (N_9346,N_6522,N_7080);
nand U9347 (N_9347,N_7463,N_6244);
or U9348 (N_9348,N_6513,N_6223);
and U9349 (N_9349,N_6077,N_5622);
and U9350 (N_9350,N_5797,N_7107);
nor U9351 (N_9351,N_7224,N_7139);
nand U9352 (N_9352,N_5552,N_5422);
or U9353 (N_9353,N_7189,N_6481);
nand U9354 (N_9354,N_7144,N_7441);
nor U9355 (N_9355,N_6867,N_5403);
or U9356 (N_9356,N_5991,N_7489);
nand U9357 (N_9357,N_7323,N_5810);
nor U9358 (N_9358,N_5135,N_6157);
nor U9359 (N_9359,N_5728,N_7013);
or U9360 (N_9360,N_6635,N_7212);
and U9361 (N_9361,N_6608,N_5088);
and U9362 (N_9362,N_5826,N_6776);
and U9363 (N_9363,N_5764,N_5713);
or U9364 (N_9364,N_6482,N_5895);
nor U9365 (N_9365,N_7472,N_6642);
nand U9366 (N_9366,N_5883,N_6925);
nor U9367 (N_9367,N_6795,N_6822);
or U9368 (N_9368,N_5091,N_6825);
nand U9369 (N_9369,N_5306,N_6953);
nor U9370 (N_9370,N_7279,N_6345);
nor U9371 (N_9371,N_5137,N_6132);
or U9372 (N_9372,N_7370,N_5269);
and U9373 (N_9373,N_6424,N_7294);
nor U9374 (N_9374,N_6389,N_6764);
nand U9375 (N_9375,N_6403,N_6085);
nand U9376 (N_9376,N_5538,N_5179);
nand U9377 (N_9377,N_6776,N_6897);
and U9378 (N_9378,N_6592,N_5773);
nand U9379 (N_9379,N_5229,N_6809);
nor U9380 (N_9380,N_6272,N_6578);
or U9381 (N_9381,N_6724,N_5818);
or U9382 (N_9382,N_5616,N_5758);
nor U9383 (N_9383,N_5225,N_7106);
and U9384 (N_9384,N_7286,N_6560);
nand U9385 (N_9385,N_5976,N_6012);
nor U9386 (N_9386,N_6433,N_7044);
nand U9387 (N_9387,N_5739,N_6122);
nand U9388 (N_9388,N_6740,N_5977);
nor U9389 (N_9389,N_5895,N_6123);
nor U9390 (N_9390,N_5579,N_5064);
nand U9391 (N_9391,N_5572,N_5757);
or U9392 (N_9392,N_7291,N_5909);
nand U9393 (N_9393,N_5860,N_5859);
nand U9394 (N_9394,N_6586,N_5856);
and U9395 (N_9395,N_6668,N_6656);
nand U9396 (N_9396,N_5708,N_6795);
nand U9397 (N_9397,N_5446,N_5462);
or U9398 (N_9398,N_5276,N_7486);
nor U9399 (N_9399,N_6417,N_6183);
nand U9400 (N_9400,N_5722,N_5423);
and U9401 (N_9401,N_6446,N_6153);
or U9402 (N_9402,N_7328,N_6003);
and U9403 (N_9403,N_5697,N_5700);
and U9404 (N_9404,N_7035,N_5497);
or U9405 (N_9405,N_6283,N_6628);
and U9406 (N_9406,N_5044,N_7272);
nor U9407 (N_9407,N_6266,N_6445);
nand U9408 (N_9408,N_5537,N_5320);
nor U9409 (N_9409,N_6698,N_5486);
nor U9410 (N_9410,N_5685,N_5712);
and U9411 (N_9411,N_6580,N_6914);
nor U9412 (N_9412,N_5140,N_5879);
or U9413 (N_9413,N_6395,N_6868);
and U9414 (N_9414,N_6182,N_5080);
and U9415 (N_9415,N_5512,N_6495);
nand U9416 (N_9416,N_5029,N_7499);
nand U9417 (N_9417,N_5744,N_6114);
nand U9418 (N_9418,N_7359,N_6531);
nand U9419 (N_9419,N_6595,N_6814);
xor U9420 (N_9420,N_5453,N_5913);
and U9421 (N_9421,N_6866,N_6709);
or U9422 (N_9422,N_5420,N_6328);
or U9423 (N_9423,N_7311,N_6744);
nand U9424 (N_9424,N_6097,N_6722);
and U9425 (N_9425,N_6500,N_6315);
or U9426 (N_9426,N_6660,N_5253);
and U9427 (N_9427,N_6561,N_5513);
nor U9428 (N_9428,N_5732,N_6164);
nand U9429 (N_9429,N_5995,N_6148);
and U9430 (N_9430,N_6728,N_6925);
nor U9431 (N_9431,N_5940,N_5040);
nor U9432 (N_9432,N_5383,N_6819);
nand U9433 (N_9433,N_5408,N_7092);
or U9434 (N_9434,N_6218,N_5256);
nand U9435 (N_9435,N_5684,N_7458);
and U9436 (N_9436,N_5324,N_6079);
and U9437 (N_9437,N_6232,N_6951);
nor U9438 (N_9438,N_6434,N_6170);
nor U9439 (N_9439,N_5767,N_6254);
nand U9440 (N_9440,N_6448,N_6589);
nor U9441 (N_9441,N_5545,N_6128);
nand U9442 (N_9442,N_5998,N_6542);
or U9443 (N_9443,N_5440,N_5706);
or U9444 (N_9444,N_7481,N_6828);
or U9445 (N_9445,N_5608,N_7393);
and U9446 (N_9446,N_6405,N_6315);
or U9447 (N_9447,N_5398,N_6914);
or U9448 (N_9448,N_7012,N_6286);
or U9449 (N_9449,N_5918,N_6014);
or U9450 (N_9450,N_5241,N_6630);
nor U9451 (N_9451,N_5417,N_6746);
or U9452 (N_9452,N_6367,N_6766);
and U9453 (N_9453,N_5877,N_5026);
or U9454 (N_9454,N_5402,N_5870);
and U9455 (N_9455,N_6865,N_5120);
and U9456 (N_9456,N_5826,N_6654);
nand U9457 (N_9457,N_6205,N_5588);
and U9458 (N_9458,N_7293,N_7368);
nand U9459 (N_9459,N_5406,N_5610);
nor U9460 (N_9460,N_7118,N_5595);
nor U9461 (N_9461,N_5311,N_5977);
and U9462 (N_9462,N_6876,N_7379);
nor U9463 (N_9463,N_6115,N_5051);
nand U9464 (N_9464,N_5979,N_6173);
and U9465 (N_9465,N_6639,N_6342);
nand U9466 (N_9466,N_6898,N_7407);
nor U9467 (N_9467,N_6397,N_5604);
nor U9468 (N_9468,N_6159,N_6837);
nor U9469 (N_9469,N_6845,N_5718);
and U9470 (N_9470,N_6514,N_6933);
nand U9471 (N_9471,N_5026,N_6678);
nor U9472 (N_9472,N_6948,N_7449);
and U9473 (N_9473,N_5793,N_5129);
nor U9474 (N_9474,N_5060,N_5907);
or U9475 (N_9475,N_6278,N_5297);
and U9476 (N_9476,N_7333,N_6423);
nand U9477 (N_9477,N_6154,N_6968);
nand U9478 (N_9478,N_5747,N_5262);
and U9479 (N_9479,N_5542,N_5849);
or U9480 (N_9480,N_6040,N_7400);
nor U9481 (N_9481,N_5946,N_6923);
nor U9482 (N_9482,N_5171,N_5495);
nand U9483 (N_9483,N_5000,N_6034);
and U9484 (N_9484,N_6095,N_5102);
nand U9485 (N_9485,N_6047,N_6422);
nor U9486 (N_9486,N_5778,N_5407);
nand U9487 (N_9487,N_5521,N_7089);
and U9488 (N_9488,N_7289,N_6101);
nor U9489 (N_9489,N_5176,N_6742);
and U9490 (N_9490,N_5977,N_6177);
and U9491 (N_9491,N_7390,N_5020);
nand U9492 (N_9492,N_6424,N_6471);
and U9493 (N_9493,N_5938,N_5385);
nor U9494 (N_9494,N_7325,N_7241);
and U9495 (N_9495,N_6422,N_5563);
or U9496 (N_9496,N_6810,N_6498);
nand U9497 (N_9497,N_5975,N_5217);
or U9498 (N_9498,N_7419,N_5716);
nand U9499 (N_9499,N_6495,N_5344);
and U9500 (N_9500,N_5479,N_5347);
nand U9501 (N_9501,N_6415,N_6742);
or U9502 (N_9502,N_6644,N_6057);
and U9503 (N_9503,N_5478,N_6623);
nand U9504 (N_9504,N_5664,N_7111);
nor U9505 (N_9505,N_5724,N_5654);
or U9506 (N_9506,N_5474,N_5266);
or U9507 (N_9507,N_5080,N_5428);
nand U9508 (N_9508,N_5026,N_5956);
and U9509 (N_9509,N_5188,N_7201);
and U9510 (N_9510,N_6974,N_5130);
and U9511 (N_9511,N_6458,N_5381);
or U9512 (N_9512,N_6309,N_6613);
or U9513 (N_9513,N_6978,N_5076);
or U9514 (N_9514,N_5867,N_5410);
nor U9515 (N_9515,N_7489,N_5973);
nand U9516 (N_9516,N_6892,N_7377);
or U9517 (N_9517,N_5063,N_6460);
nand U9518 (N_9518,N_6531,N_6510);
nand U9519 (N_9519,N_5352,N_5560);
or U9520 (N_9520,N_5009,N_5210);
or U9521 (N_9521,N_5199,N_6395);
nand U9522 (N_9522,N_7447,N_5978);
or U9523 (N_9523,N_6103,N_5242);
and U9524 (N_9524,N_5260,N_6647);
and U9525 (N_9525,N_6269,N_6009);
and U9526 (N_9526,N_5622,N_5251);
and U9527 (N_9527,N_6560,N_6578);
nand U9528 (N_9528,N_6689,N_5193);
or U9529 (N_9529,N_6163,N_5353);
nor U9530 (N_9530,N_5967,N_5783);
nor U9531 (N_9531,N_6228,N_5861);
nor U9532 (N_9532,N_5764,N_5555);
nand U9533 (N_9533,N_5648,N_6774);
nor U9534 (N_9534,N_5988,N_6366);
nor U9535 (N_9535,N_6386,N_6508);
and U9536 (N_9536,N_5548,N_5561);
nand U9537 (N_9537,N_5635,N_6227);
nor U9538 (N_9538,N_5722,N_5404);
and U9539 (N_9539,N_5545,N_7184);
or U9540 (N_9540,N_6687,N_6475);
and U9541 (N_9541,N_6094,N_7368);
nand U9542 (N_9542,N_7033,N_6331);
nor U9543 (N_9543,N_5699,N_5421);
and U9544 (N_9544,N_5755,N_6572);
nor U9545 (N_9545,N_5534,N_6810);
and U9546 (N_9546,N_5803,N_7429);
nand U9547 (N_9547,N_6097,N_6278);
or U9548 (N_9548,N_5613,N_7495);
nand U9549 (N_9549,N_6797,N_6320);
or U9550 (N_9550,N_7244,N_5777);
nor U9551 (N_9551,N_5230,N_6803);
and U9552 (N_9552,N_5462,N_6239);
and U9553 (N_9553,N_7100,N_5091);
nand U9554 (N_9554,N_7126,N_5981);
nand U9555 (N_9555,N_6361,N_5230);
nand U9556 (N_9556,N_6588,N_7213);
nand U9557 (N_9557,N_6792,N_7119);
and U9558 (N_9558,N_5913,N_6570);
and U9559 (N_9559,N_5781,N_6973);
nor U9560 (N_9560,N_7147,N_6125);
nand U9561 (N_9561,N_7065,N_7337);
or U9562 (N_9562,N_5248,N_5774);
nand U9563 (N_9563,N_5603,N_7166);
and U9564 (N_9564,N_7163,N_6725);
nor U9565 (N_9565,N_5908,N_5804);
nand U9566 (N_9566,N_5766,N_6102);
or U9567 (N_9567,N_5362,N_6186);
nor U9568 (N_9568,N_6568,N_7447);
xor U9569 (N_9569,N_5664,N_6416);
nor U9570 (N_9570,N_5337,N_7488);
or U9571 (N_9571,N_6525,N_6876);
nor U9572 (N_9572,N_6044,N_6710);
nand U9573 (N_9573,N_6445,N_5994);
nor U9574 (N_9574,N_6707,N_5273);
nand U9575 (N_9575,N_7077,N_7182);
and U9576 (N_9576,N_6668,N_5591);
and U9577 (N_9577,N_6152,N_5069);
or U9578 (N_9578,N_5019,N_6515);
nand U9579 (N_9579,N_6040,N_7463);
and U9580 (N_9580,N_6070,N_6948);
nand U9581 (N_9581,N_6002,N_5477);
nand U9582 (N_9582,N_5890,N_7370);
nor U9583 (N_9583,N_5526,N_6944);
and U9584 (N_9584,N_6198,N_5386);
nor U9585 (N_9585,N_5636,N_5664);
and U9586 (N_9586,N_5172,N_7246);
or U9587 (N_9587,N_6960,N_5117);
and U9588 (N_9588,N_5222,N_6690);
xor U9589 (N_9589,N_5664,N_5211);
nand U9590 (N_9590,N_6207,N_6757);
and U9591 (N_9591,N_6905,N_6418);
nand U9592 (N_9592,N_6609,N_5035);
and U9593 (N_9593,N_7227,N_6846);
nand U9594 (N_9594,N_6838,N_7458);
and U9595 (N_9595,N_6941,N_6877);
nand U9596 (N_9596,N_7094,N_5666);
or U9597 (N_9597,N_5695,N_7385);
nor U9598 (N_9598,N_5750,N_5713);
nand U9599 (N_9599,N_5115,N_5106);
nand U9600 (N_9600,N_5233,N_5635);
or U9601 (N_9601,N_6884,N_5393);
nand U9602 (N_9602,N_5815,N_6289);
nand U9603 (N_9603,N_7468,N_6076);
nand U9604 (N_9604,N_6984,N_5511);
or U9605 (N_9605,N_5473,N_7016);
nand U9606 (N_9606,N_6135,N_6694);
or U9607 (N_9607,N_7404,N_7344);
nand U9608 (N_9608,N_6136,N_6542);
nor U9609 (N_9609,N_7123,N_5418);
or U9610 (N_9610,N_6605,N_7321);
nand U9611 (N_9611,N_7458,N_7451);
or U9612 (N_9612,N_5726,N_7102);
nor U9613 (N_9613,N_5110,N_6358);
nor U9614 (N_9614,N_5786,N_5821);
and U9615 (N_9615,N_5289,N_7121);
or U9616 (N_9616,N_7200,N_5067);
nor U9617 (N_9617,N_6132,N_6689);
nand U9618 (N_9618,N_5869,N_6815);
nor U9619 (N_9619,N_5549,N_6100);
nor U9620 (N_9620,N_6018,N_6182);
and U9621 (N_9621,N_6481,N_6981);
or U9622 (N_9622,N_6538,N_5342);
nand U9623 (N_9623,N_5848,N_7184);
nand U9624 (N_9624,N_5994,N_7068);
nand U9625 (N_9625,N_6412,N_5890);
and U9626 (N_9626,N_5852,N_6346);
nand U9627 (N_9627,N_5509,N_6677);
or U9628 (N_9628,N_5605,N_6909);
nor U9629 (N_9629,N_5585,N_7247);
nand U9630 (N_9630,N_7239,N_6216);
nand U9631 (N_9631,N_7432,N_6084);
and U9632 (N_9632,N_5064,N_6988);
or U9633 (N_9633,N_7372,N_6593);
and U9634 (N_9634,N_7064,N_5373);
nand U9635 (N_9635,N_6170,N_5302);
or U9636 (N_9636,N_6965,N_5099);
nor U9637 (N_9637,N_7049,N_6109);
or U9638 (N_9638,N_7141,N_5850);
or U9639 (N_9639,N_6432,N_6563);
and U9640 (N_9640,N_5499,N_6414);
nor U9641 (N_9641,N_7439,N_6242);
nand U9642 (N_9642,N_7317,N_5788);
nor U9643 (N_9643,N_5310,N_6274);
or U9644 (N_9644,N_5227,N_7410);
or U9645 (N_9645,N_5130,N_5775);
or U9646 (N_9646,N_6421,N_6246);
nand U9647 (N_9647,N_6771,N_5511);
nand U9648 (N_9648,N_5317,N_5241);
or U9649 (N_9649,N_5110,N_5123);
nor U9650 (N_9650,N_7485,N_6913);
nand U9651 (N_9651,N_6805,N_5973);
or U9652 (N_9652,N_7374,N_7395);
nand U9653 (N_9653,N_5549,N_6752);
or U9654 (N_9654,N_7469,N_7430);
nor U9655 (N_9655,N_5640,N_6428);
and U9656 (N_9656,N_7196,N_6252);
or U9657 (N_9657,N_5588,N_5526);
or U9658 (N_9658,N_5785,N_5682);
nor U9659 (N_9659,N_7096,N_5800);
or U9660 (N_9660,N_6640,N_6325);
and U9661 (N_9661,N_6346,N_5487);
and U9662 (N_9662,N_5301,N_5044);
or U9663 (N_9663,N_5835,N_5728);
or U9664 (N_9664,N_6563,N_5488);
nand U9665 (N_9665,N_6947,N_7085);
and U9666 (N_9666,N_5803,N_5758);
nand U9667 (N_9667,N_6326,N_7089);
nand U9668 (N_9668,N_6073,N_6336);
and U9669 (N_9669,N_5169,N_6229);
or U9670 (N_9670,N_5625,N_6094);
or U9671 (N_9671,N_5895,N_6848);
nand U9672 (N_9672,N_5154,N_5345);
nand U9673 (N_9673,N_6781,N_7178);
or U9674 (N_9674,N_6219,N_7463);
nand U9675 (N_9675,N_5126,N_7438);
nand U9676 (N_9676,N_5690,N_7201);
and U9677 (N_9677,N_6144,N_5786);
nor U9678 (N_9678,N_6968,N_5647);
and U9679 (N_9679,N_6810,N_6196);
and U9680 (N_9680,N_6312,N_6338);
or U9681 (N_9681,N_5676,N_5493);
or U9682 (N_9682,N_6064,N_6061);
and U9683 (N_9683,N_7246,N_7203);
nand U9684 (N_9684,N_6360,N_5490);
nand U9685 (N_9685,N_5366,N_7115);
and U9686 (N_9686,N_5734,N_7318);
nand U9687 (N_9687,N_6446,N_6923);
and U9688 (N_9688,N_5822,N_6045);
or U9689 (N_9689,N_7440,N_5776);
nand U9690 (N_9690,N_7381,N_6440);
or U9691 (N_9691,N_6084,N_6558);
nand U9692 (N_9692,N_7382,N_6734);
nor U9693 (N_9693,N_7391,N_6685);
xor U9694 (N_9694,N_6677,N_5452);
and U9695 (N_9695,N_5854,N_6470);
and U9696 (N_9696,N_7289,N_6454);
and U9697 (N_9697,N_5279,N_7123);
and U9698 (N_9698,N_5629,N_5938);
and U9699 (N_9699,N_5826,N_5358);
nor U9700 (N_9700,N_6705,N_7425);
nand U9701 (N_9701,N_5127,N_5820);
nor U9702 (N_9702,N_7091,N_7379);
nand U9703 (N_9703,N_5416,N_5439);
or U9704 (N_9704,N_5576,N_6443);
nand U9705 (N_9705,N_5727,N_7093);
and U9706 (N_9706,N_7118,N_5148);
nor U9707 (N_9707,N_6921,N_6514);
and U9708 (N_9708,N_6088,N_7436);
nor U9709 (N_9709,N_7314,N_5778);
nor U9710 (N_9710,N_7001,N_5259);
nor U9711 (N_9711,N_6214,N_5039);
or U9712 (N_9712,N_6778,N_5162);
and U9713 (N_9713,N_5039,N_5489);
nand U9714 (N_9714,N_6482,N_5737);
nand U9715 (N_9715,N_7386,N_6874);
and U9716 (N_9716,N_7181,N_5268);
nor U9717 (N_9717,N_6142,N_7047);
nand U9718 (N_9718,N_7355,N_5623);
and U9719 (N_9719,N_5756,N_7259);
nand U9720 (N_9720,N_6197,N_7181);
nor U9721 (N_9721,N_6675,N_6157);
and U9722 (N_9722,N_6092,N_6102);
or U9723 (N_9723,N_5887,N_7140);
xor U9724 (N_9724,N_6329,N_6698);
nor U9725 (N_9725,N_5034,N_5166);
nor U9726 (N_9726,N_5326,N_7285);
nor U9727 (N_9727,N_6471,N_5164);
and U9728 (N_9728,N_5127,N_5633);
nor U9729 (N_9729,N_6842,N_6196);
or U9730 (N_9730,N_7271,N_6071);
nor U9731 (N_9731,N_6769,N_6188);
and U9732 (N_9732,N_5406,N_5991);
xnor U9733 (N_9733,N_7296,N_5294);
or U9734 (N_9734,N_6609,N_6726);
nor U9735 (N_9735,N_7250,N_5762);
or U9736 (N_9736,N_6005,N_6758);
and U9737 (N_9737,N_7112,N_5179);
nand U9738 (N_9738,N_5233,N_6112);
and U9739 (N_9739,N_6512,N_6043);
or U9740 (N_9740,N_6052,N_6915);
nor U9741 (N_9741,N_5036,N_6750);
nand U9742 (N_9742,N_7400,N_6562);
and U9743 (N_9743,N_7191,N_6154);
and U9744 (N_9744,N_5446,N_6143);
nand U9745 (N_9745,N_5521,N_5437);
and U9746 (N_9746,N_5092,N_6063);
nor U9747 (N_9747,N_5733,N_6721);
or U9748 (N_9748,N_6750,N_6404);
nor U9749 (N_9749,N_6383,N_5115);
and U9750 (N_9750,N_5710,N_5853);
or U9751 (N_9751,N_6520,N_6386);
nor U9752 (N_9752,N_5587,N_5597);
and U9753 (N_9753,N_6604,N_5655);
nand U9754 (N_9754,N_6874,N_7294);
nor U9755 (N_9755,N_7373,N_5938);
nand U9756 (N_9756,N_6781,N_5889);
and U9757 (N_9757,N_6958,N_6379);
and U9758 (N_9758,N_7118,N_7499);
nand U9759 (N_9759,N_5724,N_6124);
and U9760 (N_9760,N_7026,N_6677);
nand U9761 (N_9761,N_7156,N_6870);
and U9762 (N_9762,N_5294,N_7486);
or U9763 (N_9763,N_6270,N_5649);
and U9764 (N_9764,N_7290,N_6926);
or U9765 (N_9765,N_6791,N_5935);
nor U9766 (N_9766,N_7359,N_5757);
nor U9767 (N_9767,N_6137,N_7002);
and U9768 (N_9768,N_5883,N_6470);
and U9769 (N_9769,N_6840,N_6315);
nand U9770 (N_9770,N_5220,N_5057);
or U9771 (N_9771,N_5770,N_5758);
nor U9772 (N_9772,N_6017,N_5002);
and U9773 (N_9773,N_6698,N_6432);
nand U9774 (N_9774,N_5480,N_6063);
nand U9775 (N_9775,N_5053,N_5755);
nor U9776 (N_9776,N_7469,N_7263);
or U9777 (N_9777,N_6847,N_6322);
nor U9778 (N_9778,N_5288,N_5635);
or U9779 (N_9779,N_6077,N_6884);
nor U9780 (N_9780,N_6228,N_6445);
and U9781 (N_9781,N_5311,N_5983);
nand U9782 (N_9782,N_7187,N_6871);
or U9783 (N_9783,N_6862,N_6403);
nand U9784 (N_9784,N_6937,N_5600);
or U9785 (N_9785,N_5136,N_5016);
or U9786 (N_9786,N_6432,N_6387);
and U9787 (N_9787,N_6972,N_7128);
or U9788 (N_9788,N_7059,N_5896);
and U9789 (N_9789,N_6670,N_6000);
nor U9790 (N_9790,N_6492,N_7308);
or U9791 (N_9791,N_7415,N_7356);
and U9792 (N_9792,N_5284,N_5886);
and U9793 (N_9793,N_7152,N_7381);
nand U9794 (N_9794,N_6116,N_5233);
or U9795 (N_9795,N_5246,N_7342);
or U9796 (N_9796,N_5344,N_6593);
or U9797 (N_9797,N_6568,N_6062);
nor U9798 (N_9798,N_5345,N_6500);
nor U9799 (N_9799,N_6314,N_6188);
or U9800 (N_9800,N_7338,N_6809);
and U9801 (N_9801,N_5130,N_6681);
and U9802 (N_9802,N_5062,N_5275);
nand U9803 (N_9803,N_7341,N_7236);
nand U9804 (N_9804,N_7112,N_5748);
and U9805 (N_9805,N_5043,N_6383);
or U9806 (N_9806,N_6491,N_5130);
or U9807 (N_9807,N_6719,N_6967);
nand U9808 (N_9808,N_6146,N_7241);
nor U9809 (N_9809,N_5043,N_6789);
or U9810 (N_9810,N_6532,N_5932);
and U9811 (N_9811,N_7362,N_6436);
nor U9812 (N_9812,N_6730,N_6438);
nand U9813 (N_9813,N_6418,N_5291);
or U9814 (N_9814,N_5768,N_7452);
nor U9815 (N_9815,N_6800,N_6010);
and U9816 (N_9816,N_5787,N_5978);
and U9817 (N_9817,N_5398,N_6177);
nor U9818 (N_9818,N_6842,N_6198);
or U9819 (N_9819,N_5040,N_6113);
or U9820 (N_9820,N_6751,N_5264);
and U9821 (N_9821,N_5269,N_5055);
or U9822 (N_9822,N_6201,N_5554);
or U9823 (N_9823,N_6781,N_5370);
nor U9824 (N_9824,N_7065,N_5903);
nand U9825 (N_9825,N_6044,N_5598);
and U9826 (N_9826,N_5825,N_7174);
nand U9827 (N_9827,N_5891,N_6717);
or U9828 (N_9828,N_6792,N_5524);
nand U9829 (N_9829,N_7389,N_7448);
and U9830 (N_9830,N_7409,N_7088);
nand U9831 (N_9831,N_6218,N_6086);
nand U9832 (N_9832,N_5520,N_7256);
nand U9833 (N_9833,N_6981,N_7423);
and U9834 (N_9834,N_5300,N_6028);
and U9835 (N_9835,N_7455,N_5934);
or U9836 (N_9836,N_6490,N_6101);
nand U9837 (N_9837,N_6837,N_7312);
or U9838 (N_9838,N_6982,N_5684);
nand U9839 (N_9839,N_5893,N_6654);
or U9840 (N_9840,N_5406,N_5317);
nand U9841 (N_9841,N_5096,N_5240);
and U9842 (N_9842,N_5122,N_7372);
nor U9843 (N_9843,N_5973,N_6345);
or U9844 (N_9844,N_6954,N_6051);
nand U9845 (N_9845,N_7360,N_7001);
or U9846 (N_9846,N_7269,N_7134);
or U9847 (N_9847,N_6969,N_5336);
nand U9848 (N_9848,N_5679,N_7170);
nor U9849 (N_9849,N_6044,N_5139);
nand U9850 (N_9850,N_5365,N_5681);
nand U9851 (N_9851,N_6201,N_6379);
nor U9852 (N_9852,N_6437,N_5227);
or U9853 (N_9853,N_7086,N_5501);
or U9854 (N_9854,N_6468,N_6439);
nor U9855 (N_9855,N_5572,N_5318);
nor U9856 (N_9856,N_6185,N_6642);
nor U9857 (N_9857,N_5688,N_5421);
or U9858 (N_9858,N_6337,N_6595);
nor U9859 (N_9859,N_5574,N_5204);
or U9860 (N_9860,N_6190,N_6929);
nand U9861 (N_9861,N_6012,N_6513);
and U9862 (N_9862,N_6729,N_5538);
nand U9863 (N_9863,N_7133,N_5288);
nor U9864 (N_9864,N_6181,N_6629);
and U9865 (N_9865,N_5666,N_6291);
nand U9866 (N_9866,N_7238,N_6012);
or U9867 (N_9867,N_5816,N_6762);
nand U9868 (N_9868,N_6628,N_5251);
nor U9869 (N_9869,N_7108,N_5719);
nand U9870 (N_9870,N_5754,N_5475);
and U9871 (N_9871,N_6508,N_7010);
nand U9872 (N_9872,N_7030,N_5188);
nand U9873 (N_9873,N_5164,N_5331);
or U9874 (N_9874,N_6052,N_6014);
or U9875 (N_9875,N_6151,N_6832);
nor U9876 (N_9876,N_5141,N_7429);
nand U9877 (N_9877,N_5317,N_5927);
or U9878 (N_9878,N_5129,N_7064);
nand U9879 (N_9879,N_5390,N_7317);
nand U9880 (N_9880,N_6259,N_6842);
and U9881 (N_9881,N_6145,N_5509);
or U9882 (N_9882,N_7029,N_5196);
and U9883 (N_9883,N_5105,N_6602);
or U9884 (N_9884,N_5724,N_6520);
and U9885 (N_9885,N_5851,N_5495);
and U9886 (N_9886,N_6540,N_5320);
and U9887 (N_9887,N_6234,N_5810);
nand U9888 (N_9888,N_6207,N_6652);
nor U9889 (N_9889,N_5778,N_6740);
or U9890 (N_9890,N_5841,N_6285);
nor U9891 (N_9891,N_7388,N_5964);
xnor U9892 (N_9892,N_6692,N_6346);
or U9893 (N_9893,N_5620,N_6494);
or U9894 (N_9894,N_6947,N_7260);
nor U9895 (N_9895,N_7142,N_5956);
nor U9896 (N_9896,N_6355,N_7393);
or U9897 (N_9897,N_5685,N_5782);
nand U9898 (N_9898,N_5483,N_6859);
and U9899 (N_9899,N_5146,N_7292);
and U9900 (N_9900,N_6516,N_5859);
or U9901 (N_9901,N_5577,N_5298);
or U9902 (N_9902,N_7376,N_6625);
nor U9903 (N_9903,N_7485,N_6258);
and U9904 (N_9904,N_6791,N_5519);
or U9905 (N_9905,N_5193,N_5402);
and U9906 (N_9906,N_6714,N_5155);
nor U9907 (N_9907,N_5245,N_6192);
nor U9908 (N_9908,N_6536,N_6145);
and U9909 (N_9909,N_6538,N_6204);
nor U9910 (N_9910,N_5065,N_6241);
nor U9911 (N_9911,N_6431,N_7224);
or U9912 (N_9912,N_7386,N_5899);
or U9913 (N_9913,N_6687,N_5787);
and U9914 (N_9914,N_6250,N_7430);
and U9915 (N_9915,N_6636,N_5578);
or U9916 (N_9916,N_5495,N_6667);
and U9917 (N_9917,N_5057,N_6145);
nor U9918 (N_9918,N_5470,N_7445);
nand U9919 (N_9919,N_6023,N_5781);
nand U9920 (N_9920,N_5267,N_5659);
or U9921 (N_9921,N_7043,N_5650);
nor U9922 (N_9922,N_5140,N_6770);
nand U9923 (N_9923,N_7239,N_5771);
nor U9924 (N_9924,N_5205,N_5937);
or U9925 (N_9925,N_6152,N_5948);
nor U9926 (N_9926,N_5104,N_6483);
nand U9927 (N_9927,N_5244,N_5262);
or U9928 (N_9928,N_6074,N_5875);
nor U9929 (N_9929,N_5741,N_7032);
and U9930 (N_9930,N_7476,N_5793);
nand U9931 (N_9931,N_5458,N_6164);
or U9932 (N_9932,N_5947,N_7160);
nor U9933 (N_9933,N_5879,N_7272);
nand U9934 (N_9934,N_7123,N_7455);
nand U9935 (N_9935,N_7376,N_6272);
nand U9936 (N_9936,N_6278,N_7356);
or U9937 (N_9937,N_6103,N_6772);
xnor U9938 (N_9938,N_5816,N_6146);
and U9939 (N_9939,N_5976,N_6443);
nor U9940 (N_9940,N_6166,N_7074);
nand U9941 (N_9941,N_5758,N_6347);
nor U9942 (N_9942,N_6191,N_5222);
and U9943 (N_9943,N_6329,N_7384);
or U9944 (N_9944,N_6225,N_6233);
nor U9945 (N_9945,N_5389,N_6721);
nor U9946 (N_9946,N_7400,N_7390);
and U9947 (N_9947,N_5387,N_5846);
or U9948 (N_9948,N_5473,N_7020);
nand U9949 (N_9949,N_5353,N_6380);
nand U9950 (N_9950,N_6193,N_5696);
xor U9951 (N_9951,N_6892,N_6911);
nand U9952 (N_9952,N_5445,N_6933);
and U9953 (N_9953,N_5973,N_5056);
or U9954 (N_9954,N_5195,N_6869);
nor U9955 (N_9955,N_5512,N_5396);
and U9956 (N_9956,N_5127,N_5602);
or U9957 (N_9957,N_5947,N_5142);
and U9958 (N_9958,N_6292,N_5930);
and U9959 (N_9959,N_6552,N_6469);
nor U9960 (N_9960,N_5223,N_6919);
nor U9961 (N_9961,N_5808,N_7130);
or U9962 (N_9962,N_6226,N_6065);
nor U9963 (N_9963,N_7005,N_7294);
or U9964 (N_9964,N_6710,N_6368);
or U9965 (N_9965,N_6862,N_6615);
and U9966 (N_9966,N_6638,N_5162);
nand U9967 (N_9967,N_6615,N_7341);
or U9968 (N_9968,N_6956,N_6529);
or U9969 (N_9969,N_6211,N_7435);
nor U9970 (N_9970,N_5361,N_6363);
nor U9971 (N_9971,N_6063,N_6682);
and U9972 (N_9972,N_5750,N_7358);
nor U9973 (N_9973,N_6808,N_5212);
and U9974 (N_9974,N_7489,N_7251);
or U9975 (N_9975,N_6072,N_6471);
or U9976 (N_9976,N_6887,N_5577);
nand U9977 (N_9977,N_7445,N_6075);
or U9978 (N_9978,N_6611,N_7143);
nand U9979 (N_9979,N_6048,N_6849);
nand U9980 (N_9980,N_7370,N_5550);
nor U9981 (N_9981,N_6569,N_5850);
nor U9982 (N_9982,N_5919,N_5383);
or U9983 (N_9983,N_7466,N_7461);
and U9984 (N_9984,N_7183,N_6487);
or U9985 (N_9985,N_5747,N_6807);
nand U9986 (N_9986,N_5079,N_6485);
nor U9987 (N_9987,N_5717,N_6321);
and U9988 (N_9988,N_6770,N_7119);
and U9989 (N_9989,N_5790,N_5268);
nand U9990 (N_9990,N_6631,N_6042);
and U9991 (N_9991,N_6233,N_6399);
or U9992 (N_9992,N_6189,N_6239);
and U9993 (N_9993,N_5583,N_6381);
nand U9994 (N_9994,N_6254,N_7437);
nor U9995 (N_9995,N_6865,N_7211);
nand U9996 (N_9996,N_5459,N_5774);
nand U9997 (N_9997,N_6020,N_5584);
nand U9998 (N_9998,N_5713,N_5872);
and U9999 (N_9999,N_5286,N_7376);
nand UO_0 (O_0,N_8802,N_9064);
nor UO_1 (O_1,N_7821,N_8022);
and UO_2 (O_2,N_9657,N_8431);
or UO_3 (O_3,N_9871,N_8807);
nand UO_4 (O_4,N_8051,N_9327);
nor UO_5 (O_5,N_8767,N_7527);
and UO_6 (O_6,N_7914,N_8904);
nor UO_7 (O_7,N_8706,N_8787);
or UO_8 (O_8,N_7731,N_9085);
nor UO_9 (O_9,N_7912,N_8662);
nand UO_10 (O_10,N_8135,N_8997);
nand UO_11 (O_11,N_8960,N_9671);
nor UO_12 (O_12,N_7689,N_8038);
nor UO_13 (O_13,N_7622,N_7817);
xor UO_14 (O_14,N_7795,N_8832);
or UO_15 (O_15,N_9666,N_8836);
and UO_16 (O_16,N_7812,N_9922);
nor UO_17 (O_17,N_8373,N_8837);
or UO_18 (O_18,N_7707,N_7909);
and UO_19 (O_19,N_7803,N_9945);
or UO_20 (O_20,N_9323,N_8446);
nor UO_21 (O_21,N_8217,N_8284);
nand UO_22 (O_22,N_7726,N_7587);
or UO_23 (O_23,N_8275,N_8303);
nor UO_24 (O_24,N_7678,N_9895);
nor UO_25 (O_25,N_8930,N_8118);
or UO_26 (O_26,N_8131,N_8660);
nor UO_27 (O_27,N_8870,N_8577);
nor UO_28 (O_28,N_7719,N_8633);
and UO_29 (O_29,N_9599,N_7672);
and UO_30 (O_30,N_9620,N_9449);
nor UO_31 (O_31,N_9114,N_8067);
nor UO_32 (O_32,N_9097,N_7528);
nor UO_33 (O_33,N_8472,N_8138);
or UO_34 (O_34,N_8008,N_9157);
or UO_35 (O_35,N_7789,N_9083);
nand UO_36 (O_36,N_9023,N_7907);
nand UO_37 (O_37,N_7950,N_8567);
nor UO_38 (O_38,N_9569,N_9631);
and UO_39 (O_39,N_8996,N_7946);
or UO_40 (O_40,N_8913,N_7603);
and UO_41 (O_41,N_7582,N_8682);
and UO_42 (O_42,N_7893,N_7694);
or UO_43 (O_43,N_8495,N_9742);
or UO_44 (O_44,N_8911,N_8085);
xor UO_45 (O_45,N_8484,N_7586);
or UO_46 (O_46,N_8849,N_9744);
or UO_47 (O_47,N_9564,N_8490);
or UO_48 (O_48,N_7598,N_9681);
xor UO_49 (O_49,N_8784,N_9234);
nand UO_50 (O_50,N_7976,N_7576);
nand UO_51 (O_51,N_9302,N_9081);
nand UO_52 (O_52,N_8745,N_7855);
nand UO_53 (O_53,N_9904,N_8600);
and UO_54 (O_54,N_9825,N_7787);
and UO_55 (O_55,N_9534,N_8690);
nor UO_56 (O_56,N_9557,N_9929);
nor UO_57 (O_57,N_8089,N_9916);
nor UO_58 (O_58,N_9288,N_8300);
nor UO_59 (O_59,N_9044,N_7616);
nor UO_60 (O_60,N_9866,N_8331);
nor UO_61 (O_61,N_8024,N_9978);
nor UO_62 (O_62,N_9504,N_8047);
nand UO_63 (O_63,N_8114,N_9455);
nor UO_64 (O_64,N_8732,N_9458);
and UO_65 (O_65,N_7838,N_8740);
nand UO_66 (O_66,N_8090,N_8675);
nand UO_67 (O_67,N_7670,N_8841);
or UO_68 (O_68,N_7693,N_7686);
nand UO_69 (O_69,N_9646,N_8729);
nand UO_70 (O_70,N_8752,N_7846);
and UO_71 (O_71,N_9988,N_8888);
and UO_72 (O_72,N_8921,N_9964);
and UO_73 (O_73,N_9493,N_8358);
nand UO_74 (O_74,N_8687,N_9628);
or UO_75 (O_75,N_8272,N_8670);
nor UO_76 (O_76,N_8599,N_9851);
nor UO_77 (O_77,N_9275,N_8795);
nor UO_78 (O_78,N_8834,N_9863);
nor UO_79 (O_79,N_9315,N_8769);
nand UO_80 (O_80,N_8334,N_8892);
and UO_81 (O_81,N_8553,N_8189);
nand UO_82 (O_82,N_8467,N_7891);
nand UO_83 (O_83,N_8780,N_7905);
and UO_84 (O_84,N_7700,N_9622);
or UO_85 (O_85,N_9185,N_8560);
or UO_86 (O_86,N_9210,N_9954);
nor UO_87 (O_87,N_7965,N_7602);
or UO_88 (O_88,N_8658,N_8698);
nor UO_89 (O_89,N_8361,N_8853);
nor UO_90 (O_90,N_7948,N_8678);
and UO_91 (O_91,N_9475,N_9959);
nand UO_92 (O_92,N_9498,N_8129);
and UO_93 (O_93,N_8520,N_9103);
nor UO_94 (O_94,N_8514,N_7865);
nor UO_95 (O_95,N_8044,N_9618);
or UO_96 (O_96,N_9838,N_8323);
nor UO_97 (O_97,N_7649,N_8954);
or UO_98 (O_98,N_9295,N_8677);
nand UO_99 (O_99,N_9247,N_7966);
or UO_100 (O_100,N_9764,N_8269);
nand UO_101 (O_101,N_9193,N_8449);
nor UO_102 (O_102,N_9052,N_8301);
nand UO_103 (O_103,N_9716,N_8153);
and UO_104 (O_104,N_9365,N_9071);
or UO_105 (O_105,N_9518,N_7796);
nor UO_106 (O_106,N_8348,N_8518);
or UO_107 (O_107,N_8052,N_9488);
nand UO_108 (O_108,N_8053,N_7880);
or UO_109 (O_109,N_9382,N_9481);
and UO_110 (O_110,N_9746,N_9484);
nand UO_111 (O_111,N_7816,N_7645);
nor UO_112 (O_112,N_8015,N_8861);
and UO_113 (O_113,N_8844,N_9651);
nor UO_114 (O_114,N_8639,N_9086);
or UO_115 (O_115,N_7975,N_9099);
nor UO_116 (O_116,N_8213,N_8032);
nor UO_117 (O_117,N_8757,N_8883);
or UO_118 (O_118,N_8572,N_7922);
and UO_119 (O_119,N_7878,N_8042);
nand UO_120 (O_120,N_8215,N_7799);
or UO_121 (O_121,N_9093,N_8187);
nor UO_122 (O_122,N_8266,N_7577);
nand UO_123 (O_123,N_7804,N_8880);
and UO_124 (O_124,N_8483,N_9819);
nor UO_125 (O_125,N_8686,N_7684);
nand UO_126 (O_126,N_7537,N_8626);
nor UO_127 (O_127,N_7571,N_9600);
nand UO_128 (O_128,N_8978,N_8447);
and UO_129 (O_129,N_9139,N_9537);
and UO_130 (O_130,N_7579,N_8414);
and UO_131 (O_131,N_9870,N_9669);
nand UO_132 (O_132,N_8357,N_9722);
or UO_133 (O_133,N_7859,N_7725);
or UO_134 (O_134,N_9374,N_9563);
and UO_135 (O_135,N_8970,N_9240);
or UO_136 (O_136,N_8655,N_9667);
and UO_137 (O_137,N_7779,N_8456);
nor UO_138 (O_138,N_7839,N_9642);
and UO_139 (O_139,N_9732,N_7657);
nand UO_140 (O_140,N_9508,N_7546);
nor UO_141 (O_141,N_7911,N_8010);
or UO_142 (O_142,N_9963,N_8260);
nor UO_143 (O_143,N_9440,N_9340);
and UO_144 (O_144,N_9334,N_7944);
or UO_145 (O_145,N_9252,N_9843);
nand UO_146 (O_146,N_7674,N_8276);
or UO_147 (O_147,N_9554,N_9796);
nor UO_148 (O_148,N_8859,N_8661);
or UO_149 (O_149,N_9645,N_9282);
nand UO_150 (O_150,N_9689,N_8758);
and UO_151 (O_151,N_8250,N_7933);
nand UO_152 (O_152,N_9845,N_9806);
nand UO_153 (O_153,N_9899,N_9224);
or UO_154 (O_154,N_9468,N_8195);
or UO_155 (O_155,N_9349,N_9360);
or UO_156 (O_156,N_9443,N_9042);
and UO_157 (O_157,N_8799,N_8879);
or UO_158 (O_158,N_9636,N_7718);
nor UO_159 (O_159,N_8214,N_8207);
and UO_160 (O_160,N_9026,N_9354);
nand UO_161 (O_161,N_8221,N_9972);
nor UO_162 (O_162,N_8916,N_8541);
and UO_163 (O_163,N_9608,N_9406);
and UO_164 (O_164,N_7745,N_7849);
nor UO_165 (O_165,N_7815,N_9239);
or UO_166 (O_166,N_9731,N_9723);
nand UO_167 (O_167,N_9160,N_8155);
nor UO_168 (O_168,N_7900,N_9080);
nand UO_169 (O_169,N_8905,N_8606);
nor UO_170 (O_170,N_7740,N_8491);
nand UO_171 (O_171,N_9319,N_8143);
and UO_172 (O_172,N_7814,N_9505);
nand UO_173 (O_173,N_9528,N_7723);
nand UO_174 (O_174,N_7947,N_7942);
and UO_175 (O_175,N_7737,N_9907);
nor UO_176 (O_176,N_7675,N_8124);
and UO_177 (O_177,N_9982,N_9359);
and UO_178 (O_178,N_7998,N_9820);
nor UO_179 (O_179,N_9930,N_8239);
nand UO_180 (O_180,N_8561,N_8501);
or UO_181 (O_181,N_8427,N_7570);
nand UO_182 (O_182,N_8545,N_8866);
and UO_183 (O_183,N_8352,N_9206);
or UO_184 (O_184,N_9420,N_9459);
or UO_185 (O_185,N_8112,N_8186);
nand UO_186 (O_186,N_9673,N_8528);
nor UO_187 (O_187,N_7962,N_9803);
or UO_188 (O_188,N_7877,N_7507);
nand UO_189 (O_189,N_9719,N_9092);
nor UO_190 (O_190,N_9311,N_9865);
and UO_191 (O_191,N_9523,N_9637);
nor UO_192 (O_192,N_8665,N_9704);
and UO_193 (O_193,N_8333,N_8324);
or UO_194 (O_194,N_9290,N_8666);
xor UO_195 (O_195,N_9626,N_9441);
nand UO_196 (O_196,N_8393,N_7643);
and UO_197 (O_197,N_9258,N_7663);
and UO_198 (O_198,N_8671,N_8336);
or UO_199 (O_199,N_8152,N_9204);
xnor UO_200 (O_200,N_8293,N_9521);
nor UO_201 (O_201,N_9011,N_9379);
or UO_202 (O_202,N_9771,N_8234);
and UO_203 (O_203,N_8909,N_9708);
nor UO_204 (O_204,N_9678,N_8014);
or UO_205 (O_205,N_8631,N_8533);
nand UO_206 (O_206,N_8183,N_9770);
nor UO_207 (O_207,N_9222,N_9602);
or UO_208 (O_208,N_7646,N_7956);
or UO_209 (O_209,N_7770,N_8689);
nor UO_210 (O_210,N_7851,N_8081);
nand UO_211 (O_211,N_9718,N_8181);
nor UO_212 (O_212,N_8382,N_8874);
nor UO_213 (O_213,N_8307,N_9874);
nand UO_214 (O_214,N_8851,N_9022);
nor UO_215 (O_215,N_8165,N_9684);
and UO_216 (O_216,N_8951,N_9353);
and UO_217 (O_217,N_9800,N_8615);
and UO_218 (O_218,N_8522,N_9386);
or UO_219 (O_219,N_9162,N_8313);
nand UO_220 (O_220,N_9355,N_9680);
nand UO_221 (O_221,N_9749,N_8783);
nand UO_222 (O_222,N_8095,N_9824);
or UO_223 (O_223,N_9159,N_9546);
and UO_224 (O_224,N_8873,N_9077);
nand UO_225 (O_225,N_9107,N_8203);
xnor UO_226 (O_226,N_7664,N_8236);
or UO_227 (O_227,N_8901,N_9171);
and UO_228 (O_228,N_9695,N_8317);
and UO_229 (O_229,N_8728,N_8206);
and UO_230 (O_230,N_9853,N_8999);
or UO_231 (O_231,N_9691,N_8977);
nand UO_232 (O_232,N_9402,N_9585);
and UO_233 (O_233,N_9809,N_7682);
nor UO_234 (O_234,N_9961,N_9289);
or UO_235 (O_235,N_7943,N_9203);
or UO_236 (O_236,N_7692,N_9209);
nand UO_237 (O_237,N_9404,N_8725);
nor UO_238 (O_238,N_8992,N_9738);
nand UO_239 (O_239,N_7773,N_8254);
nand UO_240 (O_240,N_9492,N_8136);
nand UO_241 (O_241,N_9520,N_9432);
nand UO_242 (O_242,N_8743,N_7919);
nand UO_243 (O_243,N_9140,N_9860);
and UO_244 (O_244,N_7983,N_8942);
nand UO_245 (O_245,N_8228,N_8180);
and UO_246 (O_246,N_7504,N_9677);
or UO_247 (O_247,N_7801,N_9358);
and UO_248 (O_248,N_9109,N_8605);
and UO_249 (O_249,N_7769,N_9532);
or UO_250 (O_250,N_9967,N_9592);
and UO_251 (O_251,N_9775,N_8676);
and UO_252 (O_252,N_8416,N_9456);
or UO_253 (O_253,N_7797,N_8209);
and UO_254 (O_254,N_8641,N_8077);
nand UO_255 (O_255,N_9872,N_7721);
nand UO_256 (O_256,N_8157,N_7824);
nand UO_257 (O_257,N_9605,N_7930);
nand UO_258 (O_258,N_9105,N_9448);
nand UO_259 (O_259,N_7753,N_9074);
nand UO_260 (O_260,N_7613,N_9952);
nor UO_261 (O_261,N_8184,N_7658);
and UO_262 (O_262,N_8342,N_8391);
and UO_263 (O_263,N_9877,N_7977);
and UO_264 (O_264,N_9989,N_9477);
nor UO_265 (O_265,N_7829,N_9012);
nor UO_266 (O_266,N_7755,N_8499);
nor UO_267 (O_267,N_8268,N_8292);
xnor UO_268 (O_268,N_9245,N_9920);
nand UO_269 (O_269,N_8691,N_9510);
nor UO_270 (O_270,N_8154,N_8094);
nor UO_271 (O_271,N_9141,N_9451);
and UO_272 (O_272,N_7677,N_7756);
nor UO_273 (O_273,N_9313,N_9652);
nand UO_274 (O_274,N_9471,N_8482);
or UO_275 (O_275,N_8309,N_8111);
nand UO_276 (O_276,N_9367,N_9474);
nand UO_277 (O_277,N_8488,N_7805);
nand UO_278 (O_278,N_7866,N_8814);
or UO_279 (O_279,N_8616,N_8684);
nand UO_280 (O_280,N_8473,N_8471);
nand UO_281 (O_281,N_7713,N_8233);
and UO_282 (O_282,N_8506,N_7539);
nand UO_283 (O_283,N_8969,N_9985);
nand UO_284 (O_284,N_9342,N_8701);
and UO_285 (O_285,N_7802,N_9163);
or UO_286 (O_286,N_9479,N_7863);
and UO_287 (O_287,N_8663,N_8882);
nand UO_288 (O_288,N_8881,N_7701);
or UO_289 (O_289,N_9392,N_8647);
nand UO_290 (O_290,N_9390,N_7705);
or UO_291 (O_291,N_7923,N_8311);
nor UO_292 (O_292,N_9197,N_9987);
or UO_293 (O_293,N_8602,N_9395);
and UO_294 (O_294,N_8959,N_9951);
nand UO_295 (O_295,N_9547,N_7985);
and UO_296 (O_296,N_8164,N_9403);
and UO_297 (O_297,N_8542,N_8995);
nand UO_298 (O_298,N_7786,N_9060);
nand UO_299 (O_299,N_7808,N_9005);
nor UO_300 (O_300,N_7955,N_9867);
and UO_301 (O_301,N_9164,N_9836);
or UO_302 (O_302,N_8731,N_7704);
nor UO_303 (O_303,N_7973,N_9960);
nand UO_304 (O_304,N_8903,N_9507);
nor UO_305 (O_305,N_8127,N_9303);
and UO_306 (O_306,N_9047,N_8394);
and UO_307 (O_307,N_9030,N_9352);
and UO_308 (O_308,N_9388,N_8243);
nand UO_309 (O_309,N_8188,N_9729);
xnor UO_310 (O_310,N_8279,N_9229);
nand UO_311 (O_311,N_9970,N_9807);
nand UO_312 (O_312,N_8212,N_7784);
or UO_313 (O_313,N_8737,N_8068);
nand UO_314 (O_314,N_8305,N_9199);
nand UO_315 (O_315,N_9277,N_9172);
nor UO_316 (O_316,N_7515,N_8420);
and UO_317 (O_317,N_8265,N_9580);
and UO_318 (O_318,N_8840,N_9152);
nor UO_319 (O_319,N_8764,N_8249);
and UO_320 (O_320,N_8825,N_9454);
or UO_321 (O_321,N_9055,N_8497);
nand UO_322 (O_322,N_7848,N_8101);
or UO_323 (O_323,N_8544,N_8381);
nor UO_324 (O_324,N_9401,N_8778);
or UO_325 (O_325,N_8494,N_7563);
nand UO_326 (O_326,N_7999,N_9413);
or UO_327 (O_327,N_7621,N_7592);
and UO_328 (O_328,N_9274,N_7992);
or UO_329 (O_329,N_8173,N_9848);
or UO_330 (O_330,N_8286,N_7883);
nand UO_331 (O_331,N_9726,N_7596);
nand UO_332 (O_332,N_7666,N_9552);
and UO_333 (O_333,N_9123,N_8906);
or UO_334 (O_334,N_7500,N_9869);
nor UO_335 (O_335,N_9514,N_8838);
nand UO_336 (O_336,N_9984,N_8256);
nor UO_337 (O_337,N_9511,N_8868);
nor UO_338 (O_338,N_9006,N_7888);
and UO_339 (O_339,N_8355,N_9018);
nand UO_340 (O_340,N_8592,N_7588);
nand UO_341 (O_341,N_9994,N_7858);
nor UO_342 (O_342,N_9227,N_8711);
and UO_343 (O_343,N_9572,N_8339);
nand UO_344 (O_344,N_9291,N_8232);
nand UO_345 (O_345,N_8974,N_9950);
xnor UO_346 (O_346,N_8412,N_7655);
nand UO_347 (O_347,N_8770,N_8283);
nor UO_348 (O_348,N_9378,N_7780);
xor UO_349 (O_349,N_7869,N_7629);
nor UO_350 (O_350,N_8399,N_9721);
nand UO_351 (O_351,N_8466,N_8811);
nand UO_352 (O_352,N_9625,N_9371);
and UO_353 (O_353,N_8822,N_8925);
nand UO_354 (O_354,N_9331,N_8445);
nor UO_355 (O_355,N_9177,N_8299);
nand UO_356 (O_356,N_8823,N_8009);
or UO_357 (O_357,N_9442,N_8980);
nor UO_358 (O_358,N_8877,N_8894);
nor UO_359 (O_359,N_8216,N_7642);
nand UO_360 (O_360,N_7825,N_9329);
or UO_361 (O_361,N_8429,N_8798);
xor UO_362 (O_362,N_8280,N_7970);
nor UO_363 (O_363,N_9898,N_8989);
nand UO_364 (O_364,N_8549,N_9834);
or UO_365 (O_365,N_8063,N_9001);
xnor UO_366 (O_366,N_9629,N_9846);
or UO_367 (O_367,N_9915,N_9849);
nor UO_368 (O_368,N_9408,N_7766);
nand UO_369 (O_369,N_9128,N_8340);
nor UO_370 (O_370,N_7777,N_9814);
nor UO_371 (O_371,N_7757,N_7525);
nor UO_372 (O_372,N_9059,N_9641);
nor UO_373 (O_373,N_8197,N_8168);
or UO_374 (O_374,N_7548,N_8296);
or UO_375 (O_375,N_9529,N_8789);
nand UO_376 (O_376,N_8958,N_7867);
and UO_377 (O_377,N_7688,N_9790);
nand UO_378 (O_378,N_7860,N_8120);
nor UO_379 (O_379,N_9188,N_9316);
or UO_380 (O_380,N_9590,N_8507);
nor UO_381 (O_381,N_9754,N_9253);
nand UO_382 (O_382,N_8613,N_8792);
or UO_383 (O_383,N_8573,N_7533);
and UO_384 (O_384,N_8657,N_9463);
nor UO_385 (O_385,N_7750,N_8707);
and UO_386 (O_386,N_9362,N_8222);
or UO_387 (O_387,N_9079,N_9527);
or UO_388 (O_388,N_8177,N_9276);
nor UO_389 (O_389,N_8788,N_8235);
nand UO_390 (O_390,N_9142,N_9453);
and UO_391 (O_391,N_9539,N_9427);
and UO_392 (O_392,N_8934,N_8946);
and UO_393 (O_393,N_8607,N_9430);
or UO_394 (O_394,N_9394,N_8779);
or UO_395 (O_395,N_9595,N_9896);
and UO_396 (O_396,N_9412,N_9804);
and UO_397 (O_397,N_8765,N_9926);
and UO_398 (O_398,N_7857,N_9658);
nor UO_399 (O_399,N_7772,N_9762);
nor UO_400 (O_400,N_8257,N_7641);
or UO_401 (O_401,N_9842,N_7882);
nand UO_402 (O_402,N_9400,N_7640);
and UO_403 (O_403,N_8200,N_7547);
and UO_404 (O_404,N_9810,N_9501);
and UO_405 (O_405,N_7526,N_8441);
nor UO_406 (O_406,N_9668,N_9217);
and UO_407 (O_407,N_7996,N_8629);
or UO_408 (O_408,N_7538,N_9126);
xor UO_409 (O_409,N_8774,N_9573);
and UO_410 (O_410,N_8454,N_7845);
nand UO_411 (O_411,N_9343,N_9815);
nor UO_412 (O_412,N_9397,N_8656);
and UO_413 (O_413,N_9616,N_9181);
and UO_414 (O_414,N_8536,N_8872);
and UO_415 (O_415,N_9158,N_8371);
nor UO_416 (O_416,N_7782,N_8386);
nand UO_417 (O_417,N_9170,N_9272);
or UO_418 (O_418,N_9470,N_9567);
nand UO_419 (O_419,N_9783,N_7873);
nor UO_420 (O_420,N_8869,N_8023);
nor UO_421 (O_421,N_9971,N_8049);
and UO_422 (O_422,N_9761,N_9757);
or UO_423 (O_423,N_8018,N_7968);
nor UO_424 (O_424,N_9482,N_9231);
or UO_425 (O_425,N_9997,N_7562);
and UO_426 (O_426,N_9587,N_8793);
and UO_427 (O_427,N_9610,N_9320);
nor UO_428 (O_428,N_9917,N_8363);
nor UO_429 (O_429,N_7768,N_7842);
nand UO_430 (O_430,N_9750,N_7583);
nor UO_431 (O_431,N_9812,N_7578);
nor UO_432 (O_432,N_9073,N_8074);
nor UO_433 (O_433,N_7758,N_8163);
nand UO_434 (O_434,N_9736,N_8896);
nor UO_435 (O_435,N_9875,N_9974);
nor UO_436 (O_436,N_8178,N_9324);
or UO_437 (O_437,N_8130,N_7555);
nor UO_438 (O_438,N_7699,N_8845);
or UO_439 (O_439,N_7729,N_8121);
or UO_440 (O_440,N_7987,N_9647);
nor UO_441 (O_441,N_7508,N_9249);
and UO_442 (O_442,N_8083,N_8462);
and UO_443 (O_443,N_8404,N_9782);
or UO_444 (O_444,N_9020,N_8408);
and UO_445 (O_445,N_8683,N_7650);
and UO_446 (O_446,N_8620,N_9751);
or UO_447 (O_447,N_8436,N_9486);
nor UO_448 (O_448,N_9986,N_9462);
or UO_449 (O_449,N_9698,N_9476);
nand UO_450 (O_450,N_9586,N_8100);
or UO_451 (O_451,N_8571,N_9908);
nand UO_452 (O_452,N_7903,N_7518);
nand UO_453 (O_453,N_8985,N_9017);
nor UO_454 (O_454,N_9983,N_9603);
and UO_455 (O_455,N_9061,N_9781);
or UO_456 (O_456,N_7886,N_8295);
nand UO_457 (O_457,N_9497,N_9644);
nand UO_458 (O_458,N_7775,N_7607);
nor UO_459 (O_459,N_9279,N_8673);
or UO_460 (O_460,N_7519,N_9553);
nand UO_461 (O_461,N_9992,N_9385);
nor UO_462 (O_462,N_8563,N_9799);
nand UO_463 (O_463,N_8538,N_9174);
nand UO_464 (O_464,N_9098,N_7852);
and UO_465 (O_465,N_8517,N_7516);
nand UO_466 (O_466,N_9134,N_9176);
and UO_467 (O_467,N_8891,N_9146);
and UO_468 (O_468,N_7549,N_9912);
nor UO_469 (O_469,N_9542,N_7568);
nand UO_470 (O_470,N_8418,N_9213);
nor UO_471 (O_471,N_8277,N_8547);
xnor UO_472 (O_472,N_7819,N_9014);
and UO_473 (O_473,N_8744,N_7744);
nor UO_474 (O_474,N_8413,N_8423);
nor UO_475 (O_475,N_8829,N_9921);
nand UO_476 (O_476,N_8804,N_9007);
nand UO_477 (O_477,N_7589,N_7634);
and UO_478 (O_478,N_7899,N_9701);
and UO_479 (O_479,N_9832,N_8835);
or UO_480 (O_480,N_9594,N_8559);
or UO_481 (O_481,N_9794,N_9422);
nand UO_482 (O_482,N_9269,N_9743);
and UO_483 (O_483,N_9377,N_8659);
nand UO_484 (O_484,N_7632,N_8947);
and UO_485 (O_485,N_9178,N_9145);
or UO_486 (O_486,N_9472,N_8580);
nor UO_487 (O_487,N_9632,N_8259);
or UO_488 (O_488,N_9568,N_7931);
nor UO_489 (O_489,N_7558,N_9087);
nand UO_490 (O_490,N_8335,N_9286);
or UO_491 (O_491,N_9541,N_7894);
nand UO_492 (O_492,N_8900,N_9082);
and UO_493 (O_493,N_8952,N_7826);
nand UO_494 (O_494,N_8718,N_9363);
or UO_495 (O_495,N_7542,N_8043);
and UO_496 (O_496,N_8551,N_8172);
nand UO_497 (O_497,N_8253,N_8037);
nand UO_498 (O_498,N_9094,N_9410);
nand UO_499 (O_499,N_7614,N_9307);
nor UO_500 (O_500,N_9469,N_8278);
nand UO_501 (O_501,N_9583,N_9955);
and UO_502 (O_502,N_9318,N_9856);
xor UO_503 (O_503,N_8123,N_7920);
nand UO_504 (O_504,N_9619,N_7742);
nand UO_505 (O_505,N_9000,N_9376);
or UO_506 (O_506,N_9067,N_8006);
and UO_507 (O_507,N_8858,N_7834);
and UO_508 (O_508,N_8050,N_7654);
or UO_509 (O_509,N_8990,N_9655);
nor UO_510 (O_510,N_8424,N_9236);
and UO_511 (O_511,N_8475,N_7567);
nor UO_512 (O_512,N_7844,N_8007);
and UO_513 (O_513,N_8442,N_9298);
and UO_514 (O_514,N_9991,N_8612);
or UO_515 (O_515,N_9381,N_9889);
nor UO_516 (O_516,N_8161,N_9076);
nand UO_517 (O_517,N_7599,N_7952);
and UO_518 (O_518,N_9127,N_9745);
nand UO_519 (O_519,N_7961,N_9341);
nand UO_520 (O_520,N_8438,N_9882);
nand UO_521 (O_521,N_8017,N_9980);
nor UO_522 (O_522,N_9256,N_9862);
or UO_523 (O_523,N_9649,N_7806);
or UO_524 (O_524,N_9223,N_8987);
nand UO_525 (O_525,N_9424,N_8046);
nand UO_526 (O_526,N_9075,N_8627);
and UO_527 (O_527,N_8550,N_7875);
nor UO_528 (O_528,N_9167,N_8889);
nand UO_529 (O_529,N_9335,N_8529);
or UO_530 (O_530,N_7653,N_8714);
nand UO_531 (O_531,N_7511,N_9522);
nor UO_532 (O_532,N_7902,N_7778);
and UO_533 (O_533,N_8332,N_8957);
nand UO_534 (O_534,N_8805,N_8712);
nor UO_535 (O_535,N_8219,N_9308);
and UO_536 (O_536,N_9688,N_7506);
or UO_537 (O_537,N_8622,N_9027);
nand UO_538 (O_538,N_7637,N_9788);
and UO_539 (O_539,N_7932,N_9571);
nor UO_540 (O_540,N_7874,N_8011);
nor UO_541 (O_541,N_8871,N_9190);
and UO_542 (O_542,N_8940,N_7695);
and UO_543 (O_543,N_8531,N_8512);
and UO_544 (O_544,N_9133,N_9839);
and UO_545 (O_545,N_7529,N_7597);
and UO_546 (O_546,N_8530,N_9122);
nor UO_547 (O_547,N_9503,N_9426);
nor UO_548 (O_548,N_9664,N_9570);
nand UO_549 (O_549,N_8918,N_7556);
and UO_550 (O_550,N_9995,N_7680);
nor UO_551 (O_551,N_8667,N_7584);
nor UO_552 (O_552,N_8407,N_7544);
and UO_553 (O_553,N_7792,N_9473);
or UO_554 (O_554,N_8555,N_7934);
nor UO_555 (O_555,N_8831,N_9201);
or UO_556 (O_556,N_8621,N_7671);
or UO_557 (O_557,N_8149,N_9822);
nand UO_558 (O_558,N_8320,N_9830);
or UO_559 (O_559,N_8349,N_9478);
nand UO_560 (O_560,N_8099,N_8966);
and UO_561 (O_561,N_9840,N_8579);
and UO_562 (O_562,N_8857,N_9251);
nor UO_563 (O_563,N_9697,N_8196);
and UO_564 (O_564,N_8813,N_8398);
nor UO_565 (O_565,N_8587,N_9460);
nor UO_566 (O_566,N_7747,N_9883);
nor UO_567 (O_567,N_7502,N_9002);
and UO_568 (O_568,N_8469,N_8617);
and UO_569 (O_569,N_8425,N_7590);
nand UO_570 (O_570,N_9888,N_7557);
nand UO_571 (O_571,N_8762,N_8029);
or UO_572 (O_572,N_8158,N_9137);
nand UO_573 (O_573,N_7881,N_9264);
and UO_574 (O_574,N_9670,N_9648);
and UO_575 (O_575,N_8890,N_8298);
nand UO_576 (O_576,N_9901,N_9357);
nand UO_577 (O_577,N_8117,N_9990);
and UO_578 (O_578,N_9558,N_9593);
or UO_579 (O_579,N_7608,N_9965);
or UO_580 (O_580,N_9156,N_8182);
and UO_581 (O_581,N_7938,N_9576);
and UO_582 (O_582,N_9633,N_8144);
nor UO_583 (O_583,N_7536,N_8915);
or UO_584 (O_584,N_9581,N_8941);
nor UO_585 (O_585,N_8148,N_7990);
or UO_586 (O_586,N_9306,N_8948);
and UO_587 (O_587,N_9450,N_9333);
and UO_588 (O_588,N_7836,N_9271);
and UO_589 (O_589,N_7505,N_8230);
nand UO_590 (O_590,N_8886,N_8460);
or UO_591 (O_591,N_9465,N_8492);
nand UO_592 (O_592,N_9675,N_9149);
or UO_593 (O_593,N_7788,N_9769);
and UO_594 (O_594,N_9310,N_9421);
nand UO_595 (O_595,N_9265,N_7609);
nor UO_596 (O_596,N_8045,N_8922);
nor UO_597 (O_597,N_8937,N_8532);
or UO_598 (O_598,N_7785,N_9638);
and UO_599 (O_599,N_8082,N_9878);
or UO_600 (O_600,N_9847,N_8039);
nand UO_601 (O_601,N_9423,N_9737);
nor UO_602 (O_602,N_7870,N_9634);
or UO_603 (O_603,N_8596,N_8887);
nor UO_604 (O_604,N_8353,N_8422);
or UO_605 (O_605,N_8723,N_7709);
nand UO_606 (O_606,N_7639,N_8034);
nor UO_607 (O_607,N_8036,N_9639);
or UO_608 (O_608,N_9262,N_9759);
nor UO_609 (O_609,N_9207,N_9297);
nand UO_610 (O_610,N_9063,N_8322);
or UO_611 (O_611,N_8150,N_7960);
nor UO_612 (O_612,N_9347,N_7651);
and UO_613 (O_613,N_8761,N_8931);
or UO_614 (O_614,N_8463,N_8634);
nor UO_615 (O_615,N_7746,N_7921);
or UO_616 (O_616,N_9332,N_8345);
or UO_617 (O_617,N_8643,N_9235);
nand UO_618 (O_618,N_8202,N_8035);
nand UO_619 (O_619,N_8697,N_9548);
or UO_620 (O_620,N_9433,N_7512);
and UO_621 (O_621,N_8343,N_9161);
or UO_622 (O_622,N_9692,N_8703);
nor UO_623 (O_623,N_8385,N_8508);
nor UO_624 (O_624,N_8078,N_9147);
nor UO_625 (O_625,N_8554,N_9280);
and UO_626 (O_626,N_8708,N_8091);
or UO_627 (O_627,N_9516,N_8511);
and UO_628 (O_628,N_7916,N_9939);
nor UO_629 (O_629,N_8070,N_9036);
nand UO_630 (O_630,N_8176,N_8500);
nand UO_631 (O_631,N_8064,N_9419);
nor UO_632 (O_632,N_8610,N_9601);
or UO_633 (O_633,N_8623,N_7954);
nand UO_634 (O_634,N_8086,N_8920);
and UO_635 (O_635,N_8344,N_9555);
nand UO_636 (O_636,N_7604,N_8817);
nand UO_637 (O_637,N_8485,N_8694);
and UO_638 (O_638,N_8493,N_8630);
and UO_639 (O_639,N_8653,N_9205);
and UO_640 (O_640,N_8395,N_8956);
or UO_641 (O_641,N_9057,N_8405);
nand UO_642 (O_642,N_8654,N_9911);
nor UO_643 (O_643,N_8417,N_9730);
nor UO_644 (O_644,N_8751,N_8972);
nand UO_645 (O_645,N_8991,N_8437);
nand UO_646 (O_646,N_9130,N_8674);
nand UO_647 (O_647,N_8597,N_9066);
nor UO_648 (O_648,N_8411,N_9884);
and UO_649 (O_649,N_9941,N_7550);
or UO_650 (O_650,N_8105,N_8820);
or UO_651 (O_651,N_7734,N_8601);
or UO_652 (O_652,N_8924,N_9538);
nor UO_653 (O_653,N_8368,N_9437);
and UO_654 (O_654,N_8939,N_8696);
or UO_655 (O_655,N_7906,N_8267);
nand UO_656 (O_656,N_7601,N_8108);
nand UO_657 (O_657,N_9813,N_9380);
nand UO_658 (O_658,N_8772,N_9973);
xnor UO_659 (O_659,N_9998,N_8928);
nand UO_660 (O_660,N_9182,N_9132);
nor UO_661 (O_661,N_7676,N_8646);
nor UO_662 (O_662,N_9215,N_9574);
nand UO_663 (O_663,N_7915,N_8341);
nand UO_664 (O_664,N_8863,N_9106);
nor UO_665 (O_665,N_9793,N_9577);
nand UO_666 (O_666,N_9735,N_7971);
and UO_667 (O_667,N_7561,N_8428);
and UO_668 (O_668,N_8867,N_9038);
nand UO_669 (O_669,N_8722,N_7591);
nand UO_670 (O_670,N_9949,N_7898);
and UO_671 (O_671,N_9054,N_8073);
or UO_672 (O_672,N_9089,N_7868);
nand UO_673 (O_673,N_8263,N_9927);
and UO_674 (O_674,N_8569,N_9763);
and UO_675 (O_675,N_9243,N_9976);
xor UO_676 (O_676,N_9084,N_8830);
or UO_677 (O_677,N_9364,N_7687);
nand UO_678 (O_678,N_9125,N_8314);
nor UO_679 (O_679,N_7617,N_9278);
nor UO_680 (O_680,N_8548,N_9499);
nand UO_681 (O_681,N_8933,N_8464);
nor UO_682 (O_682,N_9446,N_7509);
nor UO_683 (O_683,N_8330,N_9414);
nor UO_684 (O_684,N_8797,N_7809);
and UO_685 (O_685,N_8727,N_8261);
and UO_686 (O_686,N_7928,N_9344);
nand UO_687 (O_687,N_9411,N_7781);
and UO_688 (O_688,N_8384,N_9962);
and UO_689 (O_689,N_8801,N_7953);
and UO_690 (O_690,N_7913,N_8862);
or UO_691 (O_691,N_9445,N_8584);
or UO_692 (O_692,N_9640,N_7514);
or UO_693 (O_693,N_7522,N_9189);
and UO_694 (O_694,N_9808,N_8973);
nand UO_695 (O_695,N_8651,N_9707);
or UO_696 (O_696,N_8122,N_9894);
nand UO_697 (O_697,N_7994,N_7830);
nor UO_698 (O_698,N_8664,N_9776);
nor UO_699 (O_699,N_8962,N_9119);
nand UO_700 (O_700,N_9356,N_7940);
and UO_701 (O_701,N_9187,N_9436);
nand UO_702 (O_702,N_7748,N_9979);
and UO_703 (O_703,N_9409,N_8833);
nand UO_704 (O_704,N_9712,N_8069);
nand UO_705 (O_705,N_8534,N_8963);
or UO_706 (O_706,N_9301,N_9791);
nand UO_707 (O_707,N_9428,N_8803);
nor UO_708 (O_708,N_9923,N_8282);
and UO_709 (O_709,N_9946,N_8318);
nand UO_710 (O_710,N_8927,N_8109);
and UO_711 (O_711,N_7831,N_9533);
nor UO_712 (O_712,N_8146,N_7585);
or UO_713 (O_713,N_9513,N_7733);
and UO_714 (O_714,N_8402,N_7690);
nand UO_715 (O_715,N_9337,N_9702);
nor UO_716 (O_716,N_9273,N_9905);
or UO_717 (O_717,N_9837,N_9758);
nor UO_718 (O_718,N_9536,N_8162);
and UO_719 (O_719,N_8392,N_8756);
or UO_720 (O_720,N_9049,N_9609);
and UO_721 (O_721,N_8246,N_7569);
or UO_722 (O_722,N_8644,N_9208);
nand UO_723 (O_723,N_8062,N_8988);
nor UO_724 (O_724,N_9257,N_9056);
nand UO_725 (O_725,N_9635,N_8198);
nand UO_726 (O_726,N_7926,N_8258);
nor UO_727 (O_727,N_7981,N_9679);
or UO_728 (O_728,N_9665,N_9494);
nand UO_729 (O_729,N_8251,N_9598);
and UO_730 (O_730,N_9218,N_8848);
nor UO_731 (O_731,N_8480,N_8586);
and UO_732 (O_732,N_7841,N_8350);
nor UO_733 (O_733,N_8430,N_8056);
nand UO_734 (O_734,N_9031,N_9944);
or UO_735 (O_735,N_8557,N_9789);
or UO_736 (O_736,N_9198,N_9784);
and UO_737 (O_737,N_9425,N_9496);
and UO_738 (O_738,N_8072,N_7728);
nor UO_739 (O_739,N_8588,N_9173);
nand UO_740 (O_740,N_9418,N_8961);
and UO_741 (O_741,N_8071,N_8489);
and UO_742 (O_742,N_9168,N_9861);
nand UO_743 (O_743,N_9328,N_9095);
nand UO_744 (O_744,N_9841,N_7862);
nand UO_745 (O_745,N_9614,N_9739);
nand UO_746 (O_746,N_8955,N_7711);
nor UO_747 (O_747,N_8426,N_9051);
nand UO_748 (O_748,N_9774,N_8294);
or UO_749 (O_749,N_9175,N_7850);
or UO_750 (O_750,N_9760,N_9756);
or UO_751 (O_751,N_8796,N_9727);
or UO_752 (O_752,N_8084,N_8583);
nand UO_753 (O_753,N_8503,N_9384);
or UO_754 (O_754,N_9956,N_9039);
or UO_755 (O_755,N_8448,N_9797);
nor UO_756 (O_756,N_7945,N_8210);
and UO_757 (O_757,N_8899,N_8245);
and UO_758 (O_758,N_7984,N_8252);
nand UO_759 (O_759,N_8274,N_7626);
or UO_760 (O_760,N_8194,N_7683);
nor UO_761 (O_761,N_8021,N_7660);
nand UO_762 (O_762,N_8000,N_8306);
or UO_763 (O_763,N_8818,N_7534);
nor UO_764 (O_764,N_9387,N_8125);
nor UO_765 (O_765,N_8581,N_7991);
and UO_766 (O_766,N_8496,N_9116);
and UO_767 (O_767,N_7794,N_8115);
and UO_768 (O_768,N_7566,N_7988);
nor UO_769 (O_769,N_9447,N_7763);
or UO_770 (O_770,N_8054,N_9078);
nand UO_771 (O_771,N_7967,N_9857);
nand UO_772 (O_772,N_9611,N_7908);
or UO_773 (O_773,N_9715,N_7652);
nand UO_774 (O_774,N_7800,N_9650);
and UO_775 (O_775,N_8790,N_9336);
and UO_776 (O_776,N_9035,N_8169);
or UO_777 (O_777,N_7738,N_7861);
nor UO_778 (O_778,N_9958,N_8611);
or UO_779 (O_779,N_8895,N_9407);
nor UO_780 (O_780,N_9226,N_7716);
and UO_781 (O_781,N_9897,N_8360);
and UO_782 (O_782,N_9351,N_8865);
nor UO_783 (O_783,N_9506,N_9019);
or UO_784 (O_784,N_8741,N_8025);
nor UO_785 (O_785,N_9118,N_9893);
nor UO_786 (O_786,N_8379,N_8461);
or UO_787 (O_787,N_9562,N_8435);
nand UO_788 (O_788,N_8288,N_8713);
nand UO_789 (O_789,N_8552,N_8208);
nor UO_790 (O_790,N_7612,N_8884);
and UO_791 (O_791,N_8730,N_8810);
and UO_792 (O_792,N_9773,N_9798);
nand UO_793 (O_793,N_8170,N_8815);
or UO_794 (O_794,N_9464,N_9467);
and UO_795 (O_795,N_8238,N_9623);
nand UO_796 (O_796,N_8364,N_9549);
nand UO_797 (O_797,N_8964,N_9886);
nand UO_798 (O_798,N_9596,N_9373);
nand UO_799 (O_799,N_9993,N_9858);
nor UO_800 (O_800,N_8328,N_9880);
nor UO_801 (O_801,N_8619,N_9879);
and UO_802 (O_802,N_9065,N_9292);
xnor UO_803 (O_803,N_9008,N_9703);
and UO_804 (O_804,N_7611,N_7774);
nand UO_805 (O_805,N_7741,N_8147);
nor UO_806 (O_806,N_8628,N_8004);
nand UO_807 (O_807,N_9627,N_8028);
and UO_808 (O_808,N_8981,N_9165);
nand UO_809 (O_809,N_7630,N_8668);
nor UO_810 (O_810,N_7668,N_7530);
or UO_811 (O_811,N_8096,N_9817);
or UO_812 (O_812,N_8603,N_8079);
nand UO_813 (O_813,N_9515,N_8700);
or UO_814 (O_814,N_8066,N_8327);
and UO_815 (O_815,N_8852,N_8443);
and UO_816 (O_816,N_7736,N_9519);
and UO_817 (O_817,N_9630,N_8458);
nand UO_818 (O_818,N_7958,N_8749);
nand UO_819 (O_819,N_7997,N_7624);
or UO_820 (O_820,N_9579,N_9270);
nand UO_821 (O_821,N_9135,N_9827);
or UO_822 (O_822,N_7635,N_9366);
nand UO_823 (O_823,N_9415,N_7872);
or UO_824 (O_824,N_9710,N_8516);
nor UO_825 (O_825,N_8110,N_9805);
nand UO_826 (O_826,N_8929,N_8031);
nand UO_827 (O_827,N_7935,N_7895);
nand UO_828 (O_828,N_7644,N_9578);
nor UO_829 (O_829,N_8001,N_9267);
or UO_830 (O_830,N_7535,N_9699);
and UO_831 (O_831,N_7820,N_8636);
nor UO_832 (O_832,N_9021,N_8087);
nand UO_833 (O_833,N_8938,N_9968);
nand UO_834 (O_834,N_9582,N_9399);
or UO_835 (O_835,N_9309,N_9220);
or UO_836 (O_836,N_8504,N_7897);
nand UO_837 (O_837,N_8816,N_7939);
nand UO_838 (O_838,N_9643,N_9136);
and UO_839 (O_839,N_7510,N_8809);
nand UO_840 (O_840,N_8897,N_9748);
and UO_841 (O_841,N_7717,N_9765);
nand UO_842 (O_842,N_9046,N_9933);
xor UO_843 (O_843,N_8308,N_9143);
nand UO_844 (O_844,N_7856,N_8346);
or UO_845 (O_845,N_8791,N_7545);
nand UO_846 (O_846,N_8539,N_9540);
nand UO_847 (O_847,N_7714,N_9524);
nand UO_848 (O_848,N_8748,N_8002);
or UO_849 (O_849,N_9966,N_9891);
nand UO_850 (O_850,N_9823,N_9591);
or UO_851 (O_851,N_9195,N_9237);
nand UO_852 (O_852,N_9102,N_7969);
or UO_853 (O_853,N_8415,N_8564);
nand UO_854 (O_854,N_8618,N_9674);
or UO_855 (O_855,N_9069,N_9550);
or UO_856 (O_856,N_8325,N_8546);
or UO_857 (O_857,N_7901,N_9714);
nor UO_858 (O_858,N_8876,N_9296);
or UO_859 (O_859,N_8166,N_9892);
or UO_860 (O_860,N_9914,N_9821);
and UO_861 (O_861,N_8505,N_8224);
nor UO_862 (O_862,N_8794,N_7818);
nor UO_863 (O_863,N_8359,N_9100);
nor UO_864 (O_864,N_8672,N_8967);
and UO_865 (O_865,N_8470,N_7697);
nand UO_866 (O_866,N_7832,N_9439);
or UO_867 (O_867,N_8570,N_8808);
and UO_868 (O_868,N_7659,N_9438);
nand UO_869 (O_869,N_9003,N_8474);
nand UO_870 (O_870,N_8692,N_9034);
or UO_871 (O_871,N_9855,N_8388);
and UO_872 (O_872,N_8637,N_9466);
nor UO_873 (O_873,N_8179,N_9948);
and UO_874 (O_874,N_8827,N_8773);
and UO_875 (O_875,N_7656,N_7673);
nor UO_876 (O_876,N_8374,N_8106);
and UO_877 (O_877,N_8598,N_9248);
or UO_878 (O_878,N_8440,N_8847);
or UO_879 (O_879,N_8098,N_9487);
and UO_880 (O_880,N_8058,N_9480);
nor UO_881 (O_881,N_8609,N_8377);
or UO_882 (O_882,N_9260,N_8632);
nand UO_883 (O_883,N_7679,N_8406);
or UO_884 (O_884,N_8116,N_8720);
and UO_885 (O_885,N_8585,N_8453);
and UO_886 (O_886,N_7937,N_7524);
and UO_887 (O_887,N_9452,N_8191);
nand UO_888 (O_888,N_8645,N_7696);
nand UO_889 (O_889,N_7625,N_7554);
nor UO_890 (O_890,N_8576,N_8242);
nor UO_891 (O_891,N_9868,N_9685);
and UO_892 (O_892,N_7827,N_8540);
and UO_893 (O_893,N_9778,N_9225);
or UO_894 (O_894,N_8434,N_9705);
nor UO_895 (O_895,N_9918,N_8145);
nor UO_896 (O_896,N_7638,N_8747);
xor UO_897 (O_897,N_8369,N_8401);
or UO_898 (O_898,N_8885,N_8821);
nor UO_899 (O_899,N_8487,N_8635);
nand UO_900 (O_900,N_8695,N_9090);
and UO_901 (O_901,N_8367,N_9033);
nand UO_902 (O_902,N_9700,N_8227);
and UO_903 (O_903,N_8574,N_8315);
nor UO_904 (O_904,N_8211,N_9150);
nor UO_905 (O_905,N_9656,N_9138);
nand UO_906 (O_906,N_7791,N_9013);
and UO_907 (O_907,N_8075,N_9940);
and UO_908 (O_908,N_8160,N_7936);
nor UO_909 (O_909,N_8593,N_9934);
nand UO_910 (O_910,N_9396,N_9500);
and UO_911 (O_911,N_9304,N_8855);
or UO_912 (O_912,N_9314,N_9525);
nand UO_913 (O_913,N_9155,N_9509);
and UO_914 (O_914,N_9131,N_8614);
nand UO_915 (O_915,N_7924,N_9202);
and UO_916 (O_916,N_8513,N_8033);
nor UO_917 (O_917,N_8819,N_8193);
and UO_918 (O_918,N_9728,N_8201);
and UO_919 (O_919,N_9300,N_8140);
and UO_920 (O_920,N_9368,N_9864);
and UO_921 (O_921,N_8608,N_9887);
nor UO_922 (O_922,N_8220,N_9975);
nor UO_923 (O_923,N_9321,N_7681);
nand UO_924 (O_924,N_9179,N_7995);
nand UO_925 (O_925,N_7807,N_8704);
nand UO_926 (O_926,N_8240,N_9242);
and UO_927 (O_927,N_9711,N_9828);
and UO_928 (O_928,N_7669,N_9259);
or UO_929 (O_929,N_8702,N_8223);
nor UO_930 (O_930,N_7843,N_8156);
nand UO_931 (O_931,N_8979,N_8624);
nand UO_932 (O_932,N_8968,N_7619);
nand UO_933 (O_933,N_8457,N_8397);
and UO_934 (O_934,N_8409,N_8478);
and UO_935 (O_935,N_8126,N_7703);
nor UO_936 (O_936,N_8486,N_9266);
nand UO_937 (O_937,N_8681,N_8760);
or UO_938 (O_938,N_7595,N_9391);
nor UO_939 (O_939,N_9108,N_7885);
or UO_940 (O_940,N_9435,N_9676);
nand UO_941 (O_941,N_8604,N_7665);
and UO_942 (O_942,N_8943,N_7765);
and UO_943 (O_943,N_7618,N_7560);
and UO_944 (O_944,N_9232,N_8174);
or UO_945 (O_945,N_8768,N_7759);
nand UO_946 (O_946,N_9393,N_9687);
nor UO_947 (O_947,N_8060,N_7835);
nor UO_948 (O_948,N_9148,N_9653);
nand UO_949 (O_949,N_9686,N_7712);
nor UO_950 (O_950,N_9104,N_8945);
nor UO_951 (O_951,N_7662,N_9943);
nor UO_952 (O_952,N_8926,N_9683);
nor UO_953 (O_953,N_8142,N_8750);
nand UO_954 (O_954,N_8137,N_8648);
or UO_955 (O_955,N_8128,N_9713);
and UO_956 (O_956,N_9584,N_8316);
or UO_957 (O_957,N_8362,N_7565);
and UO_958 (O_958,N_8468,N_8568);
and UO_959 (O_959,N_9305,N_9909);
and UO_960 (O_960,N_7887,N_7811);
and UO_961 (O_961,N_8878,N_8289);
nand UO_962 (O_962,N_9370,N_8465);
or UO_963 (O_963,N_7929,N_9777);
xnor UO_964 (O_964,N_8225,N_7581);
nor UO_965 (O_965,N_8735,N_9566);
nand UO_966 (O_966,N_9416,N_8983);
or UO_967 (O_967,N_8419,N_7986);
nand UO_968 (O_968,N_8290,N_7540);
nor UO_969 (O_969,N_8403,N_9350);
and UO_970 (O_970,N_7523,N_9854);
nor UO_971 (O_971,N_9490,N_7823);
and UO_972 (O_972,N_8459,N_8917);
and UO_973 (O_973,N_8650,N_8244);
nand UO_974 (O_974,N_7837,N_8652);
nor UO_975 (O_975,N_8102,N_8986);
nand UO_976 (O_976,N_8719,N_8241);
or UO_977 (O_977,N_7896,N_8061);
nand UO_978 (O_978,N_7520,N_9169);
nor UO_979 (O_979,N_8030,N_8566);
or UO_980 (O_980,N_7871,N_9906);
and UO_981 (O_981,N_9517,N_8226);
nor UO_982 (O_982,N_9281,N_8151);
nor UO_983 (O_983,N_9792,N_9244);
and UO_984 (O_984,N_8383,N_9556);
and UO_985 (O_985,N_8262,N_8828);
or UO_986 (O_986,N_8746,N_7949);
nor UO_987 (O_987,N_9330,N_7879);
or UO_988 (O_988,N_9682,N_9795);
nand UO_989 (O_989,N_8354,N_8975);
nand UO_990 (O_990,N_9028,N_7989);
nand UO_991 (O_991,N_9752,N_7661);
or UO_992 (O_992,N_8558,N_8476);
nor UO_993 (O_993,N_7580,N_9016);
nor UO_994 (O_994,N_9969,N_9228);
or UO_995 (O_995,N_8537,N_9873);
nor UO_996 (O_996,N_7620,N_9200);
and UO_997 (O_997,N_8763,N_7559);
nand UO_998 (O_998,N_9062,N_7749);
nand UO_999 (O_999,N_9859,N_9345);
and UO_1000 (O_1000,N_8378,N_9902);
or UO_1001 (O_1001,N_9925,N_9551);
nor UO_1002 (O_1002,N_9191,N_8824);
nor UO_1003 (O_1003,N_7573,N_9931);
nand UO_1004 (O_1004,N_9913,N_9942);
and UO_1005 (O_1005,N_8755,N_9530);
xnor UO_1006 (O_1006,N_9233,N_9772);
nor UO_1007 (O_1007,N_9040,N_8119);
nand UO_1008 (O_1008,N_9876,N_9230);
or UO_1009 (O_1009,N_9740,N_8771);
nand UO_1010 (O_1010,N_9151,N_9346);
nor UO_1011 (O_1011,N_7706,N_8535);
nand UO_1012 (O_1012,N_8013,N_9535);
or UO_1013 (O_1013,N_8133,N_7715);
or UO_1014 (O_1014,N_8826,N_8839);
and UO_1015 (O_1015,N_8842,N_9560);
and UO_1016 (O_1016,N_7951,N_7980);
xnor UO_1017 (O_1017,N_9015,N_9221);
and UO_1018 (O_1018,N_8271,N_7889);
and UO_1019 (O_1019,N_8040,N_9461);
or UO_1020 (O_1020,N_9129,N_8521);
and UO_1021 (O_1021,N_7776,N_8510);
and UO_1022 (O_1022,N_8270,N_9753);
or UO_1023 (O_1023,N_9375,N_9254);
nand UO_1024 (O_1024,N_9890,N_9431);
or UO_1025 (O_1025,N_9043,N_9660);
nor UO_1026 (O_1026,N_8347,N_7754);
or UO_1027 (O_1027,N_7876,N_7793);
and UO_1028 (O_1028,N_8724,N_9919);
or UO_1029 (O_1029,N_9050,N_8366);
nand UO_1030 (O_1030,N_8141,N_8338);
nand UO_1031 (O_1031,N_9429,N_7925);
or UO_1032 (O_1032,N_8281,N_7941);
and UO_1033 (O_1033,N_9246,N_9121);
nor UO_1034 (O_1034,N_9531,N_8027);
nand UO_1035 (O_1035,N_9621,N_9690);
or UO_1036 (O_1036,N_8380,N_7884);
and UO_1037 (O_1037,N_8782,N_9489);
and UO_1038 (O_1038,N_8455,N_9900);
nand UO_1039 (O_1039,N_7764,N_8132);
nand UO_1040 (O_1040,N_9787,N_9559);
nand UO_1041 (O_1041,N_8843,N_9212);
and UO_1042 (O_1042,N_7771,N_9372);
or UO_1043 (O_1043,N_8291,N_8591);
and UO_1044 (O_1044,N_8594,N_9733);
nand UO_1045 (O_1045,N_7600,N_8781);
nand UO_1046 (O_1046,N_9068,N_9417);
nor UO_1047 (O_1047,N_8304,N_8575);
and UO_1048 (O_1048,N_7979,N_9924);
or UO_1049 (O_1049,N_7972,N_7982);
nand UO_1050 (O_1050,N_9785,N_9589);
nand UO_1051 (O_1051,N_9194,N_8481);
or UO_1052 (O_1052,N_8753,N_7783);
nand UO_1053 (O_1053,N_8875,N_8104);
or UO_1054 (O_1054,N_9885,N_8734);
nor UO_1055 (O_1055,N_8107,N_8097);
or UO_1056 (O_1056,N_9096,N_9826);
nor UO_1057 (O_1057,N_8297,N_9317);
and UO_1058 (O_1058,N_9910,N_7963);
or UO_1059 (O_1059,N_8372,N_9048);
nor UO_1060 (O_1060,N_9383,N_7720);
nor UO_1061 (O_1061,N_8638,N_7918);
nor UO_1062 (O_1062,N_9444,N_8971);
and UO_1063 (O_1063,N_8994,N_7628);
nand UO_1064 (O_1064,N_9312,N_8582);
nor UO_1065 (O_1065,N_8914,N_9010);
nor UO_1066 (O_1066,N_9434,N_8998);
nand UO_1067 (O_1067,N_7917,N_8736);
nor UO_1068 (O_1068,N_7564,N_9936);
or UO_1069 (O_1069,N_8860,N_7702);
nand UO_1070 (O_1070,N_8984,N_9338);
and UO_1071 (O_1071,N_9485,N_9935);
or UO_1072 (O_1072,N_9624,N_8721);
nor UO_1073 (O_1073,N_9196,N_9741);
and UO_1074 (O_1074,N_9238,N_9144);
nand UO_1075 (O_1075,N_8337,N_8949);
or UO_1076 (O_1076,N_9607,N_9299);
and UO_1077 (O_1077,N_9706,N_8526);
nand UO_1078 (O_1078,N_8649,N_9709);
nand UO_1079 (O_1079,N_8229,N_8680);
nor UO_1080 (O_1080,N_9348,N_7521);
or UO_1081 (O_1081,N_7959,N_9457);
and UO_1082 (O_1082,N_9725,N_7517);
nor UO_1083 (O_1083,N_9575,N_8139);
and UO_1084 (O_1084,N_8679,N_8302);
nor UO_1085 (O_1085,N_8329,N_8237);
nor UO_1086 (O_1086,N_7593,N_9101);
nor UO_1087 (O_1087,N_9717,N_8310);
nand UO_1088 (O_1088,N_9831,N_9766);
nor UO_1089 (O_1089,N_8255,N_8451);
or UO_1090 (O_1090,N_8432,N_7761);
nand UO_1091 (O_1091,N_8590,N_9661);
or UO_1092 (O_1092,N_9786,N_7594);
and UO_1093 (O_1093,N_8688,N_7691);
nand UO_1094 (O_1094,N_7732,N_8982);
nand UO_1095 (O_1095,N_9285,N_7572);
nand UO_1096 (O_1096,N_9811,N_9113);
nor UO_1097 (O_1097,N_8519,N_9072);
nand UO_1098 (O_1098,N_9025,N_8850);
and UO_1099 (O_1099,N_8525,N_9881);
nor UO_1100 (O_1100,N_8048,N_8854);
nand UO_1101 (O_1101,N_8134,N_8932);
or UO_1102 (O_1102,N_7636,N_8976);
nand UO_1103 (O_1103,N_8375,N_7730);
and UO_1104 (O_1104,N_8993,N_8450);
and UO_1105 (O_1105,N_8965,N_9545);
nand UO_1106 (O_1106,N_8041,N_7553);
or UO_1107 (O_1107,N_8351,N_8204);
nor UO_1108 (O_1108,N_8726,N_8776);
and UO_1109 (O_1109,N_8312,N_7685);
nor UO_1110 (O_1110,N_7735,N_9693);
nand UO_1111 (O_1111,N_9180,N_9091);
and UO_1112 (O_1112,N_7910,N_9495);
nor UO_1113 (O_1113,N_9154,N_9041);
or UO_1114 (O_1114,N_7767,N_8012);
nand UO_1115 (O_1115,N_8786,N_8543);
nand UO_1116 (O_1116,N_8936,N_7551);
or UO_1117 (O_1117,N_8019,N_8733);
nor UO_1118 (O_1118,N_8923,N_8248);
or UO_1119 (O_1119,N_8775,N_7503);
and UO_1120 (O_1120,N_8185,N_9565);
nand UO_1121 (O_1121,N_7606,N_8093);
or UO_1122 (O_1122,N_8950,N_7615);
nor UO_1123 (O_1123,N_8365,N_7541);
and UO_1124 (O_1124,N_8190,N_9326);
or UO_1125 (O_1125,N_7854,N_8264);
and UO_1126 (O_1126,N_7631,N_9502);
and UO_1127 (O_1127,N_8055,N_9981);
nor UO_1128 (O_1128,N_8026,N_9768);
nand UO_1129 (O_1129,N_7847,N_7698);
and UO_1130 (O_1130,N_9214,N_9604);
nand UO_1131 (O_1131,N_8287,N_8806);
and UO_1132 (O_1132,N_9322,N_8433);
and UO_1133 (O_1133,N_9543,N_7798);
nand UO_1134 (O_1134,N_8717,N_9009);
or UO_1135 (O_1135,N_9662,N_9483);
nor UO_1136 (O_1136,N_8080,N_9615);
or UO_1137 (O_1137,N_8444,N_8812);
and UO_1138 (O_1138,N_9659,N_8766);
nor UO_1139 (O_1139,N_8715,N_8710);
or UO_1140 (O_1140,N_8759,N_9293);
nand UO_1141 (O_1141,N_9112,N_9283);
nor UO_1142 (O_1142,N_8205,N_9903);
or UO_1143 (O_1143,N_8556,N_8524);
nor UO_1144 (O_1144,N_8742,N_9045);
or UO_1145 (O_1145,N_8192,N_7724);
and UO_1146 (O_1146,N_9117,N_9361);
and UO_1147 (O_1147,N_8400,N_9937);
or UO_1148 (O_1148,N_8705,N_9835);
nor UO_1149 (O_1149,N_7648,N_8800);
nand UO_1150 (O_1150,N_7647,N_9938);
nor UO_1151 (O_1151,N_9953,N_9124);
nand UO_1152 (O_1152,N_8410,N_9284);
nand UO_1153 (O_1153,N_9287,N_9389);
nand UO_1154 (O_1154,N_7833,N_9999);
and UO_1155 (O_1155,N_7853,N_8387);
nand UO_1156 (O_1156,N_8376,N_8919);
and UO_1157 (O_1157,N_8159,N_7552);
nor UO_1158 (O_1158,N_7710,N_9816);
nand UO_1159 (O_1159,N_9617,N_7722);
nand UO_1160 (O_1160,N_9829,N_9720);
or UO_1161 (O_1161,N_8777,N_8910);
nor UO_1162 (O_1162,N_8175,N_8092);
nand UO_1163 (O_1163,N_8477,N_8319);
nor UO_1164 (O_1164,N_8565,N_8562);
nor UO_1165 (O_1165,N_9780,N_8247);
nor UO_1166 (O_1166,N_9928,N_7708);
nand UO_1167 (O_1167,N_7575,N_7727);
and UO_1168 (O_1168,N_9802,N_9216);
nor UO_1169 (O_1169,N_9029,N_8912);
nand UO_1170 (O_1170,N_9192,N_9037);
or UO_1171 (O_1171,N_8709,N_8509);
or UO_1172 (O_1172,N_7739,N_9767);
or UO_1173 (O_1173,N_8285,N_9672);
nand UO_1174 (O_1174,N_7627,N_8088);
nand UO_1175 (O_1175,N_8396,N_8699);
nand UO_1176 (O_1176,N_7574,N_8527);
nor UO_1177 (O_1177,N_8893,N_7822);
nand UO_1178 (O_1178,N_9398,N_8640);
nor UO_1179 (O_1179,N_7751,N_9339);
nor UO_1180 (O_1180,N_8113,N_8935);
nor UO_1181 (O_1181,N_8785,N_9255);
or UO_1182 (O_1182,N_8065,N_9544);
and UO_1183 (O_1183,N_9250,N_9241);
or UO_1184 (O_1184,N_9512,N_9526);
xor UO_1185 (O_1185,N_9058,N_8578);
or UO_1186 (O_1186,N_9263,N_8390);
nand UO_1187 (O_1187,N_7531,N_8273);
or UO_1188 (O_1188,N_9696,N_7605);
nor UO_1189 (O_1189,N_9491,N_8907);
nand UO_1190 (O_1190,N_8171,N_8523);
and UO_1191 (O_1191,N_9186,N_9612);
nand UO_1192 (O_1192,N_8864,N_9211);
nor UO_1193 (O_1193,N_9957,N_9325);
or UO_1194 (O_1194,N_8479,N_9747);
nor UO_1195 (O_1195,N_7790,N_8003);
and UO_1196 (O_1196,N_8076,N_8693);
or UO_1197 (O_1197,N_8515,N_8716);
and UO_1198 (O_1198,N_9183,N_9947);
nor UO_1199 (O_1199,N_9588,N_9932);
or UO_1200 (O_1200,N_9663,N_8020);
nand UO_1201 (O_1201,N_9184,N_9597);
nand UO_1202 (O_1202,N_8944,N_7978);
nand UO_1203 (O_1203,N_8754,N_9833);
nor UO_1204 (O_1204,N_8642,N_8856);
and UO_1205 (O_1205,N_9111,N_9977);
nor UO_1206 (O_1206,N_7813,N_9779);
nor UO_1207 (O_1207,N_9755,N_9405);
nor UO_1208 (O_1208,N_7532,N_8356);
or UO_1209 (O_1209,N_8326,N_7667);
nor UO_1210 (O_1210,N_7610,N_8953);
or UO_1211 (O_1211,N_7760,N_7752);
and UO_1212 (O_1212,N_8685,N_9613);
or UO_1213 (O_1213,N_7623,N_8908);
or UO_1214 (O_1214,N_9219,N_9268);
and UO_1215 (O_1215,N_7810,N_9850);
nor UO_1216 (O_1216,N_9724,N_8589);
nor UO_1217 (O_1217,N_9115,N_7513);
nor UO_1218 (O_1218,N_7762,N_7904);
nand UO_1219 (O_1219,N_9032,N_8738);
or UO_1220 (O_1220,N_9369,N_9606);
and UO_1221 (O_1221,N_7927,N_9110);
nand UO_1222 (O_1222,N_7864,N_9654);
and UO_1223 (O_1223,N_7964,N_9053);
nand UO_1224 (O_1224,N_8421,N_9004);
nor UO_1225 (O_1225,N_8502,N_8059);
or UO_1226 (O_1226,N_7633,N_9261);
nor UO_1227 (O_1227,N_9070,N_9166);
nor UO_1228 (O_1228,N_7743,N_9734);
or UO_1229 (O_1229,N_8103,N_8321);
and UO_1230 (O_1230,N_8625,N_8595);
nor UO_1231 (O_1231,N_9153,N_8389);
and UO_1232 (O_1232,N_8218,N_9088);
or UO_1233 (O_1233,N_8057,N_8898);
nand UO_1234 (O_1234,N_7957,N_8498);
and UO_1235 (O_1235,N_7974,N_8167);
and UO_1236 (O_1236,N_8199,N_8739);
and UO_1237 (O_1237,N_9996,N_7828);
nor UO_1238 (O_1238,N_9294,N_8669);
and UO_1239 (O_1239,N_9120,N_8452);
nor UO_1240 (O_1240,N_9024,N_8016);
and UO_1241 (O_1241,N_9694,N_8439);
and UO_1242 (O_1242,N_7892,N_8902);
and UO_1243 (O_1243,N_9801,N_9844);
nand UO_1244 (O_1244,N_7543,N_7993);
or UO_1245 (O_1245,N_7840,N_8231);
nor UO_1246 (O_1246,N_7890,N_7501);
nor UO_1247 (O_1247,N_8370,N_8005);
or UO_1248 (O_1248,N_9818,N_8846);
nand UO_1249 (O_1249,N_9852,N_9561);
nor UO_1250 (O_1250,N_8859,N_8440);
nand UO_1251 (O_1251,N_7962,N_8645);
nand UO_1252 (O_1252,N_8906,N_8279);
and UO_1253 (O_1253,N_8261,N_8231);
nor UO_1254 (O_1254,N_8594,N_8379);
and UO_1255 (O_1255,N_9048,N_8221);
nor UO_1256 (O_1256,N_7693,N_8122);
and UO_1257 (O_1257,N_9102,N_7582);
nor UO_1258 (O_1258,N_7663,N_8704);
nor UO_1259 (O_1259,N_9632,N_7666);
nor UO_1260 (O_1260,N_7577,N_9329);
or UO_1261 (O_1261,N_9784,N_9437);
nand UO_1262 (O_1262,N_8700,N_9568);
or UO_1263 (O_1263,N_8547,N_9721);
and UO_1264 (O_1264,N_7733,N_9710);
nor UO_1265 (O_1265,N_9841,N_9973);
nor UO_1266 (O_1266,N_9505,N_7654);
nand UO_1267 (O_1267,N_9082,N_8689);
nor UO_1268 (O_1268,N_8399,N_8180);
nand UO_1269 (O_1269,N_7601,N_9240);
nor UO_1270 (O_1270,N_8997,N_9659);
xnor UO_1271 (O_1271,N_7653,N_8891);
and UO_1272 (O_1272,N_8501,N_9123);
or UO_1273 (O_1273,N_9140,N_7789);
nand UO_1274 (O_1274,N_9362,N_8826);
or UO_1275 (O_1275,N_7545,N_9859);
or UO_1276 (O_1276,N_8828,N_8562);
nor UO_1277 (O_1277,N_7881,N_8584);
nand UO_1278 (O_1278,N_9679,N_8542);
or UO_1279 (O_1279,N_9826,N_8118);
or UO_1280 (O_1280,N_8504,N_9206);
or UO_1281 (O_1281,N_8762,N_9046);
nand UO_1282 (O_1282,N_8226,N_8358);
nor UO_1283 (O_1283,N_8227,N_8142);
nor UO_1284 (O_1284,N_8833,N_8766);
or UO_1285 (O_1285,N_9622,N_9157);
nor UO_1286 (O_1286,N_9747,N_8311);
xor UO_1287 (O_1287,N_9311,N_8865);
nor UO_1288 (O_1288,N_7519,N_9232);
or UO_1289 (O_1289,N_8493,N_9254);
xnor UO_1290 (O_1290,N_7525,N_8741);
nor UO_1291 (O_1291,N_7935,N_9635);
or UO_1292 (O_1292,N_9494,N_7850);
nor UO_1293 (O_1293,N_7981,N_8076);
nor UO_1294 (O_1294,N_7545,N_9326);
xnor UO_1295 (O_1295,N_7868,N_8734);
nand UO_1296 (O_1296,N_9537,N_9655);
and UO_1297 (O_1297,N_8058,N_9119);
or UO_1298 (O_1298,N_8726,N_9489);
nor UO_1299 (O_1299,N_8110,N_7848);
nand UO_1300 (O_1300,N_8941,N_7567);
xnor UO_1301 (O_1301,N_8883,N_8711);
nand UO_1302 (O_1302,N_9161,N_9570);
and UO_1303 (O_1303,N_9101,N_9172);
or UO_1304 (O_1304,N_9484,N_8898);
nor UO_1305 (O_1305,N_9820,N_9283);
nor UO_1306 (O_1306,N_8876,N_8430);
nand UO_1307 (O_1307,N_9646,N_9932);
or UO_1308 (O_1308,N_9323,N_7909);
nand UO_1309 (O_1309,N_7570,N_8041);
or UO_1310 (O_1310,N_9410,N_8440);
and UO_1311 (O_1311,N_7835,N_7790);
or UO_1312 (O_1312,N_8973,N_8332);
or UO_1313 (O_1313,N_8881,N_8541);
xnor UO_1314 (O_1314,N_8825,N_9602);
nor UO_1315 (O_1315,N_9640,N_8470);
and UO_1316 (O_1316,N_9776,N_8351);
nand UO_1317 (O_1317,N_8395,N_8139);
nor UO_1318 (O_1318,N_9861,N_9134);
and UO_1319 (O_1319,N_9060,N_8383);
and UO_1320 (O_1320,N_8278,N_8443);
nor UO_1321 (O_1321,N_8170,N_9715);
nor UO_1322 (O_1322,N_7530,N_9331);
or UO_1323 (O_1323,N_7548,N_9880);
xor UO_1324 (O_1324,N_9593,N_7649);
or UO_1325 (O_1325,N_9693,N_8429);
and UO_1326 (O_1326,N_9303,N_8844);
nand UO_1327 (O_1327,N_8646,N_9030);
nor UO_1328 (O_1328,N_8165,N_7936);
and UO_1329 (O_1329,N_8981,N_8676);
xor UO_1330 (O_1330,N_9810,N_9420);
nand UO_1331 (O_1331,N_9959,N_8927);
nand UO_1332 (O_1332,N_8618,N_9544);
and UO_1333 (O_1333,N_8755,N_9347);
and UO_1334 (O_1334,N_8271,N_8768);
nand UO_1335 (O_1335,N_7960,N_7581);
or UO_1336 (O_1336,N_8620,N_9106);
or UO_1337 (O_1337,N_8741,N_9540);
and UO_1338 (O_1338,N_9220,N_9013);
and UO_1339 (O_1339,N_9011,N_8239);
and UO_1340 (O_1340,N_7895,N_8756);
xnor UO_1341 (O_1341,N_8424,N_9445);
nand UO_1342 (O_1342,N_8041,N_8192);
or UO_1343 (O_1343,N_9828,N_9910);
nand UO_1344 (O_1344,N_9916,N_8269);
or UO_1345 (O_1345,N_8604,N_8560);
nor UO_1346 (O_1346,N_8558,N_9169);
nand UO_1347 (O_1347,N_9645,N_9314);
nor UO_1348 (O_1348,N_9087,N_8609);
nand UO_1349 (O_1349,N_8539,N_9100);
and UO_1350 (O_1350,N_7880,N_9949);
nor UO_1351 (O_1351,N_8082,N_8998);
and UO_1352 (O_1352,N_9822,N_9797);
or UO_1353 (O_1353,N_9374,N_8440);
nand UO_1354 (O_1354,N_9679,N_9304);
nor UO_1355 (O_1355,N_9183,N_7553);
nand UO_1356 (O_1356,N_8324,N_7852);
nand UO_1357 (O_1357,N_8905,N_8239);
nand UO_1358 (O_1358,N_9788,N_8657);
nor UO_1359 (O_1359,N_8591,N_9067);
or UO_1360 (O_1360,N_9236,N_7712);
nand UO_1361 (O_1361,N_9689,N_9906);
nor UO_1362 (O_1362,N_9856,N_9461);
nor UO_1363 (O_1363,N_7882,N_9499);
nand UO_1364 (O_1364,N_9582,N_8108);
nand UO_1365 (O_1365,N_8539,N_7798);
or UO_1366 (O_1366,N_7515,N_8173);
and UO_1367 (O_1367,N_7585,N_7973);
nand UO_1368 (O_1368,N_8783,N_8364);
or UO_1369 (O_1369,N_7614,N_9417);
and UO_1370 (O_1370,N_7963,N_7753);
nor UO_1371 (O_1371,N_8880,N_9319);
and UO_1372 (O_1372,N_7660,N_8263);
and UO_1373 (O_1373,N_9347,N_9040);
or UO_1374 (O_1374,N_8959,N_8378);
or UO_1375 (O_1375,N_7567,N_8087);
or UO_1376 (O_1376,N_9372,N_9515);
or UO_1377 (O_1377,N_7738,N_8236);
or UO_1378 (O_1378,N_7818,N_8955);
or UO_1379 (O_1379,N_9420,N_9591);
nand UO_1380 (O_1380,N_9411,N_8549);
and UO_1381 (O_1381,N_9839,N_8599);
and UO_1382 (O_1382,N_9151,N_8730);
nand UO_1383 (O_1383,N_8138,N_8322);
nor UO_1384 (O_1384,N_8758,N_7808);
nor UO_1385 (O_1385,N_9731,N_8335);
nor UO_1386 (O_1386,N_8951,N_7590);
nor UO_1387 (O_1387,N_9924,N_9563);
nand UO_1388 (O_1388,N_9817,N_8485);
and UO_1389 (O_1389,N_7967,N_7878);
nand UO_1390 (O_1390,N_9350,N_9293);
nand UO_1391 (O_1391,N_8786,N_9162);
xor UO_1392 (O_1392,N_8955,N_9760);
nor UO_1393 (O_1393,N_9082,N_9466);
nor UO_1394 (O_1394,N_8130,N_8458);
or UO_1395 (O_1395,N_8852,N_9590);
or UO_1396 (O_1396,N_9521,N_8900);
and UO_1397 (O_1397,N_8786,N_7555);
nor UO_1398 (O_1398,N_8401,N_7925);
and UO_1399 (O_1399,N_8280,N_7758);
or UO_1400 (O_1400,N_8161,N_9608);
or UO_1401 (O_1401,N_8260,N_9393);
nor UO_1402 (O_1402,N_9266,N_9016);
or UO_1403 (O_1403,N_9279,N_9861);
nand UO_1404 (O_1404,N_8479,N_7978);
or UO_1405 (O_1405,N_8905,N_7686);
nor UO_1406 (O_1406,N_8740,N_7884);
and UO_1407 (O_1407,N_9763,N_8615);
nand UO_1408 (O_1408,N_8344,N_9900);
and UO_1409 (O_1409,N_8692,N_7975);
or UO_1410 (O_1410,N_8424,N_9624);
nor UO_1411 (O_1411,N_9529,N_8914);
nand UO_1412 (O_1412,N_7897,N_9154);
nor UO_1413 (O_1413,N_8738,N_9714);
nand UO_1414 (O_1414,N_8461,N_8823);
nand UO_1415 (O_1415,N_9672,N_9153);
or UO_1416 (O_1416,N_7529,N_7862);
and UO_1417 (O_1417,N_8681,N_7631);
nand UO_1418 (O_1418,N_7872,N_7531);
and UO_1419 (O_1419,N_9547,N_9607);
nand UO_1420 (O_1420,N_9769,N_9809);
nand UO_1421 (O_1421,N_9792,N_9391);
nand UO_1422 (O_1422,N_9316,N_9618);
and UO_1423 (O_1423,N_9915,N_9421);
nor UO_1424 (O_1424,N_8659,N_9973);
and UO_1425 (O_1425,N_9277,N_9673);
and UO_1426 (O_1426,N_9971,N_8637);
or UO_1427 (O_1427,N_8731,N_9865);
or UO_1428 (O_1428,N_8674,N_8387);
and UO_1429 (O_1429,N_8281,N_8768);
nor UO_1430 (O_1430,N_9587,N_9451);
nand UO_1431 (O_1431,N_8340,N_9735);
nor UO_1432 (O_1432,N_9308,N_8670);
or UO_1433 (O_1433,N_8591,N_9233);
or UO_1434 (O_1434,N_8437,N_8445);
nor UO_1435 (O_1435,N_7993,N_8338);
or UO_1436 (O_1436,N_7769,N_7633);
nand UO_1437 (O_1437,N_9981,N_8480);
or UO_1438 (O_1438,N_9604,N_8089);
and UO_1439 (O_1439,N_9663,N_8050);
nor UO_1440 (O_1440,N_9920,N_8861);
or UO_1441 (O_1441,N_7896,N_7708);
nand UO_1442 (O_1442,N_9612,N_9097);
nor UO_1443 (O_1443,N_7708,N_8949);
nor UO_1444 (O_1444,N_9481,N_7590);
nor UO_1445 (O_1445,N_9269,N_8168);
nor UO_1446 (O_1446,N_8422,N_8510);
nor UO_1447 (O_1447,N_8359,N_9494);
nor UO_1448 (O_1448,N_9932,N_9911);
nand UO_1449 (O_1449,N_8532,N_9601);
nand UO_1450 (O_1450,N_8541,N_9288);
nor UO_1451 (O_1451,N_9081,N_7550);
and UO_1452 (O_1452,N_7862,N_8320);
nand UO_1453 (O_1453,N_8199,N_9833);
nand UO_1454 (O_1454,N_7568,N_8604);
or UO_1455 (O_1455,N_9860,N_8789);
and UO_1456 (O_1456,N_8720,N_9544);
and UO_1457 (O_1457,N_9553,N_8803);
or UO_1458 (O_1458,N_8713,N_8078);
and UO_1459 (O_1459,N_8738,N_8727);
nor UO_1460 (O_1460,N_9260,N_9563);
and UO_1461 (O_1461,N_8601,N_9187);
or UO_1462 (O_1462,N_9640,N_9763);
nand UO_1463 (O_1463,N_7829,N_8317);
or UO_1464 (O_1464,N_7897,N_9207);
nand UO_1465 (O_1465,N_9769,N_9783);
nand UO_1466 (O_1466,N_8096,N_8688);
nor UO_1467 (O_1467,N_9705,N_9647);
nand UO_1468 (O_1468,N_8600,N_8001);
and UO_1469 (O_1469,N_9352,N_9696);
nand UO_1470 (O_1470,N_7932,N_8335);
or UO_1471 (O_1471,N_8810,N_7968);
nand UO_1472 (O_1472,N_7664,N_9300);
nand UO_1473 (O_1473,N_9028,N_8001);
nor UO_1474 (O_1474,N_8548,N_8630);
nand UO_1475 (O_1475,N_8133,N_8950);
nor UO_1476 (O_1476,N_9465,N_8250);
nand UO_1477 (O_1477,N_8975,N_9717);
nand UO_1478 (O_1478,N_9977,N_7784);
nand UO_1479 (O_1479,N_8552,N_8771);
and UO_1480 (O_1480,N_7778,N_8461);
or UO_1481 (O_1481,N_9769,N_8838);
and UO_1482 (O_1482,N_8468,N_8028);
and UO_1483 (O_1483,N_9941,N_9359);
nand UO_1484 (O_1484,N_8830,N_8328);
nand UO_1485 (O_1485,N_8845,N_8930);
nor UO_1486 (O_1486,N_9299,N_8643);
nor UO_1487 (O_1487,N_9885,N_8539);
or UO_1488 (O_1488,N_9829,N_8961);
nand UO_1489 (O_1489,N_9297,N_8453);
or UO_1490 (O_1490,N_8317,N_9141);
and UO_1491 (O_1491,N_9711,N_8470);
or UO_1492 (O_1492,N_8442,N_7882);
nand UO_1493 (O_1493,N_7925,N_7738);
nand UO_1494 (O_1494,N_9522,N_7979);
or UO_1495 (O_1495,N_8455,N_7802);
nand UO_1496 (O_1496,N_9285,N_9414);
and UO_1497 (O_1497,N_9295,N_9742);
nor UO_1498 (O_1498,N_8248,N_9223);
nor UO_1499 (O_1499,N_8265,N_7894);
endmodule