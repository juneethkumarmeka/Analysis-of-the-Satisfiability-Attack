module basic_5000_50000_5000_50_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nand U0 (N_0,In_4023,In_4448);
or U1 (N_1,In_2399,In_1943);
or U2 (N_2,In_1221,In_2248);
and U3 (N_3,In_2470,In_1680);
nor U4 (N_4,In_3362,In_4796);
or U5 (N_5,In_35,In_1069);
nor U6 (N_6,In_2060,In_4325);
nand U7 (N_7,In_2245,In_1972);
nor U8 (N_8,In_4976,In_2390);
nor U9 (N_9,In_980,In_3083);
or U10 (N_10,In_2334,In_1116);
nand U11 (N_11,In_2154,In_850);
nor U12 (N_12,In_4447,In_2387);
xnor U13 (N_13,In_909,In_2364);
nand U14 (N_14,In_1510,In_3385);
nor U15 (N_15,In_4660,In_1306);
xor U16 (N_16,In_2478,In_203);
nor U17 (N_17,In_1840,In_2176);
and U18 (N_18,In_527,In_1173);
and U19 (N_19,In_4633,In_3842);
nor U20 (N_20,In_4729,In_3940);
nor U21 (N_21,In_207,In_4792);
or U22 (N_22,In_4133,In_3269);
nor U23 (N_23,In_4460,In_1531);
xor U24 (N_24,In_4743,In_795);
or U25 (N_25,In_3224,In_3790);
nand U26 (N_26,In_2772,In_2589);
xor U27 (N_27,In_4859,In_4140);
nand U28 (N_28,In_4569,In_962);
xor U29 (N_29,In_1697,In_1974);
nor U30 (N_30,In_2474,In_4587);
or U31 (N_31,In_4457,In_4258);
nor U32 (N_32,In_3204,In_907);
xnor U33 (N_33,In_2845,In_1477);
nor U34 (N_34,In_4229,In_1311);
nor U35 (N_35,In_3939,In_1548);
or U36 (N_36,In_3371,In_2183);
or U37 (N_37,In_1071,In_2613);
nand U38 (N_38,In_357,In_3636);
or U39 (N_39,In_2902,In_743);
or U40 (N_40,In_4402,In_3921);
and U41 (N_41,In_1616,In_4194);
nand U42 (N_42,In_4847,In_2750);
xnor U43 (N_43,In_2029,In_393);
and U44 (N_44,In_3581,In_2832);
nand U45 (N_45,In_1657,In_1091);
xnor U46 (N_46,In_3469,In_3446);
nor U47 (N_47,In_653,In_1471);
nand U48 (N_48,In_2409,In_275);
xor U49 (N_49,In_330,In_2538);
and U50 (N_50,In_564,In_2310);
nor U51 (N_51,In_934,In_4478);
nand U52 (N_52,In_3955,In_1379);
nor U53 (N_53,In_3756,In_4445);
xnor U54 (N_54,In_3030,In_2624);
nand U55 (N_55,In_2635,In_3085);
xnor U56 (N_56,In_4648,In_2304);
or U57 (N_57,In_591,In_2989);
nand U58 (N_58,In_4345,In_4008);
nand U59 (N_59,In_1220,In_4012);
nand U60 (N_60,In_4938,In_800);
or U61 (N_61,In_2629,In_4236);
and U62 (N_62,In_3867,In_2429);
xor U63 (N_63,In_1746,In_4499);
and U64 (N_64,In_3548,In_610);
nor U65 (N_65,In_1107,In_2526);
nand U66 (N_66,In_4339,In_1600);
nor U67 (N_67,In_3070,In_2214);
nor U68 (N_68,In_3065,In_3498);
nor U69 (N_69,In_2561,In_3615);
and U70 (N_70,In_1518,In_938);
or U71 (N_71,In_2567,In_3344);
nor U72 (N_72,In_183,In_2352);
or U73 (N_73,In_2256,In_2386);
nor U74 (N_74,In_2884,In_484);
nor U75 (N_75,In_4746,In_3494);
nor U76 (N_76,In_4466,In_4246);
nand U77 (N_77,In_2223,In_2863);
xor U78 (N_78,In_3832,In_4990);
and U79 (N_79,In_4241,In_4987);
nand U80 (N_80,In_530,In_3984);
nand U81 (N_81,In_170,In_620);
or U82 (N_82,In_173,In_186);
xor U83 (N_83,In_2554,In_4021);
xor U84 (N_84,In_2422,In_1060);
and U85 (N_85,In_3057,In_3052);
or U86 (N_86,In_4034,In_2228);
nor U87 (N_87,In_4252,In_4242);
or U88 (N_88,In_3364,In_3858);
and U89 (N_89,In_3338,In_4210);
or U90 (N_90,In_2405,In_331);
or U91 (N_91,In_231,In_640);
nand U92 (N_92,In_2499,In_4605);
nor U93 (N_93,In_210,In_3482);
nand U94 (N_94,In_1403,In_954);
and U95 (N_95,In_2141,In_178);
nor U96 (N_96,In_3692,In_3243);
or U97 (N_97,In_3035,In_3992);
nand U98 (N_98,In_3181,In_4579);
and U99 (N_99,In_3209,In_4738);
nand U100 (N_100,In_4393,In_4259);
nand U101 (N_101,In_2109,In_1268);
and U102 (N_102,In_3886,In_3399);
or U103 (N_103,In_288,In_1307);
xor U104 (N_104,In_433,In_2614);
nand U105 (N_105,In_4214,In_115);
nor U106 (N_106,In_3105,In_4476);
nand U107 (N_107,In_2047,In_1170);
and U108 (N_108,In_3782,In_2385);
nand U109 (N_109,In_2511,In_3848);
xor U110 (N_110,In_1519,In_619);
xor U111 (N_111,In_3409,In_3320);
nor U112 (N_112,In_4949,In_1997);
or U113 (N_113,In_4881,In_3899);
nand U114 (N_114,In_2115,In_2855);
xor U115 (N_115,In_2804,In_3542);
nor U116 (N_116,In_1289,In_2394);
nor U117 (N_117,In_3324,In_3936);
or U118 (N_118,In_3755,In_1290);
or U119 (N_119,In_2934,In_3720);
nand U120 (N_120,In_2320,In_1909);
xor U121 (N_121,In_1635,In_2257);
xnor U122 (N_122,In_2682,In_4335);
and U123 (N_123,In_628,In_2950);
nand U124 (N_124,In_2150,In_2790);
nand U125 (N_125,In_4737,In_1993);
xnor U126 (N_126,In_243,In_4365);
xnor U127 (N_127,In_117,In_3862);
and U128 (N_128,In_1467,In_2233);
xnor U129 (N_129,In_3563,In_1749);
and U130 (N_130,In_3981,In_4216);
and U131 (N_131,In_4040,In_4751);
nand U132 (N_132,In_3968,In_2264);
nor U133 (N_133,In_2292,In_3944);
and U134 (N_134,In_156,In_2846);
xnor U135 (N_135,In_595,In_1312);
and U136 (N_136,In_3217,In_2053);
and U137 (N_137,In_4652,In_1364);
xnor U138 (N_138,In_2945,In_461);
or U139 (N_139,In_1688,In_2737);
and U140 (N_140,In_603,In_617);
and U141 (N_141,In_580,In_1725);
xor U142 (N_142,In_3235,In_815);
xnor U143 (N_143,In_3343,In_404);
or U144 (N_144,In_2618,In_4718);
nor U145 (N_145,In_342,In_3810);
nand U146 (N_146,In_4344,In_1862);
xor U147 (N_147,In_4495,In_65);
nor U148 (N_148,In_2034,In_363);
xor U149 (N_149,In_1924,In_3174);
xnor U150 (N_150,In_3986,In_3258);
nor U151 (N_151,In_1250,In_2609);
nor U152 (N_152,In_1503,In_3716);
nand U153 (N_153,In_4189,In_3503);
nor U154 (N_154,In_4175,In_3547);
or U155 (N_155,In_996,In_1171);
nor U156 (N_156,In_1570,In_1131);
nor U157 (N_157,In_4653,In_1070);
or U158 (N_158,In_1959,In_1757);
and U159 (N_159,In_1406,In_4673);
nor U160 (N_160,In_859,In_1331);
and U161 (N_161,In_3046,In_1123);
or U162 (N_162,In_623,In_4692);
nor U163 (N_163,In_3643,In_3748);
or U164 (N_164,In_139,In_3207);
and U165 (N_165,In_3851,In_2717);
xor U166 (N_166,In_553,In_3613);
nand U167 (N_167,In_4015,In_1685);
nor U168 (N_168,In_1397,In_3397);
and U169 (N_169,In_2578,In_2254);
nor U170 (N_170,In_3496,In_2199);
nand U171 (N_171,In_974,In_3620);
xor U172 (N_172,In_2780,In_634);
or U173 (N_173,In_4665,In_1283);
xnor U174 (N_174,In_3987,In_1447);
nand U175 (N_175,In_1017,In_4176);
xnor U176 (N_176,In_2961,In_1217);
nor U177 (N_177,In_4109,In_1335);
or U178 (N_178,In_4994,In_3552);
nand U179 (N_179,In_939,In_4085);
and U180 (N_180,In_616,In_3737);
nor U181 (N_181,In_2755,In_2539);
xnor U182 (N_182,In_4999,In_1249);
or U183 (N_183,In_4761,In_626);
nand U184 (N_184,In_1555,In_625);
nor U185 (N_185,In_1147,In_3516);
nor U186 (N_186,In_1314,In_1229);
xnor U187 (N_187,In_4267,In_545);
nor U188 (N_188,In_3526,In_965);
and U189 (N_189,In_3917,In_4644);
or U190 (N_190,In_336,In_1851);
and U191 (N_191,In_2639,In_28);
nand U192 (N_192,In_2679,In_2419);
nand U193 (N_193,In_4060,In_2374);
or U194 (N_194,In_3771,In_1281);
or U195 (N_195,In_2827,In_2128);
or U196 (N_196,In_1969,In_985);
and U197 (N_197,In_1885,In_2496);
and U198 (N_198,In_4668,In_3360);
or U199 (N_199,In_720,In_57);
xor U200 (N_200,In_2032,In_2082);
and U201 (N_201,In_2423,In_4814);
nor U202 (N_202,In_2312,In_2500);
nand U203 (N_203,In_1489,In_507);
xnor U204 (N_204,In_4186,In_3798);
xor U205 (N_205,In_473,In_2503);
nand U206 (N_206,In_1549,In_3021);
xnor U207 (N_207,In_249,In_3830);
and U208 (N_208,In_1037,In_1243);
nor U209 (N_209,In_3437,In_892);
nor U210 (N_210,In_95,In_2987);
or U211 (N_211,In_3964,In_1636);
or U212 (N_212,In_1665,In_3127);
xor U213 (N_213,In_3805,In_4101);
or U214 (N_214,In_1910,In_2779);
nor U215 (N_215,In_3265,In_2046);
or U216 (N_216,In_1882,In_1753);
nor U217 (N_217,In_2074,In_3453);
and U218 (N_218,In_1563,In_3670);
and U219 (N_219,In_2709,In_926);
nand U220 (N_220,In_4563,In_3793);
or U221 (N_221,In_2969,In_2628);
and U222 (N_222,In_3017,In_3606);
nor U223 (N_223,In_4975,In_3892);
xnor U224 (N_224,In_1901,In_2973);
or U225 (N_225,In_1855,In_2145);
nand U226 (N_226,In_4209,In_3759);
xnor U227 (N_227,In_1423,In_4159);
or U228 (N_228,In_4177,In_2897);
nand U229 (N_229,In_1102,In_989);
and U230 (N_230,In_3534,In_4968);
nand U231 (N_231,In_3395,In_3504);
or U232 (N_232,In_4560,In_3704);
nand U233 (N_233,In_161,In_3998);
and U234 (N_234,In_1837,In_4360);
or U235 (N_235,In_1568,In_2163);
and U236 (N_236,In_882,In_2955);
and U237 (N_237,In_2565,In_3241);
nand U238 (N_238,In_3604,In_3567);
xnor U239 (N_239,In_4052,In_2105);
or U240 (N_240,In_2239,In_1767);
and U241 (N_241,In_2660,In_4399);
nor U242 (N_242,In_3172,In_3202);
and U243 (N_243,In_1922,In_4559);
and U244 (N_244,In_3531,In_4473);
or U245 (N_245,In_4786,In_284);
or U246 (N_246,In_1858,In_1968);
or U247 (N_247,In_2742,In_2446);
and U248 (N_248,In_2348,In_4157);
and U249 (N_249,In_74,In_2889);
nand U250 (N_250,In_2646,In_3304);
and U251 (N_251,In_4982,In_1611);
xor U252 (N_252,In_2625,In_4619);
nor U253 (N_253,In_4535,In_3432);
xor U254 (N_254,In_2774,In_3836);
nor U255 (N_255,In_108,In_1146);
xor U256 (N_256,In_3551,In_3633);
and U257 (N_257,In_495,In_63);
nand U258 (N_258,In_3835,In_3739);
xor U259 (N_259,In_2174,In_1230);
or U260 (N_260,In_344,In_3253);
nor U261 (N_261,In_2959,In_3513);
nand U262 (N_262,In_1770,In_2276);
nor U263 (N_263,In_3141,In_752);
nor U264 (N_264,In_3512,In_2021);
nand U265 (N_265,In_3777,In_438);
nor U266 (N_266,In_4725,In_563);
and U267 (N_267,In_1575,In_578);
or U268 (N_268,In_2020,In_596);
or U269 (N_269,In_2229,In_62);
nor U270 (N_270,In_1309,In_1906);
nand U271 (N_271,In_4863,In_2181);
xnor U272 (N_272,In_3530,In_2694);
and U273 (N_273,In_912,In_3452);
xor U274 (N_274,In_4519,In_3045);
nand U275 (N_275,In_2497,In_4921);
xnor U276 (N_276,In_4791,In_898);
xor U277 (N_277,In_4268,In_552);
and U278 (N_278,In_4285,In_4493);
and U279 (N_279,In_2842,In_3495);
or U280 (N_280,In_1743,In_3760);
xor U281 (N_281,In_4778,In_2549);
and U282 (N_282,In_152,In_787);
and U283 (N_283,In_1983,In_2017);
nand U284 (N_284,In_1584,In_4637);
or U285 (N_285,In_528,In_2358);
and U286 (N_286,In_3278,In_1917);
xor U287 (N_287,In_4527,In_3658);
xnor U288 (N_288,In_3322,In_3673);
or U289 (N_289,In_4817,In_592);
and U290 (N_290,In_2043,In_2913);
nor U291 (N_291,In_2761,In_1106);
and U292 (N_292,In_4542,In_2393);
xnor U293 (N_293,In_4699,In_2977);
or U294 (N_294,In_4632,In_4822);
and U295 (N_295,In_2070,In_82);
xor U296 (N_296,In_2805,In_2570);
or U297 (N_297,In_2551,In_3508);
xor U298 (N_298,In_128,In_4378);
or U299 (N_299,In_305,In_599);
and U300 (N_300,In_684,In_109);
or U301 (N_301,In_995,In_3525);
nand U302 (N_302,In_2990,In_784);
nand U303 (N_303,In_2739,In_1041);
nand U304 (N_304,In_4671,In_669);
and U305 (N_305,In_467,In_881);
nand U306 (N_306,In_455,In_4000);
nand U307 (N_307,In_4768,In_126);
xor U308 (N_308,In_940,In_4130);
xnor U309 (N_309,In_4301,In_3838);
nor U310 (N_310,In_4302,In_4931);
and U311 (N_311,In_1918,In_1165);
nand U312 (N_312,In_2548,In_3683);
and U313 (N_313,In_897,In_1682);
nand U314 (N_314,In_823,In_33);
xnor U315 (N_315,In_1588,In_2472);
nand U316 (N_316,In_1235,In_1145);
and U317 (N_317,In_4386,In_2330);
nand U318 (N_318,In_4150,In_2258);
or U319 (N_319,In_3655,In_761);
or U320 (N_320,In_4523,In_1092);
nor U321 (N_321,In_215,In_3979);
nor U322 (N_322,In_2930,In_2791);
nand U323 (N_323,In_4510,In_690);
and U324 (N_324,In_3303,In_4249);
and U325 (N_325,In_2674,In_321);
or U326 (N_326,In_4002,In_4405);
and U327 (N_327,In_42,In_749);
nor U328 (N_328,In_4414,In_1646);
nor U329 (N_329,In_4275,In_97);
or U330 (N_330,In_1552,In_4889);
xor U331 (N_331,In_1506,In_1088);
and U332 (N_332,In_85,In_3259);
and U333 (N_333,In_3069,In_2956);
xnor U334 (N_334,In_781,In_4962);
and U335 (N_335,In_4094,In_1940);
and U336 (N_336,In_8,In_2187);
and U337 (N_337,In_3593,In_2090);
xor U338 (N_338,In_2220,In_2061);
and U339 (N_339,In_4926,In_2958);
and U340 (N_340,In_1272,In_2058);
nor U341 (N_341,In_3292,In_1828);
nand U342 (N_342,In_3001,In_153);
nor U343 (N_343,In_1026,In_4946);
nand U344 (N_344,In_1315,In_2130);
xnor U345 (N_345,In_4811,In_2160);
and U346 (N_346,In_2180,In_833);
or U347 (N_347,In_4296,In_2974);
nand U348 (N_348,In_1726,In_3652);
nand U349 (N_349,In_1543,In_3485);
or U350 (N_350,In_2782,In_4907);
xor U351 (N_351,In_338,In_3162);
xor U352 (N_352,In_349,In_1606);
nor U353 (N_353,In_3691,In_3417);
or U354 (N_354,In_1777,In_3337);
nand U355 (N_355,In_3648,In_1354);
or U356 (N_356,In_3128,In_424);
or U357 (N_357,In_2366,In_2424);
or U358 (N_358,In_1532,In_4701);
and U359 (N_359,In_3428,In_3730);
nor U360 (N_360,In_4061,In_2408);
or U361 (N_361,In_4385,In_2718);
nand U362 (N_362,In_4440,In_3698);
xor U363 (N_363,In_2978,In_1556);
nand U364 (N_364,In_4888,In_510);
nand U365 (N_365,In_2313,In_3558);
or U366 (N_366,In_4276,In_4337);
nand U367 (N_367,In_4031,In_542);
nor U368 (N_368,In_1179,In_1167);
xnor U369 (N_369,In_2649,In_1948);
xor U370 (N_370,In_38,In_9);
nor U371 (N_371,In_1053,In_4058);
nor U372 (N_372,In_1628,In_3356);
nor U373 (N_373,In_4838,In_4369);
nor U374 (N_374,In_3455,In_2107);
or U375 (N_375,In_3628,In_4427);
nor U376 (N_376,In_612,In_947);
or U377 (N_377,In_796,In_3048);
nand U378 (N_378,In_4767,In_1202);
and U379 (N_379,In_4996,In_1946);
nor U380 (N_380,In_3837,In_1117);
or U381 (N_381,In_1133,In_2912);
nor U382 (N_382,In_1232,In_1476);
nand U383 (N_383,In_4118,In_2579);
or U384 (N_384,In_4721,In_4639);
and U385 (N_385,In_1027,In_2234);
nand U386 (N_386,In_1957,In_2170);
or U387 (N_387,In_4469,In_448);
or U388 (N_388,In_4145,In_537);
or U389 (N_389,In_1143,In_4240);
nand U390 (N_390,In_16,In_253);
nand U391 (N_391,In_1899,In_4954);
nand U392 (N_392,In_3664,In_858);
or U393 (N_393,In_3195,In_4465);
xor U394 (N_394,In_2415,In_2935);
nor U395 (N_395,In_1180,In_1747);
and U396 (N_396,In_34,In_301);
or U397 (N_397,In_3155,In_4195);
or U398 (N_398,In_2617,In_257);
and U399 (N_399,In_2018,In_1754);
nor U400 (N_400,In_751,In_638);
and U401 (N_401,In_3173,In_4022);
xor U402 (N_402,In_4463,In_1497);
nand U403 (N_403,In_1878,In_779);
nand U404 (N_404,In_3194,In_4797);
or U405 (N_405,In_3568,In_3486);
xnor U406 (N_406,In_3275,In_1595);
nand U407 (N_407,In_1648,In_1369);
xnor U408 (N_408,In_3123,In_3923);
nor U409 (N_409,In_67,In_1775);
nor U410 (N_410,In_4389,In_2230);
nor U411 (N_411,In_2598,In_2010);
xnor U412 (N_412,In_1293,In_1207);
and U413 (N_413,In_1010,In_482);
and U414 (N_414,In_392,In_3138);
nand U415 (N_415,In_1987,In_1008);
nor U416 (N_416,In_4269,In_4583);
xnor U417 (N_417,In_4849,In_4496);
or U418 (N_418,In_4902,In_4742);
or U419 (N_419,In_1119,In_2608);
nor U420 (N_420,In_138,In_1277);
or U421 (N_421,In_4215,In_1614);
nor U422 (N_422,In_1717,In_521);
nand U423 (N_423,In_1122,In_4411);
nand U424 (N_424,In_25,In_1100);
nor U425 (N_425,In_852,In_1561);
nand U426 (N_426,In_1325,In_1298);
and U427 (N_427,In_268,In_1134);
or U428 (N_428,In_2678,In_547);
nor U429 (N_429,In_4011,In_816);
nor U430 (N_430,In_343,In_3520);
or U431 (N_431,In_397,In_764);
xnor U432 (N_432,In_1615,In_2633);
nor U433 (N_433,In_4437,In_1474);
xor U434 (N_434,In_2916,In_355);
nand U435 (N_435,In_3796,In_2983);
nand U436 (N_436,In_3631,In_1154);
nor U437 (N_437,In_2114,In_1321);
and U438 (N_438,In_4409,In_1197);
or U439 (N_439,In_3521,In_1572);
xnor U440 (N_440,In_2896,In_3533);
nand U441 (N_441,In_4418,In_664);
nand U442 (N_442,In_2921,In_2789);
nor U443 (N_443,In_670,In_381);
nor U444 (N_444,In_2657,In_2477);
or U445 (N_445,In_2836,In_3477);
xor U446 (N_446,In_4073,In_1057);
or U447 (N_447,In_4037,In_799);
xnor U448 (N_448,In_2868,In_2926);
or U449 (N_449,In_2857,In_3640);
xnor U450 (N_450,In_2283,In_3646);
xor U451 (N_451,In_179,In_2568);
or U452 (N_452,In_4354,In_4691);
or U453 (N_453,In_4033,In_4831);
and U454 (N_454,In_883,In_925);
xnor U455 (N_455,In_4439,In_3822);
nand U456 (N_456,In_479,In_1334);
or U457 (N_457,In_1,In_3982);
nand U458 (N_458,In_59,In_4089);
and U459 (N_459,In_3843,In_4818);
or U460 (N_460,In_3367,In_747);
or U461 (N_461,In_1661,In_3994);
and U462 (N_462,In_1256,In_3676);
or U463 (N_463,In_4867,In_4205);
nand U464 (N_464,In_3348,In_2534);
and U465 (N_465,In_4969,In_1114);
or U466 (N_466,In_3497,In_1086);
and U467 (N_467,In_3560,In_2416);
or U468 (N_468,In_2373,In_4945);
nor U469 (N_469,In_4218,In_3727);
xor U470 (N_470,In_2049,In_141);
nor U471 (N_471,In_695,In_3200);
nand U472 (N_472,In_632,In_4840);
or U473 (N_473,In_3614,In_2778);
and U474 (N_474,In_4826,In_3970);
and U475 (N_475,In_2986,In_4076);
or U476 (N_476,In_3500,In_1536);
xor U477 (N_477,In_3925,In_233);
xor U478 (N_478,In_3783,In_2224);
xnor U479 (N_479,In_2997,In_683);
or U480 (N_480,In_1950,In_1149);
or U481 (N_481,In_2225,In_2980);
nand U482 (N_482,In_2807,In_529);
nand U483 (N_483,In_295,In_4942);
xor U484 (N_484,In_4048,In_147);
or U485 (N_485,In_2585,In_347);
nand U486 (N_486,In_4993,In_1527);
nor U487 (N_487,In_2166,In_23);
or U488 (N_488,In_1966,In_2489);
nor U489 (N_489,In_494,In_2108);
nand U490 (N_490,In_2361,In_4486);
nor U491 (N_491,In_2573,In_227);
or U492 (N_492,In_1675,In_586);
and U493 (N_493,In_3708,In_3487);
nand U494 (N_494,In_3059,In_4142);
or U495 (N_495,In_915,In_4717);
xnor U496 (N_496,In_333,In_636);
nor U497 (N_497,In_4425,In_4462);
or U498 (N_498,In_4041,In_3294);
or U499 (N_499,In_1720,In_3564);
nand U500 (N_500,In_2471,In_1356);
nor U501 (N_501,In_959,In_1514);
xnor U502 (N_502,In_575,In_1792);
or U503 (N_503,In_3430,In_1407);
and U504 (N_504,In_2445,In_255);
or U505 (N_505,In_630,In_474);
nand U506 (N_506,In_4715,In_2574);
nor U507 (N_507,In_990,In_2000);
nand U508 (N_508,In_4810,In_2533);
nand U509 (N_509,In_2915,In_4965);
and U510 (N_510,In_780,In_1327);
or U511 (N_511,In_3168,In_3869);
nand U512 (N_512,In_3185,In_4667);
xnor U513 (N_513,In_4050,In_1059);
xor U514 (N_514,In_1787,In_3119);
or U515 (N_515,In_4078,In_4524);
nor U516 (N_516,In_3330,In_1209);
nand U517 (N_517,In_871,In_4138);
or U518 (N_518,In_2865,In_4852);
or U519 (N_519,In_2881,In_3957);
or U520 (N_520,In_900,In_1935);
and U521 (N_521,In_4026,In_185);
or U522 (N_522,In_2748,In_76);
xor U523 (N_523,In_4117,In_1495);
nand U524 (N_524,In_4207,In_3107);
or U525 (N_525,In_2521,In_1558);
or U526 (N_526,In_2347,In_4063);
nor U527 (N_527,In_4179,In_4596);
nand U528 (N_528,In_1883,In_26);
nor U529 (N_529,In_3574,In_1623);
nand U530 (N_530,In_2133,In_2289);
xnor U531 (N_531,In_3177,In_2135);
xor U532 (N_532,In_2767,In_857);
or U533 (N_533,In_1694,In_125);
xnor U534 (N_534,In_92,In_677);
nand U535 (N_535,In_2508,In_1501);
nor U536 (N_536,In_237,In_3295);
nand U537 (N_537,In_4575,In_1727);
nor U538 (N_538,In_4707,In_4682);
nor U539 (N_539,In_3841,In_713);
nand U540 (N_540,In_2299,In_569);
or U541 (N_541,In_3008,In_2377);
nand U542 (N_542,In_150,In_3055);
or U543 (N_543,In_3301,In_4410);
and U544 (N_544,In_89,In_1206);
and U545 (N_545,In_557,In_4485);
nand U546 (N_546,In_2369,In_4772);
xor U547 (N_547,In_3493,In_3726);
xor U548 (N_548,In_860,In_902);
or U549 (N_549,In_2763,In_961);
nand U550 (N_550,In_1096,In_3819);
nor U551 (N_551,In_773,In_844);
xnor U552 (N_552,In_480,In_1005);
xor U553 (N_553,In_3511,In_1932);
nor U554 (N_554,In_1706,In_658);
xnor U555 (N_555,In_3199,In_2586);
nand U556 (N_556,In_3701,In_609);
or U557 (N_557,In_1319,In_2557);
nand U558 (N_558,In_4940,In_4517);
or U559 (N_559,In_4578,In_3038);
or U560 (N_560,In_4655,In_195);
nor U561 (N_561,In_1098,In_1827);
or U562 (N_562,In_4260,In_2713);
nand U563 (N_563,In_4766,In_1591);
xnor U564 (N_564,In_2077,In_223);
xor U565 (N_565,In_2901,In_4959);
nor U566 (N_566,In_3995,In_2644);
or U567 (N_567,In_2134,In_3668);
or U568 (N_568,In_3634,In_1819);
or U569 (N_569,In_1704,In_3281);
nor U570 (N_570,In_4158,In_368);
xor U571 (N_571,In_1362,In_4225);
and U572 (N_572,In_3018,In_4532);
nand U573 (N_573,In_4864,In_2452);
or U574 (N_574,In_309,In_3813);
and U575 (N_575,In_3596,In_4630);
nand U576 (N_576,In_3879,In_1265);
nor U577 (N_577,In_3966,In_2253);
and U578 (N_578,In_2363,In_308);
nor U579 (N_579,In_1211,In_2869);
or U580 (N_580,In_577,In_2685);
nand U581 (N_581,In_3074,In_4985);
nor U582 (N_582,In_3229,In_281);
xor U583 (N_583,In_4515,In_2443);
or U584 (N_584,In_514,In_407);
and U585 (N_585,In_1144,In_4839);
nand U586 (N_586,In_2498,In_1834);
nand U587 (N_587,In_420,In_3588);
xnor U588 (N_588,In_4776,In_1104);
and U589 (N_589,In_2421,In_4088);
xor U590 (N_590,In_3557,In_2431);
xor U591 (N_591,In_372,In_738);
and U592 (N_592,In_228,In_272);
nor U593 (N_593,In_2726,In_2116);
nand U594 (N_594,In_3027,In_4028);
or U595 (N_595,In_4357,In_3150);
and U596 (N_596,In_519,In_601);
or U597 (N_597,In_711,In_2417);
nor U598 (N_598,In_2206,In_2475);
xor U599 (N_599,In_2023,In_3930);
and U600 (N_600,In_2155,In_3456);
xnor U601 (N_601,In_4025,In_3143);
nand U602 (N_602,In_4310,In_1454);
and U603 (N_603,In_4873,In_2963);
or U604 (N_604,In_3422,In_2985);
nor U605 (N_605,In_730,In_2014);
nand U606 (N_606,In_4262,In_4533);
or U607 (N_607,In_3189,In_606);
or U608 (N_608,In_2904,In_1266);
or U609 (N_609,In_3806,In_496);
xnor U610 (N_610,In_2113,In_1234);
xnor U611 (N_611,In_2252,In_4657);
nand U612 (N_612,In_4509,In_4054);
or U613 (N_613,In_259,In_2825);
nand U614 (N_614,In_2542,In_1825);
xor U615 (N_615,In_2100,In_1835);
and U616 (N_616,In_4290,In_1358);
nand U617 (N_617,In_3461,In_1683);
nand U618 (N_618,In_3663,In_4212);
nor U619 (N_619,In_775,In_1587);
nand U620 (N_620,In_2714,In_188);
xnor U621 (N_621,In_3570,In_4016);
nor U622 (N_622,In_498,In_2964);
and U623 (N_623,In_3090,In_2208);
or U624 (N_624,In_1879,In_200);
nand U625 (N_625,In_250,In_2522);
and U626 (N_626,In_2880,In_2981);
xor U627 (N_627,In_4829,In_1748);
nor U628 (N_628,In_4607,In_3764);
or U629 (N_629,In_1003,In_4808);
and U630 (N_630,In_3616,In_1439);
nor U631 (N_631,In_341,In_2900);
nor U632 (N_632,In_4392,In_1077);
or U633 (N_633,In_3948,In_2516);
xor U634 (N_634,In_434,In_3678);
or U635 (N_635,In_376,In_4638);
nor U636 (N_636,In_4170,In_2623);
xor U637 (N_637,In_2878,In_4979);
nand U638 (N_638,In_3580,In_4317);
xor U639 (N_639,In_1426,In_1286);
or U640 (N_640,In_2177,In_3230);
or U641 (N_641,In_380,In_1547);
xor U642 (N_642,In_4238,In_908);
and U643 (N_643,In_4400,In_517);
or U644 (N_644,In_2595,In_3696);
and U645 (N_645,In_3945,In_2262);
nand U646 (N_646,In_2888,In_3778);
nand U647 (N_647,In_4745,In_4910);
and U648 (N_648,In_283,In_310);
and U649 (N_649,In_3478,In_1524);
nand U650 (N_650,In_4507,In_1006);
nand U651 (N_651,In_2126,In_2911);
nand U652 (N_652,In_1911,In_383);
and U653 (N_653,In_2341,In_957);
nand U654 (N_654,In_2059,In_270);
and U655 (N_655,In_4629,In_4421);
or U656 (N_656,In_1303,In_361);
or U657 (N_657,In_874,In_4067);
xor U658 (N_658,In_1864,In_1956);
xor U659 (N_659,In_73,In_3688);
or U660 (N_660,In_2441,In_2831);
nand U661 (N_661,In_1415,In_2757);
and U662 (N_662,In_388,In_3009);
and U663 (N_663,In_2502,In_337);
and U664 (N_664,In_2490,In_3388);
nand U665 (N_665,In_3167,In_4482);
xnor U666 (N_666,In_4373,In_3444);
xor U667 (N_667,In_1908,In_4464);
xor U668 (N_668,In_4628,In_1024);
nand U669 (N_669,In_866,In_3219);
nor U670 (N_670,In_4434,In_3523);
or U671 (N_671,In_4548,In_801);
nor U672 (N_672,In_3738,In_3942);
and U673 (N_673,In_4627,In_2270);
or U674 (N_674,In_4501,In_1046);
and U675 (N_675,In_3152,In_566);
nor U676 (N_676,In_2122,In_364);
nand U677 (N_677,In_1869,In_1094);
nor U678 (N_678,In_4143,In_3946);
or U679 (N_679,In_3321,In_721);
nor U680 (N_680,In_2687,In_2209);
nand U681 (N_681,In_3577,In_2575);
nand U682 (N_682,In_2263,In_1451);
nand U683 (N_683,In_1915,In_1581);
and U684 (N_684,In_199,In_375);
nand U685 (N_685,In_219,In_1464);
and U686 (N_686,In_4916,In_1544);
xor U687 (N_687,In_4760,In_4939);
nor U688 (N_688,In_1079,In_4227);
and U689 (N_689,In_802,In_1112);
xor U690 (N_690,In_457,In_3479);
or U691 (N_691,In_4570,In_704);
xnor U692 (N_692,In_373,In_825);
and U693 (N_693,In_136,In_1590);
nand U694 (N_694,In_2346,In_1498);
xnor U695 (N_695,In_2776,In_2792);
and U696 (N_696,In_1703,In_1631);
xnor U697 (N_697,In_1538,In_1928);
and U698 (N_698,In_2219,In_3111);
nor U699 (N_699,In_2661,In_4991);
xor U700 (N_700,In_1241,In_1388);
and U701 (N_701,In_4521,In_1845);
and U702 (N_702,In_572,In_2129);
and U703 (N_703,In_3250,In_861);
or U704 (N_704,In_3435,In_378);
and U705 (N_705,In_1607,In_4304);
and U706 (N_706,In_3073,In_3507);
or U707 (N_707,In_576,In_114);
nand U708 (N_708,In_3571,In_1773);
nand U709 (N_709,In_734,In_4273);
xor U710 (N_710,In_2432,In_4973);
nand U711 (N_711,In_2102,In_3585);
xnor U712 (N_712,In_4248,In_3876);
nor U713 (N_713,In_2716,In_54);
nand U714 (N_714,In_2221,In_3261);
and U715 (N_715,In_1420,In_3821);
or U716 (N_716,In_1264,In_2929);
xnor U717 (N_717,In_2928,In_278);
or U718 (N_718,In_1417,In_4773);
nand U719 (N_719,In_1019,In_429);
nor U720 (N_720,In_2652,In_1875);
or U721 (N_721,In_2291,In_3950);
and U722 (N_722,In_2924,In_69);
nand U723 (N_723,In_1301,In_2272);
or U724 (N_724,In_2351,In_2294);
nand U725 (N_725,In_1660,In_3784);
and U726 (N_726,In_4753,In_1789);
xor U727 (N_727,In_3402,In_741);
and U728 (N_728,In_1038,In_1267);
nor U729 (N_729,In_639,In_4292);
nor U730 (N_730,In_1353,In_2089);
nand U731 (N_731,In_1345,In_820);
or U732 (N_732,In_159,In_4804);
nor U733 (N_733,In_0,In_1986);
nor U734 (N_734,In_4219,In_2282);
nor U735 (N_735,In_2537,In_3887);
or U736 (N_736,In_4787,In_3618);
xor U737 (N_737,In_3084,In_3094);
or U738 (N_738,In_244,In_2430);
nor U739 (N_739,In_3905,In_29);
or U740 (N_740,In_4609,In_1372);
xnor U741 (N_741,In_1732,In_2406);
xnor U742 (N_742,In_960,In_4204);
and U743 (N_743,In_756,In_3377);
nor U744 (N_744,In_2201,In_2356);
nand U745 (N_745,In_700,In_1686);
xor U746 (N_746,In_2844,In_4862);
and U747 (N_747,In_4278,In_3963);
and U748 (N_748,In_3144,In_318);
nor U749 (N_749,In_1184,In_1594);
and U750 (N_750,In_408,In_4914);
or U751 (N_751,In_2597,In_2946);
xor U752 (N_752,In_4475,In_2698);
nor U753 (N_753,In_2922,In_4494);
nor U754 (N_754,In_1955,In_2465);
xor U755 (N_755,In_1651,In_1790);
xnor U756 (N_756,In_2188,In_1484);
and U757 (N_757,In_674,In_4762);
or U758 (N_758,In_1239,In_1148);
nor U759 (N_759,In_2035,In_4103);
nand U760 (N_760,In_4346,In_760);
xnor U761 (N_761,In_2893,In_2797);
nand U762 (N_762,In_2231,In_2079);
nor U763 (N_763,In_3514,In_4472);
nor U764 (N_764,In_762,In_2031);
nand U765 (N_765,In_3425,In_4305);
nor U766 (N_766,In_3319,In_2488);
or U767 (N_767,In_4740,In_826);
nor U768 (N_768,In_3136,In_3158);
nor U769 (N_769,In_719,In_1130);
or U770 (N_770,In_531,In_4963);
or U771 (N_771,In_2138,In_748);
nand U772 (N_772,In_1684,In_2607);
nand U773 (N_773,In_1516,In_3549);
or U774 (N_774,In_4315,In_835);
or U775 (N_775,In_2309,In_269);
or U776 (N_776,In_3365,In_587);
and U777 (N_777,In_1624,In_3392);
or U778 (N_778,In_3025,In_4953);
nor U779 (N_779,In_2664,In_1811);
or U780 (N_780,In_4126,In_4664);
nand U781 (N_781,In_4903,In_2464);
nand U782 (N_782,In_3179,In_405);
or U783 (N_783,In_266,In_2627);
or U784 (N_784,In_1210,In_1733);
nand U785 (N_785,In_4869,In_1437);
xor U786 (N_786,In_1049,In_2991);
xnor U787 (N_787,In_1689,In_123);
or U788 (N_788,In_3175,In_3491);
nand U789 (N_789,In_1813,In_4531);
nand U790 (N_790,In_4441,In_4280);
nand U791 (N_791,In_1701,In_4522);
nor U792 (N_792,In_2571,In_1296);
and U793 (N_793,In_30,In_3214);
or U794 (N_794,In_4952,In_2747);
or U795 (N_795,In_4880,In_1934);
xnor U796 (N_796,In_329,In_3579);
or U797 (N_797,In_2634,In_2011);
xor U798 (N_798,In_4358,In_3166);
nor U799 (N_799,In_1832,In_1801);
nor U800 (N_800,In_1389,In_265);
and U801 (N_801,In_1255,In_1893);
nand U802 (N_802,In_2295,In_2765);
and U803 (N_803,In_1759,In_4430);
or U804 (N_804,In_2708,In_4857);
or U805 (N_805,In_2012,In_3433);
nand U806 (N_806,In_1157,In_3731);
and U807 (N_807,In_1853,In_846);
nor U808 (N_808,In_3058,In_621);
nor U809 (N_809,In_2481,In_3140);
xor U810 (N_810,In_2411,In_2729);
nor U811 (N_811,In_3856,In_53);
or U812 (N_812,In_1346,In_1505);
and U813 (N_813,In_1347,In_1621);
or U814 (N_814,In_196,In_3104);
nand U815 (N_815,In_3161,In_546);
and U816 (N_816,In_1333,In_681);
xor U817 (N_817,In_3681,In_4468);
xor U818 (N_818,In_3576,In_2907);
nor U819 (N_819,In_80,In_3662);
or U820 (N_820,In_4536,In_3789);
or U821 (N_821,In_4898,In_4592);
nor U822 (N_822,In_1434,In_706);
xnor U823 (N_823,In_277,In_4771);
nand U824 (N_824,In_3116,In_3007);
nor U825 (N_825,In_2493,In_2454);
and U826 (N_826,In_4923,In_518);
nor U827 (N_827,In_718,In_27);
and U828 (N_828,In_44,In_2359);
or U829 (N_829,In_691,In_2322);
nor U830 (N_830,In_3232,In_4514);
and U831 (N_831,In_3770,In_1936);
and U832 (N_832,In_3993,In_4380);
nor U833 (N_833,In_2759,In_3222);
nand U834 (N_834,In_4970,In_4534);
or U835 (N_835,In_225,In_3375);
and U836 (N_836,In_4297,In_1463);
and U837 (N_837,In_1478,In_1338);
nor U838 (N_838,In_2494,In_2057);
or U839 (N_839,In_4634,In_4913);
nor U840 (N_840,In_923,In_1502);
nor U841 (N_841,In_3012,In_1742);
and U842 (N_842,In_2121,In_3752);
nor U843 (N_843,In_4622,In_699);
or U844 (N_844,In_3449,In_4169);
xor U845 (N_845,In_3325,In_4211);
nand U846 (N_846,In_3592,In_1557);
or U847 (N_847,In_2676,In_3927);
xnor U848 (N_848,In_4577,In_1343);
and U849 (N_849,In_3584,In_4049);
xnor U850 (N_850,In_948,In_289);
and U851 (N_851,In_4844,In_4858);
or U852 (N_852,In_1190,In_2783);
nor U853 (N_853,In_534,In_1838);
xnor U854 (N_854,In_3527,In_1473);
xnor U855 (N_855,In_1965,In_2384);
nor U856 (N_856,In_955,In_2051);
and U857 (N_857,In_60,In_1750);
nand U858 (N_858,In_2738,In_516);
nand U859 (N_859,In_590,In_4193);
nor U860 (N_860,In_1424,In_3715);
or U861 (N_861,In_3255,In_2864);
nand U862 (N_862,In_2487,In_3226);
xor U863 (N_863,In_951,In_742);
nand U864 (N_864,In_4500,In_3416);
or U865 (N_865,In_745,In_51);
xor U866 (N_866,In_3263,In_3541);
nand U867 (N_867,In_3900,In_4199);
nand U868 (N_868,In_1714,In_2119);
and U869 (N_869,In_2532,In_1652);
and U870 (N_870,In_4754,In_2327);
nor U871 (N_871,In_3180,In_1626);
xor U872 (N_872,In_3221,In_2288);
nor U873 (N_873,In_622,In_1921);
xor U874 (N_874,In_2169,In_3191);
xor U875 (N_875,In_4823,In_2655);
or U876 (N_876,In_998,In_581);
or U877 (N_877,In_3539,In_2479);
nand U878 (N_878,In_3949,In_2036);
and U879 (N_879,In_4313,In_1669);
nand U880 (N_880,In_4749,In_746);
nor U881 (N_881,In_582,In_3273);
nor U882 (N_882,In_3903,In_3674);
and U883 (N_883,In_444,In_2143);
xor U884 (N_884,In_3854,In_1080);
or U885 (N_885,In_1709,In_367);
xor U886 (N_886,In_4636,In_4384);
nand U887 (N_887,In_771,In_1674);
xnor U888 (N_888,In_2442,In_1392);
xnor U889 (N_889,In_1857,In_4178);
nand U890 (N_890,In_2232,In_94);
nand U891 (N_891,In_7,In_3318);
nand U892 (N_892,In_4528,In_4780);
xor U893 (N_893,In_4573,In_4890);
or U894 (N_894,In_2178,In_4735);
or U895 (N_895,In_4783,In_1492);
nor U896 (N_896,In_4068,In_1888);
xor U897 (N_897,In_2948,In_2005);
and U898 (N_898,In_1162,In_602);
nand U899 (N_899,In_4220,In_3501);
nand U900 (N_900,In_3724,In_856);
nor U901 (N_901,In_464,In_2601);
nand U902 (N_902,In_3352,In_3866);
nand U903 (N_903,In_3019,In_4336);
nor U904 (N_904,In_352,In_2541);
nor U905 (N_905,In_895,In_2426);
nor U906 (N_906,In_827,In_113);
xor U907 (N_907,In_1127,In_1018);
or U908 (N_908,In_2695,In_428);
nor U909 (N_909,In_2546,In_1933);
nor U910 (N_910,In_1200,In_4226);
xnor U911 (N_911,In_4723,In_3201);
nand U912 (N_912,In_2891,In_3280);
or U913 (N_913,In_991,In_371);
or U914 (N_914,In_1647,In_793);
and U915 (N_915,In_2569,In_379);
xnor U916 (N_916,In_3800,In_3205);
and U917 (N_917,In_4988,In_3355);
and U918 (N_918,In_4620,In_3244);
nor U919 (N_919,In_3227,In_2111);
nor U920 (N_920,In_4245,In_4454);
or U921 (N_921,In_2962,In_166);
and U922 (N_922,In_3718,In_43);
and U923 (N_923,In_3068,In_3543);
nand U924 (N_924,In_3812,In_1493);
nor U925 (N_925,In_4082,In_508);
and U926 (N_926,In_4332,In_1292);
nand U927 (N_927,In_292,In_3093);
xnor U928 (N_928,In_332,In_3575);
or U929 (N_929,In_2117,In_4989);
or U930 (N_930,In_983,In_3713);
nor U931 (N_931,In_441,In_4815);
nand U932 (N_932,In_659,In_1795);
nor U933 (N_933,In_3170,In_2159);
and U934 (N_934,In_4974,In_4918);
xor U935 (N_935,In_1755,In_2843);
or U936 (N_936,In_631,In_1422);
nor U937 (N_937,In_3300,In_2787);
and U938 (N_938,In_2545,In_487);
nand U939 (N_939,In_322,In_4353);
and U940 (N_940,In_4003,In_1638);
and U941 (N_941,In_2202,In_4153);
nand U942 (N_942,In_1452,In_1259);
xnor U943 (N_943,In_2458,In_4470);
or U944 (N_944,In_2319,In_3290);
nand U945 (N_945,In_2547,In_184);
xor U946 (N_946,In_2999,In_4901);
xor U947 (N_947,In_1964,In_4111);
xor U948 (N_948,In_971,In_2918);
xor U949 (N_949,In_2298,In_2467);
or U950 (N_950,In_513,In_1215);
xor U951 (N_951,In_4618,In_2081);
xnor U952 (N_952,In_2673,In_2087);
xnor U953 (N_953,In_1960,In_4825);
nor U954 (N_954,In_1654,In_328);
or U955 (N_955,In_1208,In_500);
and U956 (N_956,In_4398,In_1592);
and U957 (N_957,In_2274,In_3814);
or U958 (N_958,In_4144,In_4306);
and U959 (N_959,In_4412,In_2275);
nand U960 (N_960,In_4413,In_1199);
xor U961 (N_961,In_1831,In_3036);
or U962 (N_962,In_451,In_1978);
nand U963 (N_963,In_133,In_2982);
xnor U964 (N_964,In_3404,In_2383);
or U965 (N_965,In_3476,In_2872);
or U966 (N_966,In_4005,In_4802);
or U967 (N_967,In_470,In_187);
xnor U968 (N_968,In_4104,In_3834);
and U969 (N_969,In_3096,In_2267);
or U970 (N_970,In_1938,In_3287);
and U971 (N_971,In_202,In_2942);
and U972 (N_972,In_1262,In_1291);
nand U973 (N_973,In_2297,In_3298);
xnor U974 (N_974,In_4066,In_1330);
nor U975 (N_975,In_4925,In_3171);
nand U976 (N_976,In_2684,In_1810);
or U977 (N_977,In_4719,In_2173);
or U978 (N_978,In_2103,In_389);
nor U979 (N_979,In_476,In_600);
and U980 (N_980,In_3928,In_665);
nand U981 (N_981,In_688,In_4567);
or U982 (N_982,In_4239,In_22);
or U983 (N_983,In_2434,In_1336);
or U984 (N_984,In_3550,In_1895);
nor U985 (N_985,In_1168,In_4803);
nor U986 (N_986,In_2505,In_1342);
nor U987 (N_987,In_3918,In_1023);
or U988 (N_988,In_2142,In_515);
nor U989 (N_989,In_3100,In_4631);
nor U990 (N_990,In_3153,In_3561);
nand U991 (N_991,In_3751,In_2697);
or U992 (N_992,In_1981,In_2834);
xor U993 (N_993,In_4449,In_1944);
or U994 (N_994,In_4821,In_1541);
or U995 (N_995,In_3828,In_104);
nor U996 (N_996,In_78,In_1876);
nor U997 (N_997,In_1873,In_2576);
nor U998 (N_998,In_1063,In_2951);
xnor U999 (N_999,In_458,In_20);
and U1000 (N_1000,N_527,In_1378);
and U1001 (N_1001,N_307,N_655);
or U1002 (N_1002,In_143,In_2833);
xor U1003 (N_1003,In_4656,In_3573);
or U1004 (N_1004,N_6,N_219);
or U1005 (N_1005,In_2631,In_2786);
xor U1006 (N_1006,In_2839,In_87);
nor U1007 (N_1007,In_2371,In_941);
xnor U1008 (N_1008,N_640,In_1438);
xnor U1009 (N_1009,N_672,In_2317);
nand U1010 (N_1010,N_153,In_4255);
xnor U1011 (N_1011,In_1779,In_1166);
nor U1012 (N_1012,In_2611,In_1185);
nor U1013 (N_1013,In_1128,In_2810);
nor U1014 (N_1014,In_230,In_1115);
xnor U1015 (N_1015,N_190,N_616);
or U1016 (N_1016,In_4237,In_3914);
and U1017 (N_1017,In_1441,N_856);
and U1018 (N_1018,In_1399,In_2457);
or U1019 (N_1019,In_2688,In_3882);
or U1020 (N_1020,In_2453,In_2604);
xor U1021 (N_1021,In_1530,In_3427);
and U1022 (N_1022,N_209,In_180);
xnor U1023 (N_1023,In_3931,In_2391);
nand U1024 (N_1024,N_455,In_1650);
xnor U1025 (N_1025,In_4489,N_124);
or U1026 (N_1026,In_2853,N_269);
and U1027 (N_1027,In_3736,In_1515);
and U1028 (N_1028,In_3299,In_449);
and U1029 (N_1029,In_570,In_4446);
nor U1030 (N_1030,N_955,N_531);
nand U1031 (N_1031,In_789,N_709);
xnor U1032 (N_1032,In_416,In_2886);
nor U1033 (N_1033,In_2360,In_2849);
nor U1034 (N_1034,In_417,N_397);
nand U1035 (N_1035,N_932,In_1176);
xnor U1036 (N_1036,In_4147,In_3599);
and U1037 (N_1037,In_2563,N_923);
or U1038 (N_1038,In_661,In_807);
nor U1039 (N_1039,In_2146,In_302);
nor U1040 (N_1040,In_556,In_4328);
nand U1041 (N_1041,In_4093,In_158);
or U1042 (N_1042,In_3684,In_837);
and U1043 (N_1043,In_944,In_1337);
and U1044 (N_1044,N_907,N_113);
and U1045 (N_1045,In_4467,In_2727);
and U1046 (N_1046,In_2734,In_3601);
xnor U1047 (N_1047,In_759,In_3883);
nor U1048 (N_1048,In_4243,N_440);
xnor U1049 (N_1049,In_3457,In_4213);
nand U1050 (N_1050,N_93,In_4192);
xor U1051 (N_1051,In_3654,N_964);
xnor U1052 (N_1052,In_3792,N_39);
xor U1053 (N_1053,In_3605,N_881);
and U1054 (N_1054,In_4474,N_811);
or U1055 (N_1055,In_662,In_1812);
nand U1056 (N_1056,In_1328,In_1559);
nor U1057 (N_1057,In_154,In_37);
xor U1058 (N_1058,In_1798,N_456);
or U1059 (N_1059,In_627,N_88);
and U1060 (N_1060,In_3407,In_4750);
nor U1061 (N_1061,In_3536,In_3438);
nor U1062 (N_1062,N_216,N_719);
or U1063 (N_1063,N_762,In_4348);
or U1064 (N_1064,In_554,N_419);
or U1065 (N_1065,N_538,In_4057);
nor U1066 (N_1066,N_847,In_2529);
nand U1067 (N_1067,N_780,In_2998);
xor U1068 (N_1068,In_1445,In_4404);
nand U1069 (N_1069,In_2015,In_1487);
or U1070 (N_1070,N_497,In_2340);
or U1071 (N_1071,In_400,In_1485);
and U1072 (N_1072,In_783,In_1566);
xnor U1073 (N_1073,In_1460,In_1160);
and U1074 (N_1074,In_3983,In_698);
or U1075 (N_1075,In_1310,In_4621);
and U1076 (N_1076,In_1877,N_742);
nand U1077 (N_1077,In_663,In_1368);
and U1078 (N_1078,In_3872,In_144);
and U1079 (N_1079,In_2544,In_3260);
or U1080 (N_1080,N_810,In_2450);
nor U1081 (N_1081,In_2515,N_250);
nand U1082 (N_1082,In_1520,N_976);
nand U1083 (N_1083,In_2016,N_974);
nand U1084 (N_1084,In_2581,N_169);
xnor U1085 (N_1085,N_750,N_155);
or U1086 (N_1086,N_90,N_673);
nand U1087 (N_1087,In_4505,N_801);
nand U1088 (N_1088,In_3623,N_692);
xor U1089 (N_1089,In_3028,N_574);
nor U1090 (N_1090,N_122,In_849);
nand U1091 (N_1091,In_1085,In_1048);
nor U1092 (N_1092,N_592,In_1045);
nand U1093 (N_1093,In_2979,In_1137);
xor U1094 (N_1094,In_3878,In_1737);
nor U1095 (N_1095,In_696,N_466);
nand U1096 (N_1096,In_252,In_3370);
or U1097 (N_1097,In_4502,In_2837);
nor U1098 (N_1098,In_2268,In_1011);
nand U1099 (N_1099,In_920,In_3003);
nor U1100 (N_1100,N_464,In_2476);
xor U1101 (N_1101,In_3092,In_1796);
or U1102 (N_1102,N_959,In_2645);
and U1103 (N_1103,N_285,In_1700);
nor U1104 (N_1104,N_520,In_2044);
nand U1105 (N_1105,In_3728,In_3729);
nor U1106 (N_1106,N_436,In_239);
or U1107 (N_1107,In_345,In_1545);
and U1108 (N_1108,In_647,In_2491);
or U1109 (N_1109,In_608,N_559);
xor U1110 (N_1110,In_2504,In_3602);
nor U1111 (N_1111,In_1850,In_1824);
nor U1112 (N_1112,In_1715,In_1341);
or U1113 (N_1113,In_1078,In_1248);
or U1114 (N_1114,In_2302,In_2048);
and U1115 (N_1115,In_4643,In_4540);
xnor U1116 (N_1116,N_805,In_4900);
or U1117 (N_1117,N_532,N_808);
or U1118 (N_1118,In_1126,In_1317);
nor U1119 (N_1119,N_611,N_568);
and U1120 (N_1120,In_573,In_3908);
or U1121 (N_1121,N_385,In_1678);
xnor U1122 (N_1122,In_4429,In_1867);
and U1123 (N_1123,N_885,N_373);
nand U1124 (N_1124,N_546,N_913);
nand U1125 (N_1125,In_884,In_4294);
nand U1126 (N_1126,In_1761,N_984);
xnor U1127 (N_1127,In_682,In_851);
or U1128 (N_1128,N_933,In_4820);
and U1129 (N_1129,In_4891,In_1025);
nand U1130 (N_1130,N_60,In_151);
or U1131 (N_1131,In_4388,In_267);
nor U1132 (N_1132,In_3657,N_499);
nand U1133 (N_1133,N_380,In_1847);
xnor U1134 (N_1134,In_351,N_96);
xnor U1135 (N_1135,In_4027,In_932);
nand U1136 (N_1136,In_3305,In_2894);
nor U1137 (N_1137,N_752,In_558);
nor U1138 (N_1138,In_1673,In_949);
nand U1139 (N_1139,In_4289,In_3022);
and U1140 (N_1140,In_3125,In_45);
or U1141 (N_1141,In_4125,N_601);
nand U1142 (N_1142,In_2378,In_1695);
and U1143 (N_1143,N_235,N_165);
nand U1144 (N_1144,In_4708,N_251);
xor U1145 (N_1145,In_1995,In_3441);
and U1146 (N_1146,In_472,N_883);
nor U1147 (N_1147,In_817,In_1132);
nor U1148 (N_1148,In_4435,N_144);
or U1149 (N_1149,In_1462,In_2485);
nand U1150 (N_1150,N_143,In_2943);
or U1151 (N_1151,In_4964,In_2892);
xor U1152 (N_1152,In_4883,In_3975);
or U1153 (N_1153,N_706,In_2899);
nor U1154 (N_1154,In_4616,In_1870);
and U1155 (N_1155,N_308,N_733);
nor U1156 (N_1156,N_320,In_263);
nor U1157 (N_1157,N_569,In_2731);
or U1158 (N_1158,In_685,N_596);
nor U1159 (N_1159,N_189,N_431);
nand U1160 (N_1160,N_214,In_1138);
and U1161 (N_1161,N_51,In_3288);
nor U1162 (N_1162,In_4298,In_1366);
nand U1163 (N_1163,In_2156,In_4247);
or U1164 (N_1164,In_3972,In_3060);
xnor U1165 (N_1165,In_2610,In_1409);
or U1166 (N_1166,In_1348,N_316);
nand U1167 (N_1167,In_4574,In_1039);
or U1168 (N_1168,In_120,N_184);
nand U1169 (N_1169,In_1990,In_3124);
and U1170 (N_1170,In_1550,In_293);
xnor U1171 (N_1171,N_712,In_2802);
nor U1172 (N_1172,In_3985,In_3667);
nand U1173 (N_1173,In_1735,In_235);
and U1174 (N_1174,N_727,N_880);
xor U1175 (N_1175,In_1365,In_93);
nor U1176 (N_1176,In_1554,N_852);
nor U1177 (N_1177,In_1391,N_5);
xor U1178 (N_1178,In_218,N_409);
xor U1179 (N_1179,In_1939,In_924);
and U1180 (N_1180,In_1486,N_340);
nand U1181 (N_1181,In_3907,In_421);
xor U1182 (N_1182,In_1431,In_3988);
and U1183 (N_1183,N_44,In_968);
nand U1184 (N_1184,In_4915,In_1984);
xor U1185 (N_1185,N_25,In_299);
nor U1186 (N_1186,N_998,N_840);
xor U1187 (N_1187,In_3653,In_735);
and U1188 (N_1188,In_3359,In_459);
nor U1189 (N_1189,In_728,In_1930);
and U1190 (N_1190,N_481,In_3795);
nand U1191 (N_1191,In_1393,In_317);
and U1192 (N_1192,In_3874,In_2939);
and U1193 (N_1193,N_820,In_4650);
nand U1194 (N_1194,N_943,In_4283);
and U1195 (N_1195,N_675,In_3387);
or U1196 (N_1196,In_3974,In_4805);
and U1197 (N_1197,In_4264,In_1618);
nor U1198 (N_1198,N_106,In_2191);
nand U1199 (N_1199,In_1730,In_486);
and U1200 (N_1200,In_2720,N_685);
nor U1201 (N_1201,In_2518,In_2462);
xnor U1202 (N_1202,In_1305,In_2413);
nor U1203 (N_1203,In_1040,In_2062);
nor U1204 (N_1204,In_242,In_3742);
nand U1205 (N_1205,In_3953,In_1054);
or U1206 (N_1206,In_4543,N_570);
nor U1207 (N_1207,N_595,In_145);
xnor U1208 (N_1208,In_2344,In_524);
xor U1209 (N_1209,In_4001,In_611);
or U1210 (N_1210,In_370,N_565);
xor U1211 (N_1211,In_2510,N_662);
nor U1212 (N_1212,N_54,In_1419);
xor U1213 (N_1213,N_857,In_4978);
and U1214 (N_1214,In_137,In_3350);
nor U1215 (N_1215,N_623,In_776);
and U1216 (N_1216,N_364,N_507);
nor U1217 (N_1217,N_3,In_4045);
or U1218 (N_1218,N_687,In_4758);
and U1219 (N_1219,In_2553,In_568);
nor U1220 (N_1220,N_295,In_3089);
nor U1221 (N_1221,In_4784,N_748);
xnor U1222 (N_1222,In_2088,In_414);
xor U1223 (N_1223,In_50,In_2022);
nand U1224 (N_1224,N_954,In_4702);
or U1225 (N_1225,N_916,N_107);
xor U1226 (N_1226,In_593,In_3372);
nor U1227 (N_1227,N_294,In_3458);
or U1228 (N_1228,In_4106,In_1028);
nor U1229 (N_1229,In_1380,In_1302);
nand U1230 (N_1230,In_4600,In_297);
xor U1231 (N_1231,In_49,In_1427);
xnor U1232 (N_1232,N_23,N_521);
nand U1233 (N_1233,In_4261,In_2392);
nand U1234 (N_1234,In_1808,In_1370);
nor U1235 (N_1235,N_783,In_4);
nand U1236 (N_1236,N_690,In_3656);
and U1237 (N_1237,N_550,N_383);
xor U1238 (N_1238,In_103,N_65);
and U1239 (N_1239,In_2195,In_2751);
xnor U1240 (N_1240,In_3894,In_2817);
nand U1241 (N_1241,In_3245,In_1705);
xnor U1242 (N_1242,In_4403,N_560);
and U1243 (N_1243,In_1108,N_183);
nor U1244 (N_1244,N_966,In_1072);
and U1245 (N_1245,In_3316,In_2153);
or U1246 (N_1246,In_3888,In_1999);
nand U1247 (N_1247,In_2861,In_1030);
and U1248 (N_1248,N_819,In_4617);
xnor U1249 (N_1249,N_254,In_499);
nor U1250 (N_1250,In_3638,In_2279);
nor U1251 (N_1251,N_127,In_4576);
nand U1252 (N_1252,In_1067,In_2743);
and U1253 (N_1253,In_3031,In_2281);
xnor U1254 (N_1254,In_3345,In_2650);
or U1255 (N_1255,In_306,In_2562);
xnor U1256 (N_1256,In_1785,N_779);
or U1257 (N_1257,In_4056,In_251);
nand U1258 (N_1258,In_1976,In_3612);
xnor U1259 (N_1259,In_929,In_2512);
and U1260 (N_1260,N_32,In_2306);
nand U1261 (N_1261,In_2075,N_563);
nor U1262 (N_1262,In_4308,N_835);
and U1263 (N_1263,In_765,In_3234);
nand U1264 (N_1264,In_2067,In_1639);
or U1265 (N_1265,N_602,In_2455);
nand U1266 (N_1266,In_2486,In_1124);
and U1267 (N_1267,N_248,N_704);
nor U1268 (N_1268,In_2397,In_4366);
xnor U1269 (N_1269,In_1905,In_411);
or U1270 (N_1270,In_189,In_2919);
and U1271 (N_1271,In_340,In_171);
nor U1272 (N_1272,In_1820,In_3611);
xnor U1273 (N_1273,N_937,N_628);
and U1274 (N_1274,In_1711,In_705);
nand U1275 (N_1275,In_676,N_141);
and U1276 (N_1276,N_781,In_4957);
and U1277 (N_1277,In_4998,In_1136);
or U1278 (N_1278,In_4137,In_2923);
and U1279 (N_1279,In_935,N_751);
nand U1280 (N_1280,N_629,N_961);
and U1281 (N_1281,N_757,In_2396);
or U1282 (N_1282,In_4173,In_769);
nand U1283 (N_1283,N_161,In_3881);
xnor U1284 (N_1284,In_644,In_3473);
nand U1285 (N_1285,N_555,In_943);
xor U1286 (N_1286,N_731,In_2732);
or U1287 (N_1287,In_116,In_81);
xnor U1288 (N_1288,In_1055,N_989);
or U1289 (N_1289,In_11,In_1523);
or U1290 (N_1290,In_2866,In_4124);
nor U1291 (N_1291,In_129,In_880);
nor U1292 (N_1292,In_100,In_565);
nor U1293 (N_1293,N_30,In_3271);
xor U1294 (N_1294,In_1082,In_236);
xnor U1295 (N_1295,In_3340,N_562);
xor U1296 (N_1296,In_1951,In_492);
and U1297 (N_1297,In_1926,In_813);
nand U1298 (N_1298,In_4709,In_1152);
or U1299 (N_1299,N_771,In_4554);
xor U1300 (N_1300,In_1201,In_1142);
or U1301 (N_1301,N_583,In_3266);
or U1302 (N_1302,N_505,N_558);
and U1303 (N_1303,In_2095,In_641);
nand U1304 (N_1304,In_386,N_667);
nor U1305 (N_1305,In_4168,In_2640);
nand U1306 (N_1306,In_4782,N_877);
nor U1307 (N_1307,In_2085,N_809);
nor U1308 (N_1308,N_10,In_656);
xor U1309 (N_1309,In_2580,In_3064);
xnor U1310 (N_1310,In_1821,In_2278);
or U1311 (N_1311,In_456,In_4908);
nor U1312 (N_1312,N_18,In_1799);
or U1313 (N_1313,N_914,In_3218);
xor U1314 (N_1314,In_736,In_1450);
or U1315 (N_1315,In_4417,In_4334);
xnor U1316 (N_1316,In_1394,In_1833);
nor U1317 (N_1317,N_174,In_4871);
nor U1318 (N_1318,In_1195,In_1871);
xnor U1319 (N_1319,In_3368,In_271);
nand U1320 (N_1320,In_1852,In_4611);
and U1321 (N_1321,In_3831,In_1823);
nand U1322 (N_1322,In_3246,In_1672);
and U1323 (N_1323,In_770,In_585);
xor U1324 (N_1324,In_3208,In_2577);
nor U1325 (N_1325,In_4490,N_747);
nand U1326 (N_1326,In_3098,In_3423);
nand U1327 (N_1327,In_4079,In_1880);
nor U1328 (N_1328,N_561,In_3697);
and U1329 (N_1329,N_357,In_325);
nor U1330 (N_1330,In_2314,In_4895);
xor U1331 (N_1331,In_2995,N_607);
or U1332 (N_1332,In_3797,In_1500);
or U1333 (N_1333,In_4042,In_2401);
and U1334 (N_1334,In_4597,In_1181);
or U1335 (N_1335,In_2840,N_305);
nand U1336 (N_1336,In_3470,In_4842);
nand U1337 (N_1337,In_3460,In_1535);
nand U1338 (N_1338,In_70,In_3791);
nand U1339 (N_1339,In_319,In_1095);
and U1340 (N_1340,In_3582,In_3706);
nor U1341 (N_1341,In_2096,In_2637);
xnor U1342 (N_1342,In_2910,In_906);
nor U1343 (N_1343,N_591,In_1402);
and U1344 (N_1344,N_797,In_4539);
nand U1345 (N_1345,N_59,In_4947);
and U1346 (N_1346,In_4770,In_4161);
or U1347 (N_1347,In_3565,N_547);
or U1348 (N_1348,N_231,In_320);
nor U1349 (N_1349,In_4674,N_256);
or U1350 (N_1350,N_82,N_898);
xnor U1351 (N_1351,In_4967,In_1349);
nor U1352 (N_1352,In_4550,In_4662);
nand U1353 (N_1353,In_4491,In_3313);
xor U1354 (N_1354,N_130,In_1350);
nand U1355 (N_1355,In_3213,In_4039);
nand U1356 (N_1356,In_4557,In_3391);
or U1357 (N_1357,In_2204,In_2859);
or U1358 (N_1358,N_921,In_4135);
nand U1359 (N_1359,In_3117,In_3562);
or U1360 (N_1360,In_1603,In_2324);
nor U1361 (N_1361,In_1947,In_1446);
nor U1362 (N_1362,N_730,N_872);
xnor U1363 (N_1363,In_4906,In_4983);
or U1364 (N_1364,In_3609,In_589);
and U1365 (N_1365,N_273,In_1942);
nor U1366 (N_1366,N_416,In_3076);
xor U1367 (N_1367,In_4424,N_228);
nor U1368 (N_1368,N_633,In_286);
and U1369 (N_1369,In_1783,In_2954);
nor U1370 (N_1370,In_88,In_3133);
xnor U1371 (N_1371,In_3544,In_3846);
or U1372 (N_1372,N_879,In_2781);
and U1373 (N_1373,In_3312,In_3956);
and U1374 (N_1374,In_369,In_1533);
xnor U1375 (N_1375,In_594,In_4253);
xor U1376 (N_1376,In_2572,In_1769);
nand U1377 (N_1377,In_3711,N_545);
nor U1378 (N_1378,N_405,In_3489);
nand U1379 (N_1379,In_4009,In_1756);
xnor U1380 (N_1380,In_2704,In_4316);
and U1381 (N_1381,In_475,N_834);
xnor U1382 (N_1382,N_996,N_204);
nand U1383 (N_1383,N_571,In_1881);
and U1384 (N_1384,In_3033,N_417);
nand U1385 (N_1385,In_1270,In_1308);
nand U1386 (N_1386,In_2337,In_2860);
nor U1387 (N_1387,In_4256,In_2139);
xor U1388 (N_1388,N_420,N_206);
or U1389 (N_1389,N_516,N_679);
nor U1390 (N_1390,In_2045,In_613);
and U1391 (N_1391,In_4565,In_4703);
nor U1392 (N_1392,N_803,In_1585);
and U1393 (N_1393,In_1499,N_551);
nor U1394 (N_1394,In_1919,N_999);
nor U1395 (N_1395,In_1352,In_1194);
nor U1396 (N_1396,In_4588,N_215);
xnor U1397 (N_1397,In_4764,In_3649);
xor U1398 (N_1398,In_1158,In_3398);
nor U1399 (N_1399,N_586,In_3211);
xor U1400 (N_1400,In_387,N_718);
nor U1401 (N_1401,In_18,N_37);
nor U1402 (N_1402,In_3677,In_3624);
nand U1403 (N_1403,In_701,In_2395);
and U1404 (N_1404,N_399,N_537);
nor U1405 (N_1405,In_4363,In_913);
nor U1406 (N_1406,In_463,In_4508);
nor U1407 (N_1407,In_4875,In_4984);
nor U1408 (N_1408,In_3323,In_4571);
xnor U1409 (N_1409,In_4487,In_2600);
nand U1410 (N_1410,In_1288,N_864);
nor U1411 (N_1411,In_928,In_356);
nor U1412 (N_1412,In_4171,In_3559);
or U1413 (N_1413,In_1929,In_3590);
and U1414 (N_1414,In_276,In_3754);
or U1415 (N_1415,In_1562,N_787);
nand U1416 (N_1416,N_928,In_4059);
nor U1417 (N_1417,N_263,In_4928);
and U1418 (N_1418,In_1483,In_3447);
and U1419 (N_1419,N_140,In_4733);
nor U1420 (N_1420,In_3091,In_2466);
xor U1421 (N_1421,In_4228,In_3965);
or U1422 (N_1422,In_4309,In_1465);
nand U1423 (N_1423,In_4443,N_151);
or U1424 (N_1424,N_297,In_3426);
and U1425 (N_1425,N_300,In_3522);
and U1426 (N_1426,In_3000,In_2632);
or U1427 (N_1427,N_776,In_3190);
xor U1428 (N_1428,N_985,N_175);
xnor U1429 (N_1429,In_4511,In_3935);
xor U1430 (N_1430,In_3617,In_4156);
and U1431 (N_1431,In_4134,In_2813);
nand U1432 (N_1432,In_1625,N_888);
or U1433 (N_1433,In_4422,In_1892);
and U1434 (N_1434,In_1219,In_1036);
nor U1435 (N_1435,In_2265,In_4484);
xnor U1436 (N_1436,In_645,In_4795);
or U1437 (N_1437,N_965,In_1613);
and U1438 (N_1438,In_3644,In_2728);
and U1439 (N_1439,In_2418,In_31);
and U1440 (N_1440,In_2941,N_262);
nor U1441 (N_1441,In_2131,In_2593);
nand U1442 (N_1442,In_3101,In_4912);
or U1443 (N_1443,In_3619,In_1630);
and U1444 (N_1444,In_4364,In_1914);
or U1445 (N_1445,In_2994,In_4165);
xnor U1446 (N_1446,In_1610,In_649);
xor U1447 (N_1447,N_8,In_2460);
or U1448 (N_1448,In_1509,In_3901);
nand U1449 (N_1449,N_56,In_1470);
or U1450 (N_1450,In_4566,In_966);
nor U1451 (N_1451,In_3445,In_2469);
nand U1452 (N_1452,In_1593,In_1836);
xnor U1453 (N_1453,In_2144,N_387);
nand U1454 (N_1454,In_1375,In_2350);
or U1455 (N_1455,In_4459,In_262);
and U1456 (N_1456,N_170,In_2883);
and U1457 (N_1457,N_353,In_3741);
or U1458 (N_1458,N_275,In_3198);
and U1459 (N_1459,N_246,In_2769);
xor U1460 (N_1460,In_426,In_4971);
nor U1461 (N_1461,In_4801,In_212);
nand U1462 (N_1462,N_674,N_242);
nor U1463 (N_1463,In_3014,In_1373);
xnor U1464 (N_1464,N_548,In_176);
nand U1465 (N_1465,N_171,In_2818);
nand U1466 (N_1466,In_1768,In_2848);
xnor U1467 (N_1467,In_240,In_1359);
nand U1468 (N_1468,In_3043,In_3139);
xnor U1469 (N_1469,In_1605,In_2237);
xnor U1470 (N_1470,N_841,N_166);
nand U1471 (N_1471,In_4032,In_4850);
and U1472 (N_1472,N_871,In_4303);
xnor U1473 (N_1473,In_282,In_1604);
or U1474 (N_1474,N_823,In_4684);
xor U1475 (N_1475,In_1252,In_4654);
nand U1476 (N_1476,In_312,In_4713);
nor U1477 (N_1477,In_987,In_2651);
xnor U1478 (N_1478,N_281,In_149);
nand U1479 (N_1479,In_19,N_9);
nor U1480 (N_1480,In_3827,N_14);
nor U1481 (N_1481,In_119,In_879);
and U1482 (N_1482,N_230,In_3113);
nand U1483 (N_1483,In_4785,In_1829);
or U1484 (N_1484,In_3102,In_522);
or U1485 (N_1485,In_1294,In_477);
and U1486 (N_1486,N_716,In_539);
and U1487 (N_1487,In_2456,In_4091);
xnor U1488 (N_1488,In_4433,In_2285);
xnor U1489 (N_1489,In_2733,In_1192);
and U1490 (N_1490,In_3707,In_4217);
xor U1491 (N_1491,In_2492,In_2438);
and U1492 (N_1492,In_1261,In_162);
xnor U1493 (N_1493,In_3257,In_2203);
and U1494 (N_1494,In_1135,In_4943);
nor U1495 (N_1495,N_552,In_2200);
or U1496 (N_1496,In_1776,N_142);
and U1497 (N_1497,In_3379,In_1118);
and U1498 (N_1498,In_3115,N_613);
xnor U1499 (N_1499,N_227,In_3871);
and U1500 (N_1500,In_1087,In_2137);
xor U1501 (N_1501,In_2824,In_4922);
nand U1502 (N_1502,In_3112,In_2599);
and U1503 (N_1503,N_150,In_3635);
or U1504 (N_1504,N_579,N_72);
or U1505 (N_1505,In_2531,N_429);
or U1506 (N_1506,In_1247,In_1329);
nor U1507 (N_1507,In_3971,N_77);
nor U1508 (N_1508,In_2970,In_425);
or U1509 (N_1509,In_2484,In_3758);
and U1510 (N_1510,In_2328,N_473);
or U1511 (N_1511,In_3434,N_600);
xor U1512 (N_1512,N_393,In_3037);
nand U1513 (N_1513,In_4318,In_2794);
and U1514 (N_1514,In_2098,In_4834);
nor U1515 (N_1515,In_1728,In_3448);
xor U1516 (N_1516,N_766,In_848);
nor U1517 (N_1517,In_493,In_2815);
nor U1518 (N_1518,In_3969,In_2519);
or U1519 (N_1519,In_2968,N_181);
or U1520 (N_1520,In_1937,In_1035);
nand U1521 (N_1521,N_442,In_3695);
nand U1522 (N_1522,N_770,In_168);
and U1523 (N_1523,In_1141,In_447);
xor U1524 (N_1524,In_2701,N_953);
nor U1525 (N_1525,In_4582,In_2001);
or U1526 (N_1526,N_482,In_3220);
nand U1527 (N_1527,In_1849,N_22);
nor U1528 (N_1528,In_3047,In_2909);
xnor U1529 (N_1529,In_812,In_1843);
or U1530 (N_1530,N_698,In_3762);
or U1531 (N_1531,In_2353,In_4586);
or U1532 (N_1532,In_2867,N_372);
nand U1533 (N_1533,In_3004,N_12);
nand U1534 (N_1534,N_103,In_1433);
nand U1535 (N_1535,N_990,In_3394);
or U1536 (N_1536,N_110,In_509);
xnor U1537 (N_1537,In_3256,In_680);
xor U1538 (N_1538,In_4152,In_4841);
and U1539 (N_1539,In_523,In_3400);
nand U1540 (N_1540,In_3976,N_451);
or U1541 (N_1541,N_237,In_3151);
or U1542 (N_1542,In_167,In_1781);
xnor U1543 (N_1543,In_2033,In_4950);
xor U1544 (N_1544,In_559,In_3666);
nand U1545 (N_1545,N_902,In_300);
xnor U1546 (N_1546,In_2536,In_1396);
nor U1547 (N_1547,In_3675,In_315);
or U1548 (N_1548,In_3108,N_443);
nor U1549 (N_1549,N_193,In_3472);
and U1550 (N_1550,In_3165,In_2746);
and U1551 (N_1551,In_17,N_188);
xnor U1552 (N_1552,In_2217,N_968);
xnor U1553 (N_1553,N_314,In_1076);
xor U1554 (N_1554,In_3775,N_632);
nand U1555 (N_1555,In_520,In_3462);
xor U1556 (N_1556,In_754,N_71);
or U1557 (N_1557,In_3661,N_102);
and U1558 (N_1558,N_525,In_1598);
and U1559 (N_1559,In_2596,In_4870);
nor U1560 (N_1560,In_3829,N_524);
nand U1561 (N_1561,N_799,In_4113);
nor U1562 (N_1562,N_511,In_2816);
and U1563 (N_1563,In_1528,N_891);
nand U1564 (N_1564,In_2616,In_4141);
nor U1565 (N_1565,In_4329,N_498);
or U1566 (N_1566,In_4120,In_4166);
nand U1567 (N_1567,In_876,N_361);
and U1568 (N_1568,In_2184,In_201);
and U1569 (N_1569,In_4845,N_556);
xor U1570 (N_1570,In_4541,In_1367);
and U1571 (N_1571,N_768,In_945);
and U1572 (N_1572,In_4591,N_549);
nand U1573 (N_1573,In_3336,In_1442);
and U1574 (N_1574,In_1609,In_2459);
xor U1575 (N_1575,In_423,In_2104);
xor U1576 (N_1576,In_4286,N_858);
and U1577 (N_1577,In_4635,In_506);
or U1578 (N_1578,In_4452,In_2770);
nor U1579 (N_1579,In_4603,In_2286);
nor U1580 (N_1580,In_1068,In_1269);
and U1581 (N_1581,In_588,N_729);
and U1582 (N_1582,In_4568,In_1927);
nor U1583 (N_1583,In_956,In_1043);
nor U1584 (N_1584,N_925,In_3254);
xnor U1585 (N_1585,In_834,In_1699);
nand U1586 (N_1586,In_4909,In_2691);
and U1587 (N_1587,N_207,In_3475);
or U1588 (N_1588,N_622,N_839);
and U1589 (N_1589,In_399,In_651);
nand U1590 (N_1590,In_3721,N_484);
or U1591 (N_1591,In_4704,In_1061);
and U1592 (N_1592,In_1772,N_988);
xnor U1593 (N_1593,N_859,N_109);
and U1594 (N_1594,In_3589,In_2530);
or U1595 (N_1595,In_4669,In_1797);
and U1596 (N_1596,N_371,In_3540);
and U1597 (N_1597,In_4123,In_102);
xnor U1598 (N_1598,N_806,In_2175);
nor U1599 (N_1599,In_4203,In_3239);
and U1600 (N_1600,In_525,In_1642);
nand U1601 (N_1601,N_477,N_986);
and U1602 (N_1602,In_2325,In_2171);
nand U1603 (N_1603,In_1860,In_4287);
nand U1604 (N_1604,In_4314,In_4790);
nor U1605 (N_1605,In_3884,In_2777);
nor U1606 (N_1606,In_560,In_3973);
and U1607 (N_1607,In_1022,In_1920);
or U1608 (N_1608,In_3122,In_3980);
nand U1609 (N_1609,In_4606,N_738);
nor U1610 (N_1610,In_2540,In_135);
or U1611 (N_1611,N_195,In_843);
or U1612 (N_1612,In_3630,In_1182);
and U1613 (N_1613,N_394,In_1617);
nor U1614 (N_1614,In_869,In_1996);
and U1615 (N_1615,N_408,In_2311);
and U1616 (N_1616,In_192,In_2681);
or U1617 (N_1617,In_2799,In_3103);
and U1618 (N_1618,In_3169,In_3310);
or U1619 (N_1619,In_2403,In_4872);
or U1620 (N_1620,In_4549,In_1282);
nand U1621 (N_1621,In_3097,In_3390);
or U1622 (N_1622,In_3897,N_55);
nor U1623 (N_1623,In_1741,In_1564);
nand U1624 (N_1624,N_331,In_3373);
nand U1625 (N_1625,In_3049,In_4714);
xor U1626 (N_1626,In_805,In_3769);
or U1627 (N_1627,In_2700,N_410);
nand U1628 (N_1628,N_354,In_744);
and U1629 (N_1629,In_3188,In_3077);
and U1630 (N_1630,In_1109,In_2162);
and U1631 (N_1631,In_4765,In_2841);
and U1632 (N_1632,N_638,In_937);
and U1633 (N_1633,In_229,In_4375);
xor U1634 (N_1634,N_922,N_697);
and U1635 (N_1635,In_3772,In_1677);
and U1636 (N_1636,In_2966,In_290);
and U1637 (N_1637,In_4670,N_356);
xnor U1638 (N_1638,N_824,In_4920);
xnor U1639 (N_1639,N_352,In_2501);
and U1640 (N_1640,In_2677,In_3403);
and U1641 (N_1641,In_1839,In_3844);
and U1642 (N_1642,In_339,In_3132);
nand U1643 (N_1643,In_2379,N_260);
nor U1644 (N_1644,In_2251,N_617);
nor U1645 (N_1645,In_1140,In_2041);
xnor U1646 (N_1646,N_179,In_2659);
and U1647 (N_1647,N_605,N_379);
nand U1648 (N_1648,N_401,In_3135);
nand U1649 (N_1649,N_542,In_4911);
and U1650 (N_1650,N_413,In_1084);
nand U1651 (N_1651,In_1313,N_763);
xnor U1652 (N_1652,N_350,In_2444);
nand U1653 (N_1653,In_4706,N_910);
xor U1654 (N_1654,In_55,In_2711);
nor U1655 (N_1655,In_4382,In_2636);
or U1656 (N_1656,In_2240,N_904);
or U1657 (N_1657,In_2744,In_931);
and U1658 (N_1658,In_105,In_440);
xnor U1659 (N_1659,In_131,N_15);
and U1660 (N_1660,In_1320,In_3745);
nand U1661 (N_1661,N_501,N_434);
xnor U1662 (N_1662,In_4453,In_4679);
nand U1663 (N_1663,N_469,N_620);
xor U1664 (N_1664,In_1416,N_973);
nand U1665 (N_1665,In_2339,In_3182);
nor U1666 (N_1666,N_745,In_750);
nor U1667 (N_1667,N_97,In_4288);
xor U1668 (N_1668,In_4585,In_4525);
and U1669 (N_1669,In_997,In_2756);
and U1670 (N_1670,In_165,In_205);
nor U1671 (N_1671,In_3146,In_1339);
nor U1672 (N_1672,N_800,N_43);
and U1673 (N_1673,N_319,In_2099);
or U1674 (N_1674,N_543,In_1954);
or U1675 (N_1675,In_3660,In_2895);
nor U1676 (N_1676,In_821,In_4327);
and U1677 (N_1677,In_1565,In_3148);
xor U1678 (N_1678,N_838,In_1198);
xnor U1679 (N_1679,In_460,In_3223);
or U1680 (N_1680,In_4307,N_681);
or U1681 (N_1681,In_1596,N_172);
nor U1682 (N_1682,In_714,In_2495);
nand U1683 (N_1683,N_773,N_120);
nand U1684 (N_1684,In_224,N_288);
and U1685 (N_1685,In_3262,N_323);
nor U1686 (N_1686,In_3509,In_1963);
xnor U1687 (N_1687,In_4102,In_106);
or U1688 (N_1688,In_555,N_983);
xnor U1689 (N_1689,In_4929,In_3679);
and U1690 (N_1690,In_2066,In_4397);
and U1691 (N_1691,In_1050,N_822);
or U1692 (N_1692,In_2898,N_981);
xnor U1693 (N_1693,In_3196,In_3086);
and U1694 (N_1694,In_4601,In_1090);
nand U1695 (N_1695,N_941,In_3898);
nand U1696 (N_1696,In_1051,In_2437);
nor U1697 (N_1697,In_36,In_4824);
or U1698 (N_1698,N_444,In_1299);
or U1699 (N_1699,In_4520,N_956);
nor U1700 (N_1700,N_837,In_1712);
nand U1701 (N_1701,In_4649,In_2157);
and U1702 (N_1702,N_705,In_4355);
xnor U1703 (N_1703,In_2375,In_3237);
xnor U1704 (N_1704,In_3311,N_412);
and U1705 (N_1705,N_274,In_4865);
and U1706 (N_1706,N_682,In_177);
nor U1707 (N_1707,N_627,In_256);
nand U1708 (N_1708,In_1029,In_2026);
nor U1709 (N_1709,In_3860,In_1582);
or U1710 (N_1710,In_90,In_1988);
and U1711 (N_1711,In_864,In_221);
and U1712 (N_1712,In_1316,In_3502);
or U1713 (N_1713,In_2333,In_2852);
nor U1714 (N_1714,In_842,In_2760);
and U1715 (N_1715,In_40,In_1189);
xnor U1716 (N_1716,In_2680,N_696);
xnor U1717 (N_1717,N_83,In_3961);
nand U1718 (N_1718,In_1975,In_4856);
nor U1719 (N_1719,In_4395,In_1679);
and U1720 (N_1720,In_3873,N_490);
or U1721 (N_1721,In_642,In_4813);
nand U1722 (N_1722,N_530,In_1224);
nor U1723 (N_1723,In_2436,In_2094);
nor U1724 (N_1724,In_2305,In_888);
and U1725 (N_1725,In_431,In_2235);
nor U1726 (N_1726,In_3011,In_489);
xor U1727 (N_1727,N_395,N_744);
and U1728 (N_1728,In_1062,In_174);
nor U1729 (N_1729,In_2084,In_1649);
nor U1730 (N_1730,N_286,In_1401);
or U1731 (N_1731,In_285,In_3411);
nand U1732 (N_1732,In_413,In_2967);
xnor U1733 (N_1733,N_47,In_385);
and U1734 (N_1734,In_366,In_845);
xnor U1735 (N_1735,N_915,In_56);
or U1736 (N_1736,N_790,N_654);
xor U1737 (N_1737,In_3386,In_1760);
or U1738 (N_1738,In_2696,In_4284);
nor U1739 (N_1739,In_3277,In_2823);
nand U1740 (N_1740,In_2643,In_198);
nand U1741 (N_1741,In_1475,In_21);
and U1742 (N_1742,In_2937,In_3622);
nor U1743 (N_1743,In_2261,In_346);
nor U1744 (N_1744,N_651,N_671);
nand U1745 (N_1745,In_3594,In_3600);
and U1746 (N_1746,In_2380,N_435);
or U1747 (N_1747,In_3538,In_4010);
xor U1748 (N_1748,In_314,N_869);
and U1749 (N_1749,In_2775,In_83);
or U1750 (N_1750,In_618,In_1632);
or U1751 (N_1751,In_4036,In_3481);
nand U1752 (N_1752,In_2447,In_1567);
xnor U1753 (N_1753,N_185,In_1156);
nor U1754 (N_1754,In_2821,In_3941);
nand U1755 (N_1755,In_1542,In_689);
xnor U1756 (N_1756,In_291,In_1698);
xnor U1757 (N_1757,N_258,N_512);
nor U1758 (N_1758,N_753,N_755);
or U1759 (N_1759,N_119,In_958);
xor U1760 (N_1760,In_122,N_794);
or U1761 (N_1761,In_726,In_4185);
or U1762 (N_1762,In_3820,In_146);
xor U1763 (N_1763,In_2801,In_4349);
nand U1764 (N_1764,N_802,In_2136);
nand U1765 (N_1765,In_946,In_4537);
or U1766 (N_1766,In_110,In_194);
and U1767 (N_1767,In_2795,In_4513);
nor U1768 (N_1768,In_4072,In_2246);
or U1769 (N_1769,In_4331,In_2365);
or U1770 (N_1770,In_878,In_1175);
or U1771 (N_1771,In_1663,In_633);
nor U1772 (N_1772,N_414,N_201);
nand U1773 (N_1773,In_2400,In_4231);
or U1774 (N_1774,N_582,In_1150);
nand U1775 (N_1775,In_3079,In_1793);
nand U1776 (N_1776,N_13,In_1902);
nor U1777 (N_1777,In_2552,In_3361);
and U1778 (N_1778,In_1016,In_450);
and U1779 (N_1779,In_3,In_2745);
nor U1780 (N_1780,In_3865,In_3671);
nor U1781 (N_1781,In_2972,In_2196);
nor U1782 (N_1782,In_1110,N_268);
and U1783 (N_1783,In_855,In_4018);
or U1784 (N_1784,In_2148,N_573);
or U1785 (N_1785,In_1073,In_3641);
nand U1786 (N_1786,In_2336,In_1216);
xnor U1787 (N_1787,In_767,N_929);
and U1788 (N_1788,In_264,In_2788);
xor U1789 (N_1789,In_4432,In_2996);
and U1790 (N_1790,In_4798,N_987);
xnor U1791 (N_1791,In_2028,In_241);
nand U1792 (N_1792,N_793,In_2342);
nor U1793 (N_1793,In_3685,In_1390);
xor U1794 (N_1794,In_2410,In_1645);
nand U1795 (N_1795,In_1729,N_133);
or U1796 (N_1796,N_767,In_862);
and U1797 (N_1797,N_454,In_2019);
nand U1798 (N_1798,In_220,In_4878);
nor U1799 (N_1799,In_3719,In_2514);
and U1800 (N_1800,N_257,In_1872);
or U1801 (N_1801,In_942,In_247);
xnor U1802 (N_1802,In_2198,In_4370);
xnor U1803 (N_1803,In_2588,In_1065);
nand U1804 (N_1804,N_899,In_124);
nor U1805 (N_1805,N_658,N_35);
nor U1806 (N_1806,In_2933,In_1846);
and U1807 (N_1807,In_2758,In_2693);
and U1808 (N_1808,N_322,N_508);
and U1809 (N_1809,In_1257,In_3024);
nand U1810 (N_1810,In_692,In_2349);
nor U1811 (N_1811,In_1227,N_798);
nor U1812 (N_1812,In_1539,N_528);
and U1813 (N_1813,In_4160,In_1816);
xnor U1814 (N_1814,In_2603,In_4167);
and U1815 (N_1815,N_407,In_3023);
or U1816 (N_1816,N_636,In_1923);
nand U1817 (N_1817,In_2168,In_2768);
xnor U1818 (N_1818,N_758,In_1904);
xor U1819 (N_1819,In_3274,In_504);
or U1820 (N_1820,N_686,N_854);
and U1821 (N_1821,In_3922,N_303);
nand U1822 (N_1822,In_1738,In_3415);
or U1823 (N_1823,In_134,N_526);
or U1824 (N_1824,In_4368,In_2675);
xor U1825 (N_1825,N_139,In_4069);
nor U1826 (N_1826,In_3807,In_3317);
nor U1827 (N_1827,In_148,In_2152);
and U1828 (N_1828,In_2665,N_116);
nor U1829 (N_1829,In_3824,N_298);
nand U1830 (N_1830,In_1815,In_3951);
nor U1831 (N_1831,In_2944,In_1246);
xnor U1832 (N_1832,In_2009,In_667);
xor U1833 (N_1833,In_2093,In_4154);
nor U1834 (N_1834,N_642,In_279);
nand U1835 (N_1835,In_2280,In_3553);
nor U1836 (N_1836,In_280,In_2689);
nand U1837 (N_1837,N_439,In_1865);
and U1838 (N_1838,In_967,N_895);
and U1839 (N_1839,N_325,In_3121);
nand U1840 (N_1840,In_1640,In_3410);
or U1841 (N_1841,N_588,In_4710);
nor U1842 (N_1842,In_1994,N_365);
xnor U1843 (N_1843,In_3248,N_495);
nand U1844 (N_1844,In_3131,N_20);
xnor U1845 (N_1845,In_2710,In_4222);
xor U1846 (N_1846,In_3904,In_1508);
xnor U1847 (N_1847,In_2024,In_4352);
nand U1848 (N_1848,In_4087,N_680);
or U1849 (N_1849,In_2584,N_330);
nor U1850 (N_1850,In_164,In_1637);
and U1851 (N_1851,In_716,In_490);
and U1852 (N_1852,In_3072,In_988);
nand U1853 (N_1853,In_3958,In_3910);
and U1854 (N_1854,In_4206,In_2723);
and U1855 (N_1855,N_468,In_2647);
nor U1856 (N_1856,In_4924,In_96);
and U1857 (N_1857,In_2161,In_1982);
and U1858 (N_1858,In_3960,N_69);
nor U1859 (N_1859,N_874,In_541);
or U1860 (N_1860,In_2835,In_3463);
or U1861 (N_1861,N_875,In_4894);
xor U1862 (N_1862,In_1009,N_934);
nor U1863 (N_1863,N_863,In_4367);
xor U1864 (N_1864,In_4401,In_2641);
nand U1865 (N_1865,In_660,In_2555);
nand U1866 (N_1866,In_2216,In_790);
or U1867 (N_1867,N_192,In_3817);
xor U1868 (N_1868,N_346,In_4233);
or U1869 (N_1869,In_2468,In_1800);
or U1870 (N_1870,In_2523,N_513);
and U1871 (N_1871,N_376,In_1886);
nand U1872 (N_1872,In_708,N_433);
or U1873 (N_1873,N_882,In_4221);
nand U1874 (N_1874,In_3996,In_3703);
nor U1875 (N_1875,In_548,In_4934);
xor U1876 (N_1876,In_4980,N_944);
nand U1877 (N_1877,N_453,In_4677);
xor U1878 (N_1878,In_4981,In_2211);
nor U1879 (N_1879,In_3753,In_360);
nor U1880 (N_1880,N_639,In_952);
xor U1881 (N_1881,In_2670,In_4112);
and U1882 (N_1882,In_1687,N_167);
or U1883 (N_1883,In_410,N_221);
or U1884 (N_1884,In_502,In_724);
nor U1885 (N_1885,In_1710,In_3554);
xnor U1886 (N_1886,In_1736,In_2362);
and U1887 (N_1887,In_2407,In_4270);
xnor U1888 (N_1888,In_1172,In_1745);
xor U1889 (N_1889,In_118,In_2903);
and U1890 (N_1890,In_1734,In_3249);
or U1891 (N_1891,In_4356,N_518);
and U1892 (N_1892,In_4793,N_21);
nor U1893 (N_1893,N_98,N_791);
xnor U1894 (N_1894,In_2164,In_1662);
nor U1895 (N_1895,In_2812,N_615);
or U1896 (N_1896,In_4663,In_4379);
xnor U1897 (N_1897,In_3147,In_3891);
nand U1898 (N_1898,In_4266,In_4647);
xor U1899 (N_1899,N_91,In_3268);
nor U1900 (N_1900,In_2762,N_191);
nand U1901 (N_1901,N_363,In_4726);
and U1902 (N_1902,N_386,In_1774);
and U1903 (N_1903,In_4688,In_1251);
or U1904 (N_1904,In_3054,N_321);
and U1905 (N_1905,N_772,In_1517);
or U1906 (N_1906,In_2167,In_4272);
and U1907 (N_1907,In_2798,In_2055);
or U1908 (N_1908,In_2092,N_402);
xnor U1909 (N_1909,In_4046,N_860);
nand U1910 (N_1910,N_580,In_2269);
nand U1911 (N_1911,In_1491,In_3912);
or U1912 (N_1912,In_1681,In_978);
xnor U1913 (N_1913,In_1304,N_339);
xnor U1914 (N_1914,In_2273,In_2343);
or U1915 (N_1915,In_3451,In_2398);
nand U1916 (N_1916,N_566,N_514);
xor U1917 (N_1917,In_2357,In_3467);
or U1918 (N_1918,In_1448,N_74);
and U1919 (N_1919,N_522,In_646);
or U1920 (N_1920,In_4966,In_2847);
nand U1921 (N_1921,In_2086,In_975);
nor U1922 (N_1922,In_4343,In_1690);
nand U1923 (N_1923,In_604,N_108);
or U1924 (N_1924,In_1332,N_533);
and U1925 (N_1925,In_3694,N_128);
nand U1926 (N_1926,N_868,N_897);
xnor U1927 (N_1927,In_865,In_1139);
and U1928 (N_1928,In_1355,In_1765);
and U1929 (N_1929,In_1896,In_4897);
xor U1930 (N_1930,In_3788,In_785);
xnor U1931 (N_1931,N_994,In_208);
and U1932 (N_1932,In_964,In_1722);
nor U1933 (N_1933,N_912,N_449);
or U1934 (N_1934,N_722,In_61);
or U1935 (N_1935,N_909,N_725);
or U1936 (N_1936,N_403,In_873);
and U1937 (N_1937,In_3505,In_3528);
xnor U1938 (N_1938,In_3099,N_931);
nor U1939 (N_1939,In_2829,In_2118);
or U1940 (N_1940,In_1826,In_84);
or U1941 (N_1941,In_2874,In_4456);
and U1942 (N_1942,In_4128,In_3607);
xnor U1943 (N_1943,In_3488,In_2927);
nand U1944 (N_1944,In_777,In_1014);
and U1945 (N_1945,N_567,In_3868);
nor U1946 (N_1946,In_142,In_1242);
and U1947 (N_1947,In_4724,In_2244);
xor U1948 (N_1948,In_2838,N_180);
xnor U1949 (N_1949,In_1784,In_4381);
nand U1950 (N_1950,In_66,In_4330);
and U1951 (N_1951,In_1033,N_381);
and U1952 (N_1952,In_936,N_79);
nor U1953 (N_1953,N_664,In_2830);
nor U1954 (N_1954,N_448,N_377);
nand U1955 (N_1955,In_3163,In_3746);
xnor U1956 (N_1956,In_4853,In_1034);
or U1957 (N_1957,In_1763,N_147);
nor U1958 (N_1958,In_3328,In_2038);
xor U1959 (N_1959,In_3238,In_854);
or U1960 (N_1960,In_2803,In_197);
xor U1961 (N_1961,N_426,N_125);
nor U1962 (N_1962,N_903,In_3947);
nand U1963 (N_1963,In_3937,N_670);
nor U1964 (N_1964,In_2506,In_1791);
and U1965 (N_1965,In_832,In_4341);
and U1966 (N_1966,N_259,N_111);
nand U1967 (N_1967,In_1258,N_997);
or U1968 (N_1968,In_2885,In_1692);
or U1969 (N_1969,In_2509,In_910);
nand U1970 (N_1970,In_3381,N_240);
or U1971 (N_1971,In_501,In_3780);
and U1972 (N_1972,In_418,N_876);
and U1973 (N_1973,In_4498,In_4951);
xnor U1974 (N_1974,In_766,In_4376);
and U1975 (N_1975,In_2875,In_2315);
nor U1976 (N_1976,In_4282,In_3413);
xor U1977 (N_1977,In_853,In_2433);
nor U1978 (N_1978,In_13,In_650);
nand U1979 (N_1979,N_255,In_4084);
and U1980 (N_1980,N_782,In_1374);
nor U1981 (N_1981,N_164,In_4861);
xnor U1982 (N_1982,In_571,In_3006);
or U1983 (N_1983,In_3406,In_4458);
or U1984 (N_1984,In_1412,In_48);
nand U1985 (N_1985,In_3366,In_412);
or U1986 (N_1986,In_4555,In_3929);
nand U1987 (N_1987,N_411,In_350);
or U1988 (N_1988,In_3967,N_749);
nand U1989 (N_1989,N_485,In_3785);
nand U1990 (N_1990,In_4190,In_436);
nand U1991 (N_1991,In_1576,In_4326);
or U1992 (N_1992,In_2215,In_3757);
or U1993 (N_1993,In_485,In_4700);
nand U1994 (N_1994,In_3431,In_4696);
and U1995 (N_1995,In_2793,In_1410);
xor U1996 (N_1996,N_479,In_3346);
and U1997 (N_1997,In_2882,N_450);
nand U1998 (N_1998,In_3572,In_1275);
nor U1999 (N_1999,In_3954,In_819);
xor U2000 (N_2000,In_3282,In_2091);
nand U2001 (N_2001,In_4848,N_1252);
nand U2002 (N_2002,N_1422,In_3412);
nand U2003 (N_2003,N_1086,In_2106);
xnor U2004 (N_2004,N_821,N_701);
and U2005 (N_2005,N_84,N_1504);
or U2006 (N_2006,In_75,In_3767);
or U2007 (N_2007,N_1283,N_540);
xor U2008 (N_2008,N_1312,In_3159);
nor U2009 (N_2009,In_722,N_1717);
xor U2010 (N_2010,In_1771,In_1854);
and U2011 (N_2011,N_534,N_1154);
nor U2012 (N_2012,N_825,In_2483);
or U2013 (N_2013,N_1964,In_2402);
or U2014 (N_2014,In_4879,N_1265);
and U2015 (N_2015,N_1448,N_135);
nor U2016 (N_2016,N_1505,N_554);
nand U2017 (N_2017,In_4958,N_1495);
nor U2018 (N_2018,In_3517,N_1880);
nand U2019 (N_2019,In_3699,N_348);
nor U2020 (N_2020,In_4728,In_324);
nor U2021 (N_2021,In_2858,In_3335);
nand U2022 (N_2022,N_1889,In_1318);
or U2023 (N_2023,N_1409,In_4092);
nor U2024 (N_2024,N_252,N_1529);
xor U2025 (N_2025,N_1179,N_187);
xnor U2026 (N_2026,In_1925,N_247);
or U2027 (N_2027,In_4396,N_152);
and U2028 (N_2028,N_272,In_550);
and U2029 (N_2029,N_1815,In_46);
nand U2030 (N_2030,N_1580,N_1721);
and U2031 (N_2031,N_1562,In_4450);
nand U2032 (N_2032,N_1888,N_33);
nand U2033 (N_2033,N_703,In_2367);
nand U2034 (N_2034,In_4613,N_1614);
nand U2035 (N_2035,In_4320,In_3450);
or U2036 (N_2036,N_129,In_1083);
xnor U2037 (N_2037,N_1483,In_4666);
nor U2038 (N_2038,N_1359,N_1539);
xor U2039 (N_2039,In_1125,In_1627);
and U2040 (N_2040,In_4789,N_1156);
nand U2041 (N_2041,In_2931,N_1989);
nand U2042 (N_2042,N_368,N_1057);
or U2043 (N_2043,N_1548,In_512);
nand U2044 (N_2044,In_1435,In_132);
xnor U2045 (N_2045,In_1898,N_1783);
or U2046 (N_2046,In_3880,In_4589);
nand U2047 (N_2047,In_1634,In_4121);
nand U2048 (N_2048,In_1377,In_3877);
or U2049 (N_2049,N_1433,In_1271);
and U2050 (N_2050,In_4562,N_1510);
nand U2051 (N_2051,In_3811,In_1818);
nor U2052 (N_2052,N_1387,N_1511);
nor U2053 (N_2053,N_467,In_1425);
or U2054 (N_2054,In_2873,N_1402);
and U2055 (N_2055,In_1977,In_1042);
xnor U2056 (N_2056,N_1257,N_1371);
xor U2057 (N_2057,In_1597,N_1241);
nand U2058 (N_2058,In_904,In_3378);
xor U2059 (N_2059,In_1890,N_936);
or U2060 (N_2060,In_2949,In_4556);
and U2061 (N_2061,N_1078,N_224);
or U2062 (N_2062,In_979,N_1111);
nor U2063 (N_2063,N_355,N_1464);
and U2064 (N_2064,In_1324,N_1667);
and U2065 (N_2065,In_3556,In_3823);
xor U2066 (N_2066,N_1437,N_1406);
and U2067 (N_2067,N_715,In_3761);
nand U2068 (N_2068,N_1027,N_1706);
nand U2069 (N_2069,N_1776,N_317);
and U2070 (N_2070,In_4182,N_1000);
nor U2071 (N_2071,In_4200,In_358);
nor U2072 (N_2072,In_3293,In_2259);
or U2073 (N_2073,N_1943,N_678);
nand U2074 (N_2074,N_333,In_3546);
nand U2075 (N_2075,In_4748,In_4774);
or U2076 (N_2076,N_427,N_1249);
xnor U2077 (N_2077,In_4020,N_1701);
or U2078 (N_2078,In_4055,N_1442);
or U2079 (N_2079,N_1879,In_1468);
or U2080 (N_2080,In_2811,N_1986);
nor U2081 (N_2081,N_1054,N_437);
nor U2082 (N_2082,N_1863,N_1236);
nor U2083 (N_2083,In_121,N_980);
xor U2084 (N_2084,N_1954,In_3852);
nor U2085 (N_2085,N_422,In_2558);
or U2086 (N_2086,N_1907,In_2785);
nand U2087 (N_2087,In_2439,In_4835);
xnor U2088 (N_2088,In_3034,In_4099);
nand U2089 (N_2089,N_1635,In_809);
nor U2090 (N_2090,N_1196,In_3934);
nor U2091 (N_2091,N_1881,In_4311);
nand U2092 (N_2092,In_4271,In_3743);
and U2093 (N_2093,N_1244,N_36);
nand U2094 (N_2094,In_1529,In_2686);
or U2095 (N_2095,N_337,In_2752);
or U2096 (N_2096,In_394,In_887);
xnor U2097 (N_2097,In_181,In_891);
nor U2098 (N_2098,In_1120,In_3524);
xnor U2099 (N_2099,In_246,N_1146);
nor U2100 (N_2100,N_40,In_922);
and U2101 (N_2101,In_893,N_1756);
xnor U2102 (N_2102,N_1396,In_3902);
xor U2103 (N_2103,In_1599,N_818);
or U2104 (N_2104,N_1360,N_575);
nor U2105 (N_2105,N_1499,In_1884);
nor U2106 (N_2106,N_707,N_1810);
nand U2107 (N_2107,N_1586,In_4544);
and U2108 (N_2108,In_1047,N_594);
and U2109 (N_2109,In_99,In_4132);
nor U2110 (N_2110,N_1291,N_1090);
xor U2111 (N_2111,In_2952,N_1043);
xor U2112 (N_2112,N_764,In_2025);
nor U2113 (N_2113,In_1064,In_1449);
nand U2114 (N_2114,N_1475,In_2642);
xnor U2115 (N_2115,N_648,In_1163);
or U2116 (N_2116,N_630,In_2151);
nand U2117 (N_2117,In_4071,N_1737);
nor U2118 (N_2118,N_34,In_4868);
nor U2119 (N_2119,N_1945,N_198);
nand U2120 (N_2120,N_1215,In_1641);
and U2121 (N_2121,N_1622,In_1174);
nor U2122 (N_2122,In_204,N_500);
or U2123 (N_2123,In_2448,N_1024);
and U2124 (N_2124,N_75,In_4836);
nand U2125 (N_2125,In_3401,N_1573);
xnor U2126 (N_2126,N_1260,N_446);
and U2127 (N_2127,N_1276,N_85);
nor U2128 (N_2128,N_1138,In_1496);
nor U2129 (N_2129,N_1797,N_249);
nor U2130 (N_2130,In_4716,N_1715);
nor U2131 (N_2131,In_2197,In_4479);
and U2132 (N_2132,N_1020,In_2389);
nand U2133 (N_2133,N_1178,In_4604);
and U2134 (N_2134,N_1055,N_236);
and U2135 (N_2135,In_3236,N_349);
xor U2136 (N_2136,In_2887,In_1351);
and U2137 (N_2137,N_1824,N_1093);
xnor U2138 (N_2138,N_1627,N_1826);
nor U2139 (N_2139,In_2820,In_3710);
nand U2140 (N_2140,N_1710,N_1662);
and U2141 (N_2141,In_3997,N_911);
xor U2142 (N_2142,N_1632,In_2027);
nor U2143 (N_2143,In_4917,In_2730);
xor U2144 (N_2144,N_1125,In_1361);
nor U2145 (N_2145,N_1526,In_2480);
nor U2146 (N_2146,N_489,In_803);
or U2147 (N_2147,In_2427,In_1859);
nor U2148 (N_2148,In_1945,In_4312);
nand U2149 (N_2149,N_1143,In_3283);
and U2150 (N_2150,In_1205,N_388);
or U2151 (N_2151,In_3439,N_1861);
or U2152 (N_2152,N_1332,N_1224);
or U2153 (N_2153,N_1267,N_1533);
and U2154 (N_2154,N_1344,N_1554);
nor U2155 (N_2155,In_1203,In_2854);
or U2156 (N_2156,In_1900,In_867);
nand U2157 (N_2157,In_4100,In_2658);
and U2158 (N_2158,In_130,In_1244);
nor U2159 (N_2159,In_4948,N_1399);
nor U2160 (N_2160,In_4406,In_1223);
and U2161 (N_2161,N_1150,In_157);
nor U2162 (N_2162,In_1571,In_4162);
or U2163 (N_2163,N_1915,In_4291);
or U2164 (N_2164,N_223,In_2332);
and U2165 (N_2165,N_168,N_576);
or U2166 (N_2166,In_4187,In_260);
and U2167 (N_2167,In_2920,N_332);
and U2168 (N_2168,N_1001,N_1115);
nand U2169 (N_2169,In_901,N_1349);
xnor U2170 (N_2170,In_693,N_478);
nand U2171 (N_2171,In_3709,N_739);
xor U2172 (N_2172,N_1624,N_1765);
nor U2173 (N_2173,N_1234,N_1922);
or U2174 (N_2174,In_4646,In_1159);
or U2175 (N_2175,In_377,In_4232);
nor U2176 (N_2176,N_1050,In_1764);
or U2177 (N_2177,In_4426,N_1992);
xnor U2178 (N_2178,In_3733,N_1255);
xor U2179 (N_2179,N_523,In_4598);
and U2180 (N_2180,N_94,In_2667);
and U2181 (N_2181,In_841,N_908);
or U2182 (N_2182,N_603,In_3095);
and U2183 (N_2183,N_1767,N_19);
nand U2184 (N_2184,N_1525,N_1820);
or U2185 (N_2185,In_4295,N_695);
nor U2186 (N_2186,N_1859,N_1550);
nand U2187 (N_2187,In_657,N_1802);
or U2188 (N_2188,N_900,In_2120);
and U2189 (N_2189,N_1925,N_1900);
xor U2190 (N_2190,N_593,N_1910);
and U2191 (N_2191,N_1488,N_1673);
or U2192 (N_2192,N_406,In_1021);
xnor U2193 (N_2193,N_282,In_2037);
nor U2194 (N_2194,In_1786,N_1430);
nor U2195 (N_2195,In_12,In_2851);
xnor U2196 (N_2196,In_2764,In_1015);
or U2197 (N_2197,N_1872,N_398);
nor U2198 (N_2198,In_3279,N_1970);
nor U2199 (N_2199,N_459,N_27);
nand U2200 (N_2200,N_1254,In_3251);
xor U2201 (N_2201,In_2796,N_289);
nor U2202 (N_2202,N_492,N_784);
xor U2203 (N_2203,N_1741,N_1242);
nor U2204 (N_2204,In_4035,In_3855);
nor U2205 (N_2205,N_1939,N_614);
and U2206 (N_2206,In_2323,N_1308);
nand U2207 (N_2207,In_2870,In_3518);
nand U2208 (N_2208,N_105,N_1984);
xnor U2209 (N_2209,N_304,N_1192);
and U2210 (N_2210,In_1363,In_3825);
or U2211 (N_2211,N_1432,N_1731);
xnor U2212 (N_2212,N_1769,In_3864);
nand U2213 (N_2213,In_4504,N_1290);
nor U2214 (N_2214,N_1512,N_1659);
nor U2215 (N_2215,N_1343,N_159);
nor U2216 (N_2216,In_213,N_1571);
xor U2217 (N_2217,In_3471,N_241);
or U2218 (N_2218,In_930,In_2724);
nor U2219 (N_2219,In_3529,In_478);
and U2220 (N_2220,In_2149,N_1415);
or U2221 (N_2221,In_3637,In_3555);
or U2222 (N_2222,N_796,In_4747);
or U2223 (N_2223,N_625,N_1743);
or U2224 (N_2224,N_535,N_539);
and U2225 (N_2225,In_551,N_850);
and U2226 (N_2226,In_831,In_4017);
nor U2227 (N_2227,In_1398,In_911);
or U2228 (N_2228,N_1560,N_203);
and U2229 (N_2229,In_1007,In_994);
or U2230 (N_2230,In_729,In_673);
and U2231 (N_2231,N_1167,In_4362);
or U2232 (N_2232,N_1137,N_1210);
and U2233 (N_2233,In_439,In_2819);
nor U2234 (N_2234,N_1366,N_1800);
and U2235 (N_2235,N_1012,In_3659);
and U2236 (N_2236,In_2370,In_2277);
or U2237 (N_2237,In_1429,In_3492);
nor U2238 (N_2238,In_2587,N_1948);
or U2239 (N_2239,N_726,In_3845);
nand U2240 (N_2240,In_2003,N_1033);
xor U2241 (N_2241,In_1058,In_287);
nor U2242 (N_2242,N_1240,N_1968);
xnor U2243 (N_2243,N_73,In_3815);
xnor U2244 (N_2244,N_1098,N_720);
or U2245 (N_2245,N_945,N_1849);
and U2246 (N_2246,In_2725,N_1509);
nand U2247 (N_2247,In_4064,N_1830);
nand U2248 (N_2248,N_1613,In_326);
or U2249 (N_2249,In_1031,N_1487);
nand U2250 (N_2250,In_2227,N_1041);
nand U2251 (N_2251,In_607,In_3156);
nand U2252 (N_2252,In_2213,N_735);
nor U2253 (N_2253,N_1320,N_700);
or U2254 (N_2254,In_2076,In_4004);
and U2255 (N_2255,In_4201,N_1246);
or U2256 (N_2256,N_1718,In_3781);
and U2257 (N_2257,N_1957,N_1353);
nand U2258 (N_2258,N_1916,In_2940);
nand U2259 (N_2259,In_2602,N_1132);
nor U2260 (N_2260,In_3621,In_1731);
or U2261 (N_2261,N_1069,In_3669);
nand U2262 (N_2262,In_1718,N_1672);
or U2263 (N_2263,N_553,N_447);
nand U2264 (N_2264,N_1117,In_727);
and U2265 (N_2265,N_1819,N_1577);
nand U2266 (N_2266,N_979,In_1802);
nand U2267 (N_2267,N_893,N_1102);
and U2268 (N_2268,N_1858,N_154);
xor U2269 (N_2269,N_1191,In_2182);
nor U2270 (N_2270,In_4610,In_3225);
xor U2271 (N_2271,In_3808,In_811);
xnor U2272 (N_2272,N_1205,In_1204);
and U2273 (N_2273,In_2212,In_1371);
xor U2274 (N_2274,N_775,In_403);
or U2275 (N_2275,In_3419,In_304);
and U2276 (N_2276,In_1344,In_2877);
and U2277 (N_2277,In_2205,In_2582);
xnor U2278 (N_2278,N_362,N_112);
nor U2279 (N_2279,N_1142,N_163);
nor U2280 (N_2280,In_4752,N_647);
xnor U2281 (N_2281,In_740,In_1481);
and U2282 (N_2282,In_4799,N_1887);
and U2283 (N_2283,In_4497,N_1232);
xnor U2284 (N_2284,In_4043,N_1282);
and U2285 (N_2285,N_1048,In_2321);
nor U2286 (N_2286,N_1517,In_4198);
xnor U2287 (N_2287,N_1336,In_3187);
nor U2288 (N_2288,In_2564,In_245);
and U2289 (N_2289,N_1008,In_3672);
nor U2290 (N_2290,In_1032,N_1019);
xnor U2291 (N_2291,In_2354,In_3126);
nand U2292 (N_2292,N_1202,N_1745);
or U2293 (N_2293,N_1874,N_1325);
or U2294 (N_2294,In_4806,In_2473);
xor U2295 (N_2295,N_265,N_1788);
nand U2296 (N_2296,N_136,N_24);
nor U2297 (N_2297,N_1583,In_2124);
nor U2298 (N_2298,In_4590,In_3184);
nand U2299 (N_2299,N_1380,In_1667);
or U2300 (N_2300,N_1891,N_375);
or U2301 (N_2301,N_1237,N_1658);
xor U2302 (N_2302,N_1626,In_1480);
xnor U2303 (N_2303,In_91,N_1034);
xor U2304 (N_2304,In_3766,N_1022);
nor U2305 (N_2305,In_3603,In_3285);
and U2306 (N_2306,In_1153,N_1816);
nand U2307 (N_2307,In_4110,N_1193);
nor U2308 (N_2308,In_2715,N_608);
nor U2309 (N_2309,In_1739,In_3420);
nand U2310 (N_2310,In_3349,N_1705);
nor U2311 (N_2311,N_1966,In_206);
and U2312 (N_2312,In_3765,In_2326);
nor U2313 (N_2313,In_1056,In_430);
xnor U2314 (N_2314,In_3702,N_1481);
xor U2315 (N_2315,N_1683,In_973);
and U2316 (N_2316,N_684,N_1870);
or U2317 (N_2317,N_1306,In_598);
and U2318 (N_2318,N_92,In_1897);
or U2319 (N_2319,N_1952,In_1782);
or U2320 (N_2320,In_3786,In_4955);
nand U2321 (N_2321,N_173,N_1846);
nor U2322 (N_2322,In_3233,In_2355);
xnor U2323 (N_2323,N_1397,In_1762);
or U2324 (N_2324,N_1963,N_1498);
or U2325 (N_2325,N_1477,N_1644);
and U2326 (N_2326,In_4148,In_4739);
nand U2327 (N_2327,N_1878,N_1960);
xor U2328 (N_2328,N_1173,In_4807);
xnor U2329 (N_2329,N_1670,N_1231);
nand U2330 (N_2330,In_1907,N_310);
nor U2331 (N_2331,N_957,N_1274);
nor U2332 (N_2332,In_4705,In_2063);
or U2333 (N_2333,In_359,N_1829);
and U2334 (N_2334,N_1460,In_2284);
and U2335 (N_2335,In_3799,N_343);
xnor U2336 (N_2336,N_101,In_258);
or U2337 (N_2337,In_2039,N_1998);
or U2338 (N_2338,In_1479,N_400);
xnor U2339 (N_2339,N_1961,In_182);
nand U2340 (N_2340,In_1461,In_79);
nand U2341 (N_2341,N_438,In_2528);
nand U2342 (N_2342,N_683,In_2784);
nand U2343 (N_2343,In_3749,N_846);
and U2344 (N_2344,N_1303,In_4854);
nand U2345 (N_2345,In_2719,In_4415);
xnor U2346 (N_2346,In_453,In_4293);
xor U2347 (N_2347,N_1541,N_66);
or U2348 (N_2348,N_1748,In_4518);
nor U2349 (N_2349,In_4846,In_1218);
and U2350 (N_2350,N_1735,In_3289);
or U2351 (N_2351,In_1280,In_4442);
xor U2352 (N_2352,In_4075,N_359);
and U2353 (N_2353,N_1886,In_731);
xnor U2354 (N_2354,N_1625,In_1012);
nand U2355 (N_2355,In_2656,N_1198);
or U2356 (N_2356,N_1393,In_532);
nand U2357 (N_2357,In_4777,In_712);
nand U2358 (N_2358,In_2626,N_1734);
nor U2359 (N_2359,N_313,N_1785);
or U2360 (N_2360,In_2525,N_1163);
nor U2361 (N_2361,N_334,N_1120);
xnor U2362 (N_2362,In_2566,N_1565);
nor U2363 (N_2363,N_626,N_867);
or U2364 (N_2364,N_1134,N_1982);
or U2365 (N_2365,In_3178,N_843);
or U2366 (N_2366,In_872,N_1987);
nor U2367 (N_2367,N_225,N_415);
or U2368 (N_2368,N_1787,N_1850);
and U2369 (N_2369,N_1194,In_4108);
nor U2370 (N_2370,N_1088,N_1059);
or U2371 (N_2371,N_1133,In_671);
nand U2372 (N_2372,N_1139,N_1074);
or U2373 (N_2373,N_1678,In_3051);
xnor U2374 (N_2374,N_1355,In_4547);
xor U2375 (N_2375,N_699,N_515);
xnor U2376 (N_2376,In_3466,In_435);
and U2377 (N_2377,In_2620,N_1615);
xor U2378 (N_2378,In_3809,N_1831);
nand U2379 (N_2379,In_3920,N_1890);
xor U2380 (N_2380,In_921,In_1980);
or U2381 (N_2381,N_1558,N_1722);
nor U2382 (N_2382,In_562,N_728);
xnor U2383 (N_2383,In_1620,In_1457);
and U2384 (N_2384,N_1148,N_1775);
or U2385 (N_2385,In_1967,N_1927);
nand U2386 (N_2386,N_828,N_792);
xor U2387 (N_2387,In_1608,In_4164);
nand U2388 (N_2388,In_4371,N_1131);
nand U2389 (N_2389,N_1211,In_4680);
nand U2390 (N_2390,In_446,N_50);
xor U2391 (N_2391,In_4899,In_254);
nor U2392 (N_2392,In_4122,N_1697);
nor U2393 (N_2393,N_1347,In_4377);
nand U2394 (N_2394,N_1334,In_6);
or U2395 (N_2395,N_149,N_1919);
and U2396 (N_2396,In_4788,In_2013);
and U2397 (N_2397,In_2218,N_1207);
nand U2398 (N_2398,N_243,N_612);
nor U2399 (N_2399,N_529,In_4564);
nor U2400 (N_2400,In_1578,N_870);
and U2401 (N_2401,In_2,In_3118);
nand U2402 (N_2402,In_217,In_2703);
and U2403 (N_2403,N_1990,N_123);
nor U2404 (N_2404,N_1594,N_1983);
nand U2405 (N_2405,N_1287,In_71);
nor U2406 (N_2406,N_1996,N_1578);
nor U2407 (N_2407,In_1276,N_946);
nand U2408 (N_2408,N_1489,In_2266);
or U2409 (N_2409,In_1360,N_1168);
and U2410 (N_2410,N_851,In_1093);
nor U2411 (N_2411,In_3499,In_4516);
xnor U2412 (N_2412,N_1155,In_3357);
and U2413 (N_2413,In_886,In_190);
xor U2414 (N_2414,N_1243,N_827);
and U2415 (N_2415,N_1354,N_199);
or U2416 (N_2416,In_739,In_4438);
and U2417 (N_2417,N_475,In_2242);
xor U2418 (N_2418,In_3284,N_653);
xor U2419 (N_2419,In_953,In_3389);
xor U2420 (N_2420,In_3252,In_679);
nor U2421 (N_2421,In_629,In_4019);
or U2422 (N_2422,N_329,N_509);
nor U2423 (N_2423,N_1462,In_3454);
nand U2424 (N_2424,N_1993,In_4886);
and U2425 (N_2425,In_1903,In_2666);
and U2426 (N_2426,In_4184,In_3768);
nor U2427 (N_2427,N_1369,N_1373);
nor U2428 (N_2428,In_3916,In_1322);
nand U2429 (N_2429,N_1637,N_619);
nand U2430 (N_2430,N_830,In_2303);
xnor U2431 (N_2431,N_1724,In_1240);
nand U2432 (N_2432,N_1825,In_3326);
xnor U2433 (N_2433,In_4736,In_1413);
nor U2434 (N_2434,In_1121,N_1608);
nor U2435 (N_2435,N_1105,In_2440);
xnor U2436 (N_2436,N_1025,N_474);
and U2437 (N_2437,N_1867,In_3595);
and U2438 (N_2438,In_3627,N_1923);
nand U2439 (N_2439,In_3106,In_3645);
and U2440 (N_2440,N_1530,N_1956);
nand U2441 (N_2441,In_1894,In_3203);
nand U2442 (N_2442,N_1251,In_4727);
nor U2443 (N_2443,In_2735,N_1839);
and U2444 (N_2444,N_1546,In_3714);
xnor U2445 (N_2445,N_1296,In_3519);
xnor U2446 (N_2446,In_4506,In_672);
xor U2447 (N_2447,N_1174,N_577);
xnor U2448 (N_2448,N_1314,In_2908);
xnor U2449 (N_2449,In_3911,In_1513);
nor U2450 (N_2450,N_676,In_1560);
or U2451 (N_2451,N_239,N_1732);
nor U2452 (N_2452,N_1857,N_1844);
and U2453 (N_2453,N_0,In_804);
and U2454 (N_2454,N_635,N_1451);
and U2455 (N_2455,N_1619,In_768);
nor U2456 (N_2456,In_1716,In_1668);
nand U2457 (N_2457,In_2524,In_2654);
and U2458 (N_2458,In_4816,In_3535);
or U2459 (N_2459,In_4698,N_1421);
nand U2460 (N_2460,N_1912,N_1564);
or U2461 (N_2461,N_1818,N_1270);
xnor U2462 (N_2462,N_1738,In_2808);
xnor U2463 (N_2463,In_1400,In_4481);
nor U2464 (N_2464,N_1206,In_927);
xnor U2465 (N_2465,N_1937,N_1754);
xor U2466 (N_2466,In_1074,In_2260);
nor U2467 (N_2467,N_1582,N_1157);
or U2468 (N_2468,N_1304,N_1704);
or U2469 (N_2469,In_654,In_1263);
and U2470 (N_2470,N_1566,In_4024);
xor U2471 (N_2471,N_1129,N_162);
xor U2472 (N_2472,N_1083,N_1407);
xnor U2473 (N_2473,In_1326,N_1491);
xnor U2474 (N_2474,In_111,In_717);
and U2475 (N_2475,N_1450,N_157);
and U2476 (N_2476,In_4149,N_131);
nand U2477 (N_2477,N_1110,N_1418);
xor U2478 (N_2478,In_1089,In_1521);
xnor U2479 (N_2479,N_1188,N_736);
and U2480 (N_2480,In_4651,In_1228);
nand U2481 (N_2481,In_3192,In_3210);
nor U2482 (N_2482,In_1658,N_1405);
xor U2483 (N_2483,In_1889,In_903);
nor U2484 (N_2484,N_1484,In_2071);
or U2485 (N_2485,In_1992,N_833);
or U2486 (N_2486,In_4812,N_1376);
or U2487 (N_2487,N_1799,N_378);
xor U2488 (N_2488,In_2290,N_1962);
and U2489 (N_2489,In_32,N_1106);
nor U2490 (N_2490,N_1809,In_3779);
nor U2491 (N_2491,In_1455,N_1128);
nand U2492 (N_2492,In_4383,In_963);
nor U2493 (N_2493,N_1384,In_2638);
and U2494 (N_2494,In_4892,N_1492);
xor U2495 (N_2495,In_1659,In_839);
xor U2496 (N_2496,N_564,In_2158);
xor U2497 (N_2497,In_2064,In_3537);
nor U2498 (N_2498,In_465,In_2550);
nor U2499 (N_2499,In_1842,In_2008);
nor U2500 (N_2500,N_1749,In_2101);
nand U2501 (N_2501,In_294,N_743);
xnor U2502 (N_2502,In_437,N_351);
nor U2503 (N_2503,In_4545,In_916);
and U2504 (N_2504,In_1691,In_981);
and U2505 (N_2505,In_4775,In_1744);
or U2506 (N_2506,N_296,In_2040);
nor U2507 (N_2507,N_1272,In_709);
and U2508 (N_2508,N_1634,In_2773);
or U2509 (N_2509,N_370,In_445);
nor U2510 (N_2510,N_849,In_2463);
nor U2511 (N_2511,N_1663,In_3082);
nor U2512 (N_2512,N_1478,In_3732);
nand U2513 (N_2513,In_3384,In_3689);
nand U2514 (N_2514,In_4794,In_2936);
nor U2515 (N_2515,N_1746,N_1713);
nor U2516 (N_2516,In_4553,N_318);
nand U2517 (N_2517,N_1792,N_1794);
nand U2518 (N_2518,N_1166,N_1985);
and U2519 (N_2519,N_41,N_1062);
or U2520 (N_2520,In_1949,In_4672);
nand U2521 (N_2521,In_1357,In_3875);
or U2522 (N_2522,In_1013,In_2412);
nor U2523 (N_2523,In_2042,N_1476);
and U2524 (N_2524,N_1018,N_1002);
nand U2525 (N_2525,In_2905,In_127);
xnor U2526 (N_2526,N_1159,In_4584);
nor U2527 (N_2527,N_1786,In_1806);
and U2528 (N_2528,N_1908,N_1108);
nor U2529 (N_2529,In_4300,In_4096);
or U2530 (N_2530,N_291,In_3142);
or U2531 (N_2531,N_1268,In_697);
xor U2532 (N_2532,N_1248,N_1162);
and U2533 (N_2533,In_875,N_465);
nor U2534 (N_2534,In_3608,N_1639);
and U2535 (N_2535,N_1759,N_587);
nand U2536 (N_2536,In_3212,N_1092);
nor U2537 (N_2537,In_1183,N_267);
nand U2538 (N_2538,In_1724,In_2590);
nand U2539 (N_2539,N_1445,N_1289);
or U2540 (N_2540,In_972,N_432);
nor U2541 (N_2541,N_598,N_1941);
nand U2542 (N_2542,In_2984,N_982);
or U2543 (N_2543,N_1363,In_3583);
xnor U2544 (N_2544,In_1436,In_1574);
or U2545 (N_2545,In_982,N_1991);
xnor U2546 (N_2546,N_114,In_2612);
nor U2547 (N_2547,In_3041,In_395);
nand U2548 (N_2548,N_1333,N_1536);
nand U2549 (N_2549,In_1408,In_4827);
nor U2550 (N_2550,N_604,N_1720);
nor U2551 (N_2551,In_1381,N_1250);
and U2552 (N_2552,In_1670,In_3840);
xnor U2553 (N_2553,In_1238,In_4694);
nor U2554 (N_2554,In_782,In_870);
nand U2555 (N_2555,In_4602,In_2449);
nand U2556 (N_2556,In_3081,N_1753);
or U2557 (N_2557,In_543,N_1124);
or U2558 (N_2558,N_1444,In_3818);
nand U2559 (N_2559,N_1350,In_1619);
or U2560 (N_2560,N_335,N_1288);
and U2561 (N_2561,In_3853,In_3314);
nand U2562 (N_2562,In_4722,N_384);
xnor U2563 (N_2563,In_353,N_480);
and U2564 (N_2564,In_992,In_863);
or U2565 (N_2565,N_1918,N_382);
xnor U2566 (N_2566,In_4594,In_536);
nand U2567 (N_2567,N_1218,N_1865);
nand U2568 (N_2568,In_1805,N_1523);
xnor U2569 (N_2569,In_3291,In_316);
xor U2570 (N_2570,In_1000,N_61);
xnor U2571 (N_2571,In_2073,N_950);
and U2572 (N_2572,N_991,N_1855);
and U2573 (N_2573,In_4503,N_1394);
or U2574 (N_2574,In_1579,N_284);
xnor U2575 (N_2575,In_1411,N_1838);
and U2576 (N_2576,In_4361,N_1413);
nand U2577 (N_2577,N_1623,N_445);
or U2578 (N_2578,In_469,In_396);
nand U2579 (N_2579,N_689,N_1781);
and U2580 (N_2580,In_1913,In_1586);
or U2581 (N_2581,N_1047,In_4720);
and U2582 (N_2582,In_2992,N_584);
or U2583 (N_2583,N_7,In_2372);
nand U2584 (N_2584,N_1719,N_1847);
or U2585 (N_2585,In_1721,N_1170);
xor U2586 (N_2586,N_1273,In_3700);
or U2587 (N_2587,In_2702,In_2699);
nand U2588 (N_2588,In_1788,N_1716);
xnor U2589 (N_2589,N_1557,N_1853);
or U2590 (N_2590,N_1474,In_702);
or U2591 (N_2591,In_3850,N_1221);
nor U2592 (N_2592,N_238,N_1259);
nor U2593 (N_2593,In_2127,N_220);
nor U2594 (N_2594,N_483,In_4919);
xor U2595 (N_2595,N_1171,N_502);
nor U2596 (N_2596,N_746,In_1958);
and U2597 (N_2597,In_1044,In_2705);
xor U2598 (N_2598,N_1656,In_4419);
and U2599 (N_2599,N_1229,In_4077);
nor U2600 (N_2600,In_1284,N_491);
xor U2601 (N_2601,N_1587,In_2301);
nand U2602 (N_2602,In_1458,N_1643);
nand U2603 (N_2603,In_4480,In_2287);
nand U2604 (N_2604,In_248,In_3039);
or U2605 (N_2605,In_3186,In_3909);
nor U2606 (N_2606,N_1999,N_714);
or U2607 (N_2607,In_3247,In_3665);
or U2608 (N_2608,In_3890,N_1563);
or U2609 (N_2609,In_4866,N_710);
nor U2610 (N_2610,N_1004,N_458);
and U2611 (N_2611,N_462,N_504);
xnor U2612 (N_2612,In_2736,In_3598);
xnor U2613 (N_2613,N_80,N_67);
or U2614 (N_2614,N_1934,N_1628);
nand U2615 (N_2615,N_1655,In_1405);
or U2616 (N_2616,N_197,N_788);
nand U2617 (N_2617,N_1153,In_3351);
nor U2618 (N_2618,In_3418,N_1616);
xor U2619 (N_2619,In_814,In_3342);
xor U2620 (N_2620,In_3341,N_1773);
or U2621 (N_2621,N_1630,In_648);
nor U2622 (N_2622,In_4250,In_778);
xor U2623 (N_2623,In_3859,In_3363);
xor U2624 (N_2624,In_3050,N_280);
nor U2625 (N_2625,In_4877,N_205);
nand U2626 (N_2626,N_723,In_3056);
xnor U2627 (N_2627,N_360,In_1653);
or U2628 (N_2628,N_1606,N_1645);
or U2629 (N_2629,N_1152,N_1);
xor U2630 (N_2630,In_1233,N_1590);
or U2631 (N_2631,In_2002,In_1643);
and U2632 (N_2632,In_3157,N_1607);
xor U2633 (N_2633,N_390,In_4558);
and U2634 (N_2634,N_1631,In_2226);
nor U2635 (N_2635,In_1952,N_1480);
or U2636 (N_2636,N_1337,N_48);
and U2637 (N_2637,In_1285,In_1178);
and U2638 (N_2638,N_1386,In_3393);
xor U2639 (N_2639,In_2078,In_3776);
nor U2640 (N_2640,In_788,N_1258);
and U2641 (N_2641,N_1286,In_3474);
nor U2642 (N_2642,In_226,In_4090);
nor U2643 (N_2643,N_1549,In_4882);
or U2644 (N_2644,N_156,N_1502);
nor U2645 (N_2645,In_3735,In_1278);
nor U2646 (N_2646,N_1581,In_914);
and U2647 (N_2647,In_4083,In_4013);
and U2648 (N_2648,N_1980,In_1794);
xor U2649 (N_2649,In_2706,N_1885);
and U2650 (N_2650,N_1046,In_3913);
and U2651 (N_2651,N_1230,In_1989);
nand U2652 (N_2652,In_2236,N_63);
nor U2653 (N_2653,N_644,N_606);
and U2654 (N_2654,N_1007,N_1772);
xnor U2655 (N_2655,In_4779,N_557);
or U2656 (N_2656,In_2957,In_4995);
and U2657 (N_2657,N_1199,In_890);
and U2658 (N_2658,In_4115,In_2316);
and U2659 (N_2659,In_4941,N_1496);
or U2660 (N_2660,In_2147,In_3443);
nand U2661 (N_2661,N_952,N_1835);
and U2662 (N_2662,N_1065,In_1151);
nor U2663 (N_2663,In_652,N_302);
xnor U2664 (N_2664,In_4188,N_1294);
nand U2665 (N_2665,N_717,N_1696);
xor U2666 (N_2666,In_2300,In_3740);
nor U2667 (N_2667,In_1953,In_561);
and U2668 (N_2668,N_1266,In_3744);
nand U2669 (N_2669,N_884,In_1702);
xor U2670 (N_2670,In_3374,N_486);
or U2671 (N_2671,N_1693,N_1935);
nor U2672 (N_2672,In_1707,In_2250);
nand U2673 (N_2673,In_3358,In_307);
xnor U2674 (N_2674,In_4711,N_659);
nor U2675 (N_2675,In_1577,In_3078);
nand U2676 (N_2676,In_703,N_493);
nand U2677 (N_2677,N_99,In_2672);
xor U2678 (N_2678,N_589,N_1666);
xor U2679 (N_2679,In_4961,In_1676);
and U2680 (N_2680,N_31,In_1020);
or U2681 (N_2681,N_1668,N_1096);
nand U2682 (N_2682,In_2971,N_1297);
nand U2683 (N_2683,N_1967,N_1226);
or U2684 (N_2684,N_202,In_2335);
nand U2685 (N_2685,N_1305,N_1060);
xor U2686 (N_2686,N_905,N_1493);
and U2687 (N_2687,In_1490,N_264);
nor U2688 (N_2688,N_1506,In_391);
nor U2689 (N_2689,In_3066,In_15);
or U2690 (N_2690,N_1121,N_873);
nand U2691 (N_2691,In_4695,N_1933);
xnor U2692 (N_2692,In_409,In_10);
xor U2693 (N_2693,In_794,N_1929);
and U2694 (N_2694,In_4053,N_894);
and U2695 (N_2695,In_1583,In_3424);
nor U2696 (N_2696,N_1883,In_1804);
nor U2697 (N_2697,N_1470,In_2592);
and U2698 (N_2698,In_1340,In_2069);
or U2699 (N_2699,In_1740,In_4299);
nand U2700 (N_2700,In_4876,In_1376);
xor U2701 (N_2701,N_1190,N_1877);
nand U2702 (N_2702,In_2692,N_1411);
or U2703 (N_2703,In_4641,In_3329);
or U2704 (N_2704,N_1136,In_3490);
and U2705 (N_2705,N_1761,N_1469);
nand U2706 (N_2706,N_1514,N_126);
or U2707 (N_2707,In_1817,N_95);
nor U2708 (N_2708,N_724,N_1067);
nand U2709 (N_2709,In_970,N_1280);
nor U2710 (N_2710,In_4658,In_3396);
or U2711 (N_2711,N_1271,N_1657);
nand U2712 (N_2712,N_1051,N_1736);
and U2713 (N_2713,N_1852,N_1760);
and U2714 (N_2714,N_1005,N_1681);
and U2715 (N_2715,In_3839,N_621);
and U2716 (N_2716,In_2932,In_1245);
nor U2717 (N_2717,In_4234,In_4599);
or U2718 (N_2718,In_894,N_1049);
nand U2719 (N_2719,In_3647,N_1813);
nand U2720 (N_2720,In_4172,In_605);
and U2721 (N_2721,In_3405,N_1836);
or U2722 (N_2722,N_1412,In_1164);
xor U2723 (N_2723,In_4423,In_4755);
or U2724 (N_2724,N_1160,N_1994);
nand U2725 (N_2725,N_1807,In_2190);
xor U2726 (N_2726,N_1313,In_1385);
and U2727 (N_2727,N_1723,In_2052);
xnor U2728 (N_2728,N_70,In_4992);
nor U2729 (N_2729,In_2560,N_358);
nand U2730 (N_2730,N_1135,In_4689);
nand U2731 (N_2731,N_1284,In_1656);
and U2732 (N_2732,In_4254,In_4391);
and U2733 (N_2733,N_1285,N_1058);
nand U2734 (N_2734,In_579,N_1443);
or U2735 (N_2735,N_1729,N_1950);
and U2736 (N_2736,In_2338,N_926);
and U2737 (N_2737,In_1970,N_148);
or U2738 (N_2738,In_4407,In_2953);
nand U2739 (N_2739,N_1750,N_1763);
nand U2740 (N_2740,N_1866,In_2520);
and U2741 (N_2741,N_16,N_1651);
or U2742 (N_2742,N_656,N_1680);
nand U2743 (N_2743,In_1780,N_1123);
and U2744 (N_2744,N_1076,N_118);
or U2745 (N_2745,N_1329,In_390);
or U2746 (N_2746,N_1410,In_4686);
or U2747 (N_2747,In_798,N_1003);
nor U2748 (N_2748,In_2605,In_4896);
nor U2749 (N_2749,N_661,N_210);
nand U2750 (N_2750,N_266,N_389);
and U2751 (N_2751,N_1905,In_3013);
nor U2752 (N_2752,N_1428,N_1895);
nor U2753 (N_2753,N_1574,In_1274);
and U2754 (N_2754,N_760,In_3380);
and U2755 (N_2755,N_1591,In_4552);
nand U2756 (N_2756,In_737,N_1064);
xnor U2757 (N_2757,N_1109,N_1520);
xnor U2758 (N_2758,N_1926,N_1149);
nand U2759 (N_2759,N_774,N_218);
and U2760 (N_2760,N_100,In_2482);
and U2761 (N_2761,N_1100,In_4614);
and U2762 (N_2762,N_1425,N_1942);
xor U2763 (N_2763,In_2740,In_4830);
and U2764 (N_2764,In_4763,In_1601);
and U2765 (N_2765,In_3276,N_1503);
and U2766 (N_2766,In_3906,N_1101);
or U2767 (N_2767,In_2065,In_3308);
or U2768 (N_2768,In_2938,In_4986);
nor U2769 (N_2769,In_3650,In_3483);
and U2770 (N_2770,N_1365,N_1642);
or U2771 (N_2771,In_3712,In_4065);
xor U2772 (N_2772,N_461,In_3773);
nand U2773 (N_2773,N_1161,In_1191);
and U2774 (N_2774,In_274,In_1103);
xor U2775 (N_2775,N_1650,In_4196);
or U2776 (N_2776,N_132,In_273);
and U2777 (N_2777,N_1901,In_2308);
xor U2778 (N_2778,N_1216,N_1821);
and U2779 (N_2779,N_1780,In_2507);
nor U2780 (N_2780,In_686,N_1375);
xor U2781 (N_2781,N_1543,In_2606);
xnor U2782 (N_2782,N_993,N_1367);
nand U2783 (N_2783,N_832,In_4347);
nor U2784 (N_2784,N_1408,N_1200);
xor U2785 (N_2785,In_3306,N_1116);
nand U2786 (N_2786,N_924,N_1789);
nand U2787 (N_2787,In_2630,N_1804);
nand U2788 (N_2788,N_1388,In_1002);
nor U2789 (N_2789,In_505,In_2671);
nor U2790 (N_2790,In_2222,In_1916);
nor U2791 (N_2791,N_1426,In_1868);
nor U2792 (N_2792,N_737,In_222);
and U2793 (N_2793,N_253,In_4661);
or U2794 (N_2794,N_1636,In_3863);
nor U2795 (N_2795,In_757,N_1791);
nor U2796 (N_2796,In_4257,In_4905);
nor U2797 (N_2797,In_4593,In_3183);
xnor U2798 (N_2798,In_2210,N_1130);
nand U2799 (N_2799,In_4274,In_1459);
xor U2800 (N_2800,N_1796,N_1454);
xor U2801 (N_2801,N_1665,N_1466);
nor U2802 (N_2802,N_960,In_4098);
nor U2803 (N_2803,In_868,N_1427);
xnor U2804 (N_2804,In_4014,In_4323);
or U2805 (N_2805,N_1699,N_1419);
nand U2806 (N_2806,In_1236,N_1446);
or U2807 (N_2807,In_3333,N_234);
nand U2808 (N_2808,In_3933,In_2110);
or U2809 (N_2809,In_313,N_293);
nand U2810 (N_2810,In_3130,N_544);
or U2811 (N_2811,N_177,N_45);
nor U2812 (N_2812,In_415,N_1944);
xor U2813 (N_2813,In_3687,In_2712);
and U2814 (N_2814,In_668,N_1868);
nor U2815 (N_2815,In_1297,In_1991);
or U2816 (N_2816,In_4885,N_1358);
and U2817 (N_2817,N_1845,N_146);
xnor U2818 (N_2818,In_3137,In_810);
or U2819 (N_2819,In_2451,N_1559);
nand U2820 (N_2820,In_2741,In_3369);
nand U2821 (N_2821,N_1262,N_1843);
or U2822 (N_2822,In_4420,In_2879);
xnor U2823 (N_2823,N_57,In_710);
xor U2824 (N_2824,N_1507,N_1277);
and U2825 (N_2825,N_1535,N_1770);
and U2826 (N_2826,In_2668,N_795);
nand U2827 (N_2827,N_836,In_4086);
xor U2828 (N_2828,In_1472,N_104);
or U2829 (N_2829,In_1664,N_1414);
nand U2830 (N_2830,N_807,In_1414);
xnor U2831 (N_2831,In_1891,In_3578);
xor U2832 (N_2832,In_3149,In_4529);
xnor U2833 (N_2833,N_1112,In_175);
nor U2834 (N_2834,N_1275,In_1254);
nor U2835 (N_2835,In_4685,N_1856);
and U2836 (N_2836,In_1961,In_1719);
nand U2837 (N_2837,In_77,N_935);
nand U2838 (N_2838,In_2068,N_978);
nand U2839 (N_2839,In_2381,N_1611);
nor U2840 (N_2840,In_4359,In_3421);
and U2841 (N_2841,In_4640,N_1801);
or U2842 (N_2842,N_326,In_172);
or U2843 (N_2843,N_645,N_541);
xor U2844 (N_2844,In_3042,N_581);
nand U2845 (N_2845,N_1684,N_1778);
nor U2846 (N_2846,N_702,In_791);
nor U2847 (N_2847,N_62,N_1006);
nand U2848 (N_2848,N_1040,In_2960);
nand U2849 (N_2849,N_1181,N_1107);
xor U2850 (N_2850,N_1671,N_4);
and U2851 (N_2851,In_1887,In_497);
nor U2852 (N_2852,N_1449,N_1646);
and U2853 (N_2853,N_732,In_3484);
and U2854 (N_2854,N_1177,N_1077);
nand U2855 (N_2855,N_865,N_1165);
xnor U2856 (N_2856,N_829,N_1551);
and U2857 (N_2857,N_855,In_2993);
nor U2858 (N_2858,N_1023,N_1688);
xor U2859 (N_2859,N_572,N_1752);
nand U2860 (N_2860,In_3334,In_3591);
or U2861 (N_2861,In_3833,In_4051);
and U2862 (N_2862,N_1695,N_666);
or U2863 (N_2863,In_2368,In_1430);
xnor U2864 (N_2864,N_1338,N_1690);
nor U2865 (N_2865,In_2189,N_1340);
nor U2866 (N_2866,N_217,N_1977);
and U2867 (N_2867,N_510,In_3231);
nand U2868 (N_2868,In_3309,N_1542);
or U2869 (N_2869,In_1941,N_1197);
xor U2870 (N_2870,In_3029,In_1874);
nand U2871 (N_2871,N_887,N_1764);
and U2872 (N_2872,In_2007,N_1377);
nand U2873 (N_2873,N_1080,N_1070);
or U2874 (N_2874,In_3717,In_4837);
nand U2875 (N_2875,In_1466,In_4860);
nand U2876 (N_2876,N_1534,In_1629);
xor U2877 (N_2877,In_4730,N_1911);
or U2878 (N_2878,N_1015,In_3270);
nor U2879 (N_2879,N_86,In_4851);
xnor U2880 (N_2880,In_4281,N_1127);
or U2881 (N_2881,In_4855,In_365);
and U2882 (N_2882,In_3801,In_4623);
nand U2883 (N_2883,In_3803,N_1823);
nand U2884 (N_2884,N_1378,In_4340);
xor U2885 (N_2885,In_538,In_4338);
or U2886 (N_2886,N_1610,In_2622);
xnor U2887 (N_2887,In_2414,In_1553);
or U2888 (N_2888,In_1066,In_2428);
or U2889 (N_2889,In_1809,In_3826);
nor U2890 (N_2890,In_2800,In_824);
or U2891 (N_2891,In_402,N_848);
and U2892 (N_2892,In_2123,N_487);
or U2893 (N_2893,N_425,In_3990);
or U2894 (N_2894,In_1193,In_2247);
and U2895 (N_2895,In_3774,N_1021);
and U2896 (N_2896,N_967,In_2194);
or U2897 (N_2897,N_677,N_1186);
and U2898 (N_2898,In_1612,In_3267);
nand U2899 (N_2899,N_1339,In_3896);
or U2900 (N_2900,N_1777,In_1525);
nand U2901 (N_2901,N_831,In_1196);
or U2902 (N_2902,In_101,N_1997);
xnor U2903 (N_2903,N_1758,N_845);
nor U2904 (N_2904,In_1404,N_1114);
nor U2905 (N_2905,N_1431,In_2030);
and U2906 (N_2906,In_1273,N_734);
nand U2907 (N_2907,In_1052,N_1036);
nand U2908 (N_2908,N_1219,N_1837);
and U2909 (N_2909,In_2556,N_1864);
nor U2910 (N_2910,N_1601,N_1429);
and U2911 (N_2911,N_1094,In_4183);
xor U2912 (N_2912,N_182,In_4374);
nand U2913 (N_2913,N_650,N_1370);
xor U2914 (N_2914,In_4321,N_229);
or U2915 (N_2915,N_506,In_1602);
and U2916 (N_2916,In_2594,In_1589);
xnor U2917 (N_2917,N_1828,In_3061);
nor U2918 (N_2918,In_4561,N_1892);
nor U2919 (N_2919,N_1227,In_4933);
and U2920 (N_2920,In_977,In_4372);
or U2921 (N_2921,N_1463,N_276);
nor U2922 (N_2922,N_1597,N_1331);
or U2923 (N_2923,N_1217,N_1876);
nor U2924 (N_2924,In_2850,In_3440);
nor U2925 (N_2925,N_1633,N_1805);
or U2926 (N_2926,N_1185,In_4731);
or U2927 (N_2927,In_3206,N_1301);
or U2928 (N_2928,N_1382,N_1898);
or U2929 (N_2929,In_14,N_1958);
and U2930 (N_2930,In_4263,N_366);
nor U2931 (N_2931,In_3242,N_585);
nor U2932 (N_2932,N_1235,In_2249);
nand U2933 (N_2933,N_1739,In_2862);
and U2934 (N_2934,In_1488,N_688);
or U2935 (N_2935,In_772,N_424);
nor U2936 (N_2936,In_4223,N_817);
and U2937 (N_2937,N_1902,In_4322);
xnor U2938 (N_2938,N_1183,N_1319);
xor U2939 (N_2939,In_72,In_3847);
and U2940 (N_2940,N_1417,N_1113);
or U2941 (N_2941,In_4781,In_2193);
xor U2942 (N_2942,N_1609,In_808);
nand U2943 (N_2943,In_1540,In_209);
or U2944 (N_2944,N_1456,In_1382);
nor U2945 (N_2945,N_599,In_2255);
nor U2946 (N_2946,In_822,In_4197);
nor U2947 (N_2947,In_4081,N_327);
xnor U2948 (N_2948,In_3347,In_4029);
or U2949 (N_2949,N_1187,N_283);
and U2950 (N_2950,N_1959,In_4581);
xnor U2951 (N_2951,N_878,In_2382);
and U2952 (N_2952,In_382,N_1893);
xor U2953 (N_2953,N_1328,In_1075);
or U2954 (N_2954,N_1095,N_1318);
nand U2955 (N_2955,N_1725,N_1685);
and U2956 (N_2956,N_1762,In_4538);
xnor U2957 (N_2957,In_3464,In_3747);
nor U2958 (N_2958,In_4625,N_1233);
nor U2959 (N_2959,In_3044,In_4843);
nor U2960 (N_2960,In_1708,In_540);
nor U2961 (N_2961,In_4127,N_1292);
nand U2962 (N_2962,N_328,N_939);
and U2963 (N_2963,N_1352,N_1518);
nor U2964 (N_2964,N_290,In_1300);
or U2965 (N_2965,N_1208,In_4956);
or U2966 (N_2966,N_1755,N_663);
nor U2967 (N_2967,N_200,In_3680);
nand U2968 (N_2968,N_367,In_3977);
nor U2969 (N_2969,In_1807,N_1714);
or U2970 (N_2970,In_1931,N_1545);
and U2971 (N_2971,In_3383,In_4277);
nor U2972 (N_2972,N_117,N_277);
nor U2973 (N_2973,N_232,In_933);
or U2974 (N_2974,In_1253,N_1949);
nand U2975 (N_2975,N_1316,N_1914);
or U2976 (N_2976,In_4676,N_1097);
and U2977 (N_2977,In_3002,N_1930);
and U2978 (N_2978,N_1513,N_1981);
or U2979 (N_2979,In_401,N_1742);
or U2980 (N_2980,N_1978,N_1490);
nand U2981 (N_2981,In_896,In_3943);
nor U2982 (N_2982,In_3120,N_1164);
or U2983 (N_2983,In_261,In_976);
and U2984 (N_2984,N_1494,In_323);
nor U2985 (N_2985,N_1420,In_1644);
xnor U2986 (N_2986,N_785,N_233);
and U2987 (N_2987,N_972,N_1368);
and U2988 (N_2988,N_1374,N_641);
nand U2989 (N_2989,N_1938,N_1795);
or U2990 (N_2990,N_1453,In_2707);
or U2991 (N_2991,In_3626,In_1001);
nand U2992 (N_2992,In_427,N_1508);
xor U2993 (N_2993,N_1679,In_1526);
or U2994 (N_2994,In_4114,N_1323);
and U2995 (N_2995,N_1751,In_3587);
nand U2996 (N_2996,In_4645,N_369);
nor U2997 (N_2997,N_1913,In_432);
or U2998 (N_2998,N_1532,In_3725);
nand U2999 (N_2999,In_666,In_163);
nand U3000 (N_3000,In_1440,In_2435);
xnor U3001 (N_3001,N_2946,N_2500);
or U3002 (N_3002,In_899,In_2271);
or U3003 (N_3003,N_1528,N_2109);
xor U3004 (N_3004,N_2814,N_1703);
or U3005 (N_3005,In_4451,N_2625);
or U3006 (N_3006,N_2132,N_2268);
nand U3007 (N_3007,In_755,N_2118);
nor U3008 (N_3008,N_2530,N_2590);
xor U3009 (N_3009,N_1438,In_3515);
or U3010 (N_3010,N_2977,N_2702);
nor U3011 (N_3011,N_341,N_1579);
or U3012 (N_3012,N_1068,N_2348);
xnor U3013 (N_3013,N_1014,In_107);
or U3014 (N_3014,N_1576,In_2192);
nand U3015 (N_3015,N_2362,N_2012);
and U3016 (N_3016,N_2293,In_4488);
nand U3017 (N_3017,N_1603,N_2235);
and U3018 (N_3018,N_2257,N_2954);
nand U3019 (N_3019,N_2712,N_2422);
nand U3020 (N_3020,N_2470,In_4095);
nor U3021 (N_3021,In_4151,In_4208);
xor U3022 (N_3022,N_2332,In_3959);
nand U3023 (N_3023,In_4932,In_2125);
xnor U3024 (N_3024,N_2808,N_2159);
nor U3025 (N_3025,N_2369,N_2722);
xor U3026 (N_3026,N_2713,In_238);
xor U3027 (N_3027,N_2769,N_49);
and U3028 (N_3028,In_3889,N_2577);
and U3029 (N_3029,N_2544,In_2988);
nand U3030 (N_3030,N_344,N_2);
or U3031 (N_3031,In_3506,N_2565);
and U3032 (N_3032,In_4030,N_2220);
nand U3033 (N_3033,In_4431,N_1089);
and U3034 (N_3034,N_756,N_2481);
xor U3035 (N_3035,N_2718,N_2998);
nand U3036 (N_3036,N_2630,N_2936);
and U3037 (N_3037,N_2934,N_2908);
xnor U3038 (N_3038,N_2974,In_311);
xnor U3039 (N_3039,N_392,N_2071);
nand U3040 (N_3040,N_1099,N_2401);
nor U3041 (N_3041,In_1841,N_2046);
nand U3042 (N_3042,N_814,N_1768);
xnor U3043 (N_3043,N_222,In_687);
and U3044 (N_3044,N_2709,In_4471);
xor U3045 (N_3045,In_3510,N_470);
nand U3046 (N_3046,N_2927,N_2999);
or U3047 (N_3047,N_2136,N_2069);
or U3048 (N_3048,N_2177,In_4416);
and U3049 (N_3049,N_476,N_2850);
xnor U3050 (N_3050,N_1955,N_1640);
xor U3051 (N_3051,N_2230,N_1327);
and U3052 (N_3052,In_4612,N_418);
and U3053 (N_3053,N_2346,N_2738);
or U3054 (N_3054,N_652,In_2083);
xnor U3055 (N_3055,N_2635,N_1712);
nor U3056 (N_3056,In_1866,N_2626);
nor U3057 (N_3057,N_2810,N_2823);
nor U3058 (N_3058,In_1758,N_2677);
xor U3059 (N_3059,N_2949,N_2706);
or U3060 (N_3060,N_2964,N_2110);
xnor U3061 (N_3061,N_2993,N_2940);
or U3062 (N_3062,N_1052,N_1348);
xor U3063 (N_3063,N_862,N_460);
and U3064 (N_3064,In_1444,N_634);
and U3065 (N_3065,In_3436,In_4997);
nor U3066 (N_3066,In_4960,N_2224);
xnor U3067 (N_3067,In_4675,N_741);
xnor U3068 (N_3068,N_2360,In_624);
xnor U3069 (N_3069,In_4683,N_2859);
or U3070 (N_3070,N_2131,N_1300);
and U3071 (N_3071,In_4512,N_2778);
nor U3072 (N_3072,N_2137,N_2549);
nor U3073 (N_3073,N_2863,In_1287);
nand U3074 (N_3074,N_1309,N_1126);
or U3075 (N_3075,N_2009,N_2391);
nor U3076 (N_3076,N_2407,N_2800);
and U3077 (N_3077,In_3129,N_2248);
or U3078 (N_3078,N_2700,In_3802);
and U3079 (N_3079,N_2397,In_4455);
or U3080 (N_3080,N_1808,N_2002);
and U3081 (N_3081,N_2897,In_2749);
and U3082 (N_3082,N_2414,In_3088);
nand U3083 (N_3083,N_1827,In_452);
nor U3084 (N_3084,N_2318,In_544);
nor U3085 (N_3085,N_1660,N_759);
or U3086 (N_3086,N_2689,N_2723);
and U3087 (N_3087,N_2316,N_2535);
and U3088 (N_3088,N_2729,N_2184);
and U3089 (N_3089,N_2795,N_2153);
nand U3090 (N_3090,N_2926,N_2436);
nand U3091 (N_3091,In_47,N_2523);
or U3092 (N_3092,In_4062,N_2539);
xor U3093 (N_3093,N_2796,In_574);
nand U3094 (N_3094,N_1326,In_723);
nor U3095 (N_3095,In_4224,N_2123);
and U3096 (N_3096,N_2969,N_17);
xor U3097 (N_3097,N_2553,In_140);
or U3098 (N_3098,N_2058,N_2668);
nor U3099 (N_3099,N_2849,N_777);
nor U3100 (N_3100,N_2455,N_1341);
or U3101 (N_3101,N_2840,N_2292);
nor U3102 (N_3102,N_2501,N_2653);
xor U3103 (N_3103,In_2425,N_1439);
and U3104 (N_3104,In_2207,N_2824);
xor U3105 (N_3105,N_1140,N_1556);
nand U3106 (N_3106,N_2512,N_2766);
and U3107 (N_3107,In_1395,N_597);
xnor U3108 (N_3108,N_1322,N_1924);
nor U3109 (N_3109,N_2338,N_769);
or U3110 (N_3110,N_2191,N_2865);
or U3111 (N_3111,N_1931,N_2327);
and U3112 (N_3112,N_2475,N_1600);
or U3113 (N_3113,N_311,In_2241);
nand U3114 (N_3114,N_1897,In_334);
and U3115 (N_3115,N_2065,N_2472);
nor U3116 (N_3116,N_1212,In_1863);
and U3117 (N_3117,N_1066,N_2518);
nor U3118 (N_3118,N_2606,N_2167);
and U3119 (N_3119,N_2053,N_2888);
and U3120 (N_3120,N_1575,N_2234);
and U3121 (N_3121,N_2991,N_1330);
or U3122 (N_3122,N_158,N_2531);
nor U3123 (N_3123,In_4436,N_1151);
or U3124 (N_3124,N_2413,N_2787);
xor U3125 (N_3125,N_2351,N_1988);
xnor U3126 (N_3126,In_4642,N_2979);
and U3127 (N_3127,In_1569,N_969);
xor U3128 (N_3128,In_3804,N_2820);
or U3129 (N_3129,N_2922,N_1459);
nand U3130 (N_3130,N_2243,N_2169);
xor U3131 (N_3131,N_2704,N_1379);
and U3132 (N_3132,N_2114,N_1147);
and U3133 (N_3133,N_2563,N_1011);
nor U3134 (N_3134,N_2396,In_4580);
and U3135 (N_3135,In_1177,N_2152);
and U3136 (N_3136,N_1629,N_1757);
nand U3137 (N_3137,N_115,N_2572);
xor U3138 (N_3138,In_4074,N_2048);
nor U3139 (N_3139,N_866,N_1082);
nand U3140 (N_3140,N_917,In_4202);
xor U3141 (N_3141,N_2067,In_3932);
and U3142 (N_3142,N_1652,N_2102);
and U3143 (N_3143,N_2162,N_691);
and U3144 (N_3144,N_1293,N_1245);
xnor U3145 (N_3145,N_1457,In_3080);
xnor U3146 (N_3146,N_2247,In_1511);
and U3147 (N_3147,N_2072,N_2879);
and U3148 (N_3148,N_861,In_4741);
xor U3149 (N_3149,N_2427,N_1038);
xor U3150 (N_3150,N_2404,N_1361);
or U3151 (N_3151,N_2304,N_2252);
and U3152 (N_3152,In_3286,N_2339);
xor U3153 (N_3153,In_3686,N_2930);
xor U3154 (N_3154,N_2835,N_2957);
nor U3155 (N_3155,N_1256,In_3629);
and U3156 (N_3156,N_1848,N_2774);
and U3157 (N_3157,N_1972,N_2736);
nor U3158 (N_3158,N_963,In_443);
or U3159 (N_3159,N_2955,N_2228);
nand U3160 (N_3160,N_2614,N_2128);
nand U3161 (N_3161,N_2342,In_1723);
or U3162 (N_3162,In_2722,In_4819);
and U3163 (N_3163,N_2066,N_1568);
or U3164 (N_3164,N_1975,N_2833);
or U3165 (N_3165,N_2852,N_947);
and U3166 (N_3166,N_2370,N_1598);
or U3167 (N_3167,In_4769,N_2172);
xnor U3168 (N_3168,N_2803,N_2270);
or U3169 (N_3169,N_2194,N_2694);
or U3170 (N_3170,N_2943,N_2876);
and U3171 (N_3171,N_342,N_2673);
xor U3172 (N_3172,N_1461,In_2826);
nand U3173 (N_3173,In_2559,N_970);
and U3174 (N_3174,N_2459,In_1666);
nor U3175 (N_3175,N_1182,In_3026);
nor U3176 (N_3176,N_1638,N_2749);
xnor U3177 (N_3177,In_362,N_2519);
nand U3178 (N_3178,N_2157,N_2576);
or U3179 (N_3179,In_3465,N_2463);
nor U3180 (N_3180,In_4119,In_1504);
or U3181 (N_3181,N_2621,In_2814);
or U3182 (N_3182,In_1985,N_2851);
nor U3183 (N_3183,In_3545,In_4887);
and U3184 (N_3184,N_213,N_2288);
and U3185 (N_3185,N_2564,N_2209);
nor U3186 (N_3186,N_1017,In_1693);
nor U3187 (N_3187,N_896,In_3459);
and U3188 (N_3188,N_2701,N_2520);
xnor U3189 (N_3189,In_1494,In_2669);
or U3190 (N_3190,N_270,In_1432);
or U3191 (N_3191,N_2450,N_1519);
xor U3192 (N_3192,N_1569,N_2742);
xnor U3193 (N_3193,N_2827,N_1225);
xor U3194 (N_3194,In_3053,N_1527);
nand U3195 (N_3195,N_2000,N_1661);
nor U3196 (N_3196,N_1833,In_1713);
xor U3197 (N_3197,N_2603,N_2885);
nand U3198 (N_3198,N_2403,N_2607);
and U3199 (N_3199,In_2293,N_211);
and U3200 (N_3200,N_2465,N_2959);
nor U3201 (N_3201,N_2664,N_2249);
or U3202 (N_3202,N_2135,N_2557);
or U3203 (N_3203,N_2724,N_2634);
and U3204 (N_3204,N_2924,In_2331);
or U3205 (N_3205,N_2219,N_1468);
nand U3206 (N_3206,N_1072,In_774);
xnor U3207 (N_3207,N_2757,N_2637);
nand U3208 (N_3208,N_2735,N_2570);
nor U3209 (N_3209,N_2663,N_2211);
xnor U3210 (N_3210,N_2605,N_2090);
or U3211 (N_3211,N_2025,N_2439);
and U3212 (N_3212,N_1592,N_1971);
or U3213 (N_3213,N_423,In_1456);
and U3214 (N_3214,N_2649,N_2039);
nand U3215 (N_3215,In_905,N_2035);
or U3216 (N_3216,N_1013,In_3442);
or U3217 (N_3217,N_2720,N_2218);
xor U3218 (N_3218,N_2932,N_1342);
xnor U3219 (N_3219,N_2406,In_950);
xnor U3220 (N_3220,N_2429,In_4893);
or U3221 (N_3221,N_81,N_1091);
or U3222 (N_3222,In_584,N_2585);
and U3223 (N_3223,N_2260,N_2045);
nand U3224 (N_3224,N_1803,N_2027);
nor U3225 (N_3225,N_2290,N_1357);
nor U3226 (N_3226,In_3919,N_1045);
nor U3227 (N_3227,N_2971,In_1778);
and U3228 (N_3228,N_2721,N_1298);
nand U3229 (N_3229,In_4333,N_2264);
xor U3230 (N_3230,N_740,N_2075);
and U3231 (N_3231,N_347,N_2678);
xnor U3232 (N_3232,N_975,In_1443);
nand U3233 (N_3233,N_2716,N_2903);
or U3234 (N_3234,In_2006,N_212);
nand U3235 (N_3235,N_2750,N_2405);
nor U3236 (N_3236,N_2797,N_1842);
nor U3237 (N_3237,N_2907,In_3040);
nor U3238 (N_3238,N_517,N_1702);
and U3239 (N_3239,N_951,N_2441);
nor U3240 (N_3240,N_2302,N_1472);
xnor U3241 (N_3241,N_2461,N_2692);
nor U3242 (N_3242,N_2341,N_2345);
or U3243 (N_3243,N_2811,N_2462);
and U3244 (N_3244,N_2457,N_1061);
and U3245 (N_3245,N_1522,In_4937);
nand U3246 (N_3246,N_2074,In_3015);
nand U3247 (N_3247,In_4759,In_3354);
nand U3248 (N_3248,N_2510,N_2882);
or U3249 (N_3249,N_2225,N_2997);
nor U3250 (N_3250,N_2961,N_2871);
nand U3251 (N_3251,N_2353,N_2430);
nand U3252 (N_3252,N_2313,N_2900);
and U3253 (N_3253,N_1335,N_2371);
and U3254 (N_3254,In_4444,N_2562);
and U3255 (N_3255,N_2261,N_2645);
xor U3256 (N_3256,In_4080,N_463);
nand U3257 (N_3257,N_2412,N_2415);
and U3258 (N_3258,N_786,N_1032);
and U3259 (N_3259,N_2612,N_2085);
and U3260 (N_3260,N_2845,N_2661);
or U3261 (N_3261,N_2581,N_2097);
or U3262 (N_3262,N_2493,N_2654);
nand U3263 (N_3263,In_466,N_2754);
or U3264 (N_3264,In_2112,In_2828);
and U3265 (N_3265,N_1346,N_2596);
or U3266 (N_3266,In_1998,N_2896);
nand U3267 (N_3267,N_2284,N_2502);
nor U3268 (N_3268,N_2324,N_2399);
nand U3269 (N_3269,N_844,In_4265);
nand U3270 (N_3270,N_391,N_2683);
and U3271 (N_3271,N_2005,In_4408);
nor U3272 (N_3272,N_2836,N_2988);
and U3273 (N_3273,N_244,N_2205);
or U3274 (N_3274,In_3763,N_2216);
nand U3275 (N_3275,In_3816,N_1524);
and U3276 (N_3276,N_2420,In_1522);
and U3277 (N_3277,N_2697,N_2307);
or U3278 (N_3278,N_471,In_2947);
nand U3279 (N_3279,N_1953,In_4690);
and U3280 (N_3280,N_2669,In_1507);
and U3281 (N_3281,In_4163,N_2928);
nand U3282 (N_3282,N_2315,N_2124);
nand U3283 (N_3283,N_1641,N_2024);
and U3284 (N_3284,N_2556,In_1231);
or U3285 (N_3285,N_1452,N_2972);
nand U3286 (N_3286,N_2609,N_2294);
nand U3287 (N_3287,N_789,N_1016);
and U3288 (N_3288,In_2050,N_1071);
and U3289 (N_3289,N_2918,N_1596);
or U3290 (N_3290,N_2241,N_2251);
and U3291 (N_3291,In_725,In_4756);
nand U3292 (N_3292,N_2434,In_1099);
or U3293 (N_3293,N_2948,N_1119);
nor U3294 (N_3294,N_1364,N_2745);
or U3295 (N_3295,In_3382,In_694);
and U3296 (N_3296,N_2580,N_2494);
and U3297 (N_3297,In_2766,N_2055);
nor U3298 (N_3298,N_2986,N_2431);
nor U3299 (N_3299,N_1909,In_836);
xor U3300 (N_3300,N_2113,N_2990);
or U3301 (N_3301,N_2788,N_2829);
or U3302 (N_3302,In_4927,N_2171);
or U3303 (N_3303,N_2687,N_2166);
xor U3304 (N_3304,N_2913,N_2210);
nand U3305 (N_3305,N_2286,In_2535);
xnor U3306 (N_3306,N_1436,In_4146);
or U3307 (N_3307,N_2333,In_1973);
xnor U3308 (N_3308,N_68,N_2175);
nor U3309 (N_3309,In_4477,In_889);
xor U3310 (N_3310,N_1356,N_2944);
nor U3311 (N_3311,N_2010,In_2591);
nor U3312 (N_3312,N_2263,N_2533);
or U3313 (N_3313,N_2089,N_2298);
nand U3314 (N_3314,N_2308,N_2299);
nor U3315 (N_3315,N_2041,In_1188);
xnor U3316 (N_3316,N_2376,N_1172);
and U3317 (N_3317,N_1553,N_1894);
xor U3318 (N_3318,N_1561,N_1766);
and U3319 (N_3319,N_2794,N_2658);
and U3320 (N_3320,N_2107,N_2336);
and U3321 (N_3321,N_2340,N_2579);
and U3322 (N_3322,In_3999,N_2967);
nor U3323 (N_3323,N_2213,N_1122);
nor U3324 (N_3324,N_428,N_1485);
nor U3325 (N_3325,N_901,In_3307);
nor U3326 (N_3326,N_2231,N_2834);
nand U3327 (N_3327,N_2792,In_155);
nor U3328 (N_3328,N_754,N_2133);
nor U3329 (N_3329,N_2259,N_1903);
or U3330 (N_3330,In_1546,N_2484);
nand U3331 (N_3331,In_1383,N_2468);
nor U3332 (N_3332,In_511,N_2785);
or U3333 (N_3333,In_4387,N_2756);
nand U3334 (N_3334,N_2477,In_2527);
xor U3335 (N_3335,N_2084,N_2715);
nand U3336 (N_3336,In_3063,N_2378);
xnor U3337 (N_3337,N_1213,N_1682);
nor U3338 (N_3338,In_214,N_2443);
and U3339 (N_3339,N_2509,N_2390);
and U3340 (N_3340,In_1696,N_2536);
xor U3341 (N_3341,N_2984,In_4678);
nor U3342 (N_3342,N_2920,N_2480);
and U3343 (N_3343,N_2670,N_949);
and U3344 (N_3344,N_2242,In_2917);
nand U3345 (N_3345,In_4070,N_26);
xor U3346 (N_3346,In_3915,N_2631);
nand U3347 (N_3347,N_2189,N_2269);
nand U3348 (N_3348,N_2755,N_2828);
xor U3349 (N_3349,N_2120,N_2780);
nor U3350 (N_3350,N_1026,N_2890);
or U3351 (N_3351,N_1669,N_1158);
xnor U3352 (N_3352,N_2179,N_1974);
xor U3353 (N_3353,In_847,N_1440);
and U3354 (N_3354,N_2958,N_1774);
xnor U3355 (N_3355,N_1709,In_707);
or U3356 (N_3356,N_2680,N_1299);
nor U3357 (N_3357,N_2272,N_2633);
nand U3358 (N_3358,N_2945,N_942);
or U3359 (N_3359,N_271,N_457);
nand U3360 (N_3360,N_2573,In_2906);
nand U3361 (N_3361,N_1790,N_2636);
xnor U3362 (N_3362,N_1281,N_2330);
nand U3363 (N_3363,In_1469,In_4874);
and U3364 (N_3364,N_2367,N_1947);
and U3365 (N_3365,N_2597,N_2042);
or U3366 (N_3366,In_4659,N_1920);
and U3367 (N_3367,N_472,N_2887);
or U3368 (N_3368,N_2121,N_1727);
or U3369 (N_3369,N_2916,N_2534);
nand U3370 (N_3370,N_2522,N_2188);
xor U3371 (N_3371,In_969,In_993);
or U3372 (N_3372,N_64,N_1385);
or U3373 (N_3373,N_2693,In_4732);
nand U3374 (N_3374,In_4230,In_732);
nor U3375 (N_3375,N_1195,N_2068);
nor U3376 (N_3376,N_1104,N_1317);
nor U3377 (N_3377,N_1840,N_2466);
nor U3378 (N_3378,N_2950,N_1687);
nand U3379 (N_3379,N_2178,N_2532);
xor U3380 (N_3380,N_2433,In_1537);
nand U3381 (N_3381,N_1184,N_2037);
nor U3382 (N_3382,N_1884,In_3750);
and U3383 (N_3383,N_2648,In_1551);
or U3384 (N_3384,N_1951,N_245);
xor U3385 (N_3385,N_660,N_2542);
or U3386 (N_3386,N_2273,N_2460);
or U3387 (N_3387,In_4105,N_2326);
nand U3388 (N_3388,N_338,N_1515);
or U3389 (N_3389,N_2144,N_2822);
nand U3390 (N_3390,N_2639,N_2710);
nor U3391 (N_3391,N_2176,N_2087);
or U3392 (N_3392,N_1403,In_2690);
xor U3393 (N_3393,N_2690,N_2855);
nor U3394 (N_3394,N_1201,N_2681);
or U3395 (N_3395,In_2056,In_1752);
nor U3396 (N_3396,In_216,N_2951);
nor U3397 (N_3397,In_4809,In_1822);
or U3398 (N_3398,N_2275,N_2499);
or U3399 (N_3399,N_2806,N_2321);
or U3400 (N_3400,N_2163,N_2497);
xnor U3401 (N_3401,In_3272,N_2142);
nor U3402 (N_3402,In_2809,N_2038);
or U3403 (N_3403,In_4155,N_2506);
nand U3404 (N_3404,N_2696,N_11);
or U3405 (N_3405,N_2385,In_3895);
nor U3406 (N_3406,N_1648,In_4097);
nor U3407 (N_3407,N_1832,N_2056);
nand U3408 (N_3408,In_1295,N_2377);
or U3409 (N_3409,In_1633,N_1700);
nor U3410 (N_3410,In_3586,In_3926);
nor U3411 (N_3411,N_336,N_1501);
xnor U3412 (N_3412,N_2125,N_1321);
xor U3413 (N_3413,N_2201,N_2976);
nand U3414 (N_3414,N_2296,N_2985);
nor U3415 (N_3415,N_2591,N_2914);
xnor U3416 (N_3416,N_2995,In_98);
nand U3417 (N_3417,N_2044,N_2846);
and U3418 (N_3418,In_758,N_2598);
nand U3419 (N_3419,N_1570,In_4551);
xor U3420 (N_3420,N_2095,In_4350);
nor U3421 (N_3421,N_2254,N_2064);
nand U3422 (N_3422,In_1004,N_2616);
or U3423 (N_3423,N_2650,N_1030);
nor U3424 (N_3424,N_1740,N_2070);
and U3425 (N_3425,In_3353,N_1390);
and U3426 (N_3426,N_137,In_2243);
nand U3427 (N_3427,N_2015,In_3861);
nand U3428 (N_3428,In_3302,N_2287);
and U3429 (N_3429,N_2186,In_234);
nand U3430 (N_3430,N_1324,N_2148);
nor U3431 (N_3431,In_1482,N_1497);
and U3432 (N_3432,In_4935,N_2655);
nor U3433 (N_3433,N_2350,N_2036);
or U3434 (N_3434,In_24,N_2452);
nand U3435 (N_3435,N_2947,N_2030);
nor U3436 (N_3436,N_2060,In_678);
nor U3437 (N_3437,N_2469,N_2023);
nor U3438 (N_3438,N_1473,N_2996);
nand U3439 (N_3439,In_1214,N_2200);
xnor U3440 (N_3440,N_1028,N_2875);
xor U3441 (N_3441,In_3924,In_4595);
nand U3442 (N_3442,In_4116,N_2595);
and U3443 (N_3443,N_452,N_2098);
nand U3444 (N_3444,In_4006,N_2317);
or U3445 (N_3445,N_1204,N_2380);
nor U3446 (N_3446,N_2831,N_2555);
and U3447 (N_3447,In_3989,N_1899);
and U3448 (N_3448,N_2698,N_1946);
nor U3449 (N_3449,N_2893,N_2111);
and U3450 (N_3450,N_2386,N_1381);
nand U3451 (N_3451,N_1310,N_2108);
and U3452 (N_3452,N_2881,In_2856);
and U3453 (N_3453,N_713,N_2727);
or U3454 (N_3454,N_668,N_2182);
or U3455 (N_3455,N_2022,In_3075);
nor U3456 (N_3456,N_2425,N_2762);
xnor U3457 (N_3457,N_1593,N_842);
or U3458 (N_3458,In_2648,N_2043);
nand U3459 (N_3459,N_2458,N_2357);
and U3460 (N_3460,N_2809,N_918);
nand U3461 (N_3461,In_1169,N_2740);
nand U3462 (N_3462,In_615,In_4181);
nor U3463 (N_3463,N_2325,In_2318);
nor U3464 (N_3464,N_2093,In_1418);
and U3465 (N_3465,In_3870,N_1602);
and U3466 (N_3466,N_2059,N_618);
nand U3467 (N_3467,N_2119,N_2467);
or U3468 (N_3468,N_2868,N_1691);
or U3469 (N_3469,N_2711,In_792);
and U3470 (N_3470,N_1744,N_2032);
nor U3471 (N_3471,N_2909,N_2139);
or U3472 (N_3472,N_624,In_917);
and U3473 (N_3473,N_2620,N_2016);
nand U3474 (N_3474,In_1323,N_1860);
nor U3475 (N_3475,N_590,In_3160);
xor U3476 (N_3476,In_797,N_2842);
nor U3477 (N_3477,In_3005,N_1209);
and U3478 (N_3478,N_890,N_1351);
nand U3479 (N_3479,N_2860,N_2130);
or U3480 (N_3480,N_1087,N_2244);
nor U3481 (N_3481,N_2731,N_2707);
nand U3482 (N_3482,In_468,N_2447);
nand U3483 (N_3483,In_818,N_2393);
xnor U3484 (N_3484,N_2880,N_2610);
xor U3485 (N_3485,N_2438,N_2642);
nand U3486 (N_3486,N_2743,In_3296);
and U3487 (N_3487,In_828,In_160);
xnor U3488 (N_3488,In_4244,N_2847);
nor U3489 (N_3489,N_2323,N_2980);
xor U3490 (N_3490,N_1995,In_4044);
nor U3491 (N_3491,In_4351,In_3264);
nand U3492 (N_3492,In_191,In_4180);
xnor U3493 (N_3493,N_2643,N_2485);
nor U3494 (N_3494,N_2051,N_2528);
and U3495 (N_3495,N_1084,In_3331);
xnor U3496 (N_3496,N_2578,N_2474);
nand U3497 (N_3497,In_1187,N_488);
nand U3498 (N_3498,In_1512,N_1486);
and U3499 (N_3499,N_2233,N_2839);
and U3500 (N_3500,N_1585,N_2684);
or U3501 (N_3501,N_2744,In_3087);
nor U3502 (N_3502,N_816,N_2033);
nor U3503 (N_3503,In_1111,N_2973);
nand U3504 (N_3504,N_2830,N_2117);
xor U3505 (N_3505,In_3991,N_1979);
nand U3506 (N_3506,N_1315,N_2337);
and U3507 (N_3507,N_2526,N_1261);
or U3508 (N_3508,In_3429,In_3566);
and U3509 (N_3509,N_1544,N_1779);
xnor U3510 (N_3510,N_2001,In_786);
nor U3511 (N_3511,N_1056,N_2373);
or U3512 (N_3512,In_2965,In_4884);
xor U3513 (N_3513,N_2073,N_1584);
nand U3514 (N_3514,N_2910,N_2741);
xnor U3515 (N_3515,N_2149,N_708);
nand U3516 (N_3516,N_1812,In_655);
nor U3517 (N_3517,N_2400,N_2608);
nor U3518 (N_3518,N_2552,N_2496);
and U3519 (N_3519,N_977,N_2155);
and U3520 (N_3520,N_2101,In_1213);
nor U3521 (N_3521,In_4139,N_1278);
nand U3522 (N_3522,N_1677,N_2106);
nand U3523 (N_3523,In_1260,In_3625);
and U3524 (N_3524,N_2082,N_1605);
xnor U3525 (N_3525,N_2937,In_806);
xnor U3526 (N_3526,N_2705,N_1604);
or U3527 (N_3527,N_2040,N_2300);
nor U3528 (N_3528,In_3569,In_583);
or U3529 (N_3529,N_2375,In_2721);
or U3530 (N_3530,N_938,In_58);
nor U3531 (N_3531,N_2490,In_3597);
nor U3532 (N_3532,N_2805,N_2250);
and U3533 (N_3533,N_2026,N_441);
and U3534 (N_3534,N_345,In_3632);
or U3535 (N_3535,N_930,N_761);
or U3536 (N_3536,N_2168,N_1345);
or U3537 (N_3537,N_2099,N_1075);
nor U3538 (N_3538,N_1401,N_2586);
xnor U3539 (N_3539,N_665,In_1971);
nor U3540 (N_3540,N_2894,In_488);
nand U3541 (N_3541,N_2511,N_649);
or U3542 (N_3542,In_3962,N_2495);
or U3543 (N_3543,N_2063,N_2615);
xnor U3544 (N_3544,In_3228,N_2418);
nor U3545 (N_3545,N_89,In_4235);
or U3546 (N_3546,N_2517,N_2322);
and U3547 (N_3547,In_3690,In_2186);
nand U3548 (N_3548,N_2619,N_2812);
and U3549 (N_3549,In_3240,N_1904);
and U3550 (N_3550,N_2952,N_2884);
and U3551 (N_3551,N_2568,N_2361);
xnor U3552 (N_3552,In_2054,N_812);
or U3553 (N_3553,N_2236,In_3938);
nor U3554 (N_3554,N_2214,N_2652);
nor U3555 (N_3555,In_2876,In_348);
nor U3556 (N_3556,N_1555,In_2653);
or U3557 (N_3557,N_1906,In_2165);
nor U3558 (N_3558,N_2424,N_421);
xor U3559 (N_3559,N_2238,N_226);
nand U3560 (N_3560,N_2052,N_2164);
nor U3561 (N_3561,N_2212,N_1391);
nand U3562 (N_3562,N_694,N_2145);
nor U3563 (N_3563,In_3327,N_2551);
nand U3564 (N_3564,N_2028,N_2866);
xor U3565 (N_3565,N_1169,N_324);
xnor U3566 (N_3566,In_840,N_2165);
nand U3567 (N_3567,N_1079,N_1932);
nor U3568 (N_3568,In_2376,N_2449);
or U3569 (N_3569,N_2054,In_614);
nand U3570 (N_3570,N_2725,In_1428);
and U3571 (N_3571,N_2221,N_278);
and U3572 (N_3572,N_1220,N_2277);
and U3573 (N_3573,N_2541,N_2057);
nand U3574 (N_3574,N_2328,N_2508);
nor U3575 (N_3575,N_1295,In_4461);
nor U3576 (N_3576,N_29,In_1129);
xor U3577 (N_3577,N_2686,N_2644);
nand U3578 (N_3578,N_2629,N_1203);
and U3579 (N_3579,N_2807,N_1063);
or U3580 (N_3580,N_494,N_962);
or U3581 (N_3581,N_2417,In_763);
or U3582 (N_3582,In_462,N_2207);
nand U3583 (N_3583,N_1771,In_3062);
and U3584 (N_3584,N_1552,N_1694);
xor U3585 (N_3585,N_1455,N_940);
xnor U3586 (N_3586,N_2077,N_1869);
or U3587 (N_3587,In_2179,N_2746);
nor U3588 (N_3588,N_1621,N_2180);
and U3589 (N_3589,In_4697,N_1441);
and U3590 (N_3590,N_2183,N_2994);
or U3591 (N_3591,N_1793,In_1848);
nand U3592 (N_3592,N_2173,N_430);
or U3593 (N_3593,N_2791,N_1214);
and U3594 (N_3594,N_1882,N_2771);
and U3595 (N_3595,N_2227,In_3885);
and U3596 (N_3596,N_2739,N_58);
nor U3597 (N_3597,N_2147,N_2751);
or U3598 (N_3598,N_2892,N_2187);
xor U3599 (N_3599,N_2498,N_2933);
nor U3600 (N_3600,N_1547,N_2942);
or U3601 (N_3601,N_2730,In_829);
xnor U3602 (N_3602,N_2453,In_3849);
nand U3603 (N_3603,N_2574,N_2253);
nor U3604 (N_3604,N_2199,In_1979);
or U3605 (N_3605,N_2019,N_886);
nor U3606 (N_3606,N_2622,In_1113);
and U3607 (N_3607,N_2129,N_2374);
and U3608 (N_3608,N_2657,In_3032);
or U3609 (N_3609,N_765,N_1521);
and U3610 (N_3610,N_2559,N_2618);
and U3611 (N_3611,N_2583,In_3639);
and U3612 (N_3612,N_2877,N_2343);
and U3613 (N_3613,N_2547,In_675);
or U3614 (N_3614,In_919,In_533);
or U3615 (N_3615,N_2813,N_2790);
nand U3616 (N_3616,N_1118,N_2782);
nor U3617 (N_3617,N_1811,N_2861);
nand U3618 (N_3618,N_2899,N_2312);
and U3619 (N_3619,N_2206,N_160);
nand U3620 (N_3620,In_4572,N_1538);
or U3621 (N_3621,N_2982,N_2956);
nor U3622 (N_3622,N_2347,N_1447);
xnor U3623 (N_3623,N_2765,N_2753);
nand U3624 (N_3624,N_2624,N_1180);
nand U3625 (N_3625,N_2368,N_813);
xor U3626 (N_3626,N_315,N_920);
nand U3627 (N_3627,N_1398,N_2915);
or U3628 (N_3628,N_2968,N_1871);
nand U3629 (N_3629,N_2150,N_2874);
xnor U3630 (N_3630,N_2760,In_1962);
and U3631 (N_3631,N_2309,In_1155);
and U3632 (N_3632,N_995,N_1434);
xor U3633 (N_3633,N_1689,N_2676);
and U3634 (N_3634,N_1692,N_2050);
and U3635 (N_3635,In_4279,N_2904);
nor U3636 (N_3636,N_208,N_2305);
nor U3637 (N_3637,In_4757,In_2185);
nand U3638 (N_3638,N_1467,In_1186);
nand U3639 (N_3639,N_2004,N_2978);
nand U3640 (N_3640,In_3376,In_597);
nand U3641 (N_3641,N_2529,In_2976);
or U3642 (N_3642,N_1896,In_2583);
or U3643 (N_3643,In_2132,N_2870);
xnor U3644 (N_3644,In_986,N_2297);
nor U3645 (N_3645,N_1675,N_536);
xnor U3646 (N_3646,N_1873,In_3197);
or U3647 (N_3647,In_1453,N_1389);
xor U3648 (N_3648,N_2423,In_4394);
nand U3649 (N_3649,N_2314,N_1921);
or U3650 (N_3650,N_1247,In_503);
or U3651 (N_3651,In_4828,N_2691);
and U3652 (N_3652,N_1649,N_1834);
or U3653 (N_3653,N_2931,In_3893);
nor U3654 (N_3654,N_906,N_815);
or U3655 (N_3655,N_2883,In_1237);
nand U3656 (N_3656,N_2656,In_1386);
nor U3657 (N_3657,In_211,In_4833);
xnor U3658 (N_3658,In_4626,N_2902);
and U3659 (N_3659,N_299,In_838);
xor U3660 (N_3660,N_2127,In_3297);
nor U3661 (N_3661,N_2115,N_1782);
and U3662 (N_3662,In_1105,In_2662);
or U3663 (N_3663,In_86,N_176);
nor U3664 (N_3664,N_2195,In_2619);
and U3665 (N_3665,N_2411,N_2575);
or U3666 (N_3666,N_2662,In_3693);
xnor U3667 (N_3667,N_2911,In_885);
nor U3668 (N_3668,In_1766,In_2345);
or U3669 (N_3669,N_2265,In_3705);
nand U3670 (N_3670,N_2602,N_2232);
xor U3671 (N_3671,N_2816,In_3952);
or U3672 (N_3672,N_2103,N_1965);
xor U3673 (N_3673,N_2020,N_1222);
xor U3674 (N_3674,N_2388,In_2296);
or U3675 (N_3675,N_2086,N_2492);
nand U3676 (N_3676,N_2923,In_4342);
or U3677 (N_3677,N_2772,In_1856);
xor U3678 (N_3678,N_2919,In_1212);
and U3679 (N_3679,In_2543,N_2192);
nor U3680 (N_3680,N_2446,In_3154);
nand U3681 (N_3681,N_2105,N_2862);
and U3682 (N_3682,N_2798,In_4972);
and U3683 (N_3683,In_68,N_279);
nand U3684 (N_3684,N_2003,In_1534);
and U3685 (N_3685,N_1239,In_2238);
or U3686 (N_3686,N_2047,N_2267);
xnor U3687 (N_3687,In_4047,N_2929);
or U3688 (N_3688,N_2891,In_3339);
and U3689 (N_3689,N_2594,N_87);
xor U3690 (N_3690,In_3642,In_296);
nand U3691 (N_3691,In_2420,N_2476);
nor U3692 (N_3692,N_2599,N_2156);
nand U3693 (N_3693,N_2354,In_2975);
and U3694 (N_3694,N_194,In_4483);
nand U3695 (N_3695,N_2473,In_5);
nand U3696 (N_3696,N_2215,N_2014);
and U3697 (N_3697,In_1580,N_2939);
nor U3698 (N_3698,N_2963,N_1647);
and U3699 (N_3699,N_2665,N_1372);
nand U3700 (N_3700,N_2478,N_1029);
and U3701 (N_3701,N_76,N_2767);
or U3702 (N_3702,In_2771,N_2775);
xnor U3703 (N_3703,N_2486,N_2546);
nor U3704 (N_3704,In_3134,N_1726);
and U3705 (N_3705,N_2274,In_3734);
and U3706 (N_3706,N_2632,N_2134);
nand U3707 (N_3707,N_2198,N_2143);
nor U3708 (N_3708,In_4324,In_2513);
xnor U3709 (N_3709,N_2799,N_2734);
nor U3710 (N_3710,N_519,In_3651);
nor U3711 (N_3711,N_2588,N_2256);
nor U3712 (N_3712,N_2392,In_2890);
xnor U3713 (N_3713,N_1817,In_483);
nand U3714 (N_3714,N_1081,N_2384);
xor U3715 (N_3715,N_1537,N_2258);
and U3716 (N_3716,In_526,N_374);
nor U3717 (N_3717,N_1664,In_1844);
xnor U3718 (N_3718,In_3010,In_1222);
nand U3719 (N_3719,N_2271,N_693);
or U3720 (N_3720,N_2545,N_2917);
nor U3721 (N_3721,N_2773,N_2514);
or U3722 (N_3722,N_2733,N_2515);
nor U3723 (N_3723,In_335,In_3532);
xor U3724 (N_3724,N_2857,N_2126);
nand U3725 (N_3725,N_38,N_2695);
and U3726 (N_3726,N_2094,N_2440);
nor U3727 (N_3727,In_2822,In_2925);
xor U3728 (N_3728,N_2246,N_1862);
and U3729 (N_3729,N_2049,N_1814);
and U3730 (N_3730,N_2938,N_2379);
nand U3731 (N_3731,N_2229,N_2208);
or U3732 (N_3732,N_1311,N_2752);
nand U3733 (N_3733,N_1362,N_2363);
xor U3734 (N_3734,N_2844,N_2600);
or U3735 (N_3735,In_4712,N_2593);
nand U3736 (N_3736,N_2873,In_3176);
and U3737 (N_3737,In_3020,N_2975);
or U3738 (N_3738,N_1238,N_2587);
xor U3739 (N_3739,N_1851,In_2753);
nor U3740 (N_3740,In_2004,N_2538);
or U3741 (N_3741,In_1861,N_2088);
nor U3742 (N_3742,In_1912,N_2331);
and U3743 (N_3743,N_2627,N_2062);
nor U3744 (N_3744,N_1395,N_2279);
xnor U3745 (N_3745,N_2777,In_4390);
and U3746 (N_3746,In_4832,N_2898);
nor U3747 (N_3747,N_292,N_646);
or U3748 (N_3748,N_1253,N_2301);
xnor U3749 (N_3749,N_2344,N_2146);
xor U3750 (N_3750,N_2319,N_637);
nor U3751 (N_3751,N_2826,N_1307);
or U3752 (N_3752,In_535,N_927);
nand U3753 (N_3753,N_2240,N_2779);
nor U3754 (N_3754,N_853,N_1175);
nor U3755 (N_3755,In_3067,N_889);
or U3756 (N_3756,N_610,In_39);
nor U3757 (N_3757,N_2140,N_186);
and U3758 (N_3758,N_1144,N_2445);
xnor U3759 (N_3759,N_2992,N_1010);
or U3760 (N_3760,In_830,N_2382);
or U3761 (N_3761,In_4936,N_2651);
nor U3762 (N_3762,N_2838,N_2112);
nand U3763 (N_3763,In_984,N_2516);
xnor U3764 (N_3764,N_1588,In_4428);
nand U3765 (N_3765,In_3787,In_2754);
xnor U3766 (N_3766,In_384,In_4007);
or U3767 (N_3767,In_454,N_2819);
or U3768 (N_3768,N_196,N_2245);
xor U3769 (N_3769,N_2081,N_609);
xor U3770 (N_3770,N_2306,N_1854);
and U3771 (N_3771,N_2666,In_4107);
nand U3772 (N_3772,N_804,In_4681);
xnor U3773 (N_3773,N_2647,In_4492);
and U3774 (N_3774,N_2092,N_2682);
nor U3775 (N_3775,N_992,N_2759);
or U3776 (N_3776,N_2719,N_2479);
nor U3777 (N_3777,In_999,N_2017);
xnor U3778 (N_3778,In_4038,N_1567);
and U3779 (N_3779,N_2965,N_2935);
nand U3780 (N_3780,In_2461,N_1404);
nor U3781 (N_3781,N_2255,In_753);
or U3782 (N_3782,In_3216,N_2748);
xor U3783 (N_3783,N_2372,N_1085);
nor U3784 (N_3784,N_2006,In_2871);
xnor U3785 (N_3785,N_2503,N_2703);
and U3786 (N_3786,N_2076,N_2953);
or U3787 (N_3787,N_2613,N_2561);
or U3788 (N_3788,In_2140,N_78);
and U3789 (N_3789,N_1730,N_2776);
or U3790 (N_3790,In_549,N_2571);
nor U3791 (N_3791,N_2204,N_669);
nor U3792 (N_3792,N_2100,N_1423);
nor U3793 (N_3793,N_2280,N_2688);
and U3794 (N_3794,In_4136,N_2558);
or U3795 (N_3795,In_41,N_2419);
or U3796 (N_3796,N_2283,N_1500);
nor U3797 (N_3797,N_1416,N_261);
or U3798 (N_3798,N_2410,N_1676);
nand U3799 (N_3799,N_2864,N_2442);
and U3800 (N_3800,N_2617,In_4693);
nor U3801 (N_3801,N_2770,N_2858);
and U3802 (N_3802,N_1279,N_1223);
xor U3803 (N_3803,N_631,N_2122);
nand U3804 (N_3804,In_398,N_2488);
and U3805 (N_3805,N_2837,N_2364);
xnor U3806 (N_3806,N_2349,In_4251);
xnor U3807 (N_3807,In_4734,N_1479);
nand U3808 (N_3808,In_4526,N_2141);
nand U3809 (N_3809,N_2671,N_2091);
nor U3810 (N_3810,In_2806,N_1531);
and U3811 (N_3811,In_471,In_3723);
nand U3812 (N_3812,N_2962,N_2737);
xor U3813 (N_3813,N_1073,N_1936);
nor U3814 (N_3814,N_2170,In_3332);
nand U3815 (N_3815,N_46,N_2941);
and U3816 (N_3816,In_374,N_2832);
xor U3817 (N_3817,N_1482,N_134);
nand U3818 (N_3818,N_2604,N_2239);
xnor U3819 (N_3819,N_2921,N_2640);
xnor U3820 (N_3820,In_52,N_2589);
and U3821 (N_3821,N_1516,N_778);
xor U3822 (N_3822,N_2334,N_2507);
and U3823 (N_3823,In_3193,N_53);
nand U3824 (N_3824,In_1814,N_2311);
xor U3825 (N_3825,N_1612,In_3794);
xnor U3826 (N_3826,In_1830,N_1969);
nand U3827 (N_3827,N_2646,N_2728);
nand U3828 (N_3828,N_2802,N_2660);
nand U3829 (N_3829,In_3468,N_2537);
xor U3830 (N_3830,N_2540,In_4930);
and U3831 (N_3831,N_145,In_3110);
xor U3832 (N_3832,N_1228,N_1940);
or U3833 (N_3833,N_2138,N_2487);
xor U3834 (N_3834,N_1264,N_2061);
or U3835 (N_3835,In_4546,In_3857);
xor U3836 (N_3836,N_2335,N_2291);
nor U3837 (N_3837,N_578,N_2416);
xnor U3838 (N_3838,In_4944,N_2550);
nand U3839 (N_3839,In_64,N_2793);
nor U3840 (N_3840,N_2801,N_2365);
nand U3841 (N_3841,N_2310,N_2358);
nor U3842 (N_3842,N_2783,In_4687);
and U3843 (N_3843,N_2548,N_2513);
or U3844 (N_3844,In_298,N_1841);
and U3845 (N_3845,N_2912,N_2435);
nand U3846 (N_3846,N_2747,N_1176);
and U3847 (N_3847,N_2560,N_2854);
xnor U3848 (N_3848,In_4174,N_2987);
and U3849 (N_3849,In_1803,In_1081);
and U3850 (N_3850,N_1733,N_2815);
nor U3851 (N_3851,N_1708,N_2527);
nor U3852 (N_3852,In_2097,In_354);
and U3853 (N_3853,In_4131,N_1798);
xor U3854 (N_3854,In_169,N_503);
xor U3855 (N_3855,N_2444,N_2761);
nand U3856 (N_3856,N_2160,N_404);
or U3857 (N_3857,N_138,N_2456);
nand U3858 (N_3858,N_2886,In_4615);
xor U3859 (N_3859,N_2079,N_1618);
and U3860 (N_3860,In_1655,In_3109);
and U3861 (N_3861,N_2825,N_1654);
nand U3862 (N_3862,N_2925,N_2504);
or U3863 (N_3863,In_2388,N_971);
nor U3864 (N_3864,N_2582,In_4191);
or U3865 (N_3865,N_1269,N_2080);
nand U3866 (N_3866,N_2383,N_1747);
nand U3867 (N_3867,N_2278,In_1751);
nor U3868 (N_3868,In_3016,In_567);
and U3869 (N_3869,In_3315,N_2895);
and U3870 (N_3870,N_2389,N_2601);
nand U3871 (N_3871,N_2197,In_3978);
xor U3872 (N_3872,N_1039,N_1042);
or U3873 (N_3873,N_2584,N_892);
nand U3874 (N_3874,N_1674,N_309);
nor U3875 (N_3875,N_2034,N_2464);
nor U3876 (N_3876,N_2451,N_2158);
nand U3877 (N_3877,N_958,N_2116);
xor U3878 (N_3878,N_2007,N_2018);
nor U3879 (N_3879,N_1009,N_2421);
nand U3880 (N_3880,N_1424,N_721);
nand U3881 (N_3881,N_1707,N_1302);
nand U3882 (N_3882,N_1392,In_4977);
nand U3883 (N_3883,In_2172,In_3722);
xor U3884 (N_3884,N_1044,N_2161);
nand U3885 (N_3885,N_2841,N_2717);
and U3886 (N_3886,In_643,N_1400);
nand U3887 (N_3887,N_2448,N_657);
or U3888 (N_3888,N_1263,N_1822);
nor U3889 (N_3889,In_4319,N_2856);
xnor U3890 (N_3890,In_4800,N_287);
xor U3891 (N_3891,N_2672,In_2663);
xor U3892 (N_3892,N_1465,N_2320);
xor U3893 (N_3893,In_4904,N_2818);
and U3894 (N_3894,N_948,N_2196);
xor U3895 (N_3895,N_2482,N_2008);
or U3896 (N_3896,N_2237,N_2011);
nand U3897 (N_3897,N_2352,In_3682);
nand U3898 (N_3898,N_2524,N_1973);
nor U3899 (N_3899,N_1435,N_2471);
and U3900 (N_3900,In_3408,N_1686);
xnor U3901 (N_3901,In_406,N_2029);
xnor U3902 (N_3902,In_4624,In_637);
nand U3903 (N_3903,N_2989,In_1421);
nor U3904 (N_3904,N_2381,N_643);
and U3905 (N_3905,N_312,N_2096);
xor U3906 (N_3906,N_2867,N_496);
or U3907 (N_3907,In_1384,In_3071);
and U3908 (N_3908,In_2080,In_419);
or U3909 (N_3909,N_2226,N_2402);
and U3910 (N_3910,N_2554,N_2329);
nor U3911 (N_3911,In_4129,N_2193);
nor U3912 (N_3912,N_1103,N_2303);
nand U3913 (N_3913,N_1617,In_715);
xnor U3914 (N_3914,N_2699,N_1728);
nand U3915 (N_3915,In_2404,N_2181);
nor U3916 (N_3916,N_2355,N_2366);
nand U3917 (N_3917,In_481,In_2072);
nor U3918 (N_3918,In_327,In_232);
nor U3919 (N_3919,N_2569,N_2013);
and U3920 (N_3920,In_733,N_2289);
or U3921 (N_3921,N_2202,N_1035);
or U3922 (N_3922,In_422,In_877);
xnor U3923 (N_3923,N_2432,N_2869);
and U3924 (N_3924,N_1653,N_2282);
xnor U3925 (N_3925,N_178,N_1031);
nand U3926 (N_3926,N_2768,N_2905);
or U3927 (N_3927,N_2732,In_2307);
and U3928 (N_3928,In_193,N_711);
xnor U3929 (N_3929,N_2426,N_2667);
xor U3930 (N_3930,N_2359,N_2031);
and U3931 (N_3931,N_2185,In_1573);
or U3932 (N_3932,N_2356,N_2848);
or U3933 (N_3933,In_1671,N_2151);
nand U3934 (N_3934,N_2983,N_2817);
nor U3935 (N_3935,N_2203,N_2104);
xnor U3936 (N_3936,N_2428,N_2970);
or U3937 (N_3937,N_2567,N_2889);
and U3938 (N_3938,N_2638,N_2679);
and U3939 (N_3939,In_442,In_1161);
nand U3940 (N_3940,N_1917,N_1806);
or U3941 (N_3941,N_2843,In_1387);
and U3942 (N_3942,N_2763,In_3610);
or U3943 (N_3943,In_1225,N_2174);
and U3944 (N_3944,N_2454,In_2517);
xor U3945 (N_3945,N_2804,N_301);
and U3946 (N_3946,N_2409,N_2437);
and U3947 (N_3947,N_1458,N_826);
nor U3948 (N_3948,In_3145,In_4530);
or U3949 (N_3949,In_918,N_2966);
nor U3950 (N_3950,In_112,N_2901);
xnor U3951 (N_3951,N_2505,In_4744);
or U3952 (N_3952,N_2659,In_3480);
xnor U3953 (N_3953,N_1711,N_2285);
or U3954 (N_3954,N_2223,N_1698);
nor U3955 (N_3955,N_2628,N_1595);
xnor U3956 (N_3956,N_1189,N_1928);
xor U3957 (N_3957,N_2408,N_1572);
nand U3958 (N_3958,In_3114,N_2566);
xor U3959 (N_3959,N_2784,In_2329);
xnor U3960 (N_3960,N_396,In_2683);
xnor U3961 (N_3961,In_2615,In_3215);
and U3962 (N_3962,N_2674,N_2398);
xor U3963 (N_3963,N_1620,N_2262);
and U3964 (N_3964,N_2872,In_2914);
nor U3965 (N_3965,In_303,N_2521);
or U3966 (N_3966,N_2078,N_2395);
and U3967 (N_3967,N_2491,N_1053);
xor U3968 (N_3968,N_2190,N_1976);
nor U3969 (N_3969,N_1471,N_1599);
nand U3970 (N_3970,N_306,In_2621);
or U3971 (N_3971,N_2021,N_2853);
and U3972 (N_3972,N_1141,N_2821);
nand U3973 (N_3973,N_1383,In_3164);
nand U3974 (N_3974,N_2786,N_2525);
or U3975 (N_3975,In_1226,In_491);
nand U3976 (N_3976,N_28,N_2641);
or U3977 (N_3977,N_2781,N_2154);
nand U3978 (N_3978,In_4608,N_2083);
or U3979 (N_3979,N_2764,N_2387);
xor U3980 (N_3980,N_42,N_2906);
or U3981 (N_3981,In_635,In_3414);
or U3982 (N_3982,N_2708,N_121);
or U3983 (N_3983,N_2489,N_52);
nor U3984 (N_3984,N_1875,N_2217);
nor U3985 (N_3985,N_2592,N_2726);
or U3986 (N_3986,N_2758,N_1589);
xnor U3987 (N_3987,N_1037,N_2483);
and U3988 (N_3988,N_2281,N_2611);
or U3989 (N_3989,N_2543,N_2878);
and U3990 (N_3990,N_2266,N_2394);
and U3991 (N_3991,In_1279,N_2981);
or U3992 (N_3992,N_2295,N_2960);
xnor U3993 (N_3993,N_1540,In_1622);
nand U3994 (N_3994,N_1145,N_1784);
or U3995 (N_3995,N_2623,N_2714);
and U3996 (N_3996,N_2675,N_919);
nand U3997 (N_3997,N_2276,In_1101);
nor U3998 (N_3998,N_2685,N_2789);
xnor U3999 (N_3999,In_1097,N_2222);
or U4000 (N_4000,N_3873,N_3320);
or U4001 (N_4001,N_3954,N_3761);
and U4002 (N_4002,N_3720,N_3200);
and U4003 (N_4003,N_3318,N_3924);
nand U4004 (N_4004,N_3806,N_3565);
nand U4005 (N_4005,N_3405,N_3251);
nor U4006 (N_4006,N_3957,N_3827);
and U4007 (N_4007,N_3271,N_3169);
xor U4008 (N_4008,N_3771,N_3083);
nand U4009 (N_4009,N_3423,N_3338);
and U4010 (N_4010,N_3865,N_3333);
nor U4011 (N_4011,N_3201,N_3196);
nor U4012 (N_4012,N_3014,N_3539);
or U4013 (N_4013,N_3136,N_3586);
nor U4014 (N_4014,N_3164,N_3383);
and U4015 (N_4015,N_3833,N_3507);
and U4016 (N_4016,N_3934,N_3882);
or U4017 (N_4017,N_3455,N_3080);
xnor U4018 (N_4018,N_3341,N_3813);
xor U4019 (N_4019,N_3149,N_3579);
nand U4020 (N_4020,N_3388,N_3207);
nand U4021 (N_4021,N_3028,N_3452);
and U4022 (N_4022,N_3242,N_3863);
nand U4023 (N_4023,N_3424,N_3979);
nand U4024 (N_4024,N_3160,N_3199);
xnor U4025 (N_4025,N_3835,N_3591);
nand U4026 (N_4026,N_3244,N_3727);
or U4027 (N_4027,N_3343,N_3741);
nand U4028 (N_4028,N_3130,N_3962);
nor U4029 (N_4029,N_3257,N_3362);
nand U4030 (N_4030,N_3682,N_3183);
and U4031 (N_4031,N_3548,N_3558);
nand U4032 (N_4032,N_3409,N_3768);
xnor U4033 (N_4033,N_3802,N_3787);
and U4034 (N_4034,N_3402,N_3735);
and U4035 (N_4035,N_3459,N_3557);
xor U4036 (N_4036,N_3050,N_3303);
nand U4037 (N_4037,N_3439,N_3473);
nor U4038 (N_4038,N_3992,N_3792);
xor U4039 (N_4039,N_3945,N_3245);
and U4040 (N_4040,N_3931,N_3477);
nor U4041 (N_4041,N_3564,N_3796);
nor U4042 (N_4042,N_3808,N_3901);
and U4043 (N_4043,N_3815,N_3948);
nor U4044 (N_4044,N_3941,N_3017);
nand U4045 (N_4045,N_3392,N_3536);
and U4046 (N_4046,N_3418,N_3858);
and U4047 (N_4047,N_3914,N_3620);
nand U4048 (N_4048,N_3104,N_3893);
or U4049 (N_4049,N_3029,N_3943);
nor U4050 (N_4050,N_3851,N_3230);
xor U4051 (N_4051,N_3165,N_3542);
or U4052 (N_4052,N_3268,N_3818);
nor U4053 (N_4053,N_3875,N_3346);
and U4054 (N_4054,N_3414,N_3575);
nand U4055 (N_4055,N_3492,N_3112);
nand U4056 (N_4056,N_3661,N_3755);
and U4057 (N_4057,N_3728,N_3133);
nand U4058 (N_4058,N_3148,N_3400);
nor U4059 (N_4059,N_3144,N_3457);
nor U4060 (N_4060,N_3264,N_3217);
nand U4061 (N_4061,N_3537,N_3973);
nand U4062 (N_4062,N_3184,N_3099);
nand U4063 (N_4063,N_3950,N_3631);
and U4064 (N_4064,N_3098,N_3785);
and U4065 (N_4065,N_3895,N_3134);
or U4066 (N_4066,N_3347,N_3265);
or U4067 (N_4067,N_3150,N_3514);
or U4068 (N_4068,N_3977,N_3438);
or U4069 (N_4069,N_3036,N_3225);
xnor U4070 (N_4070,N_3772,N_3316);
or U4071 (N_4071,N_3000,N_3676);
or U4072 (N_4072,N_3672,N_3479);
or U4073 (N_4073,N_3113,N_3571);
nor U4074 (N_4074,N_3351,N_3469);
xor U4075 (N_4075,N_3399,N_3730);
nand U4076 (N_4076,N_3842,N_3488);
xor U4077 (N_4077,N_3413,N_3512);
or U4078 (N_4078,N_3489,N_3419);
nand U4079 (N_4079,N_3317,N_3804);
or U4080 (N_4080,N_3870,N_3995);
nand U4081 (N_4081,N_3773,N_3018);
nor U4082 (N_4082,N_3355,N_3644);
and U4083 (N_4083,N_3953,N_3421);
nor U4084 (N_4084,N_3529,N_3092);
nand U4085 (N_4085,N_3241,N_3763);
and U4086 (N_4086,N_3697,N_3908);
and U4087 (N_4087,N_3657,N_3938);
nand U4088 (N_4088,N_3607,N_3709);
or U4089 (N_4089,N_3410,N_3064);
xor U4090 (N_4090,N_3856,N_3269);
nand U4091 (N_4091,N_3501,N_3004);
or U4092 (N_4092,N_3968,N_3260);
xnor U4093 (N_4093,N_3430,N_3609);
nor U4094 (N_4094,N_3190,N_3061);
or U4095 (N_4095,N_3103,N_3838);
nor U4096 (N_4096,N_3091,N_3449);
or U4097 (N_4097,N_3508,N_3721);
xor U4098 (N_4098,N_3222,N_3472);
and U4099 (N_4099,N_3101,N_3600);
or U4100 (N_4100,N_3956,N_3031);
or U4101 (N_4101,N_3033,N_3695);
nand U4102 (N_4102,N_3541,N_3708);
nor U4103 (N_4103,N_3275,N_3246);
nor U4104 (N_4104,N_3340,N_3593);
xnor U4105 (N_4105,N_3832,N_3700);
xor U4106 (N_4106,N_3589,N_3191);
xor U4107 (N_4107,N_3871,N_3853);
nor U4108 (N_4108,N_3496,N_3044);
and U4109 (N_4109,N_3262,N_3187);
or U4110 (N_4110,N_3606,N_3356);
or U4111 (N_4111,N_3864,N_3329);
and U4112 (N_4112,N_3497,N_3118);
or U4113 (N_4113,N_3876,N_3583);
and U4114 (N_4114,N_3905,N_3243);
or U4115 (N_4115,N_3443,N_3693);
xnor U4116 (N_4116,N_3256,N_3060);
xnor U4117 (N_4117,N_3855,N_3843);
and U4118 (N_4118,N_3012,N_3553);
nor U4119 (N_4119,N_3247,N_3587);
xor U4120 (N_4120,N_3203,N_3624);
nand U4121 (N_4121,N_3498,N_3633);
or U4122 (N_4122,N_3040,N_3667);
nand U4123 (N_4123,N_3255,N_3002);
and U4124 (N_4124,N_3051,N_3839);
nand U4125 (N_4125,N_3974,N_3016);
nand U4126 (N_4126,N_3563,N_3745);
nor U4127 (N_4127,N_3286,N_3887);
nand U4128 (N_4128,N_3592,N_3010);
nand U4129 (N_4129,N_3683,N_3528);
xor U4130 (N_4130,N_3770,N_3555);
and U4131 (N_4131,N_3543,N_3868);
nor U4132 (N_4132,N_3698,N_3546);
nor U4133 (N_4133,N_3482,N_3471);
and U4134 (N_4134,N_3862,N_3898);
nor U4135 (N_4135,N_3344,N_3518);
or U4136 (N_4136,N_3048,N_3218);
nand U4137 (N_4137,N_3909,N_3441);
or U4138 (N_4138,N_3325,N_3252);
nand U4139 (N_4139,N_3635,N_3155);
or U4140 (N_4140,N_3567,N_3213);
or U4141 (N_4141,N_3967,N_3240);
xor U4142 (N_4142,N_3677,N_3921);
nand U4143 (N_4143,N_3825,N_3699);
and U4144 (N_4144,N_3976,N_3090);
nand U4145 (N_4145,N_3550,N_3717);
or U4146 (N_4146,N_3110,N_3214);
or U4147 (N_4147,N_3581,N_3470);
nand U4148 (N_4148,N_3647,N_3532);
nor U4149 (N_4149,N_3319,N_3052);
xor U4150 (N_4150,N_3603,N_3666);
nor U4151 (N_4151,N_3637,N_3391);
or U4152 (N_4152,N_3045,N_3448);
or U4153 (N_4153,N_3896,N_3357);
or U4154 (N_4154,N_3041,N_3490);
nand U4155 (N_4155,N_3664,N_3076);
xnor U4156 (N_4156,N_3178,N_3776);
or U4157 (N_4157,N_3930,N_3739);
or U4158 (N_4158,N_3601,N_3042);
xnor U4159 (N_4159,N_3233,N_3248);
nor U4160 (N_4160,N_3481,N_3163);
nor U4161 (N_4161,N_3561,N_3812);
nand U4162 (N_4162,N_3353,N_3504);
and U4163 (N_4163,N_3142,N_3364);
and U4164 (N_4164,N_3179,N_3929);
or U4165 (N_4165,N_3038,N_3936);
or U4166 (N_4166,N_3878,N_3662);
nor U4167 (N_4167,N_3335,N_3463);
or U4168 (N_4168,N_3309,N_3749);
nand U4169 (N_4169,N_3132,N_3650);
xor U4170 (N_4170,N_3324,N_3066);
nor U4171 (N_4171,N_3281,N_3922);
and U4172 (N_4172,N_3226,N_3328);
nand U4173 (N_4173,N_3849,N_3544);
nor U4174 (N_4174,N_3003,N_3350);
nand U4175 (N_4175,N_3942,N_3928);
nor U4176 (N_4176,N_3267,N_3978);
nand U4177 (N_4177,N_3432,N_3961);
or U4178 (N_4178,N_3517,N_3069);
nand U4179 (N_4179,N_3008,N_3440);
xor U4180 (N_4180,N_3605,N_3170);
xor U4181 (N_4181,N_3752,N_3074);
nor U4182 (N_4182,N_3902,N_3520);
nand U4183 (N_4183,N_3454,N_3015);
xor U4184 (N_4184,N_3964,N_3814);
nor U4185 (N_4185,N_3846,N_3850);
nor U4186 (N_4186,N_3651,N_3366);
nor U4187 (N_4187,N_3085,N_3078);
nor U4188 (N_4188,N_3416,N_3623);
nand U4189 (N_4189,N_3991,N_3108);
nor U4190 (N_4190,N_3249,N_3969);
xor U4191 (N_4191,N_3519,N_3460);
and U4192 (N_4192,N_3228,N_3331);
xor U4193 (N_4193,N_3368,N_3186);
nand U4194 (N_4194,N_3088,N_3604);
nor U4195 (N_4195,N_3559,N_3983);
nor U4196 (N_4196,N_3830,N_3824);
nor U4197 (N_4197,N_3927,N_3554);
nand U4198 (N_4198,N_3743,N_3782);
xnor U4199 (N_4199,N_3704,N_3598);
and U4200 (N_4200,N_3861,N_3574);
nand U4201 (N_4201,N_3445,N_3465);
xor U4202 (N_4202,N_3822,N_3919);
and U4203 (N_4203,N_3713,N_3464);
or U4204 (N_4204,N_3900,N_3602);
xnor U4205 (N_4205,N_3885,N_3874);
nand U4206 (N_4206,N_3075,N_3759);
nand U4207 (N_4207,N_3612,N_3263);
xnor U4208 (N_4208,N_3451,N_3588);
nor U4209 (N_4209,N_3916,N_3363);
nand U4210 (N_4210,N_3070,N_3767);
nand U4211 (N_4211,N_3655,N_3114);
or U4212 (N_4212,N_3288,N_3807);
or U4213 (N_4213,N_3147,N_3336);
or U4214 (N_4214,N_3208,N_3857);
and U4215 (N_4215,N_3859,N_3348);
nand U4216 (N_4216,N_3775,N_3387);
nor U4217 (N_4217,N_3216,N_3616);
or U4218 (N_4218,N_3643,N_3381);
and U4219 (N_4219,N_3705,N_3877);
xnor U4220 (N_4220,N_3834,N_3793);
nor U4221 (N_4221,N_3596,N_3046);
and U4222 (N_4222,N_3852,N_3167);
or U4223 (N_4223,N_3461,N_3724);
nor U4224 (N_4224,N_3174,N_3625);
nand U4225 (N_4225,N_3744,N_3556);
xnor U4226 (N_4226,N_3946,N_3176);
nand U4227 (N_4227,N_3669,N_3784);
nand U4228 (N_4228,N_3327,N_3285);
xor U4229 (N_4229,N_3182,N_3786);
or U4230 (N_4230,N_3533,N_3011);
nor U4231 (N_4231,N_3385,N_3030);
or U4232 (N_4232,N_3013,N_3611);
nor U4233 (N_4233,N_3585,N_3466);
nand U4234 (N_4234,N_3933,N_3997);
nor U4235 (N_4235,N_3043,N_3282);
nor U4236 (N_4236,N_3671,N_3342);
and U4237 (N_4237,N_3433,N_3619);
or U4238 (N_4238,N_3648,N_3232);
nor U4239 (N_4239,N_3982,N_3211);
or U4240 (N_4240,N_3996,N_3975);
xnor U4241 (N_4241,N_3935,N_3159);
nor U4242 (N_4242,N_3685,N_3831);
and U4243 (N_4243,N_3753,N_3738);
and U4244 (N_4244,N_3370,N_3175);
or U4245 (N_4245,N_3143,N_3937);
and U4246 (N_4246,N_3458,N_3836);
or U4247 (N_4247,N_3172,N_3373);
or U4248 (N_4248,N_3157,N_3715);
xor U4249 (N_4249,N_3736,N_3963);
nor U4250 (N_4250,N_3406,N_3054);
xnor U4251 (N_4251,N_3122,N_3613);
or U4252 (N_4252,N_3139,N_3361);
xnor U4253 (N_4253,N_3379,N_3848);
xor U4254 (N_4254,N_3057,N_3748);
and U4255 (N_4255,N_3737,N_3800);
or U4256 (N_4256,N_3049,N_3516);
xnor U4257 (N_4257,N_3840,N_3560);
xnor U4258 (N_4258,N_3845,N_3189);
xor U4259 (N_4259,N_3980,N_3766);
nand U4260 (N_4260,N_3523,N_3302);
nor U4261 (N_4261,N_3193,N_3121);
nand U4262 (N_4262,N_3681,N_3531);
xor U4263 (N_4263,N_3540,N_3869);
or U4264 (N_4264,N_3298,N_3632);
xnor U4265 (N_4265,N_3126,N_3535);
and U4266 (N_4266,N_3883,N_3073);
and U4267 (N_4267,N_3272,N_3062);
or U4268 (N_4268,N_3679,N_3315);
nor U4269 (N_4269,N_3958,N_3740);
and U4270 (N_4270,N_3277,N_3146);
xor U4271 (N_4271,N_3910,N_3393);
xor U4272 (N_4272,N_3733,N_3360);
xor U4273 (N_4273,N_3947,N_3462);
nand U4274 (N_4274,N_3426,N_3289);
nand U4275 (N_4275,N_3981,N_3774);
nand U4276 (N_4276,N_3293,N_3694);
nand U4277 (N_4277,N_3788,N_3622);
nand U4278 (N_4278,N_3867,N_3483);
and U4279 (N_4279,N_3795,N_3854);
xnor U4280 (N_4280,N_3890,N_3597);
xor U4281 (N_4281,N_3194,N_3790);
nor U4282 (N_4282,N_3422,N_3939);
and U4283 (N_4283,N_3570,N_3545);
and U4284 (N_4284,N_3866,N_3135);
nor U4285 (N_4285,N_3680,N_3161);
nor U4286 (N_4286,N_3390,N_3227);
or U4287 (N_4287,N_3129,N_3499);
xnor U4288 (N_4288,N_3791,N_3109);
and U4289 (N_4289,N_3732,N_3659);
and U4290 (N_4290,N_3911,N_3221);
nand U4291 (N_4291,N_3436,N_3906);
nor U4292 (N_4292,N_3656,N_3986);
xor U4293 (N_4293,N_3847,N_3128);
and U4294 (N_4294,N_3310,N_3084);
or U4295 (N_4295,N_3365,N_3140);
and U4296 (N_4296,N_3783,N_3494);
nor U4297 (N_4297,N_3236,N_3754);
xor U4298 (N_4298,N_3641,N_3480);
and U4299 (N_4299,N_3258,N_3313);
and U4300 (N_4300,N_3089,N_3913);
nor U4301 (N_4301,N_3626,N_3229);
and U4302 (N_4302,N_3395,N_3478);
nand U4303 (N_4303,N_3185,N_3123);
nor U4304 (N_4304,N_3668,N_3491);
nor U4305 (N_4305,N_3442,N_3500);
and U4306 (N_4306,N_3897,N_3826);
xor U4307 (N_4307,N_3634,N_3311);
nor U4308 (N_4308,N_3396,N_3629);
and U4309 (N_4309,N_3025,N_3971);
or U4310 (N_4310,N_3181,N_3095);
nor U4311 (N_4311,N_3339,N_3125);
nand U4312 (N_4312,N_3446,N_3718);
or U4313 (N_4313,N_3714,N_3166);
xnor U4314 (N_4314,N_3117,N_3580);
nand U4315 (N_4315,N_3742,N_3547);
or U4316 (N_4316,N_3690,N_3837);
xor U4317 (N_4317,N_3777,N_3065);
and U4318 (N_4318,N_3872,N_3819);
or U4319 (N_4319,N_3284,N_3367);
or U4320 (N_4320,N_3841,N_3408);
xor U4321 (N_4321,N_3431,N_3314);
and U4322 (N_4322,N_3879,N_3590);
nand U4323 (N_4323,N_3502,N_3495);
nor U4324 (N_4324,N_3059,N_3710);
nand U4325 (N_4325,N_3920,N_3907);
or U4326 (N_4326,N_3349,N_3999);
nand U4327 (N_4327,N_3551,N_3035);
nor U4328 (N_4328,N_3158,N_3530);
nand U4329 (N_4329,N_3569,N_3485);
and U4330 (N_4330,N_3296,N_3308);
nor U4331 (N_4331,N_3456,N_3234);
nand U4332 (N_4332,N_3573,N_3223);
xor U4333 (N_4333,N_3747,N_3484);
and U4334 (N_4334,N_3618,N_3527);
and U4335 (N_4335,N_3617,N_3746);
nor U4336 (N_4336,N_3645,N_3034);
or U4337 (N_4337,N_3047,N_3153);
and U4338 (N_4338,N_3127,N_3096);
nand U4339 (N_4339,N_3111,N_3382);
nand U4340 (N_4340,N_3888,N_3468);
xnor U4341 (N_4341,N_3312,N_3063);
or U4342 (N_4342,N_3120,N_3703);
nor U4343 (N_4343,N_3654,N_3417);
and U4344 (N_4344,N_3972,N_3131);
or U4345 (N_4345,N_3412,N_3779);
nor U4346 (N_4346,N_3630,N_3007);
nand U4347 (N_4347,N_3572,N_3270);
nor U4348 (N_4348,N_3224,N_3917);
or U4349 (N_4349,N_3307,N_3881);
and U4350 (N_4350,N_3760,N_3621);
xor U4351 (N_4351,N_3696,N_3102);
nand U4352 (N_4352,N_3026,N_3889);
xor U4353 (N_4353,N_3162,N_3549);
nand U4354 (N_4354,N_3425,N_3354);
and U4355 (N_4355,N_3107,N_3798);
xor U4356 (N_4356,N_3926,N_3337);
nor U4357 (N_4357,N_3274,N_3156);
and U4358 (N_4358,N_3231,N_3640);
and U4359 (N_4359,N_3273,N_3506);
nand U4360 (N_4360,N_3912,N_3678);
nor U4361 (N_4361,N_3493,N_3509);
xnor U4362 (N_4362,N_3151,N_3297);
nand U4363 (N_4363,N_3524,N_3723);
nand U4364 (N_4364,N_3610,N_3447);
or U4365 (N_4365,N_3805,N_3577);
nor U4366 (N_4366,N_3940,N_3809);
nor U4367 (N_4367,N_3521,N_3023);
or U4368 (N_4368,N_3949,N_3254);
or U4369 (N_4369,N_3923,N_3615);
nor U4370 (N_4370,N_3077,N_3797);
xnor U4371 (N_4371,N_3079,N_3892);
or U4372 (N_4372,N_3769,N_3925);
and U4373 (N_4373,N_3434,N_3386);
nor U4374 (N_4374,N_3053,N_3145);
and U4375 (N_4375,N_3780,N_3067);
nor U4376 (N_4376,N_3538,N_3323);
nand U4377 (N_4377,N_3322,N_3687);
nand U4378 (N_4378,N_3420,N_3238);
and U4379 (N_4379,N_3614,N_3511);
nand U4380 (N_4380,N_3951,N_3032);
and U4381 (N_4381,N_3762,N_3087);
nor U4382 (N_4382,N_3966,N_3970);
or U4383 (N_4383,N_3398,N_3628);
xnor U4384 (N_4384,N_3450,N_3811);
nor U4385 (N_4385,N_3276,N_3932);
nand U4386 (N_4386,N_3301,N_3429);
and U4387 (N_4387,N_3692,N_3294);
xnor U4388 (N_4388,N_3192,N_3944);
nand U4389 (N_4389,N_3904,N_3056);
and U4390 (N_4390,N_3397,N_3177);
or U4391 (N_4391,N_3653,N_3326);
nor U4392 (N_4392,N_3844,N_3299);
nor U4393 (N_4393,N_3476,N_3106);
nor U4394 (N_4394,N_3415,N_3638);
nor U4395 (N_4395,N_3568,N_3860);
nand U4396 (N_4396,N_3712,N_3220);
xnor U4397 (N_4397,N_3829,N_3401);
xor U4398 (N_4398,N_3205,N_3195);
nand U4399 (N_4399,N_3994,N_3778);
nand U4400 (N_4400,N_3345,N_3670);
nor U4401 (N_4401,N_3562,N_3376);
nand U4402 (N_4402,N_3998,N_3304);
nand U4403 (N_4403,N_3375,N_3515);
and U4404 (N_4404,N_3380,N_3823);
or U4405 (N_4405,N_3321,N_3171);
nand U4406 (N_4406,N_3428,N_3435);
xor U4407 (N_4407,N_3334,N_3891);
nor U4408 (N_4408,N_3006,N_3055);
xor U4409 (N_4409,N_3801,N_3250);
or U4410 (N_4410,N_3377,N_3691);
or U4411 (N_4411,N_3686,N_3305);
and U4412 (N_4412,N_3358,N_3283);
or U4413 (N_4413,N_3803,N_3253);
xor U4414 (N_4414,N_3206,N_3711);
or U4415 (N_4415,N_3407,N_3820);
nor U4416 (N_4416,N_3526,N_3487);
or U4417 (N_4417,N_3209,N_3594);
and U4418 (N_4418,N_3475,N_3756);
and U4419 (N_4419,N_3627,N_3235);
nand U4420 (N_4420,N_3750,N_3115);
nor U4421 (N_4421,N_3734,N_3198);
or U4422 (N_4422,N_3534,N_3100);
nor U4423 (N_4423,N_3291,N_3959);
and U4424 (N_4424,N_3810,N_3684);
nand U4425 (N_4425,N_3210,N_3828);
and U4426 (N_4426,N_3082,N_3019);
nand U4427 (N_4427,N_3673,N_3037);
nand U4428 (N_4428,N_3688,N_3068);
or U4429 (N_4429,N_3378,N_3582);
nand U4430 (N_4430,N_3503,N_3212);
and U4431 (N_4431,N_3453,N_3566);
nor U4432 (N_4432,N_3188,N_3279);
and U4433 (N_4433,N_3394,N_3886);
nor U4434 (N_4434,N_3990,N_3706);
xor U4435 (N_4435,N_3725,N_3903);
and U4436 (N_4436,N_3595,N_3689);
nand U4437 (N_4437,N_3764,N_3384);
xnor U4438 (N_4438,N_3278,N_3952);
nor U4439 (N_4439,N_3141,N_3280);
xnor U4440 (N_4440,N_3215,N_3093);
nor U4441 (N_4441,N_3636,N_3024);
or U4442 (N_4442,N_3332,N_3474);
or U4443 (N_4443,N_3204,N_3352);
nand U4444 (N_4444,N_3290,N_3985);
nor U4445 (N_4445,N_3799,N_3988);
and U4446 (N_4446,N_3894,N_3137);
nand U4447 (N_4447,N_3510,N_3525);
or U4448 (N_4448,N_3072,N_3022);
nand U4449 (N_4449,N_3821,N_3915);
nand U4450 (N_4450,N_3197,N_3124);
and U4451 (N_4451,N_3639,N_3599);
xnor U4452 (N_4452,N_3467,N_3306);
nor U4453 (N_4453,N_3020,N_3330);
nor U4454 (N_4454,N_3021,N_3719);
and U4455 (N_4455,N_3918,N_3965);
nand U4456 (N_4456,N_3369,N_3663);
xnor U4457 (N_4457,N_3675,N_3731);
and U4458 (N_4458,N_3437,N_3094);
nor U4459 (N_4459,N_3295,N_3608);
nand U4460 (N_4460,N_3513,N_3729);
or U4461 (N_4461,N_3987,N_3758);
nand U4462 (N_4462,N_3665,N_3001);
and U4463 (N_4463,N_3300,N_3702);
nand U4464 (N_4464,N_3154,N_3984);
nand U4465 (N_4465,N_3584,N_3292);
and U4466 (N_4466,N_3168,N_3427);
nand U4467 (N_4467,N_3522,N_3751);
nand U4468 (N_4468,N_3505,N_3955);
xnor U4469 (N_4469,N_3649,N_3701);
xor U4470 (N_4470,N_3005,N_3173);
nand U4471 (N_4471,N_3757,N_3794);
and U4472 (N_4472,N_3726,N_3411);
xnor U4473 (N_4473,N_3372,N_3081);
nand U4474 (N_4474,N_3359,N_3105);
xnor U4475 (N_4475,N_3097,N_3707);
nor U4476 (N_4476,N_3646,N_3552);
nand U4477 (N_4477,N_3993,N_3652);
and U4478 (N_4478,N_3219,N_3444);
and U4479 (N_4479,N_3660,N_3899);
xnor U4480 (N_4480,N_3781,N_3989);
xnor U4481 (N_4481,N_3071,N_3119);
xor U4482 (N_4482,N_3817,N_3816);
xor U4483 (N_4483,N_3266,N_3039);
nor U4484 (N_4484,N_3058,N_3138);
or U4485 (N_4485,N_3086,N_3371);
xnor U4486 (N_4486,N_3259,N_3403);
nor U4487 (N_4487,N_3116,N_3180);
xor U4488 (N_4488,N_3374,N_3576);
xor U4489 (N_4489,N_3009,N_3237);
nor U4490 (N_4490,N_3486,N_3765);
nand U4491 (N_4491,N_3960,N_3239);
and U4492 (N_4492,N_3389,N_3202);
and U4493 (N_4493,N_3027,N_3880);
nor U4494 (N_4494,N_3261,N_3789);
or U4495 (N_4495,N_3404,N_3716);
and U4496 (N_4496,N_3884,N_3642);
nor U4497 (N_4497,N_3287,N_3722);
xnor U4498 (N_4498,N_3658,N_3674);
nor U4499 (N_4499,N_3578,N_3152);
nand U4500 (N_4500,N_3738,N_3125);
nor U4501 (N_4501,N_3340,N_3252);
and U4502 (N_4502,N_3230,N_3675);
or U4503 (N_4503,N_3921,N_3339);
and U4504 (N_4504,N_3804,N_3501);
and U4505 (N_4505,N_3023,N_3860);
xnor U4506 (N_4506,N_3590,N_3600);
nor U4507 (N_4507,N_3979,N_3810);
xor U4508 (N_4508,N_3405,N_3165);
xor U4509 (N_4509,N_3687,N_3149);
or U4510 (N_4510,N_3478,N_3793);
or U4511 (N_4511,N_3410,N_3919);
and U4512 (N_4512,N_3876,N_3948);
or U4513 (N_4513,N_3373,N_3847);
and U4514 (N_4514,N_3295,N_3582);
or U4515 (N_4515,N_3686,N_3610);
nand U4516 (N_4516,N_3940,N_3643);
nand U4517 (N_4517,N_3383,N_3311);
and U4518 (N_4518,N_3080,N_3602);
nand U4519 (N_4519,N_3231,N_3912);
or U4520 (N_4520,N_3518,N_3555);
nor U4521 (N_4521,N_3529,N_3523);
xor U4522 (N_4522,N_3542,N_3540);
nand U4523 (N_4523,N_3658,N_3314);
and U4524 (N_4524,N_3952,N_3640);
and U4525 (N_4525,N_3304,N_3006);
or U4526 (N_4526,N_3952,N_3767);
nor U4527 (N_4527,N_3217,N_3090);
xor U4528 (N_4528,N_3499,N_3111);
and U4529 (N_4529,N_3418,N_3296);
or U4530 (N_4530,N_3867,N_3418);
nand U4531 (N_4531,N_3588,N_3993);
nand U4532 (N_4532,N_3904,N_3736);
nand U4533 (N_4533,N_3205,N_3061);
and U4534 (N_4534,N_3661,N_3890);
nor U4535 (N_4535,N_3989,N_3685);
nand U4536 (N_4536,N_3951,N_3977);
xor U4537 (N_4537,N_3679,N_3864);
xor U4538 (N_4538,N_3312,N_3569);
or U4539 (N_4539,N_3004,N_3615);
xor U4540 (N_4540,N_3568,N_3074);
nor U4541 (N_4541,N_3674,N_3525);
and U4542 (N_4542,N_3028,N_3432);
nand U4543 (N_4543,N_3965,N_3439);
nand U4544 (N_4544,N_3971,N_3918);
nand U4545 (N_4545,N_3890,N_3161);
and U4546 (N_4546,N_3967,N_3650);
and U4547 (N_4547,N_3726,N_3186);
nor U4548 (N_4548,N_3281,N_3971);
xnor U4549 (N_4549,N_3884,N_3945);
nand U4550 (N_4550,N_3417,N_3628);
and U4551 (N_4551,N_3329,N_3441);
xor U4552 (N_4552,N_3986,N_3607);
or U4553 (N_4553,N_3874,N_3138);
or U4554 (N_4554,N_3096,N_3026);
xor U4555 (N_4555,N_3808,N_3650);
or U4556 (N_4556,N_3149,N_3613);
xor U4557 (N_4557,N_3278,N_3442);
nor U4558 (N_4558,N_3611,N_3597);
and U4559 (N_4559,N_3056,N_3846);
nand U4560 (N_4560,N_3532,N_3979);
or U4561 (N_4561,N_3946,N_3939);
xor U4562 (N_4562,N_3307,N_3917);
nand U4563 (N_4563,N_3324,N_3789);
nor U4564 (N_4564,N_3505,N_3737);
and U4565 (N_4565,N_3858,N_3594);
nand U4566 (N_4566,N_3587,N_3165);
or U4567 (N_4567,N_3251,N_3655);
nor U4568 (N_4568,N_3189,N_3805);
nor U4569 (N_4569,N_3659,N_3404);
nand U4570 (N_4570,N_3983,N_3110);
nor U4571 (N_4571,N_3991,N_3221);
xnor U4572 (N_4572,N_3905,N_3325);
nor U4573 (N_4573,N_3861,N_3970);
nand U4574 (N_4574,N_3234,N_3397);
xnor U4575 (N_4575,N_3837,N_3807);
nand U4576 (N_4576,N_3712,N_3709);
or U4577 (N_4577,N_3226,N_3495);
nand U4578 (N_4578,N_3670,N_3744);
xor U4579 (N_4579,N_3645,N_3150);
nand U4580 (N_4580,N_3911,N_3528);
nor U4581 (N_4581,N_3721,N_3452);
and U4582 (N_4582,N_3633,N_3786);
xnor U4583 (N_4583,N_3307,N_3632);
or U4584 (N_4584,N_3723,N_3741);
nor U4585 (N_4585,N_3093,N_3686);
nand U4586 (N_4586,N_3932,N_3902);
or U4587 (N_4587,N_3968,N_3151);
xor U4588 (N_4588,N_3078,N_3512);
nand U4589 (N_4589,N_3879,N_3753);
nand U4590 (N_4590,N_3406,N_3523);
and U4591 (N_4591,N_3067,N_3930);
nand U4592 (N_4592,N_3267,N_3537);
or U4593 (N_4593,N_3179,N_3358);
and U4594 (N_4594,N_3525,N_3304);
nor U4595 (N_4595,N_3610,N_3196);
nand U4596 (N_4596,N_3724,N_3485);
nand U4597 (N_4597,N_3656,N_3367);
xor U4598 (N_4598,N_3210,N_3487);
nand U4599 (N_4599,N_3701,N_3762);
nand U4600 (N_4600,N_3563,N_3270);
nor U4601 (N_4601,N_3617,N_3773);
or U4602 (N_4602,N_3588,N_3627);
nor U4603 (N_4603,N_3587,N_3624);
or U4604 (N_4604,N_3971,N_3426);
nor U4605 (N_4605,N_3431,N_3677);
nor U4606 (N_4606,N_3448,N_3445);
and U4607 (N_4607,N_3035,N_3443);
nand U4608 (N_4608,N_3695,N_3790);
xor U4609 (N_4609,N_3887,N_3742);
nand U4610 (N_4610,N_3075,N_3536);
or U4611 (N_4611,N_3689,N_3032);
or U4612 (N_4612,N_3846,N_3019);
xnor U4613 (N_4613,N_3937,N_3112);
xor U4614 (N_4614,N_3095,N_3791);
or U4615 (N_4615,N_3845,N_3390);
nor U4616 (N_4616,N_3589,N_3738);
and U4617 (N_4617,N_3235,N_3507);
nor U4618 (N_4618,N_3764,N_3763);
nor U4619 (N_4619,N_3812,N_3641);
and U4620 (N_4620,N_3363,N_3045);
xor U4621 (N_4621,N_3213,N_3140);
nor U4622 (N_4622,N_3231,N_3216);
xor U4623 (N_4623,N_3577,N_3916);
nor U4624 (N_4624,N_3762,N_3606);
xnor U4625 (N_4625,N_3294,N_3508);
or U4626 (N_4626,N_3387,N_3355);
xnor U4627 (N_4627,N_3605,N_3035);
nor U4628 (N_4628,N_3841,N_3549);
xor U4629 (N_4629,N_3451,N_3376);
and U4630 (N_4630,N_3063,N_3864);
nor U4631 (N_4631,N_3127,N_3461);
and U4632 (N_4632,N_3499,N_3653);
xor U4633 (N_4633,N_3604,N_3652);
nor U4634 (N_4634,N_3705,N_3128);
or U4635 (N_4635,N_3113,N_3715);
xnor U4636 (N_4636,N_3481,N_3988);
nor U4637 (N_4637,N_3135,N_3028);
and U4638 (N_4638,N_3483,N_3243);
and U4639 (N_4639,N_3291,N_3437);
xnor U4640 (N_4640,N_3007,N_3478);
nand U4641 (N_4641,N_3567,N_3892);
xor U4642 (N_4642,N_3290,N_3014);
and U4643 (N_4643,N_3929,N_3555);
nand U4644 (N_4644,N_3570,N_3686);
nand U4645 (N_4645,N_3400,N_3094);
xor U4646 (N_4646,N_3079,N_3405);
nor U4647 (N_4647,N_3838,N_3010);
nand U4648 (N_4648,N_3704,N_3224);
xor U4649 (N_4649,N_3288,N_3371);
nor U4650 (N_4650,N_3385,N_3324);
nor U4651 (N_4651,N_3878,N_3702);
nand U4652 (N_4652,N_3260,N_3352);
nor U4653 (N_4653,N_3048,N_3163);
and U4654 (N_4654,N_3227,N_3178);
and U4655 (N_4655,N_3051,N_3271);
or U4656 (N_4656,N_3309,N_3920);
xnor U4657 (N_4657,N_3017,N_3031);
xnor U4658 (N_4658,N_3154,N_3408);
xor U4659 (N_4659,N_3216,N_3502);
and U4660 (N_4660,N_3740,N_3133);
nor U4661 (N_4661,N_3779,N_3082);
nand U4662 (N_4662,N_3670,N_3163);
nor U4663 (N_4663,N_3565,N_3416);
or U4664 (N_4664,N_3226,N_3476);
or U4665 (N_4665,N_3430,N_3201);
nor U4666 (N_4666,N_3456,N_3710);
nand U4667 (N_4667,N_3768,N_3423);
and U4668 (N_4668,N_3929,N_3375);
and U4669 (N_4669,N_3367,N_3119);
and U4670 (N_4670,N_3195,N_3498);
or U4671 (N_4671,N_3284,N_3894);
or U4672 (N_4672,N_3729,N_3518);
and U4673 (N_4673,N_3127,N_3798);
or U4674 (N_4674,N_3340,N_3012);
and U4675 (N_4675,N_3671,N_3800);
nand U4676 (N_4676,N_3197,N_3561);
nor U4677 (N_4677,N_3162,N_3170);
or U4678 (N_4678,N_3138,N_3964);
or U4679 (N_4679,N_3501,N_3583);
nor U4680 (N_4680,N_3498,N_3964);
or U4681 (N_4681,N_3509,N_3940);
nor U4682 (N_4682,N_3146,N_3948);
nor U4683 (N_4683,N_3454,N_3220);
xnor U4684 (N_4684,N_3274,N_3349);
or U4685 (N_4685,N_3216,N_3114);
and U4686 (N_4686,N_3154,N_3559);
xnor U4687 (N_4687,N_3401,N_3995);
nand U4688 (N_4688,N_3204,N_3784);
or U4689 (N_4689,N_3626,N_3479);
and U4690 (N_4690,N_3280,N_3590);
nor U4691 (N_4691,N_3482,N_3048);
xnor U4692 (N_4692,N_3420,N_3689);
nor U4693 (N_4693,N_3318,N_3584);
nor U4694 (N_4694,N_3150,N_3208);
nand U4695 (N_4695,N_3410,N_3863);
nand U4696 (N_4696,N_3186,N_3000);
xnor U4697 (N_4697,N_3867,N_3199);
nor U4698 (N_4698,N_3604,N_3285);
nand U4699 (N_4699,N_3361,N_3462);
or U4700 (N_4700,N_3153,N_3700);
and U4701 (N_4701,N_3266,N_3660);
xnor U4702 (N_4702,N_3368,N_3124);
xor U4703 (N_4703,N_3186,N_3881);
or U4704 (N_4704,N_3454,N_3761);
nand U4705 (N_4705,N_3672,N_3015);
nand U4706 (N_4706,N_3109,N_3219);
xor U4707 (N_4707,N_3413,N_3565);
or U4708 (N_4708,N_3179,N_3112);
nor U4709 (N_4709,N_3271,N_3514);
xor U4710 (N_4710,N_3564,N_3196);
xnor U4711 (N_4711,N_3559,N_3429);
nor U4712 (N_4712,N_3495,N_3161);
xor U4713 (N_4713,N_3067,N_3100);
xnor U4714 (N_4714,N_3258,N_3296);
nand U4715 (N_4715,N_3996,N_3063);
xor U4716 (N_4716,N_3209,N_3844);
nand U4717 (N_4717,N_3916,N_3721);
and U4718 (N_4718,N_3607,N_3929);
nand U4719 (N_4719,N_3865,N_3153);
nor U4720 (N_4720,N_3298,N_3807);
and U4721 (N_4721,N_3076,N_3040);
nand U4722 (N_4722,N_3279,N_3471);
xnor U4723 (N_4723,N_3054,N_3083);
and U4724 (N_4724,N_3009,N_3371);
and U4725 (N_4725,N_3602,N_3664);
nand U4726 (N_4726,N_3141,N_3182);
xor U4727 (N_4727,N_3243,N_3643);
or U4728 (N_4728,N_3151,N_3131);
or U4729 (N_4729,N_3706,N_3121);
nand U4730 (N_4730,N_3004,N_3706);
nor U4731 (N_4731,N_3290,N_3098);
xnor U4732 (N_4732,N_3319,N_3744);
nor U4733 (N_4733,N_3989,N_3690);
and U4734 (N_4734,N_3299,N_3799);
nor U4735 (N_4735,N_3660,N_3812);
nand U4736 (N_4736,N_3981,N_3683);
nor U4737 (N_4737,N_3527,N_3023);
nor U4738 (N_4738,N_3901,N_3380);
xor U4739 (N_4739,N_3551,N_3646);
and U4740 (N_4740,N_3325,N_3362);
xnor U4741 (N_4741,N_3043,N_3044);
nor U4742 (N_4742,N_3350,N_3988);
xor U4743 (N_4743,N_3293,N_3149);
xnor U4744 (N_4744,N_3227,N_3020);
or U4745 (N_4745,N_3163,N_3360);
nor U4746 (N_4746,N_3862,N_3865);
or U4747 (N_4747,N_3814,N_3038);
nand U4748 (N_4748,N_3991,N_3081);
nor U4749 (N_4749,N_3847,N_3820);
and U4750 (N_4750,N_3528,N_3441);
nor U4751 (N_4751,N_3063,N_3059);
nor U4752 (N_4752,N_3387,N_3051);
or U4753 (N_4753,N_3559,N_3309);
and U4754 (N_4754,N_3537,N_3454);
xnor U4755 (N_4755,N_3988,N_3367);
nor U4756 (N_4756,N_3093,N_3832);
and U4757 (N_4757,N_3043,N_3754);
nor U4758 (N_4758,N_3646,N_3343);
nand U4759 (N_4759,N_3829,N_3386);
or U4760 (N_4760,N_3352,N_3172);
and U4761 (N_4761,N_3868,N_3476);
and U4762 (N_4762,N_3167,N_3088);
and U4763 (N_4763,N_3499,N_3844);
and U4764 (N_4764,N_3489,N_3755);
and U4765 (N_4765,N_3047,N_3555);
and U4766 (N_4766,N_3903,N_3342);
nand U4767 (N_4767,N_3770,N_3777);
or U4768 (N_4768,N_3255,N_3532);
and U4769 (N_4769,N_3616,N_3976);
and U4770 (N_4770,N_3993,N_3008);
or U4771 (N_4771,N_3544,N_3403);
nand U4772 (N_4772,N_3565,N_3527);
or U4773 (N_4773,N_3897,N_3091);
xor U4774 (N_4774,N_3886,N_3656);
nand U4775 (N_4775,N_3101,N_3920);
and U4776 (N_4776,N_3773,N_3082);
and U4777 (N_4777,N_3107,N_3695);
or U4778 (N_4778,N_3976,N_3204);
nand U4779 (N_4779,N_3749,N_3978);
nor U4780 (N_4780,N_3437,N_3240);
nand U4781 (N_4781,N_3933,N_3525);
or U4782 (N_4782,N_3552,N_3952);
xor U4783 (N_4783,N_3172,N_3462);
and U4784 (N_4784,N_3868,N_3395);
nor U4785 (N_4785,N_3972,N_3606);
nand U4786 (N_4786,N_3243,N_3554);
nor U4787 (N_4787,N_3570,N_3719);
and U4788 (N_4788,N_3908,N_3362);
xor U4789 (N_4789,N_3090,N_3122);
nor U4790 (N_4790,N_3036,N_3113);
and U4791 (N_4791,N_3978,N_3858);
nand U4792 (N_4792,N_3733,N_3695);
xnor U4793 (N_4793,N_3345,N_3758);
nand U4794 (N_4794,N_3321,N_3931);
xnor U4795 (N_4795,N_3374,N_3228);
nand U4796 (N_4796,N_3857,N_3731);
or U4797 (N_4797,N_3728,N_3410);
nor U4798 (N_4798,N_3673,N_3602);
xor U4799 (N_4799,N_3250,N_3764);
nand U4800 (N_4800,N_3490,N_3737);
and U4801 (N_4801,N_3553,N_3509);
or U4802 (N_4802,N_3440,N_3903);
and U4803 (N_4803,N_3393,N_3831);
nor U4804 (N_4804,N_3426,N_3942);
xor U4805 (N_4805,N_3939,N_3841);
and U4806 (N_4806,N_3194,N_3270);
or U4807 (N_4807,N_3421,N_3966);
nor U4808 (N_4808,N_3605,N_3530);
xor U4809 (N_4809,N_3719,N_3051);
and U4810 (N_4810,N_3721,N_3749);
and U4811 (N_4811,N_3292,N_3939);
nand U4812 (N_4812,N_3087,N_3562);
xor U4813 (N_4813,N_3336,N_3664);
nand U4814 (N_4814,N_3644,N_3906);
and U4815 (N_4815,N_3312,N_3623);
and U4816 (N_4816,N_3310,N_3470);
xor U4817 (N_4817,N_3812,N_3902);
nor U4818 (N_4818,N_3673,N_3003);
nor U4819 (N_4819,N_3544,N_3614);
xor U4820 (N_4820,N_3273,N_3884);
xor U4821 (N_4821,N_3274,N_3136);
nand U4822 (N_4822,N_3518,N_3509);
nor U4823 (N_4823,N_3454,N_3695);
or U4824 (N_4824,N_3027,N_3124);
xnor U4825 (N_4825,N_3122,N_3739);
xnor U4826 (N_4826,N_3073,N_3723);
nor U4827 (N_4827,N_3495,N_3214);
and U4828 (N_4828,N_3466,N_3186);
and U4829 (N_4829,N_3820,N_3530);
nor U4830 (N_4830,N_3010,N_3123);
nand U4831 (N_4831,N_3592,N_3886);
nand U4832 (N_4832,N_3517,N_3138);
nor U4833 (N_4833,N_3858,N_3191);
and U4834 (N_4834,N_3184,N_3095);
or U4835 (N_4835,N_3180,N_3912);
or U4836 (N_4836,N_3922,N_3155);
and U4837 (N_4837,N_3026,N_3884);
nand U4838 (N_4838,N_3511,N_3442);
xor U4839 (N_4839,N_3877,N_3846);
nand U4840 (N_4840,N_3439,N_3589);
and U4841 (N_4841,N_3748,N_3605);
nand U4842 (N_4842,N_3818,N_3098);
nand U4843 (N_4843,N_3592,N_3305);
nand U4844 (N_4844,N_3764,N_3059);
nor U4845 (N_4845,N_3349,N_3617);
nand U4846 (N_4846,N_3853,N_3001);
or U4847 (N_4847,N_3298,N_3468);
nand U4848 (N_4848,N_3618,N_3001);
xnor U4849 (N_4849,N_3446,N_3134);
xnor U4850 (N_4850,N_3572,N_3560);
or U4851 (N_4851,N_3141,N_3747);
or U4852 (N_4852,N_3468,N_3524);
and U4853 (N_4853,N_3979,N_3060);
and U4854 (N_4854,N_3927,N_3819);
nand U4855 (N_4855,N_3671,N_3218);
nor U4856 (N_4856,N_3311,N_3826);
and U4857 (N_4857,N_3076,N_3475);
or U4858 (N_4858,N_3707,N_3426);
or U4859 (N_4859,N_3576,N_3101);
xor U4860 (N_4860,N_3653,N_3873);
or U4861 (N_4861,N_3883,N_3831);
nand U4862 (N_4862,N_3402,N_3298);
xor U4863 (N_4863,N_3141,N_3763);
nor U4864 (N_4864,N_3017,N_3353);
nor U4865 (N_4865,N_3352,N_3297);
xor U4866 (N_4866,N_3357,N_3018);
xnor U4867 (N_4867,N_3424,N_3920);
nand U4868 (N_4868,N_3003,N_3838);
xnor U4869 (N_4869,N_3073,N_3964);
or U4870 (N_4870,N_3719,N_3897);
or U4871 (N_4871,N_3832,N_3909);
nor U4872 (N_4872,N_3581,N_3421);
or U4873 (N_4873,N_3577,N_3774);
or U4874 (N_4874,N_3634,N_3136);
xnor U4875 (N_4875,N_3176,N_3443);
nand U4876 (N_4876,N_3013,N_3402);
xor U4877 (N_4877,N_3482,N_3921);
and U4878 (N_4878,N_3369,N_3532);
or U4879 (N_4879,N_3757,N_3908);
or U4880 (N_4880,N_3764,N_3885);
xnor U4881 (N_4881,N_3851,N_3129);
nand U4882 (N_4882,N_3017,N_3225);
nor U4883 (N_4883,N_3641,N_3639);
nor U4884 (N_4884,N_3832,N_3702);
xnor U4885 (N_4885,N_3950,N_3423);
or U4886 (N_4886,N_3637,N_3226);
xnor U4887 (N_4887,N_3325,N_3966);
nor U4888 (N_4888,N_3924,N_3960);
or U4889 (N_4889,N_3433,N_3768);
xnor U4890 (N_4890,N_3694,N_3652);
and U4891 (N_4891,N_3338,N_3367);
and U4892 (N_4892,N_3930,N_3357);
nand U4893 (N_4893,N_3232,N_3216);
nor U4894 (N_4894,N_3960,N_3139);
nor U4895 (N_4895,N_3247,N_3813);
and U4896 (N_4896,N_3009,N_3339);
nand U4897 (N_4897,N_3411,N_3262);
xor U4898 (N_4898,N_3894,N_3536);
or U4899 (N_4899,N_3364,N_3775);
nor U4900 (N_4900,N_3792,N_3205);
and U4901 (N_4901,N_3756,N_3374);
nand U4902 (N_4902,N_3725,N_3928);
and U4903 (N_4903,N_3518,N_3093);
nor U4904 (N_4904,N_3747,N_3438);
or U4905 (N_4905,N_3925,N_3341);
nor U4906 (N_4906,N_3720,N_3429);
and U4907 (N_4907,N_3540,N_3875);
nor U4908 (N_4908,N_3793,N_3547);
nor U4909 (N_4909,N_3217,N_3953);
or U4910 (N_4910,N_3464,N_3467);
nand U4911 (N_4911,N_3372,N_3514);
or U4912 (N_4912,N_3069,N_3730);
nand U4913 (N_4913,N_3953,N_3963);
nor U4914 (N_4914,N_3426,N_3536);
xor U4915 (N_4915,N_3499,N_3420);
xnor U4916 (N_4916,N_3029,N_3554);
xor U4917 (N_4917,N_3960,N_3844);
xnor U4918 (N_4918,N_3029,N_3121);
or U4919 (N_4919,N_3854,N_3442);
or U4920 (N_4920,N_3346,N_3660);
and U4921 (N_4921,N_3353,N_3383);
xnor U4922 (N_4922,N_3244,N_3785);
xnor U4923 (N_4923,N_3647,N_3300);
nand U4924 (N_4924,N_3825,N_3910);
nand U4925 (N_4925,N_3107,N_3820);
or U4926 (N_4926,N_3076,N_3581);
or U4927 (N_4927,N_3450,N_3660);
nand U4928 (N_4928,N_3245,N_3220);
or U4929 (N_4929,N_3434,N_3233);
nor U4930 (N_4930,N_3085,N_3429);
or U4931 (N_4931,N_3369,N_3005);
or U4932 (N_4932,N_3862,N_3368);
nand U4933 (N_4933,N_3062,N_3864);
nor U4934 (N_4934,N_3038,N_3680);
or U4935 (N_4935,N_3689,N_3505);
or U4936 (N_4936,N_3090,N_3293);
or U4937 (N_4937,N_3666,N_3514);
nor U4938 (N_4938,N_3243,N_3039);
xnor U4939 (N_4939,N_3779,N_3623);
xnor U4940 (N_4940,N_3044,N_3066);
nor U4941 (N_4941,N_3341,N_3186);
nand U4942 (N_4942,N_3986,N_3254);
and U4943 (N_4943,N_3591,N_3277);
nor U4944 (N_4944,N_3390,N_3151);
xnor U4945 (N_4945,N_3959,N_3348);
nor U4946 (N_4946,N_3470,N_3713);
nor U4947 (N_4947,N_3228,N_3271);
nor U4948 (N_4948,N_3606,N_3129);
or U4949 (N_4949,N_3998,N_3503);
and U4950 (N_4950,N_3417,N_3776);
nor U4951 (N_4951,N_3203,N_3347);
nor U4952 (N_4952,N_3053,N_3891);
nand U4953 (N_4953,N_3935,N_3824);
nand U4954 (N_4954,N_3476,N_3848);
nor U4955 (N_4955,N_3328,N_3538);
nor U4956 (N_4956,N_3431,N_3918);
or U4957 (N_4957,N_3967,N_3555);
xnor U4958 (N_4958,N_3539,N_3628);
nand U4959 (N_4959,N_3353,N_3338);
nand U4960 (N_4960,N_3647,N_3687);
nand U4961 (N_4961,N_3430,N_3217);
xnor U4962 (N_4962,N_3801,N_3822);
nand U4963 (N_4963,N_3871,N_3163);
nand U4964 (N_4964,N_3363,N_3393);
and U4965 (N_4965,N_3363,N_3599);
or U4966 (N_4966,N_3054,N_3383);
and U4967 (N_4967,N_3960,N_3813);
nor U4968 (N_4968,N_3685,N_3614);
nand U4969 (N_4969,N_3985,N_3331);
xnor U4970 (N_4970,N_3415,N_3736);
nor U4971 (N_4971,N_3902,N_3152);
and U4972 (N_4972,N_3266,N_3595);
nor U4973 (N_4973,N_3474,N_3802);
and U4974 (N_4974,N_3611,N_3850);
and U4975 (N_4975,N_3947,N_3536);
or U4976 (N_4976,N_3955,N_3640);
nand U4977 (N_4977,N_3565,N_3356);
and U4978 (N_4978,N_3740,N_3181);
and U4979 (N_4979,N_3421,N_3798);
nor U4980 (N_4980,N_3453,N_3405);
nor U4981 (N_4981,N_3119,N_3445);
or U4982 (N_4982,N_3271,N_3707);
nand U4983 (N_4983,N_3019,N_3636);
nand U4984 (N_4984,N_3266,N_3581);
and U4985 (N_4985,N_3263,N_3069);
nor U4986 (N_4986,N_3133,N_3574);
and U4987 (N_4987,N_3216,N_3221);
nand U4988 (N_4988,N_3491,N_3123);
and U4989 (N_4989,N_3764,N_3016);
nand U4990 (N_4990,N_3680,N_3390);
nor U4991 (N_4991,N_3706,N_3643);
or U4992 (N_4992,N_3834,N_3726);
xnor U4993 (N_4993,N_3876,N_3150);
or U4994 (N_4994,N_3418,N_3945);
nand U4995 (N_4995,N_3042,N_3142);
or U4996 (N_4996,N_3263,N_3340);
xor U4997 (N_4997,N_3906,N_3422);
nand U4998 (N_4998,N_3228,N_3642);
or U4999 (N_4999,N_3960,N_3164);
or U5000 (N_5000,N_4703,N_4083);
and U5001 (N_5001,N_4678,N_4378);
or U5002 (N_5002,N_4669,N_4324);
or U5003 (N_5003,N_4437,N_4273);
nor U5004 (N_5004,N_4906,N_4836);
nor U5005 (N_5005,N_4412,N_4918);
nor U5006 (N_5006,N_4450,N_4851);
xnor U5007 (N_5007,N_4321,N_4817);
nor U5008 (N_5008,N_4980,N_4018);
xnor U5009 (N_5009,N_4650,N_4184);
xnor U5010 (N_5010,N_4861,N_4045);
nand U5011 (N_5011,N_4332,N_4300);
xnor U5012 (N_5012,N_4012,N_4544);
or U5013 (N_5013,N_4216,N_4206);
and U5014 (N_5014,N_4598,N_4341);
and U5015 (N_5015,N_4171,N_4038);
and U5016 (N_5016,N_4656,N_4722);
and U5017 (N_5017,N_4082,N_4478);
nand U5018 (N_5018,N_4144,N_4842);
nand U5019 (N_5019,N_4953,N_4863);
nor U5020 (N_5020,N_4556,N_4788);
xor U5021 (N_5021,N_4853,N_4510);
or U5022 (N_5022,N_4467,N_4183);
nor U5023 (N_5023,N_4127,N_4536);
nor U5024 (N_5024,N_4814,N_4513);
nand U5025 (N_5025,N_4696,N_4560);
nor U5026 (N_5026,N_4800,N_4545);
and U5027 (N_5027,N_4952,N_4472);
nor U5028 (N_5028,N_4626,N_4298);
nor U5029 (N_5029,N_4811,N_4525);
nand U5030 (N_5030,N_4282,N_4373);
nand U5031 (N_5031,N_4710,N_4465);
and U5032 (N_5032,N_4998,N_4652);
xnor U5033 (N_5033,N_4326,N_4864);
or U5034 (N_5034,N_4019,N_4844);
or U5035 (N_5035,N_4312,N_4926);
and U5036 (N_5036,N_4624,N_4944);
and U5037 (N_5037,N_4460,N_4674);
or U5038 (N_5038,N_4187,N_4190);
or U5039 (N_5039,N_4782,N_4035);
nor U5040 (N_5040,N_4774,N_4075);
xor U5041 (N_5041,N_4801,N_4633);
nor U5042 (N_5042,N_4812,N_4330);
xor U5043 (N_5043,N_4580,N_4494);
xnor U5044 (N_5044,N_4641,N_4399);
nor U5045 (N_5045,N_4431,N_4739);
or U5046 (N_5046,N_4573,N_4942);
or U5047 (N_5047,N_4567,N_4512);
or U5048 (N_5048,N_4319,N_4791);
and U5049 (N_5049,N_4483,N_4078);
xnor U5050 (N_5050,N_4359,N_4098);
nand U5051 (N_5051,N_4753,N_4742);
nand U5052 (N_5052,N_4167,N_4644);
nor U5053 (N_5053,N_4348,N_4284);
nand U5054 (N_5054,N_4605,N_4676);
xnor U5055 (N_5055,N_4766,N_4733);
or U5056 (N_5056,N_4162,N_4995);
or U5057 (N_5057,N_4873,N_4530);
or U5058 (N_5058,N_4455,N_4161);
xnor U5059 (N_5059,N_4013,N_4654);
nand U5060 (N_5060,N_4438,N_4526);
nand U5061 (N_5061,N_4846,N_4236);
or U5062 (N_5062,N_4961,N_4316);
and U5063 (N_5063,N_4666,N_4769);
nand U5064 (N_5064,N_4585,N_4519);
and U5065 (N_5065,N_4268,N_4921);
xnor U5066 (N_5066,N_4429,N_4854);
nor U5067 (N_5067,N_4278,N_4398);
xnor U5068 (N_5068,N_4761,N_4289);
or U5069 (N_5069,N_4349,N_4446);
nand U5070 (N_5070,N_4317,N_4142);
nor U5071 (N_5071,N_4339,N_4743);
or U5072 (N_5072,N_4571,N_4880);
and U5073 (N_5073,N_4597,N_4361);
and U5074 (N_5074,N_4988,N_4625);
nand U5075 (N_5075,N_4740,N_4306);
and U5076 (N_5076,N_4199,N_4186);
and U5077 (N_5077,N_4777,N_4476);
nand U5078 (N_5078,N_4837,N_4705);
and U5079 (N_5079,N_4415,N_4681);
or U5080 (N_5080,N_4645,N_4391);
xnor U5081 (N_5081,N_4305,N_4062);
or U5082 (N_5082,N_4139,N_4253);
nand U5083 (N_5083,N_4581,N_4719);
nand U5084 (N_5084,N_4040,N_4074);
nor U5085 (N_5085,N_4978,N_4870);
xor U5086 (N_5086,N_4749,N_4824);
or U5087 (N_5087,N_4879,N_4640);
nand U5088 (N_5088,N_4671,N_4243);
or U5089 (N_5089,N_4862,N_4516);
nand U5090 (N_5090,N_4302,N_4185);
xnor U5091 (N_5091,N_4986,N_4602);
nand U5092 (N_5092,N_4310,N_4783);
nand U5093 (N_5093,N_4693,N_4596);
and U5094 (N_5094,N_4444,N_4591);
and U5095 (N_5095,N_4132,N_4843);
xor U5096 (N_5096,N_4049,N_4754);
nand U5097 (N_5097,N_4210,N_4936);
or U5098 (N_5098,N_4535,N_4972);
nor U5099 (N_5099,N_4418,N_4343);
nand U5100 (N_5100,N_4576,N_4825);
nand U5101 (N_5101,N_4173,N_4487);
or U5102 (N_5102,N_4260,N_4785);
xnor U5103 (N_5103,N_4727,N_4159);
nor U5104 (N_5104,N_4557,N_4683);
nor U5105 (N_5105,N_4642,N_4355);
nand U5106 (N_5106,N_4432,N_4741);
nor U5107 (N_5107,N_4937,N_4331);
nor U5108 (N_5108,N_4290,N_4885);
xnor U5109 (N_5109,N_4589,N_4612);
or U5110 (N_5110,N_4393,N_4120);
and U5111 (N_5111,N_4929,N_4072);
and U5112 (N_5112,N_4107,N_4096);
xnor U5113 (N_5113,N_4820,N_4165);
nand U5114 (N_5114,N_4354,N_4639);
xnor U5115 (N_5115,N_4871,N_4225);
xor U5116 (N_5116,N_4117,N_4275);
and U5117 (N_5117,N_4932,N_4868);
nor U5118 (N_5118,N_4858,N_4473);
nand U5119 (N_5119,N_4549,N_4848);
xnor U5120 (N_5120,N_4907,N_4985);
xor U5121 (N_5121,N_4299,N_4307);
xnor U5122 (N_5122,N_4922,N_4500);
or U5123 (N_5123,N_4601,N_4070);
and U5124 (N_5124,N_4170,N_4169);
or U5125 (N_5125,N_4517,N_4927);
or U5126 (N_5126,N_4747,N_4276);
or U5127 (N_5127,N_4659,N_4638);
and U5128 (N_5128,N_4118,N_4583);
and U5129 (N_5129,N_4518,N_4720);
or U5130 (N_5130,N_4689,N_4283);
and U5131 (N_5131,N_4826,N_4352);
and U5132 (N_5132,N_4750,N_4439);
or U5133 (N_5133,N_4179,N_4541);
or U5134 (N_5134,N_4505,N_4706);
nand U5135 (N_5135,N_4149,N_4288);
xnor U5136 (N_5136,N_4262,N_4130);
nor U5137 (N_5137,N_4376,N_4657);
nand U5138 (N_5138,N_4277,N_4246);
xor U5139 (N_5139,N_4265,N_4385);
xor U5140 (N_5140,N_4529,N_4895);
nand U5141 (N_5141,N_4835,N_4579);
and U5142 (N_5142,N_4039,N_4548);
nor U5143 (N_5143,N_4708,N_4396);
and U5144 (N_5144,N_4053,N_4292);
nor U5145 (N_5145,N_4435,N_4353);
or U5146 (N_5146,N_4014,N_4030);
or U5147 (N_5147,N_4114,N_4469);
xnor U5148 (N_5148,N_4663,N_4409);
xnor U5149 (N_5149,N_4925,N_4136);
and U5150 (N_5150,N_4798,N_4402);
nand U5151 (N_5151,N_4152,N_4109);
xor U5152 (N_5152,N_4617,N_4570);
or U5153 (N_5153,N_4255,N_4017);
or U5154 (N_5154,N_4397,N_4784);
or U5155 (N_5155,N_4872,N_4966);
xor U5156 (N_5156,N_4023,N_4866);
nor U5157 (N_5157,N_4508,N_4347);
xnor U5158 (N_5158,N_4630,N_4375);
nor U5159 (N_5159,N_4911,N_4955);
xnor U5160 (N_5160,N_4827,N_4293);
nor U5161 (N_5161,N_4211,N_4055);
nand U5162 (N_5162,N_4855,N_4713);
and U5163 (N_5163,N_4259,N_4226);
and U5164 (N_5164,N_4884,N_4314);
nand U5165 (N_5165,N_4110,N_4101);
xnor U5166 (N_5166,N_4809,N_4538);
nor U5167 (N_5167,N_4830,N_4463);
nor U5168 (N_5168,N_4767,N_4247);
xnor U5169 (N_5169,N_4680,N_4213);
nor U5170 (N_5170,N_4458,N_4857);
and U5171 (N_5171,N_4943,N_4725);
nor U5172 (N_5172,N_4176,N_4406);
and U5173 (N_5173,N_4905,N_4655);
and U5174 (N_5174,N_4155,N_4087);
and U5175 (N_5175,N_4815,N_4094);
nand U5176 (N_5176,N_4203,N_4987);
nand U5177 (N_5177,N_4577,N_4968);
nand U5178 (N_5178,N_4464,N_4090);
or U5179 (N_5179,N_4896,N_4231);
nor U5180 (N_5180,N_4021,N_4894);
nand U5181 (N_5181,N_4540,N_4294);
or U5182 (N_5182,N_4672,N_4636);
nor U5183 (N_5183,N_4658,N_4502);
nor U5184 (N_5184,N_4603,N_4550);
or U5185 (N_5185,N_4223,N_4521);
xor U5186 (N_5186,N_4939,N_4474);
xnor U5187 (N_5187,N_4917,N_4759);
nor U5188 (N_5188,N_4252,N_4578);
xnor U5189 (N_5189,N_4876,N_4982);
nand U5190 (N_5190,N_4615,N_4191);
and U5191 (N_5191,N_4366,N_4551);
nor U5192 (N_5192,N_4042,N_4441);
xor U5193 (N_5193,N_4177,N_4200);
and U5194 (N_5194,N_4228,N_4008);
nand U5195 (N_5195,N_4893,N_4790);
or U5196 (N_5196,N_4215,N_4734);
nor U5197 (N_5197,N_4239,N_4037);
xor U5198 (N_5198,N_4643,N_4924);
nor U5199 (N_5199,N_4054,N_4606);
nor U5200 (N_5200,N_4420,N_4569);
nor U5201 (N_5201,N_4491,N_4287);
nand U5202 (N_5202,N_4621,N_4524);
nor U5203 (N_5203,N_4975,N_4224);
nand U5204 (N_5204,N_4852,N_4977);
xnor U5205 (N_5205,N_4609,N_4908);
nor U5206 (N_5206,N_4841,N_4338);
xor U5207 (N_5207,N_4729,N_4202);
xor U5208 (N_5208,N_4003,N_4765);
xnor U5209 (N_5209,N_4448,N_4095);
nand U5210 (N_5210,N_4555,N_4220);
nor U5211 (N_5211,N_4970,N_4468);
xor U5212 (N_5212,N_4974,N_4000);
xnor U5213 (N_5213,N_4610,N_4964);
nor U5214 (N_5214,N_4065,N_4954);
and U5215 (N_5215,N_4414,N_4794);
nor U5216 (N_5216,N_4073,N_4365);
and U5217 (N_5217,N_4963,N_4157);
nand U5218 (N_5218,N_4384,N_4553);
or U5219 (N_5219,N_4335,N_4103);
and U5220 (N_5220,N_4533,N_4562);
or U5221 (N_5221,N_4682,N_4482);
and U5222 (N_5222,N_4377,N_4543);
nor U5223 (N_5223,N_4140,N_4303);
nand U5224 (N_5224,N_4261,N_4833);
xnor U5225 (N_5225,N_4614,N_4697);
or U5226 (N_5226,N_4245,N_4229);
nor U5227 (N_5227,N_4126,N_4822);
or U5228 (N_5228,N_4803,N_4718);
nor U5229 (N_5229,N_4208,N_4297);
nand U5230 (N_5230,N_4272,N_4058);
nand U5231 (N_5231,N_4956,N_4492);
or U5232 (N_5232,N_4732,N_4388);
or U5233 (N_5233,N_4582,N_4285);
nand U5234 (N_5234,N_4156,N_4691);
and U5235 (N_5235,N_4763,N_4269);
nand U5236 (N_5236,N_4207,N_4586);
nor U5237 (N_5237,N_4235,N_4909);
xor U5238 (N_5238,N_4537,N_4622);
xnor U5239 (N_5239,N_4209,N_4411);
xor U5240 (N_5240,N_4821,N_4504);
nand U5241 (N_5241,N_4592,N_4426);
xnor U5242 (N_5242,N_4600,N_4296);
and U5243 (N_5243,N_4068,N_4634);
and U5244 (N_5244,N_4534,N_4877);
and U5245 (N_5245,N_4813,N_4695);
and U5246 (N_5246,N_4238,N_4775);
xor U5247 (N_5247,N_4395,N_4079);
or U5248 (N_5248,N_4903,N_4527);
or U5249 (N_5249,N_4996,N_4829);
and U5250 (N_5250,N_4242,N_4340);
nor U5251 (N_5251,N_4145,N_4370);
and U5252 (N_5252,N_4506,N_4198);
nand U5253 (N_5253,N_4383,N_4020);
nand U5254 (N_5254,N_4459,N_4707);
xor U5255 (N_5255,N_4400,N_4499);
nand U5256 (N_5256,N_4475,N_4607);
nand U5257 (N_5257,N_4313,N_4892);
nor U5258 (N_5258,N_4781,N_4434);
xnor U5259 (N_5259,N_4367,N_4889);
xor U5260 (N_5260,N_4805,N_4041);
or U5261 (N_5261,N_4291,N_4709);
and U5262 (N_5262,N_4337,N_4687);
xnor U5263 (N_5263,N_4670,N_4845);
or U5264 (N_5264,N_4133,N_4883);
xor U5265 (N_5265,N_4227,N_4838);
or U5266 (N_5266,N_4738,N_4479);
nor U5267 (N_5267,N_4009,N_4685);
xor U5268 (N_5268,N_4731,N_4452);
or U5269 (N_5269,N_4430,N_4699);
nor U5270 (N_5270,N_4890,N_4280);
nand U5271 (N_5271,N_4566,N_4802);
xnor U5272 (N_5272,N_4758,N_4902);
and U5273 (N_5273,N_4150,N_4116);
or U5274 (N_5274,N_4688,N_4250);
and U5275 (N_5275,N_4528,N_4135);
and U5276 (N_5276,N_4881,N_4613);
and U5277 (N_5277,N_4451,N_4865);
nor U5278 (N_5278,N_4005,N_4967);
and U5279 (N_5279,N_4686,N_4477);
xor U5280 (N_5280,N_4050,N_4333);
and U5281 (N_5281,N_4847,N_4181);
and U5282 (N_5282,N_4559,N_4588);
or U5283 (N_5283,N_4962,N_4714);
or U5284 (N_5284,N_4919,N_4983);
or U5285 (N_5285,N_4401,N_4295);
and U5286 (N_5286,N_4979,N_4445);
and U5287 (N_5287,N_4113,N_4819);
nor U5288 (N_5288,N_4369,N_4867);
nand U5289 (N_5289,N_4026,N_4665);
or U5290 (N_5290,N_4997,N_4322);
and U5291 (N_5291,N_4102,N_4793);
nor U5292 (N_5292,N_4172,N_4311);
and U5293 (N_5293,N_4016,N_4115);
nor U5294 (N_5294,N_4795,N_4490);
and U5295 (N_5295,N_4141,N_4823);
and U5296 (N_5296,N_4351,N_4147);
and U5297 (N_5297,N_4219,N_4779);
and U5298 (N_5298,N_4770,N_4515);
xor U5299 (N_5299,N_4148,N_4859);
xor U5300 (N_5300,N_4485,N_4044);
nor U5301 (N_5301,N_4520,N_4736);
and U5302 (N_5302,N_4694,N_4047);
nor U5303 (N_5303,N_4060,N_4461);
nor U5304 (N_5304,N_4635,N_4850);
nand U5305 (N_5305,N_4933,N_4561);
or U5306 (N_5306,N_4522,N_4104);
or U5307 (N_5307,N_4704,N_4345);
or U5308 (N_5308,N_4002,N_4608);
nand U5309 (N_5309,N_4711,N_4941);
and U5310 (N_5310,N_4668,N_4945);
or U5311 (N_5311,N_4488,N_4584);
and U5312 (N_5312,N_4724,N_4427);
xnor U5313 (N_5313,N_4503,N_4489);
xnor U5314 (N_5314,N_4137,N_4542);
or U5315 (N_5315,N_4721,N_4799);
nor U5316 (N_5316,N_4028,N_4368);
or U5317 (N_5317,N_4604,N_4684);
nor U5318 (N_5318,N_4886,N_4574);
and U5319 (N_5319,N_4234,N_4390);
xnor U5320 (N_5320,N_4737,N_4957);
nor U5321 (N_5321,N_4898,N_4660);
or U5322 (N_5322,N_4565,N_4723);
or U5323 (N_5323,N_4973,N_4947);
and U5324 (N_5324,N_4457,N_4934);
nor U5325 (N_5325,N_4204,N_4912);
and U5326 (N_5326,N_4218,N_4806);
xnor U5327 (N_5327,N_4100,N_4935);
and U5328 (N_5328,N_4389,N_4080);
xnor U5329 (N_5329,N_4648,N_4990);
and U5330 (N_5330,N_4931,N_4673);
or U5331 (N_5331,N_4914,N_4174);
nor U5332 (N_5332,N_4346,N_4514);
or U5333 (N_5333,N_4342,N_4221);
xor U5334 (N_5334,N_4364,N_4958);
or U5335 (N_5335,N_4256,N_4810);
or U5336 (N_5336,N_4497,N_4984);
nand U5337 (N_5337,N_4786,N_4563);
nand U5338 (N_5338,N_4304,N_4309);
nor U5339 (N_5339,N_4818,N_4436);
or U5340 (N_5340,N_4057,N_4197);
nor U5341 (N_5341,N_4279,N_4063);
nor U5342 (N_5342,N_4971,N_4632);
nor U5343 (N_5343,N_4664,N_4138);
and U5344 (N_5344,N_4748,N_4787);
or U5345 (N_5345,N_4532,N_4024);
and U5346 (N_5346,N_4547,N_4771);
nor U5347 (N_5347,N_4951,N_4920);
xor U5348 (N_5348,N_4649,N_4780);
and U5349 (N_5349,N_4735,N_4421);
nand U5350 (N_5350,N_4084,N_4052);
xnor U5351 (N_5351,N_4913,N_4946);
nand U5352 (N_5352,N_4433,N_4792);
or U5353 (N_5353,N_4010,N_4404);
xnor U5354 (N_5354,N_4362,N_4616);
or U5355 (N_5355,N_4493,N_4046);
and U5356 (N_5356,N_4056,N_4381);
nand U5357 (N_5357,N_4976,N_4158);
or U5358 (N_5358,N_4363,N_4027);
xnor U5359 (N_5359,N_4904,N_4992);
or U5360 (N_5360,N_4981,N_4051);
nand U5361 (N_5361,N_4900,N_4281);
and U5362 (N_5362,N_4011,N_4007);
nand U5363 (N_5363,N_4594,N_4356);
nor U5364 (N_5364,N_4745,N_4214);
and U5365 (N_5365,N_4081,N_4778);
and U5366 (N_5366,N_4129,N_4048);
nor U5367 (N_5367,N_4923,N_4568);
xnor U5368 (N_5368,N_4112,N_4440);
or U5369 (N_5369,N_4372,N_4274);
and U5370 (N_5370,N_4241,N_4222);
or U5371 (N_5371,N_4590,N_4428);
xnor U5372 (N_5372,N_4496,N_4085);
xor U5373 (N_5373,N_4449,N_4507);
or U5374 (N_5374,N_4205,N_4064);
nor U5375 (N_5375,N_4358,N_4267);
or U5376 (N_5376,N_4960,N_4481);
nand U5377 (N_5377,N_4646,N_4511);
xor U5378 (N_5378,N_4456,N_4106);
or U5379 (N_5379,N_4730,N_4258);
nand U5380 (N_5380,N_4611,N_4619);
nor U5381 (N_5381,N_4949,N_4772);
nand U5382 (N_5382,N_4965,N_4164);
xor U5383 (N_5383,N_4419,N_4128);
or U5384 (N_5384,N_4627,N_4856);
nor U5385 (N_5385,N_4371,N_4910);
xor U5386 (N_5386,N_4318,N_4816);
nand U5387 (N_5387,N_4797,N_4701);
or U5388 (N_5388,N_4762,N_4882);
and U5389 (N_5389,N_4595,N_4849);
nor U5390 (N_5390,N_4066,N_4599);
or U5391 (N_5391,N_4746,N_4160);
xnor U5392 (N_5392,N_4392,N_4999);
nor U5393 (N_5393,N_4755,N_4424);
xnor U5394 (N_5394,N_4264,N_4991);
nand U5395 (N_5395,N_4887,N_4938);
and U5396 (N_5396,N_4249,N_4717);
and U5397 (N_5397,N_4523,N_4334);
xor U5398 (N_5398,N_4470,N_4270);
nor U5399 (N_5399,N_4897,N_4410);
nand U5400 (N_5400,N_4061,N_4379);
or U5401 (N_5401,N_4327,N_4509);
xnor U5402 (N_5402,N_4131,N_4773);
or U5403 (N_5403,N_4558,N_4059);
and U5404 (N_5404,N_4153,N_4587);
nand U5405 (N_5405,N_4675,N_4832);
xnor U5406 (N_5406,N_4266,N_4423);
and U5407 (N_5407,N_4233,N_4989);
nor U5408 (N_5408,N_4564,N_4948);
nand U5409 (N_5409,N_4168,N_4025);
xnor U5410 (N_5410,N_4969,N_4629);
xor U5411 (N_5411,N_4325,N_4486);
or U5412 (N_5412,N_4146,N_4757);
xnor U5413 (N_5413,N_4993,N_4089);
or U5414 (N_5414,N_4768,N_4076);
nor U5415 (N_5415,N_4930,N_4618);
and U5416 (N_5416,N_4244,N_4254);
and U5417 (N_5417,N_4125,N_4143);
xnor U5418 (N_5418,N_4121,N_4099);
nand U5419 (N_5419,N_4271,N_4004);
nand U5420 (N_5420,N_4575,N_4201);
and U5421 (N_5421,N_4480,N_4928);
or U5422 (N_5422,N_4417,N_4808);
xor U5423 (N_5423,N_4552,N_4001);
and U5424 (N_5424,N_4408,N_4134);
nor U5425 (N_5425,N_4329,N_4531);
xor U5426 (N_5426,N_4006,N_4124);
and U5427 (N_5427,N_4336,N_4301);
nor U5428 (N_5428,N_4804,N_4405);
and U5429 (N_5429,N_4077,N_4036);
xnor U5430 (N_5430,N_4154,N_4495);
nand U5431 (N_5431,N_4442,N_4175);
and U5432 (N_5432,N_4623,N_4193);
nor U5433 (N_5433,N_4237,N_4069);
or U5434 (N_5434,N_4178,N_4751);
xnor U5435 (N_5435,N_4501,N_4093);
or U5436 (N_5436,N_4878,N_4031);
or U5437 (N_5437,N_4454,N_4484);
xor U5438 (N_5438,N_4915,N_4702);
xor U5439 (N_5439,N_4394,N_4959);
or U5440 (N_5440,N_4403,N_4189);
and U5441 (N_5441,N_4807,N_4471);
nand U5442 (N_5442,N_4123,N_4232);
nand U5443 (N_5443,N_4661,N_4029);
and U5444 (N_5444,N_4712,N_4443);
nand U5445 (N_5445,N_4653,N_4188);
xor U5446 (N_5446,N_4828,N_4033);
nand U5447 (N_5447,N_4539,N_4151);
xor U5448 (N_5448,N_4620,N_4180);
nor U5449 (N_5449,N_4860,N_4462);
and U5450 (N_5450,N_4756,N_4839);
and U5451 (N_5451,N_4466,N_4572);
and U5452 (N_5452,N_4899,N_4498);
and U5453 (N_5453,N_4086,N_4230);
xnor U5454 (N_5454,N_4195,N_4357);
or U5455 (N_5455,N_4088,N_4196);
xor U5456 (N_5456,N_4940,N_4308);
xnor U5457 (N_5457,N_4679,N_4840);
nand U5458 (N_5458,N_4092,N_4901);
nor U5459 (N_5459,N_4022,N_4263);
nand U5460 (N_5460,N_4163,N_4891);
nor U5461 (N_5461,N_4194,N_4067);
nor U5462 (N_5462,N_4015,N_4994);
and U5463 (N_5463,N_4108,N_4043);
xor U5464 (N_5464,N_4192,N_4760);
nand U5465 (N_5465,N_4315,N_4651);
xor U5466 (N_5466,N_4407,N_4286);
and U5467 (N_5467,N_4251,N_4764);
nor U5468 (N_5468,N_4628,N_4032);
and U5469 (N_5469,N_4119,N_4637);
or U5470 (N_5470,N_4111,N_4425);
nor U5471 (N_5471,N_4789,N_4212);
and U5472 (N_5472,N_4034,N_4320);
xor U5473 (N_5473,N_4240,N_4554);
xor U5474 (N_5474,N_4776,N_4105);
and U5475 (N_5475,N_4752,N_4667);
nor U5476 (N_5476,N_4698,N_4716);
and U5477 (N_5477,N_4182,N_4360);
nor U5478 (N_5478,N_4869,N_4453);
or U5479 (N_5479,N_4662,N_4328);
xor U5480 (N_5480,N_4374,N_4447);
nand U5481 (N_5481,N_4950,N_4631);
and U5482 (N_5482,N_4692,N_4593);
and U5483 (N_5483,N_4344,N_4690);
xnor U5484 (N_5484,N_4413,N_4916);
xor U5485 (N_5485,N_4217,N_4744);
nor U5486 (N_5486,N_4097,N_4834);
nor U5487 (N_5487,N_4796,N_4387);
or U5488 (N_5488,N_4715,N_4323);
or U5489 (N_5489,N_4071,N_4728);
xor U5490 (N_5490,N_4257,N_4874);
and U5491 (N_5491,N_4416,N_4888);
nand U5492 (N_5492,N_4700,N_4350);
xnor U5493 (N_5493,N_4677,N_4831);
and U5494 (N_5494,N_4546,N_4726);
and U5495 (N_5495,N_4422,N_4382);
and U5496 (N_5496,N_4091,N_4248);
xnor U5497 (N_5497,N_4386,N_4380);
xor U5498 (N_5498,N_4647,N_4875);
xor U5499 (N_5499,N_4122,N_4166);
and U5500 (N_5500,N_4479,N_4649);
or U5501 (N_5501,N_4312,N_4662);
nand U5502 (N_5502,N_4406,N_4993);
nand U5503 (N_5503,N_4506,N_4916);
or U5504 (N_5504,N_4640,N_4623);
or U5505 (N_5505,N_4495,N_4986);
and U5506 (N_5506,N_4554,N_4967);
xor U5507 (N_5507,N_4297,N_4594);
nor U5508 (N_5508,N_4089,N_4783);
and U5509 (N_5509,N_4136,N_4840);
xor U5510 (N_5510,N_4458,N_4309);
nand U5511 (N_5511,N_4308,N_4349);
and U5512 (N_5512,N_4107,N_4260);
and U5513 (N_5513,N_4790,N_4845);
nand U5514 (N_5514,N_4983,N_4253);
and U5515 (N_5515,N_4701,N_4282);
xor U5516 (N_5516,N_4683,N_4965);
xor U5517 (N_5517,N_4993,N_4515);
nand U5518 (N_5518,N_4822,N_4117);
nor U5519 (N_5519,N_4050,N_4936);
and U5520 (N_5520,N_4510,N_4032);
nand U5521 (N_5521,N_4022,N_4450);
nand U5522 (N_5522,N_4236,N_4980);
nor U5523 (N_5523,N_4626,N_4759);
nand U5524 (N_5524,N_4078,N_4762);
xnor U5525 (N_5525,N_4318,N_4908);
nand U5526 (N_5526,N_4269,N_4464);
xor U5527 (N_5527,N_4585,N_4738);
nand U5528 (N_5528,N_4531,N_4704);
xnor U5529 (N_5529,N_4400,N_4742);
nor U5530 (N_5530,N_4884,N_4097);
xnor U5531 (N_5531,N_4748,N_4658);
nand U5532 (N_5532,N_4258,N_4488);
nor U5533 (N_5533,N_4975,N_4910);
and U5534 (N_5534,N_4719,N_4598);
nand U5535 (N_5535,N_4721,N_4852);
and U5536 (N_5536,N_4104,N_4903);
xor U5537 (N_5537,N_4587,N_4664);
and U5538 (N_5538,N_4265,N_4195);
xnor U5539 (N_5539,N_4194,N_4886);
and U5540 (N_5540,N_4340,N_4796);
nand U5541 (N_5541,N_4850,N_4932);
or U5542 (N_5542,N_4549,N_4876);
nor U5543 (N_5543,N_4833,N_4411);
xor U5544 (N_5544,N_4376,N_4731);
or U5545 (N_5545,N_4832,N_4852);
and U5546 (N_5546,N_4712,N_4773);
or U5547 (N_5547,N_4343,N_4619);
or U5548 (N_5548,N_4972,N_4289);
nand U5549 (N_5549,N_4643,N_4517);
nor U5550 (N_5550,N_4221,N_4489);
and U5551 (N_5551,N_4830,N_4521);
and U5552 (N_5552,N_4998,N_4665);
nand U5553 (N_5553,N_4022,N_4367);
nand U5554 (N_5554,N_4962,N_4165);
nand U5555 (N_5555,N_4383,N_4378);
and U5556 (N_5556,N_4979,N_4703);
or U5557 (N_5557,N_4029,N_4395);
nand U5558 (N_5558,N_4225,N_4965);
xor U5559 (N_5559,N_4451,N_4740);
or U5560 (N_5560,N_4443,N_4388);
and U5561 (N_5561,N_4220,N_4691);
and U5562 (N_5562,N_4016,N_4894);
nand U5563 (N_5563,N_4298,N_4771);
nor U5564 (N_5564,N_4133,N_4532);
or U5565 (N_5565,N_4727,N_4228);
and U5566 (N_5566,N_4739,N_4215);
nor U5567 (N_5567,N_4365,N_4648);
and U5568 (N_5568,N_4886,N_4671);
nor U5569 (N_5569,N_4231,N_4289);
or U5570 (N_5570,N_4088,N_4913);
or U5571 (N_5571,N_4229,N_4153);
or U5572 (N_5572,N_4583,N_4739);
xnor U5573 (N_5573,N_4526,N_4897);
xor U5574 (N_5574,N_4238,N_4439);
and U5575 (N_5575,N_4199,N_4148);
nor U5576 (N_5576,N_4345,N_4944);
nand U5577 (N_5577,N_4003,N_4202);
nor U5578 (N_5578,N_4075,N_4556);
xnor U5579 (N_5579,N_4309,N_4835);
nand U5580 (N_5580,N_4517,N_4295);
and U5581 (N_5581,N_4671,N_4871);
and U5582 (N_5582,N_4454,N_4929);
or U5583 (N_5583,N_4875,N_4658);
nand U5584 (N_5584,N_4043,N_4322);
xor U5585 (N_5585,N_4001,N_4652);
or U5586 (N_5586,N_4152,N_4727);
or U5587 (N_5587,N_4217,N_4017);
nor U5588 (N_5588,N_4281,N_4897);
and U5589 (N_5589,N_4311,N_4543);
nor U5590 (N_5590,N_4073,N_4130);
xnor U5591 (N_5591,N_4595,N_4911);
and U5592 (N_5592,N_4605,N_4049);
nand U5593 (N_5593,N_4513,N_4176);
nand U5594 (N_5594,N_4565,N_4419);
xor U5595 (N_5595,N_4650,N_4461);
xor U5596 (N_5596,N_4263,N_4374);
and U5597 (N_5597,N_4664,N_4826);
and U5598 (N_5598,N_4895,N_4200);
xnor U5599 (N_5599,N_4883,N_4203);
xnor U5600 (N_5600,N_4076,N_4617);
and U5601 (N_5601,N_4700,N_4859);
or U5602 (N_5602,N_4428,N_4295);
nor U5603 (N_5603,N_4386,N_4892);
or U5604 (N_5604,N_4046,N_4049);
or U5605 (N_5605,N_4659,N_4479);
and U5606 (N_5606,N_4884,N_4456);
or U5607 (N_5607,N_4483,N_4511);
nand U5608 (N_5608,N_4728,N_4292);
nand U5609 (N_5609,N_4150,N_4751);
xnor U5610 (N_5610,N_4111,N_4082);
nand U5611 (N_5611,N_4635,N_4057);
and U5612 (N_5612,N_4961,N_4112);
nor U5613 (N_5613,N_4439,N_4772);
xor U5614 (N_5614,N_4427,N_4981);
and U5615 (N_5615,N_4793,N_4429);
and U5616 (N_5616,N_4447,N_4655);
xnor U5617 (N_5617,N_4409,N_4115);
xor U5618 (N_5618,N_4768,N_4857);
or U5619 (N_5619,N_4445,N_4588);
and U5620 (N_5620,N_4507,N_4167);
and U5621 (N_5621,N_4396,N_4913);
nor U5622 (N_5622,N_4592,N_4031);
and U5623 (N_5623,N_4583,N_4089);
and U5624 (N_5624,N_4937,N_4207);
and U5625 (N_5625,N_4460,N_4670);
and U5626 (N_5626,N_4928,N_4116);
and U5627 (N_5627,N_4510,N_4396);
and U5628 (N_5628,N_4567,N_4211);
and U5629 (N_5629,N_4235,N_4057);
and U5630 (N_5630,N_4049,N_4688);
nand U5631 (N_5631,N_4536,N_4643);
and U5632 (N_5632,N_4455,N_4784);
nor U5633 (N_5633,N_4501,N_4230);
nand U5634 (N_5634,N_4950,N_4537);
nor U5635 (N_5635,N_4517,N_4449);
or U5636 (N_5636,N_4228,N_4209);
nor U5637 (N_5637,N_4133,N_4361);
nor U5638 (N_5638,N_4805,N_4405);
or U5639 (N_5639,N_4839,N_4901);
and U5640 (N_5640,N_4190,N_4684);
nor U5641 (N_5641,N_4921,N_4143);
or U5642 (N_5642,N_4189,N_4524);
nand U5643 (N_5643,N_4146,N_4506);
nor U5644 (N_5644,N_4117,N_4284);
or U5645 (N_5645,N_4393,N_4907);
or U5646 (N_5646,N_4328,N_4560);
xnor U5647 (N_5647,N_4687,N_4805);
or U5648 (N_5648,N_4031,N_4352);
nand U5649 (N_5649,N_4588,N_4233);
nand U5650 (N_5650,N_4651,N_4510);
xnor U5651 (N_5651,N_4977,N_4456);
nor U5652 (N_5652,N_4283,N_4652);
nor U5653 (N_5653,N_4717,N_4079);
nand U5654 (N_5654,N_4103,N_4725);
or U5655 (N_5655,N_4084,N_4381);
or U5656 (N_5656,N_4275,N_4564);
nand U5657 (N_5657,N_4834,N_4429);
nor U5658 (N_5658,N_4342,N_4508);
or U5659 (N_5659,N_4694,N_4864);
xor U5660 (N_5660,N_4807,N_4212);
nor U5661 (N_5661,N_4961,N_4163);
or U5662 (N_5662,N_4055,N_4259);
nor U5663 (N_5663,N_4686,N_4636);
or U5664 (N_5664,N_4595,N_4517);
or U5665 (N_5665,N_4210,N_4897);
nand U5666 (N_5666,N_4465,N_4451);
nand U5667 (N_5667,N_4597,N_4939);
nor U5668 (N_5668,N_4606,N_4274);
and U5669 (N_5669,N_4600,N_4046);
nor U5670 (N_5670,N_4870,N_4248);
xor U5671 (N_5671,N_4843,N_4116);
and U5672 (N_5672,N_4319,N_4442);
nand U5673 (N_5673,N_4924,N_4269);
nor U5674 (N_5674,N_4062,N_4782);
xor U5675 (N_5675,N_4849,N_4955);
or U5676 (N_5676,N_4238,N_4491);
or U5677 (N_5677,N_4300,N_4855);
xor U5678 (N_5678,N_4309,N_4276);
or U5679 (N_5679,N_4571,N_4740);
nand U5680 (N_5680,N_4778,N_4806);
nor U5681 (N_5681,N_4433,N_4199);
nand U5682 (N_5682,N_4646,N_4175);
or U5683 (N_5683,N_4061,N_4350);
xnor U5684 (N_5684,N_4709,N_4267);
nand U5685 (N_5685,N_4525,N_4819);
or U5686 (N_5686,N_4811,N_4869);
or U5687 (N_5687,N_4281,N_4509);
and U5688 (N_5688,N_4747,N_4308);
nor U5689 (N_5689,N_4221,N_4614);
xnor U5690 (N_5690,N_4134,N_4695);
xor U5691 (N_5691,N_4675,N_4206);
or U5692 (N_5692,N_4724,N_4400);
or U5693 (N_5693,N_4834,N_4733);
nand U5694 (N_5694,N_4108,N_4573);
xnor U5695 (N_5695,N_4747,N_4550);
and U5696 (N_5696,N_4828,N_4737);
nand U5697 (N_5697,N_4700,N_4242);
nand U5698 (N_5698,N_4237,N_4583);
nor U5699 (N_5699,N_4103,N_4402);
xor U5700 (N_5700,N_4633,N_4623);
and U5701 (N_5701,N_4793,N_4485);
nand U5702 (N_5702,N_4432,N_4676);
and U5703 (N_5703,N_4992,N_4317);
or U5704 (N_5704,N_4384,N_4425);
nand U5705 (N_5705,N_4054,N_4148);
nand U5706 (N_5706,N_4263,N_4297);
nand U5707 (N_5707,N_4340,N_4641);
nor U5708 (N_5708,N_4510,N_4786);
nor U5709 (N_5709,N_4159,N_4859);
nand U5710 (N_5710,N_4952,N_4328);
nand U5711 (N_5711,N_4438,N_4296);
and U5712 (N_5712,N_4181,N_4754);
nand U5713 (N_5713,N_4392,N_4799);
nand U5714 (N_5714,N_4391,N_4216);
nand U5715 (N_5715,N_4282,N_4059);
and U5716 (N_5716,N_4593,N_4441);
or U5717 (N_5717,N_4198,N_4587);
nor U5718 (N_5718,N_4217,N_4891);
and U5719 (N_5719,N_4377,N_4751);
and U5720 (N_5720,N_4148,N_4335);
or U5721 (N_5721,N_4654,N_4606);
nor U5722 (N_5722,N_4941,N_4246);
or U5723 (N_5723,N_4309,N_4362);
nor U5724 (N_5724,N_4073,N_4819);
nor U5725 (N_5725,N_4782,N_4180);
or U5726 (N_5726,N_4762,N_4380);
and U5727 (N_5727,N_4629,N_4192);
and U5728 (N_5728,N_4068,N_4522);
and U5729 (N_5729,N_4346,N_4021);
nor U5730 (N_5730,N_4679,N_4426);
nand U5731 (N_5731,N_4283,N_4386);
nand U5732 (N_5732,N_4182,N_4141);
and U5733 (N_5733,N_4548,N_4563);
nand U5734 (N_5734,N_4584,N_4765);
xnor U5735 (N_5735,N_4007,N_4452);
nand U5736 (N_5736,N_4040,N_4085);
or U5737 (N_5737,N_4934,N_4859);
xor U5738 (N_5738,N_4595,N_4855);
nand U5739 (N_5739,N_4163,N_4686);
or U5740 (N_5740,N_4398,N_4332);
xnor U5741 (N_5741,N_4419,N_4900);
and U5742 (N_5742,N_4335,N_4620);
and U5743 (N_5743,N_4774,N_4137);
nor U5744 (N_5744,N_4080,N_4997);
nand U5745 (N_5745,N_4145,N_4701);
or U5746 (N_5746,N_4715,N_4739);
or U5747 (N_5747,N_4263,N_4132);
and U5748 (N_5748,N_4693,N_4538);
or U5749 (N_5749,N_4481,N_4095);
or U5750 (N_5750,N_4528,N_4323);
nand U5751 (N_5751,N_4897,N_4035);
xnor U5752 (N_5752,N_4410,N_4422);
nor U5753 (N_5753,N_4131,N_4712);
and U5754 (N_5754,N_4933,N_4213);
xnor U5755 (N_5755,N_4374,N_4423);
xnor U5756 (N_5756,N_4924,N_4371);
and U5757 (N_5757,N_4641,N_4410);
nor U5758 (N_5758,N_4252,N_4021);
and U5759 (N_5759,N_4066,N_4865);
nor U5760 (N_5760,N_4105,N_4626);
nand U5761 (N_5761,N_4790,N_4887);
xor U5762 (N_5762,N_4858,N_4921);
and U5763 (N_5763,N_4979,N_4252);
and U5764 (N_5764,N_4095,N_4501);
xor U5765 (N_5765,N_4034,N_4988);
or U5766 (N_5766,N_4524,N_4794);
or U5767 (N_5767,N_4514,N_4522);
nand U5768 (N_5768,N_4322,N_4344);
nand U5769 (N_5769,N_4431,N_4398);
nor U5770 (N_5770,N_4913,N_4495);
xor U5771 (N_5771,N_4855,N_4276);
or U5772 (N_5772,N_4109,N_4473);
nand U5773 (N_5773,N_4247,N_4173);
or U5774 (N_5774,N_4911,N_4536);
nor U5775 (N_5775,N_4638,N_4108);
xor U5776 (N_5776,N_4386,N_4511);
nand U5777 (N_5777,N_4305,N_4218);
nand U5778 (N_5778,N_4387,N_4898);
or U5779 (N_5779,N_4467,N_4560);
and U5780 (N_5780,N_4799,N_4534);
and U5781 (N_5781,N_4477,N_4727);
and U5782 (N_5782,N_4153,N_4540);
or U5783 (N_5783,N_4465,N_4990);
nor U5784 (N_5784,N_4515,N_4084);
nor U5785 (N_5785,N_4710,N_4653);
nand U5786 (N_5786,N_4255,N_4266);
and U5787 (N_5787,N_4157,N_4816);
and U5788 (N_5788,N_4592,N_4996);
nor U5789 (N_5789,N_4348,N_4806);
and U5790 (N_5790,N_4169,N_4990);
or U5791 (N_5791,N_4648,N_4828);
nand U5792 (N_5792,N_4663,N_4854);
nand U5793 (N_5793,N_4375,N_4193);
nor U5794 (N_5794,N_4275,N_4375);
and U5795 (N_5795,N_4845,N_4203);
or U5796 (N_5796,N_4439,N_4336);
nor U5797 (N_5797,N_4722,N_4004);
xor U5798 (N_5798,N_4864,N_4618);
xnor U5799 (N_5799,N_4797,N_4247);
xnor U5800 (N_5800,N_4235,N_4784);
nor U5801 (N_5801,N_4583,N_4178);
or U5802 (N_5802,N_4591,N_4335);
and U5803 (N_5803,N_4049,N_4666);
nand U5804 (N_5804,N_4017,N_4000);
or U5805 (N_5805,N_4604,N_4970);
and U5806 (N_5806,N_4887,N_4059);
xor U5807 (N_5807,N_4959,N_4471);
xnor U5808 (N_5808,N_4290,N_4540);
or U5809 (N_5809,N_4601,N_4935);
nor U5810 (N_5810,N_4172,N_4026);
xnor U5811 (N_5811,N_4684,N_4647);
or U5812 (N_5812,N_4038,N_4036);
nand U5813 (N_5813,N_4334,N_4739);
nor U5814 (N_5814,N_4867,N_4749);
and U5815 (N_5815,N_4833,N_4735);
nand U5816 (N_5816,N_4678,N_4563);
xnor U5817 (N_5817,N_4113,N_4913);
or U5818 (N_5818,N_4964,N_4617);
or U5819 (N_5819,N_4543,N_4816);
nand U5820 (N_5820,N_4513,N_4827);
and U5821 (N_5821,N_4347,N_4390);
nor U5822 (N_5822,N_4073,N_4463);
nor U5823 (N_5823,N_4429,N_4197);
or U5824 (N_5824,N_4381,N_4749);
or U5825 (N_5825,N_4067,N_4875);
nand U5826 (N_5826,N_4956,N_4062);
or U5827 (N_5827,N_4969,N_4962);
or U5828 (N_5828,N_4810,N_4025);
nand U5829 (N_5829,N_4492,N_4658);
nor U5830 (N_5830,N_4264,N_4002);
or U5831 (N_5831,N_4559,N_4632);
and U5832 (N_5832,N_4613,N_4633);
or U5833 (N_5833,N_4892,N_4390);
or U5834 (N_5834,N_4292,N_4392);
and U5835 (N_5835,N_4654,N_4664);
and U5836 (N_5836,N_4410,N_4253);
or U5837 (N_5837,N_4702,N_4793);
nand U5838 (N_5838,N_4466,N_4740);
nor U5839 (N_5839,N_4976,N_4771);
or U5840 (N_5840,N_4185,N_4398);
nand U5841 (N_5841,N_4763,N_4474);
xnor U5842 (N_5842,N_4697,N_4917);
nand U5843 (N_5843,N_4136,N_4573);
nand U5844 (N_5844,N_4862,N_4342);
and U5845 (N_5845,N_4071,N_4551);
xnor U5846 (N_5846,N_4820,N_4471);
and U5847 (N_5847,N_4049,N_4993);
and U5848 (N_5848,N_4301,N_4043);
nand U5849 (N_5849,N_4777,N_4457);
nor U5850 (N_5850,N_4485,N_4959);
or U5851 (N_5851,N_4672,N_4577);
or U5852 (N_5852,N_4086,N_4054);
nor U5853 (N_5853,N_4417,N_4747);
xor U5854 (N_5854,N_4623,N_4455);
or U5855 (N_5855,N_4004,N_4212);
nand U5856 (N_5856,N_4025,N_4450);
and U5857 (N_5857,N_4952,N_4048);
xnor U5858 (N_5858,N_4749,N_4684);
or U5859 (N_5859,N_4006,N_4919);
nor U5860 (N_5860,N_4274,N_4538);
xor U5861 (N_5861,N_4651,N_4310);
or U5862 (N_5862,N_4782,N_4226);
nor U5863 (N_5863,N_4469,N_4656);
and U5864 (N_5864,N_4720,N_4324);
xnor U5865 (N_5865,N_4409,N_4434);
nand U5866 (N_5866,N_4855,N_4957);
and U5867 (N_5867,N_4462,N_4453);
nand U5868 (N_5868,N_4724,N_4745);
xnor U5869 (N_5869,N_4163,N_4536);
and U5870 (N_5870,N_4583,N_4902);
nor U5871 (N_5871,N_4701,N_4345);
or U5872 (N_5872,N_4959,N_4894);
and U5873 (N_5873,N_4100,N_4194);
and U5874 (N_5874,N_4749,N_4571);
xnor U5875 (N_5875,N_4281,N_4903);
nor U5876 (N_5876,N_4188,N_4040);
nand U5877 (N_5877,N_4078,N_4142);
xnor U5878 (N_5878,N_4983,N_4432);
xor U5879 (N_5879,N_4562,N_4573);
and U5880 (N_5880,N_4696,N_4536);
nand U5881 (N_5881,N_4718,N_4498);
xnor U5882 (N_5882,N_4425,N_4641);
or U5883 (N_5883,N_4557,N_4520);
nor U5884 (N_5884,N_4035,N_4154);
xnor U5885 (N_5885,N_4771,N_4895);
or U5886 (N_5886,N_4594,N_4075);
nor U5887 (N_5887,N_4784,N_4225);
and U5888 (N_5888,N_4721,N_4436);
nor U5889 (N_5889,N_4334,N_4465);
nor U5890 (N_5890,N_4911,N_4825);
nor U5891 (N_5891,N_4888,N_4940);
or U5892 (N_5892,N_4472,N_4247);
nand U5893 (N_5893,N_4422,N_4131);
and U5894 (N_5894,N_4887,N_4783);
nor U5895 (N_5895,N_4273,N_4052);
xor U5896 (N_5896,N_4002,N_4079);
or U5897 (N_5897,N_4233,N_4234);
and U5898 (N_5898,N_4266,N_4730);
nor U5899 (N_5899,N_4301,N_4271);
and U5900 (N_5900,N_4405,N_4672);
nor U5901 (N_5901,N_4691,N_4435);
nand U5902 (N_5902,N_4266,N_4269);
nor U5903 (N_5903,N_4473,N_4991);
and U5904 (N_5904,N_4414,N_4531);
nand U5905 (N_5905,N_4532,N_4318);
or U5906 (N_5906,N_4033,N_4362);
xnor U5907 (N_5907,N_4936,N_4233);
and U5908 (N_5908,N_4110,N_4657);
and U5909 (N_5909,N_4393,N_4976);
xnor U5910 (N_5910,N_4170,N_4156);
nand U5911 (N_5911,N_4322,N_4250);
and U5912 (N_5912,N_4103,N_4732);
nor U5913 (N_5913,N_4951,N_4554);
xnor U5914 (N_5914,N_4683,N_4163);
nor U5915 (N_5915,N_4857,N_4233);
or U5916 (N_5916,N_4121,N_4980);
or U5917 (N_5917,N_4235,N_4935);
xnor U5918 (N_5918,N_4965,N_4478);
nor U5919 (N_5919,N_4781,N_4387);
nand U5920 (N_5920,N_4585,N_4996);
xnor U5921 (N_5921,N_4013,N_4204);
nand U5922 (N_5922,N_4567,N_4192);
or U5923 (N_5923,N_4022,N_4176);
nand U5924 (N_5924,N_4037,N_4027);
xnor U5925 (N_5925,N_4147,N_4591);
or U5926 (N_5926,N_4101,N_4602);
nand U5927 (N_5927,N_4542,N_4270);
and U5928 (N_5928,N_4299,N_4720);
xor U5929 (N_5929,N_4479,N_4169);
xor U5930 (N_5930,N_4053,N_4987);
nand U5931 (N_5931,N_4011,N_4394);
or U5932 (N_5932,N_4624,N_4664);
xnor U5933 (N_5933,N_4950,N_4733);
or U5934 (N_5934,N_4746,N_4960);
or U5935 (N_5935,N_4109,N_4460);
nand U5936 (N_5936,N_4122,N_4802);
xor U5937 (N_5937,N_4632,N_4884);
or U5938 (N_5938,N_4372,N_4802);
and U5939 (N_5939,N_4864,N_4405);
or U5940 (N_5940,N_4980,N_4965);
xor U5941 (N_5941,N_4143,N_4888);
xor U5942 (N_5942,N_4105,N_4694);
nor U5943 (N_5943,N_4708,N_4990);
nor U5944 (N_5944,N_4667,N_4893);
nor U5945 (N_5945,N_4503,N_4864);
and U5946 (N_5946,N_4741,N_4124);
xnor U5947 (N_5947,N_4138,N_4317);
nand U5948 (N_5948,N_4656,N_4204);
xnor U5949 (N_5949,N_4510,N_4395);
or U5950 (N_5950,N_4520,N_4749);
nor U5951 (N_5951,N_4704,N_4770);
and U5952 (N_5952,N_4106,N_4440);
and U5953 (N_5953,N_4992,N_4312);
nand U5954 (N_5954,N_4175,N_4757);
or U5955 (N_5955,N_4542,N_4971);
and U5956 (N_5956,N_4334,N_4563);
nor U5957 (N_5957,N_4762,N_4389);
nand U5958 (N_5958,N_4899,N_4524);
xnor U5959 (N_5959,N_4050,N_4257);
xor U5960 (N_5960,N_4342,N_4386);
or U5961 (N_5961,N_4164,N_4845);
or U5962 (N_5962,N_4091,N_4687);
nand U5963 (N_5963,N_4597,N_4382);
or U5964 (N_5964,N_4037,N_4542);
xor U5965 (N_5965,N_4816,N_4312);
xor U5966 (N_5966,N_4998,N_4245);
nor U5967 (N_5967,N_4295,N_4412);
nand U5968 (N_5968,N_4145,N_4497);
nor U5969 (N_5969,N_4061,N_4849);
nand U5970 (N_5970,N_4936,N_4940);
nor U5971 (N_5971,N_4697,N_4839);
nor U5972 (N_5972,N_4384,N_4703);
nor U5973 (N_5973,N_4953,N_4056);
and U5974 (N_5974,N_4714,N_4175);
or U5975 (N_5975,N_4889,N_4604);
and U5976 (N_5976,N_4522,N_4443);
or U5977 (N_5977,N_4647,N_4247);
and U5978 (N_5978,N_4307,N_4683);
nand U5979 (N_5979,N_4953,N_4971);
nand U5980 (N_5980,N_4394,N_4546);
or U5981 (N_5981,N_4068,N_4428);
xnor U5982 (N_5982,N_4791,N_4987);
nor U5983 (N_5983,N_4095,N_4258);
or U5984 (N_5984,N_4576,N_4253);
xnor U5985 (N_5985,N_4732,N_4583);
or U5986 (N_5986,N_4952,N_4679);
xnor U5987 (N_5987,N_4739,N_4993);
nand U5988 (N_5988,N_4936,N_4180);
nand U5989 (N_5989,N_4773,N_4551);
nand U5990 (N_5990,N_4468,N_4923);
and U5991 (N_5991,N_4659,N_4371);
nand U5992 (N_5992,N_4434,N_4822);
nor U5993 (N_5993,N_4994,N_4852);
and U5994 (N_5994,N_4412,N_4260);
nor U5995 (N_5995,N_4959,N_4098);
nor U5996 (N_5996,N_4457,N_4427);
nand U5997 (N_5997,N_4822,N_4209);
nor U5998 (N_5998,N_4205,N_4572);
and U5999 (N_5999,N_4146,N_4116);
nand U6000 (N_6000,N_5779,N_5701);
and U6001 (N_6001,N_5782,N_5274);
nor U6002 (N_6002,N_5875,N_5840);
nand U6003 (N_6003,N_5823,N_5648);
nand U6004 (N_6004,N_5477,N_5959);
nand U6005 (N_6005,N_5932,N_5075);
nand U6006 (N_6006,N_5235,N_5391);
xor U6007 (N_6007,N_5677,N_5272);
or U6008 (N_6008,N_5957,N_5880);
and U6009 (N_6009,N_5681,N_5127);
nand U6010 (N_6010,N_5461,N_5578);
or U6011 (N_6011,N_5383,N_5514);
nor U6012 (N_6012,N_5104,N_5700);
and U6013 (N_6013,N_5270,N_5397);
and U6014 (N_6014,N_5971,N_5451);
nand U6015 (N_6015,N_5663,N_5449);
and U6016 (N_6016,N_5828,N_5532);
nand U6017 (N_6017,N_5365,N_5122);
nand U6018 (N_6018,N_5258,N_5588);
xor U6019 (N_6019,N_5485,N_5721);
nor U6020 (N_6020,N_5496,N_5966);
and U6021 (N_6021,N_5610,N_5032);
and U6022 (N_6022,N_5209,N_5371);
and U6023 (N_6023,N_5605,N_5819);
and U6024 (N_6024,N_5878,N_5997);
xnor U6025 (N_6025,N_5557,N_5215);
nand U6026 (N_6026,N_5635,N_5482);
or U6027 (N_6027,N_5415,N_5232);
and U6028 (N_6028,N_5498,N_5084);
xnor U6029 (N_6029,N_5435,N_5945);
or U6030 (N_6030,N_5389,N_5969);
xor U6031 (N_6031,N_5034,N_5597);
nand U6032 (N_6032,N_5708,N_5968);
nand U6033 (N_6033,N_5749,N_5406);
nor U6034 (N_6034,N_5248,N_5191);
nor U6035 (N_6035,N_5128,N_5664);
nor U6036 (N_6036,N_5832,N_5695);
and U6037 (N_6037,N_5768,N_5506);
xnor U6038 (N_6038,N_5806,N_5714);
and U6039 (N_6039,N_5273,N_5647);
xor U6040 (N_6040,N_5107,N_5336);
or U6041 (N_6041,N_5289,N_5737);
nand U6042 (N_6042,N_5401,N_5702);
or U6043 (N_6043,N_5531,N_5847);
and U6044 (N_6044,N_5956,N_5527);
xnor U6045 (N_6045,N_5599,N_5261);
nand U6046 (N_6046,N_5329,N_5903);
and U6047 (N_6047,N_5891,N_5427);
nand U6048 (N_6048,N_5373,N_5432);
xor U6049 (N_6049,N_5207,N_5990);
nor U6050 (N_6050,N_5805,N_5355);
xor U6051 (N_6051,N_5291,N_5546);
nor U6052 (N_6052,N_5019,N_5511);
nor U6053 (N_6053,N_5279,N_5091);
nor U6054 (N_6054,N_5547,N_5707);
xnor U6055 (N_6055,N_5830,N_5214);
nand U6056 (N_6056,N_5103,N_5035);
xnor U6057 (N_6057,N_5755,N_5581);
or U6058 (N_6058,N_5484,N_5697);
nand U6059 (N_6059,N_5181,N_5739);
and U6060 (N_6060,N_5404,N_5410);
nor U6061 (N_6061,N_5295,N_5234);
or U6062 (N_6062,N_5278,N_5897);
nand U6063 (N_6063,N_5316,N_5481);
and U6064 (N_6064,N_5812,N_5226);
nand U6065 (N_6065,N_5748,N_5448);
and U6066 (N_6066,N_5740,N_5160);
nand U6067 (N_6067,N_5671,N_5572);
nor U6068 (N_6068,N_5333,N_5981);
nor U6069 (N_6069,N_5420,N_5256);
or U6070 (N_6070,N_5003,N_5871);
or U6071 (N_6071,N_5185,N_5146);
and U6072 (N_6072,N_5993,N_5650);
nand U6073 (N_6073,N_5447,N_5396);
and U6074 (N_6074,N_5044,N_5239);
xor U6075 (N_6075,N_5352,N_5725);
and U6076 (N_6076,N_5587,N_5766);
or U6077 (N_6077,N_5179,N_5972);
nor U6078 (N_6078,N_5910,N_5607);
xnor U6079 (N_6079,N_5370,N_5281);
nand U6080 (N_6080,N_5935,N_5149);
nand U6081 (N_6081,N_5787,N_5536);
xor U6082 (N_6082,N_5901,N_5752);
xnor U6083 (N_6083,N_5203,N_5504);
xnor U6084 (N_6084,N_5023,N_5326);
xnor U6085 (N_6085,N_5985,N_5328);
and U6086 (N_6086,N_5624,N_5706);
and U6087 (N_6087,N_5783,N_5462);
nand U6088 (N_6088,N_5066,N_5907);
xnor U6089 (N_6089,N_5839,N_5723);
or U6090 (N_6090,N_5342,N_5954);
nor U6091 (N_6091,N_5201,N_5573);
and U6092 (N_6092,N_5369,N_5976);
nand U6093 (N_6093,N_5764,N_5940);
and U6094 (N_6094,N_5458,N_5117);
nand U6095 (N_6095,N_5387,N_5006);
xnor U6096 (N_6096,N_5444,N_5184);
or U6097 (N_6097,N_5612,N_5366);
and U6098 (N_6098,N_5998,N_5363);
xor U6099 (N_6099,N_5260,N_5595);
or U6100 (N_6100,N_5896,N_5924);
xor U6101 (N_6101,N_5808,N_5013);
xnor U6102 (N_6102,N_5139,N_5645);
or U6103 (N_6103,N_5865,N_5487);
nand U6104 (N_6104,N_5180,N_5322);
nand U6105 (N_6105,N_5223,N_5499);
and U6106 (N_6106,N_5175,N_5958);
nand U6107 (N_6107,N_5821,N_5960);
and U6108 (N_6108,N_5379,N_5727);
nand U6109 (N_6109,N_5095,N_5439);
nand U6110 (N_6110,N_5086,N_5872);
and U6111 (N_6111,N_5964,N_5257);
nor U6112 (N_6112,N_5822,N_5000);
and U6113 (N_6113,N_5978,N_5125);
nand U6114 (N_6114,N_5186,N_5815);
and U6115 (N_6115,N_5984,N_5790);
or U6116 (N_6116,N_5220,N_5989);
or U6117 (N_6117,N_5111,N_5227);
nand U6118 (N_6118,N_5705,N_5965);
and U6119 (N_6119,N_5918,N_5569);
nand U6120 (N_6120,N_5466,N_5539);
or U6121 (N_6121,N_5844,N_5360);
or U6122 (N_6122,N_5080,N_5187);
nor U6123 (N_6123,N_5742,N_5134);
nand U6124 (N_6124,N_5771,N_5726);
or U6125 (N_6125,N_5123,N_5249);
nor U6126 (N_6126,N_5516,N_5548);
xor U6127 (N_6127,N_5293,N_5618);
nor U6128 (N_6128,N_5744,N_5194);
xnor U6129 (N_6129,N_5105,N_5753);
nand U6130 (N_6130,N_5300,N_5320);
and U6131 (N_6131,N_5582,N_5251);
xor U6132 (N_6132,N_5108,N_5064);
and U6133 (N_6133,N_5154,N_5887);
nand U6134 (N_6134,N_5537,N_5133);
and U6135 (N_6135,N_5094,N_5362);
or U6136 (N_6136,N_5649,N_5407);
nor U6137 (N_6137,N_5070,N_5102);
nor U6138 (N_6138,N_5277,N_5090);
or U6139 (N_6139,N_5565,N_5497);
xnor U6140 (N_6140,N_5789,N_5062);
or U6141 (N_6141,N_5561,N_5245);
or U6142 (N_6142,N_5926,N_5294);
xnor U6143 (N_6143,N_5970,N_5265);
nor U6144 (N_6144,N_5793,N_5076);
xor U6145 (N_6145,N_5949,N_5719);
nor U6146 (N_6146,N_5413,N_5393);
xor U6147 (N_6147,N_5563,N_5315);
and U6148 (N_6148,N_5746,N_5361);
and U6149 (N_6149,N_5987,N_5049);
nand U6150 (N_6150,N_5522,N_5130);
or U6151 (N_6151,N_5040,N_5479);
xnor U6152 (N_6152,N_5282,N_5304);
nand U6153 (N_6153,N_5164,N_5343);
nand U6154 (N_6154,N_5729,N_5325);
or U6155 (N_6155,N_5350,N_5698);
nor U6156 (N_6156,N_5512,N_5905);
or U6157 (N_6157,N_5859,N_5858);
and U6158 (N_6158,N_5577,N_5335);
nor U6159 (N_6159,N_5218,N_5120);
nor U6160 (N_6160,N_5135,N_5252);
or U6161 (N_6161,N_5598,N_5955);
or U6162 (N_6162,N_5622,N_5794);
nor U6163 (N_6163,N_5067,N_5033);
nor U6164 (N_6164,N_5047,N_5613);
xnor U6165 (N_6165,N_5637,N_5703);
nor U6166 (N_6166,N_5301,N_5381);
and U6167 (N_6167,N_5921,N_5367);
nor U6168 (N_6168,N_5640,N_5895);
and U6169 (N_6169,N_5491,N_5051);
xor U6170 (N_6170,N_5132,N_5089);
and U6171 (N_6171,N_5583,N_5240);
xor U6172 (N_6172,N_5165,N_5099);
nand U6173 (N_6173,N_5809,N_5161);
and U6174 (N_6174,N_5018,N_5724);
or U6175 (N_6175,N_5081,N_5619);
xor U6176 (N_6176,N_5318,N_5623);
nand U6177 (N_6177,N_5069,N_5082);
xor U6178 (N_6178,N_5585,N_5824);
nand U6179 (N_6179,N_5029,N_5473);
nand U6180 (N_6180,N_5621,N_5911);
xor U6181 (N_6181,N_5509,N_5306);
nor U6182 (N_6182,N_5378,N_5026);
and U6183 (N_6183,N_5217,N_5776);
xor U6184 (N_6184,N_5741,N_5684);
nor U6185 (N_6185,N_5596,N_5225);
and U6186 (N_6186,N_5673,N_5314);
xor U6187 (N_6187,N_5906,N_5110);
nand U6188 (N_6188,N_5429,N_5941);
or U6189 (N_6189,N_5097,N_5797);
or U6190 (N_6190,N_5192,N_5112);
or U6191 (N_6191,N_5486,N_5653);
and U6192 (N_6192,N_5348,N_5382);
nor U6193 (N_6193,N_5093,N_5733);
nand U6194 (N_6194,N_5087,N_5060);
nand U6195 (N_6195,N_5422,N_5309);
nor U6196 (N_6196,N_5254,N_5303);
nand U6197 (N_6197,N_5762,N_5178);
nand U6198 (N_6198,N_5399,N_5686);
xor U6199 (N_6199,N_5894,N_5559);
xor U6200 (N_6200,N_5608,N_5529);
and U6201 (N_6201,N_5041,N_5781);
nor U6202 (N_6202,N_5364,N_5551);
nand U6203 (N_6203,N_5627,N_5826);
xnor U6204 (N_6204,N_5501,N_5045);
nand U6205 (N_6205,N_5507,N_5230);
or U6206 (N_6206,N_5408,N_5025);
xor U6207 (N_6207,N_5827,N_5508);
and U6208 (N_6208,N_5210,N_5963);
nor U6209 (N_6209,N_5961,N_5224);
and U6210 (N_6210,N_5324,N_5228);
nor U6211 (N_6211,N_5813,N_5208);
or U6212 (N_6212,N_5944,N_5475);
nand U6213 (N_6213,N_5153,N_5525);
and U6214 (N_6214,N_5667,N_5377);
nand U6215 (N_6215,N_5829,N_5109);
xnor U6216 (N_6216,N_5158,N_5057);
nand U6217 (N_6217,N_5151,N_5403);
xor U6218 (N_6218,N_5678,N_5390);
xor U6219 (N_6219,N_5680,N_5005);
and U6220 (N_6220,N_5053,N_5953);
and U6221 (N_6221,N_5331,N_5713);
and U6222 (N_6222,N_5709,N_5480);
xnor U6223 (N_6223,N_5116,N_5943);
xor U6224 (N_6224,N_5777,N_5975);
or U6225 (N_6225,N_5031,N_5734);
xnor U6226 (N_6226,N_5020,N_5835);
xor U6227 (N_6227,N_5211,N_5884);
xor U6228 (N_6228,N_5155,N_5216);
nor U6229 (N_6229,N_5298,N_5290);
and U6230 (N_6230,N_5834,N_5384);
or U6231 (N_6231,N_5433,N_5515);
nand U6232 (N_6232,N_5747,N_5873);
nand U6233 (N_6233,N_5716,N_5357);
nand U6234 (N_6234,N_5933,N_5974);
and U6235 (N_6235,N_5919,N_5242);
nand U6236 (N_6236,N_5927,N_5063);
xor U6237 (N_6237,N_5756,N_5874);
nand U6238 (N_6238,N_5068,N_5675);
or U6239 (N_6239,N_5562,N_5570);
and U6240 (N_6240,N_5693,N_5876);
nor U6241 (N_6241,N_5398,N_5411);
nor U6242 (N_6242,N_5544,N_5048);
and U6243 (N_6243,N_5517,N_5995);
nor U6244 (N_6244,N_5296,N_5061);
and U6245 (N_6245,N_5323,N_5478);
xnor U6246 (N_6246,N_5140,N_5205);
or U6247 (N_6247,N_5474,N_5869);
nand U6248 (N_6248,N_5579,N_5758);
and U6249 (N_6249,N_5131,N_5098);
and U6250 (N_6250,N_5732,N_5540);
nor U6251 (N_6251,N_5615,N_5784);
nor U6252 (N_6252,N_5330,N_5172);
nor U6253 (N_6253,N_5440,N_5785);
xnor U6254 (N_6254,N_5977,N_5358);
xor U6255 (N_6255,N_5213,N_5002);
nand U6256 (N_6256,N_5030,N_5386);
nand U6257 (N_6257,N_5520,N_5244);
or U6258 (N_6258,N_5145,N_5024);
xor U6259 (N_6259,N_5879,N_5631);
xor U6260 (N_6260,N_5688,N_5503);
and U6261 (N_6261,N_5850,N_5077);
nor U6262 (N_6262,N_5419,N_5881);
and U6263 (N_6263,N_5246,N_5780);
and U6264 (N_6264,N_5021,N_5126);
nand U6265 (N_6265,N_5564,N_5890);
nand U6266 (N_6266,N_5803,N_5124);
xor U6267 (N_6267,N_5027,N_5791);
and U6268 (N_6268,N_5908,N_5524);
xnor U6269 (N_6269,N_5247,N_5982);
and U6270 (N_6270,N_5168,N_5374);
xor U6271 (N_6271,N_5825,N_5354);
nor U6272 (N_6272,N_5037,N_5351);
xnor U6273 (N_6273,N_5302,N_5804);
nor U6274 (N_6274,N_5575,N_5696);
nand U6275 (N_6275,N_5848,N_5345);
and U6276 (N_6276,N_5778,N_5883);
xor U6277 (N_6277,N_5425,N_5483);
xor U6278 (N_6278,N_5630,N_5672);
or U6279 (N_6279,N_5936,N_5255);
and U6280 (N_6280,N_5886,N_5450);
or U6281 (N_6281,N_5772,N_5065);
nand U6282 (N_6282,N_5909,N_5666);
or U6283 (N_6283,N_5414,N_5321);
xnor U6284 (N_6284,N_5861,N_5639);
and U6285 (N_6285,N_5556,N_5584);
and U6286 (N_6286,N_5923,N_5202);
nor U6287 (N_6287,N_5690,N_5728);
nor U6288 (N_6288,N_5088,N_5129);
nand U6289 (N_6289,N_5549,N_5676);
nor U6290 (N_6290,N_5510,N_5014);
nor U6291 (N_6291,N_5231,N_5052);
xnor U6292 (N_6292,N_5900,N_5799);
xor U6293 (N_6293,N_5428,N_5297);
and U6294 (N_6294,N_5204,N_5200);
nor U6295 (N_6295,N_5400,N_5939);
and U6296 (N_6296,N_5632,N_5773);
or U6297 (N_6297,N_5173,N_5455);
and U6298 (N_6298,N_5453,N_5288);
nand U6299 (N_6299,N_5502,N_5530);
or U6300 (N_6300,N_5817,N_5337);
nor U6301 (N_6301,N_5533,N_5616);
nand U6302 (N_6302,N_5851,N_5054);
xnor U6303 (N_6303,N_5913,N_5885);
and U6304 (N_6304,N_5931,N_5920);
nor U6305 (N_6305,N_5016,N_5807);
nand U6306 (N_6306,N_5317,N_5558);
nor U6307 (N_6307,N_5849,N_5658);
xor U6308 (N_6308,N_5442,N_5948);
and U6309 (N_6309,N_5385,N_5937);
nand U6310 (N_6310,N_5182,N_5001);
nor U6311 (N_6311,N_5628,N_5250);
and U6312 (N_6312,N_5687,N_5567);
and U6313 (N_6313,N_5898,N_5763);
or U6314 (N_6314,N_5346,N_5356);
and U6315 (N_6315,N_5864,N_5388);
and U6316 (N_6316,N_5668,N_5115);
nand U6317 (N_6317,N_5183,N_5611);
nand U6318 (N_6318,N_5136,N_5083);
nand U6319 (N_6319,N_5468,N_5718);
nand U6320 (N_6320,N_5991,N_5162);
nor U6321 (N_6321,N_5198,N_5892);
or U6322 (N_6322,N_5163,N_5229);
nand U6323 (N_6323,N_5142,N_5012);
xor U6324 (N_6324,N_5545,N_5096);
xor U6325 (N_6325,N_5902,N_5602);
nand U6326 (N_6326,N_5757,N_5170);
xnor U6327 (N_6327,N_5877,N_5452);
nand U6328 (N_6328,N_5854,N_5056);
nor U6329 (N_6329,N_5603,N_5917);
nor U6330 (N_6330,N_5994,N_5731);
xor U6331 (N_6331,N_5816,N_5138);
nand U6332 (N_6332,N_5190,N_5011);
nor U6333 (N_6333,N_5712,N_5662);
nor U6334 (N_6334,N_5661,N_5008);
xor U6335 (N_6335,N_5767,N_5863);
nand U6336 (N_6336,N_5340,N_5625);
xnor U6337 (N_6337,N_5405,N_5464);
and U6338 (N_6338,N_5592,N_5169);
and U6339 (N_6339,N_5685,N_5143);
or U6340 (N_6340,N_5176,N_5691);
and U6341 (N_6341,N_5820,N_5617);
xor U6342 (N_6342,N_5079,N_5078);
or U6343 (N_6343,N_5836,N_5541);
or U6344 (N_6344,N_5553,N_5802);
or U6345 (N_6345,N_5465,N_5262);
and U6346 (N_6346,N_5119,N_5456);
nor U6347 (N_6347,N_5243,N_5928);
or U6348 (N_6348,N_5426,N_5795);
and U6349 (N_6349,N_5505,N_5730);
nor U6350 (N_6350,N_5534,N_5445);
nand U6351 (N_6351,N_5171,N_5188);
xnor U6352 (N_6352,N_5845,N_5574);
nand U6353 (N_6353,N_5470,N_5743);
nand U6354 (N_6354,N_5715,N_5528);
nand U6355 (N_6355,N_5983,N_5538);
and U6356 (N_6356,N_5962,N_5838);
nand U6357 (N_6357,N_5904,N_5308);
nor U6358 (N_6358,N_5638,N_5986);
and U6359 (N_6359,N_5652,N_5555);
xnor U6360 (N_6360,N_5866,N_5930);
or U6361 (N_6361,N_5152,N_5434);
and U6362 (N_6362,N_5853,N_5280);
xor U6363 (N_6363,N_5028,N_5810);
nand U6364 (N_6364,N_5349,N_5141);
xnor U6365 (N_6365,N_5999,N_5311);
xor U6366 (N_6366,N_5144,N_5967);
xnor U6367 (N_6367,N_5055,N_5438);
or U6368 (N_6368,N_5852,N_5568);
nand U6369 (N_6369,N_5237,N_5899);
nand U6370 (N_6370,N_5626,N_5704);
and U6371 (N_6371,N_5916,N_5513);
nor U6372 (N_6372,N_5471,N_5100);
and U6373 (N_6373,N_5299,N_5284);
and U6374 (N_6374,N_5518,N_5915);
or U6375 (N_6375,N_5980,N_5046);
nor U6376 (N_6376,N_5837,N_5285);
xor U6377 (N_6377,N_5368,N_5147);
or U6378 (N_6378,N_5492,N_5979);
and U6379 (N_6379,N_5436,N_5275);
nand U6380 (N_6380,N_5846,N_5039);
nor U6381 (N_6381,N_5754,N_5167);
xnor U6382 (N_6382,N_5058,N_5380);
and U6383 (N_6383,N_5629,N_5253);
nor U6384 (N_6384,N_5009,N_5775);
and U6385 (N_6385,N_5593,N_5268);
and U6386 (N_6386,N_5292,N_5694);
and U6387 (N_6387,N_5341,N_5437);
nor U6388 (N_6388,N_5774,N_5893);
or U6389 (N_6389,N_5973,N_5798);
xor U6390 (N_6390,N_5106,N_5269);
or U6391 (N_6391,N_5118,N_5860);
xnor U6392 (N_6392,N_5566,N_5038);
nor U6393 (N_6393,N_5736,N_5500);
nor U6394 (N_6394,N_5017,N_5811);
nor U6395 (N_6395,N_5988,N_5085);
nand U6396 (N_6396,N_5488,N_5922);
or U6397 (N_6397,N_5590,N_5022);
and U6398 (N_6398,N_5494,N_5460);
or U6399 (N_6399,N_5344,N_5870);
nor U6400 (N_6400,N_5007,N_5651);
nand U6401 (N_6401,N_5431,N_5818);
nand U6402 (N_6402,N_5889,N_5770);
and U6403 (N_6403,N_5942,N_5489);
nand U6404 (N_6404,N_5594,N_5454);
nand U6405 (N_6405,N_5843,N_5659);
or U6406 (N_6406,N_5042,N_5267);
xor U6407 (N_6407,N_5313,N_5283);
nand U6408 (N_6408,N_5868,N_5786);
nand U6409 (N_6409,N_5327,N_5157);
nor U6410 (N_6410,N_5761,N_5660);
nand U6411 (N_6411,N_5833,N_5073);
nand U6412 (N_6412,N_5550,N_5472);
nor U6413 (N_6413,N_5862,N_5219);
and U6414 (N_6414,N_5189,N_5699);
nand U6415 (N_6415,N_5526,N_5166);
or U6416 (N_6416,N_5856,N_5855);
xnor U6417 (N_6417,N_5586,N_5751);
and U6418 (N_6418,N_5416,N_5769);
nor U6419 (N_6419,N_5121,N_5004);
or U6420 (N_6420,N_5286,N_5159);
nor U6421 (N_6421,N_5043,N_5319);
or U6422 (N_6422,N_5476,N_5882);
or U6423 (N_6423,N_5842,N_5347);
nor U6424 (N_6424,N_5552,N_5402);
nor U6425 (N_6425,N_5375,N_5417);
xnor U6426 (N_6426,N_5457,N_5222);
xor U6427 (N_6427,N_5951,N_5796);
nor U6428 (N_6428,N_5925,N_5424);
or U6429 (N_6429,N_5950,N_5888);
nor U6430 (N_6430,N_5654,N_5212);
nor U6431 (N_6431,N_5236,N_5670);
nor U6432 (N_6432,N_5199,N_5992);
xor U6433 (N_6433,N_5646,N_5312);
nand U6434 (N_6434,N_5711,N_5679);
or U6435 (N_6435,N_5519,N_5841);
or U6436 (N_6436,N_5929,N_5745);
nor U6437 (N_6437,N_5765,N_5412);
or U6438 (N_6438,N_5722,N_5010);
or U6439 (N_6439,N_5376,N_5441);
nor U6440 (N_6440,N_5113,N_5946);
or U6441 (N_6441,N_5600,N_5554);
nor U6442 (N_6442,N_5177,N_5287);
nor U6443 (N_6443,N_5469,N_5193);
xor U6444 (N_6444,N_5601,N_5036);
and U6445 (N_6445,N_5339,N_5542);
nor U6446 (N_6446,N_5307,N_5353);
and U6447 (N_6447,N_5535,N_5392);
nand U6448 (N_6448,N_5644,N_5792);
nor U6449 (N_6449,N_5634,N_5359);
or U6450 (N_6450,N_5137,N_5669);
or U6451 (N_6451,N_5443,N_5683);
nand U6452 (N_6452,N_5614,N_5710);
nor U6453 (N_6453,N_5760,N_5050);
and U6454 (N_6454,N_5310,N_5642);
or U6455 (N_6455,N_5015,N_5523);
nor U6456 (N_6456,N_5521,N_5276);
xnor U6457 (N_6457,N_5657,N_5241);
xor U6458 (N_6458,N_5338,N_5150);
xnor U6459 (N_6459,N_5759,N_5446);
or U6460 (N_6460,N_5071,N_5156);
xnor U6461 (N_6461,N_5334,N_5238);
xnor U6462 (N_6462,N_5750,N_5857);
nand U6463 (N_6463,N_5233,N_5266);
nand U6464 (N_6464,N_5682,N_5800);
nor U6465 (N_6465,N_5259,N_5490);
or U6466 (N_6466,N_5589,N_5571);
and U6467 (N_6467,N_5655,N_5264);
or U6468 (N_6468,N_5914,N_5463);
or U6469 (N_6469,N_5395,N_5665);
and U6470 (N_6470,N_5735,N_5114);
xnor U6471 (N_6471,N_5206,N_5195);
nand U6472 (N_6472,N_5196,N_5717);
or U6473 (N_6473,N_5305,N_5423);
or U6474 (N_6474,N_5606,N_5467);
xnor U6475 (N_6475,N_5609,N_5421);
nand U6476 (N_6476,N_5372,N_5934);
and U6477 (N_6477,N_5689,N_5148);
nand U6478 (N_6478,N_5072,N_5459);
or U6479 (N_6479,N_5604,N_5720);
nand U6480 (N_6480,N_5263,N_5656);
nor U6481 (N_6481,N_5801,N_5788);
nor U6482 (N_6482,N_5938,N_5738);
nor U6483 (N_6483,N_5636,N_5394);
or U6484 (N_6484,N_5641,N_5409);
or U6485 (N_6485,N_5620,N_5543);
xnor U6486 (N_6486,N_5633,N_5947);
nand U6487 (N_6487,N_5418,N_5271);
nand U6488 (N_6488,N_5643,N_5174);
or U6489 (N_6489,N_5332,N_5867);
nor U6490 (N_6490,N_5814,N_5074);
nand U6491 (N_6491,N_5674,N_5591);
nor U6492 (N_6492,N_5580,N_5221);
nor U6493 (N_6493,N_5831,N_5912);
and U6494 (N_6494,N_5996,N_5430);
xor U6495 (N_6495,N_5576,N_5560);
nand U6496 (N_6496,N_5692,N_5952);
nand U6497 (N_6497,N_5197,N_5493);
nor U6498 (N_6498,N_5092,N_5495);
and U6499 (N_6499,N_5059,N_5101);
or U6500 (N_6500,N_5115,N_5906);
xnor U6501 (N_6501,N_5530,N_5936);
nor U6502 (N_6502,N_5234,N_5402);
or U6503 (N_6503,N_5109,N_5341);
or U6504 (N_6504,N_5463,N_5930);
and U6505 (N_6505,N_5213,N_5129);
xnor U6506 (N_6506,N_5744,N_5219);
and U6507 (N_6507,N_5547,N_5766);
nand U6508 (N_6508,N_5163,N_5757);
or U6509 (N_6509,N_5543,N_5707);
xor U6510 (N_6510,N_5285,N_5818);
or U6511 (N_6511,N_5690,N_5568);
or U6512 (N_6512,N_5901,N_5707);
and U6513 (N_6513,N_5632,N_5888);
nand U6514 (N_6514,N_5301,N_5166);
xor U6515 (N_6515,N_5429,N_5361);
nor U6516 (N_6516,N_5862,N_5880);
nand U6517 (N_6517,N_5966,N_5248);
nand U6518 (N_6518,N_5396,N_5278);
xnor U6519 (N_6519,N_5624,N_5888);
and U6520 (N_6520,N_5617,N_5592);
or U6521 (N_6521,N_5466,N_5891);
and U6522 (N_6522,N_5934,N_5561);
and U6523 (N_6523,N_5811,N_5335);
nand U6524 (N_6524,N_5308,N_5344);
and U6525 (N_6525,N_5539,N_5135);
nand U6526 (N_6526,N_5806,N_5354);
nor U6527 (N_6527,N_5144,N_5499);
or U6528 (N_6528,N_5429,N_5116);
and U6529 (N_6529,N_5375,N_5517);
nand U6530 (N_6530,N_5382,N_5684);
or U6531 (N_6531,N_5694,N_5586);
nor U6532 (N_6532,N_5381,N_5336);
xnor U6533 (N_6533,N_5667,N_5354);
or U6534 (N_6534,N_5917,N_5444);
nor U6535 (N_6535,N_5519,N_5330);
xnor U6536 (N_6536,N_5019,N_5971);
and U6537 (N_6537,N_5823,N_5810);
xnor U6538 (N_6538,N_5947,N_5034);
and U6539 (N_6539,N_5359,N_5716);
or U6540 (N_6540,N_5935,N_5612);
xor U6541 (N_6541,N_5200,N_5146);
xnor U6542 (N_6542,N_5802,N_5042);
nand U6543 (N_6543,N_5112,N_5390);
nor U6544 (N_6544,N_5075,N_5441);
xnor U6545 (N_6545,N_5509,N_5609);
xnor U6546 (N_6546,N_5002,N_5308);
and U6547 (N_6547,N_5536,N_5948);
xor U6548 (N_6548,N_5946,N_5090);
nand U6549 (N_6549,N_5694,N_5101);
and U6550 (N_6550,N_5465,N_5580);
or U6551 (N_6551,N_5589,N_5679);
nor U6552 (N_6552,N_5104,N_5135);
nand U6553 (N_6553,N_5122,N_5439);
nor U6554 (N_6554,N_5454,N_5722);
xor U6555 (N_6555,N_5341,N_5495);
nand U6556 (N_6556,N_5914,N_5368);
and U6557 (N_6557,N_5799,N_5703);
and U6558 (N_6558,N_5106,N_5911);
xor U6559 (N_6559,N_5438,N_5563);
and U6560 (N_6560,N_5914,N_5230);
xnor U6561 (N_6561,N_5620,N_5165);
nand U6562 (N_6562,N_5671,N_5250);
or U6563 (N_6563,N_5264,N_5044);
xnor U6564 (N_6564,N_5485,N_5230);
xor U6565 (N_6565,N_5751,N_5935);
nor U6566 (N_6566,N_5411,N_5294);
or U6567 (N_6567,N_5994,N_5814);
and U6568 (N_6568,N_5283,N_5859);
and U6569 (N_6569,N_5627,N_5759);
xnor U6570 (N_6570,N_5051,N_5399);
or U6571 (N_6571,N_5930,N_5039);
and U6572 (N_6572,N_5350,N_5526);
nor U6573 (N_6573,N_5823,N_5150);
nor U6574 (N_6574,N_5307,N_5536);
nor U6575 (N_6575,N_5953,N_5096);
and U6576 (N_6576,N_5972,N_5680);
and U6577 (N_6577,N_5742,N_5582);
and U6578 (N_6578,N_5337,N_5175);
and U6579 (N_6579,N_5991,N_5124);
and U6580 (N_6580,N_5116,N_5903);
xnor U6581 (N_6581,N_5649,N_5705);
nor U6582 (N_6582,N_5576,N_5691);
nand U6583 (N_6583,N_5140,N_5525);
or U6584 (N_6584,N_5377,N_5872);
nor U6585 (N_6585,N_5001,N_5539);
xor U6586 (N_6586,N_5311,N_5379);
and U6587 (N_6587,N_5936,N_5178);
and U6588 (N_6588,N_5740,N_5289);
xor U6589 (N_6589,N_5679,N_5798);
nor U6590 (N_6590,N_5918,N_5496);
xor U6591 (N_6591,N_5207,N_5955);
nor U6592 (N_6592,N_5926,N_5226);
nand U6593 (N_6593,N_5453,N_5142);
or U6594 (N_6594,N_5857,N_5934);
xor U6595 (N_6595,N_5545,N_5263);
nor U6596 (N_6596,N_5919,N_5189);
xor U6597 (N_6597,N_5688,N_5761);
nand U6598 (N_6598,N_5690,N_5290);
and U6599 (N_6599,N_5917,N_5423);
nand U6600 (N_6600,N_5638,N_5084);
and U6601 (N_6601,N_5638,N_5777);
or U6602 (N_6602,N_5216,N_5265);
or U6603 (N_6603,N_5749,N_5904);
nor U6604 (N_6604,N_5372,N_5785);
or U6605 (N_6605,N_5254,N_5689);
nand U6606 (N_6606,N_5996,N_5618);
nor U6607 (N_6607,N_5874,N_5109);
xnor U6608 (N_6608,N_5886,N_5801);
xnor U6609 (N_6609,N_5329,N_5239);
nand U6610 (N_6610,N_5527,N_5723);
and U6611 (N_6611,N_5406,N_5331);
nand U6612 (N_6612,N_5077,N_5119);
xnor U6613 (N_6613,N_5920,N_5690);
and U6614 (N_6614,N_5059,N_5926);
nor U6615 (N_6615,N_5215,N_5535);
and U6616 (N_6616,N_5722,N_5230);
nand U6617 (N_6617,N_5572,N_5527);
or U6618 (N_6618,N_5044,N_5027);
nand U6619 (N_6619,N_5129,N_5893);
nor U6620 (N_6620,N_5961,N_5614);
xor U6621 (N_6621,N_5016,N_5338);
nand U6622 (N_6622,N_5099,N_5078);
nor U6623 (N_6623,N_5631,N_5682);
and U6624 (N_6624,N_5711,N_5420);
or U6625 (N_6625,N_5380,N_5081);
nand U6626 (N_6626,N_5064,N_5277);
nand U6627 (N_6627,N_5970,N_5909);
xnor U6628 (N_6628,N_5312,N_5255);
nor U6629 (N_6629,N_5341,N_5283);
or U6630 (N_6630,N_5030,N_5724);
and U6631 (N_6631,N_5158,N_5895);
xnor U6632 (N_6632,N_5310,N_5761);
nand U6633 (N_6633,N_5989,N_5750);
nand U6634 (N_6634,N_5122,N_5216);
nor U6635 (N_6635,N_5929,N_5167);
nor U6636 (N_6636,N_5747,N_5374);
or U6637 (N_6637,N_5852,N_5239);
xnor U6638 (N_6638,N_5897,N_5289);
and U6639 (N_6639,N_5517,N_5979);
nand U6640 (N_6640,N_5509,N_5571);
nand U6641 (N_6641,N_5414,N_5065);
and U6642 (N_6642,N_5433,N_5125);
nor U6643 (N_6643,N_5614,N_5933);
nand U6644 (N_6644,N_5351,N_5935);
or U6645 (N_6645,N_5136,N_5151);
xor U6646 (N_6646,N_5549,N_5475);
nand U6647 (N_6647,N_5287,N_5409);
xnor U6648 (N_6648,N_5734,N_5810);
nor U6649 (N_6649,N_5674,N_5814);
and U6650 (N_6650,N_5410,N_5511);
and U6651 (N_6651,N_5653,N_5286);
nand U6652 (N_6652,N_5437,N_5039);
nand U6653 (N_6653,N_5675,N_5028);
or U6654 (N_6654,N_5047,N_5572);
and U6655 (N_6655,N_5923,N_5220);
and U6656 (N_6656,N_5818,N_5836);
and U6657 (N_6657,N_5318,N_5665);
nor U6658 (N_6658,N_5197,N_5273);
and U6659 (N_6659,N_5157,N_5045);
nand U6660 (N_6660,N_5801,N_5338);
nand U6661 (N_6661,N_5651,N_5674);
xnor U6662 (N_6662,N_5191,N_5008);
nor U6663 (N_6663,N_5494,N_5936);
nor U6664 (N_6664,N_5035,N_5633);
xnor U6665 (N_6665,N_5649,N_5867);
nand U6666 (N_6666,N_5711,N_5508);
and U6667 (N_6667,N_5851,N_5678);
nand U6668 (N_6668,N_5545,N_5615);
and U6669 (N_6669,N_5554,N_5217);
and U6670 (N_6670,N_5369,N_5351);
or U6671 (N_6671,N_5702,N_5613);
nand U6672 (N_6672,N_5620,N_5356);
xnor U6673 (N_6673,N_5039,N_5863);
xor U6674 (N_6674,N_5572,N_5714);
nor U6675 (N_6675,N_5476,N_5665);
xnor U6676 (N_6676,N_5608,N_5889);
and U6677 (N_6677,N_5628,N_5278);
nand U6678 (N_6678,N_5325,N_5334);
xnor U6679 (N_6679,N_5917,N_5548);
nor U6680 (N_6680,N_5205,N_5352);
or U6681 (N_6681,N_5452,N_5483);
nand U6682 (N_6682,N_5066,N_5021);
or U6683 (N_6683,N_5841,N_5935);
nor U6684 (N_6684,N_5424,N_5473);
xnor U6685 (N_6685,N_5095,N_5930);
and U6686 (N_6686,N_5430,N_5722);
and U6687 (N_6687,N_5840,N_5523);
nor U6688 (N_6688,N_5682,N_5339);
xor U6689 (N_6689,N_5531,N_5947);
xnor U6690 (N_6690,N_5230,N_5247);
and U6691 (N_6691,N_5459,N_5846);
nor U6692 (N_6692,N_5838,N_5958);
and U6693 (N_6693,N_5844,N_5953);
xor U6694 (N_6694,N_5194,N_5947);
nor U6695 (N_6695,N_5512,N_5068);
xor U6696 (N_6696,N_5668,N_5199);
or U6697 (N_6697,N_5986,N_5724);
nand U6698 (N_6698,N_5745,N_5001);
nor U6699 (N_6699,N_5264,N_5946);
xnor U6700 (N_6700,N_5144,N_5292);
or U6701 (N_6701,N_5995,N_5017);
nand U6702 (N_6702,N_5480,N_5528);
xnor U6703 (N_6703,N_5732,N_5822);
and U6704 (N_6704,N_5163,N_5559);
xnor U6705 (N_6705,N_5802,N_5407);
xnor U6706 (N_6706,N_5210,N_5390);
xor U6707 (N_6707,N_5110,N_5380);
and U6708 (N_6708,N_5012,N_5731);
and U6709 (N_6709,N_5206,N_5146);
and U6710 (N_6710,N_5186,N_5383);
nor U6711 (N_6711,N_5792,N_5860);
nor U6712 (N_6712,N_5556,N_5555);
nand U6713 (N_6713,N_5759,N_5925);
xor U6714 (N_6714,N_5077,N_5280);
or U6715 (N_6715,N_5264,N_5189);
or U6716 (N_6716,N_5277,N_5879);
nand U6717 (N_6717,N_5014,N_5546);
or U6718 (N_6718,N_5525,N_5364);
or U6719 (N_6719,N_5769,N_5797);
xor U6720 (N_6720,N_5671,N_5847);
or U6721 (N_6721,N_5387,N_5257);
nand U6722 (N_6722,N_5158,N_5583);
nand U6723 (N_6723,N_5217,N_5699);
nor U6724 (N_6724,N_5949,N_5871);
and U6725 (N_6725,N_5310,N_5182);
or U6726 (N_6726,N_5750,N_5362);
or U6727 (N_6727,N_5720,N_5265);
nand U6728 (N_6728,N_5162,N_5993);
nor U6729 (N_6729,N_5972,N_5472);
nor U6730 (N_6730,N_5500,N_5425);
and U6731 (N_6731,N_5521,N_5045);
and U6732 (N_6732,N_5668,N_5070);
xnor U6733 (N_6733,N_5016,N_5330);
xnor U6734 (N_6734,N_5449,N_5439);
nor U6735 (N_6735,N_5722,N_5439);
and U6736 (N_6736,N_5077,N_5195);
or U6737 (N_6737,N_5709,N_5860);
nor U6738 (N_6738,N_5290,N_5007);
nand U6739 (N_6739,N_5661,N_5243);
xor U6740 (N_6740,N_5871,N_5620);
nand U6741 (N_6741,N_5913,N_5467);
or U6742 (N_6742,N_5198,N_5919);
or U6743 (N_6743,N_5619,N_5476);
xnor U6744 (N_6744,N_5795,N_5485);
nand U6745 (N_6745,N_5374,N_5198);
and U6746 (N_6746,N_5223,N_5274);
xor U6747 (N_6747,N_5241,N_5635);
nand U6748 (N_6748,N_5402,N_5584);
xnor U6749 (N_6749,N_5847,N_5788);
or U6750 (N_6750,N_5401,N_5591);
nor U6751 (N_6751,N_5600,N_5055);
nand U6752 (N_6752,N_5000,N_5977);
and U6753 (N_6753,N_5053,N_5285);
nand U6754 (N_6754,N_5255,N_5948);
nor U6755 (N_6755,N_5427,N_5746);
nor U6756 (N_6756,N_5311,N_5733);
or U6757 (N_6757,N_5685,N_5655);
and U6758 (N_6758,N_5315,N_5360);
or U6759 (N_6759,N_5438,N_5761);
nand U6760 (N_6760,N_5261,N_5966);
and U6761 (N_6761,N_5663,N_5617);
nor U6762 (N_6762,N_5423,N_5539);
xor U6763 (N_6763,N_5849,N_5521);
or U6764 (N_6764,N_5779,N_5223);
xor U6765 (N_6765,N_5829,N_5857);
nor U6766 (N_6766,N_5085,N_5577);
xor U6767 (N_6767,N_5146,N_5051);
nand U6768 (N_6768,N_5128,N_5057);
and U6769 (N_6769,N_5519,N_5591);
nand U6770 (N_6770,N_5127,N_5753);
or U6771 (N_6771,N_5642,N_5359);
and U6772 (N_6772,N_5318,N_5228);
and U6773 (N_6773,N_5582,N_5157);
and U6774 (N_6774,N_5475,N_5745);
or U6775 (N_6775,N_5640,N_5490);
or U6776 (N_6776,N_5776,N_5758);
nor U6777 (N_6777,N_5558,N_5243);
nor U6778 (N_6778,N_5948,N_5285);
xnor U6779 (N_6779,N_5250,N_5062);
nor U6780 (N_6780,N_5753,N_5952);
nor U6781 (N_6781,N_5930,N_5499);
nor U6782 (N_6782,N_5737,N_5306);
or U6783 (N_6783,N_5220,N_5901);
or U6784 (N_6784,N_5696,N_5918);
or U6785 (N_6785,N_5914,N_5611);
or U6786 (N_6786,N_5073,N_5477);
nand U6787 (N_6787,N_5212,N_5434);
or U6788 (N_6788,N_5297,N_5955);
nor U6789 (N_6789,N_5523,N_5051);
or U6790 (N_6790,N_5042,N_5487);
nand U6791 (N_6791,N_5649,N_5201);
nor U6792 (N_6792,N_5156,N_5873);
nor U6793 (N_6793,N_5903,N_5415);
xnor U6794 (N_6794,N_5858,N_5566);
nor U6795 (N_6795,N_5215,N_5213);
nand U6796 (N_6796,N_5502,N_5880);
xnor U6797 (N_6797,N_5826,N_5521);
nand U6798 (N_6798,N_5939,N_5466);
xnor U6799 (N_6799,N_5291,N_5281);
or U6800 (N_6800,N_5016,N_5752);
and U6801 (N_6801,N_5966,N_5106);
nand U6802 (N_6802,N_5705,N_5885);
nand U6803 (N_6803,N_5162,N_5378);
and U6804 (N_6804,N_5755,N_5939);
and U6805 (N_6805,N_5235,N_5437);
nand U6806 (N_6806,N_5853,N_5965);
and U6807 (N_6807,N_5516,N_5821);
nand U6808 (N_6808,N_5486,N_5375);
or U6809 (N_6809,N_5084,N_5358);
and U6810 (N_6810,N_5792,N_5019);
and U6811 (N_6811,N_5519,N_5418);
xor U6812 (N_6812,N_5915,N_5142);
nand U6813 (N_6813,N_5680,N_5581);
nor U6814 (N_6814,N_5289,N_5837);
and U6815 (N_6815,N_5215,N_5292);
and U6816 (N_6816,N_5614,N_5529);
or U6817 (N_6817,N_5402,N_5136);
xor U6818 (N_6818,N_5795,N_5514);
xnor U6819 (N_6819,N_5253,N_5146);
and U6820 (N_6820,N_5737,N_5356);
xnor U6821 (N_6821,N_5715,N_5527);
nand U6822 (N_6822,N_5356,N_5137);
and U6823 (N_6823,N_5174,N_5417);
and U6824 (N_6824,N_5904,N_5268);
or U6825 (N_6825,N_5100,N_5846);
nor U6826 (N_6826,N_5743,N_5701);
or U6827 (N_6827,N_5208,N_5419);
nand U6828 (N_6828,N_5628,N_5782);
or U6829 (N_6829,N_5439,N_5435);
xnor U6830 (N_6830,N_5798,N_5824);
or U6831 (N_6831,N_5003,N_5757);
nand U6832 (N_6832,N_5411,N_5141);
nor U6833 (N_6833,N_5724,N_5889);
nand U6834 (N_6834,N_5605,N_5108);
xor U6835 (N_6835,N_5385,N_5492);
xor U6836 (N_6836,N_5627,N_5797);
nand U6837 (N_6837,N_5905,N_5637);
xor U6838 (N_6838,N_5951,N_5482);
xnor U6839 (N_6839,N_5510,N_5987);
nor U6840 (N_6840,N_5077,N_5738);
or U6841 (N_6841,N_5270,N_5063);
xor U6842 (N_6842,N_5965,N_5225);
and U6843 (N_6843,N_5628,N_5984);
nor U6844 (N_6844,N_5934,N_5323);
and U6845 (N_6845,N_5694,N_5778);
nor U6846 (N_6846,N_5811,N_5136);
or U6847 (N_6847,N_5098,N_5464);
and U6848 (N_6848,N_5792,N_5862);
or U6849 (N_6849,N_5125,N_5846);
and U6850 (N_6850,N_5645,N_5886);
and U6851 (N_6851,N_5924,N_5184);
or U6852 (N_6852,N_5281,N_5642);
nor U6853 (N_6853,N_5862,N_5446);
nor U6854 (N_6854,N_5504,N_5322);
and U6855 (N_6855,N_5179,N_5999);
nand U6856 (N_6856,N_5782,N_5106);
nand U6857 (N_6857,N_5175,N_5729);
xnor U6858 (N_6858,N_5145,N_5810);
nor U6859 (N_6859,N_5406,N_5015);
xnor U6860 (N_6860,N_5006,N_5555);
xor U6861 (N_6861,N_5613,N_5209);
and U6862 (N_6862,N_5562,N_5845);
nor U6863 (N_6863,N_5386,N_5230);
nand U6864 (N_6864,N_5641,N_5040);
nor U6865 (N_6865,N_5145,N_5669);
xnor U6866 (N_6866,N_5974,N_5419);
nand U6867 (N_6867,N_5885,N_5846);
and U6868 (N_6868,N_5271,N_5096);
nor U6869 (N_6869,N_5863,N_5880);
and U6870 (N_6870,N_5527,N_5454);
or U6871 (N_6871,N_5135,N_5492);
xnor U6872 (N_6872,N_5863,N_5516);
or U6873 (N_6873,N_5371,N_5257);
nand U6874 (N_6874,N_5100,N_5613);
or U6875 (N_6875,N_5517,N_5205);
nand U6876 (N_6876,N_5405,N_5063);
nor U6877 (N_6877,N_5735,N_5579);
or U6878 (N_6878,N_5989,N_5897);
and U6879 (N_6879,N_5422,N_5012);
xor U6880 (N_6880,N_5641,N_5770);
or U6881 (N_6881,N_5774,N_5815);
and U6882 (N_6882,N_5899,N_5341);
xor U6883 (N_6883,N_5095,N_5566);
nand U6884 (N_6884,N_5998,N_5298);
nor U6885 (N_6885,N_5878,N_5567);
nor U6886 (N_6886,N_5188,N_5943);
and U6887 (N_6887,N_5628,N_5648);
nor U6888 (N_6888,N_5904,N_5761);
and U6889 (N_6889,N_5622,N_5782);
nor U6890 (N_6890,N_5116,N_5862);
or U6891 (N_6891,N_5523,N_5474);
or U6892 (N_6892,N_5768,N_5943);
nand U6893 (N_6893,N_5399,N_5358);
nand U6894 (N_6894,N_5130,N_5092);
xor U6895 (N_6895,N_5470,N_5045);
nor U6896 (N_6896,N_5519,N_5641);
and U6897 (N_6897,N_5189,N_5397);
or U6898 (N_6898,N_5742,N_5129);
and U6899 (N_6899,N_5280,N_5646);
and U6900 (N_6900,N_5776,N_5305);
nand U6901 (N_6901,N_5174,N_5168);
nand U6902 (N_6902,N_5211,N_5491);
nand U6903 (N_6903,N_5372,N_5714);
or U6904 (N_6904,N_5453,N_5848);
and U6905 (N_6905,N_5294,N_5644);
nand U6906 (N_6906,N_5375,N_5003);
or U6907 (N_6907,N_5968,N_5742);
xnor U6908 (N_6908,N_5390,N_5313);
nor U6909 (N_6909,N_5878,N_5260);
or U6910 (N_6910,N_5591,N_5521);
or U6911 (N_6911,N_5353,N_5279);
xor U6912 (N_6912,N_5134,N_5388);
xnor U6913 (N_6913,N_5669,N_5096);
and U6914 (N_6914,N_5081,N_5716);
or U6915 (N_6915,N_5711,N_5957);
or U6916 (N_6916,N_5502,N_5545);
nand U6917 (N_6917,N_5899,N_5304);
xor U6918 (N_6918,N_5206,N_5760);
xnor U6919 (N_6919,N_5069,N_5670);
and U6920 (N_6920,N_5432,N_5609);
nand U6921 (N_6921,N_5761,N_5945);
nor U6922 (N_6922,N_5026,N_5113);
and U6923 (N_6923,N_5478,N_5961);
nand U6924 (N_6924,N_5142,N_5593);
nor U6925 (N_6925,N_5769,N_5306);
nor U6926 (N_6926,N_5576,N_5640);
and U6927 (N_6927,N_5382,N_5300);
or U6928 (N_6928,N_5816,N_5546);
nand U6929 (N_6929,N_5625,N_5010);
nor U6930 (N_6930,N_5476,N_5155);
nand U6931 (N_6931,N_5826,N_5522);
or U6932 (N_6932,N_5762,N_5242);
nand U6933 (N_6933,N_5803,N_5144);
nand U6934 (N_6934,N_5554,N_5995);
and U6935 (N_6935,N_5138,N_5731);
and U6936 (N_6936,N_5402,N_5197);
or U6937 (N_6937,N_5286,N_5656);
and U6938 (N_6938,N_5336,N_5816);
nor U6939 (N_6939,N_5290,N_5655);
xor U6940 (N_6940,N_5271,N_5976);
and U6941 (N_6941,N_5233,N_5041);
nor U6942 (N_6942,N_5977,N_5851);
or U6943 (N_6943,N_5153,N_5031);
xnor U6944 (N_6944,N_5618,N_5832);
or U6945 (N_6945,N_5294,N_5679);
or U6946 (N_6946,N_5568,N_5899);
nor U6947 (N_6947,N_5016,N_5501);
xnor U6948 (N_6948,N_5625,N_5110);
nor U6949 (N_6949,N_5461,N_5021);
nand U6950 (N_6950,N_5714,N_5927);
nor U6951 (N_6951,N_5261,N_5477);
or U6952 (N_6952,N_5417,N_5471);
xor U6953 (N_6953,N_5899,N_5216);
and U6954 (N_6954,N_5097,N_5745);
or U6955 (N_6955,N_5580,N_5039);
xnor U6956 (N_6956,N_5420,N_5193);
xor U6957 (N_6957,N_5290,N_5671);
or U6958 (N_6958,N_5583,N_5736);
and U6959 (N_6959,N_5762,N_5896);
or U6960 (N_6960,N_5892,N_5118);
or U6961 (N_6961,N_5365,N_5798);
nor U6962 (N_6962,N_5366,N_5793);
and U6963 (N_6963,N_5683,N_5213);
nand U6964 (N_6964,N_5783,N_5866);
nand U6965 (N_6965,N_5009,N_5925);
xor U6966 (N_6966,N_5872,N_5066);
nor U6967 (N_6967,N_5944,N_5910);
or U6968 (N_6968,N_5305,N_5445);
and U6969 (N_6969,N_5558,N_5682);
nor U6970 (N_6970,N_5398,N_5275);
nor U6971 (N_6971,N_5849,N_5258);
nand U6972 (N_6972,N_5362,N_5491);
nor U6973 (N_6973,N_5698,N_5318);
and U6974 (N_6974,N_5942,N_5691);
xnor U6975 (N_6975,N_5753,N_5714);
or U6976 (N_6976,N_5018,N_5139);
xor U6977 (N_6977,N_5760,N_5341);
or U6978 (N_6978,N_5546,N_5749);
xnor U6979 (N_6979,N_5783,N_5332);
and U6980 (N_6980,N_5676,N_5812);
xor U6981 (N_6981,N_5468,N_5095);
xnor U6982 (N_6982,N_5433,N_5677);
or U6983 (N_6983,N_5367,N_5525);
nor U6984 (N_6984,N_5089,N_5629);
xnor U6985 (N_6985,N_5896,N_5622);
xnor U6986 (N_6986,N_5649,N_5037);
nand U6987 (N_6987,N_5283,N_5217);
nor U6988 (N_6988,N_5029,N_5941);
or U6989 (N_6989,N_5028,N_5534);
or U6990 (N_6990,N_5100,N_5325);
or U6991 (N_6991,N_5452,N_5863);
nor U6992 (N_6992,N_5687,N_5226);
nor U6993 (N_6993,N_5631,N_5079);
or U6994 (N_6994,N_5885,N_5183);
and U6995 (N_6995,N_5264,N_5336);
xor U6996 (N_6996,N_5907,N_5078);
and U6997 (N_6997,N_5926,N_5813);
xor U6998 (N_6998,N_5244,N_5081);
or U6999 (N_6999,N_5549,N_5232);
and U7000 (N_7000,N_6142,N_6426);
xnor U7001 (N_7001,N_6988,N_6655);
and U7002 (N_7002,N_6631,N_6137);
xor U7003 (N_7003,N_6567,N_6397);
or U7004 (N_7004,N_6084,N_6888);
nand U7005 (N_7005,N_6623,N_6317);
xor U7006 (N_7006,N_6972,N_6902);
nand U7007 (N_7007,N_6000,N_6369);
nand U7008 (N_7008,N_6678,N_6923);
or U7009 (N_7009,N_6189,N_6575);
nor U7010 (N_7010,N_6285,N_6372);
and U7011 (N_7011,N_6277,N_6813);
xnor U7012 (N_7012,N_6169,N_6699);
or U7013 (N_7013,N_6519,N_6584);
or U7014 (N_7014,N_6625,N_6498);
nor U7015 (N_7015,N_6634,N_6136);
nand U7016 (N_7016,N_6957,N_6176);
and U7017 (N_7017,N_6515,N_6722);
or U7018 (N_7018,N_6913,N_6804);
or U7019 (N_7019,N_6344,N_6047);
xor U7020 (N_7020,N_6436,N_6246);
or U7021 (N_7021,N_6561,N_6032);
nor U7022 (N_7022,N_6266,N_6154);
nand U7023 (N_7023,N_6379,N_6129);
nor U7024 (N_7024,N_6670,N_6205);
and U7025 (N_7025,N_6012,N_6537);
xnor U7026 (N_7026,N_6718,N_6256);
nand U7027 (N_7027,N_6881,N_6357);
nand U7028 (N_7028,N_6693,N_6126);
and U7029 (N_7029,N_6072,N_6423);
nor U7030 (N_7030,N_6761,N_6121);
or U7031 (N_7031,N_6080,N_6829);
and U7032 (N_7032,N_6089,N_6076);
nand U7033 (N_7033,N_6273,N_6816);
xnor U7034 (N_7034,N_6139,N_6723);
nor U7035 (N_7035,N_6654,N_6769);
xor U7036 (N_7036,N_6952,N_6918);
and U7037 (N_7037,N_6029,N_6735);
nor U7038 (N_7038,N_6803,N_6251);
xor U7039 (N_7039,N_6242,N_6924);
nand U7040 (N_7040,N_6335,N_6061);
or U7041 (N_7041,N_6647,N_6102);
nor U7042 (N_7042,N_6823,N_6013);
and U7043 (N_7043,N_6527,N_6059);
nor U7044 (N_7044,N_6460,N_6598);
and U7045 (N_7045,N_6283,N_6330);
nand U7046 (N_7046,N_6314,N_6604);
and U7047 (N_7047,N_6481,N_6190);
nor U7048 (N_7048,N_6275,N_6444);
xor U7049 (N_7049,N_6721,N_6704);
xnor U7050 (N_7050,N_6088,N_6668);
xnor U7051 (N_7051,N_6925,N_6135);
nor U7052 (N_7052,N_6238,N_6999);
nor U7053 (N_7053,N_6067,N_6499);
nor U7054 (N_7054,N_6024,N_6635);
and U7055 (N_7055,N_6705,N_6280);
nand U7056 (N_7056,N_6254,N_6627);
nor U7057 (N_7057,N_6962,N_6869);
nand U7058 (N_7058,N_6795,N_6740);
nand U7059 (N_7059,N_6572,N_6733);
nor U7060 (N_7060,N_6853,N_6683);
or U7061 (N_7061,N_6752,N_6742);
and U7062 (N_7062,N_6812,N_6783);
or U7063 (N_7063,N_6198,N_6440);
and U7064 (N_7064,N_6800,N_6381);
or U7065 (N_7065,N_6094,N_6518);
nand U7066 (N_7066,N_6628,N_6115);
or U7067 (N_7067,N_6196,N_6520);
nand U7068 (N_7068,N_6931,N_6960);
and U7069 (N_7069,N_6597,N_6681);
nand U7070 (N_7070,N_6430,N_6062);
xnor U7071 (N_7071,N_6151,N_6428);
or U7072 (N_7072,N_6031,N_6383);
nor U7073 (N_7073,N_6150,N_6548);
or U7074 (N_7074,N_6739,N_6832);
xor U7075 (N_7075,N_6941,N_6595);
and U7076 (N_7076,N_6221,N_6864);
and U7077 (N_7077,N_6282,N_6375);
and U7078 (N_7078,N_6020,N_6979);
nor U7079 (N_7079,N_6741,N_6160);
nand U7080 (N_7080,N_6791,N_6004);
xor U7081 (N_7081,N_6491,N_6778);
nor U7082 (N_7082,N_6985,N_6920);
xor U7083 (N_7083,N_6075,N_6915);
xor U7084 (N_7084,N_6078,N_6616);
or U7085 (N_7085,N_6991,N_6908);
xnor U7086 (N_7086,N_6351,N_6746);
and U7087 (N_7087,N_6123,N_6649);
nand U7088 (N_7088,N_6715,N_6037);
nand U7089 (N_7089,N_6431,N_6919);
or U7090 (N_7090,N_6318,N_6390);
xnor U7091 (N_7091,N_6069,N_6364);
and U7092 (N_7092,N_6987,N_6157);
or U7093 (N_7093,N_6865,N_6663);
or U7094 (N_7094,N_6014,N_6406);
or U7095 (N_7095,N_6103,N_6806);
xnor U7096 (N_7096,N_6578,N_6914);
xor U7097 (N_7097,N_6212,N_6085);
xnor U7098 (N_7098,N_6672,N_6762);
nand U7099 (N_7099,N_6880,N_6992);
nand U7100 (N_7100,N_6976,N_6451);
nor U7101 (N_7101,N_6097,N_6564);
nand U7102 (N_7102,N_6720,N_6544);
nand U7103 (N_7103,N_6732,N_6772);
nor U7104 (N_7104,N_6834,N_6862);
nand U7105 (N_7105,N_6922,N_6686);
or U7106 (N_7106,N_6230,N_6429);
xor U7107 (N_7107,N_6008,N_6214);
xor U7108 (N_7108,N_6099,N_6710);
xnor U7109 (N_7109,N_6901,N_6326);
nand U7110 (N_7110,N_6022,N_6213);
nand U7111 (N_7111,N_6294,N_6437);
nor U7112 (N_7112,N_6724,N_6226);
nand U7113 (N_7113,N_6898,N_6438);
nand U7114 (N_7114,N_6409,N_6968);
and U7115 (N_7115,N_6361,N_6378);
or U7116 (N_7116,N_6837,N_6588);
or U7117 (N_7117,N_6325,N_6808);
and U7118 (N_7118,N_6779,N_6897);
nor U7119 (N_7119,N_6973,N_6509);
nor U7120 (N_7120,N_6677,N_6691);
nand U7121 (N_7121,N_6458,N_6768);
and U7122 (N_7122,N_6650,N_6737);
nor U7123 (N_7123,N_6646,N_6497);
nor U7124 (N_7124,N_6141,N_6109);
xnor U7125 (N_7125,N_6130,N_6817);
and U7126 (N_7126,N_6959,N_6091);
xor U7127 (N_7127,N_6180,N_6336);
or U7128 (N_7128,N_6906,N_6760);
xnor U7129 (N_7129,N_6970,N_6673);
xnor U7130 (N_7130,N_6144,N_6688);
and U7131 (N_7131,N_6514,N_6026);
and U7132 (N_7132,N_6638,N_6844);
xor U7133 (N_7133,N_6048,N_6944);
nand U7134 (N_7134,N_6863,N_6872);
or U7135 (N_7135,N_6156,N_6349);
xnor U7136 (N_7136,N_6455,N_6104);
and U7137 (N_7137,N_6263,N_6164);
nor U7138 (N_7138,N_6482,N_6674);
nand U7139 (N_7139,N_6797,N_6174);
nand U7140 (N_7140,N_6017,N_6172);
or U7141 (N_7141,N_6131,N_6310);
or U7142 (N_7142,N_6521,N_6259);
or U7143 (N_7143,N_6331,N_6081);
nor U7144 (N_7144,N_6776,N_6558);
and U7145 (N_7145,N_6750,N_6755);
nor U7146 (N_7146,N_6111,N_6240);
nand U7147 (N_7147,N_6354,N_6554);
nand U7148 (N_7148,N_6652,N_6193);
nor U7149 (N_7149,N_6353,N_6249);
nand U7150 (N_7150,N_6453,N_6241);
nand U7151 (N_7151,N_6134,N_6942);
or U7152 (N_7152,N_6642,N_6821);
nand U7153 (N_7153,N_6516,N_6402);
nand U7154 (N_7154,N_6245,N_6624);
and U7155 (N_7155,N_6904,N_6345);
nor U7156 (N_7156,N_6528,N_6106);
and U7157 (N_7157,N_6267,N_6984);
nand U7158 (N_7158,N_6165,N_6689);
xnor U7159 (N_7159,N_6609,N_6873);
xnor U7160 (N_7160,N_6511,N_6660);
xor U7161 (N_7161,N_6220,N_6861);
nor U7162 (N_7162,N_6261,N_6830);
nand U7163 (N_7163,N_6030,N_6478);
nand U7164 (N_7164,N_6443,N_6152);
nor U7165 (N_7165,N_6422,N_6745);
or U7166 (N_7166,N_6706,N_6289);
xor U7167 (N_7167,N_6207,N_6237);
nor U7168 (N_7168,N_6889,N_6921);
and U7169 (N_7169,N_6794,N_6435);
or U7170 (N_7170,N_6917,N_6405);
nor U7171 (N_7171,N_6702,N_6868);
and U7172 (N_7172,N_6337,N_6512);
and U7173 (N_7173,N_6155,N_6063);
nor U7174 (N_7174,N_6708,N_6333);
nor U7175 (N_7175,N_6506,N_6954);
and U7176 (N_7176,N_6122,N_6328);
nor U7177 (N_7177,N_6876,N_6346);
xnor U7178 (N_7178,N_6199,N_6937);
or U7179 (N_7179,N_6786,N_6477);
nor U7180 (N_7180,N_6309,N_6990);
and U7181 (N_7181,N_6807,N_6362);
nor U7182 (N_7182,N_6989,N_6223);
xnor U7183 (N_7183,N_6614,N_6640);
xor U7184 (N_7184,N_6279,N_6162);
xnor U7185 (N_7185,N_6473,N_6117);
nor U7186 (N_7186,N_6608,N_6975);
nor U7187 (N_7187,N_6433,N_6981);
or U7188 (N_7188,N_6216,N_6371);
xor U7189 (N_7189,N_6982,N_6879);
and U7190 (N_7190,N_6194,N_6793);
nand U7191 (N_7191,N_6083,N_6645);
xnor U7192 (N_7192,N_6252,N_6260);
and U7193 (N_7193,N_6270,N_6943);
and U7194 (N_7194,N_6736,N_6095);
nor U7195 (N_7195,N_6234,N_6185);
nand U7196 (N_7196,N_6653,N_6232);
nand U7197 (N_7197,N_6492,N_6055);
xor U7198 (N_7198,N_6826,N_6068);
xor U7199 (N_7199,N_6747,N_6993);
nand U7200 (N_7200,N_6296,N_6233);
xnor U7201 (N_7201,N_6946,N_6639);
xnor U7202 (N_7202,N_6530,N_6239);
xnor U7203 (N_7203,N_6738,N_6936);
nor U7204 (N_7204,N_6470,N_6073);
nor U7205 (N_7205,N_6712,N_6394);
nand U7206 (N_7206,N_6366,N_6171);
or U7207 (N_7207,N_6050,N_6229);
nand U7208 (N_7208,N_6562,N_6630);
nand U7209 (N_7209,N_6219,N_6949);
xnor U7210 (N_7210,N_6827,N_6044);
and U7211 (N_7211,N_6494,N_6201);
xnor U7212 (N_7212,N_6694,N_6651);
xor U7213 (N_7213,N_6556,N_6552);
nor U7214 (N_7214,N_6603,N_6235);
xor U7215 (N_7215,N_6687,N_6666);
nor U7216 (N_7216,N_6933,N_6334);
xor U7217 (N_7217,N_6049,N_6713);
or U7218 (N_7218,N_6996,N_6421);
xor U7219 (N_7219,N_6596,N_6555);
and U7220 (N_7220,N_6483,N_6767);
nor U7221 (N_7221,N_6637,N_6502);
nor U7222 (N_7222,N_6633,N_6836);
xor U7223 (N_7223,N_6028,N_6843);
xor U7224 (N_7224,N_6855,N_6472);
and U7225 (N_7225,N_6348,N_6204);
nand U7226 (N_7226,N_6404,N_6560);
nor U7227 (N_7227,N_6181,N_6066);
nor U7228 (N_7228,N_6002,N_6485);
or U7229 (N_7229,N_6659,N_6360);
and U7230 (N_7230,N_6664,N_6247);
nand U7231 (N_7231,N_6716,N_6612);
xnor U7232 (N_7232,N_6680,N_6754);
nand U7233 (N_7233,N_6187,N_6505);
xor U7234 (N_7234,N_6538,N_6057);
xor U7235 (N_7235,N_6711,N_6227);
xor U7236 (N_7236,N_6785,N_6182);
or U7237 (N_7237,N_6591,N_6311);
xnor U7238 (N_7238,N_6475,N_6539);
and U7239 (N_7239,N_6468,N_6676);
and U7240 (N_7240,N_6629,N_6041);
nand U7241 (N_7241,N_6846,N_6493);
or U7242 (N_7242,N_6657,N_6601);
nor U7243 (N_7243,N_6671,N_6413);
and U7244 (N_7244,N_6276,N_6600);
nand U7245 (N_7245,N_6299,N_6025);
and U7246 (N_7246,N_6743,N_6526);
and U7247 (N_7247,N_6753,N_6425);
xnor U7248 (N_7248,N_6692,N_6395);
nor U7249 (N_7249,N_6023,N_6585);
or U7250 (N_7250,N_6964,N_6531);
or U7251 (N_7251,N_6814,N_6582);
or U7252 (N_7252,N_6236,N_6313);
and U7253 (N_7253,N_6107,N_6839);
nor U7254 (N_7254,N_6570,N_6293);
nand U7255 (N_7255,N_6248,N_6669);
nor U7256 (N_7256,N_6452,N_6576);
or U7257 (N_7257,N_6305,N_6714);
and U7258 (N_7258,N_6018,N_6679);
nor U7259 (N_7259,N_6449,N_6120);
nor U7260 (N_7260,N_6748,N_6860);
and U7261 (N_7261,N_6035,N_6599);
and U7262 (N_7262,N_6329,N_6698);
or U7263 (N_7263,N_6304,N_6347);
and U7264 (N_7264,N_6978,N_6594);
nand U7265 (N_7265,N_6665,N_6274);
nand U7266 (N_7266,N_6658,N_6690);
nor U7267 (N_7267,N_6054,N_6052);
and U7268 (N_7268,N_6940,N_6153);
nand U7269 (N_7269,N_6114,N_6454);
and U7270 (N_7270,N_6938,N_6818);
nand U7271 (N_7271,N_6163,N_6859);
or U7272 (N_7272,N_6466,N_6963);
nor U7273 (N_7273,N_6352,N_6302);
nor U7274 (N_7274,N_6132,N_6019);
xnor U7275 (N_7275,N_6424,N_6935);
xor U7276 (N_7276,N_6376,N_6534);
nor U7277 (N_7277,N_6819,N_6847);
nor U7278 (N_7278,N_6191,N_6272);
or U7279 (N_7279,N_6667,N_6765);
and U7280 (N_7280,N_6995,N_6866);
xor U7281 (N_7281,N_6811,N_6587);
nand U7282 (N_7282,N_6503,N_6086);
or U7283 (N_7283,N_6341,N_6486);
xnor U7284 (N_7284,N_6684,N_6148);
nor U7285 (N_7285,N_6757,N_6893);
nor U7286 (N_7286,N_6065,N_6374);
nand U7287 (N_7287,N_6469,N_6224);
and U7288 (N_7288,N_6725,N_6589);
or U7289 (N_7289,N_6950,N_6320);
nor U7290 (N_7290,N_6340,N_6384);
nand U7291 (N_7291,N_6077,N_6557);
or U7292 (N_7292,N_6119,N_6877);
xnor U7293 (N_7293,N_6926,N_6580);
nor U7294 (N_7294,N_6766,N_6618);
and U7295 (N_7295,N_6231,N_6202);
and U7296 (N_7296,N_6391,N_6489);
and U7297 (N_7297,N_6380,N_6418);
and U7298 (N_7298,N_6675,N_6851);
or U7299 (N_7299,N_6363,N_6036);
nor U7300 (N_7300,N_6894,N_6291);
or U7301 (N_7301,N_6886,N_6206);
nand U7302 (N_7302,N_6143,N_6961);
or U7303 (N_7303,N_6188,N_6271);
nand U7304 (N_7304,N_6178,N_6415);
nor U7305 (N_7305,N_6524,N_6756);
nor U7306 (N_7306,N_6719,N_6849);
nor U7307 (N_7307,N_6034,N_6884);
or U7308 (N_7308,N_6316,N_6411);
nor U7309 (N_7309,N_6900,N_6420);
nor U7310 (N_7310,N_6464,N_6764);
nor U7311 (N_7311,N_6883,N_6845);
and U7312 (N_7312,N_6459,N_6112);
nor U7313 (N_7313,N_6749,N_6593);
xnor U7314 (N_7314,N_6324,N_6321);
nor U7315 (N_7315,N_6441,N_6396);
and U7316 (N_7316,N_6140,N_6244);
nor U7317 (N_7317,N_6367,N_6096);
nand U7318 (N_7318,N_6474,N_6278);
nor U7319 (N_7319,N_6533,N_6726);
and U7320 (N_7320,N_6222,N_6432);
and U7321 (N_7321,N_6265,N_6382);
nor U7322 (N_7322,N_6264,N_6090);
nand U7323 (N_7323,N_6298,N_6701);
xor U7324 (N_7324,N_6930,N_6001);
nand U7325 (N_7325,N_6166,N_6541);
nand U7326 (N_7326,N_6445,N_6308);
or U7327 (N_7327,N_6798,N_6997);
nand U7328 (N_7328,N_6602,N_6773);
nand U7329 (N_7329,N_6332,N_6504);
nor U7330 (N_7330,N_6038,N_6934);
nand U7331 (N_7331,N_6365,N_6110);
or U7332 (N_7332,N_6288,N_6398);
nand U7333 (N_7333,N_6911,N_6442);
xor U7334 (N_7334,N_6403,N_6401);
xnor U7335 (N_7335,N_6709,N_6955);
nand U7336 (N_7336,N_6033,N_6540);
nand U7337 (N_7337,N_6118,N_6858);
nor U7338 (N_7338,N_6508,N_6281);
nor U7339 (N_7339,N_6532,N_6983);
or U7340 (N_7340,N_6565,N_6895);
nand U7341 (N_7341,N_6007,N_6899);
and U7342 (N_7342,N_6043,N_6356);
or U7343 (N_7343,N_6461,N_6124);
xnor U7344 (N_7344,N_6446,N_6292);
nand U7345 (N_7345,N_6801,N_6301);
nand U7346 (N_7346,N_6703,N_6799);
nand U7347 (N_7347,N_6286,N_6543);
xor U7348 (N_7348,N_6974,N_6300);
nand U7349 (N_7349,N_6948,N_6087);
nor U7350 (N_7350,N_6700,N_6416);
nor U7351 (N_7351,N_6805,N_6101);
or U7352 (N_7352,N_6912,N_6082);
nand U7353 (N_7353,N_6734,N_6343);
and U7354 (N_7354,N_6542,N_6175);
and U7355 (N_7355,N_6427,N_6338);
and U7356 (N_7356,N_6586,N_6792);
or U7357 (N_7357,N_6070,N_6967);
or U7358 (N_7358,N_6450,N_6809);
nand U7359 (N_7359,N_6850,N_6622);
or U7360 (N_7360,N_6513,N_6006);
and U7361 (N_7361,N_6891,N_6463);
and U7362 (N_7362,N_6496,N_6177);
and U7363 (N_7363,N_6547,N_6759);
and U7364 (N_7364,N_6966,N_6389);
and U7365 (N_7365,N_6414,N_6787);
nand U7366 (N_7366,N_6225,N_6021);
or U7367 (N_7367,N_6731,N_6183);
or U7368 (N_7368,N_6476,N_6751);
or U7369 (N_7369,N_6951,N_6928);
nor U7370 (N_7370,N_6385,N_6763);
and U7371 (N_7371,N_6268,N_6312);
nor U7372 (N_7372,N_6386,N_6856);
nand U7373 (N_7373,N_6887,N_6566);
or U7374 (N_7374,N_6200,N_6867);
nand U7375 (N_7375,N_6857,N_6824);
nand U7376 (N_7376,N_6071,N_6848);
or U7377 (N_7377,N_6835,N_6074);
xnor U7378 (N_7378,N_6841,N_6517);
nor U7379 (N_7379,N_6387,N_6656);
and U7380 (N_7380,N_6620,N_6977);
nand U7381 (N_7381,N_6456,N_6146);
or U7382 (N_7382,N_6307,N_6810);
or U7383 (N_7383,N_6885,N_6412);
or U7384 (N_7384,N_6854,N_6648);
and U7385 (N_7385,N_6255,N_6831);
nor U7386 (N_7386,N_6133,N_6100);
nor U7387 (N_7387,N_6661,N_6011);
xnor U7388 (N_7388,N_6003,N_6697);
or U7389 (N_7389,N_6770,N_6319);
and U7390 (N_7390,N_6563,N_6480);
and U7391 (N_7391,N_6833,N_6501);
nor U7392 (N_7392,N_6388,N_6253);
nand U7393 (N_7393,N_6632,N_6549);
xnor U7394 (N_7394,N_6125,N_6790);
nor U7395 (N_7395,N_6568,N_6315);
or U7396 (N_7396,N_6053,N_6641);
nand U7397 (N_7397,N_6257,N_6434);
and U7398 (N_7398,N_6579,N_6471);
xor U7399 (N_7399,N_6870,N_6553);
and U7400 (N_7400,N_6909,N_6728);
and U7401 (N_7401,N_6287,N_6744);
or U7402 (N_7402,N_6243,N_6487);
xnor U7403 (N_7403,N_6467,N_6145);
nor U7404 (N_7404,N_6010,N_6215);
nor U7405 (N_7405,N_6878,N_6621);
xnor U7406 (N_7406,N_6815,N_6173);
and U7407 (N_7407,N_6350,N_6258);
xor U7408 (N_7408,N_6262,N_6092);
nor U7409 (N_7409,N_6611,N_6184);
or U7410 (N_7410,N_6550,N_6500);
xor U7411 (N_7411,N_6535,N_6373);
nand U7412 (N_7412,N_6939,N_6758);
nand U7413 (N_7413,N_6462,N_6027);
or U7414 (N_7414,N_6820,N_6905);
or U7415 (N_7415,N_6852,N_6626);
nand U7416 (N_7416,N_6377,N_6781);
nor U7417 (N_7417,N_6788,N_6186);
or U7418 (N_7418,N_6158,N_6203);
xnor U7419 (N_7419,N_6980,N_6170);
or U7420 (N_7420,N_6370,N_6965);
or U7421 (N_7421,N_6577,N_6060);
nand U7422 (N_7422,N_6932,N_6093);
and U7423 (N_7423,N_6945,N_6840);
xnor U7424 (N_7424,N_6573,N_6610);
nor U7425 (N_7425,N_6005,N_6392);
or U7426 (N_7426,N_6168,N_6210);
nor U7427 (N_7427,N_6771,N_6228);
nor U7428 (N_7428,N_6465,N_6882);
xnor U7429 (N_7429,N_6128,N_6559);
and U7430 (N_7430,N_6998,N_6399);
nand U7431 (N_7431,N_6479,N_6167);
and U7432 (N_7432,N_6323,N_6994);
xnor U7433 (N_7433,N_6617,N_6571);
and U7434 (N_7434,N_6009,N_6605);
or U7435 (N_7435,N_6147,N_6907);
xor U7436 (N_7436,N_6197,N_6507);
or U7437 (N_7437,N_6211,N_6953);
and U7438 (N_7438,N_6583,N_6838);
or U7439 (N_7439,N_6138,N_6777);
nor U7440 (N_7440,N_6495,N_6490);
xnor U7441 (N_7441,N_6149,N_6417);
xor U7442 (N_7442,N_6042,N_6510);
nor U7443 (N_7443,N_6297,N_6545);
nand U7444 (N_7444,N_6682,N_6016);
or U7445 (N_7445,N_6729,N_6208);
and U7446 (N_7446,N_6569,N_6929);
and U7447 (N_7447,N_6040,N_6615);
xnor U7448 (N_7448,N_6971,N_6113);
nor U7449 (N_7449,N_6339,N_6916);
nand U7450 (N_7450,N_6956,N_6051);
or U7451 (N_7451,N_6796,N_6046);
and U7452 (N_7452,N_6116,N_6717);
nand U7453 (N_7453,N_6546,N_6613);
xor U7454 (N_7454,N_6662,N_6368);
or U7455 (N_7455,N_6488,N_6161);
xor U7456 (N_7456,N_6407,N_6727);
nor U7457 (N_7457,N_6643,N_6782);
and U7458 (N_7458,N_6192,N_6400);
or U7459 (N_7459,N_6056,N_6523);
and U7460 (N_7460,N_6484,N_6695);
and U7461 (N_7461,N_6574,N_6636);
or U7462 (N_7462,N_6355,N_6871);
or U7463 (N_7463,N_6875,N_6306);
and U7464 (N_7464,N_6775,N_6322);
xnor U7465 (N_7465,N_6696,N_6015);
and U7466 (N_7466,N_6079,N_6303);
and U7467 (N_7467,N_6927,N_6619);
xnor U7468 (N_7468,N_6269,N_6410);
nand U7469 (N_7469,N_6903,N_6098);
nand U7470 (N_7470,N_6892,N_6290);
xor U7471 (N_7471,N_6457,N_6969);
and U7472 (N_7472,N_6986,N_6536);
nand U7473 (N_7473,N_6707,N_6685);
and U7474 (N_7474,N_6780,N_6359);
and U7475 (N_7475,N_6342,N_6393);
and U7476 (N_7476,N_6644,N_6408);
and U7477 (N_7477,N_6284,N_6295);
and U7478 (N_7478,N_6058,N_6179);
and U7479 (N_7479,N_6802,N_6606);
and U7480 (N_7480,N_6947,N_6958);
nor U7481 (N_7481,N_6195,N_6828);
nand U7482 (N_7482,N_6159,N_6127);
xor U7483 (N_7483,N_6250,N_6825);
nor U7484 (N_7484,N_6064,N_6217);
nor U7485 (N_7485,N_6525,N_6730);
xor U7486 (N_7486,N_6842,N_6039);
xnor U7487 (N_7487,N_6874,N_6551);
and U7488 (N_7488,N_6896,N_6774);
xor U7489 (N_7489,N_6592,N_6358);
nor U7490 (N_7490,N_6822,N_6581);
and U7491 (N_7491,N_6590,N_6108);
nor U7492 (N_7492,N_6209,N_6419);
xnor U7493 (N_7493,N_6784,N_6522);
and U7494 (N_7494,N_6529,N_6607);
or U7495 (N_7495,N_6910,N_6890);
xor U7496 (N_7496,N_6218,N_6447);
nor U7497 (N_7497,N_6439,N_6045);
or U7498 (N_7498,N_6789,N_6105);
xnor U7499 (N_7499,N_6327,N_6448);
nand U7500 (N_7500,N_6514,N_6471);
xor U7501 (N_7501,N_6760,N_6162);
nand U7502 (N_7502,N_6448,N_6070);
xnor U7503 (N_7503,N_6286,N_6311);
nand U7504 (N_7504,N_6214,N_6097);
nor U7505 (N_7505,N_6867,N_6391);
xor U7506 (N_7506,N_6206,N_6875);
or U7507 (N_7507,N_6966,N_6610);
and U7508 (N_7508,N_6107,N_6983);
nor U7509 (N_7509,N_6547,N_6715);
xnor U7510 (N_7510,N_6445,N_6318);
xor U7511 (N_7511,N_6464,N_6127);
nand U7512 (N_7512,N_6773,N_6365);
and U7513 (N_7513,N_6570,N_6229);
or U7514 (N_7514,N_6975,N_6261);
nor U7515 (N_7515,N_6288,N_6035);
or U7516 (N_7516,N_6437,N_6277);
xnor U7517 (N_7517,N_6101,N_6566);
nand U7518 (N_7518,N_6964,N_6031);
nor U7519 (N_7519,N_6600,N_6931);
or U7520 (N_7520,N_6390,N_6947);
nand U7521 (N_7521,N_6765,N_6771);
nor U7522 (N_7522,N_6336,N_6565);
nor U7523 (N_7523,N_6259,N_6082);
xor U7524 (N_7524,N_6516,N_6202);
and U7525 (N_7525,N_6497,N_6050);
nand U7526 (N_7526,N_6850,N_6267);
or U7527 (N_7527,N_6763,N_6138);
nand U7528 (N_7528,N_6883,N_6432);
xnor U7529 (N_7529,N_6838,N_6883);
and U7530 (N_7530,N_6151,N_6209);
or U7531 (N_7531,N_6837,N_6620);
nand U7532 (N_7532,N_6152,N_6280);
xor U7533 (N_7533,N_6067,N_6296);
nand U7534 (N_7534,N_6460,N_6905);
or U7535 (N_7535,N_6145,N_6262);
or U7536 (N_7536,N_6056,N_6356);
or U7537 (N_7537,N_6654,N_6861);
nor U7538 (N_7538,N_6130,N_6905);
or U7539 (N_7539,N_6266,N_6607);
xor U7540 (N_7540,N_6265,N_6432);
xor U7541 (N_7541,N_6309,N_6031);
nand U7542 (N_7542,N_6542,N_6552);
nand U7543 (N_7543,N_6386,N_6507);
and U7544 (N_7544,N_6615,N_6345);
nor U7545 (N_7545,N_6498,N_6063);
nand U7546 (N_7546,N_6093,N_6823);
and U7547 (N_7547,N_6795,N_6135);
and U7548 (N_7548,N_6756,N_6499);
nand U7549 (N_7549,N_6533,N_6932);
xor U7550 (N_7550,N_6825,N_6925);
nor U7551 (N_7551,N_6696,N_6678);
nand U7552 (N_7552,N_6892,N_6564);
or U7553 (N_7553,N_6276,N_6611);
nand U7554 (N_7554,N_6515,N_6786);
or U7555 (N_7555,N_6592,N_6472);
and U7556 (N_7556,N_6781,N_6037);
and U7557 (N_7557,N_6659,N_6563);
xor U7558 (N_7558,N_6295,N_6932);
nor U7559 (N_7559,N_6975,N_6615);
nand U7560 (N_7560,N_6315,N_6051);
nor U7561 (N_7561,N_6720,N_6944);
or U7562 (N_7562,N_6890,N_6423);
nand U7563 (N_7563,N_6996,N_6412);
or U7564 (N_7564,N_6909,N_6515);
and U7565 (N_7565,N_6911,N_6807);
nor U7566 (N_7566,N_6768,N_6631);
and U7567 (N_7567,N_6224,N_6839);
xor U7568 (N_7568,N_6249,N_6718);
or U7569 (N_7569,N_6924,N_6922);
or U7570 (N_7570,N_6654,N_6562);
xor U7571 (N_7571,N_6450,N_6333);
or U7572 (N_7572,N_6239,N_6003);
nor U7573 (N_7573,N_6678,N_6673);
and U7574 (N_7574,N_6797,N_6036);
nand U7575 (N_7575,N_6819,N_6822);
nor U7576 (N_7576,N_6157,N_6915);
and U7577 (N_7577,N_6097,N_6122);
nor U7578 (N_7578,N_6549,N_6628);
nor U7579 (N_7579,N_6743,N_6831);
nor U7580 (N_7580,N_6628,N_6607);
nand U7581 (N_7581,N_6460,N_6632);
or U7582 (N_7582,N_6792,N_6843);
and U7583 (N_7583,N_6596,N_6171);
nand U7584 (N_7584,N_6204,N_6514);
xnor U7585 (N_7585,N_6349,N_6832);
nand U7586 (N_7586,N_6343,N_6574);
or U7587 (N_7587,N_6311,N_6564);
and U7588 (N_7588,N_6949,N_6101);
xnor U7589 (N_7589,N_6372,N_6198);
nor U7590 (N_7590,N_6348,N_6357);
nor U7591 (N_7591,N_6450,N_6484);
or U7592 (N_7592,N_6444,N_6425);
or U7593 (N_7593,N_6432,N_6261);
and U7594 (N_7594,N_6670,N_6331);
xnor U7595 (N_7595,N_6008,N_6939);
and U7596 (N_7596,N_6775,N_6908);
nand U7597 (N_7597,N_6483,N_6516);
or U7598 (N_7598,N_6293,N_6816);
or U7599 (N_7599,N_6902,N_6745);
nor U7600 (N_7600,N_6229,N_6023);
xnor U7601 (N_7601,N_6411,N_6106);
xnor U7602 (N_7602,N_6867,N_6467);
xnor U7603 (N_7603,N_6330,N_6535);
or U7604 (N_7604,N_6580,N_6838);
and U7605 (N_7605,N_6285,N_6262);
xnor U7606 (N_7606,N_6669,N_6767);
nand U7607 (N_7607,N_6077,N_6454);
and U7608 (N_7608,N_6713,N_6469);
nor U7609 (N_7609,N_6036,N_6050);
and U7610 (N_7610,N_6867,N_6622);
nor U7611 (N_7611,N_6866,N_6337);
nand U7612 (N_7612,N_6754,N_6540);
nor U7613 (N_7613,N_6526,N_6178);
nand U7614 (N_7614,N_6336,N_6067);
nand U7615 (N_7615,N_6722,N_6635);
or U7616 (N_7616,N_6284,N_6376);
xor U7617 (N_7617,N_6271,N_6328);
or U7618 (N_7618,N_6544,N_6156);
or U7619 (N_7619,N_6932,N_6483);
or U7620 (N_7620,N_6072,N_6672);
nor U7621 (N_7621,N_6883,N_6614);
and U7622 (N_7622,N_6694,N_6537);
or U7623 (N_7623,N_6496,N_6792);
xor U7624 (N_7624,N_6361,N_6701);
and U7625 (N_7625,N_6110,N_6085);
and U7626 (N_7626,N_6997,N_6255);
nand U7627 (N_7627,N_6621,N_6466);
or U7628 (N_7628,N_6625,N_6954);
nand U7629 (N_7629,N_6180,N_6006);
nor U7630 (N_7630,N_6893,N_6445);
or U7631 (N_7631,N_6360,N_6972);
xnor U7632 (N_7632,N_6439,N_6062);
and U7633 (N_7633,N_6222,N_6732);
nor U7634 (N_7634,N_6883,N_6344);
and U7635 (N_7635,N_6119,N_6434);
xnor U7636 (N_7636,N_6825,N_6995);
nand U7637 (N_7637,N_6018,N_6364);
nand U7638 (N_7638,N_6973,N_6958);
nand U7639 (N_7639,N_6436,N_6811);
xnor U7640 (N_7640,N_6241,N_6972);
and U7641 (N_7641,N_6491,N_6021);
xor U7642 (N_7642,N_6942,N_6744);
or U7643 (N_7643,N_6463,N_6980);
nand U7644 (N_7644,N_6060,N_6354);
nand U7645 (N_7645,N_6698,N_6292);
xnor U7646 (N_7646,N_6417,N_6281);
xor U7647 (N_7647,N_6714,N_6527);
nor U7648 (N_7648,N_6328,N_6427);
xnor U7649 (N_7649,N_6047,N_6271);
and U7650 (N_7650,N_6995,N_6762);
and U7651 (N_7651,N_6998,N_6745);
and U7652 (N_7652,N_6051,N_6518);
xor U7653 (N_7653,N_6415,N_6242);
nand U7654 (N_7654,N_6670,N_6184);
nor U7655 (N_7655,N_6272,N_6209);
nor U7656 (N_7656,N_6332,N_6750);
nor U7657 (N_7657,N_6852,N_6218);
nor U7658 (N_7658,N_6184,N_6479);
nor U7659 (N_7659,N_6493,N_6523);
nor U7660 (N_7660,N_6662,N_6009);
and U7661 (N_7661,N_6805,N_6340);
xnor U7662 (N_7662,N_6340,N_6514);
xnor U7663 (N_7663,N_6219,N_6082);
and U7664 (N_7664,N_6165,N_6030);
and U7665 (N_7665,N_6934,N_6674);
xor U7666 (N_7666,N_6770,N_6681);
and U7667 (N_7667,N_6512,N_6915);
and U7668 (N_7668,N_6754,N_6548);
or U7669 (N_7669,N_6972,N_6508);
nand U7670 (N_7670,N_6529,N_6077);
or U7671 (N_7671,N_6074,N_6347);
nand U7672 (N_7672,N_6908,N_6451);
or U7673 (N_7673,N_6131,N_6248);
xor U7674 (N_7674,N_6422,N_6533);
nand U7675 (N_7675,N_6735,N_6360);
or U7676 (N_7676,N_6699,N_6748);
and U7677 (N_7677,N_6326,N_6677);
nand U7678 (N_7678,N_6917,N_6464);
or U7679 (N_7679,N_6325,N_6968);
nand U7680 (N_7680,N_6013,N_6493);
xnor U7681 (N_7681,N_6880,N_6818);
nand U7682 (N_7682,N_6474,N_6852);
nand U7683 (N_7683,N_6490,N_6606);
nand U7684 (N_7684,N_6203,N_6360);
nor U7685 (N_7685,N_6088,N_6603);
nor U7686 (N_7686,N_6749,N_6201);
nand U7687 (N_7687,N_6537,N_6116);
nand U7688 (N_7688,N_6780,N_6639);
nor U7689 (N_7689,N_6785,N_6159);
xor U7690 (N_7690,N_6497,N_6292);
xor U7691 (N_7691,N_6431,N_6623);
or U7692 (N_7692,N_6339,N_6366);
and U7693 (N_7693,N_6583,N_6370);
nor U7694 (N_7694,N_6921,N_6544);
or U7695 (N_7695,N_6595,N_6567);
xor U7696 (N_7696,N_6093,N_6554);
xnor U7697 (N_7697,N_6099,N_6414);
and U7698 (N_7698,N_6070,N_6441);
or U7699 (N_7699,N_6246,N_6565);
nor U7700 (N_7700,N_6767,N_6674);
or U7701 (N_7701,N_6416,N_6355);
nor U7702 (N_7702,N_6871,N_6763);
and U7703 (N_7703,N_6906,N_6512);
xor U7704 (N_7704,N_6199,N_6662);
xnor U7705 (N_7705,N_6320,N_6273);
xnor U7706 (N_7706,N_6902,N_6619);
nor U7707 (N_7707,N_6210,N_6146);
nor U7708 (N_7708,N_6714,N_6755);
nor U7709 (N_7709,N_6694,N_6846);
or U7710 (N_7710,N_6398,N_6166);
and U7711 (N_7711,N_6311,N_6996);
xnor U7712 (N_7712,N_6306,N_6318);
and U7713 (N_7713,N_6552,N_6561);
or U7714 (N_7714,N_6775,N_6114);
nor U7715 (N_7715,N_6010,N_6778);
or U7716 (N_7716,N_6233,N_6424);
or U7717 (N_7717,N_6143,N_6182);
nor U7718 (N_7718,N_6835,N_6052);
xnor U7719 (N_7719,N_6654,N_6220);
or U7720 (N_7720,N_6686,N_6422);
or U7721 (N_7721,N_6652,N_6709);
nor U7722 (N_7722,N_6602,N_6377);
or U7723 (N_7723,N_6994,N_6953);
nor U7724 (N_7724,N_6381,N_6243);
and U7725 (N_7725,N_6759,N_6651);
and U7726 (N_7726,N_6604,N_6829);
and U7727 (N_7727,N_6847,N_6069);
xor U7728 (N_7728,N_6979,N_6003);
nor U7729 (N_7729,N_6647,N_6844);
or U7730 (N_7730,N_6894,N_6530);
xnor U7731 (N_7731,N_6798,N_6925);
xnor U7732 (N_7732,N_6385,N_6289);
nand U7733 (N_7733,N_6032,N_6616);
and U7734 (N_7734,N_6396,N_6733);
nor U7735 (N_7735,N_6947,N_6136);
nand U7736 (N_7736,N_6920,N_6515);
xnor U7737 (N_7737,N_6662,N_6342);
xnor U7738 (N_7738,N_6544,N_6676);
xor U7739 (N_7739,N_6113,N_6427);
xor U7740 (N_7740,N_6022,N_6849);
nor U7741 (N_7741,N_6117,N_6138);
nor U7742 (N_7742,N_6183,N_6543);
nor U7743 (N_7743,N_6527,N_6267);
nand U7744 (N_7744,N_6232,N_6159);
and U7745 (N_7745,N_6209,N_6252);
xnor U7746 (N_7746,N_6551,N_6238);
or U7747 (N_7747,N_6158,N_6402);
and U7748 (N_7748,N_6918,N_6379);
and U7749 (N_7749,N_6164,N_6301);
or U7750 (N_7750,N_6091,N_6084);
nor U7751 (N_7751,N_6711,N_6036);
or U7752 (N_7752,N_6534,N_6005);
xor U7753 (N_7753,N_6682,N_6137);
and U7754 (N_7754,N_6247,N_6102);
and U7755 (N_7755,N_6102,N_6761);
and U7756 (N_7756,N_6818,N_6299);
nand U7757 (N_7757,N_6051,N_6904);
or U7758 (N_7758,N_6985,N_6393);
and U7759 (N_7759,N_6513,N_6137);
or U7760 (N_7760,N_6632,N_6986);
nor U7761 (N_7761,N_6521,N_6003);
xor U7762 (N_7762,N_6378,N_6808);
xnor U7763 (N_7763,N_6053,N_6027);
and U7764 (N_7764,N_6202,N_6160);
and U7765 (N_7765,N_6742,N_6591);
and U7766 (N_7766,N_6250,N_6635);
or U7767 (N_7767,N_6670,N_6790);
or U7768 (N_7768,N_6936,N_6679);
and U7769 (N_7769,N_6625,N_6109);
nor U7770 (N_7770,N_6687,N_6510);
nor U7771 (N_7771,N_6554,N_6250);
nand U7772 (N_7772,N_6700,N_6534);
xor U7773 (N_7773,N_6019,N_6909);
nor U7774 (N_7774,N_6084,N_6113);
xnor U7775 (N_7775,N_6330,N_6022);
and U7776 (N_7776,N_6920,N_6852);
nor U7777 (N_7777,N_6835,N_6480);
nand U7778 (N_7778,N_6285,N_6602);
nand U7779 (N_7779,N_6622,N_6988);
and U7780 (N_7780,N_6681,N_6923);
nand U7781 (N_7781,N_6956,N_6379);
or U7782 (N_7782,N_6694,N_6603);
xnor U7783 (N_7783,N_6153,N_6327);
and U7784 (N_7784,N_6094,N_6533);
nor U7785 (N_7785,N_6024,N_6937);
xnor U7786 (N_7786,N_6722,N_6636);
nor U7787 (N_7787,N_6559,N_6440);
and U7788 (N_7788,N_6831,N_6503);
and U7789 (N_7789,N_6820,N_6536);
or U7790 (N_7790,N_6318,N_6190);
nand U7791 (N_7791,N_6696,N_6280);
or U7792 (N_7792,N_6339,N_6273);
or U7793 (N_7793,N_6972,N_6122);
nor U7794 (N_7794,N_6254,N_6821);
and U7795 (N_7795,N_6598,N_6356);
or U7796 (N_7796,N_6814,N_6051);
and U7797 (N_7797,N_6665,N_6612);
and U7798 (N_7798,N_6856,N_6852);
nand U7799 (N_7799,N_6028,N_6827);
or U7800 (N_7800,N_6025,N_6254);
nor U7801 (N_7801,N_6371,N_6584);
and U7802 (N_7802,N_6186,N_6711);
or U7803 (N_7803,N_6732,N_6579);
or U7804 (N_7804,N_6501,N_6330);
nor U7805 (N_7805,N_6404,N_6065);
or U7806 (N_7806,N_6218,N_6573);
nor U7807 (N_7807,N_6542,N_6155);
nor U7808 (N_7808,N_6002,N_6029);
or U7809 (N_7809,N_6407,N_6332);
xor U7810 (N_7810,N_6456,N_6590);
nand U7811 (N_7811,N_6775,N_6563);
or U7812 (N_7812,N_6766,N_6403);
nand U7813 (N_7813,N_6756,N_6225);
and U7814 (N_7814,N_6990,N_6177);
xor U7815 (N_7815,N_6386,N_6425);
xor U7816 (N_7816,N_6469,N_6994);
nand U7817 (N_7817,N_6097,N_6448);
nand U7818 (N_7818,N_6947,N_6659);
nand U7819 (N_7819,N_6419,N_6263);
nor U7820 (N_7820,N_6435,N_6966);
or U7821 (N_7821,N_6524,N_6283);
nand U7822 (N_7822,N_6192,N_6481);
xnor U7823 (N_7823,N_6118,N_6602);
and U7824 (N_7824,N_6205,N_6024);
nand U7825 (N_7825,N_6798,N_6384);
or U7826 (N_7826,N_6318,N_6798);
and U7827 (N_7827,N_6487,N_6110);
nand U7828 (N_7828,N_6838,N_6236);
xor U7829 (N_7829,N_6883,N_6026);
nand U7830 (N_7830,N_6649,N_6810);
nor U7831 (N_7831,N_6509,N_6409);
xnor U7832 (N_7832,N_6371,N_6041);
xnor U7833 (N_7833,N_6673,N_6914);
nand U7834 (N_7834,N_6934,N_6006);
xor U7835 (N_7835,N_6203,N_6877);
nand U7836 (N_7836,N_6492,N_6961);
and U7837 (N_7837,N_6195,N_6932);
and U7838 (N_7838,N_6117,N_6162);
nor U7839 (N_7839,N_6037,N_6284);
xnor U7840 (N_7840,N_6216,N_6965);
or U7841 (N_7841,N_6249,N_6361);
or U7842 (N_7842,N_6789,N_6778);
or U7843 (N_7843,N_6117,N_6574);
and U7844 (N_7844,N_6432,N_6568);
nand U7845 (N_7845,N_6966,N_6349);
or U7846 (N_7846,N_6949,N_6521);
nor U7847 (N_7847,N_6314,N_6131);
xnor U7848 (N_7848,N_6072,N_6860);
xor U7849 (N_7849,N_6385,N_6083);
nor U7850 (N_7850,N_6670,N_6200);
or U7851 (N_7851,N_6867,N_6130);
nor U7852 (N_7852,N_6872,N_6350);
and U7853 (N_7853,N_6006,N_6005);
xnor U7854 (N_7854,N_6649,N_6734);
nor U7855 (N_7855,N_6545,N_6228);
nor U7856 (N_7856,N_6001,N_6214);
xnor U7857 (N_7857,N_6994,N_6601);
nand U7858 (N_7858,N_6915,N_6412);
and U7859 (N_7859,N_6719,N_6751);
or U7860 (N_7860,N_6505,N_6339);
nor U7861 (N_7861,N_6378,N_6265);
or U7862 (N_7862,N_6657,N_6051);
nand U7863 (N_7863,N_6941,N_6598);
nor U7864 (N_7864,N_6596,N_6611);
and U7865 (N_7865,N_6931,N_6095);
and U7866 (N_7866,N_6008,N_6847);
nor U7867 (N_7867,N_6998,N_6474);
and U7868 (N_7868,N_6409,N_6684);
nor U7869 (N_7869,N_6703,N_6771);
nor U7870 (N_7870,N_6672,N_6028);
and U7871 (N_7871,N_6020,N_6616);
or U7872 (N_7872,N_6892,N_6028);
xnor U7873 (N_7873,N_6561,N_6795);
and U7874 (N_7874,N_6585,N_6225);
nor U7875 (N_7875,N_6647,N_6486);
and U7876 (N_7876,N_6363,N_6380);
nor U7877 (N_7877,N_6644,N_6567);
nor U7878 (N_7878,N_6773,N_6088);
or U7879 (N_7879,N_6751,N_6422);
xnor U7880 (N_7880,N_6944,N_6951);
xnor U7881 (N_7881,N_6199,N_6756);
or U7882 (N_7882,N_6342,N_6231);
nor U7883 (N_7883,N_6924,N_6970);
nor U7884 (N_7884,N_6233,N_6665);
nor U7885 (N_7885,N_6375,N_6717);
nand U7886 (N_7886,N_6745,N_6935);
or U7887 (N_7887,N_6482,N_6373);
nor U7888 (N_7888,N_6326,N_6500);
or U7889 (N_7889,N_6028,N_6407);
nand U7890 (N_7890,N_6375,N_6135);
nor U7891 (N_7891,N_6064,N_6820);
xor U7892 (N_7892,N_6407,N_6449);
and U7893 (N_7893,N_6583,N_6185);
xor U7894 (N_7894,N_6825,N_6981);
nor U7895 (N_7895,N_6264,N_6670);
and U7896 (N_7896,N_6070,N_6782);
nor U7897 (N_7897,N_6675,N_6593);
nor U7898 (N_7898,N_6336,N_6064);
or U7899 (N_7899,N_6185,N_6436);
or U7900 (N_7900,N_6409,N_6030);
and U7901 (N_7901,N_6918,N_6270);
nor U7902 (N_7902,N_6997,N_6816);
nor U7903 (N_7903,N_6483,N_6459);
and U7904 (N_7904,N_6693,N_6749);
and U7905 (N_7905,N_6034,N_6186);
or U7906 (N_7906,N_6852,N_6818);
nand U7907 (N_7907,N_6784,N_6068);
nand U7908 (N_7908,N_6127,N_6671);
or U7909 (N_7909,N_6049,N_6337);
nand U7910 (N_7910,N_6407,N_6242);
nor U7911 (N_7911,N_6914,N_6764);
nand U7912 (N_7912,N_6502,N_6184);
xor U7913 (N_7913,N_6797,N_6846);
xnor U7914 (N_7914,N_6701,N_6183);
nand U7915 (N_7915,N_6381,N_6025);
or U7916 (N_7916,N_6799,N_6812);
or U7917 (N_7917,N_6167,N_6422);
and U7918 (N_7918,N_6253,N_6295);
nand U7919 (N_7919,N_6871,N_6206);
xnor U7920 (N_7920,N_6754,N_6666);
xor U7921 (N_7921,N_6156,N_6878);
nor U7922 (N_7922,N_6818,N_6514);
xnor U7923 (N_7923,N_6887,N_6884);
or U7924 (N_7924,N_6314,N_6386);
or U7925 (N_7925,N_6604,N_6652);
or U7926 (N_7926,N_6255,N_6206);
and U7927 (N_7927,N_6939,N_6686);
nor U7928 (N_7928,N_6163,N_6861);
and U7929 (N_7929,N_6841,N_6101);
xnor U7930 (N_7930,N_6481,N_6336);
xor U7931 (N_7931,N_6249,N_6453);
or U7932 (N_7932,N_6010,N_6595);
and U7933 (N_7933,N_6628,N_6476);
nand U7934 (N_7934,N_6154,N_6368);
and U7935 (N_7935,N_6868,N_6731);
nand U7936 (N_7936,N_6626,N_6283);
xor U7937 (N_7937,N_6343,N_6508);
nand U7938 (N_7938,N_6706,N_6891);
or U7939 (N_7939,N_6396,N_6638);
and U7940 (N_7940,N_6414,N_6702);
nand U7941 (N_7941,N_6495,N_6992);
nor U7942 (N_7942,N_6004,N_6743);
and U7943 (N_7943,N_6830,N_6613);
or U7944 (N_7944,N_6272,N_6782);
nand U7945 (N_7945,N_6584,N_6514);
nand U7946 (N_7946,N_6717,N_6791);
and U7947 (N_7947,N_6531,N_6677);
or U7948 (N_7948,N_6695,N_6802);
xnor U7949 (N_7949,N_6594,N_6247);
or U7950 (N_7950,N_6862,N_6244);
xor U7951 (N_7951,N_6779,N_6912);
nand U7952 (N_7952,N_6534,N_6091);
and U7953 (N_7953,N_6143,N_6530);
nand U7954 (N_7954,N_6031,N_6826);
nand U7955 (N_7955,N_6821,N_6705);
or U7956 (N_7956,N_6934,N_6005);
nand U7957 (N_7957,N_6461,N_6326);
nand U7958 (N_7958,N_6131,N_6673);
nor U7959 (N_7959,N_6843,N_6254);
or U7960 (N_7960,N_6754,N_6598);
nand U7961 (N_7961,N_6383,N_6773);
xnor U7962 (N_7962,N_6831,N_6837);
xor U7963 (N_7963,N_6231,N_6349);
and U7964 (N_7964,N_6047,N_6421);
or U7965 (N_7965,N_6516,N_6131);
or U7966 (N_7966,N_6037,N_6126);
nor U7967 (N_7967,N_6218,N_6878);
nor U7968 (N_7968,N_6733,N_6523);
nor U7969 (N_7969,N_6311,N_6978);
and U7970 (N_7970,N_6132,N_6629);
xnor U7971 (N_7971,N_6613,N_6258);
nor U7972 (N_7972,N_6489,N_6967);
and U7973 (N_7973,N_6145,N_6285);
or U7974 (N_7974,N_6844,N_6728);
nor U7975 (N_7975,N_6153,N_6577);
xor U7976 (N_7976,N_6241,N_6049);
nand U7977 (N_7977,N_6069,N_6922);
nor U7978 (N_7978,N_6570,N_6574);
and U7979 (N_7979,N_6699,N_6210);
nor U7980 (N_7980,N_6406,N_6090);
or U7981 (N_7981,N_6995,N_6158);
and U7982 (N_7982,N_6935,N_6517);
xor U7983 (N_7983,N_6770,N_6005);
nor U7984 (N_7984,N_6629,N_6548);
or U7985 (N_7985,N_6729,N_6408);
nand U7986 (N_7986,N_6820,N_6551);
or U7987 (N_7987,N_6734,N_6209);
and U7988 (N_7988,N_6835,N_6589);
or U7989 (N_7989,N_6794,N_6123);
or U7990 (N_7990,N_6441,N_6460);
nand U7991 (N_7991,N_6853,N_6655);
nand U7992 (N_7992,N_6927,N_6632);
xnor U7993 (N_7993,N_6422,N_6479);
xor U7994 (N_7994,N_6912,N_6214);
xnor U7995 (N_7995,N_6091,N_6386);
nand U7996 (N_7996,N_6090,N_6669);
and U7997 (N_7997,N_6042,N_6684);
nor U7998 (N_7998,N_6397,N_6014);
and U7999 (N_7999,N_6729,N_6464);
nand U8000 (N_8000,N_7670,N_7556);
xor U8001 (N_8001,N_7313,N_7405);
xor U8002 (N_8002,N_7363,N_7237);
nor U8003 (N_8003,N_7141,N_7090);
nand U8004 (N_8004,N_7402,N_7617);
xnor U8005 (N_8005,N_7020,N_7289);
nor U8006 (N_8006,N_7825,N_7856);
or U8007 (N_8007,N_7462,N_7377);
xnor U8008 (N_8008,N_7959,N_7282);
or U8009 (N_8009,N_7263,N_7126);
or U8010 (N_8010,N_7780,N_7474);
and U8011 (N_8011,N_7874,N_7470);
nand U8012 (N_8012,N_7445,N_7458);
or U8013 (N_8013,N_7213,N_7568);
xor U8014 (N_8014,N_7695,N_7937);
xnor U8015 (N_8015,N_7444,N_7156);
nor U8016 (N_8016,N_7211,N_7083);
and U8017 (N_8017,N_7492,N_7956);
and U8018 (N_8018,N_7654,N_7688);
nand U8019 (N_8019,N_7966,N_7390);
and U8020 (N_8020,N_7997,N_7231);
and U8021 (N_8021,N_7969,N_7953);
and U8022 (N_8022,N_7296,N_7400);
and U8023 (N_8023,N_7508,N_7901);
and U8024 (N_8024,N_7606,N_7435);
nand U8025 (N_8025,N_7732,N_7515);
nor U8026 (N_8026,N_7041,N_7702);
and U8027 (N_8027,N_7460,N_7424);
nand U8028 (N_8028,N_7721,N_7846);
nor U8029 (N_8029,N_7487,N_7802);
xnor U8030 (N_8030,N_7523,N_7095);
xor U8031 (N_8031,N_7549,N_7301);
nor U8032 (N_8032,N_7117,N_7295);
xor U8033 (N_8033,N_7504,N_7892);
nor U8034 (N_8034,N_7244,N_7833);
or U8035 (N_8035,N_7676,N_7713);
or U8036 (N_8036,N_7649,N_7246);
xor U8037 (N_8037,N_7984,N_7151);
and U8038 (N_8038,N_7740,N_7198);
nand U8039 (N_8039,N_7976,N_7148);
or U8040 (N_8040,N_7331,N_7757);
nand U8041 (N_8041,N_7316,N_7067);
nor U8042 (N_8042,N_7559,N_7728);
and U8043 (N_8043,N_7052,N_7514);
or U8044 (N_8044,N_7798,N_7337);
nor U8045 (N_8045,N_7340,N_7636);
xor U8046 (N_8046,N_7466,N_7533);
nand U8047 (N_8047,N_7043,N_7715);
and U8048 (N_8048,N_7483,N_7137);
nand U8049 (N_8049,N_7848,N_7541);
or U8050 (N_8050,N_7915,N_7480);
xnor U8051 (N_8051,N_7689,N_7123);
or U8052 (N_8052,N_7962,N_7146);
or U8053 (N_8053,N_7049,N_7397);
xor U8054 (N_8054,N_7609,N_7255);
and U8055 (N_8055,N_7871,N_7046);
nor U8056 (N_8056,N_7342,N_7744);
nand U8057 (N_8057,N_7132,N_7344);
nand U8058 (N_8058,N_7201,N_7196);
xnor U8059 (N_8059,N_7212,N_7382);
nand U8060 (N_8060,N_7028,N_7419);
nor U8061 (N_8061,N_7172,N_7527);
xnor U8062 (N_8062,N_7764,N_7298);
nand U8063 (N_8063,N_7546,N_7058);
nand U8064 (N_8064,N_7964,N_7567);
nor U8065 (N_8065,N_7980,N_7936);
xor U8066 (N_8066,N_7767,N_7598);
or U8067 (N_8067,N_7135,N_7094);
nor U8068 (N_8068,N_7248,N_7195);
nor U8069 (N_8069,N_7091,N_7938);
nor U8070 (N_8070,N_7776,N_7888);
or U8071 (N_8071,N_7588,N_7138);
nand U8072 (N_8072,N_7130,N_7849);
nor U8073 (N_8073,N_7597,N_7170);
or U8074 (N_8074,N_7017,N_7889);
or U8075 (N_8075,N_7529,N_7755);
nor U8076 (N_8076,N_7708,N_7481);
or U8077 (N_8077,N_7399,N_7409);
or U8078 (N_8078,N_7031,N_7312);
xor U8079 (N_8079,N_7810,N_7902);
and U8080 (N_8080,N_7147,N_7415);
xor U8081 (N_8081,N_7129,N_7169);
nor U8082 (N_8082,N_7866,N_7724);
and U8083 (N_8083,N_7693,N_7811);
and U8084 (N_8084,N_7574,N_7060);
or U8085 (N_8085,N_7791,N_7789);
or U8086 (N_8086,N_7729,N_7277);
and U8087 (N_8087,N_7751,N_7349);
nand U8088 (N_8088,N_7561,N_7394);
nor U8089 (N_8089,N_7421,N_7582);
nand U8090 (N_8090,N_7864,N_7291);
nor U8091 (N_8091,N_7845,N_7578);
nor U8092 (N_8092,N_7510,N_7726);
xnor U8093 (N_8093,N_7219,N_7249);
nor U8094 (N_8094,N_7865,N_7021);
nand U8095 (N_8095,N_7239,N_7253);
xnor U8096 (N_8096,N_7912,N_7827);
xnor U8097 (N_8097,N_7760,N_7684);
xnor U8098 (N_8098,N_7620,N_7573);
nor U8099 (N_8099,N_7085,N_7310);
and U8100 (N_8100,N_7018,N_7618);
nand U8101 (N_8101,N_7978,N_7600);
or U8102 (N_8102,N_7413,N_7572);
nor U8103 (N_8103,N_7704,N_7010);
xor U8104 (N_8104,N_7376,N_7380);
nor U8105 (N_8105,N_7233,N_7928);
nor U8106 (N_8106,N_7430,N_7283);
nor U8107 (N_8107,N_7711,N_7770);
and U8108 (N_8108,N_7302,N_7545);
and U8109 (N_8109,N_7725,N_7857);
or U8110 (N_8110,N_7869,N_7493);
xnor U8111 (N_8111,N_7131,N_7186);
or U8112 (N_8112,N_7700,N_7766);
and U8113 (N_8113,N_7334,N_7662);
and U8114 (N_8114,N_7524,N_7457);
nand U8115 (N_8115,N_7330,N_7660);
xor U8116 (N_8116,N_7823,N_7797);
and U8117 (N_8117,N_7242,N_7558);
and U8118 (N_8118,N_7035,N_7088);
nor U8119 (N_8119,N_7590,N_7995);
or U8120 (N_8120,N_7513,N_7407);
nor U8121 (N_8121,N_7024,N_7417);
and U8122 (N_8122,N_7652,N_7948);
and U8123 (N_8123,N_7033,N_7804);
nand U8124 (N_8124,N_7970,N_7648);
or U8125 (N_8125,N_7433,N_7179);
or U8126 (N_8126,N_7941,N_7384);
or U8127 (N_8127,N_7496,N_7175);
nor U8128 (N_8128,N_7084,N_7411);
and U8129 (N_8129,N_7484,N_7077);
nand U8130 (N_8130,N_7155,N_7476);
xor U8131 (N_8131,N_7465,N_7663);
and U8132 (N_8132,N_7197,N_7893);
or U8133 (N_8133,N_7981,N_7486);
xor U8134 (N_8134,N_7318,N_7949);
and U8135 (N_8135,N_7308,N_7473);
nand U8136 (N_8136,N_7455,N_7647);
or U8137 (N_8137,N_7200,N_7642);
nor U8138 (N_8138,N_7993,N_7038);
nand U8139 (N_8139,N_7029,N_7772);
and U8140 (N_8140,N_7322,N_7469);
nand U8141 (N_8141,N_7867,N_7734);
xnor U8142 (N_8142,N_7641,N_7595);
or U8143 (N_8143,N_7783,N_7338);
and U8144 (N_8144,N_7634,N_7743);
nor U8145 (N_8145,N_7579,N_7406);
and U8146 (N_8146,N_7064,N_7352);
nand U8147 (N_8147,N_7991,N_7139);
nand U8148 (N_8148,N_7843,N_7591);
xor U8149 (N_8149,N_7987,N_7459);
nor U8150 (N_8150,N_7208,N_7571);
or U8151 (N_8151,N_7273,N_7630);
nand U8152 (N_8152,N_7303,N_7436);
and U8153 (N_8153,N_7214,N_7485);
nor U8154 (N_8154,N_7015,N_7491);
xor U8155 (N_8155,N_7920,N_7203);
and U8156 (N_8156,N_7784,N_7069);
and U8157 (N_8157,N_7431,N_7076);
nand U8158 (N_8158,N_7860,N_7584);
or U8159 (N_8159,N_7005,N_7752);
or U8160 (N_8160,N_7961,N_7933);
nor U8161 (N_8161,N_7269,N_7055);
and U8162 (N_8162,N_7967,N_7828);
xor U8163 (N_8163,N_7144,N_7087);
nand U8164 (N_8164,N_7566,N_7741);
and U8165 (N_8165,N_7517,N_7625);
or U8166 (N_8166,N_7025,N_7383);
nor U8167 (N_8167,N_7438,N_7080);
xnor U8168 (N_8168,N_7528,N_7830);
and U8169 (N_8169,N_7503,N_7532);
xor U8170 (N_8170,N_7446,N_7222);
and U8171 (N_8171,N_7099,N_7610);
or U8172 (N_8172,N_7243,N_7542);
or U8173 (N_8173,N_7391,N_7899);
and U8174 (N_8174,N_7191,N_7145);
nor U8175 (N_8175,N_7008,N_7121);
or U8176 (N_8176,N_7906,N_7794);
xor U8177 (N_8177,N_7822,N_7051);
nor U8178 (N_8178,N_7931,N_7265);
or U8179 (N_8179,N_7544,N_7717);
and U8180 (N_8180,N_7821,N_7168);
and U8181 (N_8181,N_7034,N_7300);
or U8182 (N_8182,N_7422,N_7389);
nand U8183 (N_8183,N_7293,N_7986);
or U8184 (N_8184,N_7036,N_7963);
xor U8185 (N_8185,N_7166,N_7521);
nand U8186 (N_8186,N_7073,N_7664);
or U8187 (N_8187,N_7304,N_7488);
and U8188 (N_8188,N_7329,N_7401);
nor U8189 (N_8189,N_7615,N_7100);
nand U8190 (N_8190,N_7266,N_7489);
xor U8191 (N_8191,N_7482,N_7586);
or U8192 (N_8192,N_7898,N_7163);
nand U8193 (N_8193,N_7593,N_7682);
and U8194 (N_8194,N_7079,N_7911);
nor U8195 (N_8195,N_7926,N_7796);
xor U8196 (N_8196,N_7287,N_7536);
xnor U8197 (N_8197,N_7669,N_7305);
or U8198 (N_8198,N_7506,N_7368);
nand U8199 (N_8199,N_7426,N_7104);
or U8200 (N_8200,N_7378,N_7650);
and U8201 (N_8201,N_7498,N_7461);
nand U8202 (N_8202,N_7687,N_7120);
and U8203 (N_8203,N_7012,N_7737);
and U8204 (N_8204,N_7102,N_7904);
nand U8205 (N_8205,N_7745,N_7782);
nor U8206 (N_8206,N_7690,N_7180);
or U8207 (N_8207,N_7016,N_7133);
xnor U8208 (N_8208,N_7171,N_7861);
nand U8209 (N_8209,N_7703,N_7799);
and U8210 (N_8210,N_7350,N_7030);
nor U8211 (N_8211,N_7883,N_7440);
nand U8212 (N_8212,N_7994,N_7839);
and U8213 (N_8213,N_7501,N_7307);
and U8214 (N_8214,N_7762,N_7379);
nor U8215 (N_8215,N_7373,N_7317);
nand U8216 (N_8216,N_7940,N_7537);
nand U8217 (N_8217,N_7164,N_7686);
nand U8218 (N_8218,N_7639,N_7245);
and U8219 (N_8219,N_7332,N_7640);
nor U8220 (N_8220,N_7339,N_7074);
nand U8221 (N_8221,N_7592,N_7907);
xnor U8222 (N_8222,N_7071,N_7599);
and U8223 (N_8223,N_7927,N_7885);
or U8224 (N_8224,N_7369,N_7321);
nand U8225 (N_8225,N_7916,N_7806);
xor U8226 (N_8226,N_7900,N_7443);
nor U8227 (N_8227,N_7587,N_7831);
or U8228 (N_8228,N_7779,N_7177);
or U8229 (N_8229,N_7112,N_7832);
or U8230 (N_8230,N_7173,N_7555);
xor U8231 (N_8231,N_7190,N_7290);
or U8232 (N_8232,N_7955,N_7738);
nand U8233 (N_8233,N_7047,N_7333);
nand U8234 (N_8234,N_7420,N_7607);
nand U8235 (N_8235,N_7730,N_7013);
nand U8236 (N_8236,N_7479,N_7224);
and U8237 (N_8237,N_7306,N_7735);
or U8238 (N_8238,N_7563,N_7124);
nand U8239 (N_8239,N_7756,N_7136);
nor U8240 (N_8240,N_7814,N_7925);
nor U8241 (N_8241,N_7011,N_7775);
nand U8242 (N_8242,N_7062,N_7720);
xnor U8243 (N_8243,N_7467,N_7001);
xor U8244 (N_8244,N_7410,N_7056);
nor U8245 (N_8245,N_7267,N_7275);
xor U8246 (N_8246,N_7884,N_7603);
nor U8247 (N_8247,N_7829,N_7006);
or U8248 (N_8248,N_7229,N_7979);
nand U8249 (N_8249,N_7909,N_7736);
and U8250 (N_8250,N_7705,N_7348);
nand U8251 (N_8251,N_7990,N_7753);
nand U8252 (N_8252,N_7111,N_7449);
xor U8253 (N_8253,N_7009,N_7646);
nor U8254 (N_8254,N_7014,N_7223);
nand U8255 (N_8255,N_7539,N_7217);
nor U8256 (N_8256,N_7623,N_7260);
and U8257 (N_8257,N_7773,N_7434);
nor U8258 (N_8258,N_7922,N_7143);
nand U8259 (N_8259,N_7027,N_7820);
and U8260 (N_8260,N_7627,N_7026);
or U8261 (N_8261,N_7657,N_7818);
nor U8262 (N_8262,N_7577,N_7477);
nand U8263 (N_8263,N_7428,N_7771);
and U8264 (N_8264,N_7985,N_7256);
and U8265 (N_8265,N_7154,N_7543);
nor U8266 (N_8266,N_7530,N_7022);
nand U8267 (N_8267,N_7604,N_7280);
or U8268 (N_8268,N_7699,N_7800);
xor U8269 (N_8269,N_7975,N_7750);
nor U8270 (N_8270,N_7873,N_7957);
and U8271 (N_8271,N_7838,N_7731);
and U8272 (N_8272,N_7215,N_7355);
xnor U8273 (N_8273,N_7210,N_7945);
nor U8274 (N_8274,N_7161,N_7370);
nor U8275 (N_8275,N_7809,N_7692);
nor U8276 (N_8276,N_7793,N_7089);
or U8277 (N_8277,N_7505,N_7075);
nand U8278 (N_8278,N_7863,N_7204);
and U8279 (N_8279,N_7323,N_7661);
nor U8280 (N_8280,N_7418,N_7362);
xor U8281 (N_8281,N_7176,N_7932);
xor U8282 (N_8282,N_7950,N_7218);
or U8283 (N_8283,N_7552,N_7836);
nand U8284 (N_8284,N_7464,N_7951);
nor U8285 (N_8285,N_7557,N_7398);
and U8286 (N_8286,N_7656,N_7965);
and U8287 (N_8287,N_7097,N_7781);
xnor U8288 (N_8288,N_7448,N_7605);
nand U8289 (N_8289,N_7816,N_7375);
and U8290 (N_8290,N_7947,N_7628);
and U8291 (N_8291,N_7502,N_7292);
and U8292 (N_8292,N_7934,N_7683);
nand U8293 (N_8293,N_7238,N_7134);
xnor U8294 (N_8294,N_7790,N_7093);
nor U8295 (N_8295,N_7727,N_7739);
xor U8296 (N_8296,N_7507,N_7518);
nor U8297 (N_8297,N_7319,N_7910);
nand U8298 (N_8298,N_7115,N_7003);
and U8299 (N_8299,N_7092,N_7105);
xor U8300 (N_8300,N_7989,N_7404);
or U8301 (N_8301,N_7879,N_7601);
and U8302 (N_8302,N_7706,N_7946);
xor U8303 (N_8303,N_7812,N_7271);
nor U8304 (N_8304,N_7803,N_7054);
and U8305 (N_8305,N_7416,N_7758);
nor U8306 (N_8306,N_7761,N_7070);
nor U8307 (N_8307,N_7387,N_7982);
xor U8308 (N_8308,N_7763,N_7570);
xor U8309 (N_8309,N_7251,N_7125);
and U8310 (N_8310,N_7905,N_7877);
nor U8311 (N_8311,N_7429,N_7974);
or U8312 (N_8312,N_7913,N_7258);
or U8313 (N_8313,N_7667,N_7769);
nand U8314 (N_8314,N_7374,N_7645);
and U8315 (N_8315,N_7759,N_7127);
xnor U8316 (N_8316,N_7685,N_7851);
xor U8317 (N_8317,N_7952,N_7712);
nor U8318 (N_8318,N_7841,N_7471);
or U8319 (N_8319,N_7019,N_7635);
nand U8320 (N_8320,N_7516,N_7061);
nand U8321 (N_8321,N_7644,N_7631);
xnor U8322 (N_8322,N_7678,N_7351);
nand U8323 (N_8323,N_7673,N_7209);
nand U8324 (N_8324,N_7924,N_7569);
nor U8325 (N_8325,N_7897,N_7452);
and U8326 (N_8326,N_7903,N_7629);
nor U8327 (N_8327,N_7853,N_7813);
xor U8328 (N_8328,N_7999,N_7608);
nand U8329 (N_8329,N_7942,N_7531);
nor U8330 (N_8330,N_7519,N_7122);
and U8331 (N_8331,N_7847,N_7472);
or U8332 (N_8332,N_7327,N_7891);
or U8333 (N_8333,N_7110,N_7972);
nor U8334 (N_8334,N_7425,N_7066);
or U8335 (N_8335,N_7819,N_7257);
xor U8336 (N_8336,N_7497,N_7614);
nand U8337 (N_8337,N_7228,N_7261);
xnor U8338 (N_8338,N_7065,N_7185);
xor U8339 (N_8339,N_7451,N_7594);
and U8340 (N_8340,N_7000,N_7886);
xnor U8341 (N_8341,N_7653,N_7633);
and U8342 (N_8342,N_7553,N_7494);
xnor U8343 (N_8343,N_7106,N_7184);
nand U8344 (N_8344,N_7944,N_7254);
or U8345 (N_8345,N_7032,N_7002);
or U8346 (N_8346,N_7921,N_7742);
nand U8347 (N_8347,N_7098,N_7336);
nor U8348 (N_8348,N_7427,N_7063);
and U8349 (N_8349,N_7288,N_7453);
or U8350 (N_8350,N_7580,N_7414);
nand U8351 (N_8351,N_7500,N_7341);
xor U8352 (N_8352,N_7632,N_7326);
nor U8353 (N_8353,N_7534,N_7815);
or U8354 (N_8354,N_7658,N_7621);
nand U8355 (N_8355,N_7565,N_7252);
and U8356 (N_8356,N_7973,N_7718);
xnor U8357 (N_8357,N_7081,N_7675);
nand U8358 (N_8358,N_7103,N_7835);
xnor U8359 (N_8359,N_7680,N_7314);
xor U8360 (N_8360,N_7040,N_7343);
nand U8361 (N_8361,N_7826,N_7876);
and U8362 (N_8362,N_7114,N_7643);
and U8363 (N_8363,N_7596,N_7939);
nor U8364 (N_8364,N_7194,N_7923);
nor U8365 (N_8365,N_7881,N_7988);
nor U8366 (N_8366,N_7240,N_7777);
and U8367 (N_8367,N_7236,N_7392);
and U8368 (N_8368,N_7691,N_7917);
nand U8369 (N_8369,N_7181,N_7954);
xnor U8370 (N_8370,N_7311,N_7616);
nor U8371 (N_8371,N_7585,N_7749);
xnor U8372 (N_8372,N_7395,N_7178);
and U8373 (N_8373,N_7057,N_7371);
or U8374 (N_8374,N_7309,N_7150);
and U8375 (N_8375,N_7862,N_7535);
xor U8376 (N_8376,N_7345,N_7442);
and U8377 (N_8377,N_7361,N_7059);
nand U8378 (N_8378,N_7393,N_7837);
xor U8379 (N_8379,N_7241,N_7206);
xor U8380 (N_8380,N_7441,N_7358);
and U8381 (N_8381,N_7581,N_7808);
xor U8382 (N_8382,N_7250,N_7220);
or U8383 (N_8383,N_7612,N_7285);
and U8384 (N_8384,N_7281,N_7372);
nor U8385 (N_8385,N_7423,N_7844);
nand U8386 (N_8386,N_7205,N_7840);
nand U8387 (N_8387,N_7674,N_7589);
or U8388 (N_8388,N_7672,N_7562);
nor U8389 (N_8389,N_7247,N_7787);
nor U8390 (N_8390,N_7272,N_7677);
and U8391 (N_8391,N_7914,N_7895);
or U8392 (N_8392,N_7335,N_7386);
nand U8393 (N_8393,N_7068,N_7512);
and U8394 (N_8394,N_7560,N_7929);
xor U8395 (N_8395,N_7174,N_7786);
or U8396 (N_8396,N_7403,N_7230);
or U8397 (N_8397,N_7575,N_7276);
xor U8398 (N_8398,N_7454,N_7490);
or U8399 (N_8399,N_7520,N_7671);
xor U8400 (N_8400,N_7943,N_7325);
nor U8401 (N_8401,N_7119,N_7227);
nand U8402 (N_8402,N_7364,N_7037);
and U8403 (N_8403,N_7187,N_7044);
nand U8404 (N_8404,N_7048,N_7096);
and U8405 (N_8405,N_7365,N_7709);
nand U8406 (N_8406,N_7522,N_7234);
xnor U8407 (N_8407,N_7188,N_7360);
and U8408 (N_8408,N_7270,N_7412);
and U8409 (N_8409,N_7294,N_7665);
nand U8410 (N_8410,N_7202,N_7896);
nor U8411 (N_8411,N_7128,N_7004);
xor U8412 (N_8412,N_7153,N_7919);
nor U8413 (N_8413,N_7118,N_7659);
xor U8414 (N_8414,N_7437,N_7538);
nand U8415 (N_8415,N_7158,N_7698);
nand U8416 (N_8416,N_7754,N_7447);
nand U8417 (N_8417,N_7697,N_7651);
xnor U8418 (N_8418,N_7199,N_7347);
or U8419 (N_8419,N_7045,N_7540);
and U8420 (N_8420,N_7554,N_7747);
nor U8421 (N_8421,N_7259,N_7805);
or U8422 (N_8422,N_7996,N_7408);
nor U8423 (N_8423,N_7279,N_7116);
nor U8424 (N_8424,N_7226,N_7576);
nand U8425 (N_8425,N_7284,N_7550);
nor U8426 (N_8426,N_7381,N_7101);
and U8427 (N_8427,N_7894,N_7007);
nor U8428 (N_8428,N_7694,N_7511);
or U8429 (N_8429,N_7960,N_7908);
and U8430 (N_8430,N_7707,N_7880);
nor U8431 (N_8431,N_7346,N_7774);
nand U8432 (N_8432,N_7320,N_7824);
nand U8433 (N_8433,N_7792,N_7189);
nor U8434 (N_8434,N_7354,N_7357);
and U8435 (N_8435,N_7870,N_7324);
nand U8436 (N_8436,N_7152,N_7109);
and U8437 (N_8437,N_7450,N_7748);
nand U8438 (N_8438,N_7149,N_7958);
xnor U8439 (N_8439,N_7525,N_7859);
nor U8440 (N_8440,N_7278,N_7082);
xnor U8441 (N_8441,N_7432,N_7356);
nand U8442 (N_8442,N_7722,N_7834);
nand U8443 (N_8443,N_7286,N_7983);
and U8444 (N_8444,N_7353,N_7638);
nor U8445 (N_8445,N_7785,N_7078);
or U8446 (N_8446,N_7053,N_7162);
xor U8447 (N_8447,N_7396,N_7701);
nand U8448 (N_8448,N_7872,N_7232);
nor U8449 (N_8449,N_7714,N_7626);
nor U8450 (N_8450,N_7681,N_7666);
nand U8451 (N_8451,N_7850,N_7930);
or U8452 (N_8452,N_7733,N_7868);
or U8453 (N_8453,N_7548,N_7315);
or U8454 (N_8454,N_7108,N_7468);
xnor U8455 (N_8455,N_7622,N_7042);
nor U8456 (N_8456,N_7366,N_7768);
and U8457 (N_8457,N_7359,N_7268);
and U8458 (N_8458,N_7696,N_7890);
nand U8459 (N_8459,N_7182,N_7439);
nand U8460 (N_8460,N_7328,N_7723);
and U8461 (N_8461,N_7478,N_7107);
or U8462 (N_8462,N_7264,N_7655);
nor U8463 (N_8463,N_7039,N_7216);
nand U8464 (N_8464,N_7637,N_7475);
and U8465 (N_8465,N_7801,N_7619);
xor U8466 (N_8466,N_7971,N_7817);
nor U8467 (N_8467,N_7274,N_7854);
and U8468 (N_8468,N_7778,N_7388);
nand U8469 (N_8469,N_7142,N_7602);
nor U8470 (N_8470,N_7297,N_7719);
xnor U8471 (N_8471,N_7193,N_7262);
or U8472 (N_8472,N_7852,N_7564);
xor U8473 (N_8473,N_7977,N_7140);
and U8474 (N_8474,N_7795,N_7160);
and U8475 (N_8475,N_7998,N_7716);
nor U8476 (N_8476,N_7807,N_7157);
nor U8477 (N_8477,N_7385,N_7765);
xnor U8478 (N_8478,N_7526,N_7456);
nor U8479 (N_8479,N_7499,N_7495);
nand U8480 (N_8480,N_7882,N_7842);
or U8481 (N_8481,N_7624,N_7551);
and U8482 (N_8482,N_7935,N_7072);
xor U8483 (N_8483,N_7710,N_7611);
xnor U8484 (N_8484,N_7583,N_7235);
xnor U8485 (N_8485,N_7050,N_7547);
xnor U8486 (N_8486,N_7299,N_7225);
or U8487 (N_8487,N_7221,N_7679);
xor U8488 (N_8488,N_7746,N_7509);
nor U8489 (N_8489,N_7183,N_7165);
xnor U8490 (N_8490,N_7463,N_7613);
nor U8491 (N_8491,N_7918,N_7023);
or U8492 (N_8492,N_7668,N_7858);
xor U8493 (N_8493,N_7207,N_7992);
xnor U8494 (N_8494,N_7887,N_7788);
xnor U8495 (N_8495,N_7878,N_7113);
or U8496 (N_8496,N_7367,N_7159);
nor U8497 (N_8497,N_7086,N_7968);
or U8498 (N_8498,N_7875,N_7855);
nor U8499 (N_8499,N_7167,N_7192);
or U8500 (N_8500,N_7171,N_7829);
or U8501 (N_8501,N_7772,N_7847);
nand U8502 (N_8502,N_7951,N_7613);
nor U8503 (N_8503,N_7547,N_7563);
or U8504 (N_8504,N_7371,N_7582);
and U8505 (N_8505,N_7193,N_7382);
nand U8506 (N_8506,N_7329,N_7945);
nand U8507 (N_8507,N_7867,N_7192);
or U8508 (N_8508,N_7407,N_7830);
and U8509 (N_8509,N_7308,N_7581);
nor U8510 (N_8510,N_7512,N_7746);
xor U8511 (N_8511,N_7517,N_7887);
nor U8512 (N_8512,N_7074,N_7134);
nor U8513 (N_8513,N_7940,N_7418);
nand U8514 (N_8514,N_7292,N_7826);
or U8515 (N_8515,N_7884,N_7520);
nand U8516 (N_8516,N_7385,N_7733);
xnor U8517 (N_8517,N_7545,N_7736);
nand U8518 (N_8518,N_7359,N_7495);
nand U8519 (N_8519,N_7109,N_7657);
nor U8520 (N_8520,N_7614,N_7139);
nor U8521 (N_8521,N_7038,N_7330);
and U8522 (N_8522,N_7619,N_7626);
nand U8523 (N_8523,N_7605,N_7678);
nand U8524 (N_8524,N_7560,N_7358);
nor U8525 (N_8525,N_7352,N_7167);
and U8526 (N_8526,N_7500,N_7961);
nand U8527 (N_8527,N_7492,N_7596);
nor U8528 (N_8528,N_7814,N_7615);
nand U8529 (N_8529,N_7107,N_7936);
nor U8530 (N_8530,N_7480,N_7376);
nor U8531 (N_8531,N_7189,N_7672);
and U8532 (N_8532,N_7038,N_7249);
nor U8533 (N_8533,N_7237,N_7037);
xor U8534 (N_8534,N_7750,N_7337);
or U8535 (N_8535,N_7228,N_7442);
or U8536 (N_8536,N_7583,N_7108);
nand U8537 (N_8537,N_7404,N_7126);
and U8538 (N_8538,N_7000,N_7040);
or U8539 (N_8539,N_7900,N_7983);
or U8540 (N_8540,N_7208,N_7578);
xor U8541 (N_8541,N_7803,N_7180);
nor U8542 (N_8542,N_7099,N_7843);
or U8543 (N_8543,N_7657,N_7193);
nand U8544 (N_8544,N_7570,N_7105);
nor U8545 (N_8545,N_7569,N_7814);
and U8546 (N_8546,N_7562,N_7401);
nand U8547 (N_8547,N_7387,N_7520);
nor U8548 (N_8548,N_7348,N_7794);
nor U8549 (N_8549,N_7192,N_7256);
and U8550 (N_8550,N_7182,N_7662);
nor U8551 (N_8551,N_7336,N_7173);
xnor U8552 (N_8552,N_7214,N_7274);
xnor U8553 (N_8553,N_7542,N_7865);
and U8554 (N_8554,N_7318,N_7488);
or U8555 (N_8555,N_7185,N_7504);
nor U8556 (N_8556,N_7855,N_7318);
nand U8557 (N_8557,N_7254,N_7463);
nor U8558 (N_8558,N_7172,N_7331);
and U8559 (N_8559,N_7684,N_7624);
xnor U8560 (N_8560,N_7506,N_7489);
nand U8561 (N_8561,N_7994,N_7731);
xnor U8562 (N_8562,N_7675,N_7640);
nor U8563 (N_8563,N_7799,N_7716);
nand U8564 (N_8564,N_7856,N_7807);
xor U8565 (N_8565,N_7807,N_7046);
and U8566 (N_8566,N_7500,N_7762);
and U8567 (N_8567,N_7754,N_7522);
xor U8568 (N_8568,N_7836,N_7590);
nor U8569 (N_8569,N_7190,N_7695);
xor U8570 (N_8570,N_7854,N_7486);
nand U8571 (N_8571,N_7222,N_7183);
nand U8572 (N_8572,N_7927,N_7272);
nor U8573 (N_8573,N_7427,N_7955);
and U8574 (N_8574,N_7355,N_7975);
xor U8575 (N_8575,N_7949,N_7461);
nor U8576 (N_8576,N_7938,N_7944);
nor U8577 (N_8577,N_7893,N_7120);
and U8578 (N_8578,N_7269,N_7263);
nand U8579 (N_8579,N_7438,N_7985);
and U8580 (N_8580,N_7936,N_7287);
nor U8581 (N_8581,N_7945,N_7272);
and U8582 (N_8582,N_7315,N_7196);
nand U8583 (N_8583,N_7794,N_7755);
xnor U8584 (N_8584,N_7409,N_7242);
or U8585 (N_8585,N_7975,N_7572);
xor U8586 (N_8586,N_7121,N_7670);
nor U8587 (N_8587,N_7367,N_7418);
xor U8588 (N_8588,N_7382,N_7605);
or U8589 (N_8589,N_7082,N_7457);
and U8590 (N_8590,N_7187,N_7612);
xor U8591 (N_8591,N_7025,N_7701);
xnor U8592 (N_8592,N_7525,N_7800);
nor U8593 (N_8593,N_7053,N_7832);
or U8594 (N_8594,N_7393,N_7142);
or U8595 (N_8595,N_7924,N_7361);
nand U8596 (N_8596,N_7764,N_7851);
xor U8597 (N_8597,N_7805,N_7865);
nand U8598 (N_8598,N_7525,N_7223);
nor U8599 (N_8599,N_7791,N_7118);
and U8600 (N_8600,N_7955,N_7681);
and U8601 (N_8601,N_7881,N_7779);
and U8602 (N_8602,N_7078,N_7108);
xor U8603 (N_8603,N_7846,N_7980);
nor U8604 (N_8604,N_7489,N_7981);
nor U8605 (N_8605,N_7584,N_7742);
or U8606 (N_8606,N_7538,N_7921);
and U8607 (N_8607,N_7584,N_7808);
and U8608 (N_8608,N_7491,N_7030);
nor U8609 (N_8609,N_7644,N_7821);
or U8610 (N_8610,N_7880,N_7511);
nand U8611 (N_8611,N_7360,N_7243);
nor U8612 (N_8612,N_7002,N_7641);
xor U8613 (N_8613,N_7845,N_7126);
nor U8614 (N_8614,N_7891,N_7905);
xnor U8615 (N_8615,N_7696,N_7856);
xor U8616 (N_8616,N_7006,N_7387);
or U8617 (N_8617,N_7206,N_7980);
and U8618 (N_8618,N_7879,N_7998);
or U8619 (N_8619,N_7725,N_7353);
xor U8620 (N_8620,N_7231,N_7565);
and U8621 (N_8621,N_7197,N_7544);
nand U8622 (N_8622,N_7855,N_7813);
and U8623 (N_8623,N_7216,N_7842);
nor U8624 (N_8624,N_7632,N_7066);
and U8625 (N_8625,N_7104,N_7422);
or U8626 (N_8626,N_7668,N_7874);
and U8627 (N_8627,N_7967,N_7787);
nand U8628 (N_8628,N_7852,N_7837);
nand U8629 (N_8629,N_7819,N_7404);
and U8630 (N_8630,N_7622,N_7477);
xnor U8631 (N_8631,N_7050,N_7920);
nor U8632 (N_8632,N_7512,N_7884);
xor U8633 (N_8633,N_7613,N_7662);
or U8634 (N_8634,N_7214,N_7311);
nor U8635 (N_8635,N_7909,N_7856);
nor U8636 (N_8636,N_7315,N_7195);
or U8637 (N_8637,N_7613,N_7785);
and U8638 (N_8638,N_7172,N_7732);
nor U8639 (N_8639,N_7588,N_7037);
nand U8640 (N_8640,N_7582,N_7394);
nand U8641 (N_8641,N_7888,N_7751);
and U8642 (N_8642,N_7503,N_7940);
nand U8643 (N_8643,N_7004,N_7827);
xnor U8644 (N_8644,N_7299,N_7423);
or U8645 (N_8645,N_7700,N_7399);
nor U8646 (N_8646,N_7082,N_7106);
nor U8647 (N_8647,N_7227,N_7995);
and U8648 (N_8648,N_7275,N_7602);
nand U8649 (N_8649,N_7697,N_7063);
and U8650 (N_8650,N_7339,N_7661);
nor U8651 (N_8651,N_7508,N_7137);
xnor U8652 (N_8652,N_7854,N_7066);
nor U8653 (N_8653,N_7918,N_7434);
nand U8654 (N_8654,N_7199,N_7742);
and U8655 (N_8655,N_7378,N_7433);
xnor U8656 (N_8656,N_7690,N_7276);
nand U8657 (N_8657,N_7972,N_7874);
nand U8658 (N_8658,N_7755,N_7245);
nand U8659 (N_8659,N_7342,N_7968);
and U8660 (N_8660,N_7302,N_7906);
or U8661 (N_8661,N_7408,N_7166);
nor U8662 (N_8662,N_7601,N_7155);
nand U8663 (N_8663,N_7851,N_7780);
nand U8664 (N_8664,N_7035,N_7415);
and U8665 (N_8665,N_7545,N_7338);
nor U8666 (N_8666,N_7159,N_7218);
nor U8667 (N_8667,N_7023,N_7103);
and U8668 (N_8668,N_7828,N_7604);
nand U8669 (N_8669,N_7465,N_7715);
or U8670 (N_8670,N_7133,N_7269);
xor U8671 (N_8671,N_7893,N_7732);
or U8672 (N_8672,N_7103,N_7306);
or U8673 (N_8673,N_7635,N_7761);
or U8674 (N_8674,N_7796,N_7399);
nand U8675 (N_8675,N_7311,N_7154);
nor U8676 (N_8676,N_7133,N_7274);
xor U8677 (N_8677,N_7035,N_7680);
nor U8678 (N_8678,N_7422,N_7482);
or U8679 (N_8679,N_7293,N_7855);
xnor U8680 (N_8680,N_7262,N_7582);
nand U8681 (N_8681,N_7300,N_7543);
nand U8682 (N_8682,N_7341,N_7268);
or U8683 (N_8683,N_7151,N_7357);
and U8684 (N_8684,N_7788,N_7067);
nor U8685 (N_8685,N_7168,N_7715);
or U8686 (N_8686,N_7469,N_7057);
xor U8687 (N_8687,N_7902,N_7820);
or U8688 (N_8688,N_7306,N_7934);
xnor U8689 (N_8689,N_7435,N_7497);
or U8690 (N_8690,N_7933,N_7661);
nand U8691 (N_8691,N_7736,N_7009);
xnor U8692 (N_8692,N_7307,N_7143);
and U8693 (N_8693,N_7283,N_7056);
nand U8694 (N_8694,N_7451,N_7252);
xnor U8695 (N_8695,N_7350,N_7789);
xor U8696 (N_8696,N_7993,N_7404);
nand U8697 (N_8697,N_7293,N_7512);
nand U8698 (N_8698,N_7172,N_7154);
nor U8699 (N_8699,N_7546,N_7179);
and U8700 (N_8700,N_7295,N_7263);
or U8701 (N_8701,N_7049,N_7911);
xor U8702 (N_8702,N_7369,N_7575);
nor U8703 (N_8703,N_7397,N_7028);
xnor U8704 (N_8704,N_7987,N_7206);
and U8705 (N_8705,N_7427,N_7765);
nor U8706 (N_8706,N_7154,N_7554);
nor U8707 (N_8707,N_7735,N_7410);
nand U8708 (N_8708,N_7943,N_7542);
xor U8709 (N_8709,N_7353,N_7380);
nand U8710 (N_8710,N_7713,N_7957);
xor U8711 (N_8711,N_7162,N_7287);
nor U8712 (N_8712,N_7063,N_7597);
xnor U8713 (N_8713,N_7203,N_7571);
nor U8714 (N_8714,N_7438,N_7389);
or U8715 (N_8715,N_7943,N_7831);
nand U8716 (N_8716,N_7308,N_7002);
nand U8717 (N_8717,N_7764,N_7758);
or U8718 (N_8718,N_7894,N_7316);
nor U8719 (N_8719,N_7867,N_7104);
and U8720 (N_8720,N_7067,N_7660);
nor U8721 (N_8721,N_7734,N_7401);
nor U8722 (N_8722,N_7594,N_7046);
or U8723 (N_8723,N_7695,N_7162);
nand U8724 (N_8724,N_7395,N_7066);
nand U8725 (N_8725,N_7069,N_7736);
nor U8726 (N_8726,N_7815,N_7419);
nor U8727 (N_8727,N_7742,N_7013);
and U8728 (N_8728,N_7373,N_7724);
xor U8729 (N_8729,N_7946,N_7750);
and U8730 (N_8730,N_7855,N_7610);
or U8731 (N_8731,N_7019,N_7630);
or U8732 (N_8732,N_7602,N_7022);
nor U8733 (N_8733,N_7288,N_7501);
nor U8734 (N_8734,N_7799,N_7532);
nand U8735 (N_8735,N_7377,N_7557);
and U8736 (N_8736,N_7575,N_7361);
nor U8737 (N_8737,N_7222,N_7376);
and U8738 (N_8738,N_7143,N_7442);
xnor U8739 (N_8739,N_7518,N_7957);
or U8740 (N_8740,N_7878,N_7455);
nand U8741 (N_8741,N_7231,N_7226);
nor U8742 (N_8742,N_7703,N_7760);
nand U8743 (N_8743,N_7944,N_7253);
and U8744 (N_8744,N_7617,N_7862);
xnor U8745 (N_8745,N_7484,N_7973);
nor U8746 (N_8746,N_7507,N_7891);
and U8747 (N_8747,N_7488,N_7737);
and U8748 (N_8748,N_7549,N_7272);
and U8749 (N_8749,N_7052,N_7678);
nor U8750 (N_8750,N_7143,N_7568);
xor U8751 (N_8751,N_7142,N_7388);
nand U8752 (N_8752,N_7791,N_7715);
xor U8753 (N_8753,N_7168,N_7409);
xnor U8754 (N_8754,N_7674,N_7099);
or U8755 (N_8755,N_7599,N_7312);
or U8756 (N_8756,N_7934,N_7077);
xnor U8757 (N_8757,N_7047,N_7653);
nor U8758 (N_8758,N_7007,N_7969);
xnor U8759 (N_8759,N_7436,N_7604);
xor U8760 (N_8760,N_7505,N_7759);
and U8761 (N_8761,N_7063,N_7367);
nor U8762 (N_8762,N_7508,N_7811);
and U8763 (N_8763,N_7083,N_7199);
xor U8764 (N_8764,N_7980,N_7755);
or U8765 (N_8765,N_7362,N_7402);
and U8766 (N_8766,N_7851,N_7150);
or U8767 (N_8767,N_7753,N_7915);
or U8768 (N_8768,N_7636,N_7661);
nand U8769 (N_8769,N_7281,N_7767);
xnor U8770 (N_8770,N_7334,N_7712);
and U8771 (N_8771,N_7935,N_7950);
nand U8772 (N_8772,N_7561,N_7916);
and U8773 (N_8773,N_7784,N_7385);
and U8774 (N_8774,N_7526,N_7162);
or U8775 (N_8775,N_7475,N_7540);
nand U8776 (N_8776,N_7081,N_7013);
and U8777 (N_8777,N_7340,N_7188);
or U8778 (N_8778,N_7082,N_7412);
and U8779 (N_8779,N_7171,N_7428);
nor U8780 (N_8780,N_7734,N_7350);
nand U8781 (N_8781,N_7677,N_7820);
or U8782 (N_8782,N_7365,N_7964);
or U8783 (N_8783,N_7959,N_7119);
and U8784 (N_8784,N_7681,N_7404);
nor U8785 (N_8785,N_7750,N_7614);
nand U8786 (N_8786,N_7174,N_7600);
nand U8787 (N_8787,N_7266,N_7613);
and U8788 (N_8788,N_7910,N_7483);
xnor U8789 (N_8789,N_7889,N_7255);
and U8790 (N_8790,N_7509,N_7716);
xor U8791 (N_8791,N_7207,N_7512);
or U8792 (N_8792,N_7710,N_7901);
nor U8793 (N_8793,N_7831,N_7242);
xor U8794 (N_8794,N_7712,N_7637);
xnor U8795 (N_8795,N_7123,N_7096);
xnor U8796 (N_8796,N_7549,N_7153);
or U8797 (N_8797,N_7165,N_7964);
nand U8798 (N_8798,N_7186,N_7098);
nor U8799 (N_8799,N_7893,N_7551);
and U8800 (N_8800,N_7595,N_7318);
nand U8801 (N_8801,N_7003,N_7568);
xor U8802 (N_8802,N_7404,N_7973);
and U8803 (N_8803,N_7888,N_7551);
and U8804 (N_8804,N_7035,N_7870);
or U8805 (N_8805,N_7948,N_7649);
xnor U8806 (N_8806,N_7490,N_7234);
or U8807 (N_8807,N_7588,N_7715);
and U8808 (N_8808,N_7620,N_7382);
xor U8809 (N_8809,N_7770,N_7307);
xnor U8810 (N_8810,N_7082,N_7453);
xor U8811 (N_8811,N_7002,N_7411);
xor U8812 (N_8812,N_7514,N_7925);
nor U8813 (N_8813,N_7535,N_7203);
and U8814 (N_8814,N_7982,N_7131);
xor U8815 (N_8815,N_7435,N_7659);
xor U8816 (N_8816,N_7919,N_7721);
or U8817 (N_8817,N_7180,N_7885);
xnor U8818 (N_8818,N_7569,N_7473);
nor U8819 (N_8819,N_7778,N_7089);
nand U8820 (N_8820,N_7241,N_7968);
xor U8821 (N_8821,N_7058,N_7368);
nand U8822 (N_8822,N_7680,N_7483);
or U8823 (N_8823,N_7322,N_7578);
nand U8824 (N_8824,N_7559,N_7448);
nand U8825 (N_8825,N_7424,N_7774);
xnor U8826 (N_8826,N_7620,N_7907);
and U8827 (N_8827,N_7785,N_7164);
nand U8828 (N_8828,N_7295,N_7897);
nand U8829 (N_8829,N_7423,N_7463);
nand U8830 (N_8830,N_7448,N_7326);
and U8831 (N_8831,N_7129,N_7788);
or U8832 (N_8832,N_7268,N_7391);
and U8833 (N_8833,N_7729,N_7711);
nor U8834 (N_8834,N_7297,N_7456);
or U8835 (N_8835,N_7464,N_7298);
nor U8836 (N_8836,N_7150,N_7533);
or U8837 (N_8837,N_7407,N_7360);
and U8838 (N_8838,N_7635,N_7506);
and U8839 (N_8839,N_7566,N_7304);
and U8840 (N_8840,N_7394,N_7475);
xor U8841 (N_8841,N_7491,N_7314);
and U8842 (N_8842,N_7708,N_7869);
nor U8843 (N_8843,N_7961,N_7025);
nand U8844 (N_8844,N_7038,N_7863);
nor U8845 (N_8845,N_7047,N_7963);
or U8846 (N_8846,N_7308,N_7788);
nor U8847 (N_8847,N_7984,N_7664);
or U8848 (N_8848,N_7548,N_7757);
nand U8849 (N_8849,N_7687,N_7916);
xnor U8850 (N_8850,N_7130,N_7710);
xor U8851 (N_8851,N_7401,N_7216);
nor U8852 (N_8852,N_7724,N_7245);
xnor U8853 (N_8853,N_7909,N_7207);
and U8854 (N_8854,N_7628,N_7295);
nand U8855 (N_8855,N_7822,N_7385);
and U8856 (N_8856,N_7667,N_7145);
nand U8857 (N_8857,N_7145,N_7564);
xnor U8858 (N_8858,N_7182,N_7392);
nand U8859 (N_8859,N_7955,N_7321);
xor U8860 (N_8860,N_7976,N_7972);
xnor U8861 (N_8861,N_7528,N_7145);
xor U8862 (N_8862,N_7415,N_7123);
xor U8863 (N_8863,N_7340,N_7189);
xor U8864 (N_8864,N_7840,N_7936);
xor U8865 (N_8865,N_7547,N_7496);
nor U8866 (N_8866,N_7603,N_7112);
nand U8867 (N_8867,N_7802,N_7053);
nor U8868 (N_8868,N_7379,N_7698);
and U8869 (N_8869,N_7364,N_7385);
nor U8870 (N_8870,N_7285,N_7100);
or U8871 (N_8871,N_7218,N_7888);
xor U8872 (N_8872,N_7011,N_7666);
or U8873 (N_8873,N_7691,N_7799);
or U8874 (N_8874,N_7642,N_7381);
and U8875 (N_8875,N_7474,N_7716);
nor U8876 (N_8876,N_7672,N_7356);
or U8877 (N_8877,N_7189,N_7611);
nand U8878 (N_8878,N_7801,N_7359);
or U8879 (N_8879,N_7447,N_7668);
and U8880 (N_8880,N_7744,N_7474);
and U8881 (N_8881,N_7088,N_7929);
nand U8882 (N_8882,N_7207,N_7940);
or U8883 (N_8883,N_7691,N_7905);
or U8884 (N_8884,N_7647,N_7038);
nand U8885 (N_8885,N_7807,N_7965);
and U8886 (N_8886,N_7118,N_7335);
xor U8887 (N_8887,N_7912,N_7231);
xnor U8888 (N_8888,N_7443,N_7647);
nand U8889 (N_8889,N_7244,N_7543);
and U8890 (N_8890,N_7108,N_7345);
and U8891 (N_8891,N_7694,N_7836);
nor U8892 (N_8892,N_7277,N_7407);
nor U8893 (N_8893,N_7259,N_7505);
nor U8894 (N_8894,N_7165,N_7128);
xor U8895 (N_8895,N_7703,N_7029);
and U8896 (N_8896,N_7305,N_7932);
nor U8897 (N_8897,N_7989,N_7900);
nand U8898 (N_8898,N_7579,N_7678);
or U8899 (N_8899,N_7678,N_7248);
xor U8900 (N_8900,N_7263,N_7046);
or U8901 (N_8901,N_7358,N_7114);
xnor U8902 (N_8902,N_7758,N_7763);
nand U8903 (N_8903,N_7590,N_7253);
xor U8904 (N_8904,N_7181,N_7243);
nor U8905 (N_8905,N_7366,N_7688);
xnor U8906 (N_8906,N_7831,N_7073);
or U8907 (N_8907,N_7697,N_7947);
nand U8908 (N_8908,N_7763,N_7675);
and U8909 (N_8909,N_7024,N_7892);
and U8910 (N_8910,N_7138,N_7037);
xnor U8911 (N_8911,N_7591,N_7230);
xor U8912 (N_8912,N_7275,N_7389);
nor U8913 (N_8913,N_7268,N_7810);
nand U8914 (N_8914,N_7419,N_7486);
or U8915 (N_8915,N_7732,N_7699);
nand U8916 (N_8916,N_7301,N_7953);
and U8917 (N_8917,N_7541,N_7564);
xnor U8918 (N_8918,N_7103,N_7430);
or U8919 (N_8919,N_7079,N_7659);
or U8920 (N_8920,N_7514,N_7475);
xnor U8921 (N_8921,N_7665,N_7126);
xor U8922 (N_8922,N_7322,N_7145);
or U8923 (N_8923,N_7774,N_7136);
or U8924 (N_8924,N_7556,N_7723);
and U8925 (N_8925,N_7359,N_7478);
and U8926 (N_8926,N_7274,N_7437);
and U8927 (N_8927,N_7596,N_7472);
or U8928 (N_8928,N_7345,N_7058);
nor U8929 (N_8929,N_7062,N_7188);
and U8930 (N_8930,N_7689,N_7820);
xnor U8931 (N_8931,N_7226,N_7973);
xnor U8932 (N_8932,N_7684,N_7160);
or U8933 (N_8933,N_7050,N_7803);
nand U8934 (N_8934,N_7866,N_7919);
nand U8935 (N_8935,N_7162,N_7692);
nand U8936 (N_8936,N_7176,N_7620);
and U8937 (N_8937,N_7329,N_7599);
nand U8938 (N_8938,N_7076,N_7091);
or U8939 (N_8939,N_7948,N_7289);
and U8940 (N_8940,N_7854,N_7964);
nor U8941 (N_8941,N_7879,N_7643);
nand U8942 (N_8942,N_7419,N_7078);
nand U8943 (N_8943,N_7843,N_7520);
or U8944 (N_8944,N_7112,N_7775);
nand U8945 (N_8945,N_7275,N_7996);
nor U8946 (N_8946,N_7396,N_7183);
or U8947 (N_8947,N_7113,N_7666);
nand U8948 (N_8948,N_7097,N_7798);
and U8949 (N_8949,N_7082,N_7848);
or U8950 (N_8950,N_7359,N_7729);
nand U8951 (N_8951,N_7407,N_7401);
nand U8952 (N_8952,N_7683,N_7951);
nand U8953 (N_8953,N_7092,N_7836);
or U8954 (N_8954,N_7897,N_7389);
xor U8955 (N_8955,N_7611,N_7851);
nand U8956 (N_8956,N_7615,N_7166);
nor U8957 (N_8957,N_7446,N_7507);
nand U8958 (N_8958,N_7846,N_7824);
nand U8959 (N_8959,N_7467,N_7893);
nand U8960 (N_8960,N_7886,N_7594);
nand U8961 (N_8961,N_7748,N_7482);
and U8962 (N_8962,N_7641,N_7142);
or U8963 (N_8963,N_7942,N_7423);
xor U8964 (N_8964,N_7236,N_7285);
and U8965 (N_8965,N_7514,N_7031);
nor U8966 (N_8966,N_7658,N_7949);
and U8967 (N_8967,N_7547,N_7044);
and U8968 (N_8968,N_7024,N_7361);
or U8969 (N_8969,N_7326,N_7833);
or U8970 (N_8970,N_7750,N_7938);
nand U8971 (N_8971,N_7735,N_7101);
xor U8972 (N_8972,N_7050,N_7942);
or U8973 (N_8973,N_7920,N_7157);
nand U8974 (N_8974,N_7608,N_7158);
nor U8975 (N_8975,N_7463,N_7931);
and U8976 (N_8976,N_7007,N_7385);
and U8977 (N_8977,N_7746,N_7913);
nor U8978 (N_8978,N_7929,N_7383);
xor U8979 (N_8979,N_7062,N_7508);
nor U8980 (N_8980,N_7312,N_7731);
or U8981 (N_8981,N_7097,N_7890);
or U8982 (N_8982,N_7342,N_7759);
nand U8983 (N_8983,N_7844,N_7329);
and U8984 (N_8984,N_7816,N_7429);
xor U8985 (N_8985,N_7280,N_7563);
xnor U8986 (N_8986,N_7020,N_7531);
or U8987 (N_8987,N_7461,N_7673);
nand U8988 (N_8988,N_7558,N_7888);
nor U8989 (N_8989,N_7465,N_7085);
and U8990 (N_8990,N_7357,N_7401);
nand U8991 (N_8991,N_7003,N_7645);
nor U8992 (N_8992,N_7538,N_7351);
nand U8993 (N_8993,N_7098,N_7434);
and U8994 (N_8994,N_7165,N_7762);
nand U8995 (N_8995,N_7829,N_7261);
xnor U8996 (N_8996,N_7716,N_7208);
nor U8997 (N_8997,N_7682,N_7657);
nor U8998 (N_8998,N_7547,N_7091);
and U8999 (N_8999,N_7017,N_7792);
xnor U9000 (N_9000,N_8420,N_8691);
nand U9001 (N_9001,N_8537,N_8692);
nor U9002 (N_9002,N_8595,N_8511);
or U9003 (N_9003,N_8489,N_8084);
xor U9004 (N_9004,N_8619,N_8293);
and U9005 (N_9005,N_8437,N_8988);
nor U9006 (N_9006,N_8247,N_8947);
xnor U9007 (N_9007,N_8972,N_8181);
and U9008 (N_9008,N_8409,N_8251);
nand U9009 (N_9009,N_8456,N_8562);
or U9010 (N_9010,N_8516,N_8810);
xnor U9011 (N_9011,N_8989,N_8336);
nor U9012 (N_9012,N_8152,N_8695);
or U9013 (N_9013,N_8945,N_8993);
nand U9014 (N_9014,N_8739,N_8746);
xnor U9015 (N_9015,N_8799,N_8067);
or U9016 (N_9016,N_8760,N_8559);
xor U9017 (N_9017,N_8736,N_8218);
or U9018 (N_9018,N_8494,N_8359);
nand U9019 (N_9019,N_8350,N_8341);
nand U9020 (N_9020,N_8541,N_8415);
and U9021 (N_9021,N_8862,N_8464);
nand U9022 (N_9022,N_8672,N_8698);
and U9023 (N_9023,N_8256,N_8486);
nor U9024 (N_9024,N_8786,N_8727);
nand U9025 (N_9025,N_8314,N_8596);
or U9026 (N_9026,N_8008,N_8816);
and U9027 (N_9027,N_8054,N_8878);
or U9028 (N_9028,N_8805,N_8789);
or U9029 (N_9029,N_8927,N_8756);
nand U9030 (N_9030,N_8468,N_8822);
xor U9031 (N_9031,N_8368,N_8533);
and U9032 (N_9032,N_8479,N_8225);
nor U9033 (N_9033,N_8274,N_8768);
and U9034 (N_9034,N_8890,N_8189);
nand U9035 (N_9035,N_8792,N_8949);
or U9036 (N_9036,N_8030,N_8183);
or U9037 (N_9037,N_8105,N_8809);
nor U9038 (N_9038,N_8066,N_8371);
or U9039 (N_9039,N_8542,N_8262);
or U9040 (N_9040,N_8280,N_8459);
xor U9041 (N_9041,N_8657,N_8401);
and U9042 (N_9042,N_8029,N_8937);
nand U9043 (N_9043,N_8601,N_8644);
xor U9044 (N_9044,N_8905,N_8423);
or U9045 (N_9045,N_8519,N_8773);
nand U9046 (N_9046,N_8903,N_8419);
xnor U9047 (N_9047,N_8106,N_8669);
nor U9048 (N_9048,N_8223,N_8715);
xnor U9049 (N_9049,N_8729,N_8667);
xor U9050 (N_9050,N_8246,N_8813);
nand U9051 (N_9051,N_8734,N_8110);
xor U9052 (N_9052,N_8481,N_8238);
nor U9053 (N_9053,N_8748,N_8299);
nor U9054 (N_9054,N_8770,N_8317);
and U9055 (N_9055,N_8325,N_8831);
xnor U9056 (N_9056,N_8042,N_8414);
xor U9057 (N_9057,N_8759,N_8588);
or U9058 (N_9058,N_8380,N_8120);
and U9059 (N_9059,N_8342,N_8663);
and U9060 (N_9060,N_8351,N_8565);
xor U9061 (N_9061,N_8551,N_8723);
nand U9062 (N_9062,N_8528,N_8934);
xor U9063 (N_9063,N_8178,N_8005);
and U9064 (N_9064,N_8022,N_8870);
nand U9065 (N_9065,N_8610,N_8774);
and U9066 (N_9066,N_8801,N_8257);
or U9067 (N_9067,N_8943,N_8113);
xor U9068 (N_9068,N_8253,N_8664);
xor U9069 (N_9069,N_8567,N_8035);
or U9070 (N_9070,N_8885,N_8048);
nor U9071 (N_9071,N_8072,N_8974);
and U9072 (N_9072,N_8910,N_8007);
nand U9073 (N_9073,N_8370,N_8365);
and U9074 (N_9074,N_8848,N_8031);
nor U9075 (N_9075,N_8026,N_8276);
xor U9076 (N_9076,N_8226,N_8662);
or U9077 (N_9077,N_8891,N_8170);
and U9078 (N_9078,N_8666,N_8568);
nor U9079 (N_9079,N_8821,N_8548);
nand U9080 (N_9080,N_8694,N_8016);
nor U9081 (N_9081,N_8612,N_8659);
or U9082 (N_9082,N_8130,N_8515);
nor U9083 (N_9083,N_8697,N_8177);
nand U9084 (N_9084,N_8332,N_8781);
or U9085 (N_9085,N_8097,N_8722);
xor U9086 (N_9086,N_8023,N_8269);
nor U9087 (N_9087,N_8076,N_8389);
nand U9088 (N_9088,N_8726,N_8064);
or U9089 (N_9089,N_8677,N_8779);
xnor U9090 (N_9090,N_8605,N_8263);
or U9091 (N_9091,N_8093,N_8840);
nand U9092 (N_9092,N_8791,N_8638);
or U9093 (N_9093,N_8776,N_8160);
nor U9094 (N_9094,N_8764,N_8439);
xor U9095 (N_9095,N_8915,N_8518);
nand U9096 (N_9096,N_8699,N_8900);
and U9097 (N_9097,N_8616,N_8538);
xor U9098 (N_9098,N_8711,N_8545);
or U9099 (N_9099,N_8604,N_8680);
nand U9100 (N_9100,N_8967,N_8963);
or U9101 (N_9101,N_8115,N_8427);
nor U9102 (N_9102,N_8408,N_8167);
nor U9103 (N_9103,N_8772,N_8717);
xnor U9104 (N_9104,N_8268,N_8324);
nor U9105 (N_9105,N_8544,N_8080);
nand U9106 (N_9106,N_8558,N_8941);
xor U9107 (N_9107,N_8200,N_8847);
xor U9108 (N_9108,N_8245,N_8311);
nor U9109 (N_9109,N_8556,N_8313);
and U9110 (N_9110,N_8444,N_8654);
or U9111 (N_9111,N_8865,N_8671);
xnor U9112 (N_9112,N_8385,N_8758);
xor U9113 (N_9113,N_8534,N_8109);
or U9114 (N_9114,N_8156,N_8880);
xnor U9115 (N_9115,N_8693,N_8432);
xnor U9116 (N_9116,N_8169,N_8948);
nor U9117 (N_9117,N_8001,N_8362);
or U9118 (N_9118,N_8686,N_8407);
xor U9119 (N_9119,N_8954,N_8524);
xor U9120 (N_9120,N_8172,N_8241);
and U9121 (N_9121,N_8622,N_8175);
and U9122 (N_9122,N_8580,N_8841);
and U9123 (N_9123,N_8212,N_8339);
nor U9124 (N_9124,N_8309,N_8114);
and U9125 (N_9125,N_8955,N_8122);
or U9126 (N_9126,N_8176,N_8390);
and U9127 (N_9127,N_8613,N_8981);
nand U9128 (N_9128,N_8942,N_8850);
xor U9129 (N_9129,N_8496,N_8208);
nand U9130 (N_9130,N_8907,N_8400);
nand U9131 (N_9131,N_8784,N_8828);
nand U9132 (N_9132,N_8911,N_8397);
and U9133 (N_9133,N_8431,N_8306);
xor U9134 (N_9134,N_8917,N_8171);
and U9135 (N_9135,N_8630,N_8069);
nor U9136 (N_9136,N_8146,N_8002);
or U9137 (N_9137,N_8194,N_8244);
or U9138 (N_9138,N_8625,N_8995);
xor U9139 (N_9139,N_8836,N_8300);
or U9140 (N_9140,N_8835,N_8908);
and U9141 (N_9141,N_8535,N_8021);
xor U9142 (N_9142,N_8575,N_8688);
nor U9143 (N_9143,N_8852,N_8259);
nor U9144 (N_9144,N_8708,N_8966);
nor U9145 (N_9145,N_8895,N_8233);
nor U9146 (N_9146,N_8099,N_8886);
nor U9147 (N_9147,N_8036,N_8203);
or U9148 (N_9148,N_8254,N_8976);
xnor U9149 (N_9149,N_8471,N_8034);
xor U9150 (N_9150,N_8552,N_8980);
xor U9151 (N_9151,N_8374,N_8320);
nand U9152 (N_9152,N_8348,N_8861);
and U9153 (N_9153,N_8844,N_8956);
or U9154 (N_9154,N_8703,N_8503);
and U9155 (N_9155,N_8015,N_8714);
and U9156 (N_9156,N_8383,N_8379);
and U9157 (N_9157,N_8939,N_8373);
xnor U9158 (N_9158,N_8394,N_8367);
or U9159 (N_9159,N_8217,N_8833);
xnor U9160 (N_9160,N_8514,N_8572);
or U9161 (N_9161,N_8433,N_8352);
and U9162 (N_9162,N_8088,N_8461);
or U9163 (N_9163,N_8495,N_8117);
nor U9164 (N_9164,N_8800,N_8512);
nand U9165 (N_9165,N_8957,N_8803);
or U9166 (N_9166,N_8752,N_8827);
nor U9167 (N_9167,N_8062,N_8651);
and U9168 (N_9168,N_8017,N_8057);
xor U9169 (N_9169,N_8829,N_8837);
nor U9170 (N_9170,N_8295,N_8070);
nand U9171 (N_9171,N_8402,N_8707);
nor U9172 (N_9172,N_8125,N_8753);
and U9173 (N_9173,N_8571,N_8308);
and U9174 (N_9174,N_8787,N_8484);
nor U9175 (N_9175,N_8843,N_8049);
and U9176 (N_9176,N_8287,N_8331);
nand U9177 (N_9177,N_8230,N_8975);
and U9178 (N_9178,N_8090,N_8586);
nor U9179 (N_9179,N_8215,N_8962);
and U9180 (N_9180,N_8174,N_8267);
nand U9181 (N_9181,N_8446,N_8819);
nand U9182 (N_9182,N_8141,N_8162);
nand U9183 (N_9183,N_8815,N_8425);
nor U9184 (N_9184,N_8634,N_8749);
nor U9185 (N_9185,N_8889,N_8576);
or U9186 (N_9186,N_8386,N_8121);
nor U9187 (N_9187,N_8343,N_8333);
or U9188 (N_9188,N_8702,N_8600);
or U9189 (N_9189,N_8643,N_8670);
nand U9190 (N_9190,N_8817,N_8553);
or U9191 (N_9191,N_8112,N_8597);
nand U9192 (N_9192,N_8849,N_8303);
xnor U9193 (N_9193,N_8363,N_8701);
nand U9194 (N_9194,N_8297,N_8492);
and U9195 (N_9195,N_8056,N_8639);
xor U9196 (N_9196,N_8607,N_8086);
nand U9197 (N_9197,N_8145,N_8261);
xor U9198 (N_9198,N_8690,N_8148);
xnor U9199 (N_9199,N_8138,N_8123);
nor U9200 (N_9200,N_8032,N_8965);
xnor U9201 (N_9201,N_8830,N_8679);
nor U9202 (N_9202,N_8258,N_8735);
nor U9203 (N_9203,N_8220,N_8582);
or U9204 (N_9204,N_8611,N_8971);
or U9205 (N_9205,N_8434,N_8075);
nand U9206 (N_9206,N_8617,N_8335);
xnor U9207 (N_9207,N_8978,N_8139);
and U9208 (N_9208,N_8040,N_8116);
nand U9209 (N_9209,N_8999,N_8323);
xor U9210 (N_9210,N_8609,N_8281);
and U9211 (N_9211,N_8924,N_8997);
xnor U9212 (N_9212,N_8450,N_8569);
xor U9213 (N_9213,N_8260,N_8872);
or U9214 (N_9214,N_8033,N_8213);
or U9215 (N_9215,N_8807,N_8777);
or U9216 (N_9216,N_8732,N_8232);
xnor U9217 (N_9217,N_8825,N_8140);
nand U9218 (N_9218,N_8540,N_8718);
nand U9219 (N_9219,N_8650,N_8501);
xnor U9220 (N_9220,N_8143,N_8583);
nor U9221 (N_9221,N_8738,N_8430);
xor U9222 (N_9222,N_8024,N_8104);
xor U9223 (N_9223,N_8655,N_8472);
nand U9224 (N_9224,N_8590,N_8046);
nand U9225 (N_9225,N_8500,N_8724);
xor U9226 (N_9226,N_8922,N_8593);
nand U9227 (N_9227,N_8010,N_8990);
nor U9228 (N_9228,N_8762,N_8951);
nand U9229 (N_9229,N_8202,N_8188);
or U9230 (N_9230,N_8598,N_8504);
or U9231 (N_9231,N_8710,N_8337);
nand U9232 (N_9232,N_8207,N_8881);
nor U9233 (N_9233,N_8411,N_8636);
or U9234 (N_9234,N_8438,N_8242);
xnor U9235 (N_9235,N_8823,N_8563);
and U9236 (N_9236,N_8790,N_8887);
and U9237 (N_9237,N_8307,N_8893);
and U9238 (N_9238,N_8755,N_8222);
xnor U9239 (N_9239,N_8623,N_8834);
nand U9240 (N_9240,N_8883,N_8094);
nand U9241 (N_9241,N_8526,N_8410);
nor U9242 (N_9242,N_8587,N_8027);
nor U9243 (N_9243,N_8648,N_8868);
xor U9244 (N_9244,N_8909,N_8846);
nand U9245 (N_9245,N_8190,N_8913);
xnor U9246 (N_9246,N_8327,N_8505);
or U9247 (N_9247,N_8053,N_8465);
xnor U9248 (N_9248,N_8019,N_8463);
nand U9249 (N_9249,N_8592,N_8424);
nor U9250 (N_9250,N_8038,N_8478);
or U9251 (N_9251,N_8025,N_8912);
or U9252 (N_9252,N_8522,N_8382);
nor U9253 (N_9253,N_8529,N_8457);
or U9254 (N_9254,N_8950,N_8318);
xor U9255 (N_9255,N_8338,N_8520);
and U9256 (N_9256,N_8133,N_8628);
or U9257 (N_9257,N_8931,N_8857);
and U9258 (N_9258,N_8445,N_8231);
or U9259 (N_9259,N_8531,N_8393);
and U9260 (N_9260,N_8043,N_8473);
and U9261 (N_9261,N_8863,N_8606);
xor U9262 (N_9262,N_8731,N_8301);
xnor U9263 (N_9263,N_8986,N_8157);
and U9264 (N_9264,N_8635,N_8854);
nor U9265 (N_9265,N_8992,N_8150);
and U9266 (N_9266,N_8673,N_8742);
nand U9267 (N_9267,N_8646,N_8682);
nor U9268 (N_9268,N_8391,N_8166);
or U9269 (N_9269,N_8416,N_8077);
and U9270 (N_9270,N_8685,N_8761);
nor U9271 (N_9271,N_8921,N_8375);
xor U9272 (N_9272,N_8132,N_8395);
nand U9273 (N_9273,N_8302,N_8665);
or U9274 (N_9274,N_8159,N_8369);
and U9275 (N_9275,N_8376,N_8289);
xnor U9276 (N_9276,N_8647,N_8959);
and U9277 (N_9277,N_8403,N_8346);
or U9278 (N_9278,N_8977,N_8720);
and U9279 (N_9279,N_8279,N_8284);
xor U9280 (N_9280,N_8916,N_8938);
and U9281 (N_9281,N_8871,N_8728);
nor U9282 (N_9282,N_8441,N_8102);
nor U9283 (N_9283,N_8914,N_8205);
or U9284 (N_9284,N_8340,N_8278);
and U9285 (N_9285,N_8737,N_8454);
xor U9286 (N_9286,N_8249,N_8165);
and U9287 (N_9287,N_8899,N_8923);
xor U9288 (N_9288,N_8083,N_8058);
and U9289 (N_9289,N_8901,N_8319);
nand U9290 (N_9290,N_8984,N_8633);
nand U9291 (N_9291,N_8357,N_8897);
xor U9292 (N_9292,N_8812,N_8599);
nand U9293 (N_9293,N_8209,N_8998);
nand U9294 (N_9294,N_8328,N_8676);
nand U9295 (N_9295,N_8460,N_8081);
and U9296 (N_9296,N_8620,N_8063);
or U9297 (N_9297,N_8970,N_8780);
xnor U9298 (N_9298,N_8013,N_8079);
or U9299 (N_9299,N_8050,N_8523);
and U9300 (N_9300,N_8709,N_8876);
nor U9301 (N_9301,N_8316,N_8969);
nand U9302 (N_9302,N_8168,N_8733);
nand U9303 (N_9303,N_8119,N_8092);
nor U9304 (N_9304,N_8510,N_8101);
nor U9305 (N_9305,N_8964,N_8012);
xor U9306 (N_9306,N_8236,N_8820);
nor U9307 (N_9307,N_8991,N_8184);
nand U9308 (N_9308,N_8902,N_8808);
and U9309 (N_9309,N_8273,N_8788);
or U9310 (N_9310,N_8838,N_8201);
or U9311 (N_9311,N_8045,N_8930);
and U9312 (N_9312,N_8239,N_8277);
nor U9313 (N_9313,N_8640,N_8087);
nand U9314 (N_9314,N_8888,N_8765);
or U9315 (N_9315,N_8705,N_8904);
nand U9316 (N_9316,N_8377,N_8491);
and U9317 (N_9317,N_8802,N_8487);
nor U9318 (N_9318,N_8627,N_8591);
nor U9319 (N_9319,N_8906,N_8614);
xnor U9320 (N_9320,N_8960,N_8873);
and U9321 (N_9321,N_8096,N_8349);
or U9322 (N_9322,N_8994,N_8811);
and U9323 (N_9323,N_8187,N_8874);
xor U9324 (N_9324,N_8126,N_8272);
and U9325 (N_9325,N_8039,N_8806);
xor U9326 (N_9326,N_8594,N_8014);
nor U9327 (N_9327,N_8882,N_8769);
and U9328 (N_9328,N_8451,N_8228);
nand U9329 (N_9329,N_8474,N_8961);
or U9330 (N_9330,N_8982,N_8356);
and U9331 (N_9331,N_8933,N_8388);
and U9332 (N_9332,N_8507,N_8645);
or U9333 (N_9333,N_8626,N_8154);
xnor U9334 (N_9334,N_8771,N_8129);
xnor U9335 (N_9335,N_8161,N_8783);
and U9336 (N_9336,N_8378,N_8291);
nand U9337 (N_9337,N_8135,N_8928);
xnor U9338 (N_9338,N_8716,N_8180);
nor U9339 (N_9339,N_8361,N_8447);
nand U9340 (N_9340,N_8859,N_8482);
or U9341 (N_9341,N_8134,N_8649);
or U9342 (N_9342,N_8216,N_8265);
xor U9343 (N_9343,N_8442,N_8637);
xnor U9344 (N_9344,N_8243,N_8095);
xnor U9345 (N_9345,N_8443,N_8118);
xor U9346 (N_9346,N_8641,N_8869);
nand U9347 (N_9347,N_8860,N_8071);
nand U9348 (N_9348,N_8577,N_8615);
nand U9349 (N_9349,N_8334,N_8429);
nand U9350 (N_9350,N_8877,N_8108);
nand U9351 (N_9351,N_8539,N_8824);
and U9352 (N_9352,N_8074,N_8757);
xor U9353 (N_9353,N_8275,N_8689);
or U9354 (N_9354,N_8674,N_8100);
nor U9355 (N_9355,N_8107,N_8124);
and U9356 (N_9356,N_8153,N_8098);
xor U9357 (N_9357,N_8557,N_8458);
xor U9358 (N_9358,N_8681,N_8462);
nand U9359 (N_9359,N_8197,N_8555);
xnor U9360 (N_9360,N_8149,N_8164);
and U9361 (N_9361,N_8059,N_8315);
and U9362 (N_9362,N_8578,N_8968);
nand U9363 (N_9363,N_8364,N_8485);
nor U9364 (N_9364,N_8078,N_8103);
nand U9365 (N_9365,N_8192,N_8574);
nand U9366 (N_9366,N_8550,N_8521);
nor U9367 (N_9367,N_8179,N_8292);
or U9368 (N_9368,N_8782,N_8743);
xor U9369 (N_9369,N_8683,N_8128);
and U9370 (N_9370,N_8000,N_8751);
or U9371 (N_9371,N_8678,N_8173);
and U9372 (N_9372,N_8793,N_8296);
or U9373 (N_9373,N_8499,N_8706);
nand U9374 (N_9374,N_8428,N_8490);
xnor U9375 (N_9375,N_8051,N_8421);
and U9376 (N_9376,N_8345,N_8795);
and U9377 (N_9377,N_8532,N_8266);
nor U9378 (N_9378,N_8741,N_8147);
nand U9379 (N_9379,N_8011,N_8513);
xor U9380 (N_9380,N_8794,N_8853);
and U9381 (N_9381,N_8264,N_8435);
nor U9382 (N_9382,N_8740,N_8744);
or U9383 (N_9383,N_8498,N_8856);
nor U9384 (N_9384,N_8250,N_8286);
xnor U9385 (N_9385,N_8898,N_8252);
nand U9386 (N_9386,N_8452,N_8422);
or U9387 (N_9387,N_8285,N_8466);
xor U9388 (N_9388,N_8525,N_8312);
and U9389 (N_9389,N_8399,N_8842);
or U9390 (N_9390,N_8061,N_8925);
or U9391 (N_9391,N_8602,N_8355);
and U9392 (N_9392,N_8426,N_8055);
or U9393 (N_9393,N_8003,N_8142);
and U9394 (N_9394,N_8564,N_8412);
or U9395 (N_9395,N_8204,N_8052);
and U9396 (N_9396,N_8656,N_8952);
or U9397 (N_9397,N_8298,N_8330);
xnor U9398 (N_9398,N_8725,N_8229);
nand U9399 (N_9399,N_8918,N_8721);
or U9400 (N_9400,N_8719,N_8091);
xor U9401 (N_9401,N_8483,N_8797);
or U9402 (N_9402,N_8477,N_8953);
xnor U9403 (N_9403,N_8546,N_8653);
nor U9404 (N_9404,N_8845,N_8798);
or U9405 (N_9405,N_8566,N_8502);
and U9406 (N_9406,N_8560,N_8237);
nand U9407 (N_9407,N_8449,N_8163);
nand U9408 (N_9408,N_8660,N_8182);
xor U9409 (N_9409,N_8618,N_8932);
nand U9410 (N_9410,N_8406,N_8384);
and U9411 (N_9411,N_8785,N_8006);
nand U9412 (N_9412,N_8321,N_8547);
nand U9413 (N_9413,N_8329,N_8508);
or U9414 (N_9414,N_8561,N_8398);
or U9415 (N_9415,N_8089,N_8754);
nor U9416 (N_9416,N_8936,N_8979);
and U9417 (N_9417,N_8527,N_8894);
nand U9418 (N_9418,N_8476,N_8004);
or U9419 (N_9419,N_8632,N_8127);
nor U9420 (N_9420,N_8417,N_8044);
or U9421 (N_9421,N_8131,N_8704);
xor U9422 (N_9422,N_8326,N_8283);
xnor U9423 (N_9423,N_8366,N_8235);
nor U9424 (N_9424,N_8985,N_8448);
xor U9425 (N_9425,N_8983,N_8470);
xor U9426 (N_9426,N_8440,N_8658);
xor U9427 (N_9427,N_8158,N_8661);
nor U9428 (N_9428,N_8944,N_8987);
and U9429 (N_9429,N_8920,N_8288);
nor U9430 (N_9430,N_8018,N_8536);
xnor U9431 (N_9431,N_8778,N_8271);
nor U9432 (N_9432,N_8467,N_8210);
nor U9433 (N_9433,N_8041,N_8191);
or U9434 (N_9434,N_8310,N_8137);
and U9435 (N_9435,N_8712,N_8506);
or U9436 (N_9436,N_8573,N_8392);
nand U9437 (N_9437,N_8198,N_8136);
or U9438 (N_9438,N_8240,N_8480);
or U9439 (N_9439,N_8193,N_8347);
nand U9440 (N_9440,N_8747,N_8696);
nor U9441 (N_9441,N_8372,N_8405);
and U9442 (N_9442,N_8413,N_8832);
or U9443 (N_9443,N_8621,N_8608);
nor U9444 (N_9444,N_8589,N_8322);
and U9445 (N_9445,N_8344,N_8579);
xor U9446 (N_9446,N_8935,N_8219);
nor U9447 (N_9447,N_8270,N_8196);
nand U9448 (N_9448,N_8224,N_8855);
and U9449 (N_9449,N_8554,N_8530);
or U9450 (N_9450,N_8629,N_8745);
xnor U9451 (N_9451,N_8826,N_8814);
and U9452 (N_9452,N_8221,N_8214);
and U9453 (N_9453,N_8353,N_8497);
nand U9454 (N_9454,N_8867,N_8713);
xnor U9455 (N_9455,N_8294,N_8996);
nor U9456 (N_9456,N_8926,N_8584);
nor U9457 (N_9457,N_8199,N_8940);
and U9458 (N_9458,N_8396,N_8603);
nand U9459 (N_9459,N_8700,N_8892);
or U9460 (N_9460,N_8082,N_8581);
and U9461 (N_9461,N_8958,N_8453);
or U9462 (N_9462,N_8804,N_8155);
xnor U9463 (N_9463,N_8549,N_8585);
nand U9464 (N_9464,N_8475,N_8509);
or U9465 (N_9465,N_8767,N_8304);
and U9466 (N_9466,N_8360,N_8766);
nand U9467 (N_9467,N_8851,N_8436);
nor U9468 (N_9468,N_8684,N_8642);
nand U9469 (N_9469,N_8730,N_8687);
xnor U9470 (N_9470,N_8517,N_8068);
xnor U9471 (N_9471,N_8144,N_8875);
or U9472 (N_9472,N_8282,N_8488);
nand U9473 (N_9473,N_8919,N_8186);
nor U9474 (N_9474,N_8206,N_8884);
xnor U9475 (N_9475,N_8866,N_8211);
nor U9476 (N_9476,N_8195,N_8354);
xnor U9477 (N_9477,N_8185,N_8037);
or U9478 (N_9478,N_8418,N_8020);
nand U9479 (N_9479,N_8065,N_8358);
and U9480 (N_9480,N_8111,N_8085);
and U9481 (N_9481,N_8028,N_8290);
nand U9482 (N_9482,N_8631,N_8763);
xor U9483 (N_9483,N_8543,N_8675);
and U9484 (N_9484,N_8929,N_8404);
or U9485 (N_9485,N_8227,N_8818);
nand U9486 (N_9486,N_8896,N_8387);
nand U9487 (N_9487,N_8864,N_8009);
or U9488 (N_9488,N_8624,N_8469);
xor U9489 (N_9489,N_8248,N_8652);
nor U9490 (N_9490,N_8570,N_8946);
nor U9491 (N_9491,N_8858,N_8879);
xor U9492 (N_9492,N_8305,N_8839);
and U9493 (N_9493,N_8775,N_8750);
and U9494 (N_9494,N_8796,N_8151);
nand U9495 (N_9495,N_8060,N_8234);
and U9496 (N_9496,N_8493,N_8455);
and U9497 (N_9497,N_8255,N_8073);
nor U9498 (N_9498,N_8973,N_8381);
and U9499 (N_9499,N_8047,N_8668);
xnor U9500 (N_9500,N_8204,N_8943);
xor U9501 (N_9501,N_8186,N_8103);
or U9502 (N_9502,N_8390,N_8382);
nand U9503 (N_9503,N_8424,N_8239);
or U9504 (N_9504,N_8996,N_8853);
nand U9505 (N_9505,N_8075,N_8236);
nor U9506 (N_9506,N_8217,N_8944);
or U9507 (N_9507,N_8392,N_8613);
nand U9508 (N_9508,N_8313,N_8335);
nand U9509 (N_9509,N_8664,N_8530);
nand U9510 (N_9510,N_8903,N_8388);
or U9511 (N_9511,N_8326,N_8822);
xor U9512 (N_9512,N_8098,N_8923);
xnor U9513 (N_9513,N_8610,N_8522);
and U9514 (N_9514,N_8517,N_8496);
nand U9515 (N_9515,N_8686,N_8142);
and U9516 (N_9516,N_8050,N_8608);
xor U9517 (N_9517,N_8930,N_8545);
xnor U9518 (N_9518,N_8708,N_8681);
nand U9519 (N_9519,N_8754,N_8939);
and U9520 (N_9520,N_8787,N_8278);
nand U9521 (N_9521,N_8200,N_8294);
nor U9522 (N_9522,N_8132,N_8716);
or U9523 (N_9523,N_8242,N_8628);
nand U9524 (N_9524,N_8339,N_8804);
and U9525 (N_9525,N_8704,N_8284);
or U9526 (N_9526,N_8149,N_8962);
xnor U9527 (N_9527,N_8815,N_8231);
and U9528 (N_9528,N_8565,N_8441);
and U9529 (N_9529,N_8153,N_8108);
or U9530 (N_9530,N_8786,N_8655);
and U9531 (N_9531,N_8714,N_8487);
and U9532 (N_9532,N_8359,N_8791);
and U9533 (N_9533,N_8512,N_8769);
nand U9534 (N_9534,N_8200,N_8445);
nand U9535 (N_9535,N_8342,N_8660);
and U9536 (N_9536,N_8022,N_8676);
nand U9537 (N_9537,N_8179,N_8429);
and U9538 (N_9538,N_8629,N_8878);
nand U9539 (N_9539,N_8030,N_8658);
or U9540 (N_9540,N_8147,N_8802);
nand U9541 (N_9541,N_8304,N_8257);
xor U9542 (N_9542,N_8414,N_8468);
xnor U9543 (N_9543,N_8439,N_8627);
nor U9544 (N_9544,N_8020,N_8711);
xor U9545 (N_9545,N_8805,N_8229);
xnor U9546 (N_9546,N_8296,N_8247);
or U9547 (N_9547,N_8913,N_8567);
xnor U9548 (N_9548,N_8639,N_8380);
nand U9549 (N_9549,N_8164,N_8613);
nor U9550 (N_9550,N_8582,N_8944);
nor U9551 (N_9551,N_8589,N_8513);
nor U9552 (N_9552,N_8400,N_8656);
and U9553 (N_9553,N_8763,N_8053);
nor U9554 (N_9554,N_8361,N_8793);
and U9555 (N_9555,N_8818,N_8167);
and U9556 (N_9556,N_8836,N_8571);
nor U9557 (N_9557,N_8658,N_8151);
or U9558 (N_9558,N_8900,N_8089);
nand U9559 (N_9559,N_8414,N_8868);
xnor U9560 (N_9560,N_8315,N_8400);
or U9561 (N_9561,N_8634,N_8426);
nor U9562 (N_9562,N_8958,N_8816);
nand U9563 (N_9563,N_8789,N_8273);
nor U9564 (N_9564,N_8210,N_8230);
xnor U9565 (N_9565,N_8924,N_8808);
nand U9566 (N_9566,N_8995,N_8724);
and U9567 (N_9567,N_8918,N_8581);
nand U9568 (N_9568,N_8593,N_8136);
nand U9569 (N_9569,N_8053,N_8500);
nand U9570 (N_9570,N_8897,N_8882);
or U9571 (N_9571,N_8535,N_8663);
nor U9572 (N_9572,N_8850,N_8246);
nand U9573 (N_9573,N_8514,N_8994);
xor U9574 (N_9574,N_8678,N_8291);
nor U9575 (N_9575,N_8609,N_8026);
xor U9576 (N_9576,N_8719,N_8697);
or U9577 (N_9577,N_8653,N_8517);
nand U9578 (N_9578,N_8680,N_8126);
and U9579 (N_9579,N_8684,N_8051);
nor U9580 (N_9580,N_8686,N_8795);
and U9581 (N_9581,N_8616,N_8415);
or U9582 (N_9582,N_8497,N_8437);
and U9583 (N_9583,N_8415,N_8681);
xor U9584 (N_9584,N_8853,N_8038);
nand U9585 (N_9585,N_8383,N_8206);
nor U9586 (N_9586,N_8355,N_8391);
nand U9587 (N_9587,N_8581,N_8480);
and U9588 (N_9588,N_8206,N_8398);
nor U9589 (N_9589,N_8041,N_8764);
nor U9590 (N_9590,N_8949,N_8445);
nor U9591 (N_9591,N_8820,N_8527);
xor U9592 (N_9592,N_8511,N_8245);
nand U9593 (N_9593,N_8057,N_8810);
and U9594 (N_9594,N_8898,N_8094);
nand U9595 (N_9595,N_8057,N_8107);
xor U9596 (N_9596,N_8145,N_8629);
xor U9597 (N_9597,N_8434,N_8911);
xor U9598 (N_9598,N_8969,N_8992);
or U9599 (N_9599,N_8917,N_8925);
nand U9600 (N_9600,N_8491,N_8788);
xor U9601 (N_9601,N_8822,N_8995);
or U9602 (N_9602,N_8733,N_8265);
xnor U9603 (N_9603,N_8141,N_8617);
nand U9604 (N_9604,N_8486,N_8115);
nand U9605 (N_9605,N_8589,N_8175);
xor U9606 (N_9606,N_8237,N_8249);
or U9607 (N_9607,N_8329,N_8990);
or U9608 (N_9608,N_8874,N_8448);
or U9609 (N_9609,N_8501,N_8406);
nand U9610 (N_9610,N_8323,N_8885);
nor U9611 (N_9611,N_8455,N_8627);
or U9612 (N_9612,N_8325,N_8346);
xnor U9613 (N_9613,N_8324,N_8672);
or U9614 (N_9614,N_8910,N_8642);
nor U9615 (N_9615,N_8564,N_8321);
and U9616 (N_9616,N_8353,N_8467);
and U9617 (N_9617,N_8818,N_8744);
nand U9618 (N_9618,N_8869,N_8728);
and U9619 (N_9619,N_8148,N_8354);
or U9620 (N_9620,N_8109,N_8762);
and U9621 (N_9621,N_8152,N_8844);
and U9622 (N_9622,N_8775,N_8985);
or U9623 (N_9623,N_8619,N_8437);
nand U9624 (N_9624,N_8903,N_8946);
or U9625 (N_9625,N_8081,N_8801);
or U9626 (N_9626,N_8292,N_8156);
nand U9627 (N_9627,N_8547,N_8025);
xor U9628 (N_9628,N_8195,N_8496);
nand U9629 (N_9629,N_8766,N_8898);
and U9630 (N_9630,N_8342,N_8173);
nor U9631 (N_9631,N_8170,N_8363);
nor U9632 (N_9632,N_8029,N_8084);
or U9633 (N_9633,N_8873,N_8540);
or U9634 (N_9634,N_8010,N_8591);
and U9635 (N_9635,N_8040,N_8665);
or U9636 (N_9636,N_8992,N_8451);
xor U9637 (N_9637,N_8397,N_8915);
nand U9638 (N_9638,N_8943,N_8846);
nand U9639 (N_9639,N_8895,N_8629);
nand U9640 (N_9640,N_8926,N_8140);
and U9641 (N_9641,N_8852,N_8514);
nand U9642 (N_9642,N_8642,N_8423);
nor U9643 (N_9643,N_8116,N_8701);
xnor U9644 (N_9644,N_8164,N_8100);
or U9645 (N_9645,N_8663,N_8889);
nor U9646 (N_9646,N_8306,N_8370);
and U9647 (N_9647,N_8984,N_8293);
nand U9648 (N_9648,N_8212,N_8679);
nand U9649 (N_9649,N_8395,N_8102);
and U9650 (N_9650,N_8041,N_8521);
or U9651 (N_9651,N_8060,N_8752);
nand U9652 (N_9652,N_8847,N_8145);
and U9653 (N_9653,N_8269,N_8106);
nor U9654 (N_9654,N_8982,N_8500);
and U9655 (N_9655,N_8175,N_8515);
nand U9656 (N_9656,N_8383,N_8672);
and U9657 (N_9657,N_8301,N_8591);
nor U9658 (N_9658,N_8875,N_8314);
and U9659 (N_9659,N_8938,N_8463);
and U9660 (N_9660,N_8754,N_8320);
and U9661 (N_9661,N_8735,N_8478);
nand U9662 (N_9662,N_8589,N_8614);
nor U9663 (N_9663,N_8485,N_8402);
nor U9664 (N_9664,N_8708,N_8881);
or U9665 (N_9665,N_8038,N_8863);
and U9666 (N_9666,N_8526,N_8326);
and U9667 (N_9667,N_8333,N_8885);
and U9668 (N_9668,N_8238,N_8681);
xnor U9669 (N_9669,N_8284,N_8988);
or U9670 (N_9670,N_8214,N_8124);
xor U9671 (N_9671,N_8943,N_8666);
nand U9672 (N_9672,N_8472,N_8237);
or U9673 (N_9673,N_8604,N_8261);
and U9674 (N_9674,N_8369,N_8851);
or U9675 (N_9675,N_8237,N_8091);
nor U9676 (N_9676,N_8987,N_8428);
xnor U9677 (N_9677,N_8513,N_8982);
nand U9678 (N_9678,N_8441,N_8698);
nor U9679 (N_9679,N_8294,N_8341);
xnor U9680 (N_9680,N_8044,N_8492);
nand U9681 (N_9681,N_8323,N_8480);
or U9682 (N_9682,N_8393,N_8793);
and U9683 (N_9683,N_8436,N_8162);
or U9684 (N_9684,N_8640,N_8675);
nand U9685 (N_9685,N_8572,N_8041);
xnor U9686 (N_9686,N_8997,N_8639);
and U9687 (N_9687,N_8288,N_8722);
nor U9688 (N_9688,N_8711,N_8740);
nand U9689 (N_9689,N_8564,N_8043);
xnor U9690 (N_9690,N_8350,N_8823);
nand U9691 (N_9691,N_8375,N_8156);
xnor U9692 (N_9692,N_8025,N_8053);
and U9693 (N_9693,N_8667,N_8302);
xor U9694 (N_9694,N_8998,N_8350);
xnor U9695 (N_9695,N_8806,N_8664);
or U9696 (N_9696,N_8896,N_8636);
xor U9697 (N_9697,N_8005,N_8501);
xnor U9698 (N_9698,N_8879,N_8940);
or U9699 (N_9699,N_8503,N_8656);
nor U9700 (N_9700,N_8746,N_8908);
and U9701 (N_9701,N_8120,N_8920);
nor U9702 (N_9702,N_8682,N_8135);
nand U9703 (N_9703,N_8605,N_8463);
nor U9704 (N_9704,N_8336,N_8034);
or U9705 (N_9705,N_8039,N_8558);
and U9706 (N_9706,N_8129,N_8428);
xor U9707 (N_9707,N_8397,N_8182);
xor U9708 (N_9708,N_8771,N_8300);
nand U9709 (N_9709,N_8916,N_8092);
and U9710 (N_9710,N_8439,N_8153);
nand U9711 (N_9711,N_8935,N_8427);
and U9712 (N_9712,N_8815,N_8040);
or U9713 (N_9713,N_8939,N_8683);
or U9714 (N_9714,N_8102,N_8464);
and U9715 (N_9715,N_8552,N_8397);
xor U9716 (N_9716,N_8221,N_8547);
or U9717 (N_9717,N_8904,N_8788);
or U9718 (N_9718,N_8749,N_8421);
and U9719 (N_9719,N_8274,N_8126);
nor U9720 (N_9720,N_8656,N_8948);
nor U9721 (N_9721,N_8886,N_8083);
and U9722 (N_9722,N_8510,N_8054);
or U9723 (N_9723,N_8953,N_8601);
and U9724 (N_9724,N_8442,N_8611);
nor U9725 (N_9725,N_8333,N_8474);
or U9726 (N_9726,N_8660,N_8500);
nand U9727 (N_9727,N_8890,N_8696);
and U9728 (N_9728,N_8528,N_8616);
and U9729 (N_9729,N_8124,N_8030);
xor U9730 (N_9730,N_8771,N_8202);
nand U9731 (N_9731,N_8780,N_8266);
xor U9732 (N_9732,N_8028,N_8336);
or U9733 (N_9733,N_8746,N_8096);
nand U9734 (N_9734,N_8158,N_8103);
xnor U9735 (N_9735,N_8624,N_8527);
nand U9736 (N_9736,N_8191,N_8915);
xnor U9737 (N_9737,N_8147,N_8750);
nor U9738 (N_9738,N_8087,N_8530);
nor U9739 (N_9739,N_8400,N_8442);
or U9740 (N_9740,N_8658,N_8941);
nor U9741 (N_9741,N_8181,N_8302);
or U9742 (N_9742,N_8467,N_8745);
xor U9743 (N_9743,N_8779,N_8216);
xnor U9744 (N_9744,N_8693,N_8220);
and U9745 (N_9745,N_8102,N_8294);
nor U9746 (N_9746,N_8090,N_8854);
nand U9747 (N_9747,N_8139,N_8544);
nand U9748 (N_9748,N_8744,N_8434);
xor U9749 (N_9749,N_8977,N_8098);
nand U9750 (N_9750,N_8462,N_8641);
nor U9751 (N_9751,N_8537,N_8773);
nor U9752 (N_9752,N_8351,N_8788);
or U9753 (N_9753,N_8622,N_8516);
or U9754 (N_9754,N_8994,N_8813);
or U9755 (N_9755,N_8699,N_8965);
nor U9756 (N_9756,N_8300,N_8556);
nand U9757 (N_9757,N_8483,N_8663);
and U9758 (N_9758,N_8003,N_8123);
or U9759 (N_9759,N_8642,N_8265);
nand U9760 (N_9760,N_8044,N_8242);
xnor U9761 (N_9761,N_8682,N_8449);
or U9762 (N_9762,N_8407,N_8557);
and U9763 (N_9763,N_8785,N_8454);
or U9764 (N_9764,N_8545,N_8963);
or U9765 (N_9765,N_8873,N_8247);
nand U9766 (N_9766,N_8813,N_8666);
nor U9767 (N_9767,N_8741,N_8258);
nor U9768 (N_9768,N_8178,N_8276);
xor U9769 (N_9769,N_8457,N_8635);
nand U9770 (N_9770,N_8348,N_8418);
nor U9771 (N_9771,N_8799,N_8981);
nand U9772 (N_9772,N_8544,N_8047);
nand U9773 (N_9773,N_8430,N_8359);
nand U9774 (N_9774,N_8562,N_8129);
and U9775 (N_9775,N_8018,N_8113);
and U9776 (N_9776,N_8188,N_8465);
nand U9777 (N_9777,N_8764,N_8723);
and U9778 (N_9778,N_8742,N_8227);
and U9779 (N_9779,N_8278,N_8153);
nand U9780 (N_9780,N_8303,N_8925);
and U9781 (N_9781,N_8425,N_8940);
nor U9782 (N_9782,N_8401,N_8206);
xor U9783 (N_9783,N_8152,N_8458);
or U9784 (N_9784,N_8621,N_8679);
or U9785 (N_9785,N_8890,N_8367);
xnor U9786 (N_9786,N_8863,N_8450);
nor U9787 (N_9787,N_8630,N_8114);
nor U9788 (N_9788,N_8102,N_8416);
and U9789 (N_9789,N_8575,N_8053);
nand U9790 (N_9790,N_8391,N_8965);
xor U9791 (N_9791,N_8409,N_8488);
xor U9792 (N_9792,N_8697,N_8547);
and U9793 (N_9793,N_8573,N_8173);
xnor U9794 (N_9794,N_8302,N_8837);
or U9795 (N_9795,N_8823,N_8017);
nand U9796 (N_9796,N_8063,N_8329);
nand U9797 (N_9797,N_8265,N_8387);
or U9798 (N_9798,N_8977,N_8033);
and U9799 (N_9799,N_8342,N_8642);
nor U9800 (N_9800,N_8745,N_8101);
nand U9801 (N_9801,N_8708,N_8153);
or U9802 (N_9802,N_8326,N_8346);
nand U9803 (N_9803,N_8750,N_8572);
nor U9804 (N_9804,N_8288,N_8804);
or U9805 (N_9805,N_8509,N_8491);
xnor U9806 (N_9806,N_8731,N_8520);
and U9807 (N_9807,N_8994,N_8332);
nor U9808 (N_9808,N_8093,N_8207);
nor U9809 (N_9809,N_8393,N_8240);
and U9810 (N_9810,N_8060,N_8184);
nor U9811 (N_9811,N_8291,N_8051);
xor U9812 (N_9812,N_8923,N_8582);
and U9813 (N_9813,N_8901,N_8704);
and U9814 (N_9814,N_8154,N_8684);
nand U9815 (N_9815,N_8913,N_8615);
nor U9816 (N_9816,N_8601,N_8206);
nor U9817 (N_9817,N_8558,N_8575);
and U9818 (N_9818,N_8775,N_8077);
nor U9819 (N_9819,N_8881,N_8634);
xnor U9820 (N_9820,N_8909,N_8634);
xnor U9821 (N_9821,N_8277,N_8816);
or U9822 (N_9822,N_8311,N_8467);
xnor U9823 (N_9823,N_8772,N_8831);
nand U9824 (N_9824,N_8674,N_8156);
nand U9825 (N_9825,N_8822,N_8670);
and U9826 (N_9826,N_8669,N_8405);
nor U9827 (N_9827,N_8551,N_8642);
xor U9828 (N_9828,N_8191,N_8709);
nor U9829 (N_9829,N_8863,N_8300);
nor U9830 (N_9830,N_8382,N_8276);
nor U9831 (N_9831,N_8235,N_8232);
nand U9832 (N_9832,N_8328,N_8055);
nand U9833 (N_9833,N_8499,N_8759);
nand U9834 (N_9834,N_8365,N_8420);
nand U9835 (N_9835,N_8365,N_8123);
or U9836 (N_9836,N_8069,N_8904);
and U9837 (N_9837,N_8863,N_8675);
nand U9838 (N_9838,N_8009,N_8187);
xnor U9839 (N_9839,N_8624,N_8590);
or U9840 (N_9840,N_8912,N_8095);
xnor U9841 (N_9841,N_8765,N_8408);
nor U9842 (N_9842,N_8388,N_8020);
nor U9843 (N_9843,N_8725,N_8760);
nand U9844 (N_9844,N_8508,N_8934);
nand U9845 (N_9845,N_8468,N_8234);
nor U9846 (N_9846,N_8884,N_8999);
nor U9847 (N_9847,N_8478,N_8516);
xnor U9848 (N_9848,N_8778,N_8870);
nand U9849 (N_9849,N_8009,N_8682);
xnor U9850 (N_9850,N_8485,N_8427);
nand U9851 (N_9851,N_8877,N_8844);
xor U9852 (N_9852,N_8689,N_8128);
and U9853 (N_9853,N_8880,N_8426);
xor U9854 (N_9854,N_8446,N_8667);
xor U9855 (N_9855,N_8221,N_8482);
nor U9856 (N_9856,N_8660,N_8413);
nor U9857 (N_9857,N_8178,N_8760);
xnor U9858 (N_9858,N_8676,N_8930);
or U9859 (N_9859,N_8938,N_8453);
nand U9860 (N_9860,N_8032,N_8228);
or U9861 (N_9861,N_8619,N_8943);
and U9862 (N_9862,N_8508,N_8854);
nor U9863 (N_9863,N_8211,N_8890);
xor U9864 (N_9864,N_8034,N_8296);
and U9865 (N_9865,N_8883,N_8493);
or U9866 (N_9866,N_8540,N_8435);
or U9867 (N_9867,N_8788,N_8380);
nor U9868 (N_9868,N_8180,N_8124);
or U9869 (N_9869,N_8573,N_8670);
and U9870 (N_9870,N_8419,N_8206);
and U9871 (N_9871,N_8262,N_8261);
nor U9872 (N_9872,N_8139,N_8782);
xnor U9873 (N_9873,N_8136,N_8833);
and U9874 (N_9874,N_8879,N_8932);
and U9875 (N_9875,N_8588,N_8114);
nand U9876 (N_9876,N_8559,N_8069);
nor U9877 (N_9877,N_8815,N_8924);
nor U9878 (N_9878,N_8472,N_8260);
xor U9879 (N_9879,N_8549,N_8240);
xor U9880 (N_9880,N_8848,N_8940);
or U9881 (N_9881,N_8847,N_8089);
and U9882 (N_9882,N_8539,N_8580);
xor U9883 (N_9883,N_8896,N_8046);
nand U9884 (N_9884,N_8607,N_8347);
or U9885 (N_9885,N_8500,N_8371);
and U9886 (N_9886,N_8357,N_8435);
and U9887 (N_9887,N_8362,N_8232);
and U9888 (N_9888,N_8707,N_8946);
nor U9889 (N_9889,N_8297,N_8887);
nor U9890 (N_9890,N_8917,N_8517);
nand U9891 (N_9891,N_8481,N_8278);
nand U9892 (N_9892,N_8672,N_8686);
or U9893 (N_9893,N_8692,N_8296);
and U9894 (N_9894,N_8051,N_8148);
nor U9895 (N_9895,N_8151,N_8642);
xor U9896 (N_9896,N_8246,N_8982);
xor U9897 (N_9897,N_8979,N_8034);
nor U9898 (N_9898,N_8020,N_8119);
xnor U9899 (N_9899,N_8601,N_8530);
and U9900 (N_9900,N_8518,N_8022);
and U9901 (N_9901,N_8532,N_8407);
or U9902 (N_9902,N_8526,N_8952);
and U9903 (N_9903,N_8282,N_8298);
xnor U9904 (N_9904,N_8465,N_8934);
and U9905 (N_9905,N_8496,N_8163);
or U9906 (N_9906,N_8392,N_8477);
nor U9907 (N_9907,N_8835,N_8728);
or U9908 (N_9908,N_8172,N_8825);
xnor U9909 (N_9909,N_8899,N_8034);
nor U9910 (N_9910,N_8451,N_8442);
xor U9911 (N_9911,N_8897,N_8900);
or U9912 (N_9912,N_8273,N_8930);
or U9913 (N_9913,N_8455,N_8142);
xor U9914 (N_9914,N_8447,N_8223);
or U9915 (N_9915,N_8794,N_8992);
nor U9916 (N_9916,N_8483,N_8670);
nor U9917 (N_9917,N_8734,N_8796);
xnor U9918 (N_9918,N_8843,N_8482);
nand U9919 (N_9919,N_8244,N_8339);
xor U9920 (N_9920,N_8584,N_8192);
xor U9921 (N_9921,N_8807,N_8102);
nor U9922 (N_9922,N_8813,N_8147);
xor U9923 (N_9923,N_8825,N_8937);
xnor U9924 (N_9924,N_8164,N_8241);
or U9925 (N_9925,N_8156,N_8451);
and U9926 (N_9926,N_8720,N_8986);
nor U9927 (N_9927,N_8399,N_8568);
xor U9928 (N_9928,N_8298,N_8612);
or U9929 (N_9929,N_8296,N_8584);
xor U9930 (N_9930,N_8744,N_8842);
xor U9931 (N_9931,N_8280,N_8299);
nand U9932 (N_9932,N_8279,N_8184);
and U9933 (N_9933,N_8923,N_8886);
or U9934 (N_9934,N_8160,N_8880);
or U9935 (N_9935,N_8385,N_8818);
or U9936 (N_9936,N_8019,N_8500);
xor U9937 (N_9937,N_8982,N_8940);
or U9938 (N_9938,N_8489,N_8017);
nand U9939 (N_9939,N_8722,N_8509);
and U9940 (N_9940,N_8182,N_8654);
or U9941 (N_9941,N_8624,N_8925);
or U9942 (N_9942,N_8527,N_8170);
or U9943 (N_9943,N_8823,N_8774);
or U9944 (N_9944,N_8748,N_8437);
nand U9945 (N_9945,N_8440,N_8498);
or U9946 (N_9946,N_8141,N_8648);
nand U9947 (N_9947,N_8778,N_8959);
or U9948 (N_9948,N_8930,N_8506);
and U9949 (N_9949,N_8512,N_8136);
xnor U9950 (N_9950,N_8734,N_8294);
nor U9951 (N_9951,N_8930,N_8197);
nor U9952 (N_9952,N_8201,N_8347);
nor U9953 (N_9953,N_8634,N_8082);
nand U9954 (N_9954,N_8098,N_8524);
nor U9955 (N_9955,N_8363,N_8881);
xnor U9956 (N_9956,N_8663,N_8677);
nand U9957 (N_9957,N_8019,N_8855);
xor U9958 (N_9958,N_8600,N_8778);
or U9959 (N_9959,N_8077,N_8104);
xnor U9960 (N_9960,N_8230,N_8245);
nor U9961 (N_9961,N_8770,N_8510);
nor U9962 (N_9962,N_8812,N_8714);
or U9963 (N_9963,N_8609,N_8177);
xor U9964 (N_9964,N_8117,N_8808);
and U9965 (N_9965,N_8958,N_8160);
and U9966 (N_9966,N_8651,N_8923);
or U9967 (N_9967,N_8310,N_8785);
nor U9968 (N_9968,N_8470,N_8929);
nor U9969 (N_9969,N_8544,N_8550);
xor U9970 (N_9970,N_8328,N_8910);
nand U9971 (N_9971,N_8453,N_8757);
nor U9972 (N_9972,N_8478,N_8178);
or U9973 (N_9973,N_8349,N_8785);
or U9974 (N_9974,N_8535,N_8473);
and U9975 (N_9975,N_8186,N_8035);
xnor U9976 (N_9976,N_8469,N_8937);
nand U9977 (N_9977,N_8695,N_8394);
nor U9978 (N_9978,N_8207,N_8392);
nor U9979 (N_9979,N_8558,N_8842);
nand U9980 (N_9980,N_8642,N_8699);
nor U9981 (N_9981,N_8244,N_8417);
or U9982 (N_9982,N_8663,N_8284);
nor U9983 (N_9983,N_8659,N_8892);
nand U9984 (N_9984,N_8027,N_8900);
and U9985 (N_9985,N_8848,N_8015);
xor U9986 (N_9986,N_8171,N_8369);
nor U9987 (N_9987,N_8904,N_8962);
and U9988 (N_9988,N_8724,N_8167);
nor U9989 (N_9989,N_8610,N_8751);
xor U9990 (N_9990,N_8463,N_8817);
xnor U9991 (N_9991,N_8968,N_8252);
or U9992 (N_9992,N_8896,N_8948);
nor U9993 (N_9993,N_8101,N_8724);
or U9994 (N_9994,N_8288,N_8335);
nand U9995 (N_9995,N_8182,N_8914);
and U9996 (N_9996,N_8582,N_8439);
nand U9997 (N_9997,N_8195,N_8561);
nor U9998 (N_9998,N_8476,N_8975);
or U9999 (N_9999,N_8080,N_8944);
xnor U10000 (N_10000,N_9242,N_9733);
xnor U10001 (N_10001,N_9251,N_9862);
and U10002 (N_10002,N_9457,N_9535);
and U10003 (N_10003,N_9334,N_9686);
xnor U10004 (N_10004,N_9365,N_9531);
or U10005 (N_10005,N_9904,N_9623);
nand U10006 (N_10006,N_9223,N_9064);
or U10007 (N_10007,N_9630,N_9224);
nand U10008 (N_10008,N_9451,N_9384);
nand U10009 (N_10009,N_9734,N_9758);
xnor U10010 (N_10010,N_9133,N_9414);
xor U10011 (N_10011,N_9494,N_9413);
or U10012 (N_10012,N_9958,N_9530);
nor U10013 (N_10013,N_9683,N_9346);
or U10014 (N_10014,N_9967,N_9998);
nor U10015 (N_10015,N_9625,N_9893);
and U10016 (N_10016,N_9736,N_9565);
or U10017 (N_10017,N_9276,N_9634);
nand U10018 (N_10018,N_9216,N_9737);
and U10019 (N_10019,N_9128,N_9485);
or U10020 (N_10020,N_9373,N_9676);
nand U10021 (N_10021,N_9984,N_9685);
or U10022 (N_10022,N_9790,N_9280);
or U10023 (N_10023,N_9661,N_9616);
xor U10024 (N_10024,N_9048,N_9279);
xnor U10025 (N_10025,N_9475,N_9724);
nor U10026 (N_10026,N_9288,N_9919);
and U10027 (N_10027,N_9305,N_9896);
and U10028 (N_10028,N_9627,N_9636);
xor U10029 (N_10029,N_9842,N_9932);
nand U10030 (N_10030,N_9101,N_9235);
or U10031 (N_10031,N_9441,N_9860);
xor U10032 (N_10032,N_9826,N_9997);
nor U10033 (N_10033,N_9337,N_9274);
nor U10034 (N_10034,N_9867,N_9138);
and U10035 (N_10035,N_9857,N_9117);
and U10036 (N_10036,N_9240,N_9488);
xor U10037 (N_10037,N_9411,N_9112);
xnor U10038 (N_10038,N_9241,N_9234);
and U10039 (N_10039,N_9991,N_9065);
xnor U10040 (N_10040,N_9143,N_9566);
and U10041 (N_10041,N_9186,N_9777);
nand U10042 (N_10042,N_9600,N_9921);
nor U10043 (N_10043,N_9882,N_9512);
nand U10044 (N_10044,N_9957,N_9474);
or U10045 (N_10045,N_9554,N_9730);
or U10046 (N_10046,N_9601,N_9892);
nand U10047 (N_10047,N_9521,N_9985);
or U10048 (N_10048,N_9670,N_9340);
xnor U10049 (N_10049,N_9057,N_9495);
nand U10050 (N_10050,N_9338,N_9275);
nand U10051 (N_10051,N_9778,N_9193);
or U10052 (N_10052,N_9834,N_9018);
and U10053 (N_10053,N_9110,N_9067);
or U10054 (N_10054,N_9339,N_9523);
nor U10055 (N_10055,N_9607,N_9529);
nor U10056 (N_10056,N_9420,N_9693);
xnor U10057 (N_10057,N_9575,N_9092);
and U10058 (N_10058,N_9253,N_9383);
or U10059 (N_10059,N_9157,N_9121);
xnor U10060 (N_10060,N_9788,N_9135);
or U10061 (N_10061,N_9605,N_9491);
nand U10062 (N_10062,N_9828,N_9708);
xor U10063 (N_10063,N_9401,N_9300);
and U10064 (N_10064,N_9403,N_9171);
nor U10065 (N_10065,N_9940,N_9327);
xor U10066 (N_10066,N_9850,N_9208);
and U10067 (N_10067,N_9141,N_9079);
and U10068 (N_10068,N_9701,N_9229);
or U10069 (N_10069,N_9260,N_9863);
xnor U10070 (N_10070,N_9342,N_9682);
and U10071 (N_10071,N_9810,N_9318);
and U10072 (N_10072,N_9209,N_9387);
xor U10073 (N_10073,N_9233,N_9037);
nand U10074 (N_10074,N_9363,N_9717);
nand U10075 (N_10075,N_9032,N_9221);
nor U10076 (N_10076,N_9493,N_9360);
nand U10077 (N_10077,N_9785,N_9895);
nand U10078 (N_10078,N_9651,N_9968);
nand U10079 (N_10079,N_9210,N_9688);
and U10080 (N_10080,N_9602,N_9847);
nand U10081 (N_10081,N_9422,N_9098);
or U10082 (N_10082,N_9243,N_9111);
and U10083 (N_10083,N_9646,N_9760);
xnor U10084 (N_10084,N_9027,N_9900);
or U10085 (N_10085,N_9052,N_9712);
or U10086 (N_10086,N_9839,N_9269);
or U10087 (N_10087,N_9690,N_9631);
or U10088 (N_10088,N_9739,N_9572);
xnor U10089 (N_10089,N_9144,N_9899);
xnor U10090 (N_10090,N_9538,N_9920);
and U10091 (N_10091,N_9444,N_9879);
xor U10092 (N_10092,N_9817,N_9819);
nor U10093 (N_10093,N_9119,N_9865);
or U10094 (N_10094,N_9513,N_9382);
xor U10095 (N_10095,N_9341,N_9410);
and U10096 (N_10096,N_9011,N_9519);
nand U10097 (N_10097,N_9800,N_9754);
or U10098 (N_10098,N_9801,N_9814);
or U10099 (N_10099,N_9731,N_9884);
or U10100 (N_10100,N_9324,N_9977);
nor U10101 (N_10101,N_9930,N_9296);
nor U10102 (N_10102,N_9870,N_9502);
and U10103 (N_10103,N_9447,N_9332);
nor U10104 (N_10104,N_9039,N_9239);
and U10105 (N_10105,N_9563,N_9325);
xnor U10106 (N_10106,N_9644,N_9041);
xnor U10107 (N_10107,N_9218,N_9626);
nand U10108 (N_10108,N_9752,N_9798);
xor U10109 (N_10109,N_9150,N_9725);
or U10110 (N_10110,N_9055,N_9190);
nor U10111 (N_10111,N_9431,N_9771);
xor U10112 (N_10112,N_9905,N_9207);
and U10113 (N_10113,N_9671,N_9167);
or U10114 (N_10114,N_9987,N_9608);
and U10115 (N_10115,N_9880,N_9890);
nor U10116 (N_10116,N_9955,N_9791);
and U10117 (N_10117,N_9237,N_9746);
and U10118 (N_10118,N_9090,N_9377);
xnor U10119 (N_10119,N_9938,N_9259);
xor U10120 (N_10120,N_9293,N_9165);
and U10121 (N_10121,N_9120,N_9399);
and U10122 (N_10122,N_9578,N_9936);
xnor U10123 (N_10123,N_9854,N_9748);
and U10124 (N_10124,N_9284,N_9467);
xnor U10125 (N_10125,N_9799,N_9767);
xnor U10126 (N_10126,N_9917,N_9522);
nand U10127 (N_10127,N_9182,N_9869);
or U10128 (N_10128,N_9642,N_9619);
or U10129 (N_10129,N_9553,N_9329);
and U10130 (N_10130,N_9285,N_9290);
and U10131 (N_10131,N_9499,N_9425);
nor U10132 (N_10132,N_9875,N_9544);
or U10133 (N_10133,N_9184,N_9195);
xor U10134 (N_10134,N_9206,N_9592);
xor U10135 (N_10135,N_9942,N_9331);
xnor U10136 (N_10136,N_9889,N_9170);
xnor U10137 (N_10137,N_9198,N_9976);
or U10138 (N_10138,N_9076,N_9481);
or U10139 (N_10139,N_9181,N_9489);
nor U10140 (N_10140,N_9396,N_9019);
xor U10141 (N_10141,N_9476,N_9374);
and U10142 (N_10142,N_9624,N_9035);
nand U10143 (N_10143,N_9518,N_9770);
or U10144 (N_10144,N_9965,N_9336);
nand U10145 (N_10145,N_9372,N_9705);
nor U10146 (N_10146,N_9236,N_9564);
nand U10147 (N_10147,N_9164,N_9154);
and U10148 (N_10148,N_9094,N_9871);
nand U10149 (N_10149,N_9716,N_9428);
or U10150 (N_10150,N_9833,N_9830);
and U10151 (N_10151,N_9415,N_9852);
xnor U10152 (N_10152,N_9013,N_9802);
xor U10153 (N_10153,N_9872,N_9546);
or U10154 (N_10154,N_9005,N_9527);
nand U10155 (N_10155,N_9149,N_9461);
and U10156 (N_10156,N_9125,N_9924);
or U10157 (N_10157,N_9768,N_9114);
and U10158 (N_10158,N_9855,N_9258);
nor U10159 (N_10159,N_9326,N_9104);
or U10160 (N_10160,N_9614,N_9911);
xor U10161 (N_10161,N_9292,N_9268);
nand U10162 (N_10162,N_9452,N_9007);
or U10163 (N_10163,N_9647,N_9812);
and U10164 (N_10164,N_9020,N_9949);
nand U10165 (N_10165,N_9265,N_9202);
xnor U10166 (N_10166,N_9438,N_9903);
or U10167 (N_10167,N_9764,N_9901);
nor U10168 (N_10168,N_9172,N_9694);
nor U10169 (N_10169,N_9081,N_9567);
xnor U10170 (N_10170,N_9492,N_9674);
nand U10171 (N_10171,N_9783,N_9836);
and U10172 (N_10172,N_9349,N_9838);
and U10173 (N_10173,N_9909,N_9099);
xor U10174 (N_10174,N_9972,N_9267);
or U10175 (N_10175,N_9416,N_9139);
or U10176 (N_10176,N_9883,N_9316);
nor U10177 (N_10177,N_9406,N_9700);
nor U10178 (N_10178,N_9925,N_9794);
xor U10179 (N_10179,N_9351,N_9471);
xnor U10180 (N_10180,N_9272,N_9542);
xor U10181 (N_10181,N_9740,N_9846);
nand U10182 (N_10182,N_9283,N_9562);
xor U10183 (N_10183,N_9540,N_9528);
nand U10184 (N_10184,N_9097,N_9118);
or U10185 (N_10185,N_9075,N_9044);
or U10186 (N_10186,N_9295,N_9189);
or U10187 (N_10187,N_9058,N_9595);
nor U10188 (N_10188,N_9205,N_9633);
and U10189 (N_10189,N_9262,N_9086);
xor U10190 (N_10190,N_9049,N_9918);
nor U10191 (N_10191,N_9548,N_9162);
nand U10192 (N_10192,N_9449,N_9774);
and U10193 (N_10193,N_9996,N_9806);
xnor U10194 (N_10194,N_9792,N_9136);
and U10195 (N_10195,N_9158,N_9366);
or U10196 (N_10196,N_9371,N_9796);
or U10197 (N_10197,N_9402,N_9015);
and U10198 (N_10198,N_9151,N_9187);
nand U10199 (N_10199,N_9960,N_9808);
and U10200 (N_10200,N_9761,N_9131);
xor U10201 (N_10201,N_9759,N_9657);
nor U10202 (N_10202,N_9837,N_9307);
nor U10203 (N_10203,N_9995,N_9696);
xnor U10204 (N_10204,N_9036,N_9482);
and U10205 (N_10205,N_9937,N_9950);
and U10206 (N_10206,N_9908,N_9100);
or U10207 (N_10207,N_9795,N_9277);
xnor U10208 (N_10208,N_9720,N_9439);
nand U10209 (N_10209,N_9386,N_9063);
nand U10210 (N_10210,N_9639,N_9361);
xnor U10211 (N_10211,N_9388,N_9231);
and U10212 (N_10212,N_9106,N_9071);
nor U10213 (N_10213,N_9418,N_9787);
xnor U10214 (N_10214,N_9508,N_9465);
xnor U10215 (N_10215,N_9188,N_9962);
or U10216 (N_10216,N_9050,N_9568);
and U10217 (N_10217,N_9446,N_9105);
nand U10218 (N_10218,N_9317,N_9809);
nand U10219 (N_10219,N_9174,N_9008);
nor U10220 (N_10220,N_9191,N_9082);
nand U10221 (N_10221,N_9735,N_9551);
nand U10222 (N_10222,N_9654,N_9673);
or U10223 (N_10223,N_9749,N_9881);
nor U10224 (N_10224,N_9609,N_9823);
nand U10225 (N_10225,N_9581,N_9359);
nor U10226 (N_10226,N_9948,N_9663);
xor U10227 (N_10227,N_9935,N_9813);
xor U10228 (N_10228,N_9095,N_9002);
and U10229 (N_10229,N_9313,N_9517);
xnor U10230 (N_10230,N_9156,N_9507);
xor U10231 (N_10231,N_9408,N_9257);
nor U10232 (N_10232,N_9335,N_9009);
nand U10233 (N_10233,N_9311,N_9358);
xnor U10234 (N_10234,N_9448,N_9951);
and U10235 (N_10235,N_9741,N_9460);
nor U10236 (N_10236,N_9784,N_9291);
or U10237 (N_10237,N_9811,N_9772);
and U10238 (N_10238,N_9389,N_9982);
or U10239 (N_10239,N_9776,N_9322);
or U10240 (N_10240,N_9750,N_9804);
and U10241 (N_10241,N_9532,N_9487);
xor U10242 (N_10242,N_9593,N_9238);
nand U10243 (N_10243,N_9668,N_9727);
nor U10244 (N_10244,N_9963,N_9073);
xnor U10245 (N_10245,N_9454,N_9844);
xor U10246 (N_10246,N_9468,N_9559);
and U10247 (N_10247,N_9312,N_9675);
nor U10248 (N_10248,N_9001,N_9089);
xor U10249 (N_10249,N_9480,N_9711);
xnor U10250 (N_10250,N_9115,N_9022);
and U10251 (N_10251,N_9308,N_9667);
and U10252 (N_10252,N_9321,N_9123);
xor U10253 (N_10253,N_9023,N_9684);
nand U10254 (N_10254,N_9436,N_9355);
and U10255 (N_10255,N_9282,N_9858);
and U10256 (N_10256,N_9320,N_9072);
xnor U10257 (N_10257,N_9249,N_9861);
xnor U10258 (N_10258,N_9132,N_9672);
or U10259 (N_10259,N_9988,N_9160);
or U10260 (N_10260,N_9818,N_9247);
nand U10261 (N_10261,N_9124,N_9878);
nor U10262 (N_10262,N_9228,N_9766);
or U10263 (N_10263,N_9051,N_9443);
nor U10264 (N_10264,N_9978,N_9297);
xor U10265 (N_10265,N_9315,N_9886);
nor U10266 (N_10266,N_9992,N_9763);
nand U10267 (N_10267,N_9524,N_9547);
or U10268 (N_10268,N_9113,N_9570);
and U10269 (N_10269,N_9618,N_9560);
or U10270 (N_10270,N_9367,N_9163);
and U10271 (N_10271,N_9056,N_9244);
or U10272 (N_10272,N_9829,N_9613);
and U10273 (N_10273,N_9213,N_9702);
or U10274 (N_10274,N_9440,N_9078);
xor U10275 (N_10275,N_9681,N_9573);
xor U10276 (N_10276,N_9638,N_9526);
or U10277 (N_10277,N_9289,N_9969);
nand U10278 (N_10278,N_9204,N_9219);
xor U10279 (N_10279,N_9470,N_9662);
or U10280 (N_10280,N_9273,N_9264);
and U10281 (N_10281,N_9999,N_9314);
xor U10282 (N_10282,N_9498,N_9215);
nor U10283 (N_10283,N_9472,N_9509);
and U10284 (N_10284,N_9640,N_9505);
and U10285 (N_10285,N_9456,N_9914);
nor U10286 (N_10286,N_9753,N_9589);
or U10287 (N_10287,N_9864,N_9956);
or U10288 (N_10288,N_9169,N_9127);
nand U10289 (N_10289,N_9665,N_9179);
and U10290 (N_10290,N_9703,N_9405);
nor U10291 (N_10291,N_9569,N_9729);
nor U10292 (N_10292,N_9140,N_9028);
nor U10293 (N_10293,N_9217,N_9689);
nor U10294 (N_10294,N_9506,N_9354);
xor U10295 (N_10295,N_9641,N_9458);
xnor U10296 (N_10296,N_9435,N_9888);
and U10297 (N_10297,N_9477,N_9496);
and U10298 (N_10298,N_9822,N_9427);
or U10299 (N_10299,N_9426,N_9745);
nand U10300 (N_10300,N_9738,N_9550);
and U10301 (N_10301,N_9926,N_9782);
nor U10302 (N_10302,N_9145,N_9306);
nand U10303 (N_10303,N_9453,N_9755);
nand U10304 (N_10304,N_9713,N_9343);
nand U10305 (N_10305,N_9201,N_9805);
or U10306 (N_10306,N_9769,N_9934);
or U10307 (N_10307,N_9923,N_9907);
and U10308 (N_10308,N_9347,N_9841);
or U10309 (N_10309,N_9891,N_9271);
nor U10310 (N_10310,N_9010,N_9214);
xor U10311 (N_10311,N_9356,N_9579);
nand U10312 (N_10312,N_9226,N_9678);
or U10313 (N_10313,N_9364,N_9574);
xor U10314 (N_10314,N_9859,N_9130);
or U10315 (N_10315,N_9757,N_9062);
nor U10316 (N_10316,N_9946,N_9142);
xor U10317 (N_10317,N_9679,N_9319);
nand U10318 (N_10318,N_9256,N_9699);
nor U10319 (N_10319,N_9147,N_9152);
nor U10320 (N_10320,N_9068,N_9424);
and U10321 (N_10321,N_9877,N_9323);
xor U10322 (N_10322,N_9483,N_9973);
xnor U10323 (N_10323,N_9604,N_9541);
xor U10324 (N_10324,N_9612,N_9876);
xor U10325 (N_10325,N_9016,N_9287);
or U10326 (N_10326,N_9557,N_9378);
nand U10327 (N_10327,N_9434,N_9825);
nor U10328 (N_10328,N_9677,N_9598);
nor U10329 (N_10329,N_9853,N_9412);
xor U10330 (N_10330,N_9397,N_9929);
nor U10331 (N_10331,N_9000,N_9450);
xor U10332 (N_10332,N_9014,N_9721);
or U10333 (N_10333,N_9659,N_9137);
nor U10334 (N_10334,N_9747,N_9539);
xor U10335 (N_10335,N_9248,N_9691);
nor U10336 (N_10336,N_9765,N_9585);
nand U10337 (N_10337,N_9006,N_9611);
and U10338 (N_10338,N_9466,N_9635);
nor U10339 (N_10339,N_9084,N_9344);
nor U10340 (N_10340,N_9379,N_9501);
and U10341 (N_10341,N_9252,N_9898);
nand U10342 (N_10342,N_9155,N_9835);
nor U10343 (N_10343,N_9781,N_9046);
nor U10344 (N_10344,N_9353,N_9666);
nor U10345 (N_10345,N_9629,N_9718);
or U10346 (N_10346,N_9632,N_9643);
xor U10347 (N_10347,N_9180,N_9298);
xnor U10348 (N_10348,N_9779,N_9504);
xnor U10349 (N_10349,N_9655,N_9840);
nor U10350 (N_10350,N_9419,N_9178);
and U10351 (N_10351,N_9109,N_9885);
and U10352 (N_10352,N_9161,N_9515);
nor U10353 (N_10353,N_9744,N_9328);
nor U10354 (N_10354,N_9042,N_9971);
and U10355 (N_10355,N_9912,N_9497);
and U10356 (N_10356,N_9375,N_9980);
and U10357 (N_10357,N_9851,N_9060);
and U10358 (N_10358,N_9591,N_9916);
nand U10359 (N_10359,N_9059,N_9652);
and U10360 (N_10360,N_9815,N_9168);
or U10361 (N_10361,N_9080,N_9649);
or U10362 (N_10362,N_9025,N_9093);
nor U10363 (N_10363,N_9370,N_9430);
and U10364 (N_10364,N_9617,N_9230);
nand U10365 (N_10365,N_9902,N_9096);
nor U10366 (N_10366,N_9645,N_9603);
xnor U10367 (N_10367,N_9622,N_9742);
nand U10368 (N_10368,N_9516,N_9832);
nand U10369 (N_10369,N_9196,N_9376);
and U10370 (N_10370,N_9246,N_9628);
nor U10371 (N_10371,N_9599,N_9706);
nand U10372 (N_10372,N_9719,N_9185);
or U10373 (N_10373,N_9087,N_9959);
nand U10374 (N_10374,N_9463,N_9442);
nor U10375 (N_10375,N_9989,N_9054);
xnor U10376 (N_10376,N_9966,N_9176);
and U10377 (N_10377,N_9807,N_9263);
nand U10378 (N_10378,N_9116,N_9278);
and U10379 (N_10379,N_9122,N_9393);
xnor U10380 (N_10380,N_9017,N_9897);
xor U10381 (N_10381,N_9220,N_9571);
nand U10382 (N_10382,N_9085,N_9620);
or U10383 (N_10383,N_9203,N_9192);
or U10384 (N_10384,N_9561,N_9873);
nand U10385 (N_10385,N_9459,N_9333);
or U10386 (N_10386,N_9687,N_9421);
xor U10387 (N_10387,N_9843,N_9380);
and U10388 (N_10388,N_9789,N_9074);
nor U10389 (N_10389,N_9827,N_9514);
or U10390 (N_10390,N_9077,N_9266);
nor U10391 (N_10391,N_9793,N_9146);
or U10392 (N_10392,N_9362,N_9091);
nor U10393 (N_10393,N_9927,N_9543);
nor U10394 (N_10394,N_9310,N_9715);
nand U10395 (N_10395,N_9697,N_9510);
xnor U10396 (N_10396,N_9933,N_9003);
nand U10397 (N_10397,N_9660,N_9433);
nand U10398 (N_10398,N_9395,N_9558);
or U10399 (N_10399,N_9732,N_9029);
xor U10400 (N_10400,N_9820,N_9486);
nand U10401 (N_10401,N_9525,N_9584);
nor U10402 (N_10402,N_9587,N_9610);
xor U10403 (N_10403,N_9583,N_9511);
or U10404 (N_10404,N_9874,N_9281);
nand U10405 (N_10405,N_9648,N_9615);
or U10406 (N_10406,N_9033,N_9650);
xor U10407 (N_10407,N_9866,N_9500);
xnor U10408 (N_10408,N_9582,N_9030);
nor U10409 (N_10409,N_9126,N_9473);
nor U10410 (N_10410,N_9129,N_9102);
nand U10411 (N_10411,N_9294,N_9173);
nor U10412 (N_10412,N_9576,N_9714);
nand U10413 (N_10413,N_9780,N_9432);
nand U10414 (N_10414,N_9596,N_9350);
nor U10415 (N_10415,N_9270,N_9061);
xnor U10416 (N_10416,N_9031,N_9398);
nand U10417 (N_10417,N_9148,N_9200);
or U10418 (N_10418,N_9232,N_9577);
and U10419 (N_10419,N_9990,N_9445);
and U10420 (N_10420,N_9910,N_9845);
nor U10421 (N_10421,N_9175,N_9047);
xnor U10422 (N_10422,N_9710,N_9664);
nor U10423 (N_10423,N_9250,N_9939);
xnor U10424 (N_10424,N_9944,N_9301);
or U10425 (N_10425,N_9040,N_9979);
nand U10426 (N_10426,N_9153,N_9947);
nand U10427 (N_10427,N_9107,N_9352);
nor U10428 (N_10428,N_9545,N_9212);
xnor U10429 (N_10429,N_9183,N_9345);
xnor U10430 (N_10430,N_9953,N_9304);
nor U10431 (N_10431,N_9034,N_9704);
nor U10432 (N_10432,N_9868,N_9552);
nand U10433 (N_10433,N_9381,N_9597);
or U10434 (N_10434,N_9756,N_9417);
nor U10435 (N_10435,N_9952,N_9159);
nand U10436 (N_10436,N_9222,N_9773);
nand U10437 (N_10437,N_9534,N_9722);
and U10438 (N_10438,N_9199,N_9590);
or U10439 (N_10439,N_9066,N_9821);
nand U10440 (N_10440,N_9658,N_9357);
or U10441 (N_10441,N_9194,N_9254);
xnor U10442 (N_10442,N_9537,N_9261);
or U10443 (N_10443,N_9134,N_9588);
and U10444 (N_10444,N_9922,N_9786);
and U10445 (N_10445,N_9533,N_9586);
or U10446 (N_10446,N_9394,N_9580);
and U10447 (N_10447,N_9698,N_9803);
xor U10448 (N_10448,N_9227,N_9462);
and U10449 (N_10449,N_9594,N_9954);
xor U10450 (N_10450,N_9024,N_9177);
nand U10451 (N_10451,N_9848,N_9986);
or U10452 (N_10452,N_9108,N_9069);
and U10453 (N_10453,N_9887,N_9849);
and U10454 (N_10454,N_9728,N_9775);
nand U10455 (N_10455,N_9038,N_9469);
or U10456 (N_10456,N_9103,N_9669);
xnor U10457 (N_10457,N_9831,N_9083);
xnor U10458 (N_10458,N_9520,N_9026);
and U10459 (N_10459,N_9490,N_9709);
or U10460 (N_10460,N_9981,N_9330);
and U10461 (N_10461,N_9974,N_9556);
nand U10462 (N_10462,N_9245,N_9302);
nand U10463 (N_10463,N_9983,N_9484);
or U10464 (N_10464,N_9680,N_9348);
or U10465 (N_10465,N_9906,N_9856);
and U10466 (N_10466,N_9464,N_9400);
nand U10467 (N_10467,N_9166,N_9653);
and U10468 (N_10468,N_9606,N_9409);
nand U10469 (N_10469,N_9762,N_9088);
nand U10470 (N_10470,N_9743,N_9197);
xor U10471 (N_10471,N_9816,N_9915);
nor U10472 (N_10472,N_9455,N_9385);
or U10473 (N_10473,N_9478,N_9004);
and U10474 (N_10474,N_9993,N_9931);
and U10475 (N_10475,N_9392,N_9970);
and U10476 (N_10476,N_9053,N_9656);
nand U10477 (N_10477,N_9695,N_9961);
xor U10478 (N_10478,N_9043,N_9407);
or U10479 (N_10479,N_9943,N_9369);
or U10480 (N_10480,N_9975,N_9549);
xnor U10481 (N_10481,N_9368,N_9303);
xnor U10482 (N_10482,N_9429,N_9928);
or U10483 (N_10483,N_9536,N_9045);
nand U10484 (N_10484,N_9945,N_9012);
and U10485 (N_10485,N_9423,N_9894);
nand U10486 (N_10486,N_9437,N_9391);
nor U10487 (N_10487,N_9751,N_9723);
and U10488 (N_10488,N_9964,N_9555);
nor U10489 (N_10489,N_9479,N_9021);
xor U10490 (N_10490,N_9404,N_9692);
and U10491 (N_10491,N_9225,N_9726);
or U10492 (N_10492,N_9913,N_9390);
xnor U10493 (N_10493,N_9824,N_9211);
or U10494 (N_10494,N_9994,N_9299);
or U10495 (N_10495,N_9503,N_9941);
xnor U10496 (N_10496,N_9707,N_9797);
nor U10497 (N_10497,N_9621,N_9255);
nor U10498 (N_10498,N_9637,N_9286);
xnor U10499 (N_10499,N_9309,N_9070);
xor U10500 (N_10500,N_9003,N_9707);
or U10501 (N_10501,N_9939,N_9210);
nand U10502 (N_10502,N_9266,N_9770);
or U10503 (N_10503,N_9298,N_9481);
or U10504 (N_10504,N_9589,N_9592);
and U10505 (N_10505,N_9095,N_9653);
and U10506 (N_10506,N_9327,N_9096);
and U10507 (N_10507,N_9507,N_9647);
nor U10508 (N_10508,N_9082,N_9221);
or U10509 (N_10509,N_9201,N_9631);
nand U10510 (N_10510,N_9767,N_9160);
xor U10511 (N_10511,N_9140,N_9323);
xnor U10512 (N_10512,N_9829,N_9588);
or U10513 (N_10513,N_9064,N_9606);
xor U10514 (N_10514,N_9488,N_9929);
xor U10515 (N_10515,N_9649,N_9489);
nand U10516 (N_10516,N_9085,N_9851);
nand U10517 (N_10517,N_9315,N_9448);
nand U10518 (N_10518,N_9090,N_9133);
xnor U10519 (N_10519,N_9064,N_9460);
nor U10520 (N_10520,N_9082,N_9230);
nor U10521 (N_10521,N_9558,N_9722);
xnor U10522 (N_10522,N_9288,N_9328);
nand U10523 (N_10523,N_9234,N_9372);
or U10524 (N_10524,N_9390,N_9594);
xnor U10525 (N_10525,N_9924,N_9111);
and U10526 (N_10526,N_9246,N_9092);
or U10527 (N_10527,N_9918,N_9452);
and U10528 (N_10528,N_9271,N_9006);
and U10529 (N_10529,N_9452,N_9465);
nand U10530 (N_10530,N_9958,N_9770);
or U10531 (N_10531,N_9600,N_9073);
or U10532 (N_10532,N_9173,N_9392);
and U10533 (N_10533,N_9341,N_9108);
xnor U10534 (N_10534,N_9049,N_9759);
or U10535 (N_10535,N_9191,N_9760);
nor U10536 (N_10536,N_9157,N_9322);
nand U10537 (N_10537,N_9505,N_9859);
or U10538 (N_10538,N_9413,N_9486);
xor U10539 (N_10539,N_9233,N_9167);
nand U10540 (N_10540,N_9396,N_9134);
or U10541 (N_10541,N_9034,N_9155);
and U10542 (N_10542,N_9431,N_9456);
and U10543 (N_10543,N_9091,N_9017);
nand U10544 (N_10544,N_9035,N_9217);
and U10545 (N_10545,N_9780,N_9690);
xnor U10546 (N_10546,N_9381,N_9676);
nor U10547 (N_10547,N_9734,N_9802);
nand U10548 (N_10548,N_9700,N_9977);
and U10549 (N_10549,N_9138,N_9332);
and U10550 (N_10550,N_9273,N_9359);
nor U10551 (N_10551,N_9933,N_9352);
nand U10552 (N_10552,N_9282,N_9693);
or U10553 (N_10553,N_9013,N_9264);
and U10554 (N_10554,N_9354,N_9545);
xnor U10555 (N_10555,N_9281,N_9828);
nand U10556 (N_10556,N_9553,N_9851);
nand U10557 (N_10557,N_9831,N_9504);
and U10558 (N_10558,N_9544,N_9441);
nor U10559 (N_10559,N_9836,N_9755);
and U10560 (N_10560,N_9433,N_9461);
nor U10561 (N_10561,N_9616,N_9715);
nand U10562 (N_10562,N_9478,N_9923);
and U10563 (N_10563,N_9974,N_9295);
nor U10564 (N_10564,N_9848,N_9355);
nand U10565 (N_10565,N_9784,N_9853);
or U10566 (N_10566,N_9304,N_9177);
or U10567 (N_10567,N_9926,N_9074);
xor U10568 (N_10568,N_9769,N_9645);
xor U10569 (N_10569,N_9251,N_9752);
nor U10570 (N_10570,N_9356,N_9486);
or U10571 (N_10571,N_9666,N_9988);
xnor U10572 (N_10572,N_9001,N_9515);
xnor U10573 (N_10573,N_9219,N_9075);
xnor U10574 (N_10574,N_9869,N_9054);
nand U10575 (N_10575,N_9524,N_9487);
nand U10576 (N_10576,N_9637,N_9464);
or U10577 (N_10577,N_9073,N_9261);
nand U10578 (N_10578,N_9838,N_9355);
and U10579 (N_10579,N_9867,N_9605);
nor U10580 (N_10580,N_9012,N_9874);
xor U10581 (N_10581,N_9460,N_9335);
and U10582 (N_10582,N_9041,N_9460);
or U10583 (N_10583,N_9452,N_9336);
nand U10584 (N_10584,N_9517,N_9898);
xnor U10585 (N_10585,N_9794,N_9121);
or U10586 (N_10586,N_9455,N_9960);
xnor U10587 (N_10587,N_9701,N_9703);
nand U10588 (N_10588,N_9312,N_9510);
nand U10589 (N_10589,N_9695,N_9628);
nor U10590 (N_10590,N_9040,N_9650);
nor U10591 (N_10591,N_9201,N_9558);
xor U10592 (N_10592,N_9381,N_9906);
xnor U10593 (N_10593,N_9326,N_9400);
or U10594 (N_10594,N_9487,N_9423);
or U10595 (N_10595,N_9638,N_9056);
and U10596 (N_10596,N_9034,N_9221);
xor U10597 (N_10597,N_9384,N_9766);
or U10598 (N_10598,N_9713,N_9936);
nor U10599 (N_10599,N_9360,N_9118);
xnor U10600 (N_10600,N_9755,N_9216);
or U10601 (N_10601,N_9661,N_9368);
nor U10602 (N_10602,N_9295,N_9406);
nand U10603 (N_10603,N_9886,N_9180);
and U10604 (N_10604,N_9746,N_9944);
nor U10605 (N_10605,N_9374,N_9911);
xnor U10606 (N_10606,N_9066,N_9404);
and U10607 (N_10607,N_9998,N_9003);
nand U10608 (N_10608,N_9746,N_9658);
and U10609 (N_10609,N_9724,N_9629);
and U10610 (N_10610,N_9185,N_9755);
nor U10611 (N_10611,N_9775,N_9982);
nand U10612 (N_10612,N_9239,N_9472);
nor U10613 (N_10613,N_9710,N_9237);
nor U10614 (N_10614,N_9724,N_9217);
nor U10615 (N_10615,N_9787,N_9781);
and U10616 (N_10616,N_9289,N_9056);
and U10617 (N_10617,N_9461,N_9612);
and U10618 (N_10618,N_9771,N_9350);
xor U10619 (N_10619,N_9599,N_9509);
and U10620 (N_10620,N_9423,N_9810);
and U10621 (N_10621,N_9553,N_9124);
nor U10622 (N_10622,N_9573,N_9041);
nand U10623 (N_10623,N_9123,N_9956);
and U10624 (N_10624,N_9493,N_9114);
and U10625 (N_10625,N_9675,N_9631);
nand U10626 (N_10626,N_9060,N_9501);
nand U10627 (N_10627,N_9393,N_9284);
or U10628 (N_10628,N_9102,N_9318);
and U10629 (N_10629,N_9441,N_9057);
xnor U10630 (N_10630,N_9290,N_9965);
and U10631 (N_10631,N_9896,N_9150);
nor U10632 (N_10632,N_9986,N_9251);
nor U10633 (N_10633,N_9459,N_9310);
or U10634 (N_10634,N_9893,N_9174);
xnor U10635 (N_10635,N_9264,N_9215);
or U10636 (N_10636,N_9092,N_9142);
xor U10637 (N_10637,N_9094,N_9368);
or U10638 (N_10638,N_9354,N_9637);
or U10639 (N_10639,N_9119,N_9518);
or U10640 (N_10640,N_9397,N_9741);
nand U10641 (N_10641,N_9539,N_9560);
and U10642 (N_10642,N_9280,N_9609);
xnor U10643 (N_10643,N_9040,N_9897);
xor U10644 (N_10644,N_9418,N_9875);
nand U10645 (N_10645,N_9382,N_9637);
or U10646 (N_10646,N_9245,N_9636);
or U10647 (N_10647,N_9791,N_9683);
nand U10648 (N_10648,N_9120,N_9082);
xnor U10649 (N_10649,N_9291,N_9187);
or U10650 (N_10650,N_9979,N_9932);
nor U10651 (N_10651,N_9844,N_9897);
nand U10652 (N_10652,N_9208,N_9636);
nor U10653 (N_10653,N_9079,N_9336);
nand U10654 (N_10654,N_9626,N_9227);
and U10655 (N_10655,N_9554,N_9148);
nand U10656 (N_10656,N_9591,N_9403);
and U10657 (N_10657,N_9179,N_9650);
or U10658 (N_10658,N_9423,N_9986);
and U10659 (N_10659,N_9583,N_9256);
or U10660 (N_10660,N_9392,N_9966);
nor U10661 (N_10661,N_9943,N_9400);
nand U10662 (N_10662,N_9335,N_9570);
or U10663 (N_10663,N_9355,N_9981);
and U10664 (N_10664,N_9036,N_9401);
and U10665 (N_10665,N_9010,N_9402);
or U10666 (N_10666,N_9287,N_9052);
xor U10667 (N_10667,N_9282,N_9898);
xnor U10668 (N_10668,N_9514,N_9054);
or U10669 (N_10669,N_9426,N_9107);
nand U10670 (N_10670,N_9969,N_9243);
nand U10671 (N_10671,N_9200,N_9965);
nand U10672 (N_10672,N_9635,N_9644);
nand U10673 (N_10673,N_9804,N_9014);
and U10674 (N_10674,N_9763,N_9896);
xnor U10675 (N_10675,N_9489,N_9891);
and U10676 (N_10676,N_9374,N_9253);
or U10677 (N_10677,N_9120,N_9772);
xnor U10678 (N_10678,N_9420,N_9893);
and U10679 (N_10679,N_9010,N_9088);
nor U10680 (N_10680,N_9732,N_9728);
or U10681 (N_10681,N_9020,N_9688);
xor U10682 (N_10682,N_9323,N_9770);
and U10683 (N_10683,N_9252,N_9040);
and U10684 (N_10684,N_9486,N_9827);
nand U10685 (N_10685,N_9851,N_9727);
or U10686 (N_10686,N_9893,N_9607);
nand U10687 (N_10687,N_9815,N_9549);
or U10688 (N_10688,N_9043,N_9828);
xnor U10689 (N_10689,N_9594,N_9667);
or U10690 (N_10690,N_9486,N_9397);
xnor U10691 (N_10691,N_9366,N_9981);
nor U10692 (N_10692,N_9167,N_9426);
and U10693 (N_10693,N_9623,N_9621);
xnor U10694 (N_10694,N_9346,N_9147);
xor U10695 (N_10695,N_9956,N_9089);
and U10696 (N_10696,N_9282,N_9674);
and U10697 (N_10697,N_9582,N_9856);
or U10698 (N_10698,N_9258,N_9613);
and U10699 (N_10699,N_9606,N_9466);
nand U10700 (N_10700,N_9702,N_9110);
nor U10701 (N_10701,N_9755,N_9366);
and U10702 (N_10702,N_9957,N_9044);
xor U10703 (N_10703,N_9873,N_9201);
xnor U10704 (N_10704,N_9507,N_9802);
nor U10705 (N_10705,N_9589,N_9254);
and U10706 (N_10706,N_9362,N_9135);
xnor U10707 (N_10707,N_9183,N_9708);
nor U10708 (N_10708,N_9487,N_9757);
nor U10709 (N_10709,N_9370,N_9116);
xnor U10710 (N_10710,N_9734,N_9068);
or U10711 (N_10711,N_9570,N_9675);
and U10712 (N_10712,N_9781,N_9659);
nand U10713 (N_10713,N_9032,N_9683);
and U10714 (N_10714,N_9326,N_9418);
xnor U10715 (N_10715,N_9584,N_9223);
nand U10716 (N_10716,N_9039,N_9005);
nand U10717 (N_10717,N_9372,N_9325);
nand U10718 (N_10718,N_9631,N_9397);
xor U10719 (N_10719,N_9675,N_9913);
xnor U10720 (N_10720,N_9737,N_9014);
nor U10721 (N_10721,N_9240,N_9897);
xnor U10722 (N_10722,N_9668,N_9277);
or U10723 (N_10723,N_9393,N_9846);
or U10724 (N_10724,N_9785,N_9444);
nand U10725 (N_10725,N_9572,N_9183);
or U10726 (N_10726,N_9015,N_9023);
or U10727 (N_10727,N_9355,N_9657);
nor U10728 (N_10728,N_9462,N_9285);
nor U10729 (N_10729,N_9721,N_9219);
and U10730 (N_10730,N_9741,N_9585);
nand U10731 (N_10731,N_9756,N_9727);
xnor U10732 (N_10732,N_9793,N_9948);
nor U10733 (N_10733,N_9539,N_9238);
xor U10734 (N_10734,N_9909,N_9995);
and U10735 (N_10735,N_9639,N_9661);
xnor U10736 (N_10736,N_9463,N_9512);
nor U10737 (N_10737,N_9590,N_9098);
nand U10738 (N_10738,N_9493,N_9974);
and U10739 (N_10739,N_9695,N_9531);
nor U10740 (N_10740,N_9240,N_9201);
and U10741 (N_10741,N_9205,N_9535);
and U10742 (N_10742,N_9247,N_9322);
nand U10743 (N_10743,N_9552,N_9136);
nor U10744 (N_10744,N_9881,N_9903);
nor U10745 (N_10745,N_9494,N_9333);
nor U10746 (N_10746,N_9159,N_9830);
or U10747 (N_10747,N_9013,N_9389);
nand U10748 (N_10748,N_9780,N_9243);
nand U10749 (N_10749,N_9637,N_9363);
and U10750 (N_10750,N_9596,N_9321);
xnor U10751 (N_10751,N_9024,N_9856);
nor U10752 (N_10752,N_9831,N_9720);
and U10753 (N_10753,N_9207,N_9540);
and U10754 (N_10754,N_9192,N_9564);
nor U10755 (N_10755,N_9656,N_9260);
nand U10756 (N_10756,N_9825,N_9909);
and U10757 (N_10757,N_9835,N_9013);
or U10758 (N_10758,N_9328,N_9604);
and U10759 (N_10759,N_9635,N_9843);
nand U10760 (N_10760,N_9023,N_9365);
nor U10761 (N_10761,N_9120,N_9376);
and U10762 (N_10762,N_9577,N_9012);
nand U10763 (N_10763,N_9427,N_9641);
nand U10764 (N_10764,N_9543,N_9873);
nor U10765 (N_10765,N_9595,N_9813);
or U10766 (N_10766,N_9349,N_9653);
nand U10767 (N_10767,N_9285,N_9673);
or U10768 (N_10768,N_9930,N_9289);
nand U10769 (N_10769,N_9476,N_9751);
nor U10770 (N_10770,N_9482,N_9943);
xnor U10771 (N_10771,N_9988,N_9550);
and U10772 (N_10772,N_9389,N_9826);
xor U10773 (N_10773,N_9047,N_9455);
nor U10774 (N_10774,N_9991,N_9628);
or U10775 (N_10775,N_9281,N_9106);
and U10776 (N_10776,N_9043,N_9759);
or U10777 (N_10777,N_9950,N_9185);
and U10778 (N_10778,N_9710,N_9732);
and U10779 (N_10779,N_9483,N_9699);
xnor U10780 (N_10780,N_9495,N_9793);
xor U10781 (N_10781,N_9931,N_9790);
or U10782 (N_10782,N_9935,N_9613);
xor U10783 (N_10783,N_9949,N_9389);
or U10784 (N_10784,N_9572,N_9104);
or U10785 (N_10785,N_9549,N_9771);
nor U10786 (N_10786,N_9506,N_9039);
or U10787 (N_10787,N_9715,N_9789);
nor U10788 (N_10788,N_9359,N_9318);
nor U10789 (N_10789,N_9266,N_9249);
nor U10790 (N_10790,N_9681,N_9805);
nand U10791 (N_10791,N_9892,N_9839);
or U10792 (N_10792,N_9673,N_9425);
or U10793 (N_10793,N_9544,N_9101);
xnor U10794 (N_10794,N_9768,N_9128);
and U10795 (N_10795,N_9933,N_9886);
nor U10796 (N_10796,N_9422,N_9929);
nor U10797 (N_10797,N_9136,N_9752);
xor U10798 (N_10798,N_9918,N_9749);
nor U10799 (N_10799,N_9075,N_9289);
nand U10800 (N_10800,N_9520,N_9540);
xnor U10801 (N_10801,N_9660,N_9729);
and U10802 (N_10802,N_9143,N_9052);
or U10803 (N_10803,N_9361,N_9095);
and U10804 (N_10804,N_9941,N_9678);
and U10805 (N_10805,N_9872,N_9250);
or U10806 (N_10806,N_9240,N_9642);
xor U10807 (N_10807,N_9978,N_9865);
nor U10808 (N_10808,N_9068,N_9693);
or U10809 (N_10809,N_9954,N_9586);
nor U10810 (N_10810,N_9176,N_9893);
nor U10811 (N_10811,N_9341,N_9659);
and U10812 (N_10812,N_9740,N_9371);
or U10813 (N_10813,N_9215,N_9608);
nor U10814 (N_10814,N_9329,N_9811);
xnor U10815 (N_10815,N_9577,N_9690);
and U10816 (N_10816,N_9518,N_9578);
and U10817 (N_10817,N_9921,N_9176);
nand U10818 (N_10818,N_9650,N_9505);
nor U10819 (N_10819,N_9332,N_9527);
nand U10820 (N_10820,N_9877,N_9699);
and U10821 (N_10821,N_9995,N_9077);
or U10822 (N_10822,N_9934,N_9559);
nand U10823 (N_10823,N_9322,N_9104);
or U10824 (N_10824,N_9215,N_9368);
nor U10825 (N_10825,N_9012,N_9358);
and U10826 (N_10826,N_9132,N_9478);
and U10827 (N_10827,N_9466,N_9717);
or U10828 (N_10828,N_9126,N_9299);
and U10829 (N_10829,N_9165,N_9556);
or U10830 (N_10830,N_9332,N_9859);
or U10831 (N_10831,N_9298,N_9598);
xor U10832 (N_10832,N_9722,N_9261);
xnor U10833 (N_10833,N_9751,N_9973);
nor U10834 (N_10834,N_9176,N_9217);
xor U10835 (N_10835,N_9841,N_9751);
or U10836 (N_10836,N_9701,N_9112);
or U10837 (N_10837,N_9565,N_9899);
xor U10838 (N_10838,N_9087,N_9429);
nor U10839 (N_10839,N_9531,N_9352);
nand U10840 (N_10840,N_9477,N_9453);
and U10841 (N_10841,N_9545,N_9153);
xnor U10842 (N_10842,N_9153,N_9680);
or U10843 (N_10843,N_9623,N_9523);
xnor U10844 (N_10844,N_9210,N_9495);
and U10845 (N_10845,N_9019,N_9746);
nor U10846 (N_10846,N_9451,N_9323);
xnor U10847 (N_10847,N_9548,N_9419);
nand U10848 (N_10848,N_9018,N_9540);
nand U10849 (N_10849,N_9076,N_9626);
xnor U10850 (N_10850,N_9173,N_9532);
xnor U10851 (N_10851,N_9043,N_9272);
or U10852 (N_10852,N_9172,N_9868);
nand U10853 (N_10853,N_9597,N_9138);
and U10854 (N_10854,N_9191,N_9845);
and U10855 (N_10855,N_9503,N_9668);
or U10856 (N_10856,N_9049,N_9693);
xor U10857 (N_10857,N_9451,N_9846);
xor U10858 (N_10858,N_9836,N_9864);
or U10859 (N_10859,N_9945,N_9736);
and U10860 (N_10860,N_9784,N_9000);
nor U10861 (N_10861,N_9811,N_9452);
or U10862 (N_10862,N_9863,N_9608);
and U10863 (N_10863,N_9813,N_9778);
or U10864 (N_10864,N_9446,N_9113);
and U10865 (N_10865,N_9721,N_9865);
xnor U10866 (N_10866,N_9579,N_9824);
nor U10867 (N_10867,N_9225,N_9302);
and U10868 (N_10868,N_9906,N_9693);
nand U10869 (N_10869,N_9390,N_9407);
nand U10870 (N_10870,N_9469,N_9165);
nand U10871 (N_10871,N_9655,N_9899);
and U10872 (N_10872,N_9080,N_9622);
nor U10873 (N_10873,N_9159,N_9752);
xnor U10874 (N_10874,N_9123,N_9272);
xnor U10875 (N_10875,N_9683,N_9523);
and U10876 (N_10876,N_9599,N_9603);
nor U10877 (N_10877,N_9340,N_9806);
or U10878 (N_10878,N_9273,N_9586);
nor U10879 (N_10879,N_9111,N_9782);
xnor U10880 (N_10880,N_9882,N_9575);
nand U10881 (N_10881,N_9806,N_9369);
or U10882 (N_10882,N_9271,N_9398);
and U10883 (N_10883,N_9899,N_9710);
nor U10884 (N_10884,N_9555,N_9773);
or U10885 (N_10885,N_9659,N_9268);
xnor U10886 (N_10886,N_9891,N_9762);
and U10887 (N_10887,N_9859,N_9954);
or U10888 (N_10888,N_9895,N_9878);
or U10889 (N_10889,N_9203,N_9907);
nand U10890 (N_10890,N_9139,N_9120);
xor U10891 (N_10891,N_9256,N_9354);
nand U10892 (N_10892,N_9667,N_9898);
nand U10893 (N_10893,N_9599,N_9111);
nand U10894 (N_10894,N_9451,N_9063);
or U10895 (N_10895,N_9438,N_9581);
xor U10896 (N_10896,N_9679,N_9147);
or U10897 (N_10897,N_9484,N_9133);
and U10898 (N_10898,N_9955,N_9757);
nand U10899 (N_10899,N_9295,N_9298);
or U10900 (N_10900,N_9427,N_9979);
and U10901 (N_10901,N_9909,N_9067);
xor U10902 (N_10902,N_9932,N_9658);
and U10903 (N_10903,N_9455,N_9256);
nand U10904 (N_10904,N_9236,N_9543);
xnor U10905 (N_10905,N_9630,N_9088);
nand U10906 (N_10906,N_9111,N_9535);
and U10907 (N_10907,N_9466,N_9750);
xor U10908 (N_10908,N_9475,N_9043);
nor U10909 (N_10909,N_9742,N_9275);
and U10910 (N_10910,N_9853,N_9506);
nor U10911 (N_10911,N_9329,N_9619);
nand U10912 (N_10912,N_9752,N_9895);
nand U10913 (N_10913,N_9170,N_9522);
xnor U10914 (N_10914,N_9966,N_9372);
nand U10915 (N_10915,N_9881,N_9360);
or U10916 (N_10916,N_9595,N_9939);
nand U10917 (N_10917,N_9164,N_9643);
xnor U10918 (N_10918,N_9564,N_9042);
xnor U10919 (N_10919,N_9129,N_9502);
or U10920 (N_10920,N_9460,N_9483);
and U10921 (N_10921,N_9959,N_9580);
and U10922 (N_10922,N_9014,N_9837);
or U10923 (N_10923,N_9765,N_9950);
xnor U10924 (N_10924,N_9155,N_9479);
and U10925 (N_10925,N_9271,N_9472);
xor U10926 (N_10926,N_9722,N_9893);
xnor U10927 (N_10927,N_9962,N_9563);
xor U10928 (N_10928,N_9668,N_9204);
and U10929 (N_10929,N_9432,N_9593);
xnor U10930 (N_10930,N_9828,N_9259);
or U10931 (N_10931,N_9861,N_9641);
and U10932 (N_10932,N_9693,N_9308);
nor U10933 (N_10933,N_9083,N_9138);
nand U10934 (N_10934,N_9800,N_9364);
nor U10935 (N_10935,N_9540,N_9619);
nand U10936 (N_10936,N_9600,N_9755);
or U10937 (N_10937,N_9326,N_9934);
nand U10938 (N_10938,N_9663,N_9509);
nor U10939 (N_10939,N_9224,N_9115);
or U10940 (N_10940,N_9725,N_9508);
or U10941 (N_10941,N_9475,N_9542);
xor U10942 (N_10942,N_9027,N_9145);
and U10943 (N_10943,N_9807,N_9121);
nor U10944 (N_10944,N_9907,N_9389);
nand U10945 (N_10945,N_9642,N_9342);
nand U10946 (N_10946,N_9939,N_9205);
nor U10947 (N_10947,N_9570,N_9593);
and U10948 (N_10948,N_9786,N_9180);
nor U10949 (N_10949,N_9479,N_9068);
nand U10950 (N_10950,N_9673,N_9166);
nor U10951 (N_10951,N_9422,N_9116);
and U10952 (N_10952,N_9278,N_9621);
or U10953 (N_10953,N_9590,N_9217);
nand U10954 (N_10954,N_9632,N_9558);
or U10955 (N_10955,N_9188,N_9311);
nor U10956 (N_10956,N_9421,N_9064);
nand U10957 (N_10957,N_9469,N_9061);
or U10958 (N_10958,N_9156,N_9238);
nand U10959 (N_10959,N_9373,N_9557);
and U10960 (N_10960,N_9701,N_9778);
xor U10961 (N_10961,N_9323,N_9983);
nand U10962 (N_10962,N_9038,N_9736);
nand U10963 (N_10963,N_9143,N_9797);
and U10964 (N_10964,N_9297,N_9225);
xor U10965 (N_10965,N_9943,N_9104);
nand U10966 (N_10966,N_9478,N_9952);
xor U10967 (N_10967,N_9040,N_9797);
nand U10968 (N_10968,N_9007,N_9857);
nor U10969 (N_10969,N_9765,N_9305);
or U10970 (N_10970,N_9674,N_9627);
nor U10971 (N_10971,N_9422,N_9247);
nor U10972 (N_10972,N_9217,N_9800);
nand U10973 (N_10973,N_9408,N_9991);
nand U10974 (N_10974,N_9417,N_9373);
and U10975 (N_10975,N_9565,N_9454);
or U10976 (N_10976,N_9735,N_9543);
xor U10977 (N_10977,N_9681,N_9079);
nor U10978 (N_10978,N_9427,N_9813);
nor U10979 (N_10979,N_9678,N_9938);
nand U10980 (N_10980,N_9998,N_9168);
nand U10981 (N_10981,N_9871,N_9476);
nor U10982 (N_10982,N_9719,N_9276);
and U10983 (N_10983,N_9808,N_9106);
and U10984 (N_10984,N_9239,N_9340);
nor U10985 (N_10985,N_9801,N_9024);
nand U10986 (N_10986,N_9045,N_9355);
or U10987 (N_10987,N_9934,N_9170);
xor U10988 (N_10988,N_9690,N_9745);
and U10989 (N_10989,N_9675,N_9408);
nand U10990 (N_10990,N_9558,N_9569);
or U10991 (N_10991,N_9134,N_9002);
nor U10992 (N_10992,N_9682,N_9187);
or U10993 (N_10993,N_9194,N_9001);
nand U10994 (N_10994,N_9598,N_9253);
or U10995 (N_10995,N_9336,N_9369);
xnor U10996 (N_10996,N_9090,N_9336);
nand U10997 (N_10997,N_9662,N_9849);
nor U10998 (N_10998,N_9479,N_9856);
nand U10999 (N_10999,N_9483,N_9715);
and U11000 (N_11000,N_10186,N_10288);
nand U11001 (N_11001,N_10805,N_10907);
or U11002 (N_11002,N_10663,N_10716);
nor U11003 (N_11003,N_10033,N_10022);
nand U11004 (N_11004,N_10464,N_10942);
and U11005 (N_11005,N_10408,N_10654);
or U11006 (N_11006,N_10373,N_10383);
xor U11007 (N_11007,N_10324,N_10031);
or U11008 (N_11008,N_10167,N_10371);
and U11009 (N_11009,N_10447,N_10453);
nor U11010 (N_11010,N_10250,N_10061);
nand U11011 (N_11011,N_10257,N_10719);
and U11012 (N_11012,N_10018,N_10200);
nor U11013 (N_11013,N_10741,N_10897);
xor U11014 (N_11014,N_10987,N_10182);
xor U11015 (N_11015,N_10818,N_10189);
and U11016 (N_11016,N_10594,N_10670);
xnor U11017 (N_11017,N_10442,N_10041);
or U11018 (N_11018,N_10555,N_10529);
or U11019 (N_11019,N_10817,N_10019);
or U11020 (N_11020,N_10884,N_10534);
nor U11021 (N_11021,N_10160,N_10116);
xnor U11022 (N_11022,N_10432,N_10536);
xor U11023 (N_11023,N_10138,N_10227);
nor U11024 (N_11024,N_10513,N_10807);
or U11025 (N_11025,N_10332,N_10180);
nor U11026 (N_11026,N_10629,N_10397);
and U11027 (N_11027,N_10691,N_10284);
xor U11028 (N_11028,N_10633,N_10964);
nand U11029 (N_11029,N_10099,N_10561);
xnor U11030 (N_11030,N_10052,N_10708);
nand U11031 (N_11031,N_10489,N_10852);
nand U11032 (N_11032,N_10706,N_10132);
nand U11033 (N_11033,N_10007,N_10045);
nor U11034 (N_11034,N_10103,N_10488);
nor U11035 (N_11035,N_10492,N_10309);
or U11036 (N_11036,N_10532,N_10713);
nand U11037 (N_11037,N_10764,N_10806);
nor U11038 (N_11038,N_10969,N_10047);
and U11039 (N_11039,N_10171,N_10799);
xor U11040 (N_11040,N_10351,N_10552);
xnor U11041 (N_11041,N_10341,N_10715);
and U11042 (N_11042,N_10995,N_10296);
xor U11043 (N_11043,N_10692,N_10579);
or U11044 (N_11044,N_10970,N_10925);
or U11045 (N_11045,N_10350,N_10424);
nand U11046 (N_11046,N_10221,N_10889);
and U11047 (N_11047,N_10804,N_10177);
nand U11048 (N_11048,N_10725,N_10024);
nand U11049 (N_11049,N_10494,N_10270);
nor U11050 (N_11050,N_10439,N_10538);
and U11051 (N_11051,N_10123,N_10664);
and U11052 (N_11052,N_10981,N_10770);
xor U11053 (N_11053,N_10701,N_10793);
nor U11054 (N_11054,N_10300,N_10246);
nor U11055 (N_11055,N_10667,N_10237);
nand U11056 (N_11056,N_10860,N_10476);
and U11057 (N_11057,N_10172,N_10002);
nand U11058 (N_11058,N_10448,N_10611);
xnor U11059 (N_11059,N_10862,N_10721);
and U11060 (N_11060,N_10365,N_10088);
and U11061 (N_11061,N_10836,N_10185);
or U11062 (N_11062,N_10349,N_10326);
nor U11063 (N_11063,N_10990,N_10076);
xnor U11064 (N_11064,N_10812,N_10444);
xnor U11065 (N_11065,N_10802,N_10333);
nor U11066 (N_11066,N_10635,N_10268);
or U11067 (N_11067,N_10881,N_10564);
or U11068 (N_11068,N_10775,N_10891);
nor U11069 (N_11069,N_10184,N_10777);
nand U11070 (N_11070,N_10718,N_10760);
and U11071 (N_11071,N_10680,N_10780);
xnor U11072 (N_11072,N_10898,N_10584);
or U11073 (N_11073,N_10127,N_10786);
or U11074 (N_11074,N_10842,N_10146);
nand U11075 (N_11075,N_10787,N_10366);
nor U11076 (N_11076,N_10150,N_10726);
or U11077 (N_11077,N_10029,N_10866);
nor U11078 (N_11078,N_10588,N_10844);
nand U11079 (N_11079,N_10294,N_10530);
xnor U11080 (N_11080,N_10254,N_10235);
or U11081 (N_11081,N_10612,N_10875);
nand U11082 (N_11082,N_10641,N_10546);
nor U11083 (N_11083,N_10609,N_10727);
and U11084 (N_11084,N_10645,N_10559);
nand U11085 (N_11085,N_10865,N_10563);
xnor U11086 (N_11086,N_10902,N_10955);
and U11087 (N_11087,N_10650,N_10694);
nor U11088 (N_11088,N_10631,N_10810);
nand U11089 (N_11089,N_10335,N_10306);
or U11090 (N_11090,N_10414,N_10164);
and U11091 (N_11091,N_10637,N_10794);
nor U11092 (N_11092,N_10267,N_10589);
nor U11093 (N_11093,N_10143,N_10468);
or U11094 (N_11094,N_10139,N_10454);
xnor U11095 (N_11095,N_10080,N_10407);
or U11096 (N_11096,N_10573,N_10178);
nand U11097 (N_11097,N_10115,N_10443);
nor U11098 (N_11098,N_10340,N_10046);
and U11099 (N_11099,N_10560,N_10377);
or U11100 (N_11100,N_10354,N_10262);
and U11101 (N_11101,N_10642,N_10356);
or U11102 (N_11102,N_10364,N_10838);
or U11103 (N_11103,N_10922,N_10242);
and U11104 (N_11104,N_10000,N_10644);
nor U11105 (N_11105,N_10506,N_10832);
xor U11106 (N_11106,N_10361,N_10988);
nand U11107 (N_11107,N_10376,N_10370);
and U11108 (N_11108,N_10252,N_10105);
nand U11109 (N_11109,N_10910,N_10508);
xor U11110 (N_11110,N_10659,N_10077);
and U11111 (N_11111,N_10100,N_10154);
xor U11112 (N_11112,N_10729,N_10605);
and U11113 (N_11113,N_10967,N_10639);
nand U11114 (N_11114,N_10732,N_10336);
or U11115 (N_11115,N_10668,N_10089);
and U11116 (N_11116,N_10226,N_10527);
and U11117 (N_11117,N_10831,N_10916);
xnor U11118 (N_11118,N_10020,N_10820);
or U11119 (N_11119,N_10876,N_10485);
nor U11120 (N_11120,N_10429,N_10986);
nor U11121 (N_11121,N_10148,N_10894);
and U11122 (N_11122,N_10829,N_10826);
xnor U11123 (N_11123,N_10384,N_10752);
and U11124 (N_11124,N_10797,N_10434);
or U11125 (N_11125,N_10264,N_10921);
nor U11126 (N_11126,N_10827,N_10736);
and U11127 (N_11127,N_10357,N_10435);
xor U11128 (N_11128,N_10005,N_10202);
nand U11129 (N_11129,N_10582,N_10417);
nor U11130 (N_11130,N_10525,N_10369);
and U11131 (N_11131,N_10112,N_10072);
and U11132 (N_11132,N_10308,N_10545);
nor U11133 (N_11133,N_10544,N_10800);
nand U11134 (N_11134,N_10418,N_10021);
xor U11135 (N_11135,N_10950,N_10156);
nand U11136 (N_11136,N_10271,N_10325);
nor U11137 (N_11137,N_10638,N_10240);
nand U11138 (N_11138,N_10491,N_10816);
nor U11139 (N_11139,N_10445,N_10575);
nand U11140 (N_11140,N_10628,N_10699);
and U11141 (N_11141,N_10743,N_10359);
and U11142 (N_11142,N_10095,N_10220);
xor U11143 (N_11143,N_10539,N_10104);
nor U11144 (N_11144,N_10512,N_10858);
nor U11145 (N_11145,N_10859,N_10040);
and U11146 (N_11146,N_10011,N_10815);
and U11147 (N_11147,N_10710,N_10323);
or U11148 (N_11148,N_10176,N_10690);
xnor U11149 (N_11149,N_10399,N_10971);
or U11150 (N_11150,N_10431,N_10540);
nor U11151 (N_11151,N_10316,N_10574);
nor U11152 (N_11152,N_10993,N_10302);
or U11153 (N_11153,N_10460,N_10962);
xor U11154 (N_11154,N_10466,N_10170);
nand U11155 (N_11155,N_10554,N_10405);
xnor U11156 (N_11156,N_10724,N_10507);
nor U11157 (N_11157,N_10543,N_10785);
nor U11158 (N_11158,N_10600,N_10751);
xnor U11159 (N_11159,N_10303,N_10358);
nor U11160 (N_11160,N_10253,N_10697);
and U11161 (N_11161,N_10789,N_10675);
nand U11162 (N_11162,N_10698,N_10795);
and U11163 (N_11163,N_10157,N_10880);
and U11164 (N_11164,N_10051,N_10121);
nand U11165 (N_11165,N_10759,N_10854);
nand U11166 (N_11166,N_10686,N_10409);
and U11167 (N_11167,N_10017,N_10493);
nor U11168 (N_11168,N_10521,N_10678);
and U11169 (N_11169,N_10689,N_10204);
xor U11170 (N_11170,N_10839,N_10841);
xor U11171 (N_11171,N_10709,N_10965);
nor U11172 (N_11172,N_10149,N_10746);
xor U11173 (N_11173,N_10607,N_10585);
or U11174 (N_11174,N_10541,N_10661);
or U11175 (N_11175,N_10135,N_10120);
and U11176 (N_11176,N_10505,N_10931);
and U11177 (N_11177,N_10475,N_10446);
or U11178 (N_11178,N_10498,N_10763);
nor U11179 (N_11179,N_10911,N_10314);
nor U11180 (N_11180,N_10755,N_10943);
nor U11181 (N_11181,N_10030,N_10319);
nand U11182 (N_11182,N_10912,N_10671);
nand U11183 (N_11183,N_10648,N_10158);
nor U11184 (N_11184,N_10769,N_10877);
nand U11185 (N_11185,N_10878,N_10071);
xnor U11186 (N_11186,N_10627,N_10168);
xor U11187 (N_11187,N_10255,N_10307);
and U11188 (N_11188,N_10337,N_10556);
and U11189 (N_11189,N_10592,N_10963);
xor U11190 (N_11190,N_10486,N_10905);
nand U11191 (N_11191,N_10249,N_10996);
xor U11192 (N_11192,N_10700,N_10081);
and U11193 (N_11193,N_10421,N_10548);
nor U11194 (N_11194,N_10059,N_10310);
nor U11195 (N_11195,N_10871,N_10392);
nor U11196 (N_11196,N_10050,N_10433);
nor U11197 (N_11197,N_10269,N_10015);
nand U11198 (N_11198,N_10469,N_10400);
xor U11199 (N_11199,N_10590,N_10066);
and U11200 (N_11200,N_10577,N_10065);
xnor U11201 (N_11201,N_10490,N_10870);
nand U11202 (N_11202,N_10056,N_10562);
or U11203 (N_11203,N_10615,N_10390);
nor U11204 (N_11204,N_10477,N_10821);
or U11205 (N_11205,N_10145,N_10396);
or U11206 (N_11206,N_10765,N_10822);
xor U11207 (N_11207,N_10687,N_10473);
xor U11208 (N_11208,N_10274,N_10652);
nor U11209 (N_11209,N_10778,N_10796);
and U11210 (N_11210,N_10362,N_10695);
xor U11211 (N_11211,N_10212,N_10265);
nand U11212 (N_11212,N_10353,N_10133);
and U11213 (N_11213,N_10092,N_10991);
or U11214 (N_11214,N_10463,N_10461);
nor U11215 (N_11215,N_10347,N_10867);
or U11216 (N_11216,N_10224,N_10207);
xor U11217 (N_11217,N_10012,N_10956);
and U11218 (N_11218,N_10239,N_10360);
nand U11219 (N_11219,N_10944,N_10382);
nand U11220 (N_11220,N_10634,N_10228);
or U11221 (N_11221,N_10936,N_10321);
or U11222 (N_11222,N_10685,N_10756);
xnor U11223 (N_11223,N_10165,N_10317);
and U11224 (N_11224,N_10674,N_10411);
and U11225 (N_11225,N_10917,N_10613);
nand U11226 (N_11226,N_10499,N_10576);
xor U11227 (N_11227,N_10163,N_10580);
nor U11228 (N_11228,N_10487,N_10982);
or U11229 (N_11229,N_10712,N_10934);
xor U11230 (N_11230,N_10196,N_10386);
or U11231 (N_11231,N_10998,N_10295);
nor U11232 (N_11232,N_10723,N_10075);
or U11233 (N_11233,N_10125,N_10602);
xor U11234 (N_11234,N_10457,N_10372);
xnor U11235 (N_11235,N_10614,N_10924);
nor U11236 (N_11236,N_10016,N_10234);
nand U11237 (N_11237,N_10134,N_10953);
and U11238 (N_11238,N_10391,N_10984);
nor U11239 (N_11239,N_10216,N_10599);
or U11240 (N_11240,N_10049,N_10043);
or U11241 (N_11241,N_10624,N_10586);
or U11242 (N_11242,N_10482,N_10162);
or U11243 (N_11243,N_10329,N_10437);
and U11244 (N_11244,N_10110,N_10042);
nor U11245 (N_11245,N_10893,N_10923);
or U11246 (N_11246,N_10063,N_10259);
xor U11247 (N_11247,N_10304,N_10179);
xnor U11248 (N_11248,N_10245,N_10209);
and U11249 (N_11249,N_10853,N_10960);
or U11250 (N_11250,N_10501,N_10722);
or U11251 (N_11251,N_10792,N_10553);
nand U11252 (N_11252,N_10436,N_10027);
nand U11253 (N_11253,N_10683,N_10869);
and U11254 (N_11254,N_10261,N_10322);
xor U11255 (N_11255,N_10658,N_10904);
or U11256 (N_11256,N_10583,N_10684);
and U11257 (N_11257,N_10900,N_10819);
nor U11258 (N_11258,N_10291,N_10717);
xor U11259 (N_11259,N_10345,N_10846);
xor U11260 (N_11260,N_10260,N_10616);
or U11261 (N_11261,N_10828,N_10626);
and U11262 (N_11262,N_10714,N_10834);
nor U11263 (N_11263,N_10899,N_10211);
nor U11264 (N_11264,N_10951,N_10208);
xor U11265 (N_11265,N_10753,N_10484);
xor U11266 (N_11266,N_10503,N_10462);
or U11267 (N_11267,N_10620,N_10301);
or U11268 (N_11268,N_10256,N_10004);
nor U11269 (N_11269,N_10978,N_10097);
xnor U11270 (N_11270,N_10481,N_10181);
xnor U11271 (N_11271,N_10083,N_10193);
xnor U11272 (N_11272,N_10731,N_10679);
nor U11273 (N_11273,N_10281,N_10630);
or U11274 (N_11274,N_10298,N_10074);
or U11275 (N_11275,N_10772,N_10035);
or U11276 (N_11276,N_10420,N_10959);
or U11277 (N_11277,N_10008,N_10330);
and U11278 (N_11278,N_10367,N_10287);
and U11279 (N_11279,N_10976,N_10142);
and U11280 (N_11280,N_10090,N_10413);
xnor U11281 (N_11281,N_10681,N_10500);
or U11282 (N_11282,N_10161,N_10136);
xor U11283 (N_11283,N_10803,N_10060);
nor U11284 (N_11284,N_10926,N_10087);
and U11285 (N_11285,N_10096,N_10937);
or U11286 (N_11286,N_10705,N_10428);
xnor U11287 (N_11287,N_10954,N_10975);
and U11288 (N_11288,N_10379,N_10696);
nand U11289 (N_11289,N_10669,N_10283);
nand U11290 (N_11290,N_10510,N_10102);
and U11291 (N_11291,N_10915,N_10174);
nand U11292 (N_11292,N_10551,N_10604);
or U11293 (N_11293,N_10702,N_10311);
nor U11294 (N_11294,N_10666,N_10275);
nor U11295 (N_11295,N_10847,N_10655);
and U11296 (N_11296,N_10999,N_10788);
xor U11297 (N_11297,N_10130,N_10006);
nor U11298 (N_11298,N_10251,N_10968);
xor U11299 (N_11299,N_10427,N_10054);
nor U11300 (N_11300,N_10459,N_10547);
nand U11301 (N_11301,N_10974,N_10286);
xor U11302 (N_11302,N_10749,N_10825);
and U11303 (N_11303,N_10814,N_10153);
nor U11304 (N_11304,N_10032,N_10879);
and U11305 (N_11305,N_10338,N_10124);
and U11306 (N_11306,N_10273,N_10385);
xnor U11307 (N_11307,N_10791,N_10906);
and U11308 (N_11308,N_10992,N_10704);
nor U11309 (N_11309,N_10868,N_10901);
nor U11310 (N_11310,N_10219,N_10450);
xor U11311 (N_11311,N_10334,N_10522);
xnor U11312 (N_11312,N_10199,N_10243);
nand U11313 (N_11313,N_10375,N_10773);
xor U11314 (N_11314,N_10069,N_10835);
xor U11315 (N_11315,N_10416,N_10518);
nor U11316 (N_11316,N_10389,N_10619);
nand U11317 (N_11317,N_10587,N_10890);
nand U11318 (N_11318,N_10232,N_10997);
nand U11319 (N_11319,N_10079,N_10929);
nand U11320 (N_11320,N_10107,N_10531);
xor U11321 (N_11321,N_10504,N_10412);
nor U11322 (N_11322,N_10394,N_10374);
xor U11323 (N_11323,N_10151,N_10315);
nand U11324 (N_11324,N_10779,N_10528);
or U11325 (N_11325,N_10225,N_10938);
xor U11326 (N_11326,N_10423,N_10872);
xor U11327 (N_11327,N_10676,N_10214);
or U11328 (N_11328,N_10078,N_10415);
nor U11329 (N_11329,N_10744,N_10402);
or U11330 (N_11330,N_10001,N_10034);
xor U11331 (N_11331,N_10848,N_10387);
or U11332 (N_11332,N_10187,N_10567);
and U11333 (N_11333,N_10811,N_10966);
xnor U11334 (N_11334,N_10010,N_10622);
or U11335 (N_11335,N_10958,N_10989);
or U11336 (N_11336,N_10571,N_10277);
and U11337 (N_11337,N_10194,N_10569);
nand U11338 (N_11338,N_10651,N_10173);
and U11339 (N_11339,N_10057,N_10280);
and U11340 (N_11340,N_10426,N_10217);
nand U11341 (N_11341,N_10798,N_10119);
and U11342 (N_11342,N_10205,N_10578);
and U11343 (N_11343,N_10215,N_10781);
and U11344 (N_11344,N_10932,N_10738);
nor U11345 (N_11345,N_10857,N_10980);
nor U11346 (N_11346,N_10355,N_10098);
xor U11347 (N_11347,N_10688,N_10363);
nor U11348 (N_11348,N_10851,N_10550);
nor U11349 (N_11349,N_10084,N_10840);
nand U11350 (N_11350,N_10276,N_10058);
xnor U11351 (N_11351,N_10919,N_10048);
nor U11352 (N_11352,N_10159,N_10483);
or U11353 (N_11353,N_10126,N_10014);
nand U11354 (N_11354,N_10094,N_10085);
xnor U11355 (N_11355,N_10197,N_10762);
xnor U11356 (N_11356,N_10526,N_10175);
nor U11357 (N_11357,N_10597,N_10203);
nand U11358 (N_11358,N_10313,N_10013);
or U11359 (N_11359,N_10452,N_10509);
or U11360 (N_11360,N_10711,N_10758);
nand U11361 (N_11361,N_10737,N_10037);
xnor U11362 (N_11362,N_10557,N_10632);
and U11363 (N_11363,N_10470,N_10122);
xnor U11364 (N_11364,N_10598,N_10750);
nand U11365 (N_11365,N_10813,N_10909);
xnor U11366 (N_11366,N_10824,N_10983);
and U11367 (N_11367,N_10318,N_10863);
nand U11368 (N_11368,N_10038,N_10745);
xor U11369 (N_11369,N_10730,N_10946);
and U11370 (N_11370,N_10266,N_10272);
and U11371 (N_11371,N_10401,N_10113);
nand U11372 (N_11372,N_10480,N_10774);
and U11373 (N_11373,N_10728,N_10053);
xor U11374 (N_11374,N_10742,N_10026);
and U11375 (N_11375,N_10449,N_10809);
nor U11376 (N_11376,N_10368,N_10129);
and U11377 (N_11377,N_10570,N_10327);
or U11378 (N_11378,N_10673,N_10381);
or U11379 (N_11379,N_10144,N_10640);
and U11380 (N_11380,N_10662,N_10665);
nand U11381 (N_11381,N_10137,N_10948);
nand U11382 (N_11382,N_10636,N_10343);
nor U11383 (N_11383,N_10610,N_10591);
nand U11384 (N_11384,N_10918,N_10601);
xnor U11385 (N_11385,N_10395,N_10055);
or U11386 (N_11386,N_10761,N_10947);
nor U11387 (N_11387,N_10348,N_10537);
or U11388 (N_11388,N_10278,N_10896);
nor U11389 (N_11389,N_10913,N_10106);
nand U11390 (N_11390,N_10109,N_10344);
xor U11391 (N_11391,N_10198,N_10244);
nor U11392 (N_11392,N_10767,N_10352);
xor U11393 (N_11393,N_10771,N_10542);
nand U11394 (N_11394,N_10025,N_10776);
and U11395 (N_11395,N_10028,N_10398);
or U11396 (N_11396,N_10784,N_10707);
nor U11397 (N_11397,N_10801,N_10682);
nor U11398 (N_11398,N_10523,N_10617);
nor U11399 (N_11399,N_10258,N_10519);
or U11400 (N_11400,N_10908,N_10191);
nor U11401 (N_11401,N_10430,N_10843);
nand U11402 (N_11402,N_10914,N_10155);
and U11403 (N_11403,N_10141,N_10930);
nor U11404 (N_11404,N_10380,N_10419);
nand U11405 (N_11405,N_10920,N_10068);
xor U11406 (N_11406,N_10091,N_10928);
nor U11407 (N_11407,N_10720,N_10093);
xnor U11408 (N_11408,N_10593,N_10305);
and U11409 (N_11409,N_10247,N_10734);
nand U11410 (N_11410,N_10236,N_10933);
xor U11411 (N_11411,N_10703,N_10935);
nand U11412 (N_11412,N_10656,N_10263);
nor U11413 (N_11413,N_10118,N_10201);
xor U11414 (N_11414,N_10210,N_10023);
xnor U11415 (N_11415,N_10192,N_10735);
nand U11416 (N_11416,N_10036,N_10467);
nand U11417 (N_11417,N_10973,N_10478);
nand U11418 (N_11418,N_10044,N_10289);
nand U11419 (N_11419,N_10515,N_10625);
xnor U11420 (N_11420,N_10535,N_10471);
nand U11421 (N_11421,N_10874,N_10949);
xnor U11422 (N_11422,N_10647,N_10108);
nor U11423 (N_11423,N_10213,N_10297);
or U11424 (N_11424,N_10514,N_10823);
xor U11425 (N_11425,N_10623,N_10495);
nand U11426 (N_11426,N_10440,N_10549);
and U11427 (N_11427,N_10882,N_10062);
and U11428 (N_11428,N_10994,N_10524);
or U11429 (N_11429,N_10406,N_10856);
and U11430 (N_11430,N_10114,N_10873);
and U11431 (N_11431,N_10940,N_10067);
xor U11432 (N_11432,N_10086,N_10238);
and U11433 (N_11433,N_10479,N_10885);
nor U11434 (N_11434,N_10581,N_10850);
and U11435 (N_11435,N_10474,N_10320);
xnor U11436 (N_11436,N_10064,N_10282);
nor U11437 (N_11437,N_10895,N_10887);
and U11438 (N_11438,N_10608,N_10606);
nand U11439 (N_11439,N_10404,N_10248);
nor U11440 (N_11440,N_10783,N_10458);
nor U11441 (N_11441,N_10952,N_10169);
xnor U11442 (N_11442,N_10766,N_10957);
nand U11443 (N_11443,N_10101,N_10422);
or U11444 (N_11444,N_10945,N_10222);
or U11445 (N_11445,N_10861,N_10939);
xor U11446 (N_11446,N_10941,N_10190);
xor U11447 (N_11447,N_10595,N_10757);
or U11448 (N_11448,N_10497,N_10533);
nand U11449 (N_11449,N_10618,N_10339);
nor U11450 (N_11450,N_10183,N_10754);
nor U11451 (N_11451,N_10849,N_10147);
or U11452 (N_11452,N_10830,N_10603);
nor U11453 (N_11453,N_10672,N_10231);
and U11454 (N_11454,N_10128,N_10378);
nor U11455 (N_11455,N_10502,N_10566);
and U11456 (N_11456,N_10233,N_10733);
nor U11457 (N_11457,N_10790,N_10342);
or U11458 (N_11458,N_10845,N_10328);
and U11459 (N_11459,N_10388,N_10438);
xor U11460 (N_11460,N_10808,N_10410);
xor U11461 (N_11461,N_10039,N_10003);
nand U11462 (N_11462,N_10070,N_10346);
or U11463 (N_11463,N_10782,N_10596);
nand U11464 (N_11464,N_10961,N_10864);
xnor U11465 (N_11465,N_10886,N_10451);
or U11466 (N_11466,N_10568,N_10441);
and U11467 (N_11467,N_10520,N_10166);
or U11468 (N_11468,N_10140,N_10677);
and U11469 (N_11469,N_10511,N_10279);
nor U11470 (N_11470,N_10455,N_10456);
and U11471 (N_11471,N_10985,N_10855);
nand U11472 (N_11472,N_10572,N_10285);
or U11473 (N_11473,N_10747,N_10903);
or U11474 (N_11474,N_10290,N_10206);
nand U11475 (N_11475,N_10657,N_10496);
xor U11476 (N_11476,N_10565,N_10293);
or U11477 (N_11477,N_10229,N_10393);
and U11478 (N_11478,N_10517,N_10425);
nand U11479 (N_11479,N_10888,N_10465);
and U11480 (N_11480,N_10740,N_10621);
nor U11481 (N_11481,N_10837,N_10009);
or U11482 (N_11482,N_10073,N_10241);
nor U11483 (N_11483,N_10082,N_10117);
and U11484 (N_11484,N_10472,N_10748);
and U11485 (N_11485,N_10218,N_10299);
nand U11486 (N_11486,N_10312,N_10979);
and U11487 (N_11487,N_10643,N_10152);
nand U11488 (N_11488,N_10927,N_10131);
nor U11489 (N_11489,N_10649,N_10977);
xor U11490 (N_11490,N_10195,N_10558);
or U11491 (N_11491,N_10111,N_10188);
nand U11492 (N_11492,N_10768,N_10646);
or U11493 (N_11493,N_10223,N_10516);
nor U11494 (N_11494,N_10660,N_10292);
nor U11495 (N_11495,N_10972,N_10833);
or U11496 (N_11496,N_10403,N_10883);
or U11497 (N_11497,N_10739,N_10892);
and U11498 (N_11498,N_10693,N_10230);
nand U11499 (N_11499,N_10653,N_10331);
nor U11500 (N_11500,N_10852,N_10831);
and U11501 (N_11501,N_10611,N_10725);
and U11502 (N_11502,N_10226,N_10090);
nand U11503 (N_11503,N_10078,N_10955);
nand U11504 (N_11504,N_10086,N_10020);
or U11505 (N_11505,N_10306,N_10654);
or U11506 (N_11506,N_10489,N_10299);
xor U11507 (N_11507,N_10560,N_10005);
or U11508 (N_11508,N_10323,N_10921);
and U11509 (N_11509,N_10161,N_10783);
and U11510 (N_11510,N_10485,N_10566);
or U11511 (N_11511,N_10829,N_10601);
xnor U11512 (N_11512,N_10950,N_10048);
and U11513 (N_11513,N_10564,N_10068);
and U11514 (N_11514,N_10810,N_10241);
nand U11515 (N_11515,N_10922,N_10490);
nor U11516 (N_11516,N_10340,N_10604);
xor U11517 (N_11517,N_10382,N_10718);
nand U11518 (N_11518,N_10834,N_10292);
nor U11519 (N_11519,N_10668,N_10845);
and U11520 (N_11520,N_10085,N_10003);
xnor U11521 (N_11521,N_10029,N_10419);
and U11522 (N_11522,N_10439,N_10567);
nor U11523 (N_11523,N_10971,N_10404);
nand U11524 (N_11524,N_10419,N_10346);
and U11525 (N_11525,N_10583,N_10520);
and U11526 (N_11526,N_10798,N_10199);
xnor U11527 (N_11527,N_10229,N_10234);
nor U11528 (N_11528,N_10482,N_10554);
nor U11529 (N_11529,N_10699,N_10149);
nor U11530 (N_11530,N_10264,N_10520);
or U11531 (N_11531,N_10347,N_10838);
nor U11532 (N_11532,N_10182,N_10544);
xnor U11533 (N_11533,N_10265,N_10403);
nand U11534 (N_11534,N_10075,N_10822);
xnor U11535 (N_11535,N_10655,N_10587);
or U11536 (N_11536,N_10633,N_10779);
nor U11537 (N_11537,N_10905,N_10275);
and U11538 (N_11538,N_10768,N_10170);
xnor U11539 (N_11539,N_10201,N_10612);
and U11540 (N_11540,N_10954,N_10647);
nand U11541 (N_11541,N_10173,N_10370);
and U11542 (N_11542,N_10093,N_10320);
or U11543 (N_11543,N_10048,N_10069);
and U11544 (N_11544,N_10286,N_10387);
and U11545 (N_11545,N_10150,N_10566);
xor U11546 (N_11546,N_10096,N_10186);
or U11547 (N_11547,N_10163,N_10922);
xor U11548 (N_11548,N_10785,N_10122);
and U11549 (N_11549,N_10909,N_10065);
and U11550 (N_11550,N_10777,N_10073);
nor U11551 (N_11551,N_10192,N_10333);
nor U11552 (N_11552,N_10234,N_10983);
and U11553 (N_11553,N_10346,N_10113);
and U11554 (N_11554,N_10821,N_10558);
nand U11555 (N_11555,N_10096,N_10249);
xnor U11556 (N_11556,N_10020,N_10435);
nor U11557 (N_11557,N_10763,N_10883);
nand U11558 (N_11558,N_10076,N_10134);
nand U11559 (N_11559,N_10422,N_10976);
or U11560 (N_11560,N_10492,N_10192);
or U11561 (N_11561,N_10959,N_10564);
or U11562 (N_11562,N_10029,N_10601);
xnor U11563 (N_11563,N_10361,N_10453);
or U11564 (N_11564,N_10939,N_10060);
nand U11565 (N_11565,N_10532,N_10108);
nor U11566 (N_11566,N_10573,N_10082);
nand U11567 (N_11567,N_10774,N_10313);
nand U11568 (N_11568,N_10274,N_10924);
nand U11569 (N_11569,N_10515,N_10939);
and U11570 (N_11570,N_10345,N_10845);
and U11571 (N_11571,N_10491,N_10537);
nor U11572 (N_11572,N_10622,N_10718);
or U11573 (N_11573,N_10720,N_10965);
xnor U11574 (N_11574,N_10343,N_10576);
nor U11575 (N_11575,N_10141,N_10982);
and U11576 (N_11576,N_10355,N_10429);
xnor U11577 (N_11577,N_10936,N_10755);
xor U11578 (N_11578,N_10647,N_10973);
or U11579 (N_11579,N_10389,N_10878);
or U11580 (N_11580,N_10483,N_10761);
and U11581 (N_11581,N_10667,N_10045);
and U11582 (N_11582,N_10820,N_10022);
and U11583 (N_11583,N_10757,N_10079);
or U11584 (N_11584,N_10588,N_10379);
nand U11585 (N_11585,N_10554,N_10884);
and U11586 (N_11586,N_10231,N_10465);
and U11587 (N_11587,N_10009,N_10077);
nand U11588 (N_11588,N_10551,N_10928);
or U11589 (N_11589,N_10692,N_10980);
and U11590 (N_11590,N_10466,N_10641);
nor U11591 (N_11591,N_10007,N_10525);
nor U11592 (N_11592,N_10327,N_10209);
and U11593 (N_11593,N_10999,N_10863);
nand U11594 (N_11594,N_10741,N_10643);
and U11595 (N_11595,N_10914,N_10933);
xnor U11596 (N_11596,N_10424,N_10233);
xor U11597 (N_11597,N_10424,N_10275);
xor U11598 (N_11598,N_10036,N_10162);
nor U11599 (N_11599,N_10234,N_10509);
xnor U11600 (N_11600,N_10162,N_10680);
nand U11601 (N_11601,N_10727,N_10092);
or U11602 (N_11602,N_10740,N_10059);
nor U11603 (N_11603,N_10125,N_10844);
xnor U11604 (N_11604,N_10641,N_10022);
nor U11605 (N_11605,N_10050,N_10821);
nor U11606 (N_11606,N_10067,N_10910);
xnor U11607 (N_11607,N_10394,N_10858);
nor U11608 (N_11608,N_10581,N_10719);
xnor U11609 (N_11609,N_10380,N_10640);
nand U11610 (N_11610,N_10420,N_10522);
and U11611 (N_11611,N_10117,N_10883);
and U11612 (N_11612,N_10999,N_10560);
and U11613 (N_11613,N_10744,N_10623);
nor U11614 (N_11614,N_10708,N_10932);
xnor U11615 (N_11615,N_10049,N_10017);
nor U11616 (N_11616,N_10236,N_10467);
and U11617 (N_11617,N_10051,N_10808);
or U11618 (N_11618,N_10586,N_10614);
xnor U11619 (N_11619,N_10443,N_10897);
nand U11620 (N_11620,N_10848,N_10611);
xnor U11621 (N_11621,N_10624,N_10812);
or U11622 (N_11622,N_10772,N_10451);
and U11623 (N_11623,N_10215,N_10282);
nor U11624 (N_11624,N_10397,N_10093);
or U11625 (N_11625,N_10281,N_10347);
xor U11626 (N_11626,N_10262,N_10857);
or U11627 (N_11627,N_10301,N_10836);
nor U11628 (N_11628,N_10329,N_10708);
and U11629 (N_11629,N_10634,N_10282);
and U11630 (N_11630,N_10450,N_10539);
nand U11631 (N_11631,N_10335,N_10199);
nand U11632 (N_11632,N_10877,N_10534);
xnor U11633 (N_11633,N_10232,N_10950);
or U11634 (N_11634,N_10368,N_10597);
or U11635 (N_11635,N_10510,N_10250);
nor U11636 (N_11636,N_10469,N_10283);
and U11637 (N_11637,N_10123,N_10477);
or U11638 (N_11638,N_10278,N_10536);
nand U11639 (N_11639,N_10767,N_10043);
or U11640 (N_11640,N_10854,N_10886);
xor U11641 (N_11641,N_10021,N_10263);
nand U11642 (N_11642,N_10079,N_10314);
nor U11643 (N_11643,N_10413,N_10164);
and U11644 (N_11644,N_10553,N_10447);
xor U11645 (N_11645,N_10811,N_10934);
or U11646 (N_11646,N_10714,N_10156);
xor U11647 (N_11647,N_10767,N_10705);
or U11648 (N_11648,N_10419,N_10509);
xor U11649 (N_11649,N_10052,N_10183);
and U11650 (N_11650,N_10166,N_10300);
xor U11651 (N_11651,N_10821,N_10552);
or U11652 (N_11652,N_10316,N_10197);
or U11653 (N_11653,N_10375,N_10071);
and U11654 (N_11654,N_10141,N_10139);
nor U11655 (N_11655,N_10210,N_10003);
xor U11656 (N_11656,N_10217,N_10556);
xnor U11657 (N_11657,N_10157,N_10774);
and U11658 (N_11658,N_10343,N_10205);
and U11659 (N_11659,N_10133,N_10886);
or U11660 (N_11660,N_10528,N_10938);
nor U11661 (N_11661,N_10662,N_10031);
and U11662 (N_11662,N_10441,N_10252);
xor U11663 (N_11663,N_10841,N_10330);
xor U11664 (N_11664,N_10412,N_10141);
nand U11665 (N_11665,N_10100,N_10227);
and U11666 (N_11666,N_10033,N_10290);
nand U11667 (N_11667,N_10904,N_10350);
or U11668 (N_11668,N_10935,N_10461);
nor U11669 (N_11669,N_10109,N_10994);
or U11670 (N_11670,N_10394,N_10075);
nand U11671 (N_11671,N_10812,N_10219);
nand U11672 (N_11672,N_10527,N_10356);
nand U11673 (N_11673,N_10485,N_10621);
or U11674 (N_11674,N_10006,N_10820);
nand U11675 (N_11675,N_10068,N_10727);
and U11676 (N_11676,N_10928,N_10351);
xnor U11677 (N_11677,N_10620,N_10266);
nor U11678 (N_11678,N_10978,N_10992);
nor U11679 (N_11679,N_10611,N_10795);
and U11680 (N_11680,N_10810,N_10623);
nand U11681 (N_11681,N_10698,N_10767);
nor U11682 (N_11682,N_10974,N_10149);
or U11683 (N_11683,N_10575,N_10211);
nand U11684 (N_11684,N_10866,N_10043);
or U11685 (N_11685,N_10278,N_10506);
and U11686 (N_11686,N_10127,N_10759);
nand U11687 (N_11687,N_10701,N_10256);
nand U11688 (N_11688,N_10912,N_10657);
nand U11689 (N_11689,N_10803,N_10298);
nand U11690 (N_11690,N_10607,N_10435);
or U11691 (N_11691,N_10800,N_10451);
xor U11692 (N_11692,N_10073,N_10678);
nor U11693 (N_11693,N_10707,N_10618);
xor U11694 (N_11694,N_10033,N_10330);
nand U11695 (N_11695,N_10909,N_10927);
or U11696 (N_11696,N_10008,N_10851);
xor U11697 (N_11697,N_10053,N_10223);
and U11698 (N_11698,N_10925,N_10162);
nand U11699 (N_11699,N_10189,N_10284);
nor U11700 (N_11700,N_10067,N_10701);
and U11701 (N_11701,N_10005,N_10292);
and U11702 (N_11702,N_10909,N_10299);
nand U11703 (N_11703,N_10642,N_10402);
xor U11704 (N_11704,N_10462,N_10072);
and U11705 (N_11705,N_10263,N_10465);
and U11706 (N_11706,N_10882,N_10037);
or U11707 (N_11707,N_10025,N_10532);
or U11708 (N_11708,N_10507,N_10472);
and U11709 (N_11709,N_10290,N_10403);
or U11710 (N_11710,N_10406,N_10469);
or U11711 (N_11711,N_10423,N_10705);
or U11712 (N_11712,N_10423,N_10625);
and U11713 (N_11713,N_10119,N_10529);
nor U11714 (N_11714,N_10717,N_10024);
and U11715 (N_11715,N_10321,N_10244);
nor U11716 (N_11716,N_10857,N_10025);
nor U11717 (N_11717,N_10485,N_10585);
xor U11718 (N_11718,N_10483,N_10284);
nand U11719 (N_11719,N_10321,N_10586);
xor U11720 (N_11720,N_10658,N_10270);
and U11721 (N_11721,N_10860,N_10192);
nand U11722 (N_11722,N_10298,N_10207);
or U11723 (N_11723,N_10292,N_10961);
and U11724 (N_11724,N_10219,N_10308);
nor U11725 (N_11725,N_10790,N_10137);
xor U11726 (N_11726,N_10645,N_10879);
nand U11727 (N_11727,N_10907,N_10112);
or U11728 (N_11728,N_10860,N_10679);
or U11729 (N_11729,N_10349,N_10804);
or U11730 (N_11730,N_10288,N_10169);
nor U11731 (N_11731,N_10921,N_10852);
xor U11732 (N_11732,N_10150,N_10542);
or U11733 (N_11733,N_10753,N_10628);
or U11734 (N_11734,N_10563,N_10790);
and U11735 (N_11735,N_10002,N_10091);
xor U11736 (N_11736,N_10316,N_10521);
nor U11737 (N_11737,N_10907,N_10815);
and U11738 (N_11738,N_10081,N_10734);
nand U11739 (N_11739,N_10311,N_10915);
and U11740 (N_11740,N_10597,N_10779);
and U11741 (N_11741,N_10711,N_10993);
nand U11742 (N_11742,N_10906,N_10748);
xor U11743 (N_11743,N_10905,N_10392);
nor U11744 (N_11744,N_10609,N_10461);
nand U11745 (N_11745,N_10629,N_10128);
or U11746 (N_11746,N_10221,N_10337);
nand U11747 (N_11747,N_10583,N_10370);
or U11748 (N_11748,N_10399,N_10719);
nor U11749 (N_11749,N_10802,N_10756);
or U11750 (N_11750,N_10769,N_10013);
or U11751 (N_11751,N_10348,N_10401);
xnor U11752 (N_11752,N_10627,N_10913);
and U11753 (N_11753,N_10990,N_10285);
nand U11754 (N_11754,N_10011,N_10327);
or U11755 (N_11755,N_10147,N_10210);
nor U11756 (N_11756,N_10957,N_10271);
or U11757 (N_11757,N_10466,N_10964);
nor U11758 (N_11758,N_10603,N_10581);
nor U11759 (N_11759,N_10065,N_10328);
or U11760 (N_11760,N_10571,N_10094);
nor U11761 (N_11761,N_10274,N_10766);
or U11762 (N_11762,N_10876,N_10067);
nor U11763 (N_11763,N_10669,N_10058);
nor U11764 (N_11764,N_10620,N_10319);
nor U11765 (N_11765,N_10783,N_10897);
nor U11766 (N_11766,N_10106,N_10693);
nand U11767 (N_11767,N_10330,N_10032);
or U11768 (N_11768,N_10711,N_10544);
nand U11769 (N_11769,N_10410,N_10019);
xor U11770 (N_11770,N_10544,N_10479);
xor U11771 (N_11771,N_10466,N_10180);
nor U11772 (N_11772,N_10918,N_10186);
or U11773 (N_11773,N_10403,N_10591);
nand U11774 (N_11774,N_10113,N_10433);
and U11775 (N_11775,N_10340,N_10913);
xnor U11776 (N_11776,N_10304,N_10768);
nor U11777 (N_11777,N_10197,N_10162);
nand U11778 (N_11778,N_10639,N_10811);
and U11779 (N_11779,N_10757,N_10164);
or U11780 (N_11780,N_10008,N_10898);
and U11781 (N_11781,N_10519,N_10376);
xor U11782 (N_11782,N_10684,N_10666);
or U11783 (N_11783,N_10412,N_10448);
nor U11784 (N_11784,N_10003,N_10470);
and U11785 (N_11785,N_10560,N_10775);
or U11786 (N_11786,N_10828,N_10034);
xnor U11787 (N_11787,N_10195,N_10987);
xnor U11788 (N_11788,N_10212,N_10670);
xor U11789 (N_11789,N_10983,N_10734);
nand U11790 (N_11790,N_10487,N_10269);
or U11791 (N_11791,N_10871,N_10549);
xor U11792 (N_11792,N_10355,N_10395);
nor U11793 (N_11793,N_10626,N_10034);
and U11794 (N_11794,N_10904,N_10484);
and U11795 (N_11795,N_10483,N_10144);
nand U11796 (N_11796,N_10313,N_10983);
and U11797 (N_11797,N_10810,N_10116);
nor U11798 (N_11798,N_10272,N_10004);
xor U11799 (N_11799,N_10389,N_10765);
and U11800 (N_11800,N_10726,N_10085);
nor U11801 (N_11801,N_10621,N_10504);
xnor U11802 (N_11802,N_10385,N_10010);
nor U11803 (N_11803,N_10422,N_10157);
nand U11804 (N_11804,N_10623,N_10840);
or U11805 (N_11805,N_10200,N_10341);
nor U11806 (N_11806,N_10283,N_10050);
or U11807 (N_11807,N_10932,N_10003);
or U11808 (N_11808,N_10648,N_10830);
nor U11809 (N_11809,N_10635,N_10370);
nor U11810 (N_11810,N_10522,N_10764);
nand U11811 (N_11811,N_10366,N_10701);
xor U11812 (N_11812,N_10954,N_10464);
and U11813 (N_11813,N_10112,N_10915);
nor U11814 (N_11814,N_10648,N_10564);
or U11815 (N_11815,N_10992,N_10189);
or U11816 (N_11816,N_10981,N_10084);
nand U11817 (N_11817,N_10915,N_10497);
or U11818 (N_11818,N_10976,N_10607);
xnor U11819 (N_11819,N_10593,N_10548);
nor U11820 (N_11820,N_10850,N_10220);
nor U11821 (N_11821,N_10366,N_10509);
nand U11822 (N_11822,N_10688,N_10908);
or U11823 (N_11823,N_10948,N_10623);
or U11824 (N_11824,N_10330,N_10043);
or U11825 (N_11825,N_10436,N_10751);
xnor U11826 (N_11826,N_10142,N_10510);
xnor U11827 (N_11827,N_10849,N_10608);
or U11828 (N_11828,N_10524,N_10939);
nor U11829 (N_11829,N_10024,N_10307);
nand U11830 (N_11830,N_10541,N_10218);
and U11831 (N_11831,N_10607,N_10343);
or U11832 (N_11832,N_10729,N_10558);
and U11833 (N_11833,N_10922,N_10272);
nand U11834 (N_11834,N_10797,N_10725);
or U11835 (N_11835,N_10782,N_10236);
nor U11836 (N_11836,N_10349,N_10445);
nand U11837 (N_11837,N_10471,N_10757);
xnor U11838 (N_11838,N_10361,N_10640);
nor U11839 (N_11839,N_10110,N_10881);
nand U11840 (N_11840,N_10878,N_10230);
nand U11841 (N_11841,N_10547,N_10262);
nand U11842 (N_11842,N_10145,N_10810);
xnor U11843 (N_11843,N_10931,N_10377);
and U11844 (N_11844,N_10026,N_10638);
xor U11845 (N_11845,N_10079,N_10574);
nand U11846 (N_11846,N_10581,N_10398);
nand U11847 (N_11847,N_10135,N_10880);
xor U11848 (N_11848,N_10070,N_10750);
nor U11849 (N_11849,N_10851,N_10390);
and U11850 (N_11850,N_10456,N_10656);
xor U11851 (N_11851,N_10187,N_10457);
xnor U11852 (N_11852,N_10491,N_10225);
xnor U11853 (N_11853,N_10426,N_10972);
nand U11854 (N_11854,N_10520,N_10977);
nor U11855 (N_11855,N_10746,N_10080);
nor U11856 (N_11856,N_10140,N_10379);
nor U11857 (N_11857,N_10257,N_10792);
xor U11858 (N_11858,N_10204,N_10470);
or U11859 (N_11859,N_10778,N_10365);
and U11860 (N_11860,N_10381,N_10558);
xnor U11861 (N_11861,N_10834,N_10002);
or U11862 (N_11862,N_10526,N_10152);
nor U11863 (N_11863,N_10488,N_10078);
nand U11864 (N_11864,N_10219,N_10075);
and U11865 (N_11865,N_10791,N_10728);
and U11866 (N_11866,N_10239,N_10151);
and U11867 (N_11867,N_10438,N_10018);
xnor U11868 (N_11868,N_10406,N_10051);
xnor U11869 (N_11869,N_10731,N_10928);
or U11870 (N_11870,N_10801,N_10406);
and U11871 (N_11871,N_10024,N_10277);
xnor U11872 (N_11872,N_10525,N_10860);
nand U11873 (N_11873,N_10974,N_10978);
or U11874 (N_11874,N_10070,N_10828);
xor U11875 (N_11875,N_10960,N_10579);
nor U11876 (N_11876,N_10549,N_10080);
nor U11877 (N_11877,N_10940,N_10618);
xnor U11878 (N_11878,N_10583,N_10806);
and U11879 (N_11879,N_10494,N_10114);
nand U11880 (N_11880,N_10573,N_10272);
nand U11881 (N_11881,N_10479,N_10487);
and U11882 (N_11882,N_10191,N_10784);
xnor U11883 (N_11883,N_10703,N_10645);
and U11884 (N_11884,N_10791,N_10914);
and U11885 (N_11885,N_10577,N_10284);
xnor U11886 (N_11886,N_10532,N_10038);
or U11887 (N_11887,N_10506,N_10610);
nand U11888 (N_11888,N_10304,N_10835);
xnor U11889 (N_11889,N_10476,N_10989);
xnor U11890 (N_11890,N_10256,N_10499);
or U11891 (N_11891,N_10761,N_10486);
or U11892 (N_11892,N_10562,N_10475);
or U11893 (N_11893,N_10786,N_10495);
nor U11894 (N_11894,N_10002,N_10743);
and U11895 (N_11895,N_10471,N_10012);
nor U11896 (N_11896,N_10786,N_10288);
nand U11897 (N_11897,N_10940,N_10551);
xor U11898 (N_11898,N_10972,N_10625);
nor U11899 (N_11899,N_10899,N_10143);
or U11900 (N_11900,N_10103,N_10897);
nor U11901 (N_11901,N_10991,N_10353);
xnor U11902 (N_11902,N_10134,N_10351);
and U11903 (N_11903,N_10857,N_10496);
nand U11904 (N_11904,N_10323,N_10629);
or U11905 (N_11905,N_10315,N_10605);
nor U11906 (N_11906,N_10048,N_10082);
nand U11907 (N_11907,N_10660,N_10131);
nand U11908 (N_11908,N_10642,N_10079);
or U11909 (N_11909,N_10941,N_10800);
and U11910 (N_11910,N_10196,N_10783);
and U11911 (N_11911,N_10096,N_10873);
or U11912 (N_11912,N_10229,N_10461);
xnor U11913 (N_11913,N_10069,N_10990);
nand U11914 (N_11914,N_10002,N_10915);
nor U11915 (N_11915,N_10961,N_10274);
nor U11916 (N_11916,N_10054,N_10044);
nand U11917 (N_11917,N_10446,N_10734);
xor U11918 (N_11918,N_10939,N_10588);
nand U11919 (N_11919,N_10980,N_10102);
nand U11920 (N_11920,N_10481,N_10733);
nor U11921 (N_11921,N_10535,N_10170);
nor U11922 (N_11922,N_10046,N_10979);
nor U11923 (N_11923,N_10847,N_10121);
and U11924 (N_11924,N_10427,N_10619);
or U11925 (N_11925,N_10216,N_10781);
xor U11926 (N_11926,N_10680,N_10428);
and U11927 (N_11927,N_10747,N_10546);
or U11928 (N_11928,N_10930,N_10979);
or U11929 (N_11929,N_10365,N_10218);
and U11930 (N_11930,N_10972,N_10010);
nor U11931 (N_11931,N_10415,N_10456);
xor U11932 (N_11932,N_10434,N_10012);
xnor U11933 (N_11933,N_10629,N_10799);
nand U11934 (N_11934,N_10271,N_10328);
nand U11935 (N_11935,N_10198,N_10873);
xnor U11936 (N_11936,N_10955,N_10383);
nand U11937 (N_11937,N_10562,N_10371);
or U11938 (N_11938,N_10364,N_10423);
nor U11939 (N_11939,N_10630,N_10361);
xor U11940 (N_11940,N_10556,N_10355);
and U11941 (N_11941,N_10209,N_10983);
nor U11942 (N_11942,N_10492,N_10525);
or U11943 (N_11943,N_10464,N_10498);
xor U11944 (N_11944,N_10772,N_10201);
nor U11945 (N_11945,N_10353,N_10337);
xor U11946 (N_11946,N_10343,N_10289);
nor U11947 (N_11947,N_10442,N_10763);
xor U11948 (N_11948,N_10047,N_10668);
nor U11949 (N_11949,N_10197,N_10917);
or U11950 (N_11950,N_10237,N_10944);
nand U11951 (N_11951,N_10224,N_10800);
and U11952 (N_11952,N_10771,N_10505);
nor U11953 (N_11953,N_10529,N_10746);
and U11954 (N_11954,N_10732,N_10887);
xor U11955 (N_11955,N_10539,N_10748);
nand U11956 (N_11956,N_10485,N_10915);
nor U11957 (N_11957,N_10856,N_10481);
or U11958 (N_11958,N_10016,N_10867);
or U11959 (N_11959,N_10176,N_10379);
and U11960 (N_11960,N_10666,N_10226);
or U11961 (N_11961,N_10700,N_10472);
nand U11962 (N_11962,N_10139,N_10629);
xor U11963 (N_11963,N_10162,N_10822);
nor U11964 (N_11964,N_10995,N_10692);
nor U11965 (N_11965,N_10671,N_10925);
xnor U11966 (N_11966,N_10954,N_10603);
and U11967 (N_11967,N_10920,N_10137);
nor U11968 (N_11968,N_10466,N_10884);
xor U11969 (N_11969,N_10472,N_10873);
or U11970 (N_11970,N_10428,N_10442);
nand U11971 (N_11971,N_10111,N_10697);
or U11972 (N_11972,N_10851,N_10445);
nor U11973 (N_11973,N_10067,N_10361);
and U11974 (N_11974,N_10599,N_10905);
nor U11975 (N_11975,N_10878,N_10139);
and U11976 (N_11976,N_10358,N_10525);
nor U11977 (N_11977,N_10953,N_10940);
or U11978 (N_11978,N_10902,N_10068);
nand U11979 (N_11979,N_10245,N_10577);
nand U11980 (N_11980,N_10792,N_10493);
nor U11981 (N_11981,N_10015,N_10729);
and U11982 (N_11982,N_10152,N_10694);
nand U11983 (N_11983,N_10793,N_10855);
nor U11984 (N_11984,N_10390,N_10884);
nand U11985 (N_11985,N_10650,N_10988);
nand U11986 (N_11986,N_10184,N_10383);
nor U11987 (N_11987,N_10731,N_10564);
xor U11988 (N_11988,N_10098,N_10237);
xnor U11989 (N_11989,N_10763,N_10811);
or U11990 (N_11990,N_10478,N_10224);
nor U11991 (N_11991,N_10797,N_10387);
nor U11992 (N_11992,N_10396,N_10159);
or U11993 (N_11993,N_10201,N_10368);
or U11994 (N_11994,N_10065,N_10015);
xnor U11995 (N_11995,N_10744,N_10138);
or U11996 (N_11996,N_10796,N_10815);
and U11997 (N_11997,N_10855,N_10581);
nor U11998 (N_11998,N_10605,N_10155);
or U11999 (N_11999,N_10118,N_10070);
nand U12000 (N_12000,N_11071,N_11389);
nor U12001 (N_12001,N_11690,N_11770);
xnor U12002 (N_12002,N_11842,N_11253);
nor U12003 (N_12003,N_11487,N_11438);
or U12004 (N_12004,N_11707,N_11626);
and U12005 (N_12005,N_11476,N_11713);
or U12006 (N_12006,N_11296,N_11256);
and U12007 (N_12007,N_11555,N_11352);
nor U12008 (N_12008,N_11044,N_11001);
nor U12009 (N_12009,N_11233,N_11104);
or U12010 (N_12010,N_11709,N_11540);
and U12011 (N_12011,N_11114,N_11361);
and U12012 (N_12012,N_11754,N_11701);
and U12013 (N_12013,N_11580,N_11856);
or U12014 (N_12014,N_11246,N_11285);
and U12015 (N_12015,N_11163,N_11059);
nor U12016 (N_12016,N_11168,N_11174);
and U12017 (N_12017,N_11015,N_11683);
and U12018 (N_12018,N_11393,N_11244);
or U12019 (N_12019,N_11521,N_11971);
and U12020 (N_12020,N_11957,N_11167);
nor U12021 (N_12021,N_11060,N_11067);
xnor U12022 (N_12022,N_11264,N_11816);
and U12023 (N_12023,N_11217,N_11726);
xor U12024 (N_12024,N_11538,N_11194);
nand U12025 (N_12025,N_11496,N_11108);
and U12026 (N_12026,N_11807,N_11192);
or U12027 (N_12027,N_11095,N_11133);
nor U12028 (N_12028,N_11098,N_11252);
xor U12029 (N_12029,N_11960,N_11461);
and U12030 (N_12030,N_11371,N_11028);
nor U12031 (N_12031,N_11445,N_11877);
or U12032 (N_12032,N_11992,N_11922);
nor U12033 (N_12033,N_11815,N_11769);
nand U12034 (N_12034,N_11117,N_11785);
nand U12035 (N_12035,N_11828,N_11696);
or U12036 (N_12036,N_11952,N_11740);
nand U12037 (N_12037,N_11310,N_11148);
or U12038 (N_12038,N_11925,N_11145);
nor U12039 (N_12039,N_11153,N_11132);
and U12040 (N_12040,N_11717,N_11118);
or U12041 (N_12041,N_11034,N_11242);
and U12042 (N_12042,N_11169,N_11055);
xnor U12043 (N_12043,N_11358,N_11801);
xnor U12044 (N_12044,N_11719,N_11175);
xor U12045 (N_12045,N_11563,N_11229);
nor U12046 (N_12046,N_11356,N_11131);
xnor U12047 (N_12047,N_11613,N_11653);
xnor U12048 (N_12048,N_11560,N_11796);
nor U12049 (N_12049,N_11092,N_11574);
and U12050 (N_12050,N_11989,N_11534);
xor U12051 (N_12051,N_11604,N_11752);
or U12052 (N_12052,N_11147,N_11949);
nand U12053 (N_12053,N_11868,N_11031);
and U12054 (N_12054,N_11289,N_11235);
nor U12055 (N_12055,N_11418,N_11190);
nand U12056 (N_12056,N_11849,N_11646);
nand U12057 (N_12057,N_11890,N_11516);
or U12058 (N_12058,N_11263,N_11351);
nand U12059 (N_12059,N_11107,N_11585);
and U12060 (N_12060,N_11303,N_11799);
or U12061 (N_12061,N_11051,N_11552);
xor U12062 (N_12062,N_11512,N_11278);
xor U12063 (N_12063,N_11284,N_11616);
or U12064 (N_12064,N_11209,N_11206);
or U12065 (N_12065,N_11063,N_11058);
nor U12066 (N_12066,N_11017,N_11729);
xnor U12067 (N_12067,N_11057,N_11697);
xor U12068 (N_12068,N_11022,N_11293);
nand U12069 (N_12069,N_11249,N_11956);
xnor U12070 (N_12070,N_11724,N_11584);
and U12071 (N_12071,N_11066,N_11162);
and U12072 (N_12072,N_11020,N_11968);
or U12073 (N_12073,N_11985,N_11737);
nand U12074 (N_12074,N_11156,N_11495);
xor U12075 (N_12075,N_11323,N_11486);
or U12076 (N_12076,N_11692,N_11519);
nand U12077 (N_12077,N_11200,N_11795);
nand U12078 (N_12078,N_11914,N_11907);
xnor U12079 (N_12079,N_11536,N_11824);
nor U12080 (N_12080,N_11927,N_11197);
xor U12081 (N_12081,N_11834,N_11728);
and U12082 (N_12082,N_11331,N_11119);
xnor U12083 (N_12083,N_11670,N_11038);
and U12084 (N_12084,N_11775,N_11632);
and U12085 (N_12085,N_11172,N_11491);
or U12086 (N_12086,N_11301,N_11612);
or U12087 (N_12087,N_11561,N_11773);
nand U12088 (N_12088,N_11720,N_11892);
and U12089 (N_12089,N_11463,N_11084);
and U12090 (N_12090,N_11657,N_11618);
nor U12091 (N_12091,N_11976,N_11439);
nand U12092 (N_12092,N_11157,N_11847);
xor U12093 (N_12093,N_11441,N_11465);
nor U12094 (N_12094,N_11681,N_11558);
xnor U12095 (N_12095,N_11342,N_11528);
xor U12096 (N_12096,N_11312,N_11571);
xnor U12097 (N_12097,N_11798,N_11186);
or U12098 (N_12098,N_11745,N_11079);
and U12099 (N_12099,N_11648,N_11794);
or U12100 (N_12100,N_11429,N_11858);
nand U12101 (N_12101,N_11836,N_11718);
nand U12102 (N_12102,N_11549,N_11606);
nor U12103 (N_12103,N_11335,N_11788);
or U12104 (N_12104,N_11910,N_11865);
nand U12105 (N_12105,N_11499,N_11588);
and U12106 (N_12106,N_11838,N_11300);
and U12107 (N_12107,N_11756,N_11734);
and U12108 (N_12108,N_11755,N_11029);
nand U12109 (N_12109,N_11782,N_11710);
or U12110 (N_12110,N_11261,N_11041);
nor U12111 (N_12111,N_11193,N_11137);
nand U12112 (N_12112,N_11918,N_11639);
and U12113 (N_12113,N_11999,N_11941);
or U12114 (N_12114,N_11603,N_11048);
or U12115 (N_12115,N_11676,N_11617);
and U12116 (N_12116,N_11682,N_11140);
and U12117 (N_12117,N_11115,N_11570);
or U12118 (N_12118,N_11535,N_11384);
or U12119 (N_12119,N_11023,N_11583);
nand U12120 (N_12120,N_11056,N_11595);
nand U12121 (N_12121,N_11874,N_11725);
nand U12122 (N_12122,N_11428,N_11633);
nor U12123 (N_12123,N_11894,N_11311);
xor U12124 (N_12124,N_11344,N_11642);
nand U12125 (N_12125,N_11208,N_11074);
or U12126 (N_12126,N_11497,N_11282);
and U12127 (N_12127,N_11270,N_11884);
and U12128 (N_12128,N_11234,N_11446);
and U12129 (N_12129,N_11033,N_11030);
xor U12130 (N_12130,N_11078,N_11625);
and U12131 (N_12131,N_11018,N_11021);
or U12132 (N_12132,N_11972,N_11660);
or U12133 (N_12133,N_11929,N_11803);
xnor U12134 (N_12134,N_11183,N_11492);
nor U12135 (N_12135,N_11129,N_11665);
or U12136 (N_12136,N_11715,N_11061);
xor U12137 (N_12137,N_11346,N_11399);
and U12138 (N_12138,N_11589,N_11870);
nor U12139 (N_12139,N_11016,N_11708);
nor U12140 (N_12140,N_11759,N_11722);
nand U12141 (N_12141,N_11556,N_11494);
nor U12142 (N_12142,N_11332,N_11112);
xor U12143 (N_12143,N_11577,N_11267);
and U12144 (N_12144,N_11394,N_11731);
xnor U12145 (N_12145,N_11944,N_11327);
xor U12146 (N_12146,N_11869,N_11867);
nor U12147 (N_12147,N_11598,N_11677);
nand U12148 (N_12148,N_11631,N_11478);
and U12149 (N_12149,N_11567,N_11854);
or U12150 (N_12150,N_11473,N_11564);
nor U12151 (N_12151,N_11381,N_11784);
nand U12152 (N_12152,N_11501,N_11009);
or U12153 (N_12153,N_11550,N_11790);
or U12154 (N_12154,N_11341,N_11395);
xor U12155 (N_12155,N_11774,N_11508);
and U12156 (N_12156,N_11984,N_11184);
and U12157 (N_12157,N_11076,N_11382);
nor U12158 (N_12158,N_11374,N_11334);
nand U12159 (N_12159,N_11621,N_11666);
nand U12160 (N_12160,N_11664,N_11412);
or U12161 (N_12161,N_11266,N_11539);
nand U12162 (N_12162,N_11182,N_11291);
nor U12163 (N_12163,N_11468,N_11848);
nor U12164 (N_12164,N_11875,N_11548);
xor U12165 (N_12165,N_11171,N_11187);
and U12166 (N_12166,N_11080,N_11916);
xnor U12167 (N_12167,N_11364,N_11825);
and U12168 (N_12168,N_11414,N_11685);
nor U12169 (N_12169,N_11503,N_11687);
and U12170 (N_12170,N_11276,N_11629);
or U12171 (N_12171,N_11007,N_11202);
and U12172 (N_12172,N_11529,N_11850);
nor U12173 (N_12173,N_11191,N_11227);
or U12174 (N_12174,N_11693,N_11630);
or U12175 (N_12175,N_11897,N_11760);
and U12176 (N_12176,N_11297,N_11410);
nor U12177 (N_12177,N_11125,N_11780);
nand U12178 (N_12178,N_11421,N_11149);
or U12179 (N_12179,N_11742,N_11072);
nor U12180 (N_12180,N_11680,N_11248);
or U12181 (N_12181,N_11101,N_11950);
or U12182 (N_12182,N_11979,N_11562);
xnor U12183 (N_12183,N_11213,N_11967);
and U12184 (N_12184,N_11863,N_11111);
and U12185 (N_12185,N_11615,N_11305);
or U12186 (N_12186,N_11635,N_11531);
and U12187 (N_12187,N_11109,N_11593);
and U12188 (N_12188,N_11668,N_11872);
nor U12189 (N_12189,N_11337,N_11900);
nand U12190 (N_12190,N_11860,N_11299);
nor U12191 (N_12191,N_11886,N_11325);
nor U12192 (N_12192,N_11714,N_11005);
or U12193 (N_12193,N_11228,N_11039);
nand U12194 (N_12194,N_11262,N_11068);
nand U12195 (N_12195,N_11498,N_11982);
or U12196 (N_12196,N_11336,N_11934);
xor U12197 (N_12197,N_11753,N_11885);
nor U12198 (N_12198,N_11600,N_11442);
xor U12199 (N_12199,N_11601,N_11777);
nor U12200 (N_12200,N_11322,N_11006);
and U12201 (N_12201,N_11207,N_11765);
nand U12202 (N_12202,N_11970,N_11602);
xnor U12203 (N_12203,N_11391,N_11763);
xor U12204 (N_12204,N_11088,N_11308);
and U12205 (N_12205,N_11437,N_11185);
or U12206 (N_12206,N_11746,N_11573);
nor U12207 (N_12207,N_11320,N_11587);
nor U12208 (N_12208,N_11369,N_11673);
and U12209 (N_12209,N_11469,N_11459);
and U12210 (N_12210,N_11814,N_11081);
or U12211 (N_12211,N_11298,N_11045);
nor U12212 (N_12212,N_11678,N_11096);
or U12213 (N_12213,N_11113,N_11251);
nor U12214 (N_12214,N_11813,N_11581);
xor U12215 (N_12215,N_11732,N_11406);
or U12216 (N_12216,N_11908,N_11453);
nor U12217 (N_12217,N_11170,N_11636);
and U12218 (N_12218,N_11457,N_11811);
nand U12219 (N_12219,N_11402,N_11430);
and U12220 (N_12220,N_11180,N_11450);
nor U12221 (N_12221,N_11926,N_11808);
nand U12222 (N_12222,N_11597,N_11232);
nor U12223 (N_12223,N_11733,N_11937);
nor U12224 (N_12224,N_11490,N_11988);
nand U12225 (N_12225,N_11218,N_11160);
nor U12226 (N_12226,N_11517,N_11559);
or U12227 (N_12227,N_11757,N_11042);
xnor U12228 (N_12228,N_11372,N_11833);
nand U12229 (N_12229,N_11064,N_11974);
and U12230 (N_12230,N_11062,N_11330);
xor U12231 (N_12231,N_11103,N_11953);
or U12232 (N_12232,N_11343,N_11939);
nand U12233 (N_12233,N_11998,N_11786);
or U12234 (N_12234,N_11154,N_11087);
nand U12235 (N_12235,N_11345,N_11694);
and U12236 (N_12236,N_11400,N_11980);
or U12237 (N_12237,N_11318,N_11995);
and U12238 (N_12238,N_11628,N_11379);
xnor U12239 (N_12239,N_11879,N_11576);
nand U12240 (N_12240,N_11518,N_11515);
and U12241 (N_12241,N_11853,N_11655);
xnor U12242 (N_12242,N_11887,N_11951);
and U12243 (N_12243,N_11477,N_11317);
nand U12244 (N_12244,N_11650,N_11663);
nand U12245 (N_12245,N_11607,N_11688);
nand U12246 (N_12246,N_11532,N_11195);
nor U12247 (N_12247,N_11069,N_11314);
nand U12248 (N_12248,N_11306,N_11431);
and U12249 (N_12249,N_11324,N_11699);
or U12250 (N_12250,N_11996,N_11975);
nor U12251 (N_12251,N_11647,N_11889);
nor U12252 (N_12252,N_11407,N_11997);
nor U12253 (N_12253,N_11940,N_11810);
and U12254 (N_12254,N_11596,N_11032);
or U12255 (N_12255,N_11789,N_11387);
nor U12256 (N_12256,N_11983,N_11812);
xnor U12257 (N_12257,N_11943,N_11464);
xnor U12258 (N_12258,N_11791,N_11749);
and U12259 (N_12259,N_11241,N_11040);
nand U12260 (N_12260,N_11767,N_11027);
xnor U12261 (N_12261,N_11506,N_11474);
nor U12262 (N_12262,N_11935,N_11610);
nor U12263 (N_12263,N_11376,N_11488);
nor U12264 (N_12264,N_11166,N_11273);
or U12265 (N_12265,N_11097,N_11545);
xor U12266 (N_12266,N_11751,N_11422);
xor U12267 (N_12267,N_11649,N_11684);
nand U12268 (N_12268,N_11643,N_11843);
nand U12269 (N_12269,N_11019,N_11969);
xor U12270 (N_12270,N_11820,N_11435);
or U12271 (N_12271,N_11164,N_11313);
xor U12272 (N_12272,N_11010,N_11307);
nand U12273 (N_12273,N_11134,N_11638);
nand U12274 (N_12274,N_11954,N_11804);
nor U12275 (N_12275,N_11891,N_11522);
or U12276 (N_12276,N_11859,N_11036);
and U12277 (N_12277,N_11462,N_11100);
xor U12278 (N_12278,N_11189,N_11360);
xor U12279 (N_12279,N_11750,N_11240);
or U12280 (N_12280,N_11392,N_11130);
nand U12281 (N_12281,N_11482,N_11014);
nand U12282 (N_12282,N_11275,N_11472);
xnor U12283 (N_12283,N_11222,N_11268);
nor U12284 (N_12284,N_11321,N_11409);
and U12285 (N_12285,N_11365,N_11388);
xnor U12286 (N_12286,N_11155,N_11362);
or U12287 (N_12287,N_11964,N_11738);
and U12288 (N_12288,N_11766,N_11674);
and U12289 (N_12289,N_11523,N_11230);
and U12290 (N_12290,N_11827,N_11783);
and U12291 (N_12291,N_11931,N_11280);
nand U12292 (N_12292,N_11806,N_11420);
nand U12293 (N_12293,N_11739,N_11679);
xnor U12294 (N_12294,N_11199,N_11703);
and U12295 (N_12295,N_11883,N_11736);
xor U12296 (N_12296,N_11128,N_11257);
nand U12297 (N_12297,N_11281,N_11873);
xnor U12298 (N_12298,N_11622,N_11417);
or U12299 (N_12299,N_11893,N_11150);
xnor U12300 (N_12300,N_11711,N_11520);
nor U12301 (N_12301,N_11866,N_11375);
nor U12302 (N_12302,N_11198,N_11026);
xnor U12303 (N_12303,N_11141,N_11204);
or U12304 (N_12304,N_11861,N_11255);
or U12305 (N_12305,N_11835,N_11315);
and U12306 (N_12306,N_11695,N_11623);
nand U12307 (N_12307,N_11136,N_11764);
nor U12308 (N_12308,N_11530,N_11355);
xnor U12309 (N_12309,N_11047,N_11447);
nand U12310 (N_12310,N_11467,N_11743);
xor U12311 (N_12311,N_11912,N_11921);
and U12312 (N_12312,N_11178,N_11620);
and U12313 (N_12313,N_11254,N_11151);
or U12314 (N_12314,N_11640,N_11987);
nor U12315 (N_12315,N_11915,N_11928);
nand U12316 (N_12316,N_11747,N_11238);
nand U12317 (N_12317,N_11599,N_11906);
or U12318 (N_12318,N_11675,N_11510);
or U12319 (N_12319,N_11721,N_11043);
or U12320 (N_12320,N_11024,N_11146);
or U12321 (N_12321,N_11385,N_11543);
nor U12322 (N_12322,N_11158,N_11578);
nor U12323 (N_12323,N_11651,N_11424);
xnor U12324 (N_12324,N_11250,N_11123);
xnor U12325 (N_12325,N_11089,N_11460);
nor U12326 (N_12326,N_11142,N_11434);
xor U12327 (N_12327,N_11116,N_11046);
xnor U12328 (N_12328,N_11236,N_11401);
nor U12329 (N_12329,N_11433,N_11902);
nor U12330 (N_12330,N_11821,N_11913);
xor U12331 (N_12331,N_11053,N_11797);
xor U12332 (N_12332,N_11363,N_11102);
nand U12333 (N_12333,N_11698,N_11627);
xnor U12334 (N_12334,N_11923,N_11138);
and U12335 (N_12335,N_11511,N_11243);
xor U12336 (N_12336,N_11221,N_11544);
and U12337 (N_12337,N_11566,N_11667);
and U12338 (N_12338,N_11220,N_11702);
xor U12339 (N_12339,N_11106,N_11977);
or U12340 (N_12340,N_11004,N_11505);
nand U12341 (N_12341,N_11225,N_11288);
xor U12342 (N_12342,N_11386,N_11936);
nand U12343 (N_12343,N_11328,N_11735);
xnor U12344 (N_12344,N_11121,N_11700);
nand U12345 (N_12345,N_11052,N_11656);
xor U12346 (N_12346,N_11689,N_11212);
nor U12347 (N_12347,N_11269,N_11958);
and U12348 (N_12348,N_11159,N_11085);
nor U12349 (N_12349,N_11181,N_11978);
nor U12350 (N_12350,N_11479,N_11888);
or U12351 (N_12351,N_11366,N_11377);
or U12352 (N_12352,N_11509,N_11224);
and U12353 (N_12353,N_11819,N_11942);
nand U12354 (N_12354,N_11541,N_11619);
xor U12355 (N_12355,N_11294,N_11809);
nor U12356 (N_12356,N_11259,N_11373);
nor U12357 (N_12357,N_11223,N_11924);
nor U12358 (N_12358,N_11837,N_11654);
and U12359 (N_12359,N_11470,N_11126);
or U12360 (N_12360,N_11565,N_11831);
or U12361 (N_12361,N_11513,N_11727);
xnor U12362 (N_12362,N_11899,N_11339);
and U12363 (N_12363,N_11905,N_11994);
nand U12364 (N_12364,N_11608,N_11354);
nor U12365 (N_12365,N_11554,N_11955);
xor U12366 (N_12366,N_11082,N_11569);
or U12367 (N_12367,N_11237,N_11349);
nor U12368 (N_12368,N_11525,N_11127);
xor U12369 (N_12369,N_11920,N_11210);
nand U12370 (N_12370,N_11211,N_11265);
nand U12371 (N_12371,N_11761,N_11196);
nand U12372 (N_12372,N_11823,N_11338);
xor U12373 (N_12373,N_11938,N_11444);
xor U12374 (N_12374,N_11758,N_11839);
xnor U12375 (N_12375,N_11590,N_11882);
nand U12376 (N_12376,N_11611,N_11271);
and U12377 (N_12377,N_11398,N_11480);
xnor U12378 (N_12378,N_11652,N_11443);
xor U12379 (N_12379,N_11932,N_11832);
or U12380 (N_12380,N_11247,N_11449);
nor U12381 (N_12381,N_11177,N_11295);
or U12382 (N_12382,N_11933,N_11090);
and U12383 (N_12383,N_11049,N_11919);
or U12384 (N_12384,N_11686,N_11012);
nand U12385 (N_12385,N_11917,N_11353);
nor U12386 (N_12386,N_11909,N_11203);
or U12387 (N_12387,N_11120,N_11575);
nand U12388 (N_12388,N_11427,N_11542);
nor U12389 (N_12389,N_11368,N_11948);
or U12390 (N_12390,N_11852,N_11144);
xnor U12391 (N_12391,N_11986,N_11083);
or U12392 (N_12392,N_11864,N_11800);
nor U12393 (N_12393,N_11846,N_11286);
nand U12394 (N_12394,N_11105,N_11037);
xnor U12395 (N_12395,N_11579,N_11857);
nor U12396 (N_12396,N_11456,N_11704);
and U12397 (N_12397,N_11514,N_11292);
and U12398 (N_12398,N_11143,N_11075);
nand U12399 (N_12399,N_11035,N_11659);
nor U12400 (N_12400,N_11397,N_11871);
nand U12401 (N_12401,N_11484,N_11404);
or U12402 (N_12402,N_11452,N_11805);
or U12403 (N_12403,N_11277,N_11962);
and U12404 (N_12404,N_11179,N_11348);
or U12405 (N_12405,N_11471,N_11903);
nand U12406 (N_12406,N_11706,N_11396);
xor U12407 (N_12407,N_11904,N_11787);
nor U12408 (N_12408,N_11845,N_11245);
or U12409 (N_12409,N_11287,N_11881);
xor U12410 (N_12410,N_11025,N_11582);
nand U12411 (N_12411,N_11716,N_11500);
nor U12412 (N_12412,N_11319,N_11712);
or U12413 (N_12413,N_11408,N_11135);
xnor U12414 (N_12414,N_11781,N_11901);
and U12415 (N_12415,N_11862,N_11911);
nand U12416 (N_12416,N_11002,N_11440);
xnor U12417 (N_12417,N_11383,N_11527);
and U12418 (N_12418,N_11378,N_11013);
or U12419 (N_12419,N_11748,N_11214);
and U12420 (N_12420,N_11830,N_11551);
and U12421 (N_12421,N_11537,N_11416);
nand U12422 (N_12422,N_11415,N_11493);
or U12423 (N_12423,N_11993,N_11347);
or U12424 (N_12424,N_11231,N_11898);
xnor U12425 (N_12425,N_11855,N_11432);
nor U12426 (N_12426,N_11215,N_11403);
nor U12427 (N_12427,N_11771,N_11829);
nor U12428 (N_12428,N_11413,N_11594);
nor U12429 (N_12429,N_11634,N_11086);
xnor U12430 (N_12430,N_11475,N_11959);
and U12431 (N_12431,N_11624,N_11966);
or U12432 (N_12432,N_11637,N_11669);
nand U12433 (N_12433,N_11557,N_11454);
or U12434 (N_12434,N_11260,N_11723);
or U12435 (N_12435,N_11003,N_11099);
nor U12436 (N_12436,N_11091,N_11188);
nand U12437 (N_12437,N_11614,N_11645);
nand U12438 (N_12438,N_11981,N_11778);
and U12439 (N_12439,N_11844,N_11802);
nor U12440 (N_12440,N_11507,N_11274);
and U12441 (N_12441,N_11504,N_11572);
or U12442 (N_12442,N_11818,N_11772);
or U12443 (N_12443,N_11466,N_11122);
nand U12444 (N_12444,N_11946,N_11817);
xnor U12445 (N_12445,N_11451,N_11658);
xor U12446 (N_12446,N_11485,N_11093);
and U12447 (N_12447,N_11793,N_11405);
xnor U12448 (N_12448,N_11547,N_11841);
nand U12449 (N_12449,N_11973,N_11370);
and U12450 (N_12450,N_11489,N_11077);
nor U12451 (N_12451,N_11219,N_11546);
and U12452 (N_12452,N_11526,N_11533);
or U12453 (N_12453,N_11279,N_11768);
or U12454 (N_12454,N_11592,N_11930);
nand U12455 (N_12455,N_11609,N_11991);
or U12456 (N_12456,N_11359,N_11054);
nand U12457 (N_12457,N_11876,N_11304);
nand U12458 (N_12458,N_11990,N_11419);
nor U12459 (N_12459,N_11390,N_11380);
or U12460 (N_12460,N_11591,N_11880);
xnor U12461 (N_12461,N_11705,N_11050);
or U12462 (N_12462,N_11448,N_11309);
and U12463 (N_12463,N_11762,N_11216);
xnor U12464 (N_12464,N_11124,N_11483);
nand U12465 (N_12465,N_11329,N_11822);
xnor U12466 (N_12466,N_11436,N_11641);
or U12467 (N_12467,N_11011,N_11173);
xnor U12468 (N_12468,N_11455,N_11458);
and U12469 (N_12469,N_11662,N_11411);
nand U12470 (N_12470,N_11290,N_11316);
xnor U12471 (N_12471,N_11965,N_11094);
or U12472 (N_12472,N_11239,N_11779);
nor U12473 (N_12473,N_11840,N_11283);
and U12474 (N_12474,N_11776,N_11073);
and U12475 (N_12475,N_11426,N_11524);
and U12476 (N_12476,N_11851,N_11963);
nor U12477 (N_12477,N_11553,N_11272);
nor U12478 (N_12478,N_11502,N_11340);
nor U12479 (N_12479,N_11744,N_11730);
or U12480 (N_12480,N_11961,N_11481);
nand U12481 (N_12481,N_11333,N_11568);
nor U12482 (N_12482,N_11895,N_11226);
and U12483 (N_12483,N_11605,N_11672);
or U12484 (N_12484,N_11258,N_11201);
nor U12485 (N_12485,N_11065,N_11826);
nor U12486 (N_12486,N_11205,N_11586);
nand U12487 (N_12487,N_11070,N_11945);
nor U12488 (N_12488,N_11947,N_11176);
nand U12489 (N_12489,N_11661,N_11425);
xor U12490 (N_12490,N_11691,N_11008);
nand U12491 (N_12491,N_11161,N_11896);
nor U12492 (N_12492,N_11741,N_11165);
or U12493 (N_12493,N_11423,N_11350);
and U12494 (N_12494,N_11671,N_11000);
nor U12495 (N_12495,N_11367,N_11152);
nor U12496 (N_12496,N_11357,N_11644);
nand U12497 (N_12497,N_11878,N_11326);
nor U12498 (N_12498,N_11139,N_11792);
and U12499 (N_12499,N_11302,N_11110);
and U12500 (N_12500,N_11913,N_11517);
and U12501 (N_12501,N_11393,N_11839);
or U12502 (N_12502,N_11995,N_11854);
or U12503 (N_12503,N_11040,N_11576);
nand U12504 (N_12504,N_11717,N_11624);
and U12505 (N_12505,N_11918,N_11696);
xnor U12506 (N_12506,N_11896,N_11517);
nand U12507 (N_12507,N_11559,N_11084);
nor U12508 (N_12508,N_11303,N_11227);
or U12509 (N_12509,N_11769,N_11950);
xnor U12510 (N_12510,N_11635,N_11473);
and U12511 (N_12511,N_11176,N_11380);
or U12512 (N_12512,N_11427,N_11920);
nor U12513 (N_12513,N_11739,N_11472);
xnor U12514 (N_12514,N_11696,N_11203);
and U12515 (N_12515,N_11111,N_11310);
or U12516 (N_12516,N_11755,N_11534);
nor U12517 (N_12517,N_11932,N_11965);
and U12518 (N_12518,N_11132,N_11657);
xor U12519 (N_12519,N_11099,N_11605);
nand U12520 (N_12520,N_11612,N_11476);
or U12521 (N_12521,N_11961,N_11792);
or U12522 (N_12522,N_11709,N_11943);
nor U12523 (N_12523,N_11796,N_11009);
and U12524 (N_12524,N_11555,N_11844);
nand U12525 (N_12525,N_11899,N_11847);
nand U12526 (N_12526,N_11943,N_11619);
and U12527 (N_12527,N_11726,N_11810);
xnor U12528 (N_12528,N_11637,N_11044);
or U12529 (N_12529,N_11932,N_11499);
and U12530 (N_12530,N_11011,N_11225);
nand U12531 (N_12531,N_11531,N_11702);
or U12532 (N_12532,N_11047,N_11954);
nand U12533 (N_12533,N_11920,N_11386);
nor U12534 (N_12534,N_11524,N_11819);
nand U12535 (N_12535,N_11056,N_11512);
or U12536 (N_12536,N_11517,N_11030);
nand U12537 (N_12537,N_11912,N_11446);
or U12538 (N_12538,N_11422,N_11003);
xnor U12539 (N_12539,N_11174,N_11416);
nand U12540 (N_12540,N_11969,N_11592);
or U12541 (N_12541,N_11732,N_11934);
and U12542 (N_12542,N_11994,N_11629);
and U12543 (N_12543,N_11119,N_11565);
and U12544 (N_12544,N_11394,N_11379);
and U12545 (N_12545,N_11761,N_11208);
or U12546 (N_12546,N_11586,N_11689);
or U12547 (N_12547,N_11919,N_11339);
or U12548 (N_12548,N_11152,N_11848);
nand U12549 (N_12549,N_11908,N_11935);
nor U12550 (N_12550,N_11895,N_11373);
xor U12551 (N_12551,N_11904,N_11483);
nor U12552 (N_12552,N_11544,N_11911);
nor U12553 (N_12553,N_11245,N_11235);
or U12554 (N_12554,N_11478,N_11143);
xnor U12555 (N_12555,N_11037,N_11648);
nand U12556 (N_12556,N_11312,N_11351);
or U12557 (N_12557,N_11929,N_11131);
xor U12558 (N_12558,N_11559,N_11330);
nand U12559 (N_12559,N_11566,N_11041);
xnor U12560 (N_12560,N_11767,N_11422);
and U12561 (N_12561,N_11666,N_11067);
nor U12562 (N_12562,N_11251,N_11387);
or U12563 (N_12563,N_11779,N_11006);
nand U12564 (N_12564,N_11758,N_11014);
xor U12565 (N_12565,N_11278,N_11759);
nand U12566 (N_12566,N_11698,N_11278);
nand U12567 (N_12567,N_11495,N_11015);
nand U12568 (N_12568,N_11075,N_11733);
nand U12569 (N_12569,N_11553,N_11267);
or U12570 (N_12570,N_11080,N_11147);
nand U12571 (N_12571,N_11214,N_11393);
or U12572 (N_12572,N_11004,N_11001);
nor U12573 (N_12573,N_11783,N_11577);
and U12574 (N_12574,N_11146,N_11246);
or U12575 (N_12575,N_11640,N_11489);
nand U12576 (N_12576,N_11442,N_11520);
xnor U12577 (N_12577,N_11263,N_11392);
xor U12578 (N_12578,N_11374,N_11555);
nand U12579 (N_12579,N_11474,N_11794);
nand U12580 (N_12580,N_11085,N_11415);
and U12581 (N_12581,N_11550,N_11637);
nor U12582 (N_12582,N_11409,N_11069);
nand U12583 (N_12583,N_11551,N_11074);
nand U12584 (N_12584,N_11070,N_11806);
nor U12585 (N_12585,N_11967,N_11627);
nand U12586 (N_12586,N_11976,N_11581);
nand U12587 (N_12587,N_11243,N_11343);
nand U12588 (N_12588,N_11055,N_11776);
or U12589 (N_12589,N_11524,N_11933);
and U12590 (N_12590,N_11616,N_11091);
nand U12591 (N_12591,N_11676,N_11579);
and U12592 (N_12592,N_11535,N_11292);
nand U12593 (N_12593,N_11185,N_11521);
xnor U12594 (N_12594,N_11851,N_11582);
xnor U12595 (N_12595,N_11038,N_11085);
nand U12596 (N_12596,N_11022,N_11721);
xor U12597 (N_12597,N_11375,N_11897);
nand U12598 (N_12598,N_11353,N_11518);
nand U12599 (N_12599,N_11811,N_11921);
nand U12600 (N_12600,N_11957,N_11624);
nor U12601 (N_12601,N_11142,N_11737);
nor U12602 (N_12602,N_11617,N_11226);
or U12603 (N_12603,N_11318,N_11672);
and U12604 (N_12604,N_11642,N_11003);
nand U12605 (N_12605,N_11451,N_11984);
nor U12606 (N_12606,N_11947,N_11296);
xor U12607 (N_12607,N_11031,N_11407);
nand U12608 (N_12608,N_11575,N_11235);
or U12609 (N_12609,N_11957,N_11256);
nand U12610 (N_12610,N_11934,N_11582);
and U12611 (N_12611,N_11367,N_11938);
nand U12612 (N_12612,N_11368,N_11217);
xnor U12613 (N_12613,N_11794,N_11507);
xnor U12614 (N_12614,N_11515,N_11155);
nand U12615 (N_12615,N_11836,N_11274);
nand U12616 (N_12616,N_11399,N_11303);
xnor U12617 (N_12617,N_11532,N_11477);
nand U12618 (N_12618,N_11924,N_11671);
or U12619 (N_12619,N_11181,N_11515);
xnor U12620 (N_12620,N_11552,N_11928);
or U12621 (N_12621,N_11739,N_11699);
or U12622 (N_12622,N_11279,N_11041);
xor U12623 (N_12623,N_11596,N_11527);
xnor U12624 (N_12624,N_11570,N_11040);
nand U12625 (N_12625,N_11130,N_11055);
nor U12626 (N_12626,N_11939,N_11282);
and U12627 (N_12627,N_11436,N_11556);
and U12628 (N_12628,N_11069,N_11475);
nand U12629 (N_12629,N_11369,N_11223);
or U12630 (N_12630,N_11669,N_11382);
xor U12631 (N_12631,N_11437,N_11777);
or U12632 (N_12632,N_11492,N_11205);
nand U12633 (N_12633,N_11982,N_11566);
nand U12634 (N_12634,N_11974,N_11593);
xor U12635 (N_12635,N_11289,N_11389);
or U12636 (N_12636,N_11365,N_11444);
nor U12637 (N_12637,N_11454,N_11510);
nand U12638 (N_12638,N_11823,N_11670);
and U12639 (N_12639,N_11163,N_11684);
and U12640 (N_12640,N_11209,N_11055);
or U12641 (N_12641,N_11928,N_11270);
nor U12642 (N_12642,N_11182,N_11302);
nor U12643 (N_12643,N_11923,N_11937);
xor U12644 (N_12644,N_11982,N_11785);
nor U12645 (N_12645,N_11309,N_11797);
xnor U12646 (N_12646,N_11531,N_11550);
or U12647 (N_12647,N_11171,N_11882);
nand U12648 (N_12648,N_11639,N_11934);
nand U12649 (N_12649,N_11133,N_11262);
or U12650 (N_12650,N_11775,N_11190);
nor U12651 (N_12651,N_11410,N_11049);
nor U12652 (N_12652,N_11788,N_11001);
and U12653 (N_12653,N_11481,N_11097);
and U12654 (N_12654,N_11873,N_11892);
nand U12655 (N_12655,N_11090,N_11132);
xnor U12656 (N_12656,N_11988,N_11378);
nand U12657 (N_12657,N_11710,N_11661);
or U12658 (N_12658,N_11856,N_11044);
and U12659 (N_12659,N_11866,N_11464);
nor U12660 (N_12660,N_11757,N_11390);
nand U12661 (N_12661,N_11398,N_11617);
nand U12662 (N_12662,N_11667,N_11992);
nand U12663 (N_12663,N_11210,N_11913);
or U12664 (N_12664,N_11259,N_11021);
and U12665 (N_12665,N_11329,N_11794);
xnor U12666 (N_12666,N_11204,N_11196);
nand U12667 (N_12667,N_11167,N_11551);
or U12668 (N_12668,N_11221,N_11575);
nand U12669 (N_12669,N_11579,N_11860);
and U12670 (N_12670,N_11277,N_11183);
or U12671 (N_12671,N_11815,N_11275);
and U12672 (N_12672,N_11015,N_11445);
and U12673 (N_12673,N_11865,N_11302);
or U12674 (N_12674,N_11782,N_11607);
or U12675 (N_12675,N_11197,N_11478);
xor U12676 (N_12676,N_11062,N_11766);
or U12677 (N_12677,N_11683,N_11708);
nor U12678 (N_12678,N_11097,N_11822);
nand U12679 (N_12679,N_11925,N_11943);
or U12680 (N_12680,N_11478,N_11122);
and U12681 (N_12681,N_11998,N_11069);
nor U12682 (N_12682,N_11100,N_11753);
or U12683 (N_12683,N_11764,N_11481);
nand U12684 (N_12684,N_11553,N_11623);
nand U12685 (N_12685,N_11480,N_11505);
nor U12686 (N_12686,N_11446,N_11313);
nand U12687 (N_12687,N_11517,N_11414);
nand U12688 (N_12688,N_11253,N_11200);
nor U12689 (N_12689,N_11198,N_11563);
nor U12690 (N_12690,N_11869,N_11379);
xor U12691 (N_12691,N_11266,N_11661);
nand U12692 (N_12692,N_11941,N_11027);
xor U12693 (N_12693,N_11994,N_11515);
and U12694 (N_12694,N_11564,N_11052);
nand U12695 (N_12695,N_11981,N_11775);
and U12696 (N_12696,N_11342,N_11871);
nor U12697 (N_12697,N_11756,N_11515);
and U12698 (N_12698,N_11217,N_11611);
or U12699 (N_12699,N_11316,N_11144);
or U12700 (N_12700,N_11115,N_11465);
xnor U12701 (N_12701,N_11282,N_11778);
or U12702 (N_12702,N_11805,N_11548);
and U12703 (N_12703,N_11877,N_11853);
and U12704 (N_12704,N_11065,N_11690);
nor U12705 (N_12705,N_11162,N_11128);
or U12706 (N_12706,N_11490,N_11717);
xnor U12707 (N_12707,N_11787,N_11058);
or U12708 (N_12708,N_11677,N_11988);
nor U12709 (N_12709,N_11094,N_11055);
or U12710 (N_12710,N_11172,N_11528);
xor U12711 (N_12711,N_11553,N_11382);
nor U12712 (N_12712,N_11795,N_11273);
nor U12713 (N_12713,N_11813,N_11415);
nor U12714 (N_12714,N_11657,N_11649);
and U12715 (N_12715,N_11763,N_11815);
nand U12716 (N_12716,N_11881,N_11990);
or U12717 (N_12717,N_11257,N_11366);
nor U12718 (N_12718,N_11941,N_11898);
nand U12719 (N_12719,N_11793,N_11699);
xor U12720 (N_12720,N_11252,N_11913);
xor U12721 (N_12721,N_11357,N_11068);
nor U12722 (N_12722,N_11860,N_11380);
nand U12723 (N_12723,N_11589,N_11609);
nor U12724 (N_12724,N_11524,N_11063);
nand U12725 (N_12725,N_11599,N_11142);
nor U12726 (N_12726,N_11861,N_11134);
nor U12727 (N_12727,N_11077,N_11451);
or U12728 (N_12728,N_11686,N_11054);
xor U12729 (N_12729,N_11576,N_11719);
nor U12730 (N_12730,N_11758,N_11596);
nor U12731 (N_12731,N_11115,N_11474);
or U12732 (N_12732,N_11138,N_11694);
xor U12733 (N_12733,N_11107,N_11981);
xnor U12734 (N_12734,N_11803,N_11064);
nor U12735 (N_12735,N_11510,N_11321);
nor U12736 (N_12736,N_11063,N_11927);
nand U12737 (N_12737,N_11095,N_11557);
or U12738 (N_12738,N_11864,N_11950);
nand U12739 (N_12739,N_11357,N_11073);
and U12740 (N_12740,N_11066,N_11612);
nand U12741 (N_12741,N_11735,N_11338);
xor U12742 (N_12742,N_11560,N_11153);
nand U12743 (N_12743,N_11957,N_11412);
nand U12744 (N_12744,N_11548,N_11328);
nor U12745 (N_12745,N_11195,N_11384);
or U12746 (N_12746,N_11694,N_11562);
and U12747 (N_12747,N_11084,N_11609);
and U12748 (N_12748,N_11358,N_11824);
xor U12749 (N_12749,N_11071,N_11398);
xnor U12750 (N_12750,N_11353,N_11318);
nor U12751 (N_12751,N_11150,N_11788);
and U12752 (N_12752,N_11212,N_11581);
and U12753 (N_12753,N_11348,N_11015);
or U12754 (N_12754,N_11033,N_11557);
nor U12755 (N_12755,N_11623,N_11898);
nor U12756 (N_12756,N_11291,N_11306);
nand U12757 (N_12757,N_11937,N_11365);
or U12758 (N_12758,N_11552,N_11303);
and U12759 (N_12759,N_11715,N_11738);
nand U12760 (N_12760,N_11330,N_11968);
nor U12761 (N_12761,N_11380,N_11092);
nor U12762 (N_12762,N_11361,N_11181);
nand U12763 (N_12763,N_11095,N_11170);
and U12764 (N_12764,N_11906,N_11364);
nand U12765 (N_12765,N_11349,N_11501);
nand U12766 (N_12766,N_11651,N_11801);
nor U12767 (N_12767,N_11550,N_11854);
and U12768 (N_12768,N_11073,N_11806);
or U12769 (N_12769,N_11693,N_11145);
nor U12770 (N_12770,N_11551,N_11605);
or U12771 (N_12771,N_11246,N_11307);
xor U12772 (N_12772,N_11133,N_11342);
nand U12773 (N_12773,N_11758,N_11836);
nor U12774 (N_12774,N_11663,N_11608);
or U12775 (N_12775,N_11466,N_11022);
nor U12776 (N_12776,N_11720,N_11574);
or U12777 (N_12777,N_11775,N_11858);
and U12778 (N_12778,N_11658,N_11650);
nand U12779 (N_12779,N_11961,N_11222);
and U12780 (N_12780,N_11690,N_11837);
and U12781 (N_12781,N_11894,N_11673);
nor U12782 (N_12782,N_11944,N_11499);
xor U12783 (N_12783,N_11947,N_11608);
xor U12784 (N_12784,N_11529,N_11964);
nand U12785 (N_12785,N_11109,N_11474);
nand U12786 (N_12786,N_11074,N_11001);
nor U12787 (N_12787,N_11925,N_11295);
or U12788 (N_12788,N_11743,N_11310);
and U12789 (N_12789,N_11609,N_11957);
and U12790 (N_12790,N_11831,N_11313);
or U12791 (N_12791,N_11925,N_11690);
and U12792 (N_12792,N_11571,N_11516);
xnor U12793 (N_12793,N_11243,N_11856);
xor U12794 (N_12794,N_11839,N_11363);
xor U12795 (N_12795,N_11267,N_11876);
nand U12796 (N_12796,N_11891,N_11566);
and U12797 (N_12797,N_11052,N_11721);
nor U12798 (N_12798,N_11356,N_11052);
nand U12799 (N_12799,N_11931,N_11340);
and U12800 (N_12800,N_11317,N_11053);
or U12801 (N_12801,N_11976,N_11159);
and U12802 (N_12802,N_11309,N_11987);
or U12803 (N_12803,N_11173,N_11026);
nor U12804 (N_12804,N_11772,N_11596);
xnor U12805 (N_12805,N_11190,N_11970);
or U12806 (N_12806,N_11649,N_11050);
xnor U12807 (N_12807,N_11930,N_11645);
nand U12808 (N_12808,N_11547,N_11326);
nand U12809 (N_12809,N_11455,N_11770);
nand U12810 (N_12810,N_11438,N_11717);
nor U12811 (N_12811,N_11793,N_11018);
nor U12812 (N_12812,N_11262,N_11971);
or U12813 (N_12813,N_11334,N_11629);
nand U12814 (N_12814,N_11492,N_11040);
nor U12815 (N_12815,N_11331,N_11743);
xor U12816 (N_12816,N_11491,N_11319);
xor U12817 (N_12817,N_11712,N_11616);
and U12818 (N_12818,N_11428,N_11692);
xnor U12819 (N_12819,N_11141,N_11966);
xor U12820 (N_12820,N_11294,N_11000);
nand U12821 (N_12821,N_11769,N_11590);
or U12822 (N_12822,N_11091,N_11717);
nor U12823 (N_12823,N_11528,N_11350);
or U12824 (N_12824,N_11919,N_11496);
nand U12825 (N_12825,N_11258,N_11874);
and U12826 (N_12826,N_11390,N_11402);
xor U12827 (N_12827,N_11987,N_11824);
or U12828 (N_12828,N_11415,N_11855);
or U12829 (N_12829,N_11928,N_11835);
nand U12830 (N_12830,N_11033,N_11380);
or U12831 (N_12831,N_11408,N_11333);
or U12832 (N_12832,N_11343,N_11150);
nor U12833 (N_12833,N_11025,N_11565);
and U12834 (N_12834,N_11149,N_11725);
or U12835 (N_12835,N_11517,N_11667);
and U12836 (N_12836,N_11595,N_11273);
nand U12837 (N_12837,N_11263,N_11989);
and U12838 (N_12838,N_11579,N_11852);
or U12839 (N_12839,N_11508,N_11337);
nand U12840 (N_12840,N_11560,N_11392);
nand U12841 (N_12841,N_11987,N_11812);
or U12842 (N_12842,N_11734,N_11738);
and U12843 (N_12843,N_11059,N_11993);
and U12844 (N_12844,N_11066,N_11333);
and U12845 (N_12845,N_11626,N_11669);
and U12846 (N_12846,N_11057,N_11682);
nand U12847 (N_12847,N_11270,N_11555);
xnor U12848 (N_12848,N_11836,N_11793);
nand U12849 (N_12849,N_11998,N_11871);
nand U12850 (N_12850,N_11816,N_11930);
xor U12851 (N_12851,N_11385,N_11991);
and U12852 (N_12852,N_11234,N_11862);
xor U12853 (N_12853,N_11207,N_11536);
and U12854 (N_12854,N_11240,N_11281);
nor U12855 (N_12855,N_11595,N_11816);
nor U12856 (N_12856,N_11750,N_11951);
and U12857 (N_12857,N_11663,N_11142);
xnor U12858 (N_12858,N_11601,N_11857);
and U12859 (N_12859,N_11426,N_11515);
nand U12860 (N_12860,N_11048,N_11535);
and U12861 (N_12861,N_11167,N_11934);
or U12862 (N_12862,N_11885,N_11090);
and U12863 (N_12863,N_11827,N_11699);
nor U12864 (N_12864,N_11720,N_11843);
xor U12865 (N_12865,N_11803,N_11499);
xor U12866 (N_12866,N_11511,N_11694);
or U12867 (N_12867,N_11583,N_11613);
xor U12868 (N_12868,N_11210,N_11395);
nand U12869 (N_12869,N_11037,N_11777);
xnor U12870 (N_12870,N_11868,N_11163);
or U12871 (N_12871,N_11295,N_11672);
nand U12872 (N_12872,N_11120,N_11542);
or U12873 (N_12873,N_11413,N_11653);
and U12874 (N_12874,N_11097,N_11861);
nor U12875 (N_12875,N_11063,N_11328);
or U12876 (N_12876,N_11788,N_11246);
nor U12877 (N_12877,N_11602,N_11090);
nor U12878 (N_12878,N_11167,N_11273);
and U12879 (N_12879,N_11914,N_11481);
and U12880 (N_12880,N_11622,N_11619);
xor U12881 (N_12881,N_11264,N_11103);
or U12882 (N_12882,N_11407,N_11299);
xor U12883 (N_12883,N_11958,N_11011);
xor U12884 (N_12884,N_11450,N_11583);
nor U12885 (N_12885,N_11044,N_11204);
nor U12886 (N_12886,N_11500,N_11549);
xor U12887 (N_12887,N_11254,N_11981);
nor U12888 (N_12888,N_11593,N_11948);
nor U12889 (N_12889,N_11258,N_11953);
xnor U12890 (N_12890,N_11729,N_11327);
xnor U12891 (N_12891,N_11381,N_11221);
and U12892 (N_12892,N_11362,N_11173);
nand U12893 (N_12893,N_11174,N_11345);
or U12894 (N_12894,N_11811,N_11819);
xor U12895 (N_12895,N_11151,N_11669);
nand U12896 (N_12896,N_11128,N_11872);
xor U12897 (N_12897,N_11408,N_11756);
nor U12898 (N_12898,N_11125,N_11626);
or U12899 (N_12899,N_11954,N_11750);
nand U12900 (N_12900,N_11766,N_11296);
nand U12901 (N_12901,N_11565,N_11403);
nand U12902 (N_12902,N_11768,N_11756);
xnor U12903 (N_12903,N_11242,N_11618);
nand U12904 (N_12904,N_11902,N_11108);
nor U12905 (N_12905,N_11718,N_11189);
nor U12906 (N_12906,N_11704,N_11451);
nand U12907 (N_12907,N_11821,N_11986);
and U12908 (N_12908,N_11276,N_11014);
nand U12909 (N_12909,N_11775,N_11541);
xnor U12910 (N_12910,N_11769,N_11097);
or U12911 (N_12911,N_11395,N_11393);
nor U12912 (N_12912,N_11912,N_11717);
or U12913 (N_12913,N_11008,N_11430);
nand U12914 (N_12914,N_11865,N_11519);
nand U12915 (N_12915,N_11508,N_11329);
nor U12916 (N_12916,N_11816,N_11618);
nor U12917 (N_12917,N_11241,N_11482);
nor U12918 (N_12918,N_11304,N_11376);
nand U12919 (N_12919,N_11235,N_11613);
or U12920 (N_12920,N_11411,N_11063);
or U12921 (N_12921,N_11242,N_11230);
nor U12922 (N_12922,N_11143,N_11310);
or U12923 (N_12923,N_11070,N_11858);
and U12924 (N_12924,N_11535,N_11696);
xnor U12925 (N_12925,N_11834,N_11461);
xnor U12926 (N_12926,N_11707,N_11634);
nand U12927 (N_12927,N_11235,N_11220);
xnor U12928 (N_12928,N_11899,N_11598);
xnor U12929 (N_12929,N_11379,N_11336);
and U12930 (N_12930,N_11322,N_11670);
or U12931 (N_12931,N_11602,N_11829);
nand U12932 (N_12932,N_11179,N_11976);
nand U12933 (N_12933,N_11195,N_11988);
nand U12934 (N_12934,N_11248,N_11204);
or U12935 (N_12935,N_11929,N_11567);
xnor U12936 (N_12936,N_11736,N_11514);
xnor U12937 (N_12937,N_11318,N_11750);
and U12938 (N_12938,N_11532,N_11231);
and U12939 (N_12939,N_11773,N_11051);
nor U12940 (N_12940,N_11715,N_11060);
xnor U12941 (N_12941,N_11304,N_11863);
nand U12942 (N_12942,N_11704,N_11211);
nor U12943 (N_12943,N_11027,N_11776);
nor U12944 (N_12944,N_11547,N_11329);
and U12945 (N_12945,N_11879,N_11812);
xor U12946 (N_12946,N_11921,N_11425);
nor U12947 (N_12947,N_11052,N_11641);
nand U12948 (N_12948,N_11873,N_11850);
or U12949 (N_12949,N_11721,N_11714);
and U12950 (N_12950,N_11858,N_11802);
nand U12951 (N_12951,N_11495,N_11273);
nand U12952 (N_12952,N_11731,N_11463);
xor U12953 (N_12953,N_11113,N_11666);
xor U12954 (N_12954,N_11602,N_11640);
nor U12955 (N_12955,N_11045,N_11940);
and U12956 (N_12956,N_11323,N_11344);
xor U12957 (N_12957,N_11330,N_11420);
xor U12958 (N_12958,N_11285,N_11705);
xor U12959 (N_12959,N_11134,N_11605);
nand U12960 (N_12960,N_11648,N_11704);
or U12961 (N_12961,N_11361,N_11235);
and U12962 (N_12962,N_11360,N_11165);
or U12963 (N_12963,N_11139,N_11299);
nor U12964 (N_12964,N_11108,N_11500);
nor U12965 (N_12965,N_11695,N_11062);
nand U12966 (N_12966,N_11975,N_11467);
and U12967 (N_12967,N_11142,N_11461);
or U12968 (N_12968,N_11664,N_11585);
nand U12969 (N_12969,N_11214,N_11626);
xor U12970 (N_12970,N_11707,N_11623);
nand U12971 (N_12971,N_11688,N_11534);
and U12972 (N_12972,N_11847,N_11649);
nand U12973 (N_12973,N_11163,N_11973);
nand U12974 (N_12974,N_11333,N_11876);
xnor U12975 (N_12975,N_11916,N_11330);
nor U12976 (N_12976,N_11324,N_11465);
xor U12977 (N_12977,N_11161,N_11592);
and U12978 (N_12978,N_11818,N_11812);
or U12979 (N_12979,N_11439,N_11218);
nand U12980 (N_12980,N_11724,N_11654);
xor U12981 (N_12981,N_11259,N_11548);
and U12982 (N_12982,N_11188,N_11009);
nand U12983 (N_12983,N_11360,N_11050);
and U12984 (N_12984,N_11225,N_11845);
nor U12985 (N_12985,N_11969,N_11961);
xnor U12986 (N_12986,N_11897,N_11237);
xor U12987 (N_12987,N_11964,N_11332);
nor U12988 (N_12988,N_11982,N_11971);
xnor U12989 (N_12989,N_11328,N_11265);
and U12990 (N_12990,N_11921,N_11631);
and U12991 (N_12991,N_11904,N_11745);
xnor U12992 (N_12992,N_11847,N_11226);
nand U12993 (N_12993,N_11977,N_11414);
or U12994 (N_12994,N_11799,N_11546);
nor U12995 (N_12995,N_11964,N_11481);
xor U12996 (N_12996,N_11749,N_11689);
nor U12997 (N_12997,N_11173,N_11068);
nor U12998 (N_12998,N_11467,N_11783);
xnor U12999 (N_12999,N_11425,N_11913);
and U13000 (N_13000,N_12350,N_12416);
and U13001 (N_13001,N_12444,N_12618);
nor U13002 (N_13002,N_12245,N_12334);
and U13003 (N_13003,N_12167,N_12452);
nor U13004 (N_13004,N_12064,N_12472);
and U13005 (N_13005,N_12056,N_12773);
nand U13006 (N_13006,N_12593,N_12552);
and U13007 (N_13007,N_12042,N_12335);
xor U13008 (N_13008,N_12944,N_12413);
and U13009 (N_13009,N_12818,N_12759);
nor U13010 (N_13010,N_12875,N_12088);
and U13011 (N_13011,N_12981,N_12743);
and U13012 (N_13012,N_12059,N_12545);
nor U13013 (N_13013,N_12942,N_12299);
nand U13014 (N_13014,N_12694,N_12664);
and U13015 (N_13015,N_12327,N_12096);
nand U13016 (N_13016,N_12862,N_12763);
xor U13017 (N_13017,N_12557,N_12336);
and U13018 (N_13018,N_12551,N_12524);
or U13019 (N_13019,N_12548,N_12098);
nor U13020 (N_13020,N_12858,N_12440);
nor U13021 (N_13021,N_12279,N_12676);
nor U13022 (N_13022,N_12443,N_12419);
nor U13023 (N_13023,N_12190,N_12163);
or U13024 (N_13024,N_12415,N_12221);
nand U13025 (N_13025,N_12781,N_12595);
and U13026 (N_13026,N_12066,N_12263);
nor U13027 (N_13027,N_12609,N_12680);
nor U13028 (N_13028,N_12248,N_12039);
or U13029 (N_13029,N_12582,N_12038);
or U13030 (N_13030,N_12107,N_12847);
or U13031 (N_13031,N_12909,N_12142);
or U13032 (N_13032,N_12404,N_12037);
nand U13033 (N_13033,N_12176,N_12365);
xor U13034 (N_13034,N_12608,N_12705);
and U13035 (N_13035,N_12501,N_12052);
and U13036 (N_13036,N_12325,N_12271);
xor U13037 (N_13037,N_12172,N_12022);
and U13038 (N_13038,N_12250,N_12396);
or U13039 (N_13039,N_12182,N_12885);
nand U13040 (N_13040,N_12083,N_12624);
and U13041 (N_13041,N_12740,N_12202);
nand U13042 (N_13042,N_12659,N_12171);
nor U13043 (N_13043,N_12127,N_12211);
nand U13044 (N_13044,N_12326,N_12857);
and U13045 (N_13045,N_12550,N_12650);
nand U13046 (N_13046,N_12585,N_12288);
xnor U13047 (N_13047,N_12104,N_12020);
or U13048 (N_13048,N_12733,N_12891);
or U13049 (N_13049,N_12260,N_12222);
and U13050 (N_13050,N_12722,N_12840);
xor U13051 (N_13051,N_12370,N_12215);
nor U13052 (N_13052,N_12067,N_12851);
nand U13053 (N_13053,N_12837,N_12579);
nand U13054 (N_13054,N_12360,N_12724);
nor U13055 (N_13055,N_12156,N_12817);
nand U13056 (N_13056,N_12344,N_12723);
and U13057 (N_13057,N_12374,N_12235);
xnor U13058 (N_13058,N_12927,N_12183);
xnor U13059 (N_13059,N_12797,N_12751);
and U13060 (N_13060,N_12471,N_12206);
and U13061 (N_13061,N_12943,N_12785);
or U13062 (N_13062,N_12478,N_12777);
and U13063 (N_13063,N_12589,N_12109);
nand U13064 (N_13064,N_12441,N_12569);
and U13065 (N_13065,N_12941,N_12381);
xnor U13066 (N_13066,N_12813,N_12790);
xor U13067 (N_13067,N_12398,N_12760);
xor U13068 (N_13068,N_12873,N_12418);
xnor U13069 (N_13069,N_12658,N_12553);
and U13070 (N_13070,N_12446,N_12805);
xnor U13071 (N_13071,N_12735,N_12558);
nand U13072 (N_13072,N_12725,N_12379);
nor U13073 (N_13073,N_12554,N_12488);
or U13074 (N_13074,N_12389,N_12364);
and U13075 (N_13075,N_12195,N_12679);
nor U13076 (N_13076,N_12462,N_12259);
nand U13077 (N_13077,N_12314,N_12485);
or U13078 (N_13078,N_12361,N_12072);
and U13079 (N_13079,N_12187,N_12428);
nor U13080 (N_13080,N_12584,N_12613);
nor U13081 (N_13081,N_12809,N_12426);
and U13082 (N_13082,N_12542,N_12796);
nand U13083 (N_13083,N_12191,N_12863);
and U13084 (N_13084,N_12528,N_12870);
nand U13085 (N_13085,N_12332,N_12291);
nand U13086 (N_13086,N_12228,N_12673);
nor U13087 (N_13087,N_12503,N_12125);
nor U13088 (N_13088,N_12266,N_12427);
xor U13089 (N_13089,N_12216,N_12217);
xor U13090 (N_13090,N_12368,N_12371);
xor U13091 (N_13091,N_12924,N_12457);
nor U13092 (N_13092,N_12560,N_12556);
and U13093 (N_13093,N_12755,N_12407);
xnor U13094 (N_13094,N_12303,N_12516);
nand U13095 (N_13095,N_12463,N_12695);
or U13096 (N_13096,N_12752,N_12866);
or U13097 (N_13097,N_12736,N_12848);
nand U13098 (N_13098,N_12963,N_12349);
xnor U13099 (N_13099,N_12147,N_12612);
xnor U13100 (N_13100,N_12641,N_12910);
nand U13101 (N_13101,N_12160,N_12318);
or U13102 (N_13102,N_12704,N_12054);
or U13103 (N_13103,N_12449,N_12240);
nand U13104 (N_13104,N_12561,N_12274);
nor U13105 (N_13105,N_12009,N_12521);
nand U13106 (N_13106,N_12223,N_12285);
xor U13107 (N_13107,N_12513,N_12714);
nand U13108 (N_13108,N_12654,N_12635);
or U13109 (N_13109,N_12587,N_12682);
nor U13110 (N_13110,N_12091,N_12778);
and U13111 (N_13111,N_12661,N_12949);
and U13112 (N_13112,N_12945,N_12563);
and U13113 (N_13113,N_12950,N_12881);
nor U13114 (N_13114,N_12780,N_12117);
or U13115 (N_13115,N_12712,N_12055);
nand U13116 (N_13116,N_12019,N_12464);
nand U13117 (N_13117,N_12955,N_12715);
nor U13118 (N_13118,N_12006,N_12282);
nand U13119 (N_13119,N_12816,N_12166);
nand U13120 (N_13120,N_12114,N_12395);
or U13121 (N_13121,N_12456,N_12717);
xor U13122 (N_13122,N_12244,N_12935);
and U13123 (N_13123,N_12047,N_12926);
or U13124 (N_13124,N_12794,N_12912);
xnor U13125 (N_13125,N_12859,N_12205);
or U13126 (N_13126,N_12425,N_12028);
and U13127 (N_13127,N_12157,N_12132);
and U13128 (N_13128,N_12414,N_12693);
nor U13129 (N_13129,N_12776,N_12667);
nor U13130 (N_13130,N_12701,N_12339);
xnor U13131 (N_13131,N_12196,N_12233);
nand U13132 (N_13132,N_12402,N_12341);
xnor U13133 (N_13133,N_12911,N_12508);
or U13134 (N_13134,N_12892,N_12810);
xnor U13135 (N_13135,N_12957,N_12515);
nor U13136 (N_13136,N_12744,N_12313);
and U13137 (N_13137,N_12698,N_12625);
or U13138 (N_13138,N_12430,N_12934);
xor U13139 (N_13139,N_12119,N_12372);
nor U13140 (N_13140,N_12804,N_12201);
xnor U13141 (N_13141,N_12305,N_12583);
xor U13142 (N_13142,N_12353,N_12691);
xnor U13143 (N_13143,N_12198,N_12474);
nor U13144 (N_13144,N_12110,N_12380);
nor U13145 (N_13145,N_12639,N_12903);
and U13146 (N_13146,N_12771,N_12675);
nor U13147 (N_13147,N_12026,N_12242);
nor U13148 (N_13148,N_12540,N_12126);
nor U13149 (N_13149,N_12852,N_12207);
or U13150 (N_13150,N_12879,N_12237);
xor U13151 (N_13151,N_12424,N_12145);
or U13152 (N_13152,N_12665,N_12895);
or U13153 (N_13153,N_12897,N_12779);
and U13154 (N_13154,N_12657,N_12227);
and U13155 (N_13155,N_12541,N_12627);
or U13156 (N_13156,N_12189,N_12036);
and U13157 (N_13157,N_12685,N_12293);
xor U13158 (N_13158,N_12985,N_12670);
xnor U13159 (N_13159,N_12050,N_12252);
nor U13160 (N_13160,N_12023,N_12989);
nor U13161 (N_13161,N_12732,N_12533);
and U13162 (N_13162,N_12792,N_12017);
nor U13163 (N_13163,N_12502,N_12748);
and U13164 (N_13164,N_12065,N_12005);
and U13165 (N_13165,N_12388,N_12506);
and U13166 (N_13166,N_12130,N_12011);
and U13167 (N_13167,N_12729,N_12007);
and U13168 (N_13168,N_12004,N_12842);
or U13169 (N_13169,N_12092,N_12382);
and U13170 (N_13170,N_12438,N_12113);
or U13171 (N_13171,N_12041,N_12008);
or U13172 (N_13172,N_12720,N_12787);
or U13173 (N_13173,N_12466,N_12476);
nor U13174 (N_13174,N_12409,N_12820);
and U13175 (N_13175,N_12697,N_12309);
and U13176 (N_13176,N_12486,N_12304);
xor U13177 (N_13177,N_12835,N_12494);
xnor U13178 (N_13178,N_12431,N_12180);
or U13179 (N_13179,N_12174,N_12151);
or U13180 (N_13180,N_12284,N_12839);
nor U13181 (N_13181,N_12750,N_12470);
nor U13182 (N_13182,N_12432,N_12164);
or U13183 (N_13183,N_12278,N_12784);
and U13184 (N_13184,N_12965,N_12849);
xnor U13185 (N_13185,N_12721,N_12080);
or U13186 (N_13186,N_12029,N_12032);
xor U13187 (N_13187,N_12543,N_12655);
nand U13188 (N_13188,N_12060,N_12562);
xor U13189 (N_13189,N_12573,N_12971);
or U13190 (N_13190,N_12373,N_12277);
or U13191 (N_13191,N_12451,N_12692);
nor U13192 (N_13192,N_12669,N_12102);
and U13193 (N_13193,N_12865,N_12605);
or U13194 (N_13194,N_12660,N_12033);
xor U13195 (N_13195,N_12577,N_12544);
nor U13196 (N_13196,N_12684,N_12359);
nand U13197 (N_13197,N_12101,N_12638);
nor U13198 (N_13198,N_12391,N_12437);
and U13199 (N_13199,N_12491,N_12181);
nor U13200 (N_13200,N_12337,N_12024);
nand U13201 (N_13201,N_12719,N_12118);
xor U13202 (N_13202,N_12321,N_12129);
or U13203 (N_13203,N_12194,N_12296);
or U13204 (N_13204,N_12246,N_12993);
nor U13205 (N_13205,N_12013,N_12429);
nand U13206 (N_13206,N_12994,N_12890);
and U13207 (N_13207,N_12500,N_12900);
and U13208 (N_13208,N_12168,N_12634);
xnor U13209 (N_13209,N_12392,N_12153);
nand U13210 (N_13210,N_12568,N_12856);
xor U13211 (N_13211,N_12917,N_12915);
and U13212 (N_13212,N_12534,N_12018);
nor U13213 (N_13213,N_12340,N_12089);
nor U13214 (N_13214,N_12297,N_12643);
nand U13215 (N_13215,N_12086,N_12907);
or U13216 (N_13216,N_12475,N_12970);
xor U13217 (N_13217,N_12893,N_12154);
nand U13218 (N_13218,N_12651,N_12861);
nor U13219 (N_13219,N_12075,N_12880);
and U13220 (N_13220,N_12827,N_12707);
and U13221 (N_13221,N_12826,N_12281);
nor U13222 (N_13222,N_12140,N_12306);
nor U13223 (N_13223,N_12467,N_12308);
or U13224 (N_13224,N_12203,N_12058);
xnor U13225 (N_13225,N_12090,N_12869);
or U13226 (N_13226,N_12830,N_12329);
xnor U13227 (N_13227,N_12410,N_12683);
nand U13228 (N_13228,N_12517,N_12481);
nor U13229 (N_13229,N_12403,N_12238);
or U13230 (N_13230,N_12115,N_12256);
nor U13231 (N_13231,N_12433,N_12588);
nor U13232 (N_13232,N_12711,N_12769);
xnor U13233 (N_13233,N_12400,N_12298);
xor U13234 (N_13234,N_12422,N_12224);
or U13235 (N_13235,N_12034,N_12095);
nand U13236 (N_13236,N_12112,N_12954);
nand U13237 (N_13237,N_12850,N_12681);
nor U13238 (N_13238,N_12027,N_12765);
nor U13239 (N_13239,N_12600,N_12594);
xnor U13240 (N_13240,N_12001,N_12489);
or U13241 (N_13241,N_12872,N_12646);
xor U13242 (N_13242,N_12764,N_12961);
nand U13243 (N_13243,N_12962,N_12333);
xor U13244 (N_13244,N_12601,N_12864);
xnor U13245 (N_13245,N_12057,N_12363);
xor U13246 (N_13246,N_12774,N_12982);
xor U13247 (N_13247,N_12469,N_12315);
or U13248 (N_13248,N_12300,N_12808);
nand U13249 (N_13249,N_12031,N_12746);
nor U13250 (N_13250,N_12385,N_12135);
and U13251 (N_13251,N_12131,N_12783);
nor U13252 (N_13252,N_12214,N_12572);
nand U13253 (N_13253,N_12974,N_12843);
nor U13254 (N_13254,N_12726,N_12272);
xor U13255 (N_13255,N_12251,N_12570);
and U13256 (N_13256,N_12731,N_12301);
xnor U13257 (N_13257,N_12567,N_12914);
nor U13258 (N_13258,N_12571,N_12951);
xor U13259 (N_13259,N_12290,N_12234);
and U13260 (N_13260,N_12111,N_12619);
nor U13261 (N_13261,N_12716,N_12555);
and U13262 (N_13262,N_12519,N_12267);
nand U13263 (N_13263,N_12597,N_12143);
or U13264 (N_13264,N_12292,N_12012);
or U13265 (N_13265,N_12546,N_12768);
nor U13266 (N_13266,N_12980,N_12591);
xnor U13267 (N_13267,N_12045,N_12756);
or U13268 (N_13268,N_12966,N_12596);
and U13269 (N_13269,N_12832,N_12103);
and U13270 (N_13270,N_12280,N_12504);
nor U13271 (N_13271,N_12040,N_12801);
and U13272 (N_13272,N_12108,N_12718);
nor U13273 (N_13273,N_12420,N_12121);
nor U13274 (N_13274,N_12604,N_12386);
nand U13275 (N_13275,N_12188,N_12806);
and U13276 (N_13276,N_12703,N_12249);
xnor U13277 (N_13277,N_12868,N_12645);
and U13278 (N_13278,N_12621,N_12152);
or U13279 (N_13279,N_12753,N_12853);
nor U13280 (N_13280,N_12078,N_12610);
and U13281 (N_13281,N_12666,N_12208);
xnor U13282 (N_13282,N_12003,N_12071);
or U13283 (N_13283,N_12048,N_12497);
nand U13284 (N_13284,N_12068,N_12509);
or U13285 (N_13285,N_12925,N_12647);
and U13286 (N_13286,N_12406,N_12123);
xor U13287 (N_13287,N_12939,N_12254);
nand U13288 (N_13288,N_12576,N_12648);
xor U13289 (N_13289,N_12498,N_12928);
nand U13290 (N_13290,N_12439,N_12387);
or U13291 (N_13291,N_12877,N_12405);
nand U13292 (N_13292,N_12799,N_12069);
and U13293 (N_13293,N_12087,N_12739);
or U13294 (N_13294,N_12186,N_12946);
nor U13295 (N_13295,N_12975,N_12518);
xor U13296 (N_13296,N_12480,N_12459);
nor U13297 (N_13297,N_12043,N_12902);
nand U13298 (N_13298,N_12932,N_12884);
nand U13299 (N_13299,N_12197,N_12616);
nand U13300 (N_13300,N_12894,N_12770);
and U13301 (N_13301,N_12447,N_12209);
nand U13302 (N_13302,N_12757,N_12461);
xor U13303 (N_13303,N_12077,N_12922);
and U13304 (N_13304,N_12218,N_12199);
and U13305 (N_13305,N_12883,N_12986);
or U13306 (N_13306,N_12000,N_12815);
or U13307 (N_13307,N_12964,N_12825);
and U13308 (N_13308,N_12231,N_12139);
or U13309 (N_13309,N_12690,N_12793);
nor U13310 (N_13310,N_12434,N_12331);
nor U13311 (N_13311,N_12261,N_12953);
or U13312 (N_13312,N_12987,N_12495);
nand U13313 (N_13313,N_12882,N_12824);
and U13314 (N_13314,N_12905,N_12747);
nor U13315 (N_13315,N_12316,N_12737);
nor U13316 (N_13316,N_12124,N_12754);
nor U13317 (N_13317,N_12795,N_12225);
nor U13318 (N_13318,N_12378,N_12184);
and U13319 (N_13319,N_12220,N_12836);
and U13320 (N_13320,N_12514,N_12150);
xnor U13321 (N_13321,N_12454,N_12623);
xnor U13322 (N_13322,N_12526,N_12257);
or U13323 (N_13323,N_12106,N_12615);
and U13324 (N_13324,N_12273,N_12878);
and U13325 (N_13325,N_12630,N_12937);
nor U13326 (N_13326,N_12766,N_12844);
and U13327 (N_13327,N_12607,N_12901);
or U13328 (N_13328,N_12745,N_12663);
nand U13329 (N_13329,N_12838,N_12161);
or U13330 (N_13330,N_12133,N_12995);
or U13331 (N_13331,N_12969,N_12535);
or U13332 (N_13332,N_12959,N_12136);
or U13333 (N_13333,N_12979,N_12445);
or U13334 (N_13334,N_12940,N_12144);
xor U13335 (N_13335,N_12738,N_12074);
xnor U13336 (N_13336,N_12800,N_12049);
or U13337 (N_13337,N_12499,N_12734);
and U13338 (N_13338,N_12458,N_12384);
or U13339 (N_13339,N_12061,N_12831);
nand U13340 (N_13340,N_12210,N_12232);
or U13341 (N_13341,N_12626,N_12421);
or U13342 (N_13342,N_12148,N_12527);
nor U13343 (N_13343,N_12204,N_12175);
xnor U13344 (N_13344,N_12644,N_12496);
or U13345 (N_13345,N_12581,N_12170);
or U13346 (N_13346,N_12958,N_12984);
nor U13347 (N_13347,N_12319,N_12330);
nand U13348 (N_13348,N_12898,N_12442);
or U13349 (N_13349,N_12046,N_12302);
nand U13350 (N_13350,N_12348,N_12919);
nor U13351 (N_13351,N_12983,N_12845);
nor U13352 (N_13352,N_12212,N_12397);
xor U13353 (N_13353,N_12473,N_12312);
nor U13354 (N_13354,N_12178,N_12070);
xnor U13355 (N_13355,N_12484,N_12908);
nand U13356 (N_13356,N_12632,N_12617);
or U13357 (N_13357,N_12435,N_12507);
xor U13358 (N_13358,N_12120,N_12487);
nand U13359 (N_13359,N_12097,N_12702);
nor U13360 (N_13360,N_12631,N_12821);
nor U13361 (N_13361,N_12357,N_12833);
or U13362 (N_13362,N_12479,N_12358);
and U13363 (N_13363,N_12586,N_12999);
or U13364 (N_13364,N_12798,N_12493);
xor U13365 (N_13365,N_12633,N_12169);
xor U13366 (N_13366,N_12992,N_12492);
xnor U13367 (N_13367,N_12906,N_12532);
nand U13368 (N_13368,N_12149,N_12352);
and U13369 (N_13369,N_12412,N_12417);
and U13370 (N_13370,N_12367,N_12294);
or U13371 (N_13371,N_12997,N_12085);
or U13372 (N_13372,N_12592,N_12559);
and U13373 (N_13373,N_12081,N_12255);
xor U13374 (N_13374,N_12938,N_12749);
nor U13375 (N_13375,N_12867,N_12122);
nor U13376 (N_13376,N_12700,N_12383);
nor U13377 (N_13377,N_12295,N_12002);
and U13378 (N_13378,N_12342,N_12423);
nand U13379 (N_13379,N_12977,N_12791);
nand U13380 (N_13380,N_12956,N_12611);
xor U13381 (N_13381,N_12823,N_12269);
and U13382 (N_13382,N_12276,N_12450);
and U13383 (N_13383,N_12923,N_12968);
nand U13384 (N_13384,N_12162,N_12159);
xor U13385 (N_13385,N_12991,N_12270);
and U13386 (N_13386,N_12323,N_12286);
and U13387 (N_13387,N_12511,N_12345);
nor U13388 (N_13388,N_12742,N_12530);
xor U13389 (N_13389,N_12674,N_12351);
xnor U13390 (N_13390,N_12689,N_12887);
nand U13391 (N_13391,N_12510,N_12598);
and U13392 (N_13392,N_12931,N_12200);
or U13393 (N_13393,N_12141,N_12229);
nand U13394 (N_13394,N_12084,N_12165);
or U13395 (N_13395,N_12628,N_12566);
and U13396 (N_13396,N_12035,N_12761);
xnor U13397 (N_13397,N_12930,N_12854);
or U13398 (N_13398,N_12536,N_12710);
or U13399 (N_13399,N_12727,N_12565);
nor U13400 (N_13400,N_12236,N_12094);
xor U13401 (N_13401,N_12637,N_12053);
and U13402 (N_13402,N_12772,N_12063);
nand U13403 (N_13403,N_12453,N_12976);
and U13404 (N_13404,N_12874,N_12708);
nand U13405 (N_13405,N_12137,N_12247);
and U13406 (N_13406,N_12775,N_12512);
nand U13407 (N_13407,N_12529,N_12614);
nor U13408 (N_13408,N_12936,N_12622);
nand U13409 (N_13409,N_12899,N_12603);
xnor U13410 (N_13410,N_12539,N_12505);
nor U13411 (N_13411,N_12812,N_12226);
xor U13412 (N_13412,N_12871,N_12030);
or U13413 (N_13413,N_12656,N_12814);
xor U13414 (N_13414,N_12062,N_12490);
nand U13415 (N_13415,N_12310,N_12460);
or U13416 (N_13416,N_12362,N_12636);
nor U13417 (N_13417,N_12730,N_12354);
nor U13418 (N_13418,N_12967,N_12128);
and U13419 (N_13419,N_12275,N_12411);
xor U13420 (N_13420,N_12401,N_12146);
and U13421 (N_13421,N_12687,N_12929);
or U13422 (N_13422,N_12328,N_12390);
and U13423 (N_13423,N_12253,N_12741);
xor U13424 (N_13424,N_12876,N_12523);
or U13425 (N_13425,N_12662,N_12173);
or U13426 (N_13426,N_12549,N_12921);
or U13427 (N_13427,N_12155,N_12265);
or U13428 (N_13428,N_12377,N_12642);
xor U13429 (N_13429,N_12758,N_12347);
nand U13430 (N_13430,N_12978,N_12652);
and U13431 (N_13431,N_12520,N_12021);
or U13432 (N_13432,N_12564,N_12789);
and U13433 (N_13433,N_12317,N_12653);
and U13434 (N_13434,N_12366,N_12483);
xor U13435 (N_13435,N_12828,N_12016);
nor U13436 (N_13436,N_12394,N_12258);
nor U13437 (N_13437,N_12972,N_12044);
xnor U13438 (N_13438,N_12099,N_12846);
nand U13439 (N_13439,N_12010,N_12262);
or U13440 (N_13440,N_12307,N_12241);
nor U13441 (N_13441,N_12547,N_12677);
and U13442 (N_13442,N_12213,N_12960);
xnor U13443 (N_13443,N_12802,N_12620);
nand U13444 (N_13444,N_12916,N_12230);
xor U13445 (N_13445,N_12822,N_12522);
xnor U13446 (N_13446,N_12538,N_12192);
xnor U13447 (N_13447,N_12918,N_12688);
nand U13448 (N_13448,N_12287,N_12436);
nand U13449 (N_13449,N_12575,N_12578);
xnor U13450 (N_13450,N_12179,N_12606);
and U13451 (N_13451,N_12803,N_12855);
nand U13452 (N_13452,N_12324,N_12116);
nand U13453 (N_13453,N_12079,N_12015);
and U13454 (N_13454,N_12185,N_12819);
nor U13455 (N_13455,N_12376,N_12356);
or U13456 (N_13456,N_12537,N_12580);
xnor U13457 (N_13457,N_12686,N_12408);
nand U13458 (N_13458,N_12788,N_12343);
or U13459 (N_13459,N_12640,N_12629);
or U13460 (N_13460,N_12531,N_12889);
and U13461 (N_13461,N_12602,N_12355);
and U13462 (N_13462,N_12477,N_12346);
or U13463 (N_13463,N_12888,N_12590);
nor U13464 (N_13464,N_12990,N_12886);
nor U13465 (N_13465,N_12482,N_12375);
nor U13466 (N_13466,N_12672,N_12913);
nor U13467 (N_13467,N_12082,N_12713);
or U13468 (N_13468,N_12311,N_12134);
xor U13469 (N_13469,N_12025,N_12834);
and U13470 (N_13470,N_12283,N_12996);
nor U13471 (N_13471,N_12138,N_12786);
nand U13472 (N_13472,N_12952,N_12574);
xnor U13473 (N_13473,N_12807,N_12264);
xor U13474 (N_13474,N_12338,N_12322);
or U13475 (N_13475,N_12320,N_12988);
xor U13476 (N_13476,N_12105,N_12948);
xor U13477 (N_13477,N_12289,N_12369);
nand U13478 (N_13478,N_12998,N_12393);
nand U13479 (N_13479,N_12671,N_12239);
xor U13480 (N_13480,N_12696,N_12668);
or U13481 (N_13481,N_12399,N_12649);
and U13482 (N_13482,N_12599,N_12767);
and U13483 (N_13483,N_12811,N_12076);
xor U13484 (N_13484,N_12100,N_12860);
nor U13485 (N_13485,N_12678,N_12455);
xor U13486 (N_13486,N_12973,N_12947);
nor U13487 (N_13487,N_12782,N_12468);
xor U13488 (N_13488,N_12177,N_12073);
or U13489 (N_13489,N_12525,N_12933);
and U13490 (N_13490,N_12896,N_12158);
and U13491 (N_13491,N_12051,N_12841);
xor U13492 (N_13492,N_12243,N_12762);
or U13493 (N_13493,N_12904,N_12706);
or U13494 (N_13494,N_12219,N_12014);
nand U13495 (N_13495,N_12448,N_12268);
nand U13496 (N_13496,N_12699,N_12829);
or U13497 (N_13497,N_12465,N_12709);
xnor U13498 (N_13498,N_12193,N_12728);
or U13499 (N_13499,N_12093,N_12920);
and U13500 (N_13500,N_12413,N_12639);
nand U13501 (N_13501,N_12292,N_12321);
xnor U13502 (N_13502,N_12932,N_12610);
nand U13503 (N_13503,N_12391,N_12351);
nor U13504 (N_13504,N_12295,N_12937);
and U13505 (N_13505,N_12509,N_12911);
xnor U13506 (N_13506,N_12754,N_12803);
and U13507 (N_13507,N_12048,N_12933);
xor U13508 (N_13508,N_12407,N_12183);
or U13509 (N_13509,N_12862,N_12778);
or U13510 (N_13510,N_12169,N_12861);
or U13511 (N_13511,N_12183,N_12693);
and U13512 (N_13512,N_12787,N_12970);
or U13513 (N_13513,N_12662,N_12956);
xnor U13514 (N_13514,N_12378,N_12916);
and U13515 (N_13515,N_12047,N_12032);
nor U13516 (N_13516,N_12645,N_12149);
and U13517 (N_13517,N_12506,N_12356);
nor U13518 (N_13518,N_12566,N_12847);
nor U13519 (N_13519,N_12369,N_12619);
and U13520 (N_13520,N_12204,N_12631);
or U13521 (N_13521,N_12813,N_12556);
nor U13522 (N_13522,N_12069,N_12260);
nor U13523 (N_13523,N_12193,N_12839);
xnor U13524 (N_13524,N_12268,N_12293);
xnor U13525 (N_13525,N_12070,N_12760);
xnor U13526 (N_13526,N_12371,N_12310);
and U13527 (N_13527,N_12772,N_12009);
nor U13528 (N_13528,N_12495,N_12074);
or U13529 (N_13529,N_12808,N_12386);
or U13530 (N_13530,N_12049,N_12869);
and U13531 (N_13531,N_12937,N_12906);
or U13532 (N_13532,N_12672,N_12780);
nor U13533 (N_13533,N_12652,N_12458);
xor U13534 (N_13534,N_12762,N_12324);
xor U13535 (N_13535,N_12734,N_12259);
or U13536 (N_13536,N_12265,N_12867);
nand U13537 (N_13537,N_12911,N_12128);
and U13538 (N_13538,N_12050,N_12556);
and U13539 (N_13539,N_12074,N_12124);
nor U13540 (N_13540,N_12362,N_12807);
nand U13541 (N_13541,N_12385,N_12144);
or U13542 (N_13542,N_12768,N_12599);
nor U13543 (N_13543,N_12327,N_12291);
or U13544 (N_13544,N_12632,N_12810);
nor U13545 (N_13545,N_12046,N_12789);
nand U13546 (N_13546,N_12497,N_12475);
and U13547 (N_13547,N_12966,N_12704);
nor U13548 (N_13548,N_12016,N_12855);
xor U13549 (N_13549,N_12901,N_12851);
nand U13550 (N_13550,N_12812,N_12647);
xor U13551 (N_13551,N_12768,N_12830);
or U13552 (N_13552,N_12468,N_12194);
xnor U13553 (N_13553,N_12849,N_12122);
and U13554 (N_13554,N_12945,N_12141);
xnor U13555 (N_13555,N_12876,N_12009);
nand U13556 (N_13556,N_12265,N_12460);
nand U13557 (N_13557,N_12799,N_12026);
and U13558 (N_13558,N_12085,N_12483);
and U13559 (N_13559,N_12021,N_12402);
nor U13560 (N_13560,N_12959,N_12257);
and U13561 (N_13561,N_12365,N_12481);
nand U13562 (N_13562,N_12454,N_12442);
nand U13563 (N_13563,N_12714,N_12677);
and U13564 (N_13564,N_12071,N_12606);
xor U13565 (N_13565,N_12924,N_12680);
nor U13566 (N_13566,N_12080,N_12347);
and U13567 (N_13567,N_12361,N_12265);
xnor U13568 (N_13568,N_12633,N_12340);
nand U13569 (N_13569,N_12913,N_12926);
xor U13570 (N_13570,N_12793,N_12444);
and U13571 (N_13571,N_12267,N_12539);
nor U13572 (N_13572,N_12764,N_12123);
nand U13573 (N_13573,N_12642,N_12152);
nand U13574 (N_13574,N_12435,N_12424);
or U13575 (N_13575,N_12204,N_12438);
or U13576 (N_13576,N_12876,N_12530);
nor U13577 (N_13577,N_12262,N_12507);
or U13578 (N_13578,N_12348,N_12838);
or U13579 (N_13579,N_12424,N_12558);
xor U13580 (N_13580,N_12527,N_12567);
or U13581 (N_13581,N_12977,N_12297);
nand U13582 (N_13582,N_12620,N_12322);
nor U13583 (N_13583,N_12820,N_12742);
nand U13584 (N_13584,N_12512,N_12517);
xor U13585 (N_13585,N_12294,N_12097);
nor U13586 (N_13586,N_12216,N_12063);
and U13587 (N_13587,N_12259,N_12793);
xor U13588 (N_13588,N_12273,N_12760);
and U13589 (N_13589,N_12963,N_12731);
or U13590 (N_13590,N_12132,N_12707);
nand U13591 (N_13591,N_12545,N_12557);
nand U13592 (N_13592,N_12458,N_12683);
and U13593 (N_13593,N_12518,N_12680);
or U13594 (N_13594,N_12034,N_12027);
nor U13595 (N_13595,N_12608,N_12817);
or U13596 (N_13596,N_12682,N_12806);
nor U13597 (N_13597,N_12775,N_12807);
or U13598 (N_13598,N_12629,N_12658);
or U13599 (N_13599,N_12930,N_12460);
or U13600 (N_13600,N_12933,N_12790);
and U13601 (N_13601,N_12032,N_12283);
and U13602 (N_13602,N_12516,N_12296);
or U13603 (N_13603,N_12802,N_12302);
nand U13604 (N_13604,N_12645,N_12486);
nand U13605 (N_13605,N_12311,N_12230);
nor U13606 (N_13606,N_12464,N_12148);
or U13607 (N_13607,N_12026,N_12973);
xor U13608 (N_13608,N_12545,N_12797);
xnor U13609 (N_13609,N_12091,N_12879);
nand U13610 (N_13610,N_12705,N_12252);
nor U13611 (N_13611,N_12005,N_12739);
or U13612 (N_13612,N_12123,N_12339);
and U13613 (N_13613,N_12717,N_12804);
nor U13614 (N_13614,N_12860,N_12696);
or U13615 (N_13615,N_12075,N_12567);
xor U13616 (N_13616,N_12728,N_12228);
or U13617 (N_13617,N_12603,N_12564);
or U13618 (N_13618,N_12933,N_12144);
nand U13619 (N_13619,N_12069,N_12473);
nor U13620 (N_13620,N_12322,N_12385);
and U13621 (N_13621,N_12264,N_12099);
nand U13622 (N_13622,N_12436,N_12954);
and U13623 (N_13623,N_12379,N_12333);
or U13624 (N_13624,N_12869,N_12453);
or U13625 (N_13625,N_12941,N_12042);
xor U13626 (N_13626,N_12618,N_12002);
or U13627 (N_13627,N_12253,N_12094);
xor U13628 (N_13628,N_12166,N_12023);
or U13629 (N_13629,N_12802,N_12002);
nor U13630 (N_13630,N_12167,N_12073);
and U13631 (N_13631,N_12178,N_12854);
or U13632 (N_13632,N_12664,N_12921);
xor U13633 (N_13633,N_12203,N_12436);
or U13634 (N_13634,N_12263,N_12564);
nand U13635 (N_13635,N_12286,N_12890);
xor U13636 (N_13636,N_12039,N_12056);
and U13637 (N_13637,N_12865,N_12819);
xor U13638 (N_13638,N_12772,N_12909);
nor U13639 (N_13639,N_12238,N_12993);
nand U13640 (N_13640,N_12262,N_12456);
and U13641 (N_13641,N_12039,N_12424);
nand U13642 (N_13642,N_12804,N_12952);
nor U13643 (N_13643,N_12364,N_12516);
xnor U13644 (N_13644,N_12141,N_12918);
or U13645 (N_13645,N_12002,N_12243);
nor U13646 (N_13646,N_12192,N_12775);
nand U13647 (N_13647,N_12681,N_12236);
nor U13648 (N_13648,N_12610,N_12008);
and U13649 (N_13649,N_12217,N_12938);
nand U13650 (N_13650,N_12052,N_12546);
nor U13651 (N_13651,N_12143,N_12178);
nor U13652 (N_13652,N_12393,N_12481);
nand U13653 (N_13653,N_12832,N_12817);
or U13654 (N_13654,N_12540,N_12515);
and U13655 (N_13655,N_12444,N_12300);
nor U13656 (N_13656,N_12273,N_12588);
nand U13657 (N_13657,N_12119,N_12753);
nor U13658 (N_13658,N_12126,N_12627);
xnor U13659 (N_13659,N_12441,N_12030);
nand U13660 (N_13660,N_12948,N_12473);
nor U13661 (N_13661,N_12776,N_12350);
and U13662 (N_13662,N_12735,N_12631);
or U13663 (N_13663,N_12821,N_12045);
and U13664 (N_13664,N_12889,N_12381);
xnor U13665 (N_13665,N_12124,N_12601);
xnor U13666 (N_13666,N_12466,N_12904);
nand U13667 (N_13667,N_12499,N_12163);
and U13668 (N_13668,N_12714,N_12109);
and U13669 (N_13669,N_12356,N_12385);
or U13670 (N_13670,N_12244,N_12459);
xor U13671 (N_13671,N_12970,N_12116);
nand U13672 (N_13672,N_12000,N_12640);
nand U13673 (N_13673,N_12650,N_12854);
nand U13674 (N_13674,N_12858,N_12803);
and U13675 (N_13675,N_12863,N_12035);
or U13676 (N_13676,N_12868,N_12968);
nor U13677 (N_13677,N_12000,N_12141);
nand U13678 (N_13678,N_12120,N_12126);
or U13679 (N_13679,N_12707,N_12769);
nor U13680 (N_13680,N_12122,N_12125);
and U13681 (N_13681,N_12321,N_12682);
or U13682 (N_13682,N_12303,N_12163);
nand U13683 (N_13683,N_12267,N_12091);
and U13684 (N_13684,N_12293,N_12748);
nand U13685 (N_13685,N_12319,N_12884);
and U13686 (N_13686,N_12314,N_12299);
nor U13687 (N_13687,N_12096,N_12177);
and U13688 (N_13688,N_12691,N_12137);
or U13689 (N_13689,N_12505,N_12570);
nand U13690 (N_13690,N_12283,N_12828);
nand U13691 (N_13691,N_12527,N_12485);
and U13692 (N_13692,N_12153,N_12442);
or U13693 (N_13693,N_12662,N_12712);
and U13694 (N_13694,N_12152,N_12850);
and U13695 (N_13695,N_12811,N_12335);
xnor U13696 (N_13696,N_12345,N_12127);
and U13697 (N_13697,N_12770,N_12496);
and U13698 (N_13698,N_12963,N_12519);
and U13699 (N_13699,N_12433,N_12229);
xnor U13700 (N_13700,N_12016,N_12681);
xnor U13701 (N_13701,N_12080,N_12172);
xnor U13702 (N_13702,N_12714,N_12413);
xnor U13703 (N_13703,N_12453,N_12516);
nor U13704 (N_13704,N_12308,N_12337);
nor U13705 (N_13705,N_12102,N_12167);
nand U13706 (N_13706,N_12099,N_12403);
xnor U13707 (N_13707,N_12022,N_12754);
and U13708 (N_13708,N_12733,N_12910);
nor U13709 (N_13709,N_12948,N_12447);
nand U13710 (N_13710,N_12463,N_12218);
nand U13711 (N_13711,N_12506,N_12750);
nor U13712 (N_13712,N_12613,N_12390);
nor U13713 (N_13713,N_12613,N_12432);
xor U13714 (N_13714,N_12989,N_12770);
and U13715 (N_13715,N_12992,N_12013);
or U13716 (N_13716,N_12673,N_12202);
and U13717 (N_13717,N_12936,N_12387);
or U13718 (N_13718,N_12082,N_12357);
and U13719 (N_13719,N_12803,N_12149);
or U13720 (N_13720,N_12068,N_12997);
xor U13721 (N_13721,N_12574,N_12028);
or U13722 (N_13722,N_12062,N_12863);
or U13723 (N_13723,N_12213,N_12796);
xor U13724 (N_13724,N_12424,N_12738);
nor U13725 (N_13725,N_12361,N_12116);
and U13726 (N_13726,N_12764,N_12794);
and U13727 (N_13727,N_12310,N_12453);
or U13728 (N_13728,N_12736,N_12546);
xnor U13729 (N_13729,N_12830,N_12301);
and U13730 (N_13730,N_12039,N_12650);
nand U13731 (N_13731,N_12025,N_12388);
and U13732 (N_13732,N_12302,N_12134);
xor U13733 (N_13733,N_12414,N_12797);
or U13734 (N_13734,N_12268,N_12747);
nand U13735 (N_13735,N_12229,N_12354);
or U13736 (N_13736,N_12636,N_12399);
or U13737 (N_13737,N_12035,N_12507);
xnor U13738 (N_13738,N_12617,N_12081);
nor U13739 (N_13739,N_12634,N_12626);
and U13740 (N_13740,N_12746,N_12973);
and U13741 (N_13741,N_12666,N_12373);
or U13742 (N_13742,N_12344,N_12946);
or U13743 (N_13743,N_12627,N_12870);
nand U13744 (N_13744,N_12331,N_12516);
and U13745 (N_13745,N_12184,N_12716);
xor U13746 (N_13746,N_12007,N_12986);
xnor U13747 (N_13747,N_12199,N_12072);
and U13748 (N_13748,N_12691,N_12132);
and U13749 (N_13749,N_12924,N_12066);
xor U13750 (N_13750,N_12351,N_12789);
nand U13751 (N_13751,N_12760,N_12117);
nand U13752 (N_13752,N_12293,N_12439);
nor U13753 (N_13753,N_12857,N_12361);
xnor U13754 (N_13754,N_12870,N_12656);
xnor U13755 (N_13755,N_12634,N_12541);
nor U13756 (N_13756,N_12087,N_12209);
or U13757 (N_13757,N_12021,N_12685);
xor U13758 (N_13758,N_12441,N_12476);
xor U13759 (N_13759,N_12317,N_12163);
nand U13760 (N_13760,N_12030,N_12506);
nand U13761 (N_13761,N_12470,N_12479);
and U13762 (N_13762,N_12852,N_12540);
or U13763 (N_13763,N_12189,N_12592);
nand U13764 (N_13764,N_12606,N_12747);
nand U13765 (N_13765,N_12785,N_12889);
nor U13766 (N_13766,N_12920,N_12343);
nor U13767 (N_13767,N_12934,N_12062);
or U13768 (N_13768,N_12205,N_12583);
nand U13769 (N_13769,N_12126,N_12604);
or U13770 (N_13770,N_12381,N_12155);
nand U13771 (N_13771,N_12770,N_12442);
nor U13772 (N_13772,N_12722,N_12830);
and U13773 (N_13773,N_12360,N_12951);
xor U13774 (N_13774,N_12440,N_12661);
nand U13775 (N_13775,N_12041,N_12825);
nand U13776 (N_13776,N_12184,N_12642);
nor U13777 (N_13777,N_12080,N_12674);
and U13778 (N_13778,N_12647,N_12800);
or U13779 (N_13779,N_12172,N_12391);
xnor U13780 (N_13780,N_12932,N_12808);
xor U13781 (N_13781,N_12458,N_12437);
and U13782 (N_13782,N_12076,N_12407);
or U13783 (N_13783,N_12183,N_12849);
xnor U13784 (N_13784,N_12773,N_12455);
nand U13785 (N_13785,N_12415,N_12241);
xor U13786 (N_13786,N_12834,N_12696);
nand U13787 (N_13787,N_12980,N_12963);
nand U13788 (N_13788,N_12339,N_12476);
or U13789 (N_13789,N_12070,N_12617);
or U13790 (N_13790,N_12359,N_12136);
and U13791 (N_13791,N_12431,N_12721);
nand U13792 (N_13792,N_12606,N_12516);
and U13793 (N_13793,N_12479,N_12121);
nor U13794 (N_13794,N_12850,N_12333);
or U13795 (N_13795,N_12953,N_12582);
nand U13796 (N_13796,N_12773,N_12390);
xor U13797 (N_13797,N_12157,N_12514);
nand U13798 (N_13798,N_12384,N_12952);
nand U13799 (N_13799,N_12391,N_12357);
and U13800 (N_13800,N_12740,N_12543);
nor U13801 (N_13801,N_12899,N_12263);
xnor U13802 (N_13802,N_12811,N_12985);
xor U13803 (N_13803,N_12510,N_12804);
nand U13804 (N_13804,N_12567,N_12891);
xnor U13805 (N_13805,N_12191,N_12485);
xnor U13806 (N_13806,N_12755,N_12771);
and U13807 (N_13807,N_12657,N_12155);
or U13808 (N_13808,N_12208,N_12097);
nand U13809 (N_13809,N_12641,N_12697);
xnor U13810 (N_13810,N_12680,N_12490);
nand U13811 (N_13811,N_12208,N_12627);
and U13812 (N_13812,N_12144,N_12895);
or U13813 (N_13813,N_12223,N_12718);
or U13814 (N_13814,N_12449,N_12622);
and U13815 (N_13815,N_12623,N_12505);
nand U13816 (N_13816,N_12646,N_12172);
and U13817 (N_13817,N_12636,N_12893);
nand U13818 (N_13818,N_12374,N_12917);
or U13819 (N_13819,N_12123,N_12482);
and U13820 (N_13820,N_12250,N_12096);
nor U13821 (N_13821,N_12470,N_12290);
xor U13822 (N_13822,N_12769,N_12211);
nor U13823 (N_13823,N_12512,N_12915);
nor U13824 (N_13824,N_12182,N_12278);
and U13825 (N_13825,N_12801,N_12731);
xor U13826 (N_13826,N_12260,N_12194);
and U13827 (N_13827,N_12611,N_12539);
xor U13828 (N_13828,N_12498,N_12232);
xnor U13829 (N_13829,N_12687,N_12924);
nor U13830 (N_13830,N_12604,N_12980);
xor U13831 (N_13831,N_12344,N_12055);
or U13832 (N_13832,N_12365,N_12150);
nand U13833 (N_13833,N_12493,N_12327);
or U13834 (N_13834,N_12636,N_12681);
and U13835 (N_13835,N_12249,N_12032);
and U13836 (N_13836,N_12444,N_12083);
nor U13837 (N_13837,N_12669,N_12906);
nand U13838 (N_13838,N_12560,N_12137);
or U13839 (N_13839,N_12106,N_12350);
xor U13840 (N_13840,N_12581,N_12881);
nor U13841 (N_13841,N_12092,N_12190);
and U13842 (N_13842,N_12059,N_12889);
or U13843 (N_13843,N_12428,N_12921);
nor U13844 (N_13844,N_12536,N_12176);
or U13845 (N_13845,N_12477,N_12799);
nor U13846 (N_13846,N_12882,N_12241);
and U13847 (N_13847,N_12088,N_12853);
nand U13848 (N_13848,N_12645,N_12406);
xor U13849 (N_13849,N_12950,N_12607);
nand U13850 (N_13850,N_12838,N_12213);
and U13851 (N_13851,N_12899,N_12442);
xnor U13852 (N_13852,N_12016,N_12282);
nor U13853 (N_13853,N_12472,N_12470);
xnor U13854 (N_13854,N_12315,N_12058);
nand U13855 (N_13855,N_12395,N_12360);
or U13856 (N_13856,N_12124,N_12316);
nand U13857 (N_13857,N_12141,N_12848);
xnor U13858 (N_13858,N_12909,N_12706);
or U13859 (N_13859,N_12459,N_12644);
xnor U13860 (N_13860,N_12009,N_12218);
and U13861 (N_13861,N_12326,N_12033);
or U13862 (N_13862,N_12985,N_12663);
or U13863 (N_13863,N_12504,N_12693);
and U13864 (N_13864,N_12076,N_12875);
xor U13865 (N_13865,N_12043,N_12793);
xor U13866 (N_13866,N_12957,N_12874);
xor U13867 (N_13867,N_12331,N_12094);
and U13868 (N_13868,N_12023,N_12037);
nand U13869 (N_13869,N_12857,N_12965);
xor U13870 (N_13870,N_12793,N_12366);
xor U13871 (N_13871,N_12038,N_12493);
xnor U13872 (N_13872,N_12974,N_12160);
nand U13873 (N_13873,N_12586,N_12102);
or U13874 (N_13874,N_12211,N_12725);
nand U13875 (N_13875,N_12196,N_12406);
xnor U13876 (N_13876,N_12909,N_12851);
and U13877 (N_13877,N_12685,N_12263);
nand U13878 (N_13878,N_12251,N_12125);
xor U13879 (N_13879,N_12367,N_12039);
xor U13880 (N_13880,N_12165,N_12485);
and U13881 (N_13881,N_12291,N_12984);
xnor U13882 (N_13882,N_12217,N_12445);
or U13883 (N_13883,N_12951,N_12629);
xor U13884 (N_13884,N_12106,N_12078);
or U13885 (N_13885,N_12800,N_12217);
nor U13886 (N_13886,N_12849,N_12161);
nor U13887 (N_13887,N_12695,N_12825);
nor U13888 (N_13888,N_12253,N_12616);
xor U13889 (N_13889,N_12683,N_12648);
and U13890 (N_13890,N_12986,N_12725);
or U13891 (N_13891,N_12972,N_12612);
nand U13892 (N_13892,N_12169,N_12502);
or U13893 (N_13893,N_12327,N_12711);
nor U13894 (N_13894,N_12906,N_12350);
nand U13895 (N_13895,N_12450,N_12852);
nand U13896 (N_13896,N_12384,N_12477);
nor U13897 (N_13897,N_12707,N_12654);
xnor U13898 (N_13898,N_12658,N_12055);
or U13899 (N_13899,N_12695,N_12478);
or U13900 (N_13900,N_12737,N_12293);
and U13901 (N_13901,N_12063,N_12632);
xnor U13902 (N_13902,N_12290,N_12392);
or U13903 (N_13903,N_12443,N_12942);
xnor U13904 (N_13904,N_12460,N_12792);
xor U13905 (N_13905,N_12275,N_12971);
xnor U13906 (N_13906,N_12320,N_12766);
nor U13907 (N_13907,N_12926,N_12860);
xnor U13908 (N_13908,N_12867,N_12521);
nor U13909 (N_13909,N_12837,N_12149);
or U13910 (N_13910,N_12490,N_12350);
nor U13911 (N_13911,N_12094,N_12019);
nor U13912 (N_13912,N_12622,N_12782);
nor U13913 (N_13913,N_12258,N_12461);
and U13914 (N_13914,N_12835,N_12784);
xor U13915 (N_13915,N_12395,N_12895);
nor U13916 (N_13916,N_12460,N_12005);
nor U13917 (N_13917,N_12735,N_12769);
nor U13918 (N_13918,N_12671,N_12675);
nand U13919 (N_13919,N_12460,N_12541);
nor U13920 (N_13920,N_12833,N_12990);
nor U13921 (N_13921,N_12249,N_12475);
nand U13922 (N_13922,N_12100,N_12657);
and U13923 (N_13923,N_12540,N_12750);
nand U13924 (N_13924,N_12088,N_12744);
or U13925 (N_13925,N_12845,N_12228);
xnor U13926 (N_13926,N_12096,N_12631);
and U13927 (N_13927,N_12212,N_12394);
xor U13928 (N_13928,N_12317,N_12448);
nand U13929 (N_13929,N_12419,N_12687);
nor U13930 (N_13930,N_12793,N_12772);
nand U13931 (N_13931,N_12105,N_12557);
or U13932 (N_13932,N_12964,N_12758);
or U13933 (N_13933,N_12536,N_12804);
or U13934 (N_13934,N_12265,N_12142);
nor U13935 (N_13935,N_12156,N_12871);
nor U13936 (N_13936,N_12781,N_12438);
xor U13937 (N_13937,N_12831,N_12667);
xor U13938 (N_13938,N_12225,N_12640);
xnor U13939 (N_13939,N_12490,N_12646);
nand U13940 (N_13940,N_12908,N_12812);
xnor U13941 (N_13941,N_12751,N_12308);
and U13942 (N_13942,N_12838,N_12074);
xor U13943 (N_13943,N_12693,N_12013);
nor U13944 (N_13944,N_12408,N_12133);
nand U13945 (N_13945,N_12983,N_12508);
xnor U13946 (N_13946,N_12072,N_12311);
and U13947 (N_13947,N_12807,N_12152);
nor U13948 (N_13948,N_12366,N_12546);
nand U13949 (N_13949,N_12705,N_12735);
nand U13950 (N_13950,N_12428,N_12816);
nor U13951 (N_13951,N_12911,N_12337);
xor U13952 (N_13952,N_12311,N_12894);
nor U13953 (N_13953,N_12707,N_12095);
nand U13954 (N_13954,N_12787,N_12972);
and U13955 (N_13955,N_12586,N_12994);
nand U13956 (N_13956,N_12680,N_12770);
and U13957 (N_13957,N_12145,N_12152);
nand U13958 (N_13958,N_12074,N_12678);
nor U13959 (N_13959,N_12220,N_12045);
and U13960 (N_13960,N_12754,N_12208);
or U13961 (N_13961,N_12511,N_12237);
nand U13962 (N_13962,N_12900,N_12272);
nand U13963 (N_13963,N_12478,N_12126);
xnor U13964 (N_13964,N_12058,N_12599);
or U13965 (N_13965,N_12619,N_12884);
or U13966 (N_13966,N_12752,N_12258);
xor U13967 (N_13967,N_12000,N_12629);
or U13968 (N_13968,N_12435,N_12771);
nand U13969 (N_13969,N_12352,N_12262);
xor U13970 (N_13970,N_12785,N_12496);
nor U13971 (N_13971,N_12699,N_12701);
or U13972 (N_13972,N_12251,N_12862);
and U13973 (N_13973,N_12046,N_12793);
or U13974 (N_13974,N_12878,N_12629);
and U13975 (N_13975,N_12348,N_12557);
or U13976 (N_13976,N_12409,N_12221);
nand U13977 (N_13977,N_12433,N_12902);
nand U13978 (N_13978,N_12450,N_12691);
or U13979 (N_13979,N_12622,N_12722);
xnor U13980 (N_13980,N_12774,N_12349);
xor U13981 (N_13981,N_12146,N_12153);
and U13982 (N_13982,N_12745,N_12203);
xor U13983 (N_13983,N_12174,N_12382);
and U13984 (N_13984,N_12521,N_12944);
xnor U13985 (N_13985,N_12557,N_12031);
or U13986 (N_13986,N_12910,N_12340);
nand U13987 (N_13987,N_12340,N_12246);
xor U13988 (N_13988,N_12908,N_12886);
and U13989 (N_13989,N_12930,N_12005);
and U13990 (N_13990,N_12798,N_12917);
or U13991 (N_13991,N_12599,N_12628);
xnor U13992 (N_13992,N_12977,N_12347);
nor U13993 (N_13993,N_12289,N_12908);
nand U13994 (N_13994,N_12558,N_12079);
or U13995 (N_13995,N_12861,N_12444);
or U13996 (N_13996,N_12406,N_12106);
or U13997 (N_13997,N_12652,N_12164);
nand U13998 (N_13998,N_12138,N_12505);
nand U13999 (N_13999,N_12305,N_12938);
nor U14000 (N_14000,N_13844,N_13707);
or U14001 (N_14001,N_13834,N_13024);
and U14002 (N_14002,N_13162,N_13668);
nor U14003 (N_14003,N_13877,N_13709);
nand U14004 (N_14004,N_13763,N_13519);
and U14005 (N_14005,N_13388,N_13674);
xnor U14006 (N_14006,N_13405,N_13224);
nor U14007 (N_14007,N_13489,N_13087);
nand U14008 (N_14008,N_13047,N_13886);
nand U14009 (N_14009,N_13068,N_13457);
xor U14010 (N_14010,N_13464,N_13708);
and U14011 (N_14011,N_13430,N_13310);
and U14012 (N_14012,N_13357,N_13583);
xnor U14013 (N_14013,N_13157,N_13397);
and U14014 (N_14014,N_13131,N_13158);
or U14015 (N_14015,N_13728,N_13656);
nand U14016 (N_14016,N_13505,N_13203);
nand U14017 (N_14017,N_13099,N_13644);
or U14018 (N_14018,N_13662,N_13268);
and U14019 (N_14019,N_13653,N_13904);
and U14020 (N_14020,N_13978,N_13150);
xnor U14021 (N_14021,N_13968,N_13765);
and U14022 (N_14022,N_13926,N_13743);
xor U14023 (N_14023,N_13970,N_13952);
xor U14024 (N_14024,N_13727,N_13487);
xor U14025 (N_14025,N_13616,N_13138);
and U14026 (N_14026,N_13034,N_13080);
or U14027 (N_14027,N_13869,N_13642);
or U14028 (N_14028,N_13614,N_13588);
and U14029 (N_14029,N_13584,N_13379);
xnor U14030 (N_14030,N_13324,N_13547);
nand U14031 (N_14031,N_13915,N_13619);
nor U14032 (N_14032,N_13331,N_13463);
and U14033 (N_14033,N_13714,N_13658);
xor U14034 (N_14034,N_13725,N_13675);
nand U14035 (N_14035,N_13028,N_13346);
or U14036 (N_14036,N_13939,N_13330);
xor U14037 (N_14037,N_13493,N_13638);
xor U14038 (N_14038,N_13839,N_13730);
and U14039 (N_14039,N_13450,N_13998);
nand U14040 (N_14040,N_13012,N_13825);
nand U14041 (N_14041,N_13353,N_13354);
nor U14042 (N_14042,N_13782,N_13913);
xnor U14043 (N_14043,N_13842,N_13374);
xor U14044 (N_14044,N_13733,N_13462);
xor U14045 (N_14045,N_13365,N_13221);
nor U14046 (N_14046,N_13009,N_13558);
and U14047 (N_14047,N_13855,N_13222);
and U14048 (N_14048,N_13192,N_13777);
nand U14049 (N_14049,N_13267,N_13861);
or U14050 (N_14050,N_13164,N_13309);
xor U14051 (N_14051,N_13077,N_13314);
nor U14052 (N_14052,N_13671,N_13485);
xnor U14053 (N_14053,N_13492,N_13041);
nor U14054 (N_14054,N_13677,N_13279);
nand U14055 (N_14055,N_13690,N_13836);
or U14056 (N_14056,N_13303,N_13982);
xnor U14057 (N_14057,N_13731,N_13278);
or U14058 (N_14058,N_13901,N_13997);
xnor U14059 (N_14059,N_13593,N_13476);
or U14060 (N_14060,N_13459,N_13337);
xor U14061 (N_14061,N_13738,N_13928);
and U14062 (N_14062,N_13561,N_13205);
or U14063 (N_14063,N_13623,N_13121);
xor U14064 (N_14064,N_13000,N_13029);
or U14065 (N_14065,N_13076,N_13033);
nand U14066 (N_14066,N_13816,N_13191);
or U14067 (N_14067,N_13994,N_13622);
nor U14068 (N_14068,N_13061,N_13055);
nand U14069 (N_14069,N_13697,N_13103);
nand U14070 (N_14070,N_13688,N_13789);
or U14071 (N_14071,N_13413,N_13498);
and U14072 (N_14072,N_13551,N_13426);
or U14073 (N_14073,N_13914,N_13691);
and U14074 (N_14074,N_13270,N_13585);
nand U14075 (N_14075,N_13235,N_13375);
nor U14076 (N_14076,N_13764,N_13899);
and U14077 (N_14077,N_13434,N_13830);
nor U14078 (N_14078,N_13535,N_13581);
and U14079 (N_14079,N_13945,N_13894);
nand U14080 (N_14080,N_13876,N_13518);
nand U14081 (N_14081,N_13655,N_13504);
nand U14082 (N_14082,N_13387,N_13868);
and U14083 (N_14083,N_13130,N_13665);
and U14084 (N_14084,N_13862,N_13128);
xor U14085 (N_14085,N_13546,N_13654);
or U14086 (N_14086,N_13944,N_13002);
xnor U14087 (N_14087,N_13516,N_13694);
xor U14088 (N_14088,N_13921,N_13470);
nor U14089 (N_14089,N_13596,N_13762);
or U14090 (N_14090,N_13597,N_13300);
nand U14091 (N_14091,N_13373,N_13805);
or U14092 (N_14092,N_13398,N_13417);
nor U14093 (N_14093,N_13163,N_13624);
xor U14094 (N_14094,N_13758,N_13075);
or U14095 (N_14095,N_13981,N_13408);
and U14096 (N_14096,N_13005,N_13237);
or U14097 (N_14097,N_13081,N_13600);
nor U14098 (N_14098,N_13084,N_13248);
xnor U14099 (N_14099,N_13643,N_13657);
or U14100 (N_14100,N_13511,N_13955);
nor U14101 (N_14101,N_13984,N_13119);
or U14102 (N_14102,N_13992,N_13380);
nor U14103 (N_14103,N_13160,N_13885);
xor U14104 (N_14104,N_13115,N_13796);
and U14105 (N_14105,N_13768,N_13907);
xor U14106 (N_14106,N_13848,N_13385);
xnor U14107 (N_14107,N_13801,N_13679);
or U14108 (N_14108,N_13094,N_13480);
nand U14109 (N_14109,N_13338,N_13858);
xnor U14110 (N_14110,N_13019,N_13118);
nor U14111 (N_14111,N_13017,N_13503);
nor U14112 (N_14112,N_13431,N_13578);
or U14113 (N_14113,N_13917,N_13053);
nor U14114 (N_14114,N_13317,N_13537);
nor U14115 (N_14115,N_13395,N_13064);
nor U14116 (N_14116,N_13711,N_13571);
or U14117 (N_14117,N_13739,N_13481);
nor U14118 (N_14118,N_13590,N_13197);
nand U14119 (N_14119,N_13681,N_13960);
xor U14120 (N_14120,N_13420,N_13569);
and U14121 (N_14121,N_13265,N_13608);
nor U14122 (N_14122,N_13069,N_13508);
and U14123 (N_14123,N_13559,N_13227);
and U14124 (N_14124,N_13078,N_13214);
and U14125 (N_14125,N_13401,N_13308);
and U14126 (N_14126,N_13941,N_13250);
xor U14127 (N_14127,N_13467,N_13785);
and U14128 (N_14128,N_13715,N_13766);
nor U14129 (N_14129,N_13276,N_13564);
xnor U14130 (N_14130,N_13108,N_13165);
nor U14131 (N_14131,N_13294,N_13021);
or U14132 (N_14132,N_13345,N_13933);
xnor U14133 (N_14133,N_13242,N_13827);
xnor U14134 (N_14134,N_13520,N_13734);
xor U14135 (N_14135,N_13682,N_13591);
and U14136 (N_14136,N_13719,N_13996);
nand U14137 (N_14137,N_13054,N_13577);
and U14138 (N_14138,N_13183,N_13910);
or U14139 (N_14139,N_13186,N_13274);
nor U14140 (N_14140,N_13972,N_13717);
xnor U14141 (N_14141,N_13252,N_13938);
or U14142 (N_14142,N_13510,N_13700);
and U14143 (N_14143,N_13137,N_13335);
nand U14144 (N_14144,N_13234,N_13142);
nand U14145 (N_14145,N_13219,N_13924);
and U14146 (N_14146,N_13453,N_13306);
nand U14147 (N_14147,N_13211,N_13815);
nor U14148 (N_14148,N_13501,N_13740);
and U14149 (N_14149,N_13347,N_13095);
and U14150 (N_14150,N_13223,N_13529);
and U14151 (N_14151,N_13440,N_13906);
nand U14152 (N_14152,N_13849,N_13576);
nor U14153 (N_14153,N_13935,N_13446);
nor U14154 (N_14154,N_13466,N_13478);
nand U14155 (N_14155,N_13874,N_13025);
and U14156 (N_14156,N_13788,N_13987);
or U14157 (N_14157,N_13540,N_13589);
xnor U14158 (N_14158,N_13760,N_13863);
xnor U14159 (N_14159,N_13358,N_13394);
nor U14160 (N_14160,N_13311,N_13857);
or U14161 (N_14161,N_13750,N_13942);
nor U14162 (N_14162,N_13007,N_13946);
nor U14163 (N_14163,N_13079,N_13134);
and U14164 (N_14164,N_13652,N_13925);
nor U14165 (N_14165,N_13930,N_13199);
nor U14166 (N_14166,N_13436,N_13177);
nor U14167 (N_14167,N_13646,N_13524);
nand U14168 (N_14168,N_13587,N_13795);
nand U14169 (N_14169,N_13473,N_13621);
xnor U14170 (N_14170,N_13568,N_13916);
or U14171 (N_14171,N_13172,N_13692);
xor U14172 (N_14172,N_13049,N_13180);
nand U14173 (N_14173,N_13835,N_13536);
and U14174 (N_14174,N_13565,N_13898);
xnor U14175 (N_14175,N_13672,N_13947);
nand U14176 (N_14176,N_13455,N_13831);
or U14177 (N_14177,N_13297,N_13553);
or U14178 (N_14178,N_13149,N_13056);
and U14179 (N_14179,N_13141,N_13490);
and U14180 (N_14180,N_13384,N_13598);
nor U14181 (N_14181,N_13271,N_13920);
or U14182 (N_14182,N_13132,N_13684);
xor U14183 (N_14183,N_13046,N_13889);
or U14184 (N_14184,N_13555,N_13011);
or U14185 (N_14185,N_13023,N_13366);
xnor U14186 (N_14186,N_13295,N_13236);
xnor U14187 (N_14187,N_13648,N_13350);
or U14188 (N_14188,N_13231,N_13549);
nand U14189 (N_14189,N_13949,N_13631);
nand U14190 (N_14190,N_13514,N_13783);
xor U14191 (N_14191,N_13104,N_13178);
nand U14192 (N_14192,N_13040,N_13018);
nand U14193 (N_14193,N_13479,N_13402);
and U14194 (N_14194,N_13494,N_13367);
xor U14195 (N_14195,N_13666,N_13418);
nor U14196 (N_14196,N_13745,N_13291);
nor U14197 (N_14197,N_13735,N_13628);
xnor U14198 (N_14198,N_13964,N_13275);
xor U14199 (N_14199,N_13340,N_13850);
and U14200 (N_14200,N_13573,N_13723);
and U14201 (N_14201,N_13202,N_13313);
nand U14202 (N_14202,N_13477,N_13976);
or U14203 (N_14203,N_13454,N_13048);
or U14204 (N_14204,N_13841,N_13030);
nor U14205 (N_14205,N_13020,N_13167);
or U14206 (N_14206,N_13890,N_13482);
and U14207 (N_14207,N_13198,N_13441);
xor U14208 (N_14208,N_13022,N_13066);
or U14209 (N_14209,N_13107,N_13400);
nand U14210 (N_14210,N_13206,N_13190);
and U14211 (N_14211,N_13574,N_13208);
nand U14212 (N_14212,N_13074,N_13315);
nor U14213 (N_14213,N_13249,N_13264);
and U14214 (N_14214,N_13756,N_13837);
and U14215 (N_14215,N_13599,N_13154);
and U14216 (N_14216,N_13959,N_13680);
or U14217 (N_14217,N_13060,N_13209);
or U14218 (N_14218,N_13305,N_13845);
xnor U14219 (N_14219,N_13484,N_13273);
nand U14220 (N_14220,N_13355,N_13859);
or U14221 (N_14221,N_13193,N_13606);
nand U14222 (N_14222,N_13050,N_13755);
or U14223 (N_14223,N_13369,N_13932);
nor U14224 (N_14224,N_13348,N_13342);
nor U14225 (N_14225,N_13804,N_13534);
nand U14226 (N_14226,N_13423,N_13851);
nand U14227 (N_14227,N_13176,N_13336);
xnor U14228 (N_14228,N_13229,N_13749);
xnor U14229 (N_14229,N_13286,N_13098);
xor U14230 (N_14230,N_13770,N_13230);
or U14231 (N_14231,N_13184,N_13334);
nor U14232 (N_14232,N_13761,N_13406);
nor U14233 (N_14233,N_13386,N_13509);
or U14234 (N_14234,N_13109,N_13042);
or U14235 (N_14235,N_13092,N_13757);
nand U14236 (N_14236,N_13635,N_13082);
xor U14237 (N_14237,N_13262,N_13882);
nand U14238 (N_14238,N_13556,N_13327);
nand U14239 (N_14239,N_13032,N_13759);
xor U14240 (N_14240,N_13403,N_13813);
or U14241 (N_14241,N_13878,N_13567);
nor U14242 (N_14242,N_13883,N_13856);
or U14243 (N_14243,N_13775,N_13979);
nand U14244 (N_14244,N_13962,N_13895);
xnor U14245 (N_14245,N_13085,N_13751);
and U14246 (N_14246,N_13439,N_13343);
xnor U14247 (N_14247,N_13880,N_13560);
nand U14248 (N_14248,N_13152,N_13148);
nand U14249 (N_14249,N_13438,N_13116);
or U14250 (N_14250,N_13052,N_13543);
nor U14251 (N_14251,N_13840,N_13156);
xor U14252 (N_14252,N_13341,N_13687);
xnor U14253 (N_14253,N_13826,N_13531);
nor U14254 (N_14254,N_13277,N_13713);
xnor U14255 (N_14255,N_13124,N_13429);
nand U14256 (N_14256,N_13639,N_13433);
or U14257 (N_14257,N_13168,N_13371);
nand U14258 (N_14258,N_13506,N_13318);
nor U14259 (N_14259,N_13187,N_13557);
nand U14260 (N_14260,N_13604,N_13483);
or U14261 (N_14261,N_13120,N_13256);
nand U14262 (N_14262,N_13522,N_13442);
xnor U14263 (N_14263,N_13810,N_13182);
nor U14264 (N_14264,N_13062,N_13685);
xnor U14265 (N_14265,N_13961,N_13888);
and U14266 (N_14266,N_13196,N_13105);
or U14267 (N_14267,N_13144,N_13607);
nor U14268 (N_14268,N_13710,N_13281);
xnor U14269 (N_14269,N_13983,N_13189);
xor U14270 (N_14270,N_13383,N_13702);
or U14271 (N_14271,N_13974,N_13382);
xor U14272 (N_14272,N_13797,N_13865);
and U14273 (N_14273,N_13969,N_13500);
nand U14274 (N_14274,N_13111,N_13833);
and U14275 (N_14275,N_13039,N_13329);
nor U14276 (N_14276,N_13263,N_13634);
xnor U14277 (N_14277,N_13207,N_13389);
nor U14278 (N_14278,N_13891,N_13261);
and U14279 (N_14279,N_13852,N_13284);
nor U14280 (N_14280,N_13332,N_13517);
xnor U14281 (N_14281,N_13823,N_13333);
xnor U14282 (N_14282,N_13288,N_13807);
and U14283 (N_14283,N_13580,N_13404);
and U14284 (N_14284,N_13127,N_13239);
nor U14285 (N_14285,N_13471,N_13474);
xor U14286 (N_14286,N_13247,N_13747);
nor U14287 (N_14287,N_13806,N_13044);
and U14288 (N_14288,N_13488,N_13486);
or U14289 (N_14289,N_13999,N_13737);
nor U14290 (N_14290,N_13159,N_13610);
xor U14291 (N_14291,N_13732,N_13746);
and U14292 (N_14292,N_13843,N_13396);
and U14293 (N_14293,N_13004,N_13258);
nor U14294 (N_14294,N_13822,N_13122);
nand U14295 (N_14295,N_13173,N_13376);
or U14296 (N_14296,N_13633,N_13544);
xor U14297 (N_14297,N_13245,N_13563);
or U14298 (N_14298,N_13298,N_13475);
xnor U14299 (N_14299,N_13254,N_13499);
and U14300 (N_14300,N_13110,N_13013);
nor U14301 (N_14301,N_13113,N_13432);
xor U14302 (N_14302,N_13659,N_13472);
nor U14303 (N_14303,N_13465,N_13444);
nand U14304 (N_14304,N_13900,N_13582);
xnor U14305 (N_14305,N_13377,N_13650);
or U14306 (N_14306,N_13909,N_13051);
nor U14307 (N_14307,N_13502,N_13636);
nand U14308 (N_14308,N_13809,N_13447);
nor U14309 (N_14309,N_13512,N_13781);
nor U14310 (N_14310,N_13542,N_13112);
nor U14311 (N_14311,N_13716,N_13640);
nand U14312 (N_14312,N_13322,N_13927);
and U14313 (N_14313,N_13873,N_13414);
and U14314 (N_14314,N_13627,N_13545);
or U14315 (N_14315,N_13072,N_13200);
xnor U14316 (N_14316,N_13527,N_13201);
nand U14317 (N_14317,N_13670,N_13391);
or U14318 (N_14318,N_13461,N_13253);
nor U14319 (N_14319,N_13778,N_13566);
nor U14320 (N_14320,N_13696,N_13411);
and U14321 (N_14321,N_13323,N_13307);
xor U14322 (N_14322,N_13014,N_13218);
and U14323 (N_14323,N_13602,N_13325);
nor U14324 (N_14324,N_13793,N_13174);
nand U14325 (N_14325,N_13922,N_13721);
xor U14326 (N_14326,N_13101,N_13854);
xnor U14327 (N_14327,N_13609,N_13421);
or U14328 (N_14328,N_13879,N_13686);
xnor U14329 (N_14329,N_13703,N_13412);
nand U14330 (N_14330,N_13975,N_13001);
and U14331 (N_14331,N_13864,N_13817);
xnor U14332 (N_14332,N_13963,N_13695);
or U14333 (N_14333,N_13729,N_13361);
nand U14334 (N_14334,N_13896,N_13605);
xnor U14335 (N_14335,N_13067,N_13010);
nand U14336 (N_14336,N_13683,N_13272);
nor U14337 (N_14337,N_13541,N_13803);
and U14338 (N_14338,N_13993,N_13575);
or U14339 (N_14339,N_13460,N_13991);
or U14340 (N_14340,N_13289,N_13603);
or U14341 (N_14341,N_13181,N_13929);
nor U14342 (N_14342,N_13956,N_13513);
nand U14343 (N_14343,N_13045,N_13496);
xnor U14344 (N_14344,N_13892,N_13445);
and U14345 (N_14345,N_13296,N_13523);
xnor U14346 (N_14346,N_13497,N_13409);
or U14347 (N_14347,N_13615,N_13415);
nor U14348 (N_14348,N_13469,N_13748);
xor U14349 (N_14349,N_13136,N_13867);
xor U14350 (N_14350,N_13808,N_13943);
xnor U14351 (N_14351,N_13903,N_13967);
nor U14352 (N_14352,N_13706,N_13424);
nor U14353 (N_14353,N_13106,N_13086);
and U14354 (N_14354,N_13073,N_13378);
and U14355 (N_14355,N_13422,N_13918);
and U14356 (N_14356,N_13008,N_13986);
or U14357 (N_14357,N_13720,N_13491);
nor U14358 (N_14358,N_13741,N_13282);
or U14359 (N_14359,N_13003,N_13293);
and U14360 (N_14360,N_13824,N_13255);
and U14361 (N_14361,N_13170,N_13416);
and U14362 (N_14362,N_13287,N_13872);
or U14363 (N_14363,N_13973,N_13035);
and U14364 (N_14364,N_13651,N_13515);
xnor U14365 (N_14365,N_13037,N_13283);
nand U14366 (N_14366,N_13435,N_13215);
and U14367 (N_14367,N_13736,N_13526);
nand U14368 (N_14368,N_13776,N_13953);
or U14369 (N_14369,N_13989,N_13228);
and U14370 (N_14370,N_13812,N_13893);
and U14371 (N_14371,N_13292,N_13226);
nor U14372 (N_14372,N_13853,N_13951);
nand U14373 (N_14373,N_13269,N_13611);
nand U14374 (N_14374,N_13618,N_13241);
nand U14375 (N_14375,N_13027,N_13114);
or U14376 (N_14376,N_13097,N_13847);
or U14377 (N_14377,N_13990,N_13699);
nor U14378 (N_14378,N_13133,N_13507);
nand U14379 (N_14379,N_13664,N_13161);
and U14380 (N_14380,N_13673,N_13356);
nor U14381 (N_14381,N_13015,N_13320);
or U14382 (N_14382,N_13592,N_13285);
or U14383 (N_14383,N_13351,N_13135);
or U14384 (N_14384,N_13773,N_13316);
or U14385 (N_14385,N_13630,N_13179);
nor U14386 (N_14386,N_13689,N_13620);
nand U14387 (N_14387,N_13784,N_13771);
xor U14388 (N_14388,N_13821,N_13233);
xor U14389 (N_14389,N_13579,N_13767);
nand U14390 (N_14390,N_13676,N_13870);
or U14391 (N_14391,N_13971,N_13246);
xnor U14392 (N_14392,N_13667,N_13212);
nand U14393 (N_14393,N_13155,N_13220);
nand U14394 (N_14394,N_13328,N_13452);
xor U14395 (N_14395,N_13145,N_13458);
and U14396 (N_14396,N_13586,N_13065);
nand U14397 (N_14397,N_13902,N_13096);
nand U14398 (N_14398,N_13570,N_13613);
or U14399 (N_14399,N_13059,N_13923);
nor U14400 (N_14400,N_13251,N_13143);
or U14401 (N_14401,N_13931,N_13661);
or U14402 (N_14402,N_13381,N_13629);
or U14403 (N_14403,N_13985,N_13153);
xnor U14404 (N_14404,N_13393,N_13216);
xor U14405 (N_14405,N_13832,N_13299);
and U14406 (N_14406,N_13185,N_13232);
nor U14407 (N_14407,N_13742,N_13058);
nand U14408 (N_14408,N_13301,N_13139);
nand U14409 (N_14409,N_13495,N_13780);
and U14410 (N_14410,N_13779,N_13372);
and U14411 (N_14411,N_13266,N_13102);
or U14412 (N_14412,N_13147,N_13940);
nor U14413 (N_14413,N_13828,N_13213);
nand U14414 (N_14414,N_13954,N_13123);
and U14415 (N_14415,N_13753,N_13669);
or U14416 (N_14416,N_13026,N_13319);
nand U14417 (N_14417,N_13769,N_13698);
nor U14418 (N_14418,N_13911,N_13533);
or U14419 (N_14419,N_13754,N_13977);
or U14420 (N_14420,N_13399,N_13626);
and U14421 (N_14421,N_13908,N_13774);
or U14422 (N_14422,N_13070,N_13705);
nor U14423 (N_14423,N_13091,N_13090);
nor U14424 (N_14424,N_13772,N_13290);
xnor U14425 (N_14425,N_13093,N_13129);
and U14426 (N_14426,N_13359,N_13428);
xnor U14427 (N_14427,N_13194,N_13016);
xor U14428 (N_14428,N_13169,N_13649);
and U14429 (N_14429,N_13811,N_13260);
nand U14430 (N_14430,N_13663,N_13860);
or U14431 (N_14431,N_13846,N_13820);
or U14432 (N_14432,N_13410,N_13538);
and U14433 (N_14433,N_13425,N_13243);
xor U14434 (N_14434,N_13238,N_13456);
xor U14435 (N_14435,N_13304,N_13443);
and U14436 (N_14436,N_13884,N_13548);
nand U14437 (N_14437,N_13966,N_13368);
and U14438 (N_14438,N_13678,N_13038);
xnor U14439 (N_14439,N_13752,N_13125);
and U14440 (N_14440,N_13427,N_13244);
and U14441 (N_14441,N_13552,N_13521);
nand U14442 (N_14442,N_13819,N_13259);
and U14443 (N_14443,N_13724,N_13875);
xor U14444 (N_14444,N_13370,N_13140);
nor U14445 (N_14445,N_13866,N_13195);
or U14446 (N_14446,N_13031,N_13006);
and U14447 (N_14447,N_13958,N_13791);
xor U14448 (N_14448,N_13829,N_13794);
nand U14449 (N_14449,N_13595,N_13204);
nor U14450 (N_14450,N_13637,N_13530);
xor U14451 (N_14451,N_13572,N_13965);
or U14452 (N_14452,N_13802,N_13468);
and U14453 (N_14453,N_13948,N_13407);
xor U14454 (N_14454,N_13838,N_13887);
xnor U14455 (N_14455,N_13071,N_13344);
xnor U14456 (N_14456,N_13100,N_13800);
nand U14457 (N_14457,N_13449,N_13641);
and U14458 (N_14458,N_13326,N_13339);
xnor U14459 (N_14459,N_13448,N_13792);
nor U14460 (N_14460,N_13188,N_13126);
or U14461 (N_14461,N_13988,N_13704);
nand U14462 (N_14462,N_13360,N_13088);
nand U14463 (N_14463,N_13645,N_13151);
and U14464 (N_14464,N_13257,N_13722);
nor U14465 (N_14465,N_13363,N_13349);
or U14466 (N_14466,N_13043,N_13392);
nand U14467 (N_14467,N_13146,N_13647);
nand U14468 (N_14468,N_13225,N_13787);
and U14469 (N_14469,N_13818,N_13612);
and U14470 (N_14470,N_13934,N_13550);
xnor U14471 (N_14471,N_13995,N_13790);
xor U14472 (N_14472,N_13897,N_13919);
xor U14473 (N_14473,N_13217,N_13799);
nand U14474 (N_14474,N_13364,N_13210);
or U14475 (N_14475,N_13451,N_13562);
or U14476 (N_14476,N_13871,N_13718);
or U14477 (N_14477,N_13693,N_13701);
or U14478 (N_14478,N_13083,N_13390);
and U14479 (N_14479,N_13744,N_13594);
nand U14480 (N_14480,N_13280,N_13632);
and U14481 (N_14481,N_13936,N_13532);
nor U14482 (N_14482,N_13798,N_13419);
and U14483 (N_14483,N_13980,N_13117);
or U14484 (N_14484,N_13712,N_13554);
xnor U14485 (N_14485,N_13617,N_13321);
nand U14486 (N_14486,N_13312,N_13166);
nand U14487 (N_14487,N_13437,N_13171);
nor U14488 (N_14488,N_13539,N_13814);
or U14489 (N_14489,N_13786,N_13240);
xor U14490 (N_14490,N_13525,N_13528);
xor U14491 (N_14491,N_13950,N_13063);
nand U14492 (N_14492,N_13175,N_13302);
and U14493 (N_14493,N_13625,N_13937);
nand U14494 (N_14494,N_13089,N_13362);
or U14495 (N_14495,N_13957,N_13352);
xor U14496 (N_14496,N_13881,N_13905);
nor U14497 (N_14497,N_13660,N_13601);
xor U14498 (N_14498,N_13036,N_13726);
or U14499 (N_14499,N_13057,N_13912);
xor U14500 (N_14500,N_13292,N_13582);
xnor U14501 (N_14501,N_13712,N_13202);
xnor U14502 (N_14502,N_13658,N_13539);
nand U14503 (N_14503,N_13805,N_13169);
nand U14504 (N_14504,N_13590,N_13841);
xnor U14505 (N_14505,N_13710,N_13406);
and U14506 (N_14506,N_13336,N_13301);
and U14507 (N_14507,N_13341,N_13003);
xnor U14508 (N_14508,N_13585,N_13820);
nor U14509 (N_14509,N_13976,N_13664);
and U14510 (N_14510,N_13651,N_13318);
and U14511 (N_14511,N_13855,N_13309);
nand U14512 (N_14512,N_13530,N_13705);
nor U14513 (N_14513,N_13576,N_13808);
nand U14514 (N_14514,N_13998,N_13391);
and U14515 (N_14515,N_13108,N_13329);
nor U14516 (N_14516,N_13092,N_13362);
and U14517 (N_14517,N_13803,N_13859);
and U14518 (N_14518,N_13657,N_13408);
nand U14519 (N_14519,N_13111,N_13137);
and U14520 (N_14520,N_13887,N_13452);
xor U14521 (N_14521,N_13048,N_13581);
nand U14522 (N_14522,N_13650,N_13569);
xor U14523 (N_14523,N_13562,N_13075);
or U14524 (N_14524,N_13514,N_13191);
xor U14525 (N_14525,N_13237,N_13802);
nor U14526 (N_14526,N_13088,N_13097);
xnor U14527 (N_14527,N_13015,N_13715);
xnor U14528 (N_14528,N_13763,N_13308);
nand U14529 (N_14529,N_13829,N_13084);
or U14530 (N_14530,N_13209,N_13157);
or U14531 (N_14531,N_13132,N_13422);
nor U14532 (N_14532,N_13280,N_13412);
nor U14533 (N_14533,N_13164,N_13942);
nand U14534 (N_14534,N_13375,N_13933);
xnor U14535 (N_14535,N_13712,N_13128);
or U14536 (N_14536,N_13788,N_13668);
nor U14537 (N_14537,N_13168,N_13084);
nor U14538 (N_14538,N_13607,N_13279);
xnor U14539 (N_14539,N_13509,N_13910);
or U14540 (N_14540,N_13175,N_13299);
nand U14541 (N_14541,N_13046,N_13844);
nor U14542 (N_14542,N_13239,N_13523);
or U14543 (N_14543,N_13338,N_13980);
and U14544 (N_14544,N_13856,N_13297);
or U14545 (N_14545,N_13648,N_13822);
xnor U14546 (N_14546,N_13136,N_13336);
xor U14547 (N_14547,N_13972,N_13014);
nor U14548 (N_14548,N_13339,N_13225);
or U14549 (N_14549,N_13240,N_13709);
and U14550 (N_14550,N_13829,N_13403);
nand U14551 (N_14551,N_13289,N_13952);
and U14552 (N_14552,N_13840,N_13032);
and U14553 (N_14553,N_13339,N_13127);
nand U14554 (N_14554,N_13333,N_13070);
or U14555 (N_14555,N_13502,N_13023);
or U14556 (N_14556,N_13653,N_13447);
nor U14557 (N_14557,N_13483,N_13202);
nor U14558 (N_14558,N_13775,N_13033);
nor U14559 (N_14559,N_13693,N_13525);
xor U14560 (N_14560,N_13201,N_13532);
xnor U14561 (N_14561,N_13679,N_13907);
xor U14562 (N_14562,N_13810,N_13263);
or U14563 (N_14563,N_13857,N_13780);
xor U14564 (N_14564,N_13995,N_13817);
nor U14565 (N_14565,N_13635,N_13603);
nor U14566 (N_14566,N_13617,N_13969);
nor U14567 (N_14567,N_13684,N_13803);
nor U14568 (N_14568,N_13366,N_13308);
xnor U14569 (N_14569,N_13064,N_13850);
xnor U14570 (N_14570,N_13030,N_13945);
nand U14571 (N_14571,N_13604,N_13754);
and U14572 (N_14572,N_13125,N_13842);
xor U14573 (N_14573,N_13290,N_13237);
xnor U14574 (N_14574,N_13634,N_13810);
xnor U14575 (N_14575,N_13571,N_13122);
and U14576 (N_14576,N_13716,N_13215);
and U14577 (N_14577,N_13475,N_13807);
nor U14578 (N_14578,N_13464,N_13494);
xnor U14579 (N_14579,N_13230,N_13657);
nor U14580 (N_14580,N_13742,N_13036);
nand U14581 (N_14581,N_13653,N_13694);
and U14582 (N_14582,N_13870,N_13740);
or U14583 (N_14583,N_13386,N_13456);
xor U14584 (N_14584,N_13191,N_13131);
or U14585 (N_14585,N_13157,N_13088);
and U14586 (N_14586,N_13888,N_13601);
and U14587 (N_14587,N_13842,N_13393);
and U14588 (N_14588,N_13541,N_13038);
and U14589 (N_14589,N_13362,N_13456);
or U14590 (N_14590,N_13419,N_13090);
nor U14591 (N_14591,N_13064,N_13588);
and U14592 (N_14592,N_13248,N_13858);
nand U14593 (N_14593,N_13802,N_13721);
xor U14594 (N_14594,N_13555,N_13280);
nor U14595 (N_14595,N_13418,N_13452);
or U14596 (N_14596,N_13108,N_13031);
or U14597 (N_14597,N_13981,N_13698);
or U14598 (N_14598,N_13535,N_13446);
nand U14599 (N_14599,N_13103,N_13154);
or U14600 (N_14600,N_13910,N_13721);
and U14601 (N_14601,N_13041,N_13657);
and U14602 (N_14602,N_13771,N_13946);
and U14603 (N_14603,N_13229,N_13148);
nor U14604 (N_14604,N_13732,N_13607);
xor U14605 (N_14605,N_13330,N_13930);
and U14606 (N_14606,N_13077,N_13839);
or U14607 (N_14607,N_13739,N_13331);
xor U14608 (N_14608,N_13486,N_13931);
or U14609 (N_14609,N_13494,N_13322);
and U14610 (N_14610,N_13987,N_13037);
nor U14611 (N_14611,N_13611,N_13420);
nor U14612 (N_14612,N_13380,N_13549);
nand U14613 (N_14613,N_13363,N_13396);
nand U14614 (N_14614,N_13957,N_13569);
nor U14615 (N_14615,N_13628,N_13761);
nor U14616 (N_14616,N_13476,N_13704);
and U14617 (N_14617,N_13605,N_13879);
nand U14618 (N_14618,N_13078,N_13463);
nor U14619 (N_14619,N_13890,N_13860);
nor U14620 (N_14620,N_13073,N_13478);
nand U14621 (N_14621,N_13477,N_13406);
nor U14622 (N_14622,N_13807,N_13200);
xor U14623 (N_14623,N_13141,N_13189);
nand U14624 (N_14624,N_13993,N_13302);
and U14625 (N_14625,N_13127,N_13277);
xnor U14626 (N_14626,N_13147,N_13370);
nand U14627 (N_14627,N_13287,N_13931);
and U14628 (N_14628,N_13219,N_13836);
nand U14629 (N_14629,N_13435,N_13476);
or U14630 (N_14630,N_13961,N_13917);
and U14631 (N_14631,N_13372,N_13750);
nand U14632 (N_14632,N_13453,N_13102);
nand U14633 (N_14633,N_13713,N_13087);
xnor U14634 (N_14634,N_13487,N_13295);
or U14635 (N_14635,N_13337,N_13450);
nand U14636 (N_14636,N_13987,N_13443);
xor U14637 (N_14637,N_13109,N_13438);
or U14638 (N_14638,N_13239,N_13431);
or U14639 (N_14639,N_13615,N_13499);
nand U14640 (N_14640,N_13678,N_13641);
nor U14641 (N_14641,N_13442,N_13445);
or U14642 (N_14642,N_13239,N_13418);
nand U14643 (N_14643,N_13607,N_13351);
nand U14644 (N_14644,N_13820,N_13043);
or U14645 (N_14645,N_13359,N_13688);
nand U14646 (N_14646,N_13435,N_13711);
and U14647 (N_14647,N_13199,N_13664);
nand U14648 (N_14648,N_13335,N_13871);
or U14649 (N_14649,N_13757,N_13046);
xnor U14650 (N_14650,N_13958,N_13816);
nor U14651 (N_14651,N_13904,N_13271);
xor U14652 (N_14652,N_13986,N_13029);
nor U14653 (N_14653,N_13746,N_13069);
and U14654 (N_14654,N_13922,N_13944);
nor U14655 (N_14655,N_13659,N_13432);
nor U14656 (N_14656,N_13524,N_13050);
and U14657 (N_14657,N_13913,N_13936);
and U14658 (N_14658,N_13110,N_13966);
nor U14659 (N_14659,N_13828,N_13473);
xnor U14660 (N_14660,N_13111,N_13828);
or U14661 (N_14661,N_13995,N_13173);
nor U14662 (N_14662,N_13372,N_13476);
nor U14663 (N_14663,N_13124,N_13663);
xnor U14664 (N_14664,N_13649,N_13230);
or U14665 (N_14665,N_13085,N_13813);
xnor U14666 (N_14666,N_13311,N_13540);
nor U14667 (N_14667,N_13821,N_13021);
or U14668 (N_14668,N_13027,N_13359);
nor U14669 (N_14669,N_13255,N_13122);
nand U14670 (N_14670,N_13208,N_13115);
or U14671 (N_14671,N_13917,N_13470);
nand U14672 (N_14672,N_13594,N_13255);
and U14673 (N_14673,N_13832,N_13510);
xor U14674 (N_14674,N_13207,N_13117);
nand U14675 (N_14675,N_13688,N_13248);
and U14676 (N_14676,N_13225,N_13314);
and U14677 (N_14677,N_13795,N_13083);
and U14678 (N_14678,N_13307,N_13936);
nand U14679 (N_14679,N_13457,N_13322);
nor U14680 (N_14680,N_13293,N_13370);
and U14681 (N_14681,N_13459,N_13579);
or U14682 (N_14682,N_13147,N_13495);
xor U14683 (N_14683,N_13620,N_13132);
nand U14684 (N_14684,N_13774,N_13718);
and U14685 (N_14685,N_13501,N_13931);
or U14686 (N_14686,N_13513,N_13905);
nor U14687 (N_14687,N_13164,N_13706);
or U14688 (N_14688,N_13742,N_13489);
nor U14689 (N_14689,N_13950,N_13152);
and U14690 (N_14690,N_13723,N_13507);
or U14691 (N_14691,N_13270,N_13188);
nand U14692 (N_14692,N_13908,N_13915);
xor U14693 (N_14693,N_13458,N_13059);
and U14694 (N_14694,N_13496,N_13579);
or U14695 (N_14695,N_13903,N_13755);
nor U14696 (N_14696,N_13591,N_13771);
nor U14697 (N_14697,N_13774,N_13230);
nor U14698 (N_14698,N_13944,N_13247);
or U14699 (N_14699,N_13326,N_13307);
nor U14700 (N_14700,N_13297,N_13857);
nand U14701 (N_14701,N_13867,N_13331);
nor U14702 (N_14702,N_13573,N_13267);
nand U14703 (N_14703,N_13566,N_13940);
or U14704 (N_14704,N_13247,N_13164);
xnor U14705 (N_14705,N_13101,N_13668);
nor U14706 (N_14706,N_13156,N_13946);
and U14707 (N_14707,N_13412,N_13108);
xnor U14708 (N_14708,N_13624,N_13708);
nand U14709 (N_14709,N_13850,N_13917);
or U14710 (N_14710,N_13220,N_13126);
and U14711 (N_14711,N_13310,N_13951);
or U14712 (N_14712,N_13093,N_13717);
nand U14713 (N_14713,N_13102,N_13308);
or U14714 (N_14714,N_13911,N_13513);
xor U14715 (N_14715,N_13098,N_13956);
nand U14716 (N_14716,N_13758,N_13459);
nor U14717 (N_14717,N_13623,N_13142);
nand U14718 (N_14718,N_13494,N_13973);
nor U14719 (N_14719,N_13026,N_13508);
nand U14720 (N_14720,N_13931,N_13476);
nand U14721 (N_14721,N_13666,N_13636);
or U14722 (N_14722,N_13789,N_13248);
xnor U14723 (N_14723,N_13297,N_13896);
or U14724 (N_14724,N_13214,N_13971);
nand U14725 (N_14725,N_13772,N_13693);
xnor U14726 (N_14726,N_13195,N_13256);
or U14727 (N_14727,N_13387,N_13031);
xor U14728 (N_14728,N_13625,N_13610);
nor U14729 (N_14729,N_13664,N_13776);
nand U14730 (N_14730,N_13229,N_13582);
and U14731 (N_14731,N_13530,N_13263);
nor U14732 (N_14732,N_13219,N_13066);
nand U14733 (N_14733,N_13734,N_13542);
and U14734 (N_14734,N_13967,N_13045);
or U14735 (N_14735,N_13757,N_13634);
or U14736 (N_14736,N_13114,N_13871);
nor U14737 (N_14737,N_13297,N_13038);
nor U14738 (N_14738,N_13792,N_13584);
or U14739 (N_14739,N_13158,N_13724);
nand U14740 (N_14740,N_13682,N_13762);
and U14741 (N_14741,N_13160,N_13396);
xnor U14742 (N_14742,N_13799,N_13961);
nand U14743 (N_14743,N_13870,N_13282);
nand U14744 (N_14744,N_13943,N_13099);
nor U14745 (N_14745,N_13670,N_13580);
or U14746 (N_14746,N_13621,N_13452);
nor U14747 (N_14747,N_13294,N_13528);
or U14748 (N_14748,N_13109,N_13582);
nand U14749 (N_14749,N_13159,N_13980);
and U14750 (N_14750,N_13562,N_13042);
and U14751 (N_14751,N_13779,N_13251);
xnor U14752 (N_14752,N_13297,N_13719);
nor U14753 (N_14753,N_13362,N_13747);
nor U14754 (N_14754,N_13876,N_13849);
nor U14755 (N_14755,N_13479,N_13974);
nand U14756 (N_14756,N_13283,N_13338);
and U14757 (N_14757,N_13948,N_13931);
or U14758 (N_14758,N_13344,N_13041);
nand U14759 (N_14759,N_13940,N_13562);
xor U14760 (N_14760,N_13983,N_13175);
or U14761 (N_14761,N_13030,N_13004);
and U14762 (N_14762,N_13343,N_13460);
nor U14763 (N_14763,N_13980,N_13944);
nand U14764 (N_14764,N_13492,N_13702);
xor U14765 (N_14765,N_13706,N_13603);
nor U14766 (N_14766,N_13034,N_13048);
or U14767 (N_14767,N_13383,N_13306);
or U14768 (N_14768,N_13404,N_13182);
nand U14769 (N_14769,N_13813,N_13275);
or U14770 (N_14770,N_13135,N_13499);
or U14771 (N_14771,N_13929,N_13171);
nand U14772 (N_14772,N_13004,N_13970);
xnor U14773 (N_14773,N_13921,N_13399);
or U14774 (N_14774,N_13638,N_13970);
nand U14775 (N_14775,N_13405,N_13071);
xor U14776 (N_14776,N_13346,N_13870);
nand U14777 (N_14777,N_13683,N_13170);
nor U14778 (N_14778,N_13991,N_13228);
nand U14779 (N_14779,N_13838,N_13323);
and U14780 (N_14780,N_13295,N_13653);
nand U14781 (N_14781,N_13933,N_13266);
nand U14782 (N_14782,N_13581,N_13485);
xnor U14783 (N_14783,N_13773,N_13841);
and U14784 (N_14784,N_13962,N_13649);
nand U14785 (N_14785,N_13206,N_13737);
xnor U14786 (N_14786,N_13096,N_13837);
or U14787 (N_14787,N_13793,N_13263);
or U14788 (N_14788,N_13866,N_13389);
or U14789 (N_14789,N_13768,N_13881);
xnor U14790 (N_14790,N_13346,N_13461);
or U14791 (N_14791,N_13076,N_13517);
nand U14792 (N_14792,N_13571,N_13308);
nor U14793 (N_14793,N_13498,N_13028);
nor U14794 (N_14794,N_13625,N_13572);
and U14795 (N_14795,N_13787,N_13168);
nand U14796 (N_14796,N_13385,N_13525);
nand U14797 (N_14797,N_13875,N_13554);
nand U14798 (N_14798,N_13983,N_13477);
xnor U14799 (N_14799,N_13947,N_13989);
xor U14800 (N_14800,N_13015,N_13617);
or U14801 (N_14801,N_13864,N_13137);
nand U14802 (N_14802,N_13636,N_13514);
or U14803 (N_14803,N_13312,N_13257);
nor U14804 (N_14804,N_13969,N_13615);
xnor U14805 (N_14805,N_13248,N_13443);
and U14806 (N_14806,N_13364,N_13701);
nor U14807 (N_14807,N_13943,N_13211);
and U14808 (N_14808,N_13775,N_13435);
and U14809 (N_14809,N_13779,N_13034);
xor U14810 (N_14810,N_13226,N_13462);
xor U14811 (N_14811,N_13045,N_13578);
and U14812 (N_14812,N_13325,N_13894);
nand U14813 (N_14813,N_13516,N_13128);
or U14814 (N_14814,N_13954,N_13719);
xnor U14815 (N_14815,N_13383,N_13873);
and U14816 (N_14816,N_13298,N_13086);
and U14817 (N_14817,N_13064,N_13808);
nand U14818 (N_14818,N_13306,N_13319);
or U14819 (N_14819,N_13239,N_13277);
and U14820 (N_14820,N_13485,N_13932);
xnor U14821 (N_14821,N_13285,N_13329);
and U14822 (N_14822,N_13637,N_13406);
xor U14823 (N_14823,N_13917,N_13487);
xnor U14824 (N_14824,N_13205,N_13052);
and U14825 (N_14825,N_13874,N_13947);
xor U14826 (N_14826,N_13484,N_13646);
or U14827 (N_14827,N_13439,N_13727);
xnor U14828 (N_14828,N_13310,N_13031);
nand U14829 (N_14829,N_13238,N_13786);
nor U14830 (N_14830,N_13701,N_13256);
and U14831 (N_14831,N_13786,N_13548);
and U14832 (N_14832,N_13563,N_13501);
nor U14833 (N_14833,N_13020,N_13256);
and U14834 (N_14834,N_13194,N_13853);
or U14835 (N_14835,N_13968,N_13563);
or U14836 (N_14836,N_13466,N_13154);
or U14837 (N_14837,N_13812,N_13920);
nand U14838 (N_14838,N_13821,N_13763);
nand U14839 (N_14839,N_13561,N_13624);
and U14840 (N_14840,N_13549,N_13580);
xnor U14841 (N_14841,N_13361,N_13581);
nand U14842 (N_14842,N_13758,N_13884);
or U14843 (N_14843,N_13461,N_13104);
and U14844 (N_14844,N_13571,N_13163);
xor U14845 (N_14845,N_13344,N_13208);
nor U14846 (N_14846,N_13548,N_13685);
nor U14847 (N_14847,N_13553,N_13536);
nor U14848 (N_14848,N_13799,N_13936);
xnor U14849 (N_14849,N_13713,N_13456);
and U14850 (N_14850,N_13698,N_13453);
or U14851 (N_14851,N_13185,N_13985);
xor U14852 (N_14852,N_13203,N_13971);
nand U14853 (N_14853,N_13332,N_13221);
nand U14854 (N_14854,N_13218,N_13792);
or U14855 (N_14855,N_13766,N_13535);
and U14856 (N_14856,N_13277,N_13593);
or U14857 (N_14857,N_13909,N_13132);
and U14858 (N_14858,N_13251,N_13538);
and U14859 (N_14859,N_13765,N_13762);
and U14860 (N_14860,N_13418,N_13226);
xnor U14861 (N_14861,N_13584,N_13662);
or U14862 (N_14862,N_13074,N_13440);
and U14863 (N_14863,N_13455,N_13542);
xnor U14864 (N_14864,N_13722,N_13097);
and U14865 (N_14865,N_13068,N_13178);
nand U14866 (N_14866,N_13982,N_13406);
nor U14867 (N_14867,N_13830,N_13291);
and U14868 (N_14868,N_13938,N_13360);
and U14869 (N_14869,N_13055,N_13475);
nand U14870 (N_14870,N_13315,N_13756);
or U14871 (N_14871,N_13174,N_13376);
and U14872 (N_14872,N_13808,N_13408);
nor U14873 (N_14873,N_13490,N_13256);
or U14874 (N_14874,N_13603,N_13391);
xnor U14875 (N_14875,N_13208,N_13879);
nand U14876 (N_14876,N_13413,N_13761);
or U14877 (N_14877,N_13310,N_13504);
nand U14878 (N_14878,N_13843,N_13208);
and U14879 (N_14879,N_13820,N_13677);
nand U14880 (N_14880,N_13400,N_13792);
nand U14881 (N_14881,N_13789,N_13241);
or U14882 (N_14882,N_13889,N_13629);
xnor U14883 (N_14883,N_13968,N_13238);
nor U14884 (N_14884,N_13037,N_13196);
xor U14885 (N_14885,N_13505,N_13698);
and U14886 (N_14886,N_13230,N_13666);
or U14887 (N_14887,N_13934,N_13543);
or U14888 (N_14888,N_13781,N_13927);
xor U14889 (N_14889,N_13653,N_13481);
nand U14890 (N_14890,N_13777,N_13061);
nand U14891 (N_14891,N_13234,N_13727);
nand U14892 (N_14892,N_13128,N_13696);
nor U14893 (N_14893,N_13777,N_13911);
or U14894 (N_14894,N_13645,N_13374);
or U14895 (N_14895,N_13942,N_13153);
or U14896 (N_14896,N_13516,N_13597);
xnor U14897 (N_14897,N_13846,N_13061);
nand U14898 (N_14898,N_13694,N_13815);
or U14899 (N_14899,N_13422,N_13024);
xor U14900 (N_14900,N_13158,N_13257);
nand U14901 (N_14901,N_13029,N_13961);
xor U14902 (N_14902,N_13937,N_13365);
and U14903 (N_14903,N_13582,N_13979);
nand U14904 (N_14904,N_13650,N_13801);
nor U14905 (N_14905,N_13072,N_13787);
nor U14906 (N_14906,N_13723,N_13626);
nor U14907 (N_14907,N_13532,N_13402);
or U14908 (N_14908,N_13142,N_13137);
nand U14909 (N_14909,N_13378,N_13704);
nor U14910 (N_14910,N_13972,N_13452);
nor U14911 (N_14911,N_13587,N_13155);
or U14912 (N_14912,N_13059,N_13898);
nand U14913 (N_14913,N_13401,N_13060);
nand U14914 (N_14914,N_13029,N_13856);
nand U14915 (N_14915,N_13968,N_13489);
or U14916 (N_14916,N_13266,N_13201);
and U14917 (N_14917,N_13722,N_13607);
xor U14918 (N_14918,N_13561,N_13230);
and U14919 (N_14919,N_13930,N_13904);
nand U14920 (N_14920,N_13356,N_13089);
and U14921 (N_14921,N_13609,N_13840);
and U14922 (N_14922,N_13292,N_13055);
and U14923 (N_14923,N_13256,N_13113);
and U14924 (N_14924,N_13946,N_13247);
nor U14925 (N_14925,N_13111,N_13491);
nor U14926 (N_14926,N_13836,N_13895);
xnor U14927 (N_14927,N_13845,N_13809);
or U14928 (N_14928,N_13951,N_13581);
or U14929 (N_14929,N_13735,N_13206);
or U14930 (N_14930,N_13935,N_13626);
or U14931 (N_14931,N_13959,N_13077);
nand U14932 (N_14932,N_13263,N_13991);
nor U14933 (N_14933,N_13478,N_13705);
nand U14934 (N_14934,N_13161,N_13156);
nor U14935 (N_14935,N_13013,N_13851);
nand U14936 (N_14936,N_13462,N_13094);
and U14937 (N_14937,N_13258,N_13135);
or U14938 (N_14938,N_13373,N_13311);
xor U14939 (N_14939,N_13659,N_13295);
nand U14940 (N_14940,N_13535,N_13941);
nor U14941 (N_14941,N_13293,N_13248);
or U14942 (N_14942,N_13780,N_13931);
nand U14943 (N_14943,N_13977,N_13290);
nand U14944 (N_14944,N_13059,N_13650);
nand U14945 (N_14945,N_13145,N_13131);
nor U14946 (N_14946,N_13587,N_13147);
nor U14947 (N_14947,N_13783,N_13920);
and U14948 (N_14948,N_13498,N_13785);
xnor U14949 (N_14949,N_13020,N_13216);
and U14950 (N_14950,N_13887,N_13285);
xnor U14951 (N_14951,N_13656,N_13116);
nor U14952 (N_14952,N_13073,N_13864);
and U14953 (N_14953,N_13916,N_13865);
and U14954 (N_14954,N_13033,N_13819);
xor U14955 (N_14955,N_13484,N_13781);
xor U14956 (N_14956,N_13235,N_13579);
or U14957 (N_14957,N_13192,N_13627);
xnor U14958 (N_14958,N_13509,N_13681);
xnor U14959 (N_14959,N_13101,N_13272);
xor U14960 (N_14960,N_13817,N_13718);
xnor U14961 (N_14961,N_13076,N_13673);
or U14962 (N_14962,N_13738,N_13081);
and U14963 (N_14963,N_13228,N_13130);
nand U14964 (N_14964,N_13425,N_13061);
and U14965 (N_14965,N_13812,N_13010);
nor U14966 (N_14966,N_13416,N_13953);
xnor U14967 (N_14967,N_13820,N_13067);
or U14968 (N_14968,N_13083,N_13004);
nor U14969 (N_14969,N_13764,N_13540);
and U14970 (N_14970,N_13125,N_13979);
nor U14971 (N_14971,N_13668,N_13438);
xnor U14972 (N_14972,N_13766,N_13401);
nand U14973 (N_14973,N_13195,N_13390);
and U14974 (N_14974,N_13027,N_13717);
xnor U14975 (N_14975,N_13893,N_13704);
and U14976 (N_14976,N_13320,N_13597);
nand U14977 (N_14977,N_13448,N_13277);
and U14978 (N_14978,N_13379,N_13560);
xor U14979 (N_14979,N_13511,N_13099);
or U14980 (N_14980,N_13674,N_13472);
xnor U14981 (N_14981,N_13564,N_13157);
or U14982 (N_14982,N_13039,N_13800);
nand U14983 (N_14983,N_13605,N_13321);
nor U14984 (N_14984,N_13614,N_13575);
nor U14985 (N_14985,N_13300,N_13096);
nor U14986 (N_14986,N_13821,N_13297);
and U14987 (N_14987,N_13681,N_13195);
nand U14988 (N_14988,N_13220,N_13657);
nor U14989 (N_14989,N_13273,N_13759);
and U14990 (N_14990,N_13573,N_13387);
nand U14991 (N_14991,N_13741,N_13141);
and U14992 (N_14992,N_13965,N_13083);
xor U14993 (N_14993,N_13989,N_13364);
xnor U14994 (N_14994,N_13870,N_13684);
xor U14995 (N_14995,N_13774,N_13732);
or U14996 (N_14996,N_13772,N_13647);
nor U14997 (N_14997,N_13712,N_13379);
xor U14998 (N_14998,N_13857,N_13609);
or U14999 (N_14999,N_13432,N_13298);
or U15000 (N_15000,N_14822,N_14696);
and U15001 (N_15001,N_14996,N_14232);
nor U15002 (N_15002,N_14906,N_14915);
and U15003 (N_15003,N_14623,N_14757);
xnor U15004 (N_15004,N_14876,N_14719);
xor U15005 (N_15005,N_14358,N_14523);
or U15006 (N_15006,N_14040,N_14254);
and U15007 (N_15007,N_14508,N_14647);
or U15008 (N_15008,N_14433,N_14924);
and U15009 (N_15009,N_14660,N_14718);
nor U15010 (N_15010,N_14609,N_14484);
nand U15011 (N_15011,N_14051,N_14415);
xor U15012 (N_15012,N_14676,N_14751);
and U15013 (N_15013,N_14223,N_14105);
or U15014 (N_15014,N_14395,N_14429);
or U15015 (N_15015,N_14825,N_14371);
xnor U15016 (N_15016,N_14158,N_14553);
nor U15017 (N_15017,N_14313,N_14188);
and U15018 (N_15018,N_14635,N_14020);
nor U15019 (N_15019,N_14170,N_14761);
xnor U15020 (N_15020,N_14134,N_14092);
and U15021 (N_15021,N_14887,N_14971);
xor U15022 (N_15022,N_14943,N_14330);
nand U15023 (N_15023,N_14815,N_14545);
xnor U15024 (N_15024,N_14162,N_14805);
nand U15025 (N_15025,N_14893,N_14275);
and U15026 (N_15026,N_14533,N_14151);
and U15027 (N_15027,N_14240,N_14620);
nor U15028 (N_15028,N_14849,N_14382);
xor U15029 (N_15029,N_14299,N_14651);
and U15030 (N_15030,N_14550,N_14540);
and U15031 (N_15031,N_14043,N_14854);
or U15032 (N_15032,N_14695,N_14776);
nor U15033 (N_15033,N_14673,N_14074);
or U15034 (N_15034,N_14572,N_14501);
or U15035 (N_15035,N_14013,N_14820);
and U15036 (N_15036,N_14594,N_14072);
and U15037 (N_15037,N_14455,N_14000);
nand U15038 (N_15038,N_14225,N_14627);
nand U15039 (N_15039,N_14125,N_14866);
nand U15040 (N_15040,N_14454,N_14988);
xnor U15041 (N_15041,N_14301,N_14667);
xnor U15042 (N_15042,N_14704,N_14048);
and U15043 (N_15043,N_14588,N_14833);
or U15044 (N_15044,N_14009,N_14787);
or U15045 (N_15045,N_14999,N_14003);
nand U15046 (N_15046,N_14546,N_14570);
and U15047 (N_15047,N_14715,N_14894);
nand U15048 (N_15048,N_14103,N_14412);
nand U15049 (N_15049,N_14154,N_14390);
and U15050 (N_15050,N_14872,N_14184);
nor U15051 (N_15051,N_14591,N_14164);
nor U15052 (N_15052,N_14381,N_14414);
xor U15053 (N_15053,N_14802,N_14038);
and U15054 (N_15054,N_14206,N_14773);
nand U15055 (N_15055,N_14486,N_14227);
or U15056 (N_15056,N_14175,N_14099);
and U15057 (N_15057,N_14470,N_14265);
and U15058 (N_15058,N_14049,N_14474);
or U15059 (N_15059,N_14185,N_14131);
xnor U15060 (N_15060,N_14927,N_14293);
xnor U15061 (N_15061,N_14693,N_14803);
xor U15062 (N_15062,N_14913,N_14018);
or U15063 (N_15063,N_14949,N_14650);
nand U15064 (N_15064,N_14136,N_14129);
and U15065 (N_15065,N_14289,N_14441);
nor U15066 (N_15066,N_14936,N_14912);
and U15067 (N_15067,N_14375,N_14215);
and U15068 (N_15068,N_14961,N_14359);
nand U15069 (N_15069,N_14574,N_14785);
nor U15070 (N_15070,N_14211,N_14780);
nor U15071 (N_15071,N_14118,N_14080);
nand U15072 (N_15072,N_14955,N_14939);
and U15073 (N_15073,N_14919,N_14442);
xor U15074 (N_15074,N_14675,N_14644);
and U15075 (N_15075,N_14513,N_14436);
xnor U15076 (N_15076,N_14909,N_14882);
and U15077 (N_15077,N_14427,N_14604);
nand U15078 (N_15078,N_14400,N_14498);
or U15079 (N_15079,N_14034,N_14132);
or U15080 (N_15080,N_14182,N_14527);
nor U15081 (N_15081,N_14317,N_14365);
xor U15082 (N_15082,N_14333,N_14016);
nand U15083 (N_15083,N_14023,N_14662);
and U15084 (N_15084,N_14385,N_14249);
nor U15085 (N_15085,N_14189,N_14210);
nor U15086 (N_15086,N_14422,N_14257);
and U15087 (N_15087,N_14446,N_14665);
nand U15088 (N_15088,N_14898,N_14198);
nand U15089 (N_15089,N_14266,N_14236);
nand U15090 (N_15090,N_14777,N_14658);
or U15091 (N_15091,N_14139,N_14378);
nand U15092 (N_15092,N_14119,N_14838);
nor U15093 (N_15093,N_14011,N_14443);
or U15094 (N_15094,N_14711,N_14668);
and U15095 (N_15095,N_14832,N_14408);
xor U15096 (N_15096,N_14699,N_14753);
or U15097 (N_15097,N_14302,N_14810);
xnor U15098 (N_15098,N_14253,N_14113);
or U15099 (N_15099,N_14497,N_14464);
and U15100 (N_15100,N_14272,N_14672);
nor U15101 (N_15101,N_14111,N_14953);
nand U15102 (N_15102,N_14858,N_14790);
nor U15103 (N_15103,N_14307,N_14165);
and U15104 (N_15104,N_14723,N_14772);
nand U15105 (N_15105,N_14602,N_14694);
nor U15106 (N_15106,N_14143,N_14937);
and U15107 (N_15107,N_14774,N_14601);
nor U15108 (N_15108,N_14260,N_14640);
or U15109 (N_15109,N_14798,N_14179);
and U15110 (N_15110,N_14918,N_14622);
or U15111 (N_15111,N_14745,N_14027);
nor U15112 (N_15112,N_14108,N_14852);
nor U15113 (N_15113,N_14499,N_14311);
nor U15114 (N_15114,N_14053,N_14706);
nor U15115 (N_15115,N_14702,N_14507);
or U15116 (N_15116,N_14259,N_14328);
or U15117 (N_15117,N_14207,N_14794);
nand U15118 (N_15118,N_14251,N_14823);
and U15119 (N_15119,N_14713,N_14735);
nor U15120 (N_15120,N_14959,N_14697);
nand U15121 (N_15121,N_14308,N_14855);
or U15122 (N_15122,N_14922,N_14021);
or U15123 (N_15123,N_14122,N_14345);
and U15124 (N_15124,N_14703,N_14343);
and U15125 (N_15125,N_14944,N_14112);
and U15126 (N_15126,N_14933,N_14033);
and U15127 (N_15127,N_14440,N_14263);
or U15128 (N_15128,N_14298,N_14568);
nor U15129 (N_15129,N_14377,N_14710);
nor U15130 (N_15130,N_14789,N_14071);
or U15131 (N_15131,N_14459,N_14629);
nand U15132 (N_15132,N_14467,N_14914);
and U15133 (N_15133,N_14052,N_14046);
xor U15134 (N_15134,N_14290,N_14683);
and U15135 (N_15135,N_14091,N_14521);
or U15136 (N_15136,N_14727,N_14851);
nor U15137 (N_15137,N_14754,N_14584);
and U15138 (N_15138,N_14800,N_14194);
xnor U15139 (N_15139,N_14280,N_14639);
xnor U15140 (N_15140,N_14321,N_14881);
or U15141 (N_15141,N_14309,N_14434);
and U15142 (N_15142,N_14305,N_14001);
xnor U15143 (N_15143,N_14682,N_14342);
nand U15144 (N_15144,N_14892,N_14690);
xor U15145 (N_15145,N_14461,N_14234);
and U15146 (N_15146,N_14193,N_14063);
xor U15147 (N_15147,N_14654,N_14793);
xor U15148 (N_15148,N_14085,N_14191);
and U15149 (N_15149,N_14804,N_14149);
and U15150 (N_15150,N_14750,N_14039);
nor U15151 (N_15151,N_14235,N_14487);
and U15152 (N_15152,N_14144,N_14140);
nor U15153 (N_15153,N_14397,N_14760);
xnor U15154 (N_15154,N_14445,N_14929);
nor U15155 (N_15155,N_14073,N_14525);
or U15156 (N_15156,N_14784,N_14503);
or U15157 (N_15157,N_14743,N_14324);
nor U15158 (N_15158,N_14086,N_14169);
nor U15159 (N_15159,N_14161,N_14566);
or U15160 (N_15160,N_14560,N_14244);
or U15161 (N_15161,N_14109,N_14237);
or U15162 (N_15162,N_14983,N_14421);
nand U15163 (N_15163,N_14732,N_14347);
and U15164 (N_15164,N_14870,N_14628);
and U15165 (N_15165,N_14065,N_14864);
and U15166 (N_15166,N_14426,N_14625);
nor U15167 (N_15167,N_14138,N_14535);
and U15168 (N_15168,N_14469,N_14731);
nor U15169 (N_15169,N_14425,N_14576);
and U15170 (N_15170,N_14167,N_14128);
and U15171 (N_15171,N_14500,N_14734);
or U15172 (N_15172,N_14663,N_14270);
nand U15173 (N_15173,N_14981,N_14571);
nor U15174 (N_15174,N_14649,N_14782);
and U15175 (N_15175,N_14879,N_14368);
or U15176 (N_15176,N_14997,N_14173);
and U15177 (N_15177,N_14520,N_14146);
and U15178 (N_15178,N_14972,N_14895);
or U15179 (N_15179,N_14808,N_14722);
or U15180 (N_15180,N_14982,N_14351);
xor U15181 (N_15181,N_14468,N_14615);
or U15182 (N_15182,N_14819,N_14025);
nand U15183 (N_15183,N_14960,N_14813);
nor U15184 (N_15184,N_14726,N_14314);
xor U15185 (N_15185,N_14582,N_14796);
xnor U15186 (N_15186,N_14472,N_14012);
xor U15187 (N_15187,N_14712,N_14869);
and U15188 (N_15188,N_14142,N_14689);
and U15189 (N_15189,N_14202,N_14465);
or U15190 (N_15190,N_14097,N_14471);
and U15191 (N_15191,N_14495,N_14245);
or U15192 (N_15192,N_14603,N_14199);
nor U15193 (N_15193,N_14957,N_14766);
nand U15194 (N_15194,N_14453,N_14332);
and U15195 (N_15195,N_14203,N_14637);
nand U15196 (N_15196,N_14004,N_14231);
nand U15197 (N_15197,N_14995,N_14653);
nand U15198 (N_15198,N_14536,N_14386);
and U15199 (N_15199,N_14075,N_14531);
xnor U15200 (N_15200,N_14897,N_14606);
and U15201 (N_15201,N_14951,N_14352);
nand U15202 (N_15202,N_14462,N_14666);
nor U15203 (N_15203,N_14456,N_14806);
nor U15204 (N_15204,N_14764,N_14466);
nor U15205 (N_15205,N_14526,N_14172);
and U15206 (N_15206,N_14197,N_14739);
xor U15207 (N_15207,N_14567,N_14853);
nand U15208 (N_15208,N_14032,N_14014);
or U15209 (N_15209,N_14195,N_14979);
nand U15210 (N_15210,N_14066,N_14130);
or U15211 (N_15211,N_14926,N_14056);
and U15212 (N_15212,N_14857,N_14886);
xor U15213 (N_15213,N_14835,N_14076);
nor U15214 (N_15214,N_14127,N_14044);
and U15215 (N_15215,N_14600,N_14786);
xor U15216 (N_15216,N_14110,N_14084);
nand U15217 (N_15217,N_14911,N_14792);
and U15218 (N_15218,N_14423,N_14973);
xor U15219 (N_15219,N_14543,N_14967);
nor U15220 (N_15220,N_14831,N_14950);
or U15221 (N_15221,N_14476,N_14717);
and U15222 (N_15222,N_14791,N_14411);
nand U15223 (N_15223,N_14372,N_14392);
nor U15224 (N_15224,N_14241,N_14860);
nand U15225 (N_15225,N_14163,N_14827);
nor U15226 (N_15226,N_14756,N_14370);
nand U15227 (N_15227,N_14413,N_14424);
nor U15228 (N_15228,N_14532,N_14348);
nand U15229 (N_15229,N_14367,N_14990);
nor U15230 (N_15230,N_14209,N_14537);
nor U15231 (N_15231,N_14871,N_14190);
nand U15232 (N_15232,N_14511,N_14361);
xor U15233 (N_15233,N_14589,N_14363);
nand U15234 (N_15234,N_14267,N_14171);
nand U15235 (N_15235,N_14264,N_14082);
xor U15236 (N_15236,N_14376,N_14047);
or U15237 (N_15237,N_14248,N_14283);
xor U15238 (N_15238,N_14318,N_14315);
xnor U15239 (N_15239,N_14035,N_14277);
nand U15240 (N_15240,N_14002,N_14554);
and U15241 (N_15241,N_14399,N_14291);
nand U15242 (N_15242,N_14077,N_14387);
and U15243 (N_15243,N_14258,N_14181);
xor U15244 (N_15244,N_14137,N_14799);
nand U15245 (N_15245,N_14975,N_14920);
or U15246 (N_15246,N_14360,N_14222);
nand U15247 (N_15247,N_14910,N_14458);
nand U15248 (N_15248,N_14998,N_14384);
and U15249 (N_15249,N_14050,N_14389);
nand U15250 (N_15250,N_14153,N_14457);
nand U15251 (N_15251,N_14485,N_14841);
nand U15252 (N_15252,N_14610,N_14037);
nor U15253 (N_15253,N_14934,N_14707);
and U15254 (N_15254,N_14337,N_14089);
and U15255 (N_15255,N_14010,N_14948);
and U15256 (N_15256,N_14326,N_14274);
nand U15257 (N_15257,N_14709,N_14765);
xnor U15258 (N_15258,N_14678,N_14724);
nand U15259 (N_15259,N_14670,N_14573);
and U15260 (N_15260,N_14396,N_14908);
nand U15261 (N_15261,N_14017,N_14094);
or U15262 (N_15262,N_14090,N_14530);
and U15263 (N_15263,N_14705,N_14968);
nor U15264 (N_15264,N_14157,N_14217);
xor U15265 (N_15265,N_14904,N_14518);
and U15266 (N_15266,N_14221,N_14150);
xor U15267 (N_15267,N_14252,N_14821);
xnor U15268 (N_15268,N_14636,N_14312);
nor U15269 (N_15269,N_14563,N_14698);
or U15270 (N_15270,N_14681,N_14036);
or U15271 (N_15271,N_14716,N_14026);
nand U15272 (N_15272,N_14816,N_14657);
or U15273 (N_15273,N_14942,N_14155);
xnor U15274 (N_15274,N_14310,N_14515);
and U15275 (N_15275,N_14986,N_14059);
xor U15276 (N_15276,N_14133,N_14510);
and U15277 (N_15277,N_14938,N_14120);
nor U15278 (N_15278,N_14323,N_14448);
or U15279 (N_15279,N_14561,N_14394);
nor U15280 (N_15280,N_14580,N_14250);
nand U15281 (N_15281,N_14737,N_14867);
and U15282 (N_15282,N_14522,N_14256);
or U15283 (N_15283,N_14980,N_14547);
nor U15284 (N_15284,N_14325,N_14428);
nor U15285 (N_15285,N_14528,N_14230);
and U15286 (N_15286,N_14405,N_14616);
and U15287 (N_15287,N_14863,N_14512);
nor U15288 (N_15288,N_14836,N_14407);
xor U15289 (N_15289,N_14888,N_14839);
xor U15290 (N_15290,N_14555,N_14964);
xor U15291 (N_15291,N_14124,N_14339);
xor U15292 (N_15292,N_14208,N_14374);
nand U15293 (N_15293,N_14862,N_14795);
nand U15294 (N_15294,N_14941,N_14945);
nor U15295 (N_15295,N_14905,N_14954);
and U15296 (N_15296,N_14061,N_14054);
nor U15297 (N_15297,N_14204,N_14783);
or U15298 (N_15298,N_14692,N_14885);
nor U15299 (N_15299,N_14993,N_14304);
or U15300 (N_15300,N_14218,N_14874);
and U15301 (N_15301,N_14398,N_14369);
and U15302 (N_15302,N_14030,N_14549);
and U15303 (N_15303,N_14024,N_14435);
and U15304 (N_15304,N_14294,N_14115);
xor U15305 (N_15305,N_14238,N_14788);
nand U15306 (N_15306,N_14093,N_14873);
and U15307 (N_15307,N_14336,N_14509);
or U15308 (N_15308,N_14357,N_14460);
or U15309 (N_15309,N_14450,N_14444);
or U15310 (N_15310,N_14877,N_14147);
nand U15311 (N_15311,N_14192,N_14917);
nor U15312 (N_15312,N_14963,N_14978);
nor U15313 (N_15313,N_14214,N_14187);
xnor U15314 (N_15314,N_14556,N_14581);
xor U15315 (N_15315,N_14952,N_14008);
nand U15316 (N_15316,N_14341,N_14826);
and U15317 (N_15317,N_14007,N_14686);
or U15318 (N_15318,N_14220,N_14834);
nor U15319 (N_15319,N_14300,N_14814);
xor U15320 (N_15320,N_14430,N_14101);
nand U15321 (N_15321,N_14432,N_14262);
nand U15322 (N_15322,N_14356,N_14940);
nand U15323 (N_15323,N_14329,N_14552);
nand U15324 (N_15324,N_14279,N_14159);
or U15325 (N_15325,N_14327,N_14102);
nor U15326 (N_15326,N_14031,N_14233);
nand U15327 (N_15327,N_14539,N_14402);
nand U15328 (N_15328,N_14156,N_14551);
and U15329 (N_15329,N_14725,N_14742);
nand U15330 (N_15330,N_14284,N_14491);
or U15331 (N_15331,N_14664,N_14579);
nand U15332 (N_15332,N_14062,N_14504);
nor U15333 (N_15333,N_14976,N_14496);
and U15334 (N_15334,N_14614,N_14104);
and U15335 (N_15335,N_14216,N_14956);
nand U15336 (N_15336,N_14303,N_14296);
nand U15337 (N_15337,N_14344,N_14088);
nand U15338 (N_15338,N_14631,N_14516);
xor U15339 (N_15339,N_14899,N_14656);
nor U15340 (N_15340,N_14517,N_14987);
nor U15341 (N_15341,N_14379,N_14060);
or U15342 (N_15342,N_14685,N_14847);
or U15343 (N_15343,N_14564,N_14687);
and U15344 (N_15344,N_14519,N_14481);
or U15345 (N_15345,N_14648,N_14618);
and U15346 (N_15346,N_14596,N_14095);
or U15347 (N_15347,N_14067,N_14166);
xnor U15348 (N_15348,N_14482,N_14632);
and U15349 (N_15349,N_14652,N_14506);
nor U15350 (N_15350,N_14946,N_14100);
xnor U15351 (N_15351,N_14022,N_14655);
nand U15352 (N_15352,N_14684,N_14607);
and U15353 (N_15353,N_14403,N_14593);
xor U15354 (N_15354,N_14985,N_14830);
or U15355 (N_15355,N_14630,N_14592);
or U15356 (N_15356,N_14295,N_14930);
nor U15357 (N_15357,N_14542,N_14213);
nor U15358 (N_15358,N_14762,N_14078);
nand U15359 (N_15359,N_14322,N_14569);
or U15360 (N_15360,N_14598,N_14177);
nor U15361 (N_15361,N_14281,N_14057);
and U15362 (N_15362,N_14015,N_14041);
or U15363 (N_15363,N_14416,N_14451);
or U15364 (N_15364,N_14005,N_14633);
xor U15365 (N_15365,N_14107,N_14843);
and U15366 (N_15366,N_14889,N_14969);
xor U15367 (N_15367,N_14994,N_14478);
or U15368 (N_15368,N_14406,N_14900);
and U15369 (N_15369,N_14708,N_14316);
nand U15370 (N_15370,N_14276,N_14064);
nand U15371 (N_15371,N_14287,N_14224);
or U15372 (N_15372,N_14720,N_14779);
and U15373 (N_15373,N_14768,N_14931);
nand U15374 (N_15374,N_14055,N_14634);
xor U15375 (N_15375,N_14729,N_14514);
nor U15376 (N_15376,N_14587,N_14744);
and U15377 (N_15377,N_14431,N_14028);
xnor U15378 (N_15378,N_14176,N_14261);
or U15379 (N_15379,N_14247,N_14671);
nor U15380 (N_15380,N_14809,N_14770);
and U15381 (N_15381,N_14674,N_14494);
xnor U15382 (N_15382,N_14970,N_14006);
nand U15383 (N_15383,N_14868,N_14740);
and U15384 (N_15384,N_14292,N_14346);
nor U15385 (N_15385,N_14958,N_14114);
nor U15386 (N_15386,N_14680,N_14410);
nor U15387 (N_15387,N_14439,N_14180);
and U15388 (N_15388,N_14070,N_14160);
or U15389 (N_15389,N_14763,N_14388);
nor U15390 (N_15390,N_14271,N_14595);
and U15391 (N_15391,N_14965,N_14320);
nand U15392 (N_15392,N_14557,N_14558);
nor U15393 (N_15393,N_14212,N_14420);
nor U15394 (N_15394,N_14121,N_14242);
and U15395 (N_15395,N_14174,N_14452);
nand U15396 (N_15396,N_14850,N_14123);
and U15397 (N_15397,N_14349,N_14925);
xnor U15398 (N_15398,N_14087,N_14611);
or U15399 (N_15399,N_14391,N_14642);
nand U15400 (N_15400,N_14183,N_14890);
nor U15401 (N_15401,N_14880,N_14383);
and U15402 (N_15402,N_14624,N_14490);
or U15403 (N_15403,N_14083,N_14643);
nand U15404 (N_15404,N_14229,N_14449);
xor U15405 (N_15405,N_14974,N_14544);
and U15406 (N_15406,N_14688,N_14058);
xor U15407 (N_15407,N_14947,N_14338);
and U15408 (N_15408,N_14362,N_14273);
and U15409 (N_15409,N_14691,N_14529);
and U15410 (N_15410,N_14081,N_14152);
nand U15411 (N_15411,N_14818,N_14608);
and U15412 (N_15412,N_14700,N_14243);
nor U15413 (N_15413,N_14613,N_14366);
xor U15414 (N_15414,N_14483,N_14068);
nor U15415 (N_15415,N_14373,N_14538);
nor U15416 (N_15416,N_14559,N_14380);
nand U15417 (N_15417,N_14148,N_14844);
and U15418 (N_15418,N_14865,N_14896);
xnor U15419 (N_15419,N_14916,N_14923);
nor U15420 (N_15420,N_14845,N_14590);
nand U15421 (N_15421,N_14069,N_14409);
xnor U15422 (N_15422,N_14489,N_14837);
or U15423 (N_15423,N_14534,N_14646);
or U15424 (N_15424,N_14226,N_14901);
nand U15425 (N_15425,N_14106,N_14492);
or U15426 (N_15426,N_14282,N_14775);
nand U15427 (N_15427,N_14306,N_14907);
or U15428 (N_15428,N_14856,N_14884);
nand U15429 (N_15429,N_14759,N_14285);
nand U15430 (N_15430,N_14019,N_14921);
nand U15431 (N_15431,N_14859,N_14733);
and U15432 (N_15432,N_14811,N_14669);
or U15433 (N_15433,N_14848,N_14626);
nor U15434 (N_15434,N_14488,N_14145);
and U15435 (N_15435,N_14891,N_14781);
nor U15436 (N_15436,N_14875,N_14045);
xor U15437 (N_15437,N_14597,N_14029);
xor U15438 (N_15438,N_14962,N_14749);
nand U15439 (N_15439,N_14721,N_14417);
nand U15440 (N_15440,N_14393,N_14878);
xnor U15441 (N_15441,N_14991,N_14746);
xnor U15442 (N_15442,N_14126,N_14728);
and U15443 (N_15443,N_14984,N_14350);
xor U15444 (N_15444,N_14612,N_14562);
and U15445 (N_15445,N_14638,N_14246);
nand U15446 (N_15446,N_14619,N_14135);
or U15447 (N_15447,N_14659,N_14575);
xnor U15448 (N_15448,N_14771,N_14548);
nand U15449 (N_15449,N_14861,N_14168);
xnor U15450 (N_15450,N_14437,N_14541);
nor U15451 (N_15451,N_14586,N_14755);
or U15452 (N_15452,N_14319,N_14477);
nand U15453 (N_15453,N_14098,N_14677);
xnor U15454 (N_15454,N_14401,N_14042);
xnor U15455 (N_15455,N_14463,N_14178);
or U15456 (N_15456,N_14824,N_14186);
and U15457 (N_15457,N_14701,N_14205);
nand U15458 (N_15458,N_14297,N_14807);
nor U15459 (N_15459,N_14992,N_14585);
xnor U15460 (N_15460,N_14599,N_14418);
and U15461 (N_15461,N_14801,N_14340);
or U15462 (N_15462,N_14493,N_14196);
and U15463 (N_15463,N_14334,N_14447);
or U15464 (N_15464,N_14502,N_14473);
xor U15465 (N_15465,N_14935,N_14758);
xor U15466 (N_15466,N_14268,N_14736);
xnor U15467 (N_15467,N_14219,N_14747);
nor U15468 (N_15468,N_14505,N_14966);
nor U15469 (N_15469,N_14730,N_14840);
or U15470 (N_15470,N_14354,N_14621);
and U15471 (N_15471,N_14079,N_14117);
xnor U15472 (N_15472,N_14364,N_14355);
nand U15473 (N_15473,N_14977,N_14278);
or U15474 (N_15474,N_14524,N_14928);
xor U15475 (N_15475,N_14141,N_14331);
nand U15476 (N_15476,N_14565,N_14605);
nand U15477 (N_15477,N_14828,N_14989);
xor U15478 (N_15478,N_14577,N_14903);
nor U15479 (N_15479,N_14797,N_14679);
and U15480 (N_15480,N_14661,N_14812);
and U15481 (N_15481,N_14288,N_14255);
and U15482 (N_15482,N_14883,N_14778);
and U15483 (N_15483,N_14748,N_14228);
or U15484 (N_15484,N_14201,N_14842);
and U15485 (N_15485,N_14741,N_14335);
nand U15486 (N_15486,N_14829,N_14617);
nand U15487 (N_15487,N_14438,N_14479);
and U15488 (N_15488,N_14116,N_14578);
and U15489 (N_15489,N_14419,N_14583);
or U15490 (N_15490,N_14480,N_14353);
and U15491 (N_15491,N_14269,N_14738);
nand U15492 (N_15492,N_14817,N_14475);
nand U15493 (N_15493,N_14902,N_14932);
and U15494 (N_15494,N_14096,N_14714);
xor U15495 (N_15495,N_14752,N_14645);
nor U15496 (N_15496,N_14767,N_14846);
nand U15497 (N_15497,N_14286,N_14769);
or U15498 (N_15498,N_14239,N_14404);
nand U15499 (N_15499,N_14641,N_14200);
nor U15500 (N_15500,N_14778,N_14644);
and U15501 (N_15501,N_14883,N_14740);
nand U15502 (N_15502,N_14181,N_14236);
xor U15503 (N_15503,N_14378,N_14175);
nor U15504 (N_15504,N_14193,N_14861);
and U15505 (N_15505,N_14170,N_14875);
and U15506 (N_15506,N_14592,N_14768);
nand U15507 (N_15507,N_14214,N_14507);
nand U15508 (N_15508,N_14720,N_14821);
xor U15509 (N_15509,N_14839,N_14590);
or U15510 (N_15510,N_14613,N_14618);
nand U15511 (N_15511,N_14101,N_14057);
or U15512 (N_15512,N_14315,N_14227);
xor U15513 (N_15513,N_14210,N_14498);
xnor U15514 (N_15514,N_14428,N_14289);
and U15515 (N_15515,N_14615,N_14630);
or U15516 (N_15516,N_14032,N_14776);
nor U15517 (N_15517,N_14554,N_14363);
nor U15518 (N_15518,N_14393,N_14615);
or U15519 (N_15519,N_14046,N_14641);
and U15520 (N_15520,N_14040,N_14604);
xnor U15521 (N_15521,N_14640,N_14185);
and U15522 (N_15522,N_14293,N_14853);
nand U15523 (N_15523,N_14188,N_14762);
xor U15524 (N_15524,N_14200,N_14805);
and U15525 (N_15525,N_14380,N_14370);
and U15526 (N_15526,N_14482,N_14089);
or U15527 (N_15527,N_14383,N_14877);
nand U15528 (N_15528,N_14351,N_14770);
xnor U15529 (N_15529,N_14855,N_14561);
and U15530 (N_15530,N_14827,N_14213);
nor U15531 (N_15531,N_14609,N_14780);
nand U15532 (N_15532,N_14618,N_14814);
nor U15533 (N_15533,N_14784,N_14216);
or U15534 (N_15534,N_14371,N_14540);
or U15535 (N_15535,N_14154,N_14416);
or U15536 (N_15536,N_14720,N_14488);
and U15537 (N_15537,N_14227,N_14222);
and U15538 (N_15538,N_14924,N_14660);
xnor U15539 (N_15539,N_14165,N_14302);
nor U15540 (N_15540,N_14152,N_14317);
or U15541 (N_15541,N_14699,N_14148);
and U15542 (N_15542,N_14625,N_14390);
nand U15543 (N_15543,N_14346,N_14164);
nand U15544 (N_15544,N_14072,N_14592);
and U15545 (N_15545,N_14799,N_14757);
or U15546 (N_15546,N_14499,N_14116);
and U15547 (N_15547,N_14550,N_14515);
nor U15548 (N_15548,N_14260,N_14707);
and U15549 (N_15549,N_14699,N_14645);
or U15550 (N_15550,N_14864,N_14267);
and U15551 (N_15551,N_14226,N_14805);
nand U15552 (N_15552,N_14912,N_14398);
nand U15553 (N_15553,N_14715,N_14579);
nor U15554 (N_15554,N_14341,N_14525);
nand U15555 (N_15555,N_14529,N_14864);
xnor U15556 (N_15556,N_14388,N_14855);
nand U15557 (N_15557,N_14493,N_14117);
xnor U15558 (N_15558,N_14103,N_14208);
nand U15559 (N_15559,N_14567,N_14680);
nand U15560 (N_15560,N_14520,N_14098);
xor U15561 (N_15561,N_14769,N_14855);
xor U15562 (N_15562,N_14078,N_14643);
xor U15563 (N_15563,N_14314,N_14377);
xor U15564 (N_15564,N_14128,N_14186);
nor U15565 (N_15565,N_14222,N_14113);
xor U15566 (N_15566,N_14298,N_14912);
nand U15567 (N_15567,N_14444,N_14260);
or U15568 (N_15568,N_14431,N_14608);
or U15569 (N_15569,N_14020,N_14118);
nor U15570 (N_15570,N_14276,N_14324);
nand U15571 (N_15571,N_14960,N_14866);
or U15572 (N_15572,N_14339,N_14931);
nand U15573 (N_15573,N_14895,N_14940);
nor U15574 (N_15574,N_14220,N_14107);
or U15575 (N_15575,N_14803,N_14738);
nor U15576 (N_15576,N_14153,N_14460);
nor U15577 (N_15577,N_14394,N_14701);
xor U15578 (N_15578,N_14529,N_14646);
or U15579 (N_15579,N_14143,N_14176);
nand U15580 (N_15580,N_14945,N_14096);
or U15581 (N_15581,N_14881,N_14964);
xor U15582 (N_15582,N_14901,N_14194);
nand U15583 (N_15583,N_14064,N_14229);
xor U15584 (N_15584,N_14212,N_14518);
nor U15585 (N_15585,N_14186,N_14358);
nor U15586 (N_15586,N_14057,N_14147);
nand U15587 (N_15587,N_14613,N_14507);
xnor U15588 (N_15588,N_14785,N_14238);
nor U15589 (N_15589,N_14618,N_14792);
or U15590 (N_15590,N_14516,N_14960);
nor U15591 (N_15591,N_14164,N_14320);
or U15592 (N_15592,N_14493,N_14237);
xnor U15593 (N_15593,N_14739,N_14068);
or U15594 (N_15594,N_14782,N_14883);
nor U15595 (N_15595,N_14913,N_14230);
or U15596 (N_15596,N_14983,N_14031);
nand U15597 (N_15597,N_14923,N_14392);
and U15598 (N_15598,N_14434,N_14397);
and U15599 (N_15599,N_14563,N_14871);
xor U15600 (N_15600,N_14941,N_14662);
nor U15601 (N_15601,N_14874,N_14614);
nand U15602 (N_15602,N_14155,N_14367);
xnor U15603 (N_15603,N_14897,N_14880);
nor U15604 (N_15604,N_14407,N_14015);
xor U15605 (N_15605,N_14836,N_14994);
xor U15606 (N_15606,N_14326,N_14517);
xor U15607 (N_15607,N_14356,N_14674);
nor U15608 (N_15608,N_14127,N_14271);
nor U15609 (N_15609,N_14112,N_14055);
nor U15610 (N_15610,N_14795,N_14493);
and U15611 (N_15611,N_14373,N_14371);
or U15612 (N_15612,N_14222,N_14914);
or U15613 (N_15613,N_14614,N_14505);
and U15614 (N_15614,N_14856,N_14628);
nor U15615 (N_15615,N_14775,N_14468);
and U15616 (N_15616,N_14900,N_14999);
xnor U15617 (N_15617,N_14895,N_14928);
nor U15618 (N_15618,N_14097,N_14035);
or U15619 (N_15619,N_14864,N_14408);
nand U15620 (N_15620,N_14552,N_14899);
or U15621 (N_15621,N_14609,N_14452);
nor U15622 (N_15622,N_14906,N_14309);
nor U15623 (N_15623,N_14720,N_14049);
or U15624 (N_15624,N_14359,N_14532);
xor U15625 (N_15625,N_14224,N_14679);
nand U15626 (N_15626,N_14633,N_14353);
nor U15627 (N_15627,N_14657,N_14648);
or U15628 (N_15628,N_14364,N_14140);
nand U15629 (N_15629,N_14540,N_14911);
xnor U15630 (N_15630,N_14698,N_14149);
xor U15631 (N_15631,N_14177,N_14743);
nor U15632 (N_15632,N_14072,N_14116);
or U15633 (N_15633,N_14180,N_14617);
xor U15634 (N_15634,N_14404,N_14920);
nor U15635 (N_15635,N_14297,N_14438);
xor U15636 (N_15636,N_14236,N_14834);
nand U15637 (N_15637,N_14717,N_14527);
or U15638 (N_15638,N_14989,N_14933);
and U15639 (N_15639,N_14319,N_14549);
xnor U15640 (N_15640,N_14054,N_14687);
or U15641 (N_15641,N_14144,N_14108);
and U15642 (N_15642,N_14395,N_14065);
and U15643 (N_15643,N_14989,N_14231);
nand U15644 (N_15644,N_14855,N_14849);
nand U15645 (N_15645,N_14195,N_14634);
xnor U15646 (N_15646,N_14877,N_14502);
and U15647 (N_15647,N_14579,N_14079);
xor U15648 (N_15648,N_14405,N_14029);
xor U15649 (N_15649,N_14333,N_14386);
xor U15650 (N_15650,N_14395,N_14978);
xnor U15651 (N_15651,N_14576,N_14482);
xor U15652 (N_15652,N_14896,N_14693);
nor U15653 (N_15653,N_14920,N_14728);
or U15654 (N_15654,N_14028,N_14138);
xnor U15655 (N_15655,N_14828,N_14478);
nand U15656 (N_15656,N_14447,N_14252);
nand U15657 (N_15657,N_14282,N_14409);
nand U15658 (N_15658,N_14225,N_14644);
or U15659 (N_15659,N_14065,N_14110);
nand U15660 (N_15660,N_14885,N_14458);
and U15661 (N_15661,N_14260,N_14031);
and U15662 (N_15662,N_14179,N_14094);
nand U15663 (N_15663,N_14756,N_14007);
or U15664 (N_15664,N_14777,N_14082);
xor U15665 (N_15665,N_14264,N_14876);
nor U15666 (N_15666,N_14023,N_14867);
or U15667 (N_15667,N_14511,N_14009);
xor U15668 (N_15668,N_14812,N_14616);
nor U15669 (N_15669,N_14126,N_14611);
and U15670 (N_15670,N_14938,N_14003);
nor U15671 (N_15671,N_14949,N_14169);
and U15672 (N_15672,N_14982,N_14584);
nand U15673 (N_15673,N_14066,N_14926);
nand U15674 (N_15674,N_14388,N_14416);
and U15675 (N_15675,N_14588,N_14060);
nand U15676 (N_15676,N_14650,N_14795);
nand U15677 (N_15677,N_14552,N_14378);
xor U15678 (N_15678,N_14002,N_14622);
or U15679 (N_15679,N_14505,N_14399);
and U15680 (N_15680,N_14114,N_14094);
nand U15681 (N_15681,N_14219,N_14985);
nand U15682 (N_15682,N_14405,N_14194);
nand U15683 (N_15683,N_14546,N_14126);
nand U15684 (N_15684,N_14553,N_14760);
xor U15685 (N_15685,N_14254,N_14991);
nand U15686 (N_15686,N_14745,N_14989);
and U15687 (N_15687,N_14386,N_14786);
nand U15688 (N_15688,N_14552,N_14951);
and U15689 (N_15689,N_14453,N_14118);
or U15690 (N_15690,N_14689,N_14312);
or U15691 (N_15691,N_14522,N_14708);
xor U15692 (N_15692,N_14977,N_14264);
xnor U15693 (N_15693,N_14876,N_14525);
nand U15694 (N_15694,N_14717,N_14830);
nand U15695 (N_15695,N_14096,N_14731);
and U15696 (N_15696,N_14067,N_14879);
nand U15697 (N_15697,N_14160,N_14801);
nor U15698 (N_15698,N_14714,N_14970);
or U15699 (N_15699,N_14683,N_14126);
nand U15700 (N_15700,N_14664,N_14875);
nor U15701 (N_15701,N_14194,N_14195);
nor U15702 (N_15702,N_14823,N_14088);
and U15703 (N_15703,N_14729,N_14536);
nand U15704 (N_15704,N_14896,N_14036);
xor U15705 (N_15705,N_14496,N_14097);
nand U15706 (N_15706,N_14434,N_14972);
and U15707 (N_15707,N_14020,N_14880);
and U15708 (N_15708,N_14910,N_14802);
or U15709 (N_15709,N_14310,N_14930);
nor U15710 (N_15710,N_14797,N_14469);
and U15711 (N_15711,N_14419,N_14280);
and U15712 (N_15712,N_14839,N_14842);
nand U15713 (N_15713,N_14105,N_14729);
nor U15714 (N_15714,N_14044,N_14333);
xor U15715 (N_15715,N_14207,N_14284);
xnor U15716 (N_15716,N_14765,N_14801);
nor U15717 (N_15717,N_14744,N_14092);
nor U15718 (N_15718,N_14020,N_14280);
nor U15719 (N_15719,N_14170,N_14308);
and U15720 (N_15720,N_14768,N_14029);
or U15721 (N_15721,N_14410,N_14826);
and U15722 (N_15722,N_14734,N_14923);
nor U15723 (N_15723,N_14431,N_14263);
or U15724 (N_15724,N_14157,N_14863);
and U15725 (N_15725,N_14186,N_14442);
nor U15726 (N_15726,N_14315,N_14996);
and U15727 (N_15727,N_14925,N_14721);
nand U15728 (N_15728,N_14317,N_14453);
xor U15729 (N_15729,N_14019,N_14731);
xor U15730 (N_15730,N_14887,N_14557);
and U15731 (N_15731,N_14970,N_14941);
nand U15732 (N_15732,N_14788,N_14464);
xnor U15733 (N_15733,N_14831,N_14789);
and U15734 (N_15734,N_14480,N_14879);
or U15735 (N_15735,N_14567,N_14802);
nor U15736 (N_15736,N_14010,N_14282);
or U15737 (N_15737,N_14369,N_14065);
nor U15738 (N_15738,N_14890,N_14375);
or U15739 (N_15739,N_14324,N_14390);
and U15740 (N_15740,N_14522,N_14547);
and U15741 (N_15741,N_14506,N_14725);
and U15742 (N_15742,N_14997,N_14412);
nor U15743 (N_15743,N_14360,N_14267);
xor U15744 (N_15744,N_14975,N_14128);
nor U15745 (N_15745,N_14950,N_14538);
nor U15746 (N_15746,N_14214,N_14553);
nor U15747 (N_15747,N_14077,N_14997);
or U15748 (N_15748,N_14100,N_14307);
nor U15749 (N_15749,N_14182,N_14481);
or U15750 (N_15750,N_14054,N_14740);
nand U15751 (N_15751,N_14623,N_14780);
nand U15752 (N_15752,N_14551,N_14348);
xor U15753 (N_15753,N_14063,N_14821);
or U15754 (N_15754,N_14599,N_14385);
or U15755 (N_15755,N_14998,N_14039);
xor U15756 (N_15756,N_14718,N_14272);
and U15757 (N_15757,N_14197,N_14981);
nor U15758 (N_15758,N_14028,N_14236);
xnor U15759 (N_15759,N_14794,N_14979);
and U15760 (N_15760,N_14353,N_14334);
nand U15761 (N_15761,N_14262,N_14126);
xnor U15762 (N_15762,N_14230,N_14587);
and U15763 (N_15763,N_14075,N_14415);
nor U15764 (N_15764,N_14746,N_14382);
nor U15765 (N_15765,N_14451,N_14193);
nand U15766 (N_15766,N_14631,N_14064);
and U15767 (N_15767,N_14627,N_14075);
xnor U15768 (N_15768,N_14347,N_14390);
nor U15769 (N_15769,N_14725,N_14710);
nand U15770 (N_15770,N_14794,N_14364);
or U15771 (N_15771,N_14771,N_14115);
nand U15772 (N_15772,N_14857,N_14725);
xor U15773 (N_15773,N_14231,N_14248);
xor U15774 (N_15774,N_14427,N_14223);
xor U15775 (N_15775,N_14433,N_14205);
nor U15776 (N_15776,N_14332,N_14399);
nor U15777 (N_15777,N_14993,N_14528);
or U15778 (N_15778,N_14187,N_14365);
nand U15779 (N_15779,N_14091,N_14977);
nand U15780 (N_15780,N_14230,N_14274);
nand U15781 (N_15781,N_14315,N_14124);
or U15782 (N_15782,N_14413,N_14611);
nand U15783 (N_15783,N_14205,N_14216);
nor U15784 (N_15784,N_14417,N_14439);
and U15785 (N_15785,N_14754,N_14933);
nor U15786 (N_15786,N_14081,N_14778);
xor U15787 (N_15787,N_14493,N_14299);
nand U15788 (N_15788,N_14958,N_14779);
or U15789 (N_15789,N_14009,N_14883);
nand U15790 (N_15790,N_14279,N_14544);
and U15791 (N_15791,N_14691,N_14934);
nand U15792 (N_15792,N_14247,N_14447);
or U15793 (N_15793,N_14154,N_14089);
xor U15794 (N_15794,N_14996,N_14474);
or U15795 (N_15795,N_14567,N_14954);
nand U15796 (N_15796,N_14955,N_14996);
nand U15797 (N_15797,N_14678,N_14506);
nand U15798 (N_15798,N_14819,N_14667);
xnor U15799 (N_15799,N_14003,N_14522);
nand U15800 (N_15800,N_14216,N_14298);
xnor U15801 (N_15801,N_14338,N_14887);
xor U15802 (N_15802,N_14424,N_14958);
and U15803 (N_15803,N_14732,N_14643);
and U15804 (N_15804,N_14229,N_14953);
and U15805 (N_15805,N_14084,N_14262);
and U15806 (N_15806,N_14302,N_14689);
or U15807 (N_15807,N_14181,N_14439);
nand U15808 (N_15808,N_14016,N_14832);
and U15809 (N_15809,N_14613,N_14553);
or U15810 (N_15810,N_14098,N_14058);
nand U15811 (N_15811,N_14985,N_14111);
or U15812 (N_15812,N_14348,N_14414);
nand U15813 (N_15813,N_14349,N_14649);
xnor U15814 (N_15814,N_14422,N_14316);
nor U15815 (N_15815,N_14049,N_14339);
nand U15816 (N_15816,N_14948,N_14731);
nand U15817 (N_15817,N_14442,N_14321);
nor U15818 (N_15818,N_14886,N_14831);
nand U15819 (N_15819,N_14015,N_14696);
or U15820 (N_15820,N_14689,N_14126);
xnor U15821 (N_15821,N_14919,N_14668);
and U15822 (N_15822,N_14808,N_14779);
xnor U15823 (N_15823,N_14869,N_14913);
and U15824 (N_15824,N_14456,N_14638);
nor U15825 (N_15825,N_14481,N_14857);
and U15826 (N_15826,N_14003,N_14898);
nand U15827 (N_15827,N_14109,N_14659);
nand U15828 (N_15828,N_14996,N_14581);
or U15829 (N_15829,N_14940,N_14388);
or U15830 (N_15830,N_14487,N_14135);
xor U15831 (N_15831,N_14602,N_14003);
nand U15832 (N_15832,N_14367,N_14216);
xnor U15833 (N_15833,N_14207,N_14062);
nand U15834 (N_15834,N_14373,N_14055);
or U15835 (N_15835,N_14531,N_14603);
xor U15836 (N_15836,N_14112,N_14785);
or U15837 (N_15837,N_14420,N_14410);
xor U15838 (N_15838,N_14943,N_14789);
nor U15839 (N_15839,N_14760,N_14010);
nand U15840 (N_15840,N_14990,N_14754);
xnor U15841 (N_15841,N_14424,N_14749);
xor U15842 (N_15842,N_14278,N_14961);
or U15843 (N_15843,N_14531,N_14113);
nand U15844 (N_15844,N_14791,N_14373);
xnor U15845 (N_15845,N_14991,N_14864);
nor U15846 (N_15846,N_14192,N_14849);
or U15847 (N_15847,N_14582,N_14470);
nand U15848 (N_15848,N_14219,N_14355);
and U15849 (N_15849,N_14285,N_14387);
nand U15850 (N_15850,N_14651,N_14003);
and U15851 (N_15851,N_14306,N_14287);
nor U15852 (N_15852,N_14759,N_14284);
or U15853 (N_15853,N_14910,N_14851);
and U15854 (N_15854,N_14423,N_14881);
nand U15855 (N_15855,N_14052,N_14999);
nor U15856 (N_15856,N_14369,N_14591);
or U15857 (N_15857,N_14757,N_14455);
and U15858 (N_15858,N_14050,N_14675);
or U15859 (N_15859,N_14193,N_14626);
nor U15860 (N_15860,N_14858,N_14550);
nor U15861 (N_15861,N_14355,N_14974);
nor U15862 (N_15862,N_14171,N_14839);
xor U15863 (N_15863,N_14496,N_14233);
and U15864 (N_15864,N_14061,N_14226);
or U15865 (N_15865,N_14092,N_14585);
nor U15866 (N_15866,N_14474,N_14542);
xnor U15867 (N_15867,N_14110,N_14194);
nor U15868 (N_15868,N_14627,N_14086);
or U15869 (N_15869,N_14954,N_14841);
nand U15870 (N_15870,N_14514,N_14819);
or U15871 (N_15871,N_14749,N_14943);
and U15872 (N_15872,N_14229,N_14469);
or U15873 (N_15873,N_14182,N_14397);
nor U15874 (N_15874,N_14699,N_14858);
and U15875 (N_15875,N_14747,N_14048);
xor U15876 (N_15876,N_14891,N_14004);
nor U15877 (N_15877,N_14417,N_14223);
nand U15878 (N_15878,N_14303,N_14916);
xor U15879 (N_15879,N_14497,N_14746);
or U15880 (N_15880,N_14720,N_14615);
nor U15881 (N_15881,N_14690,N_14632);
nor U15882 (N_15882,N_14098,N_14891);
nor U15883 (N_15883,N_14928,N_14393);
and U15884 (N_15884,N_14214,N_14248);
and U15885 (N_15885,N_14333,N_14117);
and U15886 (N_15886,N_14585,N_14877);
nor U15887 (N_15887,N_14811,N_14234);
and U15888 (N_15888,N_14202,N_14011);
or U15889 (N_15889,N_14800,N_14880);
xor U15890 (N_15890,N_14713,N_14734);
nor U15891 (N_15891,N_14333,N_14981);
xor U15892 (N_15892,N_14884,N_14237);
or U15893 (N_15893,N_14765,N_14550);
nand U15894 (N_15894,N_14889,N_14686);
xnor U15895 (N_15895,N_14021,N_14204);
nor U15896 (N_15896,N_14506,N_14051);
and U15897 (N_15897,N_14121,N_14266);
nand U15898 (N_15898,N_14083,N_14474);
and U15899 (N_15899,N_14458,N_14913);
and U15900 (N_15900,N_14636,N_14470);
nand U15901 (N_15901,N_14983,N_14155);
or U15902 (N_15902,N_14679,N_14568);
nor U15903 (N_15903,N_14507,N_14259);
nand U15904 (N_15904,N_14095,N_14789);
and U15905 (N_15905,N_14003,N_14074);
xor U15906 (N_15906,N_14683,N_14649);
or U15907 (N_15907,N_14859,N_14946);
or U15908 (N_15908,N_14629,N_14533);
xor U15909 (N_15909,N_14815,N_14909);
nand U15910 (N_15910,N_14212,N_14308);
and U15911 (N_15911,N_14864,N_14229);
and U15912 (N_15912,N_14548,N_14112);
or U15913 (N_15913,N_14651,N_14524);
or U15914 (N_15914,N_14331,N_14675);
nor U15915 (N_15915,N_14467,N_14602);
nand U15916 (N_15916,N_14414,N_14718);
nor U15917 (N_15917,N_14642,N_14381);
nand U15918 (N_15918,N_14817,N_14119);
nand U15919 (N_15919,N_14546,N_14858);
or U15920 (N_15920,N_14209,N_14233);
xnor U15921 (N_15921,N_14484,N_14903);
xor U15922 (N_15922,N_14569,N_14306);
xnor U15923 (N_15923,N_14431,N_14356);
or U15924 (N_15924,N_14345,N_14303);
xor U15925 (N_15925,N_14780,N_14983);
or U15926 (N_15926,N_14165,N_14693);
xnor U15927 (N_15927,N_14303,N_14302);
and U15928 (N_15928,N_14818,N_14893);
and U15929 (N_15929,N_14347,N_14571);
xnor U15930 (N_15930,N_14188,N_14039);
nand U15931 (N_15931,N_14087,N_14192);
nor U15932 (N_15932,N_14211,N_14387);
nor U15933 (N_15933,N_14064,N_14533);
xnor U15934 (N_15934,N_14089,N_14454);
or U15935 (N_15935,N_14726,N_14981);
nor U15936 (N_15936,N_14229,N_14014);
nor U15937 (N_15937,N_14512,N_14503);
nor U15938 (N_15938,N_14485,N_14335);
xnor U15939 (N_15939,N_14286,N_14573);
xor U15940 (N_15940,N_14424,N_14210);
xor U15941 (N_15941,N_14987,N_14228);
and U15942 (N_15942,N_14836,N_14723);
nand U15943 (N_15943,N_14666,N_14457);
nand U15944 (N_15944,N_14914,N_14800);
xnor U15945 (N_15945,N_14325,N_14091);
or U15946 (N_15946,N_14518,N_14126);
or U15947 (N_15947,N_14962,N_14926);
or U15948 (N_15948,N_14481,N_14648);
xnor U15949 (N_15949,N_14827,N_14269);
nor U15950 (N_15950,N_14421,N_14265);
nand U15951 (N_15951,N_14422,N_14596);
nand U15952 (N_15952,N_14348,N_14619);
nor U15953 (N_15953,N_14812,N_14647);
nor U15954 (N_15954,N_14706,N_14335);
and U15955 (N_15955,N_14058,N_14723);
or U15956 (N_15956,N_14325,N_14797);
nor U15957 (N_15957,N_14409,N_14004);
or U15958 (N_15958,N_14279,N_14277);
and U15959 (N_15959,N_14729,N_14111);
nand U15960 (N_15960,N_14217,N_14106);
and U15961 (N_15961,N_14226,N_14245);
and U15962 (N_15962,N_14452,N_14142);
xor U15963 (N_15963,N_14856,N_14724);
and U15964 (N_15964,N_14414,N_14477);
or U15965 (N_15965,N_14380,N_14303);
xor U15966 (N_15966,N_14095,N_14204);
nor U15967 (N_15967,N_14364,N_14593);
and U15968 (N_15968,N_14069,N_14907);
nor U15969 (N_15969,N_14098,N_14663);
and U15970 (N_15970,N_14240,N_14640);
xor U15971 (N_15971,N_14709,N_14600);
or U15972 (N_15972,N_14512,N_14855);
or U15973 (N_15973,N_14704,N_14877);
and U15974 (N_15974,N_14094,N_14801);
xor U15975 (N_15975,N_14433,N_14561);
and U15976 (N_15976,N_14692,N_14295);
xor U15977 (N_15977,N_14608,N_14981);
nor U15978 (N_15978,N_14929,N_14462);
and U15979 (N_15979,N_14786,N_14044);
or U15980 (N_15980,N_14322,N_14615);
xor U15981 (N_15981,N_14718,N_14646);
nor U15982 (N_15982,N_14698,N_14280);
xor U15983 (N_15983,N_14560,N_14470);
nand U15984 (N_15984,N_14238,N_14617);
xor U15985 (N_15985,N_14305,N_14676);
nor U15986 (N_15986,N_14173,N_14915);
nand U15987 (N_15987,N_14088,N_14618);
xor U15988 (N_15988,N_14363,N_14641);
xnor U15989 (N_15989,N_14457,N_14669);
xnor U15990 (N_15990,N_14759,N_14057);
nor U15991 (N_15991,N_14663,N_14434);
or U15992 (N_15992,N_14824,N_14161);
and U15993 (N_15993,N_14494,N_14793);
nor U15994 (N_15994,N_14413,N_14696);
or U15995 (N_15995,N_14771,N_14267);
nor U15996 (N_15996,N_14283,N_14993);
and U15997 (N_15997,N_14598,N_14216);
nand U15998 (N_15998,N_14080,N_14012);
xor U15999 (N_15999,N_14297,N_14792);
nor U16000 (N_16000,N_15773,N_15948);
nor U16001 (N_16001,N_15081,N_15157);
nor U16002 (N_16002,N_15949,N_15801);
nor U16003 (N_16003,N_15928,N_15431);
nor U16004 (N_16004,N_15419,N_15849);
nor U16005 (N_16005,N_15272,N_15936);
nor U16006 (N_16006,N_15069,N_15664);
nand U16007 (N_16007,N_15511,N_15221);
xor U16008 (N_16008,N_15981,N_15053);
nand U16009 (N_16009,N_15754,N_15034);
or U16010 (N_16010,N_15497,N_15422);
or U16011 (N_16011,N_15152,N_15790);
nor U16012 (N_16012,N_15972,N_15971);
or U16013 (N_16013,N_15847,N_15522);
and U16014 (N_16014,N_15499,N_15114);
nor U16015 (N_16015,N_15516,N_15892);
and U16016 (N_16016,N_15534,N_15456);
or U16017 (N_16017,N_15430,N_15220);
nor U16018 (N_16018,N_15125,N_15150);
and U16019 (N_16019,N_15250,N_15357);
or U16020 (N_16020,N_15418,N_15760);
nor U16021 (N_16021,N_15787,N_15297);
nand U16022 (N_16022,N_15656,N_15321);
nor U16023 (N_16023,N_15313,N_15446);
nor U16024 (N_16024,N_15324,N_15919);
and U16025 (N_16025,N_15479,N_15194);
or U16026 (N_16026,N_15959,N_15421);
nor U16027 (N_16027,N_15043,N_15925);
and U16028 (N_16028,N_15756,N_15211);
or U16029 (N_16029,N_15531,N_15976);
nor U16030 (N_16030,N_15005,N_15672);
or U16031 (N_16031,N_15681,N_15917);
xnor U16032 (N_16032,N_15415,N_15292);
and U16033 (N_16033,N_15208,N_15484);
xnor U16034 (N_16034,N_15859,N_15390);
nand U16035 (N_16035,N_15876,N_15374);
or U16036 (N_16036,N_15101,N_15771);
xnor U16037 (N_16037,N_15269,N_15662);
xor U16038 (N_16038,N_15035,N_15602);
and U16039 (N_16039,N_15804,N_15119);
and U16040 (N_16040,N_15874,N_15857);
and U16041 (N_16041,N_15481,N_15079);
and U16042 (N_16042,N_15493,N_15837);
nand U16043 (N_16043,N_15059,N_15477);
and U16044 (N_16044,N_15625,N_15312);
and U16045 (N_16045,N_15398,N_15004);
nor U16046 (N_16046,N_15524,N_15102);
and U16047 (N_16047,N_15975,N_15750);
and U16048 (N_16048,N_15340,N_15433);
xnor U16049 (N_16049,N_15666,N_15451);
nor U16050 (N_16050,N_15749,N_15382);
or U16051 (N_16051,N_15647,N_15447);
or U16052 (N_16052,N_15748,N_15105);
nor U16053 (N_16053,N_15770,N_15118);
and U16054 (N_16054,N_15112,N_15160);
xor U16055 (N_16055,N_15448,N_15145);
nand U16056 (N_16056,N_15469,N_15097);
and U16057 (N_16057,N_15638,N_15411);
nand U16058 (N_16058,N_15805,N_15813);
and U16059 (N_16059,N_15260,N_15038);
xnor U16060 (N_16060,N_15015,N_15894);
or U16061 (N_16061,N_15768,N_15755);
or U16062 (N_16062,N_15690,N_15089);
nand U16063 (N_16063,N_15514,N_15995);
nand U16064 (N_16064,N_15199,N_15061);
nand U16065 (N_16065,N_15718,N_15802);
or U16066 (N_16066,N_15621,N_15765);
or U16067 (N_16067,N_15630,N_15589);
nand U16068 (N_16068,N_15439,N_15614);
nand U16069 (N_16069,N_15535,N_15597);
or U16070 (N_16070,N_15784,N_15624);
xor U16071 (N_16071,N_15449,N_15240);
and U16072 (N_16072,N_15007,N_15828);
nand U16073 (N_16073,N_15598,N_15686);
nand U16074 (N_16074,N_15018,N_15227);
xor U16075 (N_16075,N_15734,N_15796);
and U16076 (N_16076,N_15844,N_15402);
and U16077 (N_16077,N_15908,N_15682);
nor U16078 (N_16078,N_15716,N_15510);
or U16079 (N_16079,N_15291,N_15489);
nor U16080 (N_16080,N_15890,N_15351);
nand U16081 (N_16081,N_15488,N_15130);
nor U16082 (N_16082,N_15617,N_15338);
nor U16083 (N_16083,N_15190,N_15850);
xnor U16084 (N_16084,N_15654,N_15528);
nor U16085 (N_16085,N_15065,N_15234);
xor U16086 (N_16086,N_15370,N_15237);
nor U16087 (N_16087,N_15270,N_15769);
or U16088 (N_16088,N_15884,N_15349);
nand U16089 (N_16089,N_15717,N_15953);
and U16090 (N_16090,N_15891,N_15858);
nor U16091 (N_16091,N_15642,N_15905);
nor U16092 (N_16092,N_15336,N_15646);
xnor U16093 (N_16093,N_15281,N_15149);
and U16094 (N_16094,N_15914,N_15271);
and U16095 (N_16095,N_15473,N_15818);
nor U16096 (N_16096,N_15671,N_15546);
or U16097 (N_16097,N_15747,N_15583);
xnor U16098 (N_16098,N_15273,N_15095);
or U16099 (N_16099,N_15827,N_15315);
or U16100 (N_16100,N_15725,N_15994);
xnor U16101 (N_16101,N_15496,N_15968);
and U16102 (N_16102,N_15162,N_15545);
nand U16103 (N_16103,N_15608,N_15226);
or U16104 (N_16104,N_15577,N_15319);
xor U16105 (N_16105,N_15644,N_15204);
nor U16106 (N_16106,N_15244,N_15048);
xor U16107 (N_16107,N_15047,N_15029);
or U16108 (N_16108,N_15051,N_15856);
nand U16109 (N_16109,N_15861,N_15871);
or U16110 (N_16110,N_15955,N_15592);
or U16111 (N_16111,N_15251,N_15068);
xor U16112 (N_16112,N_15159,N_15509);
or U16113 (N_16113,N_15560,N_15816);
nand U16114 (N_16114,N_15322,N_15706);
nand U16115 (N_16115,N_15887,N_15763);
or U16116 (N_16116,N_15970,N_15262);
xnor U16117 (N_16117,N_15316,N_15628);
or U16118 (N_16118,N_15626,N_15793);
and U16119 (N_16119,N_15274,N_15361);
xnor U16120 (N_16120,N_15380,N_15229);
nor U16121 (N_16121,N_15989,N_15491);
nor U16122 (N_16122,N_15513,N_15703);
nand U16123 (N_16123,N_15569,N_15417);
nand U16124 (N_16124,N_15730,N_15457);
nor U16125 (N_16125,N_15026,N_15570);
and U16126 (N_16126,N_15426,N_15944);
and U16127 (N_16127,N_15487,N_15609);
nor U16128 (N_16128,N_15263,N_15868);
nand U16129 (N_16129,N_15788,N_15683);
and U16130 (N_16130,N_15475,N_15033);
nand U16131 (N_16131,N_15882,N_15201);
nand U16132 (N_16132,N_15169,N_15806);
or U16133 (N_16133,N_15259,N_15054);
or U16134 (N_16134,N_15261,N_15021);
nand U16135 (N_16135,N_15386,N_15287);
and U16136 (N_16136,N_15550,N_15083);
nand U16137 (N_16137,N_15979,N_15396);
nor U16138 (N_16138,N_15305,N_15500);
nand U16139 (N_16139,N_15337,N_15455);
xor U16140 (N_16140,N_15937,N_15285);
xor U16141 (N_16141,N_15778,N_15729);
nor U16142 (N_16142,N_15178,N_15333);
and U16143 (N_16143,N_15164,N_15721);
nand U16144 (N_16144,N_15699,N_15636);
and U16145 (N_16145,N_15603,N_15586);
nor U16146 (N_16146,N_15909,N_15923);
xnor U16147 (N_16147,N_15973,N_15620);
and U16148 (N_16148,N_15320,N_15854);
nand U16149 (N_16149,N_15853,N_15276);
and U16150 (N_16150,N_15358,N_15520);
xor U16151 (N_16151,N_15179,N_15895);
xnor U16152 (N_16152,N_15561,N_15512);
xnor U16153 (N_16153,N_15803,N_15031);
nor U16154 (N_16154,N_15687,N_15412);
and U16155 (N_16155,N_15978,N_15595);
or U16156 (N_16156,N_15371,N_15231);
xor U16157 (N_16157,N_15865,N_15384);
and U16158 (N_16158,N_15530,N_15565);
or U16159 (N_16159,N_15896,N_15040);
xor U16160 (N_16160,N_15282,N_15082);
nand U16161 (N_16161,N_15774,N_15132);
and U16162 (N_16162,N_15036,N_15326);
xnor U16163 (N_16163,N_15334,N_15606);
xor U16164 (N_16164,N_15407,N_15632);
nand U16165 (N_16165,N_15091,N_15506);
xnor U16166 (N_16166,N_15037,N_15677);
nor U16167 (N_16167,N_15266,N_15391);
xor U16168 (N_16168,N_15039,N_15177);
nand U16169 (N_16169,N_15104,N_15459);
or U16170 (N_16170,N_15810,N_15987);
or U16171 (N_16171,N_15071,N_15552);
or U16172 (N_16172,N_15373,N_15111);
xnor U16173 (N_16173,N_15184,N_15126);
nand U16174 (N_16174,N_15331,N_15916);
nor U16175 (N_16175,N_15317,N_15120);
xnor U16176 (N_16176,N_15964,N_15799);
xnor U16177 (N_16177,N_15924,N_15591);
xor U16178 (N_16178,N_15922,N_15008);
nor U16179 (N_16179,N_15265,N_15807);
xor U16180 (N_16180,N_15962,N_15992);
and U16181 (N_16181,N_15710,N_15127);
and U16182 (N_16182,N_15408,N_15328);
xnor U16183 (N_16183,N_15028,N_15056);
or U16184 (N_16184,N_15676,N_15575);
or U16185 (N_16185,N_15153,N_15872);
xnor U16186 (N_16186,N_15780,N_15186);
nand U16187 (N_16187,N_15820,N_15883);
or U16188 (N_16188,N_15329,N_15090);
nand U16189 (N_16189,N_15785,N_15860);
nor U16190 (N_16190,N_15367,N_15723);
xnor U16191 (N_16191,N_15840,N_15673);
and U16192 (N_16192,N_15692,N_15161);
or U16193 (N_16193,N_15501,N_15372);
or U16194 (N_16194,N_15131,N_15766);
nand U16195 (N_16195,N_15660,N_15143);
nor U16196 (N_16196,N_15888,N_15658);
and U16197 (N_16197,N_15067,N_15616);
and U16198 (N_16198,N_15913,N_15640);
xor U16199 (N_16199,N_15267,N_15022);
or U16200 (N_16200,N_15277,N_15852);
or U16201 (N_16201,N_15757,N_15578);
and U16202 (N_16202,N_15452,N_15353);
xor U16203 (N_16203,N_15425,N_15215);
nand U16204 (N_16204,N_15599,N_15834);
and U16205 (N_16205,N_15822,N_15956);
xnor U16206 (N_16206,N_15899,N_15257);
nor U16207 (N_16207,N_15783,N_15247);
nor U16208 (N_16208,N_15495,N_15232);
xnor U16209 (N_16209,N_15873,N_15841);
nand U16210 (N_16210,N_15189,N_15537);
xnor U16211 (N_16211,N_15492,N_15017);
xnor U16212 (N_16212,N_15898,N_15631);
nand U16213 (N_16213,N_15424,N_15302);
or U16214 (N_16214,N_15206,N_15318);
xor U16215 (N_16215,N_15241,N_15574);
or U16216 (N_16216,N_15951,N_15141);
nand U16217 (N_16217,N_15002,N_15738);
and U16218 (N_16218,N_15675,N_15003);
or U16219 (N_16219,N_15167,N_15669);
and U16220 (N_16220,N_15295,N_15746);
or U16221 (N_16221,N_15014,N_15001);
nor U16222 (N_16222,N_15490,N_15289);
or U16223 (N_16223,N_15420,N_15427);
or U16224 (N_16224,N_15202,N_15138);
or U16225 (N_16225,N_15436,N_15196);
or U16226 (N_16226,N_15121,N_15878);
nand U16227 (N_16227,N_15348,N_15084);
nor U16228 (N_16228,N_15180,N_15428);
nor U16229 (N_16229,N_15122,N_15693);
and U16230 (N_16230,N_15713,N_15158);
and U16231 (N_16231,N_15294,N_15668);
nor U16232 (N_16232,N_15323,N_15634);
or U16233 (N_16233,N_15182,N_15006);
nor U16234 (N_16234,N_15142,N_15238);
xnor U16235 (N_16235,N_15759,N_15044);
nor U16236 (N_16236,N_15996,N_15831);
nand U16237 (N_16237,N_15593,N_15696);
nor U16238 (N_16238,N_15183,N_15144);
nand U16239 (N_16239,N_15714,N_15657);
nor U16240 (N_16240,N_15041,N_15623);
xnor U16241 (N_16241,N_15864,N_15742);
or U16242 (N_16242,N_15405,N_15109);
and U16243 (N_16243,N_15555,N_15585);
and U16244 (N_16244,N_15982,N_15932);
nand U16245 (N_16245,N_15776,N_15210);
nand U16246 (N_16246,N_15988,N_15904);
nor U16247 (N_16247,N_15085,N_15659);
xor U16248 (N_16248,N_15532,N_15942);
nand U16249 (N_16249,N_15224,N_15508);
xor U16250 (N_16250,N_15846,N_15551);
and U16251 (N_16251,N_15918,N_15151);
nor U16252 (N_16252,N_15072,N_15191);
or U16253 (N_16253,N_15901,N_15579);
nand U16254 (N_16254,N_15377,N_15863);
nand U16255 (N_16255,N_15622,N_15503);
nor U16256 (N_16256,N_15376,N_15737);
and U16257 (N_16257,N_15306,N_15465);
xnor U16258 (N_16258,N_15910,N_15406);
and U16259 (N_16259,N_15965,N_15394);
and U16260 (N_16260,N_15688,N_15346);
nor U16261 (N_16261,N_15637,N_15576);
nor U16262 (N_16262,N_15464,N_15627);
or U16263 (N_16263,N_15443,N_15794);
xnor U16264 (N_16264,N_15526,N_15288);
or U16265 (N_16265,N_15678,N_15124);
nor U16266 (N_16266,N_15472,N_15413);
xnor U16267 (N_16267,N_15613,N_15077);
nand U16268 (N_16268,N_15379,N_15800);
nand U16269 (N_16269,N_15735,N_15934);
xor U16270 (N_16270,N_15906,N_15388);
and U16271 (N_16271,N_15325,N_15070);
xor U16272 (N_16272,N_15564,N_15870);
nand U16273 (N_16273,N_15304,N_15722);
or U16274 (N_16274,N_15467,N_15093);
xnor U16275 (N_16275,N_15092,N_15607);
nor U16276 (N_16276,N_15587,N_15568);
or U16277 (N_16277,N_15156,N_15782);
nand U16278 (N_16278,N_15155,N_15498);
nor U16279 (N_16279,N_15246,N_15571);
and U16280 (N_16280,N_15401,N_15764);
and U16281 (N_16281,N_15330,N_15521);
or U16282 (N_16282,N_15228,N_15042);
or U16283 (N_16283,N_15945,N_15057);
and U16284 (N_16284,N_15739,N_15661);
or U16285 (N_16285,N_15518,N_15911);
nor U16286 (N_16286,N_15848,N_15838);
nand U16287 (N_16287,N_15011,N_15543);
or U16288 (N_16288,N_15073,N_15612);
or U16289 (N_16289,N_15437,N_15539);
nand U16290 (N_16290,N_15680,N_15205);
nand U16291 (N_16291,N_15217,N_15605);
nand U16292 (N_16292,N_15248,N_15045);
or U16293 (N_16293,N_15663,N_15679);
xnor U16294 (N_16294,N_15429,N_15772);
xnor U16295 (N_16295,N_15767,N_15476);
nand U16296 (N_16296,N_15468,N_15298);
xor U16297 (N_16297,N_15581,N_15781);
and U16298 (N_16298,N_15080,N_15762);
and U16299 (N_16299,N_15610,N_15958);
and U16300 (N_16300,N_15470,N_15236);
or U16301 (N_16301,N_15824,N_15761);
and U16302 (N_16302,N_15980,N_15432);
and U16303 (N_16303,N_15943,N_15173);
nor U16304 (N_16304,N_15012,N_15548);
or U16305 (N_16305,N_15146,N_15135);
nand U16306 (N_16306,N_15286,N_15176);
nand U16307 (N_16307,N_15296,N_15235);
xnor U16308 (N_16308,N_15886,N_15381);
xor U16309 (N_16309,N_15024,N_15835);
and U16310 (N_16310,N_15066,N_15255);
or U16311 (N_16311,N_15639,N_15078);
and U16312 (N_16312,N_15946,N_15926);
and U16313 (N_16313,N_15998,N_15385);
and U16314 (N_16314,N_15087,N_15364);
nand U16315 (N_16315,N_15845,N_15483);
or U16316 (N_16316,N_15588,N_15020);
or U16317 (N_16317,N_15825,N_15650);
nor U16318 (N_16318,N_15219,N_15823);
nor U16319 (N_16319,N_15695,N_15795);
nor U16320 (N_16320,N_15655,N_15867);
and U16321 (N_16321,N_15740,N_15303);
nand U16322 (N_16322,N_15808,N_15618);
xnor U16323 (N_16323,N_15930,N_15016);
or U16324 (N_16324,N_15557,N_15137);
xnor U16325 (N_16325,N_15290,N_15258);
xor U16326 (N_16326,N_15615,N_15355);
or U16327 (N_16327,N_15821,N_15653);
nor U16328 (N_16328,N_15147,N_15731);
nor U16329 (N_16329,N_15529,N_15881);
nand U16330 (N_16330,N_15842,N_15486);
nor U16331 (N_16331,N_15103,N_15741);
or U16332 (N_16332,N_15517,N_15154);
nor U16333 (N_16333,N_15438,N_15967);
or U16334 (N_16334,N_15309,N_15549);
xor U16335 (N_16335,N_15921,N_15243);
nand U16336 (N_16336,N_15811,N_15544);
or U16337 (N_16337,N_15393,N_15984);
xnor U16338 (N_16338,N_15843,N_15839);
and U16339 (N_16339,N_15991,N_15245);
and U16340 (N_16340,N_15368,N_15814);
or U16341 (N_16341,N_15275,N_15563);
nor U16342 (N_16342,N_15900,N_15527);
xor U16343 (N_16343,N_15293,N_15708);
and U16344 (N_16344,N_15474,N_15175);
nor U16345 (N_16345,N_15139,N_15869);
nor U16346 (N_16346,N_15345,N_15299);
nor U16347 (N_16347,N_15086,N_15947);
nor U16348 (N_16348,N_15249,N_15013);
or U16349 (N_16349,N_15553,N_15547);
nand U16350 (N_16350,N_15099,N_15667);
nor U16351 (N_16351,N_15301,N_15985);
nor U16352 (N_16352,N_15050,N_15726);
nor U16353 (N_16353,N_15280,N_15117);
nor U16354 (N_16354,N_15986,N_15461);
nor U16355 (N_16355,N_15397,N_15728);
nand U16356 (N_16356,N_15974,N_15128);
or U16357 (N_16357,N_15075,N_15931);
and U16358 (N_16358,N_15573,N_15466);
nor U16359 (N_16359,N_15507,N_15709);
and U16360 (N_16360,N_15957,N_15233);
or U16361 (N_16361,N_15283,N_15171);
nand U16362 (N_16362,N_15594,N_15062);
nor U16363 (N_16363,N_15879,N_15440);
xnor U16364 (N_16364,N_15554,N_15567);
nand U16365 (N_16365,N_15812,N_15387);
or U16366 (N_16366,N_15343,N_15458);
xnor U16367 (N_16367,N_15023,N_15254);
xnor U16368 (N_16368,N_15363,N_15809);
xor U16369 (N_16369,N_15941,N_15880);
or U16370 (N_16370,N_15836,N_15797);
xnor U16371 (N_16371,N_15938,N_15025);
nand U16372 (N_16372,N_15933,N_15209);
nand U16373 (N_16373,N_15106,N_15792);
xor U16374 (N_16374,N_15369,N_15652);
or U16375 (N_16375,N_15665,N_15268);
nand U16376 (N_16376,N_15643,N_15030);
nor U16377 (N_16377,N_15445,N_15889);
or U16378 (N_16378,N_15253,N_15744);
and U16379 (N_16379,N_15826,N_15515);
xnor U16380 (N_16380,N_15108,N_15356);
nor U16381 (N_16381,N_15629,N_15903);
nand U16382 (N_16382,N_15195,N_15533);
or U16383 (N_16383,N_15935,N_15172);
nor U16384 (N_16384,N_15862,N_15076);
nor U16385 (N_16385,N_15218,N_15403);
nor U16386 (N_16386,N_15096,N_15743);
xnor U16387 (N_16387,N_15416,N_15187);
nand U16388 (N_16388,N_15284,N_15203);
xor U16389 (N_16389,N_15502,N_15851);
and U16390 (N_16390,N_15200,N_15929);
xor U16391 (N_16391,N_15359,N_15775);
nand U16392 (N_16392,N_15875,N_15453);
nor U16393 (N_16393,N_15727,N_15674);
nor U16394 (N_16394,N_15990,N_15758);
nor U16395 (N_16395,N_15999,N_15893);
nand U16396 (N_16396,N_15116,N_15378);
and U16397 (N_16397,N_15733,N_15752);
xor U16398 (N_16398,N_15684,N_15027);
nand U16399 (N_16399,N_15829,N_15940);
nor U16400 (N_16400,N_15482,N_15136);
nor U16401 (N_16401,N_15414,N_15327);
or U16402 (N_16402,N_15635,N_15389);
or U16403 (N_16403,N_15815,N_15966);
nor U16404 (N_16404,N_15392,N_15670);
and U16405 (N_16405,N_15166,N_15751);
nand U16406 (N_16406,N_15558,N_15601);
and U16407 (N_16407,N_15049,N_15832);
nand U16408 (N_16408,N_15129,N_15168);
nor U16409 (N_16409,N_15052,N_15736);
or U16410 (N_16410,N_15649,N_15395);
nand U16411 (N_16411,N_15480,N_15423);
nand U16412 (N_16412,N_15961,N_15633);
nor U16413 (N_16413,N_15110,N_15691);
xor U16414 (N_16414,N_15264,N_15952);
nor U16415 (N_16415,N_15559,N_15088);
and U16416 (N_16416,N_15897,N_15701);
nor U16417 (N_16417,N_15444,N_15977);
xor U16418 (N_16418,N_15566,N_15611);
or U16419 (N_16419,N_15174,N_15927);
xnor U16420 (N_16420,N_15115,N_15074);
and U16421 (N_16421,N_15055,N_15256);
and U16422 (N_16422,N_15460,N_15786);
nor U16423 (N_16423,N_15641,N_15833);
nand U16424 (N_16424,N_15185,N_15310);
nand U16425 (N_16425,N_15308,N_15198);
nand U16426 (N_16426,N_15541,N_15339);
or U16427 (N_16427,N_15058,N_15278);
nor U16428 (N_16428,N_15242,N_15645);
xor U16429 (N_16429,N_15584,N_15098);
nand U16430 (N_16430,N_15360,N_15197);
nor U16431 (N_16431,N_15170,N_15148);
and U16432 (N_16432,N_15877,N_15715);
and U16433 (N_16433,N_15193,N_15009);
and U16434 (N_16434,N_15997,N_15335);
nand U16435 (N_16435,N_15540,N_15463);
nand U16436 (N_16436,N_15332,N_15435);
nand U16437 (N_16437,N_15538,N_15399);
xnor U16438 (N_16438,N_15969,N_15700);
nand U16439 (N_16439,N_15347,N_15165);
xnor U16440 (N_16440,N_15352,N_15434);
nand U16441 (N_16441,N_15580,N_15819);
nand U16442 (N_16442,N_15983,N_15950);
xnor U16443 (N_16443,N_15712,N_15342);
and U16444 (N_16444,N_15107,N_15314);
xor U16445 (N_16445,N_15113,N_15100);
nand U16446 (N_16446,N_15753,N_15383);
or U16447 (N_16447,N_15019,N_15223);
xor U16448 (N_16448,N_15478,N_15885);
xnor U16449 (N_16449,N_15719,N_15400);
nor U16450 (N_16450,N_15365,N_15745);
or U16451 (N_16451,N_15212,N_15902);
or U16452 (N_16452,N_15562,N_15354);
xnor U16453 (N_16453,N_15404,N_15724);
nor U16454 (N_16454,N_15410,N_15707);
and U16455 (N_16455,N_15000,N_15960);
nand U16456 (N_16456,N_15344,N_15907);
xnor U16457 (N_16457,N_15720,N_15094);
nor U16458 (N_16458,N_15134,N_15462);
and U16459 (N_16459,N_15694,N_15866);
and U16460 (N_16460,N_15791,N_15525);
nor U16461 (N_16461,N_15519,N_15993);
or U16462 (N_16462,N_15123,N_15213);
and U16463 (N_16463,N_15064,N_15494);
nand U16464 (N_16464,N_15572,N_15582);
and U16465 (N_16465,N_15604,N_15920);
xnor U16466 (N_16466,N_15442,N_15192);
nand U16467 (N_16467,N_15505,N_15705);
nand U16468 (N_16468,N_15689,N_15341);
nor U16469 (N_16469,N_15225,N_15222);
nor U16470 (N_16470,N_15915,N_15450);
and U16471 (N_16471,N_15230,N_15855);
and U16472 (N_16472,N_15711,N_15648);
xor U16473 (N_16473,N_15307,N_15697);
nand U16474 (N_16474,N_15536,N_15542);
xor U16475 (N_16475,N_15912,N_15600);
and U16476 (N_16476,N_15702,N_15216);
xnor U16477 (N_16477,N_15060,N_15596);
nand U16478 (N_16478,N_15732,N_15777);
nand U16479 (N_16479,N_15556,N_15239);
xor U16480 (N_16480,N_15207,N_15032);
xor U16481 (N_16481,N_15375,N_15471);
nand U16482 (N_16482,N_15954,N_15063);
or U16483 (N_16483,N_15817,N_15685);
nor U16484 (N_16484,N_15963,N_15362);
nand U16485 (N_16485,N_15798,N_15366);
and U16486 (N_16486,N_15181,N_15619);
xnor U16487 (N_16487,N_15939,N_15252);
nand U16488 (N_16488,N_15300,N_15779);
xnor U16489 (N_16489,N_15188,N_15279);
nor U16490 (N_16490,N_15163,N_15454);
nor U16491 (N_16491,N_15590,N_15311);
or U16492 (N_16492,N_15133,N_15830);
or U16493 (N_16493,N_15485,N_15789);
nor U16494 (N_16494,N_15651,N_15214);
nand U16495 (N_16495,N_15523,N_15350);
and U16496 (N_16496,N_15698,N_15140);
or U16497 (N_16497,N_15704,N_15409);
and U16498 (N_16498,N_15010,N_15441);
and U16499 (N_16499,N_15504,N_15046);
or U16500 (N_16500,N_15037,N_15058);
and U16501 (N_16501,N_15969,N_15487);
nor U16502 (N_16502,N_15775,N_15535);
and U16503 (N_16503,N_15199,N_15897);
nor U16504 (N_16504,N_15631,N_15755);
nor U16505 (N_16505,N_15842,N_15716);
nand U16506 (N_16506,N_15212,N_15412);
nor U16507 (N_16507,N_15819,N_15470);
nand U16508 (N_16508,N_15814,N_15996);
or U16509 (N_16509,N_15662,N_15571);
and U16510 (N_16510,N_15752,N_15466);
nor U16511 (N_16511,N_15875,N_15732);
and U16512 (N_16512,N_15164,N_15747);
nor U16513 (N_16513,N_15735,N_15415);
and U16514 (N_16514,N_15788,N_15592);
or U16515 (N_16515,N_15999,N_15013);
nor U16516 (N_16516,N_15487,N_15366);
nor U16517 (N_16517,N_15197,N_15989);
nor U16518 (N_16518,N_15185,N_15679);
nand U16519 (N_16519,N_15116,N_15722);
or U16520 (N_16520,N_15344,N_15796);
and U16521 (N_16521,N_15375,N_15873);
or U16522 (N_16522,N_15397,N_15215);
or U16523 (N_16523,N_15663,N_15145);
nor U16524 (N_16524,N_15911,N_15039);
or U16525 (N_16525,N_15423,N_15123);
xnor U16526 (N_16526,N_15778,N_15295);
nor U16527 (N_16527,N_15905,N_15434);
or U16528 (N_16528,N_15462,N_15921);
nand U16529 (N_16529,N_15202,N_15778);
xnor U16530 (N_16530,N_15202,N_15671);
nand U16531 (N_16531,N_15965,N_15472);
xnor U16532 (N_16532,N_15232,N_15958);
and U16533 (N_16533,N_15643,N_15841);
xnor U16534 (N_16534,N_15785,N_15174);
nand U16535 (N_16535,N_15529,N_15615);
xor U16536 (N_16536,N_15384,N_15660);
nand U16537 (N_16537,N_15954,N_15946);
or U16538 (N_16538,N_15432,N_15887);
nor U16539 (N_16539,N_15131,N_15323);
nor U16540 (N_16540,N_15998,N_15601);
or U16541 (N_16541,N_15591,N_15024);
nor U16542 (N_16542,N_15835,N_15736);
xnor U16543 (N_16543,N_15146,N_15813);
nand U16544 (N_16544,N_15099,N_15772);
and U16545 (N_16545,N_15372,N_15191);
or U16546 (N_16546,N_15545,N_15210);
nor U16547 (N_16547,N_15126,N_15434);
nor U16548 (N_16548,N_15131,N_15609);
nor U16549 (N_16549,N_15198,N_15373);
nand U16550 (N_16550,N_15175,N_15352);
xnor U16551 (N_16551,N_15484,N_15813);
nand U16552 (N_16552,N_15306,N_15387);
nand U16553 (N_16553,N_15019,N_15348);
xor U16554 (N_16554,N_15265,N_15267);
or U16555 (N_16555,N_15038,N_15087);
xor U16556 (N_16556,N_15792,N_15002);
nand U16557 (N_16557,N_15560,N_15753);
and U16558 (N_16558,N_15268,N_15711);
nand U16559 (N_16559,N_15879,N_15522);
nand U16560 (N_16560,N_15905,N_15372);
nand U16561 (N_16561,N_15340,N_15002);
nand U16562 (N_16562,N_15291,N_15511);
nand U16563 (N_16563,N_15772,N_15519);
and U16564 (N_16564,N_15468,N_15437);
and U16565 (N_16565,N_15351,N_15649);
nor U16566 (N_16566,N_15997,N_15447);
nor U16567 (N_16567,N_15361,N_15150);
nand U16568 (N_16568,N_15824,N_15802);
nand U16569 (N_16569,N_15048,N_15899);
and U16570 (N_16570,N_15641,N_15115);
nand U16571 (N_16571,N_15010,N_15346);
nand U16572 (N_16572,N_15741,N_15643);
nand U16573 (N_16573,N_15895,N_15126);
nand U16574 (N_16574,N_15215,N_15872);
or U16575 (N_16575,N_15594,N_15100);
nor U16576 (N_16576,N_15254,N_15265);
and U16577 (N_16577,N_15421,N_15574);
nor U16578 (N_16578,N_15173,N_15623);
or U16579 (N_16579,N_15722,N_15583);
nand U16580 (N_16580,N_15863,N_15430);
and U16581 (N_16581,N_15295,N_15109);
nor U16582 (N_16582,N_15592,N_15142);
and U16583 (N_16583,N_15360,N_15599);
or U16584 (N_16584,N_15417,N_15519);
nand U16585 (N_16585,N_15958,N_15134);
or U16586 (N_16586,N_15602,N_15570);
nor U16587 (N_16587,N_15029,N_15879);
or U16588 (N_16588,N_15711,N_15753);
nor U16589 (N_16589,N_15800,N_15005);
xnor U16590 (N_16590,N_15140,N_15977);
nor U16591 (N_16591,N_15083,N_15246);
or U16592 (N_16592,N_15346,N_15498);
xor U16593 (N_16593,N_15265,N_15752);
nand U16594 (N_16594,N_15669,N_15320);
or U16595 (N_16595,N_15349,N_15063);
xor U16596 (N_16596,N_15304,N_15462);
xnor U16597 (N_16597,N_15179,N_15761);
and U16598 (N_16598,N_15392,N_15797);
nand U16599 (N_16599,N_15702,N_15710);
nand U16600 (N_16600,N_15683,N_15920);
nand U16601 (N_16601,N_15162,N_15743);
nor U16602 (N_16602,N_15378,N_15180);
xor U16603 (N_16603,N_15122,N_15280);
and U16604 (N_16604,N_15765,N_15224);
nor U16605 (N_16605,N_15502,N_15972);
nand U16606 (N_16606,N_15015,N_15217);
nor U16607 (N_16607,N_15594,N_15589);
and U16608 (N_16608,N_15288,N_15674);
and U16609 (N_16609,N_15070,N_15578);
or U16610 (N_16610,N_15428,N_15944);
nand U16611 (N_16611,N_15698,N_15037);
nor U16612 (N_16612,N_15743,N_15352);
nand U16613 (N_16613,N_15348,N_15309);
xnor U16614 (N_16614,N_15115,N_15750);
or U16615 (N_16615,N_15884,N_15522);
or U16616 (N_16616,N_15372,N_15106);
nand U16617 (N_16617,N_15362,N_15916);
or U16618 (N_16618,N_15211,N_15801);
nor U16619 (N_16619,N_15167,N_15450);
or U16620 (N_16620,N_15215,N_15264);
xor U16621 (N_16621,N_15870,N_15654);
xor U16622 (N_16622,N_15602,N_15924);
nand U16623 (N_16623,N_15364,N_15010);
xor U16624 (N_16624,N_15087,N_15800);
xor U16625 (N_16625,N_15467,N_15087);
nand U16626 (N_16626,N_15346,N_15578);
nand U16627 (N_16627,N_15799,N_15091);
or U16628 (N_16628,N_15062,N_15823);
nand U16629 (N_16629,N_15701,N_15315);
nand U16630 (N_16630,N_15478,N_15004);
nand U16631 (N_16631,N_15477,N_15072);
or U16632 (N_16632,N_15203,N_15294);
and U16633 (N_16633,N_15006,N_15776);
or U16634 (N_16634,N_15142,N_15211);
xor U16635 (N_16635,N_15693,N_15467);
nor U16636 (N_16636,N_15162,N_15365);
xnor U16637 (N_16637,N_15876,N_15139);
xnor U16638 (N_16638,N_15008,N_15252);
or U16639 (N_16639,N_15828,N_15745);
xor U16640 (N_16640,N_15369,N_15135);
nand U16641 (N_16641,N_15339,N_15688);
and U16642 (N_16642,N_15505,N_15148);
and U16643 (N_16643,N_15247,N_15428);
or U16644 (N_16644,N_15284,N_15598);
xnor U16645 (N_16645,N_15243,N_15529);
xnor U16646 (N_16646,N_15453,N_15283);
nor U16647 (N_16647,N_15436,N_15353);
or U16648 (N_16648,N_15949,N_15416);
or U16649 (N_16649,N_15169,N_15976);
nand U16650 (N_16650,N_15572,N_15842);
nand U16651 (N_16651,N_15197,N_15963);
xnor U16652 (N_16652,N_15740,N_15558);
xnor U16653 (N_16653,N_15611,N_15964);
xor U16654 (N_16654,N_15554,N_15725);
and U16655 (N_16655,N_15812,N_15460);
and U16656 (N_16656,N_15384,N_15275);
nor U16657 (N_16657,N_15465,N_15728);
or U16658 (N_16658,N_15946,N_15696);
xor U16659 (N_16659,N_15381,N_15545);
or U16660 (N_16660,N_15689,N_15265);
nor U16661 (N_16661,N_15288,N_15298);
or U16662 (N_16662,N_15138,N_15403);
nand U16663 (N_16663,N_15996,N_15562);
and U16664 (N_16664,N_15513,N_15054);
and U16665 (N_16665,N_15981,N_15499);
nand U16666 (N_16666,N_15119,N_15788);
or U16667 (N_16667,N_15509,N_15245);
and U16668 (N_16668,N_15191,N_15352);
nand U16669 (N_16669,N_15200,N_15782);
nand U16670 (N_16670,N_15896,N_15160);
or U16671 (N_16671,N_15641,N_15973);
xnor U16672 (N_16672,N_15863,N_15804);
xnor U16673 (N_16673,N_15999,N_15220);
nand U16674 (N_16674,N_15001,N_15891);
or U16675 (N_16675,N_15294,N_15523);
xnor U16676 (N_16676,N_15465,N_15323);
nor U16677 (N_16677,N_15419,N_15389);
nand U16678 (N_16678,N_15480,N_15292);
nand U16679 (N_16679,N_15413,N_15980);
nor U16680 (N_16680,N_15727,N_15997);
or U16681 (N_16681,N_15949,N_15113);
or U16682 (N_16682,N_15145,N_15532);
or U16683 (N_16683,N_15359,N_15520);
xnor U16684 (N_16684,N_15122,N_15960);
nor U16685 (N_16685,N_15152,N_15454);
nand U16686 (N_16686,N_15890,N_15669);
or U16687 (N_16687,N_15709,N_15754);
nand U16688 (N_16688,N_15214,N_15046);
and U16689 (N_16689,N_15634,N_15012);
and U16690 (N_16690,N_15023,N_15935);
xor U16691 (N_16691,N_15222,N_15145);
or U16692 (N_16692,N_15453,N_15600);
nor U16693 (N_16693,N_15737,N_15833);
or U16694 (N_16694,N_15306,N_15529);
or U16695 (N_16695,N_15695,N_15715);
nand U16696 (N_16696,N_15609,N_15878);
and U16697 (N_16697,N_15571,N_15845);
and U16698 (N_16698,N_15166,N_15653);
nor U16699 (N_16699,N_15879,N_15191);
xor U16700 (N_16700,N_15013,N_15347);
or U16701 (N_16701,N_15674,N_15075);
xor U16702 (N_16702,N_15335,N_15641);
and U16703 (N_16703,N_15112,N_15885);
xnor U16704 (N_16704,N_15040,N_15907);
nand U16705 (N_16705,N_15016,N_15106);
nor U16706 (N_16706,N_15299,N_15026);
or U16707 (N_16707,N_15843,N_15181);
or U16708 (N_16708,N_15410,N_15152);
nand U16709 (N_16709,N_15212,N_15793);
and U16710 (N_16710,N_15908,N_15419);
nand U16711 (N_16711,N_15464,N_15052);
xnor U16712 (N_16712,N_15414,N_15092);
or U16713 (N_16713,N_15580,N_15405);
nor U16714 (N_16714,N_15932,N_15439);
nor U16715 (N_16715,N_15128,N_15028);
nor U16716 (N_16716,N_15332,N_15751);
nand U16717 (N_16717,N_15584,N_15029);
xnor U16718 (N_16718,N_15905,N_15226);
nand U16719 (N_16719,N_15017,N_15696);
xor U16720 (N_16720,N_15667,N_15324);
xor U16721 (N_16721,N_15247,N_15289);
nor U16722 (N_16722,N_15406,N_15513);
nand U16723 (N_16723,N_15977,N_15078);
xnor U16724 (N_16724,N_15453,N_15952);
and U16725 (N_16725,N_15260,N_15645);
xor U16726 (N_16726,N_15112,N_15275);
nand U16727 (N_16727,N_15140,N_15745);
and U16728 (N_16728,N_15298,N_15287);
nand U16729 (N_16729,N_15583,N_15171);
nand U16730 (N_16730,N_15747,N_15857);
or U16731 (N_16731,N_15563,N_15919);
and U16732 (N_16732,N_15082,N_15742);
nand U16733 (N_16733,N_15867,N_15190);
and U16734 (N_16734,N_15229,N_15555);
or U16735 (N_16735,N_15339,N_15485);
nor U16736 (N_16736,N_15638,N_15136);
and U16737 (N_16737,N_15456,N_15763);
or U16738 (N_16738,N_15671,N_15373);
or U16739 (N_16739,N_15705,N_15304);
and U16740 (N_16740,N_15757,N_15771);
nand U16741 (N_16741,N_15687,N_15735);
xor U16742 (N_16742,N_15138,N_15812);
nand U16743 (N_16743,N_15660,N_15623);
nand U16744 (N_16744,N_15688,N_15427);
and U16745 (N_16745,N_15603,N_15174);
nand U16746 (N_16746,N_15369,N_15696);
nor U16747 (N_16747,N_15190,N_15205);
xnor U16748 (N_16748,N_15728,N_15015);
xnor U16749 (N_16749,N_15480,N_15299);
or U16750 (N_16750,N_15875,N_15346);
and U16751 (N_16751,N_15187,N_15102);
xor U16752 (N_16752,N_15333,N_15493);
nor U16753 (N_16753,N_15232,N_15796);
nor U16754 (N_16754,N_15612,N_15385);
or U16755 (N_16755,N_15638,N_15856);
and U16756 (N_16756,N_15582,N_15682);
nor U16757 (N_16757,N_15264,N_15451);
nand U16758 (N_16758,N_15825,N_15815);
and U16759 (N_16759,N_15904,N_15550);
xnor U16760 (N_16760,N_15964,N_15615);
or U16761 (N_16761,N_15440,N_15645);
xor U16762 (N_16762,N_15442,N_15895);
and U16763 (N_16763,N_15039,N_15924);
or U16764 (N_16764,N_15587,N_15888);
xnor U16765 (N_16765,N_15611,N_15560);
xor U16766 (N_16766,N_15756,N_15206);
xnor U16767 (N_16767,N_15755,N_15779);
nor U16768 (N_16768,N_15458,N_15131);
xor U16769 (N_16769,N_15407,N_15367);
or U16770 (N_16770,N_15723,N_15452);
xnor U16771 (N_16771,N_15843,N_15322);
and U16772 (N_16772,N_15425,N_15372);
nor U16773 (N_16773,N_15603,N_15017);
or U16774 (N_16774,N_15720,N_15211);
nor U16775 (N_16775,N_15044,N_15406);
nand U16776 (N_16776,N_15321,N_15144);
nand U16777 (N_16777,N_15208,N_15860);
or U16778 (N_16778,N_15833,N_15371);
nand U16779 (N_16779,N_15510,N_15104);
and U16780 (N_16780,N_15570,N_15616);
nor U16781 (N_16781,N_15761,N_15714);
and U16782 (N_16782,N_15390,N_15001);
nand U16783 (N_16783,N_15642,N_15076);
xnor U16784 (N_16784,N_15337,N_15220);
nand U16785 (N_16785,N_15028,N_15656);
nor U16786 (N_16786,N_15040,N_15748);
and U16787 (N_16787,N_15512,N_15198);
nor U16788 (N_16788,N_15444,N_15075);
nor U16789 (N_16789,N_15600,N_15796);
nand U16790 (N_16790,N_15321,N_15761);
or U16791 (N_16791,N_15186,N_15002);
and U16792 (N_16792,N_15761,N_15433);
nand U16793 (N_16793,N_15278,N_15160);
and U16794 (N_16794,N_15217,N_15608);
or U16795 (N_16795,N_15682,N_15563);
or U16796 (N_16796,N_15307,N_15553);
nand U16797 (N_16797,N_15192,N_15087);
xor U16798 (N_16798,N_15838,N_15341);
nand U16799 (N_16799,N_15578,N_15626);
xnor U16800 (N_16800,N_15991,N_15083);
xnor U16801 (N_16801,N_15432,N_15528);
nor U16802 (N_16802,N_15535,N_15668);
and U16803 (N_16803,N_15942,N_15267);
xor U16804 (N_16804,N_15000,N_15526);
nor U16805 (N_16805,N_15352,N_15676);
nand U16806 (N_16806,N_15383,N_15371);
and U16807 (N_16807,N_15925,N_15124);
nand U16808 (N_16808,N_15144,N_15721);
or U16809 (N_16809,N_15312,N_15683);
xnor U16810 (N_16810,N_15968,N_15829);
and U16811 (N_16811,N_15747,N_15990);
nor U16812 (N_16812,N_15633,N_15983);
xor U16813 (N_16813,N_15434,N_15135);
nor U16814 (N_16814,N_15389,N_15520);
or U16815 (N_16815,N_15122,N_15320);
nor U16816 (N_16816,N_15818,N_15809);
and U16817 (N_16817,N_15912,N_15024);
and U16818 (N_16818,N_15537,N_15202);
nand U16819 (N_16819,N_15466,N_15340);
xnor U16820 (N_16820,N_15451,N_15826);
or U16821 (N_16821,N_15308,N_15809);
nand U16822 (N_16822,N_15193,N_15357);
nor U16823 (N_16823,N_15912,N_15493);
nand U16824 (N_16824,N_15175,N_15579);
or U16825 (N_16825,N_15422,N_15558);
and U16826 (N_16826,N_15987,N_15336);
or U16827 (N_16827,N_15704,N_15189);
or U16828 (N_16828,N_15200,N_15855);
or U16829 (N_16829,N_15228,N_15887);
and U16830 (N_16830,N_15255,N_15536);
and U16831 (N_16831,N_15762,N_15220);
nor U16832 (N_16832,N_15677,N_15075);
xor U16833 (N_16833,N_15591,N_15861);
nor U16834 (N_16834,N_15208,N_15342);
nand U16835 (N_16835,N_15654,N_15000);
or U16836 (N_16836,N_15385,N_15056);
nor U16837 (N_16837,N_15494,N_15081);
nand U16838 (N_16838,N_15620,N_15527);
nand U16839 (N_16839,N_15059,N_15208);
nor U16840 (N_16840,N_15548,N_15856);
or U16841 (N_16841,N_15251,N_15764);
nand U16842 (N_16842,N_15353,N_15684);
and U16843 (N_16843,N_15912,N_15223);
nor U16844 (N_16844,N_15237,N_15591);
nand U16845 (N_16845,N_15249,N_15145);
xnor U16846 (N_16846,N_15158,N_15905);
nor U16847 (N_16847,N_15970,N_15117);
and U16848 (N_16848,N_15239,N_15949);
nand U16849 (N_16849,N_15826,N_15517);
or U16850 (N_16850,N_15212,N_15245);
xor U16851 (N_16851,N_15311,N_15708);
xnor U16852 (N_16852,N_15058,N_15686);
nand U16853 (N_16853,N_15702,N_15526);
nand U16854 (N_16854,N_15731,N_15365);
and U16855 (N_16855,N_15504,N_15676);
and U16856 (N_16856,N_15628,N_15115);
nor U16857 (N_16857,N_15608,N_15400);
nand U16858 (N_16858,N_15854,N_15968);
xor U16859 (N_16859,N_15401,N_15909);
or U16860 (N_16860,N_15621,N_15302);
or U16861 (N_16861,N_15009,N_15211);
nand U16862 (N_16862,N_15039,N_15625);
or U16863 (N_16863,N_15722,N_15855);
nor U16864 (N_16864,N_15351,N_15744);
nor U16865 (N_16865,N_15501,N_15661);
or U16866 (N_16866,N_15692,N_15609);
nand U16867 (N_16867,N_15502,N_15811);
xnor U16868 (N_16868,N_15589,N_15749);
and U16869 (N_16869,N_15669,N_15683);
xor U16870 (N_16870,N_15248,N_15748);
nor U16871 (N_16871,N_15311,N_15523);
xnor U16872 (N_16872,N_15106,N_15543);
or U16873 (N_16873,N_15992,N_15868);
nor U16874 (N_16874,N_15759,N_15528);
or U16875 (N_16875,N_15947,N_15605);
nor U16876 (N_16876,N_15978,N_15531);
nand U16877 (N_16877,N_15688,N_15118);
or U16878 (N_16878,N_15201,N_15258);
nor U16879 (N_16879,N_15960,N_15057);
nor U16880 (N_16880,N_15112,N_15059);
and U16881 (N_16881,N_15457,N_15462);
xor U16882 (N_16882,N_15326,N_15661);
nand U16883 (N_16883,N_15580,N_15918);
and U16884 (N_16884,N_15785,N_15773);
nor U16885 (N_16885,N_15646,N_15821);
xor U16886 (N_16886,N_15295,N_15527);
nand U16887 (N_16887,N_15893,N_15867);
or U16888 (N_16888,N_15090,N_15425);
or U16889 (N_16889,N_15710,N_15202);
nand U16890 (N_16890,N_15030,N_15315);
nand U16891 (N_16891,N_15276,N_15263);
and U16892 (N_16892,N_15171,N_15166);
nor U16893 (N_16893,N_15290,N_15893);
and U16894 (N_16894,N_15757,N_15703);
and U16895 (N_16895,N_15121,N_15308);
or U16896 (N_16896,N_15523,N_15931);
nor U16897 (N_16897,N_15760,N_15727);
nand U16898 (N_16898,N_15945,N_15437);
and U16899 (N_16899,N_15028,N_15291);
or U16900 (N_16900,N_15329,N_15820);
xor U16901 (N_16901,N_15559,N_15188);
and U16902 (N_16902,N_15303,N_15469);
or U16903 (N_16903,N_15904,N_15299);
or U16904 (N_16904,N_15772,N_15559);
nor U16905 (N_16905,N_15093,N_15152);
xnor U16906 (N_16906,N_15156,N_15906);
nor U16907 (N_16907,N_15371,N_15765);
and U16908 (N_16908,N_15400,N_15939);
and U16909 (N_16909,N_15147,N_15400);
or U16910 (N_16910,N_15616,N_15487);
nor U16911 (N_16911,N_15011,N_15188);
or U16912 (N_16912,N_15401,N_15271);
nand U16913 (N_16913,N_15364,N_15923);
nand U16914 (N_16914,N_15258,N_15518);
and U16915 (N_16915,N_15019,N_15251);
nor U16916 (N_16916,N_15882,N_15547);
xnor U16917 (N_16917,N_15033,N_15746);
xor U16918 (N_16918,N_15566,N_15363);
and U16919 (N_16919,N_15116,N_15785);
or U16920 (N_16920,N_15111,N_15173);
and U16921 (N_16921,N_15112,N_15901);
xnor U16922 (N_16922,N_15773,N_15791);
nand U16923 (N_16923,N_15198,N_15986);
nor U16924 (N_16924,N_15915,N_15128);
and U16925 (N_16925,N_15506,N_15627);
xor U16926 (N_16926,N_15047,N_15167);
nor U16927 (N_16927,N_15857,N_15482);
and U16928 (N_16928,N_15345,N_15399);
and U16929 (N_16929,N_15576,N_15631);
or U16930 (N_16930,N_15534,N_15417);
and U16931 (N_16931,N_15940,N_15397);
nor U16932 (N_16932,N_15139,N_15540);
xnor U16933 (N_16933,N_15626,N_15740);
or U16934 (N_16934,N_15368,N_15057);
and U16935 (N_16935,N_15524,N_15836);
nor U16936 (N_16936,N_15422,N_15207);
and U16937 (N_16937,N_15678,N_15573);
nor U16938 (N_16938,N_15215,N_15726);
and U16939 (N_16939,N_15069,N_15894);
nand U16940 (N_16940,N_15607,N_15333);
nor U16941 (N_16941,N_15907,N_15788);
nand U16942 (N_16942,N_15547,N_15453);
and U16943 (N_16943,N_15778,N_15722);
nand U16944 (N_16944,N_15060,N_15845);
xor U16945 (N_16945,N_15757,N_15563);
or U16946 (N_16946,N_15057,N_15098);
nor U16947 (N_16947,N_15273,N_15147);
nand U16948 (N_16948,N_15713,N_15212);
nor U16949 (N_16949,N_15302,N_15742);
and U16950 (N_16950,N_15435,N_15726);
or U16951 (N_16951,N_15141,N_15006);
nor U16952 (N_16952,N_15159,N_15179);
nand U16953 (N_16953,N_15044,N_15489);
nor U16954 (N_16954,N_15312,N_15227);
nor U16955 (N_16955,N_15202,N_15355);
and U16956 (N_16956,N_15452,N_15823);
or U16957 (N_16957,N_15310,N_15584);
nor U16958 (N_16958,N_15241,N_15033);
nor U16959 (N_16959,N_15345,N_15220);
or U16960 (N_16960,N_15805,N_15122);
or U16961 (N_16961,N_15585,N_15069);
nand U16962 (N_16962,N_15641,N_15410);
and U16963 (N_16963,N_15953,N_15291);
nand U16964 (N_16964,N_15874,N_15997);
xor U16965 (N_16965,N_15120,N_15118);
xnor U16966 (N_16966,N_15749,N_15940);
and U16967 (N_16967,N_15157,N_15470);
or U16968 (N_16968,N_15277,N_15460);
xor U16969 (N_16969,N_15911,N_15189);
xnor U16970 (N_16970,N_15809,N_15025);
and U16971 (N_16971,N_15883,N_15259);
xor U16972 (N_16972,N_15118,N_15598);
xor U16973 (N_16973,N_15128,N_15736);
xor U16974 (N_16974,N_15286,N_15957);
xnor U16975 (N_16975,N_15976,N_15283);
xor U16976 (N_16976,N_15445,N_15130);
and U16977 (N_16977,N_15168,N_15393);
nor U16978 (N_16978,N_15511,N_15842);
nand U16979 (N_16979,N_15347,N_15402);
xnor U16980 (N_16980,N_15149,N_15729);
and U16981 (N_16981,N_15540,N_15225);
and U16982 (N_16982,N_15585,N_15682);
and U16983 (N_16983,N_15754,N_15193);
xor U16984 (N_16984,N_15491,N_15175);
and U16985 (N_16985,N_15988,N_15889);
nand U16986 (N_16986,N_15561,N_15003);
nand U16987 (N_16987,N_15855,N_15843);
nand U16988 (N_16988,N_15574,N_15569);
xnor U16989 (N_16989,N_15226,N_15197);
nand U16990 (N_16990,N_15587,N_15133);
or U16991 (N_16991,N_15734,N_15221);
nor U16992 (N_16992,N_15404,N_15712);
or U16993 (N_16993,N_15772,N_15883);
and U16994 (N_16994,N_15012,N_15882);
and U16995 (N_16995,N_15948,N_15667);
or U16996 (N_16996,N_15155,N_15943);
or U16997 (N_16997,N_15853,N_15016);
or U16998 (N_16998,N_15085,N_15042);
xor U16999 (N_16999,N_15877,N_15664);
nor U17000 (N_17000,N_16282,N_16436);
and U17001 (N_17001,N_16985,N_16298);
or U17002 (N_17002,N_16536,N_16424);
or U17003 (N_17003,N_16430,N_16165);
nor U17004 (N_17004,N_16009,N_16486);
and U17005 (N_17005,N_16245,N_16541);
and U17006 (N_17006,N_16511,N_16048);
and U17007 (N_17007,N_16172,N_16716);
nor U17008 (N_17008,N_16354,N_16023);
or U17009 (N_17009,N_16262,N_16350);
and U17010 (N_17010,N_16584,N_16862);
nand U17011 (N_17011,N_16796,N_16360);
nor U17012 (N_17012,N_16326,N_16817);
and U17013 (N_17013,N_16659,N_16612);
nor U17014 (N_17014,N_16770,N_16996);
nand U17015 (N_17015,N_16701,N_16846);
or U17016 (N_17016,N_16188,N_16873);
or U17017 (N_17017,N_16807,N_16991);
or U17018 (N_17018,N_16778,N_16575);
nor U17019 (N_17019,N_16933,N_16404);
and U17020 (N_17020,N_16487,N_16446);
xnor U17021 (N_17021,N_16342,N_16173);
xor U17022 (N_17022,N_16407,N_16561);
xor U17023 (N_17023,N_16594,N_16047);
and U17024 (N_17024,N_16473,N_16027);
xor U17025 (N_17025,N_16115,N_16621);
xor U17026 (N_17026,N_16972,N_16276);
or U17027 (N_17027,N_16368,N_16864);
nand U17028 (N_17028,N_16440,N_16085);
or U17029 (N_17029,N_16415,N_16912);
nand U17030 (N_17030,N_16179,N_16832);
nor U17031 (N_17031,N_16225,N_16026);
xnor U17032 (N_17032,N_16780,N_16878);
xnor U17033 (N_17033,N_16201,N_16177);
nand U17034 (N_17034,N_16640,N_16013);
nor U17035 (N_17035,N_16031,N_16155);
or U17036 (N_17036,N_16971,N_16274);
nor U17037 (N_17037,N_16364,N_16858);
nor U17038 (N_17038,N_16740,N_16979);
and U17039 (N_17039,N_16984,N_16443);
nand U17040 (N_17040,N_16554,N_16668);
nand U17041 (N_17041,N_16944,N_16892);
and U17042 (N_17042,N_16427,N_16284);
nand U17043 (N_17043,N_16555,N_16727);
xor U17044 (N_17044,N_16344,N_16695);
and U17045 (N_17045,N_16181,N_16736);
nor U17046 (N_17046,N_16148,N_16974);
nor U17047 (N_17047,N_16628,N_16526);
and U17048 (N_17048,N_16422,N_16635);
nand U17049 (N_17049,N_16623,N_16755);
xor U17050 (N_17050,N_16825,N_16247);
nand U17051 (N_17051,N_16560,N_16098);
or U17052 (N_17052,N_16685,N_16369);
or U17053 (N_17053,N_16549,N_16291);
xnor U17054 (N_17054,N_16738,N_16302);
or U17055 (N_17055,N_16953,N_16975);
or U17056 (N_17056,N_16752,N_16634);
nor U17057 (N_17057,N_16515,N_16688);
nor U17058 (N_17058,N_16123,N_16937);
and U17059 (N_17059,N_16679,N_16116);
nand U17060 (N_17060,N_16137,N_16058);
or U17061 (N_17061,N_16559,N_16677);
nor U17062 (N_17062,N_16769,N_16929);
nand U17063 (N_17063,N_16267,N_16530);
nor U17064 (N_17064,N_16934,N_16357);
and U17065 (N_17065,N_16647,N_16228);
nand U17066 (N_17066,N_16061,N_16012);
or U17067 (N_17067,N_16168,N_16145);
and U17068 (N_17068,N_16162,N_16080);
or U17069 (N_17069,N_16133,N_16186);
xor U17070 (N_17070,N_16469,N_16429);
xor U17071 (N_17071,N_16928,N_16684);
xor U17072 (N_17072,N_16136,N_16707);
nor U17073 (N_17073,N_16987,N_16489);
nand U17074 (N_17074,N_16994,N_16845);
xor U17075 (N_17075,N_16028,N_16384);
or U17076 (N_17076,N_16884,N_16777);
xnor U17077 (N_17077,N_16843,N_16599);
nor U17078 (N_17078,N_16563,N_16750);
xor U17079 (N_17079,N_16100,N_16015);
nor U17080 (N_17080,N_16307,N_16170);
nand U17081 (N_17081,N_16243,N_16083);
xnor U17082 (N_17082,N_16951,N_16185);
and U17083 (N_17083,N_16003,N_16576);
nand U17084 (N_17084,N_16978,N_16818);
or U17085 (N_17085,N_16318,N_16721);
xor U17086 (N_17086,N_16402,N_16257);
nand U17087 (N_17087,N_16073,N_16938);
nor U17088 (N_17088,N_16724,N_16062);
xor U17089 (N_17089,N_16689,N_16508);
nor U17090 (N_17090,N_16363,N_16040);
xnor U17091 (N_17091,N_16632,N_16230);
nand U17092 (N_17092,N_16572,N_16483);
nand U17093 (N_17093,N_16596,N_16361);
xnor U17094 (N_17094,N_16507,N_16005);
nand U17095 (N_17095,N_16460,N_16798);
xor U17096 (N_17096,N_16729,N_16731);
and U17097 (N_17097,N_16479,N_16957);
and U17098 (N_17098,N_16129,N_16333);
and U17099 (N_17099,N_16319,N_16498);
and U17100 (N_17100,N_16521,N_16334);
nor U17101 (N_17101,N_16653,N_16030);
xnor U17102 (N_17102,N_16945,N_16259);
xnor U17103 (N_17103,N_16374,N_16650);
or U17104 (N_17104,N_16683,N_16558);
nor U17105 (N_17105,N_16909,N_16279);
and U17106 (N_17106,N_16140,N_16125);
and U17107 (N_17107,N_16053,N_16159);
nand U17108 (N_17108,N_16103,N_16704);
xnor U17109 (N_17109,N_16233,N_16300);
and U17110 (N_17110,N_16019,N_16849);
nor U17111 (N_17111,N_16772,N_16900);
and U17112 (N_17112,N_16657,N_16816);
nor U17113 (N_17113,N_16639,N_16138);
nand U17114 (N_17114,N_16585,N_16389);
or U17115 (N_17115,N_16006,N_16480);
and U17116 (N_17116,N_16477,N_16393);
or U17117 (N_17117,N_16034,N_16760);
xor U17118 (N_17118,N_16820,N_16540);
nand U17119 (N_17119,N_16611,N_16157);
and U17120 (N_17120,N_16304,N_16847);
nand U17121 (N_17121,N_16497,N_16841);
nor U17122 (N_17122,N_16789,N_16306);
xor U17123 (N_17123,N_16949,N_16767);
nor U17124 (N_17124,N_16703,N_16197);
nor U17125 (N_17125,N_16008,N_16128);
or U17126 (N_17126,N_16550,N_16256);
or U17127 (N_17127,N_16359,N_16255);
nand U17128 (N_17128,N_16625,N_16021);
nor U17129 (N_17129,N_16204,N_16737);
and U17130 (N_17130,N_16775,N_16468);
and U17131 (N_17131,N_16202,N_16714);
and U17132 (N_17132,N_16792,N_16371);
nor U17133 (N_17133,N_16183,N_16207);
nand U17134 (N_17134,N_16578,N_16416);
xnor U17135 (N_17135,N_16403,N_16331);
or U17136 (N_17136,N_16887,N_16305);
nand U17137 (N_17137,N_16260,N_16311);
or U17138 (N_17138,N_16602,N_16890);
nand U17139 (N_17139,N_16806,N_16340);
and U17140 (N_17140,N_16606,N_16733);
nor U17141 (N_17141,N_16581,N_16567);
nand U17142 (N_17142,N_16896,N_16224);
nor U17143 (N_17143,N_16874,N_16124);
nand U17144 (N_17144,N_16870,N_16086);
nor U17145 (N_17145,N_16449,N_16908);
and U17146 (N_17146,N_16052,N_16889);
nor U17147 (N_17147,N_16705,N_16152);
nor U17148 (N_17148,N_16014,N_16220);
nor U17149 (N_17149,N_16232,N_16451);
nor U17150 (N_17150,N_16209,N_16398);
xnor U17151 (N_17151,N_16386,N_16999);
and U17152 (N_17152,N_16840,N_16823);
xor U17153 (N_17153,N_16670,N_16029);
nand U17154 (N_17154,N_16856,N_16831);
and U17155 (N_17155,N_16438,N_16117);
xnor U17156 (N_17156,N_16665,N_16600);
xor U17157 (N_17157,N_16886,N_16902);
and U17158 (N_17158,N_16980,N_16246);
nor U17159 (N_17159,N_16502,N_16993);
and U17160 (N_17160,N_16899,N_16089);
or U17161 (N_17161,N_16312,N_16801);
nand U17162 (N_17162,N_16335,N_16463);
nor U17163 (N_17163,N_16542,N_16154);
nand U17164 (N_17164,N_16408,N_16456);
and U17165 (N_17165,N_16283,N_16166);
xor U17166 (N_17166,N_16692,N_16854);
or U17167 (N_17167,N_16761,N_16348);
and U17168 (N_17168,N_16111,N_16482);
nand U17169 (N_17169,N_16212,N_16102);
or U17170 (N_17170,N_16397,N_16271);
and U17171 (N_17171,N_16897,N_16551);
xnor U17172 (N_17172,N_16180,N_16918);
xnor U17173 (N_17173,N_16272,N_16401);
and U17174 (N_17174,N_16470,N_16317);
nand U17175 (N_17175,N_16164,N_16566);
and U17176 (N_17176,N_16211,N_16265);
nor U17177 (N_17177,N_16144,N_16339);
or U17178 (N_17178,N_16925,N_16442);
xnor U17179 (N_17179,N_16961,N_16586);
and U17180 (N_17180,N_16147,N_16804);
or U17181 (N_17181,N_16139,N_16041);
xor U17182 (N_17182,N_16658,N_16901);
or U17183 (N_17183,N_16693,N_16523);
and U17184 (N_17184,N_16349,N_16490);
and U17185 (N_17185,N_16924,N_16732);
nor U17186 (N_17186,N_16099,N_16258);
and U17187 (N_17187,N_16966,N_16643);
nand U17188 (N_17188,N_16485,N_16464);
or U17189 (N_17189,N_16289,N_16057);
nand U17190 (N_17190,N_16454,N_16046);
nor U17191 (N_17191,N_16218,N_16253);
or U17192 (N_17192,N_16503,N_16671);
nor U17193 (N_17193,N_16184,N_16939);
nor U17194 (N_17194,N_16774,N_16134);
xnor U17195 (N_17195,N_16122,N_16370);
nand U17196 (N_17196,N_16758,N_16717);
xor U17197 (N_17197,N_16394,N_16765);
or U17198 (N_17198,N_16898,N_16084);
xnor U17199 (N_17199,N_16501,N_16904);
nand U17200 (N_17200,N_16131,N_16963);
xnor U17201 (N_17201,N_16090,N_16803);
nand U17202 (N_17202,N_16756,N_16644);
nor U17203 (N_17203,N_16678,N_16160);
or U17204 (N_17204,N_16191,N_16035);
nor U17205 (N_17205,N_16645,N_16024);
xnor U17206 (N_17206,N_16263,N_16108);
or U17207 (N_17207,N_16794,N_16534);
xor U17208 (N_17208,N_16616,N_16171);
nand U17209 (N_17209,N_16753,N_16836);
and U17210 (N_17210,N_16839,N_16141);
xnor U17211 (N_17211,N_16518,N_16075);
xnor U17212 (N_17212,N_16308,N_16377);
xnor U17213 (N_17213,N_16852,N_16982);
and U17214 (N_17214,N_16327,N_16210);
or U17215 (N_17215,N_16877,N_16802);
or U17216 (N_17216,N_16434,N_16569);
and U17217 (N_17217,N_16471,N_16719);
and U17218 (N_17218,N_16713,N_16239);
and U17219 (N_17219,N_16032,N_16888);
or U17220 (N_17220,N_16663,N_16859);
xnor U17221 (N_17221,N_16995,N_16529);
nand U17222 (N_17222,N_16496,N_16728);
and U17223 (N_17223,N_16819,N_16950);
and U17224 (N_17224,N_16715,N_16747);
xnor U17225 (N_17225,N_16835,N_16396);
xor U17226 (N_17226,N_16637,N_16885);
nand U17227 (N_17227,N_16020,N_16251);
xnor U17228 (N_17228,N_16590,N_16863);
nand U17229 (N_17229,N_16146,N_16196);
nand U17230 (N_17230,N_16343,N_16051);
xnor U17231 (N_17231,N_16895,N_16301);
or U17232 (N_17232,N_16346,N_16143);
nand U17233 (N_17233,N_16506,N_16910);
nor U17234 (N_17234,N_16287,N_16379);
nor U17235 (N_17235,N_16544,N_16475);
nand U17236 (N_17236,N_16552,N_16940);
nor U17237 (N_17237,N_16269,N_16321);
nand U17238 (N_17238,N_16524,N_16067);
nand U17239 (N_17239,N_16465,N_16288);
or U17240 (N_17240,N_16722,N_16814);
or U17241 (N_17241,N_16865,N_16484);
xor U17242 (N_17242,N_16547,N_16894);
or U17243 (N_17243,N_16474,N_16231);
and U17244 (N_17244,N_16236,N_16598);
xnor U17245 (N_17245,N_16244,N_16395);
xor U17246 (N_17246,N_16399,N_16345);
nand U17247 (N_17247,N_16783,N_16786);
nor U17248 (N_17248,N_16445,N_16193);
nand U17249 (N_17249,N_16793,N_16499);
xnor U17250 (N_17250,N_16376,N_16883);
nand U17251 (N_17251,N_16176,N_16954);
nand U17252 (N_17252,N_16278,N_16223);
nor U17253 (N_17253,N_16022,N_16879);
and U17254 (N_17254,N_16564,N_16320);
nor U17255 (N_17255,N_16292,N_16294);
nand U17256 (N_17256,N_16661,N_16367);
xor U17257 (N_17257,N_16097,N_16076);
and U17258 (N_17258,N_16927,N_16771);
or U17259 (N_17259,N_16213,N_16419);
nor U17260 (N_17260,N_16592,N_16946);
xnor U17261 (N_17261,N_16094,N_16455);
or U17262 (N_17262,N_16915,N_16007);
xor U17263 (N_17263,N_16527,N_16095);
nor U17264 (N_17264,N_16983,N_16655);
and U17265 (N_17265,N_16286,N_16106);
and U17266 (N_17266,N_16532,N_16630);
nor U17267 (N_17267,N_16044,N_16893);
nand U17268 (N_17268,N_16947,N_16597);
and U17269 (N_17269,N_16505,N_16385);
xnor U17270 (N_17270,N_16548,N_16556);
nand U17271 (N_17271,N_16811,N_16881);
nor U17272 (N_17272,N_16337,N_16459);
xor U17273 (N_17273,N_16353,N_16277);
nor U17274 (N_17274,N_16355,N_16039);
and U17275 (N_17275,N_16418,N_16314);
nor U17276 (N_17276,N_16676,N_16356);
nand U17277 (N_17277,N_16425,N_16077);
and U17278 (N_17278,N_16962,N_16038);
or U17279 (N_17279,N_16025,N_16161);
nand U17280 (N_17280,N_16341,N_16358);
or U17281 (N_17281,N_16848,N_16101);
xnor U17282 (N_17282,N_16472,N_16539);
and U17283 (N_17283,N_16064,N_16214);
nor U17284 (N_17284,N_16880,N_16720);
xor U17285 (N_17285,N_16538,N_16799);
nor U17286 (N_17286,N_16735,N_16942);
nor U17287 (N_17287,N_16215,N_16054);
and U17288 (N_17288,N_16531,N_16299);
and U17289 (N_17289,N_16219,N_16654);
or U17290 (N_17290,N_16913,N_16235);
nor U17291 (N_17291,N_16981,N_16666);
xnor U17292 (N_17292,N_16433,N_16309);
or U17293 (N_17293,N_16698,N_16092);
and U17294 (N_17294,N_16280,N_16579);
xnor U17295 (N_17295,N_16608,N_16745);
or U17296 (N_17296,N_16203,N_16866);
nor U17297 (N_17297,N_16328,N_16222);
nor U17298 (N_17298,N_16613,N_16290);
or U17299 (N_17299,N_16383,N_16553);
or U17300 (N_17300,N_16620,N_16001);
or U17301 (N_17301,N_16182,N_16624);
or U17302 (N_17302,N_16296,N_16686);
nand U17303 (N_17303,N_16956,N_16821);
xor U17304 (N_17304,N_16812,N_16651);
nor U17305 (N_17305,N_16842,N_16697);
nand U17306 (N_17306,N_16426,N_16923);
nand U17307 (N_17307,N_16411,N_16467);
xor U17308 (N_17308,N_16520,N_16838);
nor U17309 (N_17309,N_16795,N_16681);
nand U17310 (N_17310,N_16457,N_16229);
xor U17311 (N_17311,N_16788,N_16672);
and U17312 (N_17312,N_16365,N_16988);
nand U17313 (N_17313,N_16512,N_16074);
nand U17314 (N_17314,N_16113,N_16535);
or U17315 (N_17315,N_16405,N_16941);
and U17316 (N_17316,N_16329,N_16248);
nand U17317 (N_17317,N_16421,N_16293);
xor U17318 (N_17318,N_16066,N_16366);
nand U17319 (N_17319,N_16509,N_16875);
or U17320 (N_17320,N_16919,N_16577);
xnor U17321 (N_17321,N_16135,N_16297);
and U17322 (N_17322,N_16412,N_16633);
or U17323 (N_17323,N_16432,N_16593);
nand U17324 (N_17324,N_16660,N_16726);
nor U17325 (N_17325,N_16332,N_16391);
or U17326 (N_17326,N_16237,N_16943);
nor U17327 (N_17327,N_16056,N_16310);
nor U17328 (N_17328,N_16615,N_16478);
nor U17329 (N_17329,N_16510,N_16565);
nor U17330 (N_17330,N_16270,N_16711);
xnor U17331 (N_17331,N_16400,N_16087);
xor U17332 (N_17332,N_16603,N_16568);
or U17333 (N_17333,N_16986,N_16680);
nor U17334 (N_17334,N_16762,N_16249);
or U17335 (N_17335,N_16936,N_16748);
xnor U17336 (N_17336,N_16631,N_16295);
nor U17337 (N_17337,N_16158,N_16533);
xor U17338 (N_17338,N_16388,N_16238);
nor U17339 (N_17339,N_16648,N_16787);
nand U17340 (N_17340,N_16917,N_16751);
or U17341 (N_17341,N_16423,N_16322);
and U17342 (N_17342,N_16822,N_16797);
xnor U17343 (N_17343,N_16266,N_16868);
xnor U17344 (N_17344,N_16096,N_16439);
nand U17345 (N_17345,N_16800,N_16528);
nand U17346 (N_17346,N_16763,N_16649);
xnor U17347 (N_17347,N_16682,N_16206);
and U17348 (N_17348,N_16045,N_16071);
nand U17349 (N_17349,N_16313,N_16617);
nor U17350 (N_17350,N_16105,N_16065);
or U17351 (N_17351,N_16907,N_16652);
or U17352 (N_17352,N_16583,N_16330);
nand U17353 (N_17353,N_16060,N_16130);
nand U17354 (N_17354,N_16861,N_16381);
nor U17355 (N_17355,N_16221,N_16757);
nand U17356 (N_17356,N_16323,N_16759);
and U17357 (N_17357,N_16033,N_16447);
and U17358 (N_17358,N_16808,N_16725);
nand U17359 (N_17359,N_16114,N_16036);
and U17360 (N_17360,N_16187,N_16517);
nand U17361 (N_17361,N_16709,N_16261);
nand U17362 (N_17362,N_16618,N_16674);
nand U17363 (N_17363,N_16642,N_16156);
nor U17364 (N_17364,N_16132,N_16827);
or U17365 (N_17365,N_16930,N_16303);
and U17366 (N_17366,N_16543,N_16718);
nand U17367 (N_17367,N_16687,N_16574);
xor U17368 (N_17368,N_16926,N_16017);
xor U17369 (N_17369,N_16601,N_16002);
or U17370 (N_17370,N_16785,N_16607);
nor U17371 (N_17371,N_16921,N_16192);
nor U17372 (N_17372,N_16557,N_16175);
and U17373 (N_17373,N_16120,N_16694);
xor U17374 (N_17374,N_16151,N_16826);
xor U17375 (N_17375,N_16452,N_16104);
xnor U17376 (N_17376,N_16948,N_16545);
nand U17377 (N_17377,N_16285,N_16142);
or U17378 (N_17378,N_16699,N_16390);
nand U17379 (N_17379,N_16240,N_16997);
or U17380 (N_17380,N_16869,N_16829);
or U17381 (N_17381,N_16779,N_16205);
and U17382 (N_17382,N_16905,N_16088);
or U17383 (N_17383,N_16037,N_16043);
and U17384 (N_17384,N_16970,N_16629);
or U17385 (N_17385,N_16466,N_16448);
and U17386 (N_17386,N_16153,N_16782);
or U17387 (N_17387,N_16234,N_16494);
nand U17388 (N_17388,N_16911,N_16042);
and U17389 (N_17389,N_16641,N_16992);
or U17390 (N_17390,N_16435,N_16871);
nor U17391 (N_17391,N_16766,N_16739);
nor U17392 (N_17392,N_16573,N_16010);
or U17393 (N_17393,N_16857,N_16189);
nand U17394 (N_17394,N_16516,N_16562);
xnor U17395 (N_17395,N_16078,N_16275);
xnor U17396 (N_17396,N_16055,N_16018);
or U17397 (N_17397,N_16488,N_16163);
or U17398 (N_17398,N_16749,N_16790);
nor U17399 (N_17399,N_16906,N_16195);
and U17400 (N_17400,N_16476,N_16000);
xor U17401 (N_17401,N_16068,N_16112);
or U17402 (N_17402,N_16595,N_16730);
or U17403 (N_17403,N_16588,N_16109);
nand U17404 (N_17404,N_16700,N_16493);
or U17405 (N_17405,N_16273,N_16990);
xnor U17406 (N_17406,N_16741,N_16706);
nand U17407 (N_17407,N_16091,N_16968);
or U17408 (N_17408,N_16764,N_16437);
nand U17409 (N_17409,N_16315,N_16582);
and U17410 (N_17410,N_16414,N_16977);
xor U17411 (N_17411,N_16920,N_16268);
nor U17412 (N_17412,N_16387,N_16431);
nand U17413 (N_17413,N_16522,N_16610);
and U17414 (N_17414,N_16636,N_16081);
xnor U17415 (N_17415,N_16217,N_16198);
nand U17416 (N_17416,N_16169,N_16495);
or U17417 (N_17417,N_16810,N_16855);
nand U17418 (N_17418,N_16410,N_16127);
xor U17419 (N_17419,N_16050,N_16960);
xor U17420 (N_17420,N_16932,N_16491);
nand U17421 (N_17421,N_16059,N_16107);
xor U17422 (N_17422,N_16069,N_16969);
and U17423 (N_17423,N_16063,N_16675);
and U17424 (N_17424,N_16891,N_16691);
nand U17425 (N_17425,N_16093,N_16622);
and U17426 (N_17426,N_16604,N_16325);
and U17427 (N_17427,N_16872,N_16004);
nand U17428 (N_17428,N_16696,N_16955);
nand U17429 (N_17429,N_16444,N_16525);
nand U17430 (N_17430,N_16702,N_16519);
nand U17431 (N_17431,N_16500,N_16605);
xnor U17432 (N_17432,N_16481,N_16011);
and U17433 (N_17433,N_16998,N_16967);
xnor U17434 (N_17434,N_16372,N_16742);
or U17435 (N_17435,N_16614,N_16952);
or U17436 (N_17436,N_16537,N_16110);
or U17437 (N_17437,N_16815,N_16850);
nand U17438 (N_17438,N_16461,N_16504);
or U17439 (N_17439,N_16254,N_16250);
nor U17440 (N_17440,N_16914,N_16809);
or U17441 (N_17441,N_16208,N_16336);
nand U17442 (N_17442,N_16453,N_16242);
xnor U17443 (N_17443,N_16362,N_16690);
nand U17444 (N_17444,N_16199,N_16830);
and U17445 (N_17445,N_16619,N_16646);
xnor U17446 (N_17446,N_16673,N_16591);
nor U17447 (N_17447,N_16669,N_16882);
nand U17448 (N_17448,N_16965,N_16546);
nor U17449 (N_17449,N_16834,N_16813);
and U17450 (N_17450,N_16458,N_16580);
and U17451 (N_17451,N_16380,N_16420);
nand U17452 (N_17452,N_16338,N_16662);
nor U17453 (N_17453,N_16082,N_16413);
nand U17454 (N_17454,N_16450,N_16178);
xnor U17455 (N_17455,N_16072,N_16776);
and U17456 (N_17456,N_16150,N_16571);
nand U17457 (N_17457,N_16958,N_16964);
nor U17458 (N_17458,N_16226,N_16781);
and U17459 (N_17459,N_16833,N_16784);
nand U17460 (N_17460,N_16805,N_16149);
and U17461 (N_17461,N_16324,N_16626);
nand U17462 (N_17462,N_16708,N_16382);
or U17463 (N_17463,N_16828,N_16281);
and U17464 (N_17464,N_16773,N_16200);
and U17465 (N_17465,N_16916,N_16851);
xor U17466 (N_17466,N_16316,N_16079);
xnor U17467 (N_17467,N_16118,N_16216);
or U17468 (N_17468,N_16406,N_16167);
or U17469 (N_17469,N_16070,N_16375);
nor U17470 (N_17470,N_16710,N_16352);
nand U17471 (N_17471,N_16049,N_16587);
xnor U17472 (N_17472,N_16754,N_16989);
nor U17473 (N_17473,N_16174,N_16241);
and U17474 (N_17474,N_16791,N_16119);
nor U17475 (N_17475,N_16194,N_16227);
or U17476 (N_17476,N_16190,N_16723);
xnor U17477 (N_17477,N_16976,N_16378);
and U17478 (N_17478,N_16922,N_16609);
and U17479 (N_17479,N_16768,N_16126);
or U17480 (N_17480,N_16428,N_16513);
and U17481 (N_17481,N_16853,N_16392);
xor U17482 (N_17482,N_16903,N_16935);
xnor U17483 (N_17483,N_16837,N_16514);
nand U17484 (N_17484,N_16860,N_16351);
or U17485 (N_17485,N_16627,N_16743);
or U17486 (N_17486,N_16417,N_16664);
or U17487 (N_17487,N_16734,N_16264);
nor U17488 (N_17488,N_16252,N_16844);
nor U17489 (N_17489,N_16959,N_16492);
and U17490 (N_17490,N_16667,N_16121);
and U17491 (N_17491,N_16876,N_16016);
or U17492 (N_17492,N_16824,N_16973);
nor U17493 (N_17493,N_16638,N_16712);
and U17494 (N_17494,N_16462,N_16656);
nand U17495 (N_17495,N_16931,N_16744);
nor U17496 (N_17496,N_16570,N_16867);
xnor U17497 (N_17497,N_16347,N_16373);
nand U17498 (N_17498,N_16589,N_16441);
and U17499 (N_17499,N_16409,N_16746);
nand U17500 (N_17500,N_16450,N_16410);
nand U17501 (N_17501,N_16556,N_16947);
nor U17502 (N_17502,N_16860,N_16513);
and U17503 (N_17503,N_16812,N_16974);
nor U17504 (N_17504,N_16440,N_16909);
nand U17505 (N_17505,N_16768,N_16330);
and U17506 (N_17506,N_16192,N_16471);
or U17507 (N_17507,N_16172,N_16346);
xor U17508 (N_17508,N_16511,N_16948);
nand U17509 (N_17509,N_16113,N_16694);
or U17510 (N_17510,N_16403,N_16638);
xnor U17511 (N_17511,N_16710,N_16724);
xnor U17512 (N_17512,N_16299,N_16000);
and U17513 (N_17513,N_16521,N_16656);
nand U17514 (N_17514,N_16016,N_16136);
and U17515 (N_17515,N_16512,N_16957);
xor U17516 (N_17516,N_16130,N_16649);
or U17517 (N_17517,N_16997,N_16281);
or U17518 (N_17518,N_16609,N_16858);
nand U17519 (N_17519,N_16501,N_16804);
nand U17520 (N_17520,N_16208,N_16069);
nand U17521 (N_17521,N_16358,N_16058);
nand U17522 (N_17522,N_16268,N_16627);
xnor U17523 (N_17523,N_16133,N_16415);
nor U17524 (N_17524,N_16604,N_16074);
xor U17525 (N_17525,N_16511,N_16401);
nor U17526 (N_17526,N_16879,N_16438);
nor U17527 (N_17527,N_16428,N_16705);
nand U17528 (N_17528,N_16384,N_16124);
or U17529 (N_17529,N_16776,N_16107);
xnor U17530 (N_17530,N_16012,N_16314);
nand U17531 (N_17531,N_16642,N_16401);
and U17532 (N_17532,N_16166,N_16268);
xor U17533 (N_17533,N_16270,N_16960);
nand U17534 (N_17534,N_16589,N_16997);
xnor U17535 (N_17535,N_16859,N_16941);
and U17536 (N_17536,N_16774,N_16072);
xor U17537 (N_17537,N_16091,N_16503);
nor U17538 (N_17538,N_16173,N_16791);
nor U17539 (N_17539,N_16175,N_16136);
xor U17540 (N_17540,N_16937,N_16299);
and U17541 (N_17541,N_16640,N_16904);
and U17542 (N_17542,N_16536,N_16476);
and U17543 (N_17543,N_16911,N_16662);
xnor U17544 (N_17544,N_16124,N_16123);
nand U17545 (N_17545,N_16084,N_16829);
nand U17546 (N_17546,N_16007,N_16857);
nor U17547 (N_17547,N_16008,N_16308);
and U17548 (N_17548,N_16260,N_16930);
xnor U17549 (N_17549,N_16504,N_16776);
nand U17550 (N_17550,N_16223,N_16696);
xor U17551 (N_17551,N_16129,N_16247);
nand U17552 (N_17552,N_16107,N_16101);
xor U17553 (N_17553,N_16186,N_16575);
or U17554 (N_17554,N_16403,N_16427);
or U17555 (N_17555,N_16001,N_16424);
nand U17556 (N_17556,N_16381,N_16280);
and U17557 (N_17557,N_16727,N_16827);
or U17558 (N_17558,N_16013,N_16525);
nor U17559 (N_17559,N_16356,N_16745);
xnor U17560 (N_17560,N_16548,N_16282);
and U17561 (N_17561,N_16161,N_16917);
nand U17562 (N_17562,N_16291,N_16605);
and U17563 (N_17563,N_16926,N_16580);
and U17564 (N_17564,N_16834,N_16346);
nor U17565 (N_17565,N_16966,N_16220);
nand U17566 (N_17566,N_16286,N_16833);
xnor U17567 (N_17567,N_16893,N_16035);
xnor U17568 (N_17568,N_16096,N_16640);
xnor U17569 (N_17569,N_16386,N_16132);
nor U17570 (N_17570,N_16804,N_16644);
and U17571 (N_17571,N_16618,N_16798);
xor U17572 (N_17572,N_16729,N_16185);
or U17573 (N_17573,N_16547,N_16757);
and U17574 (N_17574,N_16518,N_16382);
xor U17575 (N_17575,N_16938,N_16946);
and U17576 (N_17576,N_16046,N_16016);
nand U17577 (N_17577,N_16867,N_16792);
nor U17578 (N_17578,N_16861,N_16651);
nor U17579 (N_17579,N_16263,N_16745);
or U17580 (N_17580,N_16365,N_16492);
nand U17581 (N_17581,N_16343,N_16143);
nand U17582 (N_17582,N_16727,N_16733);
nor U17583 (N_17583,N_16550,N_16095);
nand U17584 (N_17584,N_16603,N_16462);
xor U17585 (N_17585,N_16097,N_16404);
and U17586 (N_17586,N_16787,N_16044);
xor U17587 (N_17587,N_16073,N_16251);
nor U17588 (N_17588,N_16892,N_16661);
nor U17589 (N_17589,N_16242,N_16089);
or U17590 (N_17590,N_16485,N_16941);
nor U17591 (N_17591,N_16370,N_16001);
and U17592 (N_17592,N_16978,N_16571);
or U17593 (N_17593,N_16386,N_16875);
or U17594 (N_17594,N_16234,N_16695);
xnor U17595 (N_17595,N_16411,N_16661);
nor U17596 (N_17596,N_16746,N_16698);
xor U17597 (N_17597,N_16453,N_16180);
or U17598 (N_17598,N_16784,N_16259);
or U17599 (N_17599,N_16656,N_16647);
xnor U17600 (N_17600,N_16263,N_16485);
xor U17601 (N_17601,N_16347,N_16194);
and U17602 (N_17602,N_16827,N_16120);
nand U17603 (N_17603,N_16264,N_16567);
nand U17604 (N_17604,N_16350,N_16912);
and U17605 (N_17605,N_16151,N_16664);
xnor U17606 (N_17606,N_16223,N_16364);
or U17607 (N_17607,N_16870,N_16928);
or U17608 (N_17608,N_16165,N_16519);
nand U17609 (N_17609,N_16274,N_16150);
or U17610 (N_17610,N_16457,N_16930);
and U17611 (N_17611,N_16611,N_16542);
nor U17612 (N_17612,N_16969,N_16119);
and U17613 (N_17613,N_16390,N_16283);
or U17614 (N_17614,N_16769,N_16407);
xor U17615 (N_17615,N_16357,N_16642);
or U17616 (N_17616,N_16778,N_16245);
xor U17617 (N_17617,N_16008,N_16657);
xnor U17618 (N_17618,N_16847,N_16343);
or U17619 (N_17619,N_16364,N_16884);
xor U17620 (N_17620,N_16543,N_16338);
nor U17621 (N_17621,N_16451,N_16022);
nand U17622 (N_17622,N_16128,N_16245);
nor U17623 (N_17623,N_16406,N_16873);
nor U17624 (N_17624,N_16122,N_16927);
xor U17625 (N_17625,N_16193,N_16366);
nand U17626 (N_17626,N_16994,N_16106);
or U17627 (N_17627,N_16567,N_16132);
and U17628 (N_17628,N_16180,N_16825);
xnor U17629 (N_17629,N_16756,N_16810);
nor U17630 (N_17630,N_16477,N_16045);
xnor U17631 (N_17631,N_16855,N_16506);
xnor U17632 (N_17632,N_16361,N_16021);
nand U17633 (N_17633,N_16787,N_16099);
nand U17634 (N_17634,N_16974,N_16786);
and U17635 (N_17635,N_16038,N_16301);
or U17636 (N_17636,N_16494,N_16572);
nand U17637 (N_17637,N_16861,N_16641);
and U17638 (N_17638,N_16252,N_16815);
nand U17639 (N_17639,N_16447,N_16001);
nor U17640 (N_17640,N_16357,N_16293);
nor U17641 (N_17641,N_16169,N_16454);
xor U17642 (N_17642,N_16588,N_16495);
and U17643 (N_17643,N_16484,N_16498);
and U17644 (N_17644,N_16370,N_16204);
nand U17645 (N_17645,N_16729,N_16094);
nand U17646 (N_17646,N_16293,N_16414);
xnor U17647 (N_17647,N_16906,N_16460);
xor U17648 (N_17648,N_16478,N_16512);
nand U17649 (N_17649,N_16838,N_16071);
and U17650 (N_17650,N_16265,N_16551);
and U17651 (N_17651,N_16823,N_16118);
nand U17652 (N_17652,N_16295,N_16637);
nor U17653 (N_17653,N_16643,N_16134);
and U17654 (N_17654,N_16250,N_16618);
xor U17655 (N_17655,N_16401,N_16076);
or U17656 (N_17656,N_16116,N_16552);
or U17657 (N_17657,N_16057,N_16034);
xor U17658 (N_17658,N_16876,N_16851);
nand U17659 (N_17659,N_16092,N_16694);
nand U17660 (N_17660,N_16856,N_16696);
nor U17661 (N_17661,N_16769,N_16884);
nor U17662 (N_17662,N_16365,N_16374);
or U17663 (N_17663,N_16203,N_16686);
and U17664 (N_17664,N_16366,N_16352);
nand U17665 (N_17665,N_16664,N_16629);
xnor U17666 (N_17666,N_16760,N_16114);
or U17667 (N_17667,N_16448,N_16417);
nor U17668 (N_17668,N_16212,N_16196);
or U17669 (N_17669,N_16201,N_16116);
and U17670 (N_17670,N_16510,N_16663);
nor U17671 (N_17671,N_16637,N_16584);
nor U17672 (N_17672,N_16771,N_16999);
xor U17673 (N_17673,N_16732,N_16157);
and U17674 (N_17674,N_16973,N_16552);
nor U17675 (N_17675,N_16064,N_16978);
nand U17676 (N_17676,N_16472,N_16133);
or U17677 (N_17677,N_16828,N_16871);
and U17678 (N_17678,N_16926,N_16055);
and U17679 (N_17679,N_16472,N_16496);
xor U17680 (N_17680,N_16952,N_16575);
and U17681 (N_17681,N_16774,N_16062);
nor U17682 (N_17682,N_16380,N_16967);
nand U17683 (N_17683,N_16555,N_16776);
or U17684 (N_17684,N_16701,N_16178);
and U17685 (N_17685,N_16360,N_16856);
nand U17686 (N_17686,N_16679,N_16294);
nand U17687 (N_17687,N_16519,N_16970);
xnor U17688 (N_17688,N_16596,N_16485);
nand U17689 (N_17689,N_16563,N_16467);
nor U17690 (N_17690,N_16423,N_16904);
nand U17691 (N_17691,N_16249,N_16472);
xor U17692 (N_17692,N_16340,N_16289);
or U17693 (N_17693,N_16761,N_16305);
or U17694 (N_17694,N_16842,N_16088);
and U17695 (N_17695,N_16219,N_16090);
nor U17696 (N_17696,N_16560,N_16891);
and U17697 (N_17697,N_16248,N_16114);
or U17698 (N_17698,N_16315,N_16433);
and U17699 (N_17699,N_16294,N_16009);
xor U17700 (N_17700,N_16569,N_16094);
xor U17701 (N_17701,N_16195,N_16863);
nor U17702 (N_17702,N_16022,N_16951);
and U17703 (N_17703,N_16883,N_16517);
nand U17704 (N_17704,N_16222,N_16708);
xnor U17705 (N_17705,N_16612,N_16831);
nor U17706 (N_17706,N_16055,N_16905);
or U17707 (N_17707,N_16772,N_16891);
or U17708 (N_17708,N_16199,N_16026);
nand U17709 (N_17709,N_16613,N_16638);
nor U17710 (N_17710,N_16130,N_16910);
or U17711 (N_17711,N_16456,N_16190);
nand U17712 (N_17712,N_16093,N_16482);
xor U17713 (N_17713,N_16049,N_16621);
and U17714 (N_17714,N_16978,N_16185);
or U17715 (N_17715,N_16215,N_16227);
nand U17716 (N_17716,N_16458,N_16819);
xnor U17717 (N_17717,N_16591,N_16517);
or U17718 (N_17718,N_16458,N_16582);
or U17719 (N_17719,N_16942,N_16407);
and U17720 (N_17720,N_16766,N_16816);
xnor U17721 (N_17721,N_16845,N_16151);
and U17722 (N_17722,N_16584,N_16062);
nand U17723 (N_17723,N_16591,N_16400);
nand U17724 (N_17724,N_16022,N_16591);
xnor U17725 (N_17725,N_16807,N_16561);
nand U17726 (N_17726,N_16676,N_16110);
xnor U17727 (N_17727,N_16876,N_16741);
and U17728 (N_17728,N_16229,N_16757);
and U17729 (N_17729,N_16546,N_16555);
nor U17730 (N_17730,N_16811,N_16769);
nor U17731 (N_17731,N_16612,N_16959);
or U17732 (N_17732,N_16295,N_16968);
xor U17733 (N_17733,N_16580,N_16917);
and U17734 (N_17734,N_16179,N_16938);
and U17735 (N_17735,N_16327,N_16083);
nor U17736 (N_17736,N_16764,N_16353);
or U17737 (N_17737,N_16045,N_16024);
nor U17738 (N_17738,N_16717,N_16837);
xnor U17739 (N_17739,N_16577,N_16023);
xor U17740 (N_17740,N_16503,N_16333);
xor U17741 (N_17741,N_16491,N_16784);
nand U17742 (N_17742,N_16597,N_16749);
and U17743 (N_17743,N_16641,N_16075);
nand U17744 (N_17744,N_16377,N_16533);
and U17745 (N_17745,N_16096,N_16291);
and U17746 (N_17746,N_16564,N_16740);
nor U17747 (N_17747,N_16000,N_16044);
and U17748 (N_17748,N_16901,N_16821);
and U17749 (N_17749,N_16564,N_16822);
nor U17750 (N_17750,N_16183,N_16720);
nor U17751 (N_17751,N_16803,N_16424);
or U17752 (N_17752,N_16062,N_16470);
nor U17753 (N_17753,N_16874,N_16899);
or U17754 (N_17754,N_16049,N_16329);
or U17755 (N_17755,N_16322,N_16665);
nor U17756 (N_17756,N_16420,N_16101);
nor U17757 (N_17757,N_16126,N_16627);
xnor U17758 (N_17758,N_16702,N_16518);
and U17759 (N_17759,N_16038,N_16081);
nand U17760 (N_17760,N_16049,N_16420);
or U17761 (N_17761,N_16298,N_16152);
xor U17762 (N_17762,N_16764,N_16438);
nand U17763 (N_17763,N_16427,N_16729);
and U17764 (N_17764,N_16689,N_16285);
nor U17765 (N_17765,N_16287,N_16520);
and U17766 (N_17766,N_16078,N_16508);
and U17767 (N_17767,N_16430,N_16934);
nand U17768 (N_17768,N_16192,N_16449);
nand U17769 (N_17769,N_16965,N_16137);
and U17770 (N_17770,N_16076,N_16881);
nand U17771 (N_17771,N_16604,N_16492);
and U17772 (N_17772,N_16106,N_16741);
nor U17773 (N_17773,N_16312,N_16291);
xor U17774 (N_17774,N_16423,N_16871);
nor U17775 (N_17775,N_16336,N_16753);
or U17776 (N_17776,N_16361,N_16585);
and U17777 (N_17777,N_16272,N_16420);
or U17778 (N_17778,N_16657,N_16271);
or U17779 (N_17779,N_16623,N_16933);
xnor U17780 (N_17780,N_16190,N_16178);
or U17781 (N_17781,N_16683,N_16908);
nand U17782 (N_17782,N_16423,N_16163);
xnor U17783 (N_17783,N_16307,N_16046);
or U17784 (N_17784,N_16062,N_16227);
or U17785 (N_17785,N_16093,N_16263);
or U17786 (N_17786,N_16585,N_16905);
nor U17787 (N_17787,N_16803,N_16981);
nor U17788 (N_17788,N_16538,N_16049);
xnor U17789 (N_17789,N_16252,N_16014);
xnor U17790 (N_17790,N_16864,N_16183);
nand U17791 (N_17791,N_16895,N_16185);
and U17792 (N_17792,N_16671,N_16234);
nand U17793 (N_17793,N_16204,N_16812);
nand U17794 (N_17794,N_16338,N_16519);
nand U17795 (N_17795,N_16577,N_16913);
nand U17796 (N_17796,N_16494,N_16142);
and U17797 (N_17797,N_16807,N_16611);
nor U17798 (N_17798,N_16356,N_16518);
xnor U17799 (N_17799,N_16933,N_16408);
and U17800 (N_17800,N_16297,N_16833);
and U17801 (N_17801,N_16932,N_16906);
and U17802 (N_17802,N_16983,N_16788);
or U17803 (N_17803,N_16158,N_16026);
or U17804 (N_17804,N_16035,N_16941);
or U17805 (N_17805,N_16879,N_16915);
or U17806 (N_17806,N_16936,N_16162);
nand U17807 (N_17807,N_16410,N_16836);
xor U17808 (N_17808,N_16873,N_16443);
and U17809 (N_17809,N_16385,N_16217);
and U17810 (N_17810,N_16825,N_16403);
nand U17811 (N_17811,N_16271,N_16019);
and U17812 (N_17812,N_16942,N_16489);
nor U17813 (N_17813,N_16082,N_16282);
xor U17814 (N_17814,N_16352,N_16208);
xor U17815 (N_17815,N_16089,N_16383);
nand U17816 (N_17816,N_16960,N_16767);
nor U17817 (N_17817,N_16222,N_16275);
nand U17818 (N_17818,N_16386,N_16834);
or U17819 (N_17819,N_16352,N_16238);
nor U17820 (N_17820,N_16292,N_16960);
and U17821 (N_17821,N_16975,N_16490);
nor U17822 (N_17822,N_16640,N_16435);
nand U17823 (N_17823,N_16094,N_16442);
and U17824 (N_17824,N_16695,N_16959);
xnor U17825 (N_17825,N_16654,N_16075);
and U17826 (N_17826,N_16526,N_16408);
nand U17827 (N_17827,N_16942,N_16741);
nor U17828 (N_17828,N_16099,N_16936);
nand U17829 (N_17829,N_16077,N_16737);
xor U17830 (N_17830,N_16239,N_16514);
xor U17831 (N_17831,N_16704,N_16129);
nor U17832 (N_17832,N_16397,N_16931);
nor U17833 (N_17833,N_16763,N_16723);
nor U17834 (N_17834,N_16594,N_16382);
nand U17835 (N_17835,N_16114,N_16887);
nand U17836 (N_17836,N_16780,N_16065);
or U17837 (N_17837,N_16406,N_16137);
or U17838 (N_17838,N_16770,N_16969);
xnor U17839 (N_17839,N_16192,N_16006);
and U17840 (N_17840,N_16117,N_16175);
nand U17841 (N_17841,N_16664,N_16558);
nor U17842 (N_17842,N_16921,N_16628);
and U17843 (N_17843,N_16658,N_16279);
nor U17844 (N_17844,N_16105,N_16716);
or U17845 (N_17845,N_16765,N_16810);
or U17846 (N_17846,N_16662,N_16125);
or U17847 (N_17847,N_16351,N_16838);
nand U17848 (N_17848,N_16533,N_16479);
or U17849 (N_17849,N_16661,N_16127);
and U17850 (N_17850,N_16556,N_16036);
or U17851 (N_17851,N_16775,N_16729);
and U17852 (N_17852,N_16017,N_16988);
or U17853 (N_17853,N_16174,N_16671);
xnor U17854 (N_17854,N_16634,N_16581);
and U17855 (N_17855,N_16499,N_16465);
nor U17856 (N_17856,N_16954,N_16715);
or U17857 (N_17857,N_16934,N_16331);
nand U17858 (N_17858,N_16902,N_16532);
nor U17859 (N_17859,N_16283,N_16831);
nor U17860 (N_17860,N_16207,N_16007);
xor U17861 (N_17861,N_16965,N_16043);
nor U17862 (N_17862,N_16690,N_16471);
nand U17863 (N_17863,N_16937,N_16507);
nor U17864 (N_17864,N_16688,N_16584);
or U17865 (N_17865,N_16012,N_16827);
or U17866 (N_17866,N_16758,N_16352);
xnor U17867 (N_17867,N_16682,N_16346);
nand U17868 (N_17868,N_16417,N_16694);
xor U17869 (N_17869,N_16100,N_16110);
xnor U17870 (N_17870,N_16809,N_16155);
xnor U17871 (N_17871,N_16834,N_16905);
xor U17872 (N_17872,N_16180,N_16173);
xnor U17873 (N_17873,N_16732,N_16672);
or U17874 (N_17874,N_16980,N_16071);
nand U17875 (N_17875,N_16358,N_16870);
xnor U17876 (N_17876,N_16722,N_16726);
nor U17877 (N_17877,N_16465,N_16266);
or U17878 (N_17878,N_16839,N_16677);
nor U17879 (N_17879,N_16685,N_16543);
xnor U17880 (N_17880,N_16387,N_16654);
nor U17881 (N_17881,N_16979,N_16015);
nand U17882 (N_17882,N_16804,N_16858);
xor U17883 (N_17883,N_16552,N_16701);
xnor U17884 (N_17884,N_16430,N_16131);
and U17885 (N_17885,N_16944,N_16641);
and U17886 (N_17886,N_16048,N_16829);
and U17887 (N_17887,N_16625,N_16404);
xor U17888 (N_17888,N_16700,N_16964);
nand U17889 (N_17889,N_16732,N_16872);
or U17890 (N_17890,N_16701,N_16460);
and U17891 (N_17891,N_16658,N_16125);
and U17892 (N_17892,N_16849,N_16671);
xor U17893 (N_17893,N_16339,N_16640);
or U17894 (N_17894,N_16615,N_16955);
or U17895 (N_17895,N_16588,N_16998);
nand U17896 (N_17896,N_16130,N_16098);
or U17897 (N_17897,N_16050,N_16410);
nor U17898 (N_17898,N_16258,N_16133);
nor U17899 (N_17899,N_16378,N_16384);
xnor U17900 (N_17900,N_16671,N_16827);
and U17901 (N_17901,N_16069,N_16086);
nand U17902 (N_17902,N_16766,N_16897);
nand U17903 (N_17903,N_16586,N_16508);
xnor U17904 (N_17904,N_16460,N_16490);
nand U17905 (N_17905,N_16597,N_16336);
nor U17906 (N_17906,N_16078,N_16519);
nor U17907 (N_17907,N_16078,N_16956);
or U17908 (N_17908,N_16139,N_16264);
and U17909 (N_17909,N_16675,N_16411);
xnor U17910 (N_17910,N_16747,N_16285);
and U17911 (N_17911,N_16688,N_16250);
xnor U17912 (N_17912,N_16680,N_16643);
or U17913 (N_17913,N_16010,N_16277);
nand U17914 (N_17914,N_16758,N_16076);
nor U17915 (N_17915,N_16443,N_16783);
xor U17916 (N_17916,N_16836,N_16725);
xnor U17917 (N_17917,N_16445,N_16761);
xnor U17918 (N_17918,N_16305,N_16347);
and U17919 (N_17919,N_16849,N_16378);
xor U17920 (N_17920,N_16267,N_16598);
nor U17921 (N_17921,N_16415,N_16094);
nand U17922 (N_17922,N_16125,N_16454);
or U17923 (N_17923,N_16290,N_16324);
or U17924 (N_17924,N_16155,N_16924);
nor U17925 (N_17925,N_16931,N_16790);
xnor U17926 (N_17926,N_16644,N_16102);
nand U17927 (N_17927,N_16554,N_16614);
xor U17928 (N_17928,N_16842,N_16730);
xor U17929 (N_17929,N_16295,N_16685);
and U17930 (N_17930,N_16497,N_16025);
nand U17931 (N_17931,N_16969,N_16435);
nor U17932 (N_17932,N_16043,N_16640);
nand U17933 (N_17933,N_16370,N_16921);
xor U17934 (N_17934,N_16997,N_16101);
nor U17935 (N_17935,N_16707,N_16462);
xnor U17936 (N_17936,N_16294,N_16317);
and U17937 (N_17937,N_16706,N_16814);
nand U17938 (N_17938,N_16887,N_16237);
nand U17939 (N_17939,N_16070,N_16970);
nand U17940 (N_17940,N_16108,N_16375);
and U17941 (N_17941,N_16944,N_16942);
nor U17942 (N_17942,N_16510,N_16970);
and U17943 (N_17943,N_16179,N_16114);
nand U17944 (N_17944,N_16983,N_16706);
xnor U17945 (N_17945,N_16587,N_16372);
or U17946 (N_17946,N_16258,N_16375);
and U17947 (N_17947,N_16265,N_16003);
nand U17948 (N_17948,N_16917,N_16450);
nand U17949 (N_17949,N_16713,N_16549);
xnor U17950 (N_17950,N_16783,N_16441);
or U17951 (N_17951,N_16178,N_16940);
xnor U17952 (N_17952,N_16458,N_16208);
xor U17953 (N_17953,N_16865,N_16978);
nor U17954 (N_17954,N_16224,N_16118);
and U17955 (N_17955,N_16076,N_16941);
nand U17956 (N_17956,N_16670,N_16413);
or U17957 (N_17957,N_16026,N_16382);
nor U17958 (N_17958,N_16185,N_16265);
xnor U17959 (N_17959,N_16546,N_16910);
and U17960 (N_17960,N_16195,N_16239);
or U17961 (N_17961,N_16737,N_16620);
xor U17962 (N_17962,N_16667,N_16291);
or U17963 (N_17963,N_16302,N_16196);
and U17964 (N_17964,N_16525,N_16745);
nand U17965 (N_17965,N_16456,N_16450);
and U17966 (N_17966,N_16219,N_16685);
nor U17967 (N_17967,N_16005,N_16455);
or U17968 (N_17968,N_16863,N_16327);
and U17969 (N_17969,N_16227,N_16979);
and U17970 (N_17970,N_16784,N_16462);
nor U17971 (N_17971,N_16686,N_16193);
and U17972 (N_17972,N_16699,N_16190);
xnor U17973 (N_17973,N_16568,N_16494);
or U17974 (N_17974,N_16273,N_16428);
nand U17975 (N_17975,N_16489,N_16705);
nand U17976 (N_17976,N_16115,N_16176);
and U17977 (N_17977,N_16379,N_16481);
xnor U17978 (N_17978,N_16386,N_16064);
xnor U17979 (N_17979,N_16462,N_16376);
and U17980 (N_17980,N_16185,N_16525);
xnor U17981 (N_17981,N_16830,N_16639);
and U17982 (N_17982,N_16160,N_16142);
nor U17983 (N_17983,N_16248,N_16738);
nor U17984 (N_17984,N_16712,N_16288);
xor U17985 (N_17985,N_16967,N_16599);
xor U17986 (N_17986,N_16209,N_16932);
nor U17987 (N_17987,N_16249,N_16367);
or U17988 (N_17988,N_16061,N_16656);
or U17989 (N_17989,N_16887,N_16661);
or U17990 (N_17990,N_16257,N_16325);
or U17991 (N_17991,N_16617,N_16998);
and U17992 (N_17992,N_16065,N_16977);
or U17993 (N_17993,N_16802,N_16194);
and U17994 (N_17994,N_16666,N_16808);
and U17995 (N_17995,N_16759,N_16862);
nor U17996 (N_17996,N_16906,N_16371);
nor U17997 (N_17997,N_16657,N_16195);
or U17998 (N_17998,N_16606,N_16061);
xor U17999 (N_17999,N_16751,N_16098);
xor U18000 (N_18000,N_17699,N_17782);
or U18001 (N_18001,N_17648,N_17797);
and U18002 (N_18002,N_17879,N_17767);
nor U18003 (N_18003,N_17590,N_17530);
nand U18004 (N_18004,N_17096,N_17633);
nor U18005 (N_18005,N_17892,N_17703);
nand U18006 (N_18006,N_17411,N_17283);
or U18007 (N_18007,N_17870,N_17627);
or U18008 (N_18008,N_17134,N_17151);
xor U18009 (N_18009,N_17152,N_17754);
nand U18010 (N_18010,N_17400,N_17551);
and U18011 (N_18011,N_17208,N_17364);
and U18012 (N_18012,N_17292,N_17576);
or U18013 (N_18013,N_17557,N_17068);
xor U18014 (N_18014,N_17030,N_17313);
xnor U18015 (N_18015,N_17671,N_17841);
and U18016 (N_18016,N_17000,N_17696);
and U18017 (N_18017,N_17658,N_17942);
nand U18018 (N_18018,N_17641,N_17715);
nor U18019 (N_18019,N_17444,N_17562);
nand U18020 (N_18020,N_17114,N_17407);
and U18021 (N_18021,N_17278,N_17631);
or U18022 (N_18022,N_17970,N_17501);
or U18023 (N_18023,N_17736,N_17693);
nand U18024 (N_18024,N_17384,N_17286);
or U18025 (N_18025,N_17630,N_17546);
or U18026 (N_18026,N_17183,N_17388);
or U18027 (N_18027,N_17695,N_17868);
xnor U18028 (N_18028,N_17135,N_17506);
nand U18029 (N_18029,N_17265,N_17498);
nand U18030 (N_18030,N_17539,N_17988);
and U18031 (N_18031,N_17670,N_17303);
and U18032 (N_18032,N_17236,N_17533);
nor U18033 (N_18033,N_17386,N_17418);
and U18034 (N_18034,N_17740,N_17429);
xnor U18035 (N_18035,N_17010,N_17651);
or U18036 (N_18036,N_17331,N_17689);
xnor U18037 (N_18037,N_17452,N_17103);
nor U18038 (N_18038,N_17713,N_17772);
nor U18039 (N_18039,N_17999,N_17849);
or U18040 (N_18040,N_17345,N_17910);
nor U18041 (N_18041,N_17322,N_17613);
xnor U18042 (N_18042,N_17416,N_17143);
xnor U18043 (N_18043,N_17535,N_17990);
nand U18044 (N_18044,N_17329,N_17674);
nand U18045 (N_18045,N_17099,N_17047);
nand U18046 (N_18046,N_17110,N_17298);
nor U18047 (N_18047,N_17887,N_17543);
and U18048 (N_18048,N_17355,N_17904);
and U18049 (N_18049,N_17802,N_17690);
nand U18050 (N_18050,N_17512,N_17734);
or U18051 (N_18051,N_17757,N_17838);
and U18052 (N_18052,N_17818,N_17202);
or U18053 (N_18053,N_17247,N_17796);
and U18054 (N_18054,N_17607,N_17759);
and U18055 (N_18055,N_17371,N_17375);
nor U18056 (N_18056,N_17780,N_17795);
or U18057 (N_18057,N_17005,N_17973);
and U18058 (N_18058,N_17336,N_17253);
and U18059 (N_18059,N_17321,N_17585);
nand U18060 (N_18060,N_17333,N_17248);
nand U18061 (N_18061,N_17428,N_17747);
and U18062 (N_18062,N_17786,N_17544);
xnor U18063 (N_18063,N_17197,N_17308);
nor U18064 (N_18064,N_17495,N_17620);
or U18065 (N_18065,N_17687,N_17864);
and U18066 (N_18066,N_17464,N_17145);
nand U18067 (N_18067,N_17271,N_17707);
nand U18068 (N_18068,N_17396,N_17514);
nor U18069 (N_18069,N_17729,N_17285);
or U18070 (N_18070,N_17097,N_17349);
and U18071 (N_18071,N_17427,N_17575);
and U18072 (N_18072,N_17160,N_17784);
or U18073 (N_18073,N_17593,N_17179);
xnor U18074 (N_18074,N_17888,N_17794);
or U18075 (N_18075,N_17803,N_17347);
nor U18076 (N_18076,N_17320,N_17601);
or U18077 (N_18077,N_17680,N_17969);
nor U18078 (N_18078,N_17367,N_17884);
and U18079 (N_18079,N_17527,N_17978);
nand U18080 (N_18080,N_17591,N_17455);
nor U18081 (N_18081,N_17812,N_17291);
or U18082 (N_18082,N_17040,N_17629);
or U18083 (N_18083,N_17877,N_17675);
nor U18084 (N_18084,N_17956,N_17581);
and U18085 (N_18085,N_17775,N_17223);
and U18086 (N_18086,N_17664,N_17288);
or U18087 (N_18087,N_17279,N_17979);
and U18088 (N_18088,N_17485,N_17661);
or U18089 (N_18089,N_17063,N_17017);
nand U18090 (N_18090,N_17635,N_17166);
xnor U18091 (N_18091,N_17305,N_17440);
or U18092 (N_18092,N_17564,N_17245);
and U18093 (N_18093,N_17339,N_17568);
and U18094 (N_18094,N_17710,N_17106);
or U18095 (N_18095,N_17259,N_17799);
nor U18096 (N_18096,N_17697,N_17177);
nand U18097 (N_18097,N_17161,N_17924);
and U18098 (N_18098,N_17597,N_17625);
nand U18099 (N_18099,N_17348,N_17943);
nand U18100 (N_18100,N_17511,N_17310);
nand U18101 (N_18101,N_17328,N_17843);
xor U18102 (N_18102,N_17857,N_17982);
nand U18103 (N_18103,N_17266,N_17914);
nand U18104 (N_18104,N_17122,N_17038);
xor U18105 (N_18105,N_17457,N_17281);
and U18106 (N_18106,N_17340,N_17876);
xor U18107 (N_18107,N_17437,N_17002);
or U18108 (N_18108,N_17256,N_17178);
and U18109 (N_18109,N_17337,N_17617);
nor U18110 (N_18110,N_17822,N_17257);
nor U18111 (N_18111,N_17450,N_17953);
xor U18112 (N_18112,N_17380,N_17078);
nand U18113 (N_18113,N_17883,N_17120);
or U18114 (N_18114,N_17940,N_17523);
xnor U18115 (N_18115,N_17750,N_17714);
and U18116 (N_18116,N_17189,N_17109);
xnor U18117 (N_18117,N_17112,N_17372);
nand U18118 (N_18118,N_17473,N_17731);
xor U18119 (N_18119,N_17569,N_17733);
or U18120 (N_18120,N_17324,N_17505);
or U18121 (N_18121,N_17126,N_17346);
nor U18122 (N_18122,N_17272,N_17301);
nor U18123 (N_18123,N_17659,N_17541);
xor U18124 (N_18124,N_17808,N_17685);
nand U18125 (N_18125,N_17837,N_17438);
or U18126 (N_18126,N_17701,N_17762);
nand U18127 (N_18127,N_17850,N_17957);
nor U18128 (N_18128,N_17077,N_17792);
and U18129 (N_18129,N_17974,N_17362);
nand U18130 (N_18130,N_17267,N_17730);
xor U18131 (N_18131,N_17052,N_17559);
nand U18132 (N_18132,N_17422,N_17600);
nand U18133 (N_18133,N_17127,N_17167);
or U18134 (N_18134,N_17069,N_17011);
nor U18135 (N_18135,N_17132,N_17018);
nand U18136 (N_18136,N_17677,N_17354);
nand U18137 (N_18137,N_17072,N_17662);
and U18138 (N_18138,N_17834,N_17828);
and U18139 (N_18139,N_17216,N_17359);
or U18140 (N_18140,N_17251,N_17948);
and U18141 (N_18141,N_17980,N_17420);
and U18142 (N_18142,N_17382,N_17073);
nor U18143 (N_18143,N_17711,N_17560);
and U18144 (N_18144,N_17954,N_17376);
and U18145 (N_18145,N_17025,N_17358);
and U18146 (N_18146,N_17261,N_17201);
nand U18147 (N_18147,N_17255,N_17862);
nor U18148 (N_18148,N_17379,N_17436);
nand U18149 (N_18149,N_17451,N_17181);
or U18150 (N_18150,N_17706,N_17724);
xnor U18151 (N_18151,N_17262,N_17162);
nand U18152 (N_18152,N_17971,N_17556);
xor U18153 (N_18153,N_17726,N_17075);
nor U18154 (N_18154,N_17447,N_17920);
nand U18155 (N_18155,N_17667,N_17091);
or U18156 (N_18156,N_17960,N_17975);
or U18157 (N_18157,N_17609,N_17213);
nor U18158 (N_18158,N_17654,N_17489);
xor U18159 (N_18159,N_17705,N_17153);
nor U18160 (N_18160,N_17592,N_17951);
nand U18161 (N_18161,N_17493,N_17555);
or U18162 (N_18162,N_17009,N_17764);
and U18163 (N_18163,N_17287,N_17570);
and U18164 (N_18164,N_17070,N_17210);
nand U18165 (N_18165,N_17242,N_17778);
and U18166 (N_18166,N_17188,N_17603);
and U18167 (N_18167,N_17963,N_17840);
nand U18168 (N_18168,N_17579,N_17475);
and U18169 (N_18169,N_17553,N_17660);
nand U18170 (N_18170,N_17871,N_17545);
and U18171 (N_18171,N_17854,N_17390);
or U18172 (N_18172,N_17300,N_17832);
nor U18173 (N_18173,N_17566,N_17826);
xnor U18174 (N_18174,N_17398,N_17098);
nor U18175 (N_18175,N_17147,N_17766);
nor U18176 (N_18176,N_17144,N_17691);
or U18177 (N_18177,N_17062,N_17855);
nor U18178 (N_18178,N_17908,N_17031);
nand U18179 (N_18179,N_17430,N_17923);
and U18180 (N_18180,N_17909,N_17852);
nor U18181 (N_18181,N_17700,N_17540);
nor U18182 (N_18182,N_17875,N_17433);
xnor U18183 (N_18183,N_17024,N_17623);
nor U18184 (N_18184,N_17995,N_17064);
nand U18185 (N_18185,N_17142,N_17155);
nor U18186 (N_18186,N_17751,N_17692);
nand U18187 (N_18187,N_17820,N_17851);
xnor U18188 (N_18188,N_17381,N_17366);
nand U18189 (N_18189,N_17182,N_17237);
nand U18190 (N_18190,N_17041,N_17967);
or U18191 (N_18191,N_17749,N_17365);
xnor U18192 (N_18192,N_17769,N_17048);
nor U18193 (N_18193,N_17829,N_17330);
and U18194 (N_18194,N_17897,N_17785);
or U18195 (N_18195,N_17352,N_17952);
nand U18196 (N_18196,N_17742,N_17946);
xnor U18197 (N_18197,N_17273,N_17720);
and U18198 (N_18198,N_17499,N_17089);
or U18199 (N_18199,N_17905,N_17642);
and U18200 (N_18200,N_17636,N_17171);
nor U18201 (N_18201,N_17094,N_17916);
and U18202 (N_18202,N_17317,N_17626);
xnor U18203 (N_18203,N_17363,N_17481);
and U18204 (N_18204,N_17141,N_17319);
or U18205 (N_18205,N_17497,N_17193);
and U18206 (N_18206,N_17831,N_17175);
nor U18207 (N_18207,N_17516,N_17578);
nand U18208 (N_18208,N_17338,N_17529);
or U18209 (N_18209,N_17415,N_17694);
nand U18210 (N_18210,N_17611,N_17244);
or U18211 (N_18211,N_17474,N_17921);
xnor U18212 (N_18212,N_17302,N_17067);
xor U18213 (N_18213,N_17977,N_17056);
xor U18214 (N_18214,N_17239,N_17774);
or U18215 (N_18215,N_17325,N_17823);
nand U18216 (N_18216,N_17001,N_17088);
and U18217 (N_18217,N_17361,N_17463);
or U18218 (N_18218,N_17824,N_17483);
xnor U18219 (N_18219,N_17140,N_17789);
or U18220 (N_18220,N_17113,N_17399);
nor U18221 (N_18221,N_17394,N_17676);
and U18222 (N_18222,N_17554,N_17655);
nand U18223 (N_18223,N_17966,N_17370);
or U18224 (N_18224,N_17218,N_17698);
nor U18225 (N_18225,N_17709,N_17863);
nand U18226 (N_18226,N_17180,N_17735);
and U18227 (N_18227,N_17421,N_17748);
and U18228 (N_18228,N_17552,N_17472);
and U18229 (N_18229,N_17962,N_17931);
xor U18230 (N_18230,N_17987,N_17881);
or U18231 (N_18231,N_17900,N_17296);
nor U18232 (N_18232,N_17318,N_17811);
nor U18233 (N_18233,N_17232,N_17486);
or U18234 (N_18234,N_17378,N_17383);
nor U18235 (N_18235,N_17023,N_17453);
or U18236 (N_18236,N_17813,N_17968);
nand U18237 (N_18237,N_17084,N_17708);
and U18238 (N_18238,N_17619,N_17174);
xnor U18239 (N_18239,N_17116,N_17487);
and U18240 (N_18240,N_17930,N_17681);
xor U18241 (N_18241,N_17217,N_17101);
or U18242 (N_18242,N_17356,N_17222);
nor U18243 (N_18243,N_17050,N_17984);
nand U18244 (N_18244,N_17814,N_17443);
or U18245 (N_18245,N_17299,N_17205);
nand U18246 (N_18246,N_17107,N_17983);
or U18247 (N_18247,N_17408,N_17426);
nand U18248 (N_18248,N_17491,N_17334);
xor U18249 (N_18249,N_17793,N_17503);
xor U18250 (N_18250,N_17462,N_17745);
nor U18251 (N_18251,N_17118,N_17332);
nand U18252 (N_18252,N_17046,N_17076);
xor U18253 (N_18253,N_17898,N_17460);
xor U18254 (N_18254,N_17466,N_17199);
xor U18255 (N_18255,N_17650,N_17950);
nand U18256 (N_18256,N_17563,N_17035);
and U18257 (N_18257,N_17583,N_17192);
nand U18258 (N_18258,N_17934,N_17304);
and U18259 (N_18259,N_17647,N_17221);
xor U18260 (N_18260,N_17246,N_17893);
and U18261 (N_18261,N_17572,N_17800);
xor U18262 (N_18262,N_17149,N_17638);
or U18263 (N_18263,N_17717,N_17233);
or U18264 (N_18264,N_17263,N_17268);
xnor U18265 (N_18265,N_17204,N_17594);
nand U18266 (N_18266,N_17728,N_17941);
or U18267 (N_18267,N_17264,N_17819);
nand U18268 (N_18268,N_17494,N_17158);
nand U18269 (N_18269,N_17917,N_17652);
nor U18270 (N_18270,N_17536,N_17341);
nand U18271 (N_18271,N_17933,N_17561);
nand U18272 (N_18272,N_17628,N_17028);
or U18273 (N_18273,N_17395,N_17816);
xor U18274 (N_18274,N_17804,N_17521);
or U18275 (N_18275,N_17458,N_17434);
nand U18276 (N_18276,N_17534,N_17200);
or U18277 (N_18277,N_17725,N_17156);
xor U18278 (N_18278,N_17859,N_17596);
nor U18279 (N_18279,N_17515,N_17848);
or U18280 (N_18280,N_17587,N_17976);
and U18281 (N_18281,N_17042,N_17615);
nand U18282 (N_18282,N_17644,N_17872);
xor U18283 (N_18283,N_17737,N_17880);
nand U18284 (N_18284,N_17935,N_17290);
nand U18285 (N_18285,N_17131,N_17079);
nor U18286 (N_18286,N_17006,N_17649);
nand U18287 (N_18287,N_17065,N_17459);
and U18288 (N_18288,N_17467,N_17889);
and U18289 (N_18289,N_17185,N_17998);
nor U18290 (N_18290,N_17809,N_17020);
or U18291 (N_18291,N_17874,N_17688);
or U18292 (N_18292,N_17518,N_17083);
or U18293 (N_18293,N_17080,N_17903);
nor U18294 (N_18294,N_17124,N_17093);
xor U18295 (N_18295,N_17741,N_17624);
or U18296 (N_18296,N_17504,N_17013);
and U18297 (N_18297,N_17856,N_17718);
nor U18298 (N_18298,N_17704,N_17643);
or U18299 (N_18299,N_17446,N_17738);
nand U18300 (N_18300,N_17215,N_17369);
or U18301 (N_18301,N_17869,N_17406);
nor U18302 (N_18302,N_17878,N_17621);
or U18303 (N_18303,N_17665,N_17249);
and U18304 (N_18304,N_17912,N_17815);
and U18305 (N_18305,N_17316,N_17805);
xnor U18306 (N_18306,N_17439,N_17776);
or U18307 (N_18307,N_17169,N_17019);
or U18308 (N_18308,N_17901,N_17085);
nor U18309 (N_18309,N_17224,N_17053);
nand U18310 (N_18310,N_17865,N_17311);
or U18311 (N_18311,N_17104,N_17582);
nand U18312 (N_18312,N_17086,N_17490);
nor U18313 (N_18313,N_17906,N_17719);
or U18314 (N_18314,N_17646,N_17393);
or U18315 (N_18315,N_17885,N_17918);
xnor U18316 (N_18316,N_17230,N_17853);
and U18317 (N_18317,N_17074,N_17139);
and U18318 (N_18318,N_17087,N_17964);
and U18319 (N_18319,N_17431,N_17618);
nand U18320 (N_18320,N_17565,N_17170);
or U18321 (N_18321,N_17986,N_17039);
xnor U18322 (N_18322,N_17022,N_17807);
xnor U18323 (N_18323,N_17274,N_17993);
nand U18324 (N_18324,N_17476,N_17732);
xor U18325 (N_18325,N_17842,N_17054);
nor U18326 (N_18326,N_17044,N_17014);
and U18327 (N_18327,N_17314,N_17225);
nand U18328 (N_18328,N_17090,N_17771);
or U18329 (N_18329,N_17913,N_17508);
and U18330 (N_18330,N_17254,N_17409);
xor U18331 (N_18331,N_17961,N_17669);
and U18332 (N_18332,N_17130,N_17833);
nor U18333 (N_18333,N_17844,N_17270);
and U18334 (N_18334,N_17666,N_17479);
xnor U18335 (N_18335,N_17907,N_17825);
or U18336 (N_18336,N_17196,N_17845);
xor U18337 (N_18337,N_17616,N_17550);
nand U18338 (N_18338,N_17435,N_17520);
nand U18339 (N_18339,N_17353,N_17972);
nor U18340 (N_18340,N_17586,N_17368);
nand U18341 (N_18341,N_17507,N_17684);
nand U18342 (N_18342,N_17277,N_17668);
and U18343 (N_18343,N_17744,N_17250);
xnor U18344 (N_18344,N_17454,N_17959);
and U18345 (N_18345,N_17276,N_17839);
or U18346 (N_18346,N_17997,N_17915);
nand U18347 (N_18347,N_17722,N_17282);
and U18348 (N_18348,N_17172,N_17401);
xnor U18349 (N_18349,N_17389,N_17716);
nand U18350 (N_18350,N_17402,N_17588);
or U18351 (N_18351,N_17936,N_17763);
or U18352 (N_18352,N_17168,N_17289);
nor U18353 (N_18353,N_17992,N_17163);
xnor U18354 (N_18354,N_17542,N_17781);
nand U18355 (N_18355,N_17866,N_17092);
nor U18356 (N_18356,N_17414,N_17351);
and U18357 (N_18357,N_17176,N_17712);
and U18358 (N_18358,N_17117,N_17821);
xor U18359 (N_18359,N_17480,N_17517);
nand U18360 (N_18360,N_17403,N_17051);
xor U18361 (N_18361,N_17243,N_17016);
and U18362 (N_18362,N_17622,N_17029);
xor U18363 (N_18363,N_17610,N_17004);
xnor U18364 (N_18364,N_17148,N_17922);
xor U18365 (N_18365,N_17297,N_17790);
xnor U18366 (N_18366,N_17656,N_17929);
and U18367 (N_18367,N_17425,N_17981);
or U18368 (N_18368,N_17788,N_17469);
and U18369 (N_18369,N_17958,N_17037);
nor U18370 (N_18370,N_17335,N_17752);
xor U18371 (N_18371,N_17723,N_17445);
or U18372 (N_18372,N_17012,N_17342);
nor U18373 (N_18373,N_17894,N_17773);
xnor U18374 (N_18374,N_17510,N_17045);
and U18375 (N_18375,N_17326,N_17284);
or U18376 (N_18376,N_17465,N_17146);
nand U18377 (N_18377,N_17584,N_17890);
xnor U18378 (N_18378,N_17639,N_17344);
xnor U18379 (N_18379,N_17121,N_17657);
or U18380 (N_18380,N_17081,N_17312);
or U18381 (N_18381,N_17327,N_17991);
nand U18382 (N_18382,N_17102,N_17496);
xor U18383 (N_18383,N_17577,N_17492);
nor U18384 (N_18384,N_17896,N_17632);
or U18385 (N_18385,N_17891,N_17835);
and U18386 (N_18386,N_17899,N_17021);
and U18387 (N_18387,N_17727,N_17810);
nor U18388 (N_18388,N_17755,N_17847);
nand U18389 (N_18389,N_17377,N_17441);
nor U18390 (N_18390,N_17468,N_17645);
xor U18391 (N_18391,N_17528,N_17059);
nor U18392 (N_18392,N_17595,N_17413);
xor U18393 (N_18393,N_17867,N_17060);
or U18394 (N_18394,N_17678,N_17484);
nand U18395 (N_18395,N_17531,N_17925);
or U18396 (N_18396,N_17129,N_17082);
or U18397 (N_18397,N_17387,N_17663);
or U18398 (N_18398,N_17173,N_17061);
nor U18399 (N_18399,N_17836,N_17911);
nor U18400 (N_18400,N_17027,N_17219);
and U18401 (N_18401,N_17071,N_17537);
and U18402 (N_18402,N_17673,N_17558);
nand U18403 (N_18403,N_17234,N_17228);
nor U18404 (N_18404,N_17258,N_17190);
and U18405 (N_18405,N_17574,N_17294);
nor U18406 (N_18406,N_17206,N_17275);
and U18407 (N_18407,N_17432,N_17034);
or U18408 (N_18408,N_17547,N_17606);
xor U18409 (N_18409,N_17599,N_17482);
nor U18410 (N_18410,N_17412,N_17756);
xnor U18411 (N_18411,N_17226,N_17191);
or U18412 (N_18412,N_17538,N_17779);
xnor U18413 (N_18413,N_17500,N_17787);
xnor U18414 (N_18414,N_17154,N_17522);
or U18415 (N_18415,N_17003,N_17614);
xnor U18416 (N_18416,N_17123,N_17955);
or U18417 (N_18417,N_17128,N_17231);
nor U18418 (N_18418,N_17309,N_17220);
or U18419 (N_18419,N_17157,N_17207);
xnor U18420 (N_18420,N_17679,N_17721);
or U18421 (N_18421,N_17830,N_17212);
nand U18422 (N_18422,N_17589,N_17526);
and U18423 (N_18423,N_17634,N_17260);
nor U18424 (N_18424,N_17612,N_17846);
or U18425 (N_18425,N_17392,N_17753);
nor U18426 (N_18426,N_17150,N_17214);
and U18427 (N_18427,N_17525,N_17026);
and U18428 (N_18428,N_17902,N_17858);
or U18429 (N_18429,N_17927,N_17442);
nor U18430 (N_18430,N_17357,N_17873);
or U18431 (N_18431,N_17937,N_17269);
nand U18432 (N_18432,N_17801,N_17391);
nand U18433 (N_18433,N_17252,N_17138);
nor U18434 (N_18434,N_17137,N_17637);
nand U18435 (N_18435,N_17861,N_17567);
or U18436 (N_18436,N_17743,N_17783);
xor U18437 (N_18437,N_17598,N_17008);
or U18438 (N_18438,N_17758,N_17198);
nand U18439 (N_18439,N_17989,N_17478);
nor U18440 (N_18440,N_17240,N_17423);
nand U18441 (N_18441,N_17448,N_17295);
nand U18442 (N_18442,N_17007,N_17768);
nand U18443 (N_18443,N_17115,N_17203);
and U18444 (N_18444,N_17949,N_17058);
and U18445 (N_18445,N_17043,N_17602);
and U18446 (N_18446,N_17928,N_17939);
and U18447 (N_18447,N_17410,N_17605);
xnor U18448 (N_18448,N_17739,N_17405);
xnor U18449 (N_18449,N_17165,N_17882);
and U18450 (N_18450,N_17100,N_17683);
xor U18451 (N_18451,N_17419,N_17791);
xnor U18452 (N_18452,N_17985,N_17374);
nor U18453 (N_18453,N_17672,N_17105);
xor U18454 (N_18454,N_17449,N_17323);
xnor U18455 (N_18455,N_17424,N_17502);
or U18456 (N_18456,N_17209,N_17095);
xor U18457 (N_18457,N_17573,N_17761);
nand U18458 (N_18458,N_17886,N_17186);
nor U18459 (N_18459,N_17108,N_17373);
nor U18460 (N_18460,N_17947,N_17211);
xor U18461 (N_18461,N_17549,N_17682);
nand U18462 (N_18462,N_17702,N_17015);
nand U18463 (N_18463,N_17760,N_17057);
and U18464 (N_18464,N_17996,N_17033);
or U18465 (N_18465,N_17119,N_17350);
nor U18466 (N_18466,N_17860,N_17519);
or U18467 (N_18467,N_17532,N_17417);
or U18468 (N_18468,N_17307,N_17770);
and U18469 (N_18469,N_17945,N_17827);
xor U18470 (N_18470,N_17238,N_17798);
nand U18471 (N_18471,N_17159,N_17360);
xor U18472 (N_18472,N_17133,N_17686);
xnor U18473 (N_18473,N_17895,N_17488);
nor U18474 (N_18474,N_17055,N_17136);
and U18475 (N_18475,N_17513,N_17315);
xnor U18476 (N_18476,N_17604,N_17164);
or U18477 (N_18477,N_17919,N_17235);
or U18478 (N_18478,N_17241,N_17229);
and U18479 (N_18479,N_17944,N_17227);
and U18480 (N_18480,N_17806,N_17184);
nand U18481 (N_18481,N_17280,N_17397);
or U18482 (N_18482,N_17548,N_17608);
xor U18483 (N_18483,N_17187,N_17817);
nor U18484 (N_18484,N_17306,N_17640);
nor U18485 (N_18485,N_17404,N_17653);
xor U18486 (N_18486,N_17471,N_17470);
xnor U18487 (N_18487,N_17477,N_17765);
nand U18488 (N_18488,N_17746,N_17111);
xnor U18489 (N_18489,N_17194,N_17524);
and U18490 (N_18490,N_17965,N_17036);
and U18491 (N_18491,N_17066,N_17049);
nor U18492 (N_18492,N_17777,N_17195);
nor U18493 (N_18493,N_17125,N_17580);
or U18494 (N_18494,N_17926,N_17461);
nand U18495 (N_18495,N_17571,N_17456);
nand U18496 (N_18496,N_17343,N_17032);
xor U18497 (N_18497,N_17994,N_17293);
or U18498 (N_18498,N_17509,N_17938);
or U18499 (N_18499,N_17385,N_17932);
or U18500 (N_18500,N_17320,N_17859);
and U18501 (N_18501,N_17668,N_17470);
xor U18502 (N_18502,N_17022,N_17071);
and U18503 (N_18503,N_17700,N_17499);
nor U18504 (N_18504,N_17309,N_17258);
or U18505 (N_18505,N_17035,N_17215);
or U18506 (N_18506,N_17760,N_17171);
and U18507 (N_18507,N_17960,N_17725);
nor U18508 (N_18508,N_17876,N_17993);
nor U18509 (N_18509,N_17206,N_17416);
xnor U18510 (N_18510,N_17498,N_17795);
xnor U18511 (N_18511,N_17711,N_17141);
or U18512 (N_18512,N_17403,N_17852);
or U18513 (N_18513,N_17606,N_17136);
nand U18514 (N_18514,N_17919,N_17700);
nand U18515 (N_18515,N_17824,N_17166);
nand U18516 (N_18516,N_17095,N_17126);
and U18517 (N_18517,N_17384,N_17029);
nand U18518 (N_18518,N_17629,N_17495);
and U18519 (N_18519,N_17786,N_17325);
and U18520 (N_18520,N_17828,N_17211);
nor U18521 (N_18521,N_17410,N_17084);
xnor U18522 (N_18522,N_17043,N_17078);
xnor U18523 (N_18523,N_17029,N_17525);
nand U18524 (N_18524,N_17175,N_17646);
nor U18525 (N_18525,N_17672,N_17209);
and U18526 (N_18526,N_17641,N_17745);
and U18527 (N_18527,N_17355,N_17962);
xor U18528 (N_18528,N_17674,N_17113);
nor U18529 (N_18529,N_17632,N_17125);
and U18530 (N_18530,N_17597,N_17607);
nor U18531 (N_18531,N_17806,N_17078);
and U18532 (N_18532,N_17584,N_17048);
xor U18533 (N_18533,N_17694,N_17407);
or U18534 (N_18534,N_17407,N_17421);
nor U18535 (N_18535,N_17281,N_17921);
nand U18536 (N_18536,N_17562,N_17136);
nor U18537 (N_18537,N_17452,N_17209);
nor U18538 (N_18538,N_17196,N_17748);
or U18539 (N_18539,N_17130,N_17192);
nor U18540 (N_18540,N_17721,N_17878);
nor U18541 (N_18541,N_17726,N_17503);
and U18542 (N_18542,N_17139,N_17286);
nor U18543 (N_18543,N_17986,N_17750);
nand U18544 (N_18544,N_17887,N_17664);
xnor U18545 (N_18545,N_17431,N_17038);
or U18546 (N_18546,N_17568,N_17032);
nand U18547 (N_18547,N_17053,N_17846);
nand U18548 (N_18548,N_17177,N_17965);
xor U18549 (N_18549,N_17645,N_17339);
nor U18550 (N_18550,N_17684,N_17061);
nor U18551 (N_18551,N_17726,N_17285);
and U18552 (N_18552,N_17487,N_17471);
nor U18553 (N_18553,N_17981,N_17198);
and U18554 (N_18554,N_17373,N_17730);
and U18555 (N_18555,N_17855,N_17006);
nand U18556 (N_18556,N_17519,N_17447);
xor U18557 (N_18557,N_17056,N_17702);
nand U18558 (N_18558,N_17259,N_17538);
or U18559 (N_18559,N_17757,N_17091);
nand U18560 (N_18560,N_17992,N_17521);
and U18561 (N_18561,N_17936,N_17436);
nor U18562 (N_18562,N_17404,N_17912);
nand U18563 (N_18563,N_17091,N_17646);
xor U18564 (N_18564,N_17810,N_17005);
xnor U18565 (N_18565,N_17130,N_17803);
or U18566 (N_18566,N_17966,N_17748);
or U18567 (N_18567,N_17918,N_17375);
xor U18568 (N_18568,N_17586,N_17598);
nor U18569 (N_18569,N_17259,N_17765);
or U18570 (N_18570,N_17474,N_17320);
or U18571 (N_18571,N_17450,N_17765);
and U18572 (N_18572,N_17970,N_17436);
or U18573 (N_18573,N_17843,N_17321);
xnor U18574 (N_18574,N_17860,N_17091);
nand U18575 (N_18575,N_17586,N_17663);
nand U18576 (N_18576,N_17928,N_17236);
or U18577 (N_18577,N_17692,N_17511);
nand U18578 (N_18578,N_17303,N_17170);
or U18579 (N_18579,N_17375,N_17388);
nand U18580 (N_18580,N_17444,N_17625);
or U18581 (N_18581,N_17767,N_17546);
nand U18582 (N_18582,N_17751,N_17518);
xnor U18583 (N_18583,N_17400,N_17623);
or U18584 (N_18584,N_17642,N_17760);
nand U18585 (N_18585,N_17174,N_17242);
or U18586 (N_18586,N_17694,N_17096);
nand U18587 (N_18587,N_17126,N_17743);
nor U18588 (N_18588,N_17498,N_17013);
nand U18589 (N_18589,N_17584,N_17984);
nor U18590 (N_18590,N_17288,N_17868);
nand U18591 (N_18591,N_17770,N_17776);
and U18592 (N_18592,N_17120,N_17436);
and U18593 (N_18593,N_17209,N_17916);
nor U18594 (N_18594,N_17334,N_17869);
xor U18595 (N_18595,N_17583,N_17208);
nand U18596 (N_18596,N_17102,N_17864);
nor U18597 (N_18597,N_17349,N_17827);
or U18598 (N_18598,N_17000,N_17072);
and U18599 (N_18599,N_17794,N_17480);
and U18600 (N_18600,N_17045,N_17422);
nand U18601 (N_18601,N_17406,N_17177);
nand U18602 (N_18602,N_17729,N_17443);
or U18603 (N_18603,N_17168,N_17791);
nand U18604 (N_18604,N_17485,N_17974);
and U18605 (N_18605,N_17851,N_17513);
nor U18606 (N_18606,N_17439,N_17292);
nor U18607 (N_18607,N_17478,N_17433);
or U18608 (N_18608,N_17532,N_17037);
nor U18609 (N_18609,N_17485,N_17593);
nand U18610 (N_18610,N_17699,N_17400);
xor U18611 (N_18611,N_17116,N_17860);
nand U18612 (N_18612,N_17937,N_17583);
nor U18613 (N_18613,N_17956,N_17768);
or U18614 (N_18614,N_17633,N_17357);
and U18615 (N_18615,N_17691,N_17586);
and U18616 (N_18616,N_17867,N_17155);
xor U18617 (N_18617,N_17796,N_17812);
and U18618 (N_18618,N_17147,N_17066);
or U18619 (N_18619,N_17459,N_17529);
or U18620 (N_18620,N_17861,N_17544);
nand U18621 (N_18621,N_17948,N_17640);
and U18622 (N_18622,N_17425,N_17034);
xor U18623 (N_18623,N_17227,N_17844);
xor U18624 (N_18624,N_17135,N_17686);
xor U18625 (N_18625,N_17495,N_17215);
nand U18626 (N_18626,N_17458,N_17422);
or U18627 (N_18627,N_17676,N_17744);
nand U18628 (N_18628,N_17376,N_17857);
and U18629 (N_18629,N_17248,N_17349);
xnor U18630 (N_18630,N_17699,N_17615);
and U18631 (N_18631,N_17547,N_17654);
nand U18632 (N_18632,N_17454,N_17057);
or U18633 (N_18633,N_17461,N_17345);
and U18634 (N_18634,N_17297,N_17914);
nor U18635 (N_18635,N_17094,N_17398);
nor U18636 (N_18636,N_17396,N_17864);
xor U18637 (N_18637,N_17507,N_17702);
or U18638 (N_18638,N_17393,N_17633);
and U18639 (N_18639,N_17995,N_17350);
and U18640 (N_18640,N_17843,N_17210);
nor U18641 (N_18641,N_17056,N_17251);
or U18642 (N_18642,N_17799,N_17018);
or U18643 (N_18643,N_17492,N_17751);
nor U18644 (N_18644,N_17329,N_17890);
nor U18645 (N_18645,N_17448,N_17205);
or U18646 (N_18646,N_17879,N_17210);
xor U18647 (N_18647,N_17459,N_17644);
xor U18648 (N_18648,N_17807,N_17763);
nand U18649 (N_18649,N_17561,N_17283);
nor U18650 (N_18650,N_17878,N_17980);
nor U18651 (N_18651,N_17980,N_17653);
and U18652 (N_18652,N_17261,N_17986);
or U18653 (N_18653,N_17675,N_17957);
nor U18654 (N_18654,N_17098,N_17893);
or U18655 (N_18655,N_17111,N_17727);
nand U18656 (N_18656,N_17691,N_17278);
nand U18657 (N_18657,N_17448,N_17334);
nand U18658 (N_18658,N_17408,N_17098);
nor U18659 (N_18659,N_17471,N_17396);
nor U18660 (N_18660,N_17050,N_17433);
nand U18661 (N_18661,N_17773,N_17634);
nand U18662 (N_18662,N_17774,N_17882);
nand U18663 (N_18663,N_17509,N_17257);
and U18664 (N_18664,N_17716,N_17415);
nand U18665 (N_18665,N_17792,N_17437);
xor U18666 (N_18666,N_17353,N_17212);
nor U18667 (N_18667,N_17235,N_17391);
or U18668 (N_18668,N_17981,N_17267);
nor U18669 (N_18669,N_17609,N_17903);
nor U18670 (N_18670,N_17656,N_17224);
and U18671 (N_18671,N_17775,N_17588);
nor U18672 (N_18672,N_17559,N_17006);
nor U18673 (N_18673,N_17210,N_17896);
nor U18674 (N_18674,N_17669,N_17505);
xnor U18675 (N_18675,N_17058,N_17425);
and U18676 (N_18676,N_17458,N_17548);
and U18677 (N_18677,N_17388,N_17363);
nand U18678 (N_18678,N_17025,N_17432);
nand U18679 (N_18679,N_17917,N_17935);
nand U18680 (N_18680,N_17154,N_17320);
nor U18681 (N_18681,N_17854,N_17727);
and U18682 (N_18682,N_17363,N_17128);
and U18683 (N_18683,N_17665,N_17355);
and U18684 (N_18684,N_17087,N_17785);
and U18685 (N_18685,N_17783,N_17129);
or U18686 (N_18686,N_17420,N_17426);
or U18687 (N_18687,N_17408,N_17031);
and U18688 (N_18688,N_17965,N_17777);
and U18689 (N_18689,N_17862,N_17950);
and U18690 (N_18690,N_17368,N_17891);
xnor U18691 (N_18691,N_17432,N_17981);
nand U18692 (N_18692,N_17728,N_17020);
nand U18693 (N_18693,N_17048,N_17743);
nor U18694 (N_18694,N_17510,N_17666);
nor U18695 (N_18695,N_17916,N_17572);
nand U18696 (N_18696,N_17230,N_17772);
xnor U18697 (N_18697,N_17505,N_17851);
xnor U18698 (N_18698,N_17780,N_17787);
or U18699 (N_18699,N_17578,N_17842);
nand U18700 (N_18700,N_17090,N_17724);
or U18701 (N_18701,N_17403,N_17374);
or U18702 (N_18702,N_17454,N_17816);
nand U18703 (N_18703,N_17477,N_17978);
or U18704 (N_18704,N_17578,N_17195);
or U18705 (N_18705,N_17756,N_17209);
or U18706 (N_18706,N_17036,N_17751);
or U18707 (N_18707,N_17736,N_17936);
nor U18708 (N_18708,N_17679,N_17374);
nand U18709 (N_18709,N_17324,N_17472);
or U18710 (N_18710,N_17283,N_17160);
xnor U18711 (N_18711,N_17242,N_17651);
and U18712 (N_18712,N_17573,N_17732);
nor U18713 (N_18713,N_17575,N_17752);
xor U18714 (N_18714,N_17123,N_17271);
or U18715 (N_18715,N_17404,N_17028);
xor U18716 (N_18716,N_17792,N_17136);
nand U18717 (N_18717,N_17608,N_17134);
nor U18718 (N_18718,N_17353,N_17271);
nand U18719 (N_18719,N_17340,N_17487);
or U18720 (N_18720,N_17764,N_17119);
or U18721 (N_18721,N_17839,N_17358);
nand U18722 (N_18722,N_17006,N_17589);
nor U18723 (N_18723,N_17976,N_17736);
nand U18724 (N_18724,N_17019,N_17961);
and U18725 (N_18725,N_17643,N_17228);
nor U18726 (N_18726,N_17674,N_17349);
and U18727 (N_18727,N_17156,N_17867);
xnor U18728 (N_18728,N_17929,N_17276);
and U18729 (N_18729,N_17657,N_17945);
xor U18730 (N_18730,N_17347,N_17249);
nand U18731 (N_18731,N_17394,N_17149);
nand U18732 (N_18732,N_17308,N_17411);
or U18733 (N_18733,N_17599,N_17230);
or U18734 (N_18734,N_17882,N_17065);
or U18735 (N_18735,N_17649,N_17091);
and U18736 (N_18736,N_17878,N_17180);
and U18737 (N_18737,N_17065,N_17067);
nor U18738 (N_18738,N_17318,N_17032);
xor U18739 (N_18739,N_17879,N_17955);
xor U18740 (N_18740,N_17977,N_17100);
nor U18741 (N_18741,N_17881,N_17063);
or U18742 (N_18742,N_17308,N_17077);
or U18743 (N_18743,N_17444,N_17936);
xor U18744 (N_18744,N_17697,N_17985);
and U18745 (N_18745,N_17306,N_17312);
and U18746 (N_18746,N_17264,N_17123);
nand U18747 (N_18747,N_17741,N_17578);
nand U18748 (N_18748,N_17775,N_17456);
and U18749 (N_18749,N_17522,N_17847);
and U18750 (N_18750,N_17098,N_17344);
nor U18751 (N_18751,N_17082,N_17228);
xnor U18752 (N_18752,N_17384,N_17904);
nand U18753 (N_18753,N_17012,N_17072);
or U18754 (N_18754,N_17908,N_17061);
and U18755 (N_18755,N_17490,N_17097);
xor U18756 (N_18756,N_17556,N_17287);
xnor U18757 (N_18757,N_17495,N_17870);
and U18758 (N_18758,N_17391,N_17217);
or U18759 (N_18759,N_17719,N_17403);
nand U18760 (N_18760,N_17077,N_17890);
nand U18761 (N_18761,N_17409,N_17968);
xnor U18762 (N_18762,N_17020,N_17825);
or U18763 (N_18763,N_17485,N_17436);
nor U18764 (N_18764,N_17430,N_17613);
nor U18765 (N_18765,N_17214,N_17617);
nand U18766 (N_18766,N_17594,N_17718);
xor U18767 (N_18767,N_17139,N_17509);
or U18768 (N_18768,N_17615,N_17349);
nand U18769 (N_18769,N_17582,N_17166);
nor U18770 (N_18770,N_17498,N_17623);
or U18771 (N_18771,N_17220,N_17473);
xnor U18772 (N_18772,N_17277,N_17070);
xnor U18773 (N_18773,N_17129,N_17548);
nand U18774 (N_18774,N_17956,N_17776);
nand U18775 (N_18775,N_17815,N_17690);
or U18776 (N_18776,N_17411,N_17412);
xnor U18777 (N_18777,N_17931,N_17815);
xnor U18778 (N_18778,N_17103,N_17755);
or U18779 (N_18779,N_17618,N_17630);
or U18780 (N_18780,N_17209,N_17726);
nor U18781 (N_18781,N_17808,N_17425);
nand U18782 (N_18782,N_17426,N_17322);
nand U18783 (N_18783,N_17314,N_17900);
nand U18784 (N_18784,N_17374,N_17253);
xnor U18785 (N_18785,N_17928,N_17349);
xor U18786 (N_18786,N_17590,N_17837);
nor U18787 (N_18787,N_17858,N_17656);
nor U18788 (N_18788,N_17290,N_17309);
and U18789 (N_18789,N_17106,N_17138);
and U18790 (N_18790,N_17972,N_17788);
nand U18791 (N_18791,N_17977,N_17114);
xnor U18792 (N_18792,N_17015,N_17128);
nor U18793 (N_18793,N_17804,N_17150);
nor U18794 (N_18794,N_17006,N_17488);
nand U18795 (N_18795,N_17914,N_17387);
or U18796 (N_18796,N_17388,N_17104);
nor U18797 (N_18797,N_17043,N_17995);
or U18798 (N_18798,N_17327,N_17776);
and U18799 (N_18799,N_17025,N_17271);
nand U18800 (N_18800,N_17600,N_17255);
xnor U18801 (N_18801,N_17454,N_17719);
nor U18802 (N_18802,N_17835,N_17458);
or U18803 (N_18803,N_17729,N_17102);
or U18804 (N_18804,N_17400,N_17548);
nor U18805 (N_18805,N_17937,N_17401);
or U18806 (N_18806,N_17805,N_17085);
nand U18807 (N_18807,N_17340,N_17413);
or U18808 (N_18808,N_17015,N_17159);
xor U18809 (N_18809,N_17690,N_17711);
or U18810 (N_18810,N_17247,N_17123);
nand U18811 (N_18811,N_17395,N_17669);
xnor U18812 (N_18812,N_17066,N_17219);
xnor U18813 (N_18813,N_17039,N_17593);
and U18814 (N_18814,N_17413,N_17616);
or U18815 (N_18815,N_17537,N_17884);
xnor U18816 (N_18816,N_17239,N_17821);
xor U18817 (N_18817,N_17709,N_17436);
nand U18818 (N_18818,N_17002,N_17630);
and U18819 (N_18819,N_17270,N_17160);
nor U18820 (N_18820,N_17998,N_17687);
and U18821 (N_18821,N_17314,N_17375);
nand U18822 (N_18822,N_17078,N_17005);
and U18823 (N_18823,N_17065,N_17203);
and U18824 (N_18824,N_17826,N_17731);
and U18825 (N_18825,N_17565,N_17420);
or U18826 (N_18826,N_17429,N_17321);
and U18827 (N_18827,N_17898,N_17545);
nor U18828 (N_18828,N_17632,N_17750);
nor U18829 (N_18829,N_17195,N_17635);
or U18830 (N_18830,N_17418,N_17104);
nand U18831 (N_18831,N_17671,N_17753);
and U18832 (N_18832,N_17309,N_17064);
and U18833 (N_18833,N_17533,N_17949);
or U18834 (N_18834,N_17446,N_17943);
nand U18835 (N_18835,N_17040,N_17748);
nor U18836 (N_18836,N_17488,N_17042);
or U18837 (N_18837,N_17019,N_17101);
nor U18838 (N_18838,N_17434,N_17138);
xnor U18839 (N_18839,N_17209,N_17189);
and U18840 (N_18840,N_17495,N_17719);
xor U18841 (N_18841,N_17573,N_17131);
or U18842 (N_18842,N_17783,N_17033);
xnor U18843 (N_18843,N_17463,N_17225);
xor U18844 (N_18844,N_17182,N_17120);
xnor U18845 (N_18845,N_17246,N_17393);
nand U18846 (N_18846,N_17494,N_17066);
and U18847 (N_18847,N_17159,N_17466);
or U18848 (N_18848,N_17579,N_17069);
nand U18849 (N_18849,N_17475,N_17410);
nor U18850 (N_18850,N_17100,N_17671);
nand U18851 (N_18851,N_17116,N_17405);
xnor U18852 (N_18852,N_17976,N_17288);
xnor U18853 (N_18853,N_17037,N_17237);
nor U18854 (N_18854,N_17379,N_17441);
nor U18855 (N_18855,N_17963,N_17660);
nand U18856 (N_18856,N_17235,N_17991);
and U18857 (N_18857,N_17041,N_17355);
nor U18858 (N_18858,N_17300,N_17284);
nand U18859 (N_18859,N_17702,N_17063);
and U18860 (N_18860,N_17003,N_17452);
xnor U18861 (N_18861,N_17243,N_17770);
nand U18862 (N_18862,N_17197,N_17685);
nor U18863 (N_18863,N_17091,N_17353);
xor U18864 (N_18864,N_17000,N_17741);
xnor U18865 (N_18865,N_17915,N_17118);
nor U18866 (N_18866,N_17633,N_17564);
and U18867 (N_18867,N_17372,N_17624);
xor U18868 (N_18868,N_17167,N_17454);
nand U18869 (N_18869,N_17487,N_17159);
nor U18870 (N_18870,N_17887,N_17707);
nor U18871 (N_18871,N_17164,N_17419);
nand U18872 (N_18872,N_17094,N_17870);
and U18873 (N_18873,N_17211,N_17226);
xor U18874 (N_18874,N_17726,N_17718);
and U18875 (N_18875,N_17340,N_17924);
or U18876 (N_18876,N_17662,N_17107);
nor U18877 (N_18877,N_17008,N_17319);
xnor U18878 (N_18878,N_17218,N_17346);
and U18879 (N_18879,N_17076,N_17372);
nor U18880 (N_18880,N_17232,N_17208);
nor U18881 (N_18881,N_17683,N_17295);
nor U18882 (N_18882,N_17248,N_17555);
nand U18883 (N_18883,N_17265,N_17367);
or U18884 (N_18884,N_17688,N_17323);
or U18885 (N_18885,N_17608,N_17942);
nor U18886 (N_18886,N_17545,N_17596);
nand U18887 (N_18887,N_17693,N_17218);
nor U18888 (N_18888,N_17601,N_17895);
and U18889 (N_18889,N_17677,N_17067);
nand U18890 (N_18890,N_17175,N_17489);
xnor U18891 (N_18891,N_17867,N_17722);
or U18892 (N_18892,N_17149,N_17468);
and U18893 (N_18893,N_17494,N_17399);
and U18894 (N_18894,N_17276,N_17283);
and U18895 (N_18895,N_17808,N_17861);
and U18896 (N_18896,N_17719,N_17455);
nor U18897 (N_18897,N_17183,N_17051);
nand U18898 (N_18898,N_17427,N_17065);
xor U18899 (N_18899,N_17119,N_17308);
or U18900 (N_18900,N_17449,N_17055);
or U18901 (N_18901,N_17567,N_17271);
nand U18902 (N_18902,N_17525,N_17249);
and U18903 (N_18903,N_17215,N_17537);
nand U18904 (N_18904,N_17236,N_17516);
nand U18905 (N_18905,N_17203,N_17233);
xor U18906 (N_18906,N_17373,N_17134);
xor U18907 (N_18907,N_17976,N_17595);
and U18908 (N_18908,N_17333,N_17135);
nand U18909 (N_18909,N_17407,N_17371);
or U18910 (N_18910,N_17463,N_17866);
and U18911 (N_18911,N_17097,N_17570);
or U18912 (N_18912,N_17344,N_17564);
nand U18913 (N_18913,N_17212,N_17922);
xor U18914 (N_18914,N_17410,N_17442);
xnor U18915 (N_18915,N_17032,N_17588);
xor U18916 (N_18916,N_17018,N_17839);
or U18917 (N_18917,N_17557,N_17131);
or U18918 (N_18918,N_17116,N_17409);
xnor U18919 (N_18919,N_17854,N_17785);
nand U18920 (N_18920,N_17226,N_17591);
xnor U18921 (N_18921,N_17533,N_17726);
xor U18922 (N_18922,N_17039,N_17434);
xnor U18923 (N_18923,N_17289,N_17114);
nand U18924 (N_18924,N_17269,N_17451);
nor U18925 (N_18925,N_17646,N_17271);
nor U18926 (N_18926,N_17792,N_17766);
or U18927 (N_18927,N_17090,N_17327);
nand U18928 (N_18928,N_17380,N_17732);
or U18929 (N_18929,N_17431,N_17690);
nand U18930 (N_18930,N_17860,N_17807);
xnor U18931 (N_18931,N_17683,N_17889);
nand U18932 (N_18932,N_17247,N_17284);
or U18933 (N_18933,N_17079,N_17928);
nand U18934 (N_18934,N_17404,N_17505);
nor U18935 (N_18935,N_17526,N_17310);
and U18936 (N_18936,N_17575,N_17319);
and U18937 (N_18937,N_17041,N_17205);
and U18938 (N_18938,N_17617,N_17650);
nand U18939 (N_18939,N_17754,N_17125);
nand U18940 (N_18940,N_17840,N_17970);
nor U18941 (N_18941,N_17729,N_17222);
nor U18942 (N_18942,N_17193,N_17328);
nand U18943 (N_18943,N_17835,N_17913);
xnor U18944 (N_18944,N_17357,N_17829);
or U18945 (N_18945,N_17273,N_17038);
nor U18946 (N_18946,N_17728,N_17268);
xnor U18947 (N_18947,N_17758,N_17348);
nor U18948 (N_18948,N_17248,N_17565);
xnor U18949 (N_18949,N_17220,N_17192);
nand U18950 (N_18950,N_17059,N_17840);
or U18951 (N_18951,N_17000,N_17287);
or U18952 (N_18952,N_17934,N_17791);
nand U18953 (N_18953,N_17836,N_17553);
and U18954 (N_18954,N_17923,N_17320);
nand U18955 (N_18955,N_17566,N_17997);
xnor U18956 (N_18956,N_17465,N_17885);
and U18957 (N_18957,N_17565,N_17697);
nor U18958 (N_18958,N_17606,N_17067);
or U18959 (N_18959,N_17982,N_17171);
and U18960 (N_18960,N_17268,N_17030);
or U18961 (N_18961,N_17203,N_17298);
and U18962 (N_18962,N_17116,N_17591);
nand U18963 (N_18963,N_17999,N_17000);
xor U18964 (N_18964,N_17955,N_17978);
or U18965 (N_18965,N_17511,N_17175);
and U18966 (N_18966,N_17091,N_17982);
and U18967 (N_18967,N_17727,N_17034);
nand U18968 (N_18968,N_17357,N_17355);
xor U18969 (N_18969,N_17901,N_17113);
nand U18970 (N_18970,N_17059,N_17677);
xor U18971 (N_18971,N_17001,N_17977);
nor U18972 (N_18972,N_17273,N_17491);
nor U18973 (N_18973,N_17240,N_17384);
and U18974 (N_18974,N_17821,N_17496);
or U18975 (N_18975,N_17398,N_17952);
nor U18976 (N_18976,N_17667,N_17479);
or U18977 (N_18977,N_17775,N_17418);
nor U18978 (N_18978,N_17639,N_17979);
or U18979 (N_18979,N_17858,N_17595);
and U18980 (N_18980,N_17677,N_17334);
nor U18981 (N_18981,N_17883,N_17864);
nand U18982 (N_18982,N_17187,N_17522);
xnor U18983 (N_18983,N_17440,N_17855);
nand U18984 (N_18984,N_17304,N_17736);
and U18985 (N_18985,N_17845,N_17847);
or U18986 (N_18986,N_17710,N_17052);
and U18987 (N_18987,N_17855,N_17349);
or U18988 (N_18988,N_17867,N_17472);
or U18989 (N_18989,N_17102,N_17609);
or U18990 (N_18990,N_17380,N_17942);
or U18991 (N_18991,N_17149,N_17751);
nand U18992 (N_18992,N_17180,N_17630);
nor U18993 (N_18993,N_17046,N_17554);
nand U18994 (N_18994,N_17372,N_17307);
or U18995 (N_18995,N_17989,N_17057);
and U18996 (N_18996,N_17972,N_17841);
and U18997 (N_18997,N_17961,N_17994);
xnor U18998 (N_18998,N_17380,N_17362);
or U18999 (N_18999,N_17101,N_17191);
xor U19000 (N_19000,N_18276,N_18950);
xnor U19001 (N_19001,N_18663,N_18130);
nand U19002 (N_19002,N_18622,N_18713);
or U19003 (N_19003,N_18913,N_18348);
xnor U19004 (N_19004,N_18387,N_18956);
or U19005 (N_19005,N_18820,N_18584);
nor U19006 (N_19006,N_18855,N_18808);
xor U19007 (N_19007,N_18044,N_18813);
nor U19008 (N_19008,N_18408,N_18945);
nor U19009 (N_19009,N_18843,N_18932);
nor U19010 (N_19010,N_18780,N_18299);
nand U19011 (N_19011,N_18419,N_18682);
nand U19012 (N_19012,N_18402,N_18849);
xnor U19013 (N_19013,N_18546,N_18582);
and U19014 (N_19014,N_18952,N_18592);
or U19015 (N_19015,N_18258,N_18962);
and U19016 (N_19016,N_18026,N_18119);
nor U19017 (N_19017,N_18372,N_18772);
nand U19018 (N_19018,N_18756,N_18303);
or U19019 (N_19019,N_18465,N_18696);
and U19020 (N_19020,N_18729,N_18087);
nand U19021 (N_19021,N_18146,N_18115);
nor U19022 (N_19022,N_18982,N_18242);
and U19023 (N_19023,N_18291,N_18818);
or U19024 (N_19024,N_18651,N_18840);
and U19025 (N_19025,N_18685,N_18270);
nand U19026 (N_19026,N_18286,N_18412);
and U19027 (N_19027,N_18698,N_18309);
or U19028 (N_19028,N_18920,N_18344);
nor U19029 (N_19029,N_18243,N_18445);
nand U19030 (N_19030,N_18547,N_18172);
nor U19031 (N_19031,N_18190,N_18846);
nor U19032 (N_19032,N_18197,N_18174);
and U19033 (N_19033,N_18168,N_18569);
and U19034 (N_19034,N_18899,N_18295);
and U19035 (N_19035,N_18936,N_18759);
or U19036 (N_19036,N_18211,N_18666);
xor U19037 (N_19037,N_18548,N_18779);
nand U19038 (N_19038,N_18004,N_18154);
nand U19039 (N_19039,N_18804,N_18383);
or U19040 (N_19040,N_18178,N_18097);
and U19041 (N_19041,N_18330,N_18468);
nor U19042 (N_19042,N_18252,N_18807);
nor U19043 (N_19043,N_18667,N_18356);
nand U19044 (N_19044,N_18156,N_18124);
nand U19045 (N_19045,N_18618,N_18670);
nand U19046 (N_19046,N_18429,N_18748);
or U19047 (N_19047,N_18781,N_18838);
or U19048 (N_19048,N_18885,N_18436);
nor U19049 (N_19049,N_18239,N_18283);
xnor U19050 (N_19050,N_18016,N_18727);
nand U19051 (N_19051,N_18300,N_18037);
or U19052 (N_19052,N_18559,N_18615);
nor U19053 (N_19053,N_18915,N_18598);
nor U19054 (N_19054,N_18573,N_18790);
and U19055 (N_19055,N_18607,N_18560);
nor U19056 (N_19056,N_18223,N_18543);
xnor U19057 (N_19057,N_18416,N_18399);
nor U19058 (N_19058,N_18853,N_18531);
nor U19059 (N_19059,N_18268,N_18279);
nor U19060 (N_19060,N_18870,N_18029);
nor U19061 (N_19061,N_18984,N_18555);
or U19062 (N_19062,N_18410,N_18095);
nor U19063 (N_19063,N_18453,N_18481);
and U19064 (N_19064,N_18933,N_18654);
nor U19065 (N_19065,N_18695,N_18248);
or U19066 (N_19066,N_18032,N_18972);
xnor U19067 (N_19067,N_18040,N_18381);
and U19068 (N_19068,N_18264,N_18414);
and U19069 (N_19069,N_18035,N_18477);
and U19070 (N_19070,N_18726,N_18519);
and U19071 (N_19071,N_18633,N_18626);
and U19072 (N_19072,N_18407,N_18676);
nor U19073 (N_19073,N_18024,N_18385);
xor U19074 (N_19074,N_18832,N_18802);
xor U19075 (N_19075,N_18012,N_18861);
nand U19076 (N_19076,N_18882,N_18486);
nor U19077 (N_19077,N_18942,N_18072);
xnor U19078 (N_19078,N_18908,N_18485);
xnor U19079 (N_19079,N_18280,N_18856);
and U19080 (N_19080,N_18815,N_18467);
nor U19081 (N_19081,N_18176,N_18823);
xnor U19082 (N_19082,N_18306,N_18020);
and U19083 (N_19083,N_18100,N_18451);
nor U19084 (N_19084,N_18162,N_18672);
xnor U19085 (N_19085,N_18123,N_18597);
nand U19086 (N_19086,N_18331,N_18797);
xor U19087 (N_19087,N_18686,N_18585);
nor U19088 (N_19088,N_18620,N_18139);
xor U19089 (N_19089,N_18549,N_18730);
xor U19090 (N_19090,N_18805,N_18974);
or U19091 (N_19091,N_18322,N_18014);
nand U19092 (N_19092,N_18221,N_18085);
or U19093 (N_19093,N_18151,N_18702);
xor U19094 (N_19094,N_18693,N_18909);
nand U19095 (N_19095,N_18938,N_18432);
nor U19096 (N_19096,N_18939,N_18405);
nand U19097 (N_19097,N_18267,N_18217);
nand U19098 (N_19098,N_18164,N_18593);
nand U19099 (N_19099,N_18017,N_18732);
nand U19100 (N_19100,N_18629,N_18490);
nor U19101 (N_19101,N_18621,N_18006);
and U19102 (N_19102,N_18210,N_18128);
nand U19103 (N_19103,N_18250,N_18894);
nand U19104 (N_19104,N_18858,N_18112);
nor U19105 (N_19105,N_18589,N_18194);
and U19106 (N_19106,N_18200,N_18101);
and U19107 (N_19107,N_18567,N_18346);
xnor U19108 (N_19108,N_18137,N_18981);
nand U19109 (N_19109,N_18627,N_18262);
or U19110 (N_19110,N_18062,N_18284);
nand U19111 (N_19111,N_18246,N_18463);
nor U19112 (N_19112,N_18249,N_18752);
or U19113 (N_19113,N_18235,N_18988);
nand U19114 (N_19114,N_18049,N_18817);
nand U19115 (N_19115,N_18907,N_18997);
or U19116 (N_19116,N_18515,N_18134);
nand U19117 (N_19117,N_18192,N_18561);
xnor U19118 (N_19118,N_18970,N_18077);
or U19119 (N_19119,N_18275,N_18847);
and U19120 (N_19120,N_18539,N_18055);
nand U19121 (N_19121,N_18816,N_18579);
nor U19122 (N_19122,N_18812,N_18528);
nand U19123 (N_19123,N_18425,N_18161);
xor U19124 (N_19124,N_18260,N_18364);
xor U19125 (N_19125,N_18513,N_18347);
and U19126 (N_19126,N_18810,N_18389);
or U19127 (N_19127,N_18000,N_18552);
or U19128 (N_19128,N_18835,N_18879);
and U19129 (N_19129,N_18891,N_18059);
and U19130 (N_19130,N_18900,N_18571);
and U19131 (N_19131,N_18664,N_18472);
or U19132 (N_19132,N_18771,N_18056);
nor U19133 (N_19133,N_18450,N_18799);
nand U19134 (N_19134,N_18474,N_18526);
nor U19135 (N_19135,N_18136,N_18341);
nor U19136 (N_19136,N_18669,N_18253);
and U19137 (N_19137,N_18690,N_18761);
xnor U19138 (N_19138,N_18090,N_18011);
or U19139 (N_19139,N_18483,N_18814);
nor U19140 (N_19140,N_18061,N_18166);
or U19141 (N_19141,N_18632,N_18129);
nor U19142 (N_19142,N_18083,N_18784);
or U19143 (N_19143,N_18754,N_18464);
and U19144 (N_19144,N_18329,N_18321);
nor U19145 (N_19145,N_18359,N_18715);
nand U19146 (N_19146,N_18497,N_18271);
nor U19147 (N_19147,N_18118,N_18707);
nand U19148 (N_19148,N_18132,N_18826);
nor U19149 (N_19149,N_18883,N_18070);
xnor U19150 (N_19150,N_18914,N_18471);
xor U19151 (N_19151,N_18825,N_18947);
or U19152 (N_19152,N_18876,N_18550);
xor U19153 (N_19153,N_18488,N_18117);
xnor U19154 (N_19154,N_18437,N_18655);
and U19155 (N_19155,N_18403,N_18110);
and U19156 (N_19156,N_18426,N_18860);
or U19157 (N_19157,N_18638,N_18206);
nor U19158 (N_19158,N_18159,N_18082);
nor U19159 (N_19159,N_18142,N_18700);
nor U19160 (N_19160,N_18841,N_18520);
xor U19161 (N_19161,N_18367,N_18361);
xnor U19162 (N_19162,N_18209,N_18019);
xnor U19163 (N_19163,N_18743,N_18572);
nor U19164 (N_19164,N_18863,N_18525);
xnor U19165 (N_19165,N_18506,N_18677);
xnor U19166 (N_19166,N_18340,N_18563);
nor U19167 (N_19167,N_18358,N_18500);
xnor U19168 (N_19168,N_18999,N_18254);
and U19169 (N_19169,N_18601,N_18777);
nand U19170 (N_19170,N_18643,N_18639);
and U19171 (N_19171,N_18333,N_18368);
nor U19172 (N_19172,N_18522,N_18189);
and U19173 (N_19173,N_18917,N_18111);
nand U19174 (N_19174,N_18951,N_18187);
and U19175 (N_19175,N_18155,N_18762);
or U19176 (N_19176,N_18971,N_18991);
or U19177 (N_19177,N_18386,N_18328);
or U19178 (N_19178,N_18739,N_18527);
or U19179 (N_19179,N_18599,N_18921);
or U19180 (N_19180,N_18273,N_18502);
and U19181 (N_19181,N_18302,N_18764);
nor U19182 (N_19182,N_18398,N_18296);
nor U19183 (N_19183,N_18957,N_18628);
nor U19184 (N_19184,N_18048,N_18400);
nand U19185 (N_19185,N_18157,N_18516);
or U19186 (N_19186,N_18930,N_18791);
nand U19187 (N_19187,N_18094,N_18641);
or U19188 (N_19188,N_18940,N_18948);
or U19189 (N_19189,N_18418,N_18766);
xor U19190 (N_19190,N_18769,N_18692);
or U19191 (N_19191,N_18906,N_18278);
nand U19192 (N_19192,N_18529,N_18365);
xor U19193 (N_19193,N_18986,N_18173);
nand U19194 (N_19194,N_18524,N_18204);
xor U19195 (N_19195,N_18057,N_18396);
xnor U19196 (N_19196,N_18659,N_18750);
nor U19197 (N_19197,N_18503,N_18728);
or U19198 (N_19198,N_18377,N_18184);
nor U19199 (N_19199,N_18648,N_18711);
or U19200 (N_19200,N_18521,N_18541);
xnor U19201 (N_19201,N_18493,N_18872);
xnor U19202 (N_19202,N_18587,N_18596);
and U19203 (N_19203,N_18195,N_18536);
nor U19204 (N_19204,N_18047,N_18289);
or U19205 (N_19205,N_18179,N_18535);
or U19206 (N_19206,N_18312,N_18786);
and U19207 (N_19207,N_18874,N_18152);
nor U19208 (N_19208,N_18723,N_18442);
nand U19209 (N_19209,N_18763,N_18869);
or U19210 (N_19210,N_18379,N_18255);
nor U19211 (N_19211,N_18608,N_18343);
nor U19212 (N_19212,N_18308,N_18036);
nor U19213 (N_19213,N_18964,N_18455);
or U19214 (N_19214,N_18704,N_18580);
nor U19215 (N_19215,N_18866,N_18323);
xor U19216 (N_19216,N_18351,N_18916);
or U19217 (N_19217,N_18339,N_18602);
nand U19218 (N_19218,N_18148,N_18269);
xor U19219 (N_19219,N_18673,N_18903);
and U19220 (N_19220,N_18009,N_18694);
nand U19221 (N_19221,N_18583,N_18697);
nand U19222 (N_19222,N_18272,N_18392);
nand U19223 (N_19223,N_18898,N_18332);
and U19224 (N_19224,N_18852,N_18979);
or U19225 (N_19225,N_18509,N_18327);
nor U19226 (N_19226,N_18428,N_18479);
nand U19227 (N_19227,N_18033,N_18795);
and U19228 (N_19228,N_18363,N_18145);
xor U19229 (N_19229,N_18191,N_18050);
nor U19230 (N_19230,N_18357,N_18417);
xor U19231 (N_19231,N_18540,N_18043);
nand U19232 (N_19232,N_18232,N_18301);
nand U19233 (N_19233,N_18030,N_18274);
xnor U19234 (N_19234,N_18440,N_18041);
or U19235 (N_19235,N_18240,N_18227);
nor U19236 (N_19236,N_18746,N_18985);
or U19237 (N_19237,N_18738,N_18466);
or U19238 (N_19238,N_18706,N_18758);
and U19239 (N_19239,N_18510,N_18806);
and U19240 (N_19240,N_18645,N_18158);
nor U19241 (N_19241,N_18703,N_18975);
or U19242 (N_19242,N_18581,N_18067);
nand U19243 (N_19243,N_18625,N_18027);
nor U19244 (N_19244,N_18656,N_18219);
nor U19245 (N_19245,N_18782,N_18845);
xor U19246 (N_19246,N_18236,N_18238);
and U19247 (N_19247,N_18013,N_18220);
or U19248 (N_19248,N_18051,N_18514);
nor U19249 (N_19249,N_18353,N_18718);
xnor U19250 (N_19250,N_18338,N_18811);
or U19251 (N_19251,N_18427,N_18854);
nand U19252 (N_19252,N_18096,N_18864);
xnor U19253 (N_19253,N_18456,N_18224);
nand U19254 (N_19254,N_18836,N_18411);
and U19255 (N_19255,N_18028,N_18491);
nand U19256 (N_19256,N_18366,N_18919);
or U19257 (N_19257,N_18544,N_18889);
nand U19258 (N_19258,N_18709,N_18773);
xnor U19259 (N_19259,N_18153,N_18753);
nand U19260 (N_19260,N_18065,N_18188);
nor U19261 (N_19261,N_18943,N_18183);
nand U19262 (N_19262,N_18310,N_18325);
xnor U19263 (N_19263,N_18298,N_18937);
nor U19264 (N_19264,N_18994,N_18446);
nor U19265 (N_19265,N_18449,N_18231);
nor U19266 (N_19266,N_18447,N_18701);
nor U19267 (N_19267,N_18577,N_18617);
and U19268 (N_19268,N_18360,N_18207);
or U19269 (N_19269,N_18163,N_18409);
nor U19270 (N_19270,N_18212,N_18553);
or U19271 (N_19271,N_18996,N_18538);
and U19272 (N_19272,N_18180,N_18518);
and U19273 (N_19273,N_18570,N_18104);
or U19274 (N_19274,N_18084,N_18614);
xor U19275 (N_19275,N_18661,N_18990);
or U19276 (N_19276,N_18494,N_18053);
and U19277 (N_19277,N_18609,N_18324);
nor U19278 (N_19278,N_18473,N_18005);
xnor U19279 (N_19279,N_18292,N_18925);
or U19280 (N_19280,N_18722,N_18443);
xor U19281 (N_19281,N_18193,N_18993);
or U19282 (N_19282,N_18374,N_18650);
and U19283 (N_19283,N_18218,N_18431);
nand U19284 (N_19284,N_18452,N_18944);
and U19285 (N_19285,N_18966,N_18557);
and U19286 (N_19286,N_18868,N_18896);
xor U19287 (N_19287,N_18352,N_18042);
and U19288 (N_19288,N_18565,N_18109);
or U19289 (N_19289,N_18106,N_18684);
xnor U19290 (N_19290,N_18745,N_18125);
nor U19291 (N_19291,N_18839,N_18430);
xnor U19292 (N_19292,N_18316,N_18665);
nor U19293 (N_19293,N_18169,N_18165);
xor U19294 (N_19294,N_18380,N_18116);
and U19295 (N_19295,N_18079,N_18370);
xnor U19296 (N_19296,N_18736,N_18147);
and U19297 (N_19297,N_18216,N_18778);
xnor U19298 (N_19298,N_18294,N_18992);
nor U19299 (N_19299,N_18963,N_18545);
nor U19300 (N_19300,N_18422,N_18681);
or U19301 (N_19301,N_18658,N_18444);
and U19302 (N_19302,N_18122,N_18788);
xnor U19303 (N_19303,N_18261,N_18613);
nor U19304 (N_19304,N_18562,N_18895);
and U19305 (N_19305,N_18099,N_18058);
xnor U19306 (N_19306,N_18803,N_18604);
and U19307 (N_19307,N_18901,N_18965);
or U19308 (N_19308,N_18461,N_18143);
or U19309 (N_19309,N_18198,N_18391);
xor U19310 (N_19310,N_18955,N_18499);
or U19311 (N_19311,N_18091,N_18290);
or U19312 (N_19312,N_18244,N_18987);
and U19313 (N_19313,N_18317,N_18859);
and U19314 (N_19314,N_18848,N_18657);
xnor U19315 (N_19315,N_18588,N_18025);
xnor U19316 (N_19316,N_18354,N_18470);
nand U19317 (N_19317,N_18458,N_18285);
or U19318 (N_19318,N_18404,N_18423);
nand U19319 (N_19319,N_18133,N_18844);
xnor U19320 (N_19320,N_18566,N_18420);
and U19321 (N_19321,N_18765,N_18946);
nor U19322 (N_19322,N_18460,N_18576);
nor U19323 (N_19323,N_18086,N_18287);
and U19324 (N_19324,N_18749,N_18787);
or U19325 (N_19325,N_18755,N_18710);
or U19326 (N_19326,N_18371,N_18640);
and U19327 (N_19327,N_18785,N_18740);
nand U19328 (N_19328,N_18689,N_18837);
nor U19329 (N_19329,N_18482,N_18871);
nand U19330 (N_19330,N_18653,N_18171);
nor U19331 (N_19331,N_18021,N_18792);
and U19332 (N_19332,N_18475,N_18880);
and U19333 (N_19333,N_18735,N_18929);
xnor U19334 (N_19334,N_18498,N_18731);
xor U19335 (N_19335,N_18649,N_18114);
nor U19336 (N_19336,N_18744,N_18088);
and U19337 (N_19337,N_18237,N_18413);
or U19338 (N_19338,N_18480,N_18010);
nand U19339 (N_19339,N_18893,N_18318);
nand U19340 (N_19340,N_18045,N_18362);
and U19341 (N_19341,N_18789,N_18725);
and U19342 (N_19342,N_18245,N_18623);
and U19343 (N_19343,N_18060,N_18668);
xnor U19344 (N_19344,N_18074,N_18958);
and U19345 (N_19345,N_18108,N_18307);
nand U19346 (N_19346,N_18135,N_18205);
or U19347 (N_19347,N_18186,N_18679);
nand U19348 (N_19348,N_18454,N_18532);
nor U19349 (N_19349,N_18199,N_18591);
xnor U19350 (N_19350,N_18107,N_18478);
nand U19351 (N_19351,N_18507,N_18170);
or U19352 (N_19352,N_18378,N_18918);
nand U19353 (N_19353,N_18234,N_18213);
nor U19354 (N_19354,N_18926,N_18675);
nand U19355 (N_19355,N_18796,N_18078);
nor U19356 (N_19356,N_18001,N_18202);
and U19357 (N_19357,N_18487,N_18121);
nor U19358 (N_19358,N_18336,N_18716);
xnor U19359 (N_19359,N_18031,N_18022);
nand U19360 (N_19360,N_18138,N_18505);
or U19361 (N_19361,N_18523,N_18558);
and U19362 (N_19362,N_18511,N_18822);
nor U19363 (N_19363,N_18457,N_18611);
or U19364 (N_19364,N_18492,N_18757);
nand U19365 (N_19365,N_18610,N_18081);
and U19366 (N_19366,N_18433,N_18369);
and U19367 (N_19367,N_18897,N_18978);
or U19368 (N_19368,N_18827,N_18373);
nor U19369 (N_19369,N_18304,N_18092);
nand U19370 (N_19370,N_18181,N_18071);
nor U19371 (N_19371,N_18508,N_18724);
or U19372 (N_19372,N_18144,N_18717);
or U19373 (N_19373,N_18265,N_18421);
and U19374 (N_19374,N_18594,N_18862);
xnor U19375 (N_19375,N_18415,N_18530);
and U19376 (N_19376,N_18439,N_18688);
and U19377 (N_19377,N_18742,N_18105);
or U19378 (N_19378,N_18881,N_18644);
nor U19379 (N_19379,N_18969,N_18120);
or U19380 (N_19380,N_18127,N_18865);
nor U19381 (N_19381,N_18647,N_18911);
xnor U19382 (N_19382,N_18775,N_18564);
xor U19383 (N_19383,N_18927,N_18424);
or U19384 (N_19384,N_18662,N_18770);
or U19385 (N_19385,N_18683,N_18397);
xor U19386 (N_19386,N_18800,N_18630);
xor U19387 (N_19387,N_18281,N_18721);
nor U19388 (N_19388,N_18241,N_18448);
nand U19389 (N_19389,N_18185,N_18039);
nand U19390 (N_19390,N_18819,N_18293);
xor U19391 (N_19391,N_18953,N_18884);
nor U19392 (N_19392,N_18776,N_18674);
xor U19393 (N_19393,N_18834,N_18063);
and U19394 (N_19394,N_18912,N_18406);
nand U19395 (N_19395,N_18828,N_18489);
and U19396 (N_19396,N_18976,N_18680);
or U19397 (N_19397,N_18501,N_18315);
or U19398 (N_19398,N_18297,N_18222);
nand U19399 (N_19399,N_18435,N_18496);
xnor U19400 (N_19400,N_18355,N_18646);
nor U19401 (N_19401,N_18968,N_18233);
xnor U19402 (N_19402,N_18829,N_18103);
or U19403 (N_19403,N_18983,N_18113);
nor U19404 (N_19404,N_18208,N_18830);
and U19405 (N_19405,N_18652,N_18388);
nand U19406 (N_19406,N_18660,N_18305);
nor U19407 (N_19407,N_18708,N_18612);
xor U19408 (N_19408,N_18783,N_18619);
nand U19409 (N_19409,N_18801,N_18551);
nor U19410 (N_19410,N_18228,N_18175);
or U19411 (N_19411,N_18384,N_18935);
nor U19412 (N_19412,N_18995,N_18824);
or U19413 (N_19413,N_18326,N_18636);
nand U19414 (N_19414,N_18977,N_18393);
nand U19415 (N_19415,N_18687,N_18167);
or U19416 (N_19416,N_18314,N_18214);
or U19417 (N_19417,N_18038,N_18476);
nor U19418 (N_19418,N_18605,N_18052);
xnor U19419 (N_19419,N_18046,N_18504);
nand U19420 (N_19420,N_18247,N_18034);
nor U19421 (N_19421,N_18350,N_18705);
xor U19422 (N_19422,N_18998,N_18699);
nor U19423 (N_19423,N_18512,N_18229);
and U19424 (N_19424,N_18959,N_18961);
and U19425 (N_19425,N_18905,N_18018);
nor U19426 (N_19426,N_18334,N_18631);
and U19427 (N_19427,N_18642,N_18578);
nor U19428 (N_19428,N_18747,N_18934);
or U19429 (N_19429,N_18989,N_18311);
xor U19430 (N_19430,N_18401,N_18691);
nand U19431 (N_19431,N_18225,N_18556);
and U19432 (N_19432,N_18678,N_18141);
xor U19433 (N_19433,N_18886,N_18201);
nor U19434 (N_19434,N_18266,N_18712);
xor U19435 (N_19435,N_18313,N_18973);
nand U19436 (N_19436,N_18089,N_18980);
nor U19437 (N_19437,N_18928,N_18337);
nor U19438 (N_19438,N_18634,N_18850);
nor U19439 (N_19439,N_18542,N_18767);
nand U19440 (N_19440,N_18960,N_18586);
and U19441 (N_19441,N_18177,N_18438);
nor U19442 (N_19442,N_18590,N_18008);
and U19443 (N_19443,N_18434,N_18595);
nand U19444 (N_19444,N_18093,N_18954);
or U19445 (N_19445,N_18887,N_18878);
nand U19446 (N_19446,N_18517,N_18320);
xor U19447 (N_19447,N_18831,N_18149);
or U19448 (N_19448,N_18066,N_18751);
nand U19449 (N_19449,N_18537,N_18288);
nor U19450 (N_19450,N_18263,N_18459);
and U19451 (N_19451,N_18256,N_18714);
and U19452 (N_19452,N_18534,N_18875);
nor U19453 (N_19453,N_18098,N_18888);
and U19454 (N_19454,N_18857,N_18259);
and U19455 (N_19455,N_18080,N_18568);
nand U19456 (N_19456,N_18890,N_18719);
xor U19457 (N_19457,N_18382,N_18734);
or U19458 (N_19458,N_18904,N_18203);
and U19459 (N_19459,N_18603,N_18574);
xor U19460 (N_19460,N_18335,N_18064);
and U19461 (N_19461,N_18150,N_18635);
and U19462 (N_19462,N_18922,N_18923);
nor U19463 (N_19463,N_18007,N_18760);
or U19464 (N_19464,N_18910,N_18390);
or U19465 (N_19465,N_18600,N_18495);
xor U19466 (N_19466,N_18251,N_18375);
and U19467 (N_19467,N_18226,N_18349);
and U19468 (N_19468,N_18877,N_18140);
nor U19469 (N_19469,N_18794,N_18394);
and U19470 (N_19470,N_18637,N_18215);
nand U19471 (N_19471,N_18774,N_18282);
or U19472 (N_19472,N_18182,N_18376);
and U19473 (N_19473,N_18533,N_18054);
and U19474 (N_19474,N_18002,N_18484);
xor U19475 (N_19475,N_18575,N_18949);
nor U19476 (N_19476,N_18131,N_18076);
nor U19477 (N_19477,N_18319,N_18741);
and U19478 (N_19478,N_18892,N_18931);
or U19479 (N_19479,N_18902,N_18345);
xnor U19480 (N_19480,N_18441,N_18821);
xnor U19481 (N_19481,N_18003,N_18257);
and U19482 (N_19482,N_18342,N_18624);
or U19483 (N_19483,N_18616,N_18768);
or U19484 (N_19484,N_18606,N_18924);
xnor U19485 (N_19485,N_18075,N_18277);
xor U19486 (N_19486,N_18196,N_18842);
xnor U19487 (N_19487,N_18015,N_18073);
nor U19488 (N_19488,N_18867,N_18793);
and U19489 (N_19489,N_18720,N_18851);
nand U19490 (N_19490,N_18126,N_18737);
or U19491 (N_19491,N_18160,N_18873);
or U19492 (N_19492,N_18462,N_18733);
nand U19493 (N_19493,N_18230,N_18395);
and U19494 (N_19494,N_18941,N_18671);
or U19495 (N_19495,N_18809,N_18798);
and U19496 (N_19496,N_18554,N_18023);
nand U19497 (N_19497,N_18967,N_18833);
or U19498 (N_19498,N_18469,N_18069);
xnor U19499 (N_19499,N_18068,N_18102);
nand U19500 (N_19500,N_18947,N_18055);
xnor U19501 (N_19501,N_18874,N_18373);
and U19502 (N_19502,N_18444,N_18342);
nor U19503 (N_19503,N_18344,N_18769);
xnor U19504 (N_19504,N_18288,N_18575);
or U19505 (N_19505,N_18365,N_18438);
and U19506 (N_19506,N_18929,N_18510);
xor U19507 (N_19507,N_18625,N_18100);
xnor U19508 (N_19508,N_18154,N_18226);
xnor U19509 (N_19509,N_18829,N_18364);
nand U19510 (N_19510,N_18010,N_18951);
nor U19511 (N_19511,N_18487,N_18181);
nand U19512 (N_19512,N_18698,N_18745);
xnor U19513 (N_19513,N_18406,N_18240);
nand U19514 (N_19514,N_18632,N_18509);
nor U19515 (N_19515,N_18783,N_18238);
nand U19516 (N_19516,N_18795,N_18741);
or U19517 (N_19517,N_18669,N_18340);
xnor U19518 (N_19518,N_18566,N_18068);
and U19519 (N_19519,N_18600,N_18653);
nor U19520 (N_19520,N_18488,N_18997);
and U19521 (N_19521,N_18746,N_18154);
nor U19522 (N_19522,N_18310,N_18817);
nor U19523 (N_19523,N_18443,N_18336);
and U19524 (N_19524,N_18472,N_18580);
nand U19525 (N_19525,N_18645,N_18244);
nand U19526 (N_19526,N_18811,N_18651);
or U19527 (N_19527,N_18243,N_18559);
nand U19528 (N_19528,N_18106,N_18597);
and U19529 (N_19529,N_18144,N_18587);
or U19530 (N_19530,N_18146,N_18583);
nand U19531 (N_19531,N_18151,N_18795);
and U19532 (N_19532,N_18954,N_18027);
and U19533 (N_19533,N_18688,N_18610);
or U19534 (N_19534,N_18928,N_18786);
xor U19535 (N_19535,N_18553,N_18973);
or U19536 (N_19536,N_18614,N_18590);
or U19537 (N_19537,N_18939,N_18203);
and U19538 (N_19538,N_18713,N_18596);
or U19539 (N_19539,N_18809,N_18258);
nor U19540 (N_19540,N_18185,N_18923);
nor U19541 (N_19541,N_18464,N_18959);
xnor U19542 (N_19542,N_18553,N_18548);
nand U19543 (N_19543,N_18317,N_18570);
nor U19544 (N_19544,N_18004,N_18713);
nand U19545 (N_19545,N_18384,N_18105);
or U19546 (N_19546,N_18487,N_18964);
and U19547 (N_19547,N_18200,N_18583);
nand U19548 (N_19548,N_18731,N_18277);
xnor U19549 (N_19549,N_18048,N_18879);
or U19550 (N_19550,N_18163,N_18743);
or U19551 (N_19551,N_18967,N_18943);
and U19552 (N_19552,N_18367,N_18779);
nor U19553 (N_19553,N_18515,N_18534);
or U19554 (N_19554,N_18526,N_18283);
xnor U19555 (N_19555,N_18300,N_18998);
or U19556 (N_19556,N_18793,N_18415);
xor U19557 (N_19557,N_18647,N_18679);
xnor U19558 (N_19558,N_18838,N_18568);
or U19559 (N_19559,N_18780,N_18366);
nor U19560 (N_19560,N_18124,N_18864);
nand U19561 (N_19561,N_18773,N_18162);
nor U19562 (N_19562,N_18636,N_18846);
nand U19563 (N_19563,N_18839,N_18185);
and U19564 (N_19564,N_18880,N_18247);
nand U19565 (N_19565,N_18321,N_18101);
xor U19566 (N_19566,N_18736,N_18424);
xor U19567 (N_19567,N_18974,N_18410);
xnor U19568 (N_19568,N_18023,N_18015);
nor U19569 (N_19569,N_18164,N_18952);
xor U19570 (N_19570,N_18823,N_18171);
nand U19571 (N_19571,N_18258,N_18194);
nand U19572 (N_19572,N_18096,N_18038);
nand U19573 (N_19573,N_18125,N_18102);
and U19574 (N_19574,N_18823,N_18440);
xnor U19575 (N_19575,N_18128,N_18005);
nand U19576 (N_19576,N_18415,N_18101);
xnor U19577 (N_19577,N_18996,N_18237);
nand U19578 (N_19578,N_18504,N_18480);
nor U19579 (N_19579,N_18654,N_18625);
or U19580 (N_19580,N_18833,N_18302);
xor U19581 (N_19581,N_18904,N_18057);
or U19582 (N_19582,N_18107,N_18850);
or U19583 (N_19583,N_18423,N_18458);
and U19584 (N_19584,N_18307,N_18488);
nand U19585 (N_19585,N_18167,N_18966);
or U19586 (N_19586,N_18296,N_18034);
xnor U19587 (N_19587,N_18802,N_18023);
nand U19588 (N_19588,N_18051,N_18331);
xnor U19589 (N_19589,N_18081,N_18004);
nand U19590 (N_19590,N_18657,N_18573);
or U19591 (N_19591,N_18623,N_18497);
and U19592 (N_19592,N_18443,N_18624);
nand U19593 (N_19593,N_18281,N_18215);
nand U19594 (N_19594,N_18196,N_18844);
xnor U19595 (N_19595,N_18167,N_18541);
and U19596 (N_19596,N_18690,N_18239);
or U19597 (N_19597,N_18027,N_18961);
or U19598 (N_19598,N_18525,N_18338);
nor U19599 (N_19599,N_18814,N_18138);
nand U19600 (N_19600,N_18029,N_18026);
nor U19601 (N_19601,N_18006,N_18497);
nor U19602 (N_19602,N_18189,N_18238);
or U19603 (N_19603,N_18816,N_18170);
nand U19604 (N_19604,N_18995,N_18075);
xor U19605 (N_19605,N_18012,N_18185);
and U19606 (N_19606,N_18911,N_18030);
and U19607 (N_19607,N_18860,N_18913);
and U19608 (N_19608,N_18492,N_18241);
nand U19609 (N_19609,N_18409,N_18606);
nand U19610 (N_19610,N_18072,N_18309);
nor U19611 (N_19611,N_18005,N_18084);
nor U19612 (N_19612,N_18078,N_18787);
or U19613 (N_19613,N_18774,N_18519);
or U19614 (N_19614,N_18666,N_18972);
xor U19615 (N_19615,N_18629,N_18193);
and U19616 (N_19616,N_18208,N_18128);
xor U19617 (N_19617,N_18477,N_18504);
xor U19618 (N_19618,N_18491,N_18406);
nor U19619 (N_19619,N_18606,N_18586);
xnor U19620 (N_19620,N_18947,N_18213);
and U19621 (N_19621,N_18421,N_18532);
and U19622 (N_19622,N_18992,N_18128);
or U19623 (N_19623,N_18014,N_18456);
and U19624 (N_19624,N_18616,N_18593);
xnor U19625 (N_19625,N_18671,N_18297);
and U19626 (N_19626,N_18891,N_18744);
or U19627 (N_19627,N_18640,N_18036);
nor U19628 (N_19628,N_18535,N_18181);
and U19629 (N_19629,N_18527,N_18616);
xnor U19630 (N_19630,N_18120,N_18268);
xor U19631 (N_19631,N_18442,N_18971);
xor U19632 (N_19632,N_18134,N_18619);
and U19633 (N_19633,N_18250,N_18245);
nor U19634 (N_19634,N_18713,N_18070);
and U19635 (N_19635,N_18329,N_18726);
xnor U19636 (N_19636,N_18144,N_18385);
or U19637 (N_19637,N_18702,N_18552);
and U19638 (N_19638,N_18421,N_18816);
and U19639 (N_19639,N_18472,N_18606);
xnor U19640 (N_19640,N_18956,N_18650);
nor U19641 (N_19641,N_18221,N_18115);
xor U19642 (N_19642,N_18608,N_18718);
xnor U19643 (N_19643,N_18099,N_18414);
or U19644 (N_19644,N_18336,N_18471);
or U19645 (N_19645,N_18121,N_18494);
or U19646 (N_19646,N_18075,N_18953);
nor U19647 (N_19647,N_18755,N_18441);
nand U19648 (N_19648,N_18698,N_18763);
nand U19649 (N_19649,N_18558,N_18951);
xnor U19650 (N_19650,N_18824,N_18777);
xnor U19651 (N_19651,N_18062,N_18417);
and U19652 (N_19652,N_18630,N_18178);
xnor U19653 (N_19653,N_18690,N_18247);
and U19654 (N_19654,N_18866,N_18570);
nor U19655 (N_19655,N_18126,N_18284);
nand U19656 (N_19656,N_18005,N_18828);
or U19657 (N_19657,N_18744,N_18598);
nor U19658 (N_19658,N_18777,N_18837);
nor U19659 (N_19659,N_18684,N_18670);
nor U19660 (N_19660,N_18279,N_18327);
or U19661 (N_19661,N_18698,N_18204);
nand U19662 (N_19662,N_18948,N_18889);
xnor U19663 (N_19663,N_18720,N_18677);
and U19664 (N_19664,N_18120,N_18580);
nor U19665 (N_19665,N_18346,N_18727);
or U19666 (N_19666,N_18273,N_18564);
or U19667 (N_19667,N_18825,N_18908);
or U19668 (N_19668,N_18709,N_18496);
or U19669 (N_19669,N_18664,N_18182);
nor U19670 (N_19670,N_18536,N_18772);
xor U19671 (N_19671,N_18912,N_18379);
xnor U19672 (N_19672,N_18071,N_18079);
nand U19673 (N_19673,N_18950,N_18658);
nor U19674 (N_19674,N_18902,N_18648);
nor U19675 (N_19675,N_18054,N_18363);
xor U19676 (N_19676,N_18065,N_18774);
and U19677 (N_19677,N_18701,N_18143);
xor U19678 (N_19678,N_18213,N_18380);
or U19679 (N_19679,N_18537,N_18252);
nor U19680 (N_19680,N_18921,N_18301);
or U19681 (N_19681,N_18605,N_18388);
nand U19682 (N_19682,N_18813,N_18595);
and U19683 (N_19683,N_18066,N_18028);
nand U19684 (N_19684,N_18325,N_18639);
nand U19685 (N_19685,N_18341,N_18496);
nor U19686 (N_19686,N_18865,N_18544);
xor U19687 (N_19687,N_18024,N_18419);
nand U19688 (N_19688,N_18851,N_18525);
and U19689 (N_19689,N_18805,N_18161);
or U19690 (N_19690,N_18509,N_18520);
xor U19691 (N_19691,N_18664,N_18393);
and U19692 (N_19692,N_18940,N_18837);
xnor U19693 (N_19693,N_18448,N_18966);
xor U19694 (N_19694,N_18234,N_18408);
nand U19695 (N_19695,N_18836,N_18716);
or U19696 (N_19696,N_18549,N_18384);
nor U19697 (N_19697,N_18402,N_18599);
nand U19698 (N_19698,N_18191,N_18812);
nor U19699 (N_19699,N_18171,N_18041);
xor U19700 (N_19700,N_18872,N_18318);
xnor U19701 (N_19701,N_18253,N_18617);
nor U19702 (N_19702,N_18703,N_18848);
nor U19703 (N_19703,N_18650,N_18619);
nor U19704 (N_19704,N_18041,N_18697);
nand U19705 (N_19705,N_18684,N_18561);
nor U19706 (N_19706,N_18075,N_18630);
and U19707 (N_19707,N_18195,N_18416);
nand U19708 (N_19708,N_18770,N_18938);
nor U19709 (N_19709,N_18513,N_18948);
nand U19710 (N_19710,N_18319,N_18085);
or U19711 (N_19711,N_18355,N_18374);
and U19712 (N_19712,N_18454,N_18626);
and U19713 (N_19713,N_18829,N_18859);
nand U19714 (N_19714,N_18067,N_18746);
or U19715 (N_19715,N_18413,N_18542);
xnor U19716 (N_19716,N_18082,N_18484);
nor U19717 (N_19717,N_18492,N_18157);
nand U19718 (N_19718,N_18781,N_18587);
or U19719 (N_19719,N_18398,N_18680);
nor U19720 (N_19720,N_18188,N_18318);
nor U19721 (N_19721,N_18133,N_18591);
and U19722 (N_19722,N_18013,N_18365);
xor U19723 (N_19723,N_18824,N_18582);
xnor U19724 (N_19724,N_18731,N_18823);
and U19725 (N_19725,N_18992,N_18216);
nor U19726 (N_19726,N_18166,N_18914);
nor U19727 (N_19727,N_18143,N_18672);
nand U19728 (N_19728,N_18873,N_18854);
nor U19729 (N_19729,N_18825,N_18736);
nand U19730 (N_19730,N_18669,N_18987);
nor U19731 (N_19731,N_18141,N_18710);
nand U19732 (N_19732,N_18292,N_18725);
nand U19733 (N_19733,N_18924,N_18055);
nor U19734 (N_19734,N_18457,N_18283);
nor U19735 (N_19735,N_18743,N_18802);
or U19736 (N_19736,N_18394,N_18503);
nor U19737 (N_19737,N_18284,N_18525);
nor U19738 (N_19738,N_18298,N_18836);
nand U19739 (N_19739,N_18833,N_18630);
xnor U19740 (N_19740,N_18227,N_18081);
or U19741 (N_19741,N_18091,N_18501);
and U19742 (N_19742,N_18924,N_18618);
nor U19743 (N_19743,N_18183,N_18510);
and U19744 (N_19744,N_18738,N_18166);
and U19745 (N_19745,N_18237,N_18852);
nor U19746 (N_19746,N_18323,N_18607);
xor U19747 (N_19747,N_18697,N_18393);
and U19748 (N_19748,N_18811,N_18124);
nand U19749 (N_19749,N_18014,N_18413);
nand U19750 (N_19750,N_18325,N_18686);
nor U19751 (N_19751,N_18164,N_18046);
or U19752 (N_19752,N_18915,N_18038);
xnor U19753 (N_19753,N_18171,N_18050);
and U19754 (N_19754,N_18274,N_18812);
and U19755 (N_19755,N_18773,N_18537);
nand U19756 (N_19756,N_18517,N_18587);
nor U19757 (N_19757,N_18766,N_18321);
or U19758 (N_19758,N_18571,N_18088);
nand U19759 (N_19759,N_18080,N_18454);
xor U19760 (N_19760,N_18202,N_18309);
nor U19761 (N_19761,N_18688,N_18172);
nand U19762 (N_19762,N_18438,N_18548);
xnor U19763 (N_19763,N_18592,N_18788);
or U19764 (N_19764,N_18785,N_18023);
xor U19765 (N_19765,N_18547,N_18196);
or U19766 (N_19766,N_18421,N_18153);
or U19767 (N_19767,N_18600,N_18060);
and U19768 (N_19768,N_18957,N_18461);
nand U19769 (N_19769,N_18131,N_18620);
xnor U19770 (N_19770,N_18483,N_18559);
or U19771 (N_19771,N_18536,N_18584);
nand U19772 (N_19772,N_18975,N_18003);
xor U19773 (N_19773,N_18259,N_18566);
or U19774 (N_19774,N_18653,N_18554);
nor U19775 (N_19775,N_18094,N_18947);
nand U19776 (N_19776,N_18983,N_18830);
or U19777 (N_19777,N_18067,N_18472);
nor U19778 (N_19778,N_18171,N_18877);
nor U19779 (N_19779,N_18173,N_18848);
xor U19780 (N_19780,N_18808,N_18465);
or U19781 (N_19781,N_18458,N_18414);
or U19782 (N_19782,N_18313,N_18252);
and U19783 (N_19783,N_18934,N_18311);
xor U19784 (N_19784,N_18413,N_18868);
xor U19785 (N_19785,N_18222,N_18758);
nand U19786 (N_19786,N_18126,N_18825);
nand U19787 (N_19787,N_18799,N_18279);
xnor U19788 (N_19788,N_18922,N_18593);
nor U19789 (N_19789,N_18010,N_18436);
and U19790 (N_19790,N_18207,N_18929);
or U19791 (N_19791,N_18582,N_18056);
and U19792 (N_19792,N_18871,N_18931);
or U19793 (N_19793,N_18673,N_18374);
xor U19794 (N_19794,N_18877,N_18257);
nor U19795 (N_19795,N_18821,N_18925);
nor U19796 (N_19796,N_18659,N_18527);
nand U19797 (N_19797,N_18050,N_18145);
or U19798 (N_19798,N_18141,N_18143);
and U19799 (N_19799,N_18420,N_18510);
and U19800 (N_19800,N_18286,N_18422);
or U19801 (N_19801,N_18125,N_18849);
xnor U19802 (N_19802,N_18714,N_18973);
nor U19803 (N_19803,N_18207,N_18494);
xor U19804 (N_19804,N_18372,N_18569);
xnor U19805 (N_19805,N_18072,N_18746);
or U19806 (N_19806,N_18110,N_18656);
nor U19807 (N_19807,N_18056,N_18458);
and U19808 (N_19808,N_18188,N_18042);
or U19809 (N_19809,N_18185,N_18471);
or U19810 (N_19810,N_18569,N_18471);
or U19811 (N_19811,N_18210,N_18693);
or U19812 (N_19812,N_18387,N_18471);
nand U19813 (N_19813,N_18237,N_18410);
and U19814 (N_19814,N_18121,N_18286);
nor U19815 (N_19815,N_18113,N_18551);
or U19816 (N_19816,N_18480,N_18850);
xnor U19817 (N_19817,N_18349,N_18350);
xor U19818 (N_19818,N_18126,N_18073);
xnor U19819 (N_19819,N_18436,N_18267);
nand U19820 (N_19820,N_18120,N_18768);
and U19821 (N_19821,N_18919,N_18330);
or U19822 (N_19822,N_18989,N_18716);
nor U19823 (N_19823,N_18599,N_18695);
nor U19824 (N_19824,N_18360,N_18251);
xnor U19825 (N_19825,N_18129,N_18958);
nor U19826 (N_19826,N_18344,N_18947);
nor U19827 (N_19827,N_18947,N_18916);
or U19828 (N_19828,N_18899,N_18889);
xnor U19829 (N_19829,N_18091,N_18421);
xnor U19830 (N_19830,N_18620,N_18647);
and U19831 (N_19831,N_18903,N_18435);
xnor U19832 (N_19832,N_18602,N_18778);
or U19833 (N_19833,N_18224,N_18365);
nand U19834 (N_19834,N_18928,N_18061);
xor U19835 (N_19835,N_18853,N_18839);
nor U19836 (N_19836,N_18058,N_18955);
nor U19837 (N_19837,N_18432,N_18657);
and U19838 (N_19838,N_18766,N_18435);
xnor U19839 (N_19839,N_18763,N_18078);
or U19840 (N_19840,N_18621,N_18994);
xor U19841 (N_19841,N_18784,N_18923);
nor U19842 (N_19842,N_18093,N_18763);
or U19843 (N_19843,N_18097,N_18753);
xor U19844 (N_19844,N_18986,N_18864);
nor U19845 (N_19845,N_18158,N_18472);
xor U19846 (N_19846,N_18117,N_18773);
and U19847 (N_19847,N_18075,N_18942);
and U19848 (N_19848,N_18712,N_18228);
and U19849 (N_19849,N_18807,N_18094);
nor U19850 (N_19850,N_18930,N_18614);
xnor U19851 (N_19851,N_18355,N_18324);
and U19852 (N_19852,N_18280,N_18041);
nand U19853 (N_19853,N_18083,N_18826);
or U19854 (N_19854,N_18499,N_18451);
or U19855 (N_19855,N_18532,N_18971);
nor U19856 (N_19856,N_18880,N_18851);
or U19857 (N_19857,N_18723,N_18201);
nand U19858 (N_19858,N_18465,N_18240);
and U19859 (N_19859,N_18257,N_18349);
or U19860 (N_19860,N_18219,N_18762);
nand U19861 (N_19861,N_18964,N_18676);
xnor U19862 (N_19862,N_18918,N_18737);
nor U19863 (N_19863,N_18064,N_18090);
or U19864 (N_19864,N_18495,N_18265);
and U19865 (N_19865,N_18429,N_18972);
nand U19866 (N_19866,N_18781,N_18441);
and U19867 (N_19867,N_18088,N_18305);
nand U19868 (N_19868,N_18140,N_18473);
nor U19869 (N_19869,N_18321,N_18182);
or U19870 (N_19870,N_18373,N_18385);
xnor U19871 (N_19871,N_18358,N_18296);
or U19872 (N_19872,N_18416,N_18353);
nand U19873 (N_19873,N_18892,N_18190);
and U19874 (N_19874,N_18305,N_18891);
or U19875 (N_19875,N_18444,N_18454);
and U19876 (N_19876,N_18075,N_18669);
and U19877 (N_19877,N_18507,N_18389);
nand U19878 (N_19878,N_18883,N_18119);
nand U19879 (N_19879,N_18469,N_18160);
or U19880 (N_19880,N_18042,N_18835);
and U19881 (N_19881,N_18148,N_18360);
and U19882 (N_19882,N_18803,N_18491);
xor U19883 (N_19883,N_18784,N_18269);
nor U19884 (N_19884,N_18569,N_18371);
or U19885 (N_19885,N_18229,N_18909);
xnor U19886 (N_19886,N_18678,N_18358);
nand U19887 (N_19887,N_18852,N_18933);
nand U19888 (N_19888,N_18191,N_18612);
xor U19889 (N_19889,N_18728,N_18100);
or U19890 (N_19890,N_18294,N_18707);
xor U19891 (N_19891,N_18484,N_18031);
nand U19892 (N_19892,N_18823,N_18902);
and U19893 (N_19893,N_18531,N_18027);
and U19894 (N_19894,N_18256,N_18863);
and U19895 (N_19895,N_18353,N_18412);
xor U19896 (N_19896,N_18849,N_18707);
and U19897 (N_19897,N_18430,N_18858);
xnor U19898 (N_19898,N_18361,N_18124);
or U19899 (N_19899,N_18626,N_18672);
or U19900 (N_19900,N_18601,N_18548);
and U19901 (N_19901,N_18107,N_18853);
xnor U19902 (N_19902,N_18547,N_18399);
xor U19903 (N_19903,N_18945,N_18505);
or U19904 (N_19904,N_18131,N_18599);
nor U19905 (N_19905,N_18580,N_18233);
and U19906 (N_19906,N_18960,N_18139);
xnor U19907 (N_19907,N_18714,N_18859);
xor U19908 (N_19908,N_18772,N_18023);
or U19909 (N_19909,N_18143,N_18113);
nand U19910 (N_19910,N_18095,N_18605);
xor U19911 (N_19911,N_18625,N_18770);
or U19912 (N_19912,N_18599,N_18198);
and U19913 (N_19913,N_18386,N_18845);
or U19914 (N_19914,N_18196,N_18267);
xor U19915 (N_19915,N_18580,N_18461);
xor U19916 (N_19916,N_18264,N_18869);
or U19917 (N_19917,N_18725,N_18614);
xnor U19918 (N_19918,N_18615,N_18239);
nor U19919 (N_19919,N_18489,N_18484);
or U19920 (N_19920,N_18482,N_18963);
or U19921 (N_19921,N_18171,N_18651);
xnor U19922 (N_19922,N_18896,N_18060);
nor U19923 (N_19923,N_18249,N_18749);
xnor U19924 (N_19924,N_18697,N_18811);
xor U19925 (N_19925,N_18960,N_18336);
xnor U19926 (N_19926,N_18666,N_18329);
xor U19927 (N_19927,N_18863,N_18411);
and U19928 (N_19928,N_18238,N_18316);
or U19929 (N_19929,N_18768,N_18585);
nand U19930 (N_19930,N_18309,N_18672);
nor U19931 (N_19931,N_18443,N_18949);
and U19932 (N_19932,N_18129,N_18117);
nand U19933 (N_19933,N_18980,N_18366);
and U19934 (N_19934,N_18513,N_18913);
or U19935 (N_19935,N_18854,N_18000);
nand U19936 (N_19936,N_18031,N_18353);
and U19937 (N_19937,N_18814,N_18275);
nor U19938 (N_19938,N_18481,N_18308);
or U19939 (N_19939,N_18808,N_18212);
and U19940 (N_19940,N_18851,N_18105);
xnor U19941 (N_19941,N_18719,N_18589);
nand U19942 (N_19942,N_18240,N_18994);
nand U19943 (N_19943,N_18951,N_18804);
and U19944 (N_19944,N_18368,N_18911);
and U19945 (N_19945,N_18200,N_18693);
or U19946 (N_19946,N_18170,N_18525);
xnor U19947 (N_19947,N_18389,N_18707);
nand U19948 (N_19948,N_18496,N_18406);
nand U19949 (N_19949,N_18834,N_18276);
nand U19950 (N_19950,N_18526,N_18531);
or U19951 (N_19951,N_18543,N_18824);
or U19952 (N_19952,N_18655,N_18961);
or U19953 (N_19953,N_18000,N_18479);
xnor U19954 (N_19954,N_18258,N_18206);
nand U19955 (N_19955,N_18884,N_18758);
and U19956 (N_19956,N_18816,N_18297);
xnor U19957 (N_19957,N_18367,N_18995);
nand U19958 (N_19958,N_18008,N_18396);
and U19959 (N_19959,N_18809,N_18379);
or U19960 (N_19960,N_18969,N_18758);
nor U19961 (N_19961,N_18586,N_18498);
nor U19962 (N_19962,N_18563,N_18296);
nand U19963 (N_19963,N_18253,N_18872);
and U19964 (N_19964,N_18294,N_18827);
nand U19965 (N_19965,N_18942,N_18055);
or U19966 (N_19966,N_18777,N_18495);
and U19967 (N_19967,N_18577,N_18734);
xnor U19968 (N_19968,N_18826,N_18631);
nor U19969 (N_19969,N_18582,N_18116);
or U19970 (N_19970,N_18200,N_18051);
xnor U19971 (N_19971,N_18996,N_18416);
or U19972 (N_19972,N_18348,N_18787);
and U19973 (N_19973,N_18166,N_18710);
nand U19974 (N_19974,N_18709,N_18358);
nor U19975 (N_19975,N_18122,N_18879);
nor U19976 (N_19976,N_18431,N_18916);
nand U19977 (N_19977,N_18355,N_18705);
xnor U19978 (N_19978,N_18497,N_18484);
nand U19979 (N_19979,N_18138,N_18029);
nand U19980 (N_19980,N_18789,N_18162);
nor U19981 (N_19981,N_18997,N_18417);
and U19982 (N_19982,N_18182,N_18738);
and U19983 (N_19983,N_18436,N_18564);
xor U19984 (N_19984,N_18544,N_18251);
xor U19985 (N_19985,N_18161,N_18607);
and U19986 (N_19986,N_18371,N_18797);
nand U19987 (N_19987,N_18307,N_18666);
and U19988 (N_19988,N_18243,N_18187);
or U19989 (N_19989,N_18057,N_18201);
nand U19990 (N_19990,N_18902,N_18983);
and U19991 (N_19991,N_18654,N_18161);
or U19992 (N_19992,N_18604,N_18748);
xor U19993 (N_19993,N_18550,N_18582);
and U19994 (N_19994,N_18418,N_18968);
and U19995 (N_19995,N_18317,N_18614);
xnor U19996 (N_19996,N_18946,N_18141);
nor U19997 (N_19997,N_18772,N_18671);
nand U19998 (N_19998,N_18219,N_18551);
nor U19999 (N_19999,N_18897,N_18673);
and U20000 (N_20000,N_19712,N_19826);
xnor U20001 (N_20001,N_19530,N_19024);
nand U20002 (N_20002,N_19103,N_19964);
or U20003 (N_20003,N_19012,N_19715);
or U20004 (N_20004,N_19172,N_19076);
or U20005 (N_20005,N_19142,N_19561);
nand U20006 (N_20006,N_19830,N_19084);
nand U20007 (N_20007,N_19909,N_19592);
xnor U20008 (N_20008,N_19202,N_19043);
nand U20009 (N_20009,N_19318,N_19697);
and U20010 (N_20010,N_19289,N_19546);
xor U20011 (N_20011,N_19124,N_19010);
nand U20012 (N_20012,N_19558,N_19719);
or U20013 (N_20013,N_19856,N_19709);
and U20014 (N_20014,N_19096,N_19746);
nor U20015 (N_20015,N_19358,N_19483);
and U20016 (N_20016,N_19920,N_19735);
nor U20017 (N_20017,N_19764,N_19571);
or U20018 (N_20018,N_19122,N_19778);
xor U20019 (N_20019,N_19685,N_19209);
xor U20020 (N_20020,N_19934,N_19452);
and U20021 (N_20021,N_19216,N_19665);
nand U20022 (N_20022,N_19528,N_19635);
or U20023 (N_20023,N_19682,N_19540);
xnor U20024 (N_20024,N_19754,N_19441);
nor U20025 (N_20025,N_19023,N_19677);
nand U20026 (N_20026,N_19393,N_19969);
xnor U20027 (N_20027,N_19505,N_19845);
and U20028 (N_20028,N_19718,N_19440);
nand U20029 (N_20029,N_19083,N_19991);
and U20030 (N_20030,N_19622,N_19354);
or U20031 (N_20031,N_19572,N_19872);
nand U20032 (N_20032,N_19721,N_19543);
or U20033 (N_20033,N_19437,N_19234);
nand U20034 (N_20034,N_19492,N_19716);
nor U20035 (N_20035,N_19935,N_19495);
nand U20036 (N_20036,N_19187,N_19097);
or U20037 (N_20037,N_19504,N_19694);
and U20038 (N_20038,N_19950,N_19650);
nor U20039 (N_20039,N_19162,N_19555);
or U20040 (N_20040,N_19183,N_19002);
xnor U20041 (N_20041,N_19156,N_19545);
or U20042 (N_20042,N_19959,N_19831);
or U20043 (N_20043,N_19021,N_19873);
nand U20044 (N_20044,N_19356,N_19229);
and U20045 (N_20045,N_19055,N_19379);
nor U20046 (N_20046,N_19725,N_19405);
and U20047 (N_20047,N_19869,N_19494);
or U20048 (N_20048,N_19863,N_19606);
nor U20049 (N_20049,N_19929,N_19008);
nor U20050 (N_20050,N_19490,N_19315);
xor U20051 (N_20051,N_19028,N_19827);
nor U20052 (N_20052,N_19154,N_19784);
nor U20053 (N_20053,N_19663,N_19302);
nand U20054 (N_20054,N_19816,N_19375);
and U20055 (N_20055,N_19502,N_19695);
nor U20056 (N_20056,N_19787,N_19348);
nor U20057 (N_20057,N_19460,N_19346);
and U20058 (N_20058,N_19705,N_19475);
or U20059 (N_20059,N_19428,N_19951);
nand U20060 (N_20060,N_19193,N_19459);
nor U20061 (N_20061,N_19423,N_19506);
and U20062 (N_20062,N_19780,N_19275);
xor U20063 (N_20063,N_19840,N_19651);
nor U20064 (N_20064,N_19400,N_19168);
nand U20065 (N_20065,N_19252,N_19353);
nor U20066 (N_20066,N_19113,N_19591);
nand U20067 (N_20067,N_19443,N_19101);
and U20068 (N_20068,N_19902,N_19066);
nor U20069 (N_20069,N_19489,N_19013);
and U20070 (N_20070,N_19563,N_19645);
xnor U20071 (N_20071,N_19064,N_19904);
or U20072 (N_20072,N_19903,N_19881);
and U20073 (N_20073,N_19107,N_19480);
xnor U20074 (N_20074,N_19847,N_19966);
nand U20075 (N_20075,N_19493,N_19818);
and U20076 (N_20076,N_19485,N_19582);
xnor U20077 (N_20077,N_19794,N_19173);
nand U20078 (N_20078,N_19415,N_19871);
xnor U20079 (N_20079,N_19453,N_19919);
nand U20080 (N_20080,N_19740,N_19262);
or U20081 (N_20081,N_19713,N_19906);
nand U20082 (N_20082,N_19549,N_19327);
or U20083 (N_20083,N_19553,N_19698);
or U20084 (N_20084,N_19300,N_19466);
nor U20085 (N_20085,N_19307,N_19538);
xnor U20086 (N_20086,N_19081,N_19511);
or U20087 (N_20087,N_19153,N_19998);
nor U20088 (N_20088,N_19377,N_19630);
xor U20089 (N_20089,N_19954,N_19636);
nand U20090 (N_20090,N_19838,N_19844);
xor U20091 (N_20091,N_19340,N_19956);
or U20092 (N_20092,N_19851,N_19771);
or U20093 (N_20093,N_19522,N_19350);
xnor U20094 (N_20094,N_19210,N_19349);
or U20095 (N_20095,N_19814,N_19503);
and U20096 (N_20096,N_19926,N_19805);
nor U20097 (N_20097,N_19184,N_19708);
nor U20098 (N_20098,N_19444,N_19821);
and U20099 (N_20099,N_19343,N_19226);
nor U20100 (N_20100,N_19603,N_19017);
xnor U20101 (N_20101,N_19638,N_19120);
nand U20102 (N_20102,N_19996,N_19696);
or U20103 (N_20103,N_19259,N_19491);
nor U20104 (N_20104,N_19781,N_19641);
nand U20105 (N_20105,N_19885,N_19086);
nor U20106 (N_20106,N_19333,N_19870);
or U20107 (N_20107,N_19027,N_19102);
nand U20108 (N_20108,N_19446,N_19512);
xor U20109 (N_20109,N_19073,N_19114);
nor U20110 (N_20110,N_19866,N_19738);
nor U20111 (N_20111,N_19999,N_19632);
nand U20112 (N_20112,N_19811,N_19848);
xnor U20113 (N_20113,N_19352,N_19949);
or U20114 (N_20114,N_19276,N_19736);
xor U20115 (N_20115,N_19237,N_19051);
or U20116 (N_20116,N_19913,N_19883);
xor U20117 (N_20117,N_19617,N_19053);
or U20118 (N_20118,N_19213,N_19843);
or U20119 (N_20119,N_19823,N_19240);
xnor U20120 (N_20120,N_19282,N_19634);
or U20121 (N_20121,N_19703,N_19834);
and U20122 (N_20122,N_19365,N_19970);
xor U20123 (N_20123,N_19457,N_19339);
xor U20124 (N_20124,N_19884,N_19230);
nor U20125 (N_20125,N_19517,N_19527);
nand U20126 (N_20126,N_19861,N_19803);
xor U20127 (N_20127,N_19813,N_19171);
and U20128 (N_20128,N_19573,N_19701);
and U20129 (N_20129,N_19133,N_19798);
nand U20130 (N_20130,N_19401,N_19940);
nand U20131 (N_20131,N_19329,N_19320);
xor U20132 (N_20132,N_19693,N_19243);
nor U20133 (N_20133,N_19141,N_19625);
nor U20134 (N_20134,N_19724,N_19316);
xnor U20135 (N_20135,N_19052,N_19192);
xnor U20136 (N_20136,N_19657,N_19468);
and U20137 (N_20137,N_19147,N_19125);
nor U20138 (N_20138,N_19983,N_19150);
or U20139 (N_20139,N_19034,N_19201);
nor U20140 (N_20140,N_19775,N_19067);
nor U20141 (N_20141,N_19305,N_19488);
and U20142 (N_20142,N_19621,N_19857);
xor U20143 (N_20143,N_19743,N_19501);
and U20144 (N_20144,N_19667,N_19879);
nor U20145 (N_20145,N_19948,N_19409);
or U20146 (N_20146,N_19600,N_19733);
xor U20147 (N_20147,N_19245,N_19808);
and U20148 (N_20148,N_19536,N_19706);
nor U20149 (N_20149,N_19464,N_19266);
nor U20150 (N_20150,N_19304,N_19456);
nor U20151 (N_20151,N_19687,N_19539);
nor U20152 (N_20152,N_19077,N_19526);
xor U20153 (N_20153,N_19601,N_19961);
or U20154 (N_20154,N_19058,N_19412);
xor U20155 (N_20155,N_19432,N_19788);
or U20156 (N_20156,N_19143,N_19106);
nor U20157 (N_20157,N_19394,N_19233);
xor U20158 (N_20158,N_19189,N_19411);
nor U20159 (N_20159,N_19299,N_19859);
xor U20160 (N_20160,N_19280,N_19268);
or U20161 (N_20161,N_19029,N_19417);
nand U20162 (N_20162,N_19551,N_19059);
nand U20163 (N_20163,N_19542,N_19197);
nand U20164 (N_20164,N_19045,N_19860);
and U20165 (N_20165,N_19242,N_19118);
nor U20166 (N_20166,N_19850,N_19577);
nor U20167 (N_20167,N_19232,N_19759);
and U20168 (N_20168,N_19837,N_19673);
xnor U20169 (N_20169,N_19054,N_19249);
nand U20170 (N_20170,N_19250,N_19430);
or U20171 (N_20171,N_19867,N_19018);
or U20172 (N_20172,N_19774,N_19825);
nor U20173 (N_20173,N_19656,N_19975);
nor U20174 (N_20174,N_19596,N_19618);
and U20175 (N_20175,N_19947,N_19758);
and U20176 (N_20176,N_19944,N_19169);
xor U20177 (N_20177,N_19541,N_19214);
nand U20178 (N_20178,N_19098,N_19777);
or U20179 (N_20179,N_19878,N_19293);
and U20180 (N_20180,N_19039,N_19410);
xor U20181 (N_20181,N_19152,N_19971);
nor U20182 (N_20182,N_19036,N_19978);
or U20183 (N_20183,N_19310,N_19416);
nand U20184 (N_20184,N_19224,N_19135);
or U20185 (N_20185,N_19565,N_19195);
or U20186 (N_20186,N_19121,N_19104);
and U20187 (N_20187,N_19567,N_19720);
and U20188 (N_20188,N_19373,N_19633);
and U20189 (N_20189,N_19616,N_19734);
xnor U20190 (N_20190,N_19014,N_19710);
and U20191 (N_20191,N_19853,N_19898);
nand U20192 (N_20192,N_19085,N_19547);
and U20193 (N_20193,N_19387,N_19313);
and U20194 (N_20194,N_19980,N_19360);
or U20195 (N_20195,N_19020,N_19936);
nor U20196 (N_20196,N_19953,N_19938);
and U20197 (N_20197,N_19439,N_19392);
and U20198 (N_20198,N_19741,N_19995);
and U20199 (N_20199,N_19131,N_19089);
xor U20200 (N_20200,N_19297,N_19513);
or U20201 (N_20201,N_19672,N_19175);
and U20202 (N_20202,N_19942,N_19281);
nor U20203 (N_20203,N_19434,N_19612);
and U20204 (N_20204,N_19855,N_19960);
xnor U20205 (N_20205,N_19351,N_19585);
and U20206 (N_20206,N_19287,N_19979);
nor U20207 (N_20207,N_19324,N_19655);
nor U20208 (N_20208,N_19939,N_19198);
nand U20209 (N_20209,N_19070,N_19060);
nand U20210 (N_20210,N_19882,N_19862);
nand U20211 (N_20211,N_19004,N_19976);
or U20212 (N_20212,N_19963,N_19742);
nor U20213 (N_20213,N_19203,N_19448);
nand U20214 (N_20214,N_19186,N_19217);
nor U20215 (N_20215,N_19537,N_19498);
nand U20216 (N_20216,N_19946,N_19127);
nor U20217 (N_20217,N_19306,N_19160);
and U20218 (N_20218,N_19091,N_19602);
or U20219 (N_20219,N_19810,N_19296);
or U20220 (N_20220,N_19075,N_19586);
nor U20221 (N_20221,N_19727,N_19574);
xor U20222 (N_20222,N_19032,N_19544);
nor U20223 (N_20223,N_19531,N_19637);
or U20224 (N_20224,N_19836,N_19005);
nand U20225 (N_20225,N_19167,N_19659);
or U20226 (N_20226,N_19450,N_19654);
nor U20227 (N_20227,N_19311,N_19690);
or U20228 (N_20228,N_19225,N_19072);
xnor U20229 (N_20229,N_19916,N_19199);
nand U20230 (N_20230,N_19381,N_19748);
and U20231 (N_20231,N_19515,N_19472);
and U20232 (N_20232,N_19436,N_19370);
xnor U20233 (N_20233,N_19852,N_19057);
and U20234 (N_20234,N_19227,N_19395);
and U20235 (N_20235,N_19368,N_19478);
or U20236 (N_20236,N_19469,N_19792);
or U20237 (N_20237,N_19977,N_19588);
xnor U20238 (N_20238,N_19328,N_19760);
and U20239 (N_20239,N_19997,N_19509);
and U20240 (N_20240,N_19425,N_19649);
or U20241 (N_20241,N_19824,N_19896);
nand U20242 (N_20242,N_19389,N_19092);
nor U20243 (N_20243,N_19974,N_19802);
nor U20244 (N_20244,N_19560,N_19769);
xnor U20245 (N_20245,N_19514,N_19148);
xor U20246 (N_20246,N_19212,N_19119);
and U20247 (N_20247,N_19144,N_19668);
or U20248 (N_20248,N_19367,N_19112);
and U20249 (N_20249,N_19181,N_19065);
nand U20250 (N_20250,N_19623,N_19404);
xor U20251 (N_20251,N_19462,N_19643);
nor U20252 (N_20252,N_19943,N_19554);
or U20253 (N_20253,N_19264,N_19548);
nor U20254 (N_20254,N_19731,N_19180);
nor U20255 (N_20255,N_19990,N_19550);
xnor U20256 (N_20256,N_19841,N_19552);
and U20257 (N_20257,N_19858,N_19000);
nand U20258 (N_20258,N_19228,N_19557);
xnor U20259 (N_20259,N_19256,N_19666);
or U20260 (N_20260,N_19793,N_19194);
xor U20261 (N_20261,N_19846,N_19797);
nand U20262 (N_20262,N_19042,N_19263);
nor U20263 (N_20263,N_19681,N_19185);
nand U20264 (N_20264,N_19080,N_19800);
nand U20265 (N_20265,N_19717,N_19179);
nor U20266 (N_20266,N_19988,N_19994);
nor U20267 (N_20267,N_19556,N_19369);
and U20268 (N_20268,N_19007,N_19383);
xnor U20269 (N_20269,N_19487,N_19191);
nor U20270 (N_20270,N_19868,N_19090);
xnor U20271 (N_20271,N_19078,N_19644);
xor U20272 (N_20272,N_19484,N_19149);
or U20273 (N_20273,N_19519,N_19279);
and U20274 (N_20274,N_19614,N_19962);
xor U20275 (N_20275,N_19615,N_19330);
nor U20276 (N_20276,N_19011,N_19905);
nor U20277 (N_20277,N_19033,N_19166);
and U20278 (N_20278,N_19178,N_19362);
nor U20279 (N_20279,N_19188,N_19100);
nor U20280 (N_20280,N_19277,N_19447);
nand U20281 (N_20281,N_19581,N_19674);
or U20282 (N_20282,N_19048,N_19757);
or U20283 (N_20283,N_19426,N_19445);
and U20284 (N_20284,N_19912,N_19965);
nor U20285 (N_20285,N_19177,N_19074);
or U20286 (N_20286,N_19454,N_19063);
or U20287 (N_20287,N_19314,N_19982);
nor U20288 (N_20288,N_19670,N_19497);
and U20289 (N_20289,N_19308,N_19116);
nor U20290 (N_20290,N_19768,N_19918);
nand U20291 (N_20291,N_19496,N_19753);
xor U20292 (N_20292,N_19533,N_19608);
nand U20293 (N_20293,N_19130,N_19886);
nor U20294 (N_20294,N_19595,N_19791);
or U20295 (N_20295,N_19006,N_19105);
and U20296 (N_20296,N_19876,N_19239);
xor U20297 (N_20297,N_19799,N_19463);
nand U20298 (N_20298,N_19499,N_19094);
xnor U20299 (N_20299,N_19875,N_19967);
and U20300 (N_20300,N_19986,N_19564);
and U20301 (N_20301,N_19255,N_19022);
nand U20302 (N_20302,N_19786,N_19474);
nand U20303 (N_20303,N_19317,N_19236);
nor U20304 (N_20304,N_19334,N_19762);
xor U20305 (N_20305,N_19516,N_19521);
or U20306 (N_20306,N_19569,N_19689);
and U20307 (N_20307,N_19985,N_19126);
and U20308 (N_20308,N_19215,N_19925);
nor U20309 (N_20309,N_19767,N_19729);
and U20310 (N_20310,N_19730,N_19190);
and U20311 (N_20311,N_19206,N_19322);
nor U20312 (N_20312,N_19639,N_19291);
or U20313 (N_20313,N_19482,N_19136);
xor U20314 (N_20314,N_19923,N_19749);
or U20315 (N_20315,N_19038,N_19278);
or U20316 (N_20316,N_19323,N_19336);
and U20317 (N_20317,N_19842,N_19839);
and U20318 (N_20318,N_19973,N_19661);
xor U20319 (N_20319,N_19772,N_19664);
nand U20320 (N_20320,N_19451,N_19807);
and U20321 (N_20321,N_19335,N_19865);
nor U20322 (N_20322,N_19272,N_19575);
or U20323 (N_20323,N_19095,N_19887);
xnor U20324 (N_20324,N_19479,N_19015);
nor U20325 (N_20325,N_19041,N_19648);
xnor U20326 (N_20326,N_19609,N_19378);
nand U20327 (N_20327,N_19221,N_19915);
or U20328 (N_20328,N_19399,N_19508);
or U20329 (N_20329,N_19200,N_19151);
or U20330 (N_20330,N_19211,N_19244);
xor U20331 (N_20331,N_19532,N_19562);
nor U20332 (N_20332,N_19429,N_19809);
or U20333 (N_20333,N_19580,N_19789);
xor U20334 (N_20334,N_19155,N_19927);
and U20335 (N_20335,N_19481,N_19675);
or U20336 (N_20336,N_19031,N_19269);
nor U20337 (N_20337,N_19751,N_19895);
nand U20338 (N_20338,N_19877,N_19908);
nor U20339 (N_20339,N_19235,N_19507);
or U20340 (N_20340,N_19955,N_19773);
nor U20341 (N_20341,N_19523,N_19653);
and U20342 (N_20342,N_19744,N_19040);
nand U20343 (N_20343,N_19026,N_19835);
and U20344 (N_20344,N_19806,N_19747);
or U20345 (N_20345,N_19363,N_19176);
or U20346 (N_20346,N_19892,N_19587);
xor U20347 (N_20347,N_19900,N_19265);
nand U20348 (N_20348,N_19833,N_19714);
or U20349 (N_20349,N_19684,N_19111);
xnor U20350 (N_20350,N_19418,N_19928);
or U20351 (N_20351,N_19110,N_19419);
xor U20352 (N_20352,N_19470,N_19607);
nor U20353 (N_20353,N_19427,N_19589);
xnor U20354 (N_20354,N_19140,N_19924);
nand U20355 (N_20355,N_19044,N_19707);
nor U20356 (N_20356,N_19099,N_19993);
or U20357 (N_20357,N_19134,N_19257);
nor U20358 (N_20358,N_19819,N_19937);
nand U20359 (N_20359,N_19880,N_19642);
nor U20360 (N_20360,N_19671,N_19247);
and U20361 (N_20361,N_19056,N_19477);
and U20362 (N_20362,N_19795,N_19750);
and U20363 (N_20363,N_19520,N_19711);
nor U20364 (N_20364,N_19286,N_19455);
nor U20365 (N_20365,N_19205,N_19598);
and U20366 (N_20366,N_19901,N_19888);
nor U20367 (N_20367,N_19783,N_19590);
and U20368 (N_20368,N_19132,N_19382);
or U20369 (N_20369,N_19261,N_19570);
nor U20370 (N_20370,N_19267,N_19309);
nor U20371 (N_20371,N_19776,N_19958);
or U20372 (N_20372,N_19828,N_19009);
and U20373 (N_20373,N_19662,N_19238);
xnor U20374 (N_20374,N_19822,N_19321);
nor U20375 (N_20375,N_19165,N_19355);
xor U20376 (N_20376,N_19431,N_19274);
xnor U20377 (N_20377,N_19597,N_19921);
nand U20378 (N_20378,N_19486,N_19108);
xnor U20379 (N_20379,N_19341,N_19380);
xor U20380 (N_20380,N_19917,N_19820);
and U20381 (N_20381,N_19815,N_19911);
nand U20382 (N_20382,N_19164,N_19298);
or U20383 (N_20383,N_19371,N_19957);
or U20384 (N_20384,N_19139,N_19204);
and U20385 (N_20385,N_19345,N_19046);
nand U20386 (N_20386,N_19326,N_19849);
nor U20387 (N_20387,N_19899,N_19500);
and U20388 (N_20388,N_19726,N_19414);
nand U20389 (N_20389,N_19295,N_19779);
or U20390 (N_20390,N_19069,N_19458);
nor U20391 (N_20391,N_19219,N_19461);
xor U20392 (N_20392,N_19312,N_19534);
xnor U20393 (N_20393,N_19241,N_19629);
xnor U20394 (N_20394,N_19163,N_19933);
nand U20395 (N_20395,N_19248,N_19471);
or U20396 (N_20396,N_19413,N_19049);
or U20397 (N_20397,N_19208,N_19421);
or U20398 (N_20398,N_19422,N_19584);
nand U20399 (N_20399,N_19071,N_19476);
xnor U20400 (N_20400,N_19932,N_19987);
or U20401 (N_20401,N_19347,N_19364);
or U20402 (N_20402,N_19220,N_19161);
xnor U20403 (N_20403,N_19337,N_19646);
nand U20404 (N_20404,N_19686,N_19218);
or U20405 (N_20405,N_19129,N_19388);
nor U20406 (N_20406,N_19145,N_19568);
nor U20407 (N_20407,N_19390,N_19782);
or U20408 (N_20408,N_19752,N_19016);
or U20409 (N_20409,N_19159,N_19231);
or U20410 (N_20410,N_19325,N_19535);
nor U20411 (N_20411,N_19068,N_19890);
or U20412 (N_20412,N_19745,N_19525);
or U20413 (N_20413,N_19403,N_19260);
nand U20414 (N_20414,N_19332,N_19763);
xor U20415 (N_20415,N_19801,N_19989);
or U20416 (N_20416,N_19251,N_19704);
nor U20417 (N_20417,N_19357,N_19001);
nor U20418 (N_20418,N_19082,N_19424);
and U20419 (N_20419,N_19384,N_19301);
or U20420 (N_20420,N_19756,N_19945);
xnor U20421 (N_20421,N_19510,N_19785);
nor U20422 (N_20422,N_19770,N_19524);
nor U20423 (N_20423,N_19579,N_19907);
nor U20424 (N_20424,N_19817,N_19442);
or U20425 (N_20425,N_19319,N_19894);
and U20426 (N_20426,N_19680,N_19376);
or U20427 (N_20427,N_19765,N_19889);
nand U20428 (N_20428,N_19473,N_19766);
nand U20429 (N_20429,N_19386,N_19683);
xnor U20430 (N_20430,N_19692,N_19660);
and U20431 (N_20431,N_19566,N_19626);
or U20432 (N_20432,N_19207,N_19366);
nand U20433 (N_20433,N_19158,N_19702);
or U20434 (N_20434,N_19435,N_19832);
xor U20435 (N_20435,N_19679,N_19361);
nand U20436 (N_20436,N_19804,N_19619);
nor U20437 (N_20437,N_19294,N_19258);
or U20438 (N_20438,N_19604,N_19449);
and U20439 (N_20439,N_19093,N_19407);
xor U20440 (N_20440,N_19790,N_19829);
nand U20441 (N_20441,N_19117,N_19196);
or U20442 (N_20442,N_19559,N_19182);
nor U20443 (N_20443,N_19406,N_19914);
nor U20444 (N_20444,N_19391,N_19128);
xnor U20445 (N_20445,N_19465,N_19594);
or U20446 (N_20446,N_19284,N_19385);
xnor U20447 (N_20447,N_19344,N_19338);
nor U20448 (N_20448,N_19398,N_19583);
or U20449 (N_20449,N_19613,N_19732);
nand U20450 (N_20450,N_19019,N_19030);
nor U20451 (N_20451,N_19138,N_19610);
nor U20452 (N_20452,N_19254,N_19611);
xnor U20453 (N_20453,N_19627,N_19930);
and U20454 (N_20454,N_19222,N_19288);
or U20455 (N_20455,N_19669,N_19420);
nand U20456 (N_20456,N_19854,N_19359);
nand U20457 (N_20457,N_19910,N_19678);
nand U20458 (N_20458,N_19984,N_19061);
nor U20459 (N_20459,N_19079,N_19864);
or U20460 (N_20460,N_19253,N_19396);
or U20461 (N_20461,N_19003,N_19891);
xnor U20462 (N_20462,N_19761,N_19658);
nand U20463 (N_20463,N_19529,N_19628);
nand U20464 (N_20464,N_19893,N_19290);
xnor U20465 (N_20465,N_19087,N_19593);
and U20466 (N_20466,N_19433,N_19408);
xor U20467 (N_20467,N_19372,N_19640);
nor U20468 (N_20468,N_19062,N_19146);
and U20469 (N_20469,N_19897,N_19438);
nand U20470 (N_20470,N_19981,N_19968);
and U20471 (N_20471,N_19952,N_19737);
xnor U20472 (N_20472,N_19972,N_19518);
nor U20473 (N_20473,N_19631,N_19270);
nor U20474 (N_20474,N_19331,N_19739);
nand U20475 (N_20475,N_19223,N_19050);
xor U20476 (N_20476,N_19273,N_19578);
and U20477 (N_20477,N_19115,N_19992);
and U20478 (N_20478,N_19691,N_19035);
or U20479 (N_20479,N_19109,N_19755);
and U20480 (N_20480,N_19652,N_19723);
xor U20481 (N_20481,N_19271,N_19285);
nand U20482 (N_20482,N_19700,N_19688);
xor U20483 (N_20483,N_19170,N_19620);
nand U20484 (N_20484,N_19283,N_19246);
nand U20485 (N_20485,N_19722,N_19922);
or U20486 (N_20486,N_19576,N_19037);
or U20487 (N_20487,N_19292,N_19374);
xnor U20488 (N_20488,N_19342,N_19467);
nand U20489 (N_20489,N_19676,N_19303);
or U20490 (N_20490,N_19157,N_19402);
or U20491 (N_20491,N_19025,N_19088);
xor U20492 (N_20492,N_19397,N_19174);
and U20493 (N_20493,N_19599,N_19647);
nand U20494 (N_20494,N_19699,N_19941);
or U20495 (N_20495,N_19137,N_19047);
xor U20496 (N_20496,N_19812,N_19796);
nor U20497 (N_20497,N_19874,N_19931);
nand U20498 (N_20498,N_19728,N_19624);
nand U20499 (N_20499,N_19605,N_19123);
and U20500 (N_20500,N_19885,N_19911);
nor U20501 (N_20501,N_19350,N_19095);
and U20502 (N_20502,N_19293,N_19395);
xor U20503 (N_20503,N_19981,N_19124);
xnor U20504 (N_20504,N_19188,N_19851);
and U20505 (N_20505,N_19976,N_19716);
nor U20506 (N_20506,N_19862,N_19619);
or U20507 (N_20507,N_19798,N_19513);
and U20508 (N_20508,N_19143,N_19117);
and U20509 (N_20509,N_19648,N_19775);
or U20510 (N_20510,N_19410,N_19296);
nor U20511 (N_20511,N_19127,N_19754);
or U20512 (N_20512,N_19981,N_19817);
nand U20513 (N_20513,N_19318,N_19722);
and U20514 (N_20514,N_19491,N_19999);
xnor U20515 (N_20515,N_19570,N_19857);
xor U20516 (N_20516,N_19132,N_19017);
or U20517 (N_20517,N_19393,N_19951);
or U20518 (N_20518,N_19593,N_19861);
or U20519 (N_20519,N_19229,N_19124);
nor U20520 (N_20520,N_19885,N_19953);
nand U20521 (N_20521,N_19226,N_19196);
and U20522 (N_20522,N_19683,N_19907);
and U20523 (N_20523,N_19540,N_19285);
xnor U20524 (N_20524,N_19746,N_19692);
and U20525 (N_20525,N_19469,N_19895);
and U20526 (N_20526,N_19759,N_19001);
or U20527 (N_20527,N_19400,N_19899);
nand U20528 (N_20528,N_19191,N_19098);
nor U20529 (N_20529,N_19507,N_19505);
and U20530 (N_20530,N_19743,N_19955);
and U20531 (N_20531,N_19757,N_19265);
xor U20532 (N_20532,N_19638,N_19213);
or U20533 (N_20533,N_19194,N_19442);
xnor U20534 (N_20534,N_19674,N_19859);
nand U20535 (N_20535,N_19859,N_19136);
or U20536 (N_20536,N_19891,N_19226);
or U20537 (N_20537,N_19013,N_19945);
xor U20538 (N_20538,N_19996,N_19533);
and U20539 (N_20539,N_19853,N_19536);
xnor U20540 (N_20540,N_19297,N_19474);
nand U20541 (N_20541,N_19061,N_19637);
nand U20542 (N_20542,N_19966,N_19729);
or U20543 (N_20543,N_19349,N_19319);
and U20544 (N_20544,N_19312,N_19651);
nand U20545 (N_20545,N_19986,N_19751);
nand U20546 (N_20546,N_19301,N_19605);
and U20547 (N_20547,N_19731,N_19010);
nand U20548 (N_20548,N_19311,N_19134);
nand U20549 (N_20549,N_19102,N_19399);
and U20550 (N_20550,N_19877,N_19868);
xor U20551 (N_20551,N_19817,N_19375);
and U20552 (N_20552,N_19839,N_19128);
and U20553 (N_20553,N_19418,N_19009);
xor U20554 (N_20554,N_19238,N_19341);
and U20555 (N_20555,N_19241,N_19694);
nand U20556 (N_20556,N_19649,N_19393);
xnor U20557 (N_20557,N_19434,N_19972);
xnor U20558 (N_20558,N_19751,N_19837);
xnor U20559 (N_20559,N_19568,N_19104);
nand U20560 (N_20560,N_19899,N_19389);
nand U20561 (N_20561,N_19588,N_19168);
nand U20562 (N_20562,N_19810,N_19821);
or U20563 (N_20563,N_19866,N_19113);
nor U20564 (N_20564,N_19648,N_19696);
or U20565 (N_20565,N_19206,N_19529);
and U20566 (N_20566,N_19679,N_19873);
or U20567 (N_20567,N_19682,N_19669);
nand U20568 (N_20568,N_19871,N_19775);
xnor U20569 (N_20569,N_19270,N_19778);
or U20570 (N_20570,N_19864,N_19938);
and U20571 (N_20571,N_19354,N_19066);
nor U20572 (N_20572,N_19954,N_19083);
nor U20573 (N_20573,N_19276,N_19227);
and U20574 (N_20574,N_19872,N_19129);
nor U20575 (N_20575,N_19689,N_19035);
nand U20576 (N_20576,N_19739,N_19309);
nand U20577 (N_20577,N_19948,N_19078);
nand U20578 (N_20578,N_19523,N_19488);
nor U20579 (N_20579,N_19650,N_19357);
nor U20580 (N_20580,N_19312,N_19832);
xor U20581 (N_20581,N_19198,N_19842);
and U20582 (N_20582,N_19524,N_19739);
or U20583 (N_20583,N_19748,N_19453);
nand U20584 (N_20584,N_19238,N_19670);
xor U20585 (N_20585,N_19551,N_19307);
and U20586 (N_20586,N_19962,N_19868);
and U20587 (N_20587,N_19178,N_19101);
and U20588 (N_20588,N_19937,N_19294);
nand U20589 (N_20589,N_19791,N_19481);
or U20590 (N_20590,N_19367,N_19591);
xor U20591 (N_20591,N_19974,N_19515);
or U20592 (N_20592,N_19367,N_19582);
and U20593 (N_20593,N_19398,N_19743);
nor U20594 (N_20594,N_19777,N_19191);
or U20595 (N_20595,N_19537,N_19278);
nand U20596 (N_20596,N_19497,N_19654);
and U20597 (N_20597,N_19283,N_19461);
nor U20598 (N_20598,N_19722,N_19331);
nor U20599 (N_20599,N_19449,N_19717);
nor U20600 (N_20600,N_19039,N_19301);
nand U20601 (N_20601,N_19841,N_19165);
or U20602 (N_20602,N_19718,N_19178);
and U20603 (N_20603,N_19960,N_19319);
xnor U20604 (N_20604,N_19732,N_19406);
or U20605 (N_20605,N_19294,N_19625);
or U20606 (N_20606,N_19218,N_19364);
nor U20607 (N_20607,N_19079,N_19268);
nand U20608 (N_20608,N_19883,N_19301);
and U20609 (N_20609,N_19183,N_19296);
nand U20610 (N_20610,N_19349,N_19045);
xnor U20611 (N_20611,N_19768,N_19238);
xor U20612 (N_20612,N_19231,N_19032);
nand U20613 (N_20613,N_19568,N_19949);
nand U20614 (N_20614,N_19973,N_19931);
nand U20615 (N_20615,N_19023,N_19558);
nor U20616 (N_20616,N_19994,N_19851);
xor U20617 (N_20617,N_19162,N_19928);
xnor U20618 (N_20618,N_19932,N_19229);
or U20619 (N_20619,N_19948,N_19263);
nor U20620 (N_20620,N_19764,N_19164);
xor U20621 (N_20621,N_19542,N_19341);
nand U20622 (N_20622,N_19063,N_19548);
nor U20623 (N_20623,N_19911,N_19430);
and U20624 (N_20624,N_19921,N_19314);
xor U20625 (N_20625,N_19391,N_19628);
nor U20626 (N_20626,N_19121,N_19708);
and U20627 (N_20627,N_19720,N_19606);
xnor U20628 (N_20628,N_19951,N_19930);
nor U20629 (N_20629,N_19426,N_19028);
xor U20630 (N_20630,N_19055,N_19007);
nand U20631 (N_20631,N_19066,N_19008);
or U20632 (N_20632,N_19975,N_19651);
or U20633 (N_20633,N_19187,N_19931);
nor U20634 (N_20634,N_19431,N_19018);
or U20635 (N_20635,N_19247,N_19103);
xor U20636 (N_20636,N_19564,N_19381);
nor U20637 (N_20637,N_19904,N_19974);
or U20638 (N_20638,N_19808,N_19390);
nor U20639 (N_20639,N_19206,N_19823);
nand U20640 (N_20640,N_19649,N_19865);
xor U20641 (N_20641,N_19234,N_19499);
xor U20642 (N_20642,N_19893,N_19912);
nand U20643 (N_20643,N_19038,N_19689);
or U20644 (N_20644,N_19139,N_19807);
nand U20645 (N_20645,N_19611,N_19157);
nand U20646 (N_20646,N_19181,N_19824);
and U20647 (N_20647,N_19881,N_19729);
and U20648 (N_20648,N_19593,N_19917);
xor U20649 (N_20649,N_19491,N_19608);
or U20650 (N_20650,N_19836,N_19460);
nor U20651 (N_20651,N_19204,N_19832);
and U20652 (N_20652,N_19265,N_19229);
xnor U20653 (N_20653,N_19517,N_19252);
nor U20654 (N_20654,N_19501,N_19832);
xnor U20655 (N_20655,N_19517,N_19388);
and U20656 (N_20656,N_19976,N_19271);
nand U20657 (N_20657,N_19522,N_19856);
nor U20658 (N_20658,N_19031,N_19257);
and U20659 (N_20659,N_19290,N_19956);
or U20660 (N_20660,N_19509,N_19552);
nand U20661 (N_20661,N_19756,N_19234);
nand U20662 (N_20662,N_19575,N_19294);
or U20663 (N_20663,N_19581,N_19715);
or U20664 (N_20664,N_19181,N_19902);
and U20665 (N_20665,N_19080,N_19204);
xor U20666 (N_20666,N_19041,N_19099);
or U20667 (N_20667,N_19382,N_19512);
nand U20668 (N_20668,N_19554,N_19909);
xnor U20669 (N_20669,N_19301,N_19962);
and U20670 (N_20670,N_19677,N_19305);
nor U20671 (N_20671,N_19301,N_19956);
and U20672 (N_20672,N_19902,N_19113);
nand U20673 (N_20673,N_19391,N_19569);
nor U20674 (N_20674,N_19909,N_19878);
xor U20675 (N_20675,N_19319,N_19594);
xnor U20676 (N_20676,N_19055,N_19161);
xnor U20677 (N_20677,N_19504,N_19233);
xnor U20678 (N_20678,N_19383,N_19443);
or U20679 (N_20679,N_19023,N_19998);
nor U20680 (N_20680,N_19595,N_19905);
or U20681 (N_20681,N_19450,N_19867);
nor U20682 (N_20682,N_19058,N_19904);
nand U20683 (N_20683,N_19272,N_19054);
or U20684 (N_20684,N_19613,N_19676);
and U20685 (N_20685,N_19732,N_19350);
or U20686 (N_20686,N_19724,N_19177);
nor U20687 (N_20687,N_19176,N_19624);
nor U20688 (N_20688,N_19803,N_19247);
xor U20689 (N_20689,N_19005,N_19380);
and U20690 (N_20690,N_19454,N_19134);
and U20691 (N_20691,N_19596,N_19923);
nor U20692 (N_20692,N_19193,N_19987);
xor U20693 (N_20693,N_19377,N_19703);
and U20694 (N_20694,N_19038,N_19058);
nor U20695 (N_20695,N_19738,N_19317);
nor U20696 (N_20696,N_19744,N_19556);
nand U20697 (N_20697,N_19436,N_19117);
nor U20698 (N_20698,N_19836,N_19247);
nand U20699 (N_20699,N_19354,N_19435);
and U20700 (N_20700,N_19905,N_19103);
or U20701 (N_20701,N_19646,N_19721);
nand U20702 (N_20702,N_19337,N_19050);
nor U20703 (N_20703,N_19967,N_19882);
and U20704 (N_20704,N_19503,N_19618);
nor U20705 (N_20705,N_19115,N_19256);
nand U20706 (N_20706,N_19580,N_19637);
or U20707 (N_20707,N_19563,N_19474);
and U20708 (N_20708,N_19503,N_19638);
xor U20709 (N_20709,N_19956,N_19637);
or U20710 (N_20710,N_19985,N_19300);
xor U20711 (N_20711,N_19679,N_19176);
and U20712 (N_20712,N_19127,N_19392);
nor U20713 (N_20713,N_19432,N_19794);
or U20714 (N_20714,N_19201,N_19728);
nor U20715 (N_20715,N_19943,N_19880);
or U20716 (N_20716,N_19592,N_19820);
or U20717 (N_20717,N_19382,N_19180);
or U20718 (N_20718,N_19212,N_19958);
and U20719 (N_20719,N_19339,N_19145);
xnor U20720 (N_20720,N_19633,N_19052);
nor U20721 (N_20721,N_19719,N_19683);
xnor U20722 (N_20722,N_19393,N_19255);
xnor U20723 (N_20723,N_19068,N_19390);
nor U20724 (N_20724,N_19462,N_19171);
xnor U20725 (N_20725,N_19476,N_19758);
nor U20726 (N_20726,N_19036,N_19472);
or U20727 (N_20727,N_19803,N_19814);
xnor U20728 (N_20728,N_19439,N_19381);
or U20729 (N_20729,N_19598,N_19039);
nor U20730 (N_20730,N_19649,N_19595);
nor U20731 (N_20731,N_19887,N_19286);
and U20732 (N_20732,N_19134,N_19933);
xnor U20733 (N_20733,N_19375,N_19823);
nor U20734 (N_20734,N_19301,N_19570);
nand U20735 (N_20735,N_19237,N_19716);
nor U20736 (N_20736,N_19196,N_19810);
nand U20737 (N_20737,N_19595,N_19049);
nand U20738 (N_20738,N_19214,N_19952);
or U20739 (N_20739,N_19043,N_19931);
nor U20740 (N_20740,N_19645,N_19973);
xnor U20741 (N_20741,N_19636,N_19056);
xor U20742 (N_20742,N_19831,N_19115);
nor U20743 (N_20743,N_19368,N_19574);
or U20744 (N_20744,N_19891,N_19394);
xor U20745 (N_20745,N_19929,N_19356);
and U20746 (N_20746,N_19524,N_19421);
nand U20747 (N_20747,N_19675,N_19497);
nand U20748 (N_20748,N_19176,N_19316);
xnor U20749 (N_20749,N_19292,N_19459);
nor U20750 (N_20750,N_19994,N_19002);
nor U20751 (N_20751,N_19970,N_19798);
or U20752 (N_20752,N_19864,N_19933);
nor U20753 (N_20753,N_19096,N_19543);
xnor U20754 (N_20754,N_19137,N_19494);
or U20755 (N_20755,N_19330,N_19770);
or U20756 (N_20756,N_19986,N_19712);
xnor U20757 (N_20757,N_19910,N_19668);
nor U20758 (N_20758,N_19080,N_19052);
and U20759 (N_20759,N_19919,N_19057);
nand U20760 (N_20760,N_19513,N_19078);
nand U20761 (N_20761,N_19474,N_19878);
or U20762 (N_20762,N_19082,N_19587);
nand U20763 (N_20763,N_19223,N_19396);
nor U20764 (N_20764,N_19577,N_19376);
xnor U20765 (N_20765,N_19623,N_19206);
nand U20766 (N_20766,N_19206,N_19108);
xnor U20767 (N_20767,N_19140,N_19317);
nor U20768 (N_20768,N_19186,N_19713);
xor U20769 (N_20769,N_19936,N_19318);
and U20770 (N_20770,N_19033,N_19122);
and U20771 (N_20771,N_19859,N_19345);
xor U20772 (N_20772,N_19191,N_19268);
nor U20773 (N_20773,N_19295,N_19541);
xnor U20774 (N_20774,N_19325,N_19454);
nand U20775 (N_20775,N_19549,N_19468);
and U20776 (N_20776,N_19499,N_19199);
nor U20777 (N_20777,N_19042,N_19277);
and U20778 (N_20778,N_19999,N_19018);
nand U20779 (N_20779,N_19838,N_19424);
xnor U20780 (N_20780,N_19040,N_19467);
nand U20781 (N_20781,N_19134,N_19833);
or U20782 (N_20782,N_19813,N_19479);
and U20783 (N_20783,N_19666,N_19600);
nor U20784 (N_20784,N_19623,N_19866);
and U20785 (N_20785,N_19629,N_19811);
xor U20786 (N_20786,N_19173,N_19602);
nor U20787 (N_20787,N_19295,N_19485);
or U20788 (N_20788,N_19187,N_19775);
nand U20789 (N_20789,N_19504,N_19221);
and U20790 (N_20790,N_19519,N_19567);
nand U20791 (N_20791,N_19118,N_19937);
and U20792 (N_20792,N_19225,N_19750);
nand U20793 (N_20793,N_19774,N_19941);
nand U20794 (N_20794,N_19587,N_19798);
nand U20795 (N_20795,N_19064,N_19133);
nand U20796 (N_20796,N_19098,N_19520);
and U20797 (N_20797,N_19214,N_19018);
and U20798 (N_20798,N_19785,N_19148);
or U20799 (N_20799,N_19294,N_19898);
or U20800 (N_20800,N_19455,N_19626);
or U20801 (N_20801,N_19618,N_19282);
and U20802 (N_20802,N_19587,N_19803);
nor U20803 (N_20803,N_19498,N_19821);
and U20804 (N_20804,N_19509,N_19516);
or U20805 (N_20805,N_19019,N_19271);
and U20806 (N_20806,N_19033,N_19263);
and U20807 (N_20807,N_19615,N_19657);
nand U20808 (N_20808,N_19505,N_19989);
nand U20809 (N_20809,N_19447,N_19275);
nor U20810 (N_20810,N_19851,N_19944);
nand U20811 (N_20811,N_19632,N_19958);
nand U20812 (N_20812,N_19022,N_19709);
xnor U20813 (N_20813,N_19187,N_19223);
or U20814 (N_20814,N_19128,N_19747);
or U20815 (N_20815,N_19263,N_19155);
and U20816 (N_20816,N_19304,N_19330);
nand U20817 (N_20817,N_19505,N_19775);
nand U20818 (N_20818,N_19061,N_19563);
xnor U20819 (N_20819,N_19890,N_19720);
and U20820 (N_20820,N_19064,N_19337);
or U20821 (N_20821,N_19847,N_19104);
or U20822 (N_20822,N_19322,N_19459);
xnor U20823 (N_20823,N_19608,N_19687);
nor U20824 (N_20824,N_19811,N_19130);
or U20825 (N_20825,N_19742,N_19197);
or U20826 (N_20826,N_19758,N_19532);
nor U20827 (N_20827,N_19795,N_19121);
or U20828 (N_20828,N_19913,N_19498);
and U20829 (N_20829,N_19928,N_19969);
nor U20830 (N_20830,N_19804,N_19664);
xnor U20831 (N_20831,N_19957,N_19106);
xor U20832 (N_20832,N_19270,N_19967);
or U20833 (N_20833,N_19210,N_19645);
and U20834 (N_20834,N_19446,N_19792);
nor U20835 (N_20835,N_19041,N_19221);
or U20836 (N_20836,N_19802,N_19344);
nor U20837 (N_20837,N_19775,N_19670);
nor U20838 (N_20838,N_19466,N_19686);
or U20839 (N_20839,N_19135,N_19861);
nor U20840 (N_20840,N_19427,N_19501);
nor U20841 (N_20841,N_19280,N_19060);
nand U20842 (N_20842,N_19192,N_19502);
xnor U20843 (N_20843,N_19493,N_19441);
nor U20844 (N_20844,N_19391,N_19941);
and U20845 (N_20845,N_19823,N_19948);
or U20846 (N_20846,N_19953,N_19620);
and U20847 (N_20847,N_19016,N_19029);
or U20848 (N_20848,N_19522,N_19786);
nand U20849 (N_20849,N_19320,N_19474);
or U20850 (N_20850,N_19062,N_19007);
xor U20851 (N_20851,N_19385,N_19153);
nand U20852 (N_20852,N_19886,N_19546);
nor U20853 (N_20853,N_19946,N_19948);
or U20854 (N_20854,N_19991,N_19177);
nand U20855 (N_20855,N_19791,N_19530);
nand U20856 (N_20856,N_19182,N_19693);
nand U20857 (N_20857,N_19509,N_19340);
and U20858 (N_20858,N_19757,N_19625);
nand U20859 (N_20859,N_19697,N_19362);
nor U20860 (N_20860,N_19434,N_19688);
nand U20861 (N_20861,N_19828,N_19908);
nor U20862 (N_20862,N_19817,N_19444);
and U20863 (N_20863,N_19051,N_19391);
nand U20864 (N_20864,N_19438,N_19050);
and U20865 (N_20865,N_19871,N_19459);
nor U20866 (N_20866,N_19616,N_19825);
nor U20867 (N_20867,N_19429,N_19405);
xnor U20868 (N_20868,N_19180,N_19372);
nor U20869 (N_20869,N_19810,N_19080);
nor U20870 (N_20870,N_19200,N_19463);
nand U20871 (N_20871,N_19733,N_19425);
nor U20872 (N_20872,N_19031,N_19852);
nand U20873 (N_20873,N_19698,N_19842);
xnor U20874 (N_20874,N_19510,N_19492);
or U20875 (N_20875,N_19005,N_19445);
nand U20876 (N_20876,N_19414,N_19257);
and U20877 (N_20877,N_19160,N_19744);
nand U20878 (N_20878,N_19997,N_19819);
and U20879 (N_20879,N_19541,N_19074);
or U20880 (N_20880,N_19129,N_19992);
or U20881 (N_20881,N_19905,N_19824);
nand U20882 (N_20882,N_19667,N_19160);
or U20883 (N_20883,N_19778,N_19879);
nand U20884 (N_20884,N_19792,N_19463);
or U20885 (N_20885,N_19406,N_19945);
xor U20886 (N_20886,N_19772,N_19536);
nor U20887 (N_20887,N_19910,N_19152);
nor U20888 (N_20888,N_19858,N_19811);
xnor U20889 (N_20889,N_19460,N_19921);
xor U20890 (N_20890,N_19668,N_19252);
and U20891 (N_20891,N_19265,N_19831);
xor U20892 (N_20892,N_19650,N_19651);
xnor U20893 (N_20893,N_19475,N_19097);
and U20894 (N_20894,N_19681,N_19750);
xor U20895 (N_20895,N_19666,N_19833);
nand U20896 (N_20896,N_19702,N_19715);
nor U20897 (N_20897,N_19459,N_19079);
xnor U20898 (N_20898,N_19821,N_19947);
xor U20899 (N_20899,N_19956,N_19653);
and U20900 (N_20900,N_19147,N_19402);
xnor U20901 (N_20901,N_19964,N_19026);
nor U20902 (N_20902,N_19904,N_19406);
nand U20903 (N_20903,N_19037,N_19405);
xnor U20904 (N_20904,N_19079,N_19866);
xor U20905 (N_20905,N_19867,N_19529);
xor U20906 (N_20906,N_19696,N_19460);
or U20907 (N_20907,N_19621,N_19595);
and U20908 (N_20908,N_19647,N_19842);
nand U20909 (N_20909,N_19500,N_19733);
or U20910 (N_20910,N_19364,N_19338);
and U20911 (N_20911,N_19430,N_19106);
xor U20912 (N_20912,N_19489,N_19956);
nand U20913 (N_20913,N_19964,N_19972);
or U20914 (N_20914,N_19423,N_19044);
nor U20915 (N_20915,N_19755,N_19444);
nand U20916 (N_20916,N_19883,N_19825);
nand U20917 (N_20917,N_19147,N_19786);
and U20918 (N_20918,N_19730,N_19913);
and U20919 (N_20919,N_19075,N_19154);
and U20920 (N_20920,N_19483,N_19368);
nand U20921 (N_20921,N_19052,N_19171);
and U20922 (N_20922,N_19944,N_19506);
nor U20923 (N_20923,N_19905,N_19665);
xnor U20924 (N_20924,N_19648,N_19171);
nor U20925 (N_20925,N_19791,N_19675);
and U20926 (N_20926,N_19132,N_19437);
xnor U20927 (N_20927,N_19338,N_19734);
nor U20928 (N_20928,N_19591,N_19037);
and U20929 (N_20929,N_19678,N_19337);
xor U20930 (N_20930,N_19515,N_19770);
nand U20931 (N_20931,N_19820,N_19795);
xor U20932 (N_20932,N_19045,N_19396);
nand U20933 (N_20933,N_19335,N_19013);
nand U20934 (N_20934,N_19945,N_19617);
nand U20935 (N_20935,N_19725,N_19882);
xnor U20936 (N_20936,N_19800,N_19594);
and U20937 (N_20937,N_19266,N_19102);
or U20938 (N_20938,N_19712,N_19910);
or U20939 (N_20939,N_19644,N_19389);
and U20940 (N_20940,N_19109,N_19609);
or U20941 (N_20941,N_19891,N_19527);
nor U20942 (N_20942,N_19338,N_19309);
nor U20943 (N_20943,N_19716,N_19330);
nand U20944 (N_20944,N_19650,N_19866);
nand U20945 (N_20945,N_19874,N_19422);
or U20946 (N_20946,N_19229,N_19446);
nand U20947 (N_20947,N_19043,N_19404);
or U20948 (N_20948,N_19728,N_19875);
and U20949 (N_20949,N_19870,N_19012);
xnor U20950 (N_20950,N_19577,N_19268);
xor U20951 (N_20951,N_19439,N_19622);
nand U20952 (N_20952,N_19123,N_19330);
xnor U20953 (N_20953,N_19907,N_19619);
xor U20954 (N_20954,N_19245,N_19513);
or U20955 (N_20955,N_19043,N_19371);
nand U20956 (N_20956,N_19410,N_19247);
nand U20957 (N_20957,N_19767,N_19273);
or U20958 (N_20958,N_19911,N_19648);
nand U20959 (N_20959,N_19168,N_19720);
or U20960 (N_20960,N_19168,N_19804);
xnor U20961 (N_20961,N_19359,N_19371);
nor U20962 (N_20962,N_19694,N_19648);
xnor U20963 (N_20963,N_19625,N_19800);
and U20964 (N_20964,N_19763,N_19004);
and U20965 (N_20965,N_19879,N_19653);
nor U20966 (N_20966,N_19413,N_19203);
xnor U20967 (N_20967,N_19487,N_19576);
nor U20968 (N_20968,N_19567,N_19866);
and U20969 (N_20969,N_19657,N_19920);
nand U20970 (N_20970,N_19496,N_19300);
nand U20971 (N_20971,N_19527,N_19248);
or U20972 (N_20972,N_19312,N_19464);
nand U20973 (N_20973,N_19972,N_19243);
nor U20974 (N_20974,N_19503,N_19947);
nand U20975 (N_20975,N_19780,N_19729);
xor U20976 (N_20976,N_19155,N_19048);
nand U20977 (N_20977,N_19977,N_19435);
and U20978 (N_20978,N_19743,N_19956);
nor U20979 (N_20979,N_19129,N_19132);
xnor U20980 (N_20980,N_19600,N_19381);
xor U20981 (N_20981,N_19677,N_19463);
or U20982 (N_20982,N_19687,N_19211);
nand U20983 (N_20983,N_19611,N_19650);
or U20984 (N_20984,N_19385,N_19111);
or U20985 (N_20985,N_19084,N_19009);
xnor U20986 (N_20986,N_19401,N_19486);
or U20987 (N_20987,N_19609,N_19500);
or U20988 (N_20988,N_19961,N_19755);
nand U20989 (N_20989,N_19184,N_19091);
or U20990 (N_20990,N_19446,N_19558);
and U20991 (N_20991,N_19548,N_19925);
xor U20992 (N_20992,N_19752,N_19755);
and U20993 (N_20993,N_19417,N_19267);
nor U20994 (N_20994,N_19128,N_19542);
or U20995 (N_20995,N_19968,N_19044);
or U20996 (N_20996,N_19281,N_19590);
nand U20997 (N_20997,N_19153,N_19900);
or U20998 (N_20998,N_19587,N_19529);
nor U20999 (N_20999,N_19381,N_19339);
and U21000 (N_21000,N_20019,N_20739);
nor U21001 (N_21001,N_20528,N_20843);
and U21002 (N_21002,N_20933,N_20507);
xor U21003 (N_21003,N_20883,N_20423);
xor U21004 (N_21004,N_20186,N_20181);
nor U21005 (N_21005,N_20666,N_20515);
xor U21006 (N_21006,N_20117,N_20301);
or U21007 (N_21007,N_20484,N_20101);
or U21008 (N_21008,N_20851,N_20300);
nor U21009 (N_21009,N_20605,N_20359);
xor U21010 (N_21010,N_20013,N_20552);
nand U21011 (N_21011,N_20789,N_20530);
or U21012 (N_21012,N_20800,N_20889);
nand U21013 (N_21013,N_20716,N_20398);
or U21014 (N_21014,N_20066,N_20505);
nor U21015 (N_21015,N_20120,N_20663);
and U21016 (N_21016,N_20430,N_20160);
and U21017 (N_21017,N_20339,N_20937);
nor U21018 (N_21018,N_20944,N_20641);
nand U21019 (N_21019,N_20306,N_20090);
nor U21020 (N_21020,N_20723,N_20224);
nand U21021 (N_21021,N_20654,N_20498);
and U21022 (N_21022,N_20676,N_20978);
nand U21023 (N_21023,N_20674,N_20499);
or U21024 (N_21024,N_20409,N_20341);
and U21025 (N_21025,N_20764,N_20936);
and U21026 (N_21026,N_20001,N_20993);
nor U21027 (N_21027,N_20111,N_20163);
nor U21028 (N_21028,N_20696,N_20023);
nand U21029 (N_21029,N_20678,N_20984);
or U21030 (N_21030,N_20620,N_20790);
xnor U21031 (N_21031,N_20832,N_20104);
or U21032 (N_21032,N_20872,N_20640);
nor U21033 (N_21033,N_20802,N_20730);
and U21034 (N_21034,N_20609,N_20879);
and U21035 (N_21035,N_20378,N_20237);
xnor U21036 (N_21036,N_20415,N_20837);
and U21037 (N_21037,N_20700,N_20814);
nand U21038 (N_21038,N_20619,N_20393);
nand U21039 (N_21039,N_20372,N_20475);
xnor U21040 (N_21040,N_20352,N_20292);
nor U21041 (N_21041,N_20154,N_20269);
xor U21042 (N_21042,N_20189,N_20848);
or U21043 (N_21043,N_20534,N_20840);
nand U21044 (N_21044,N_20895,N_20760);
xor U21045 (N_21045,N_20881,N_20436);
or U21046 (N_21046,N_20930,N_20131);
and U21047 (N_21047,N_20987,N_20769);
nor U21048 (N_21048,N_20738,N_20535);
xnor U21049 (N_21049,N_20321,N_20345);
nand U21050 (N_21050,N_20068,N_20035);
xor U21051 (N_21051,N_20860,N_20757);
or U21052 (N_21052,N_20869,N_20134);
and U21053 (N_21053,N_20586,N_20597);
xnor U21054 (N_21054,N_20956,N_20672);
nand U21055 (N_21055,N_20648,N_20222);
and U21056 (N_21056,N_20655,N_20278);
nand U21057 (N_21057,N_20329,N_20943);
and U21058 (N_21058,N_20681,N_20197);
or U21059 (N_21059,N_20839,N_20558);
nor U21060 (N_21060,N_20232,N_20245);
or U21061 (N_21061,N_20236,N_20582);
or U21062 (N_21062,N_20140,N_20317);
xor U21063 (N_21063,N_20491,N_20128);
nor U21064 (N_21064,N_20032,N_20501);
and U21065 (N_21065,N_20231,N_20756);
nor U21066 (N_21066,N_20038,N_20568);
and U21067 (N_21067,N_20497,N_20490);
nand U21068 (N_21068,N_20342,N_20434);
nand U21069 (N_21069,N_20504,N_20616);
nand U21070 (N_21070,N_20595,N_20974);
nor U21071 (N_21071,N_20272,N_20395);
nand U21072 (N_21072,N_20361,N_20809);
and U21073 (N_21073,N_20577,N_20847);
or U21074 (N_21074,N_20139,N_20334);
xor U21075 (N_21075,N_20824,N_20445);
and U21076 (N_21076,N_20218,N_20284);
xnor U21077 (N_21077,N_20366,N_20287);
nor U21078 (N_21078,N_20810,N_20248);
xor U21079 (N_21079,N_20382,N_20103);
nand U21080 (N_21080,N_20477,N_20147);
or U21081 (N_21081,N_20182,N_20752);
nand U21082 (N_21082,N_20251,N_20845);
xnor U21083 (N_21083,N_20625,N_20689);
or U21084 (N_21084,N_20755,N_20560);
xnor U21085 (N_21085,N_20375,N_20262);
xor U21086 (N_21086,N_20221,N_20999);
nor U21087 (N_21087,N_20325,N_20326);
and U21088 (N_21088,N_20673,N_20571);
or U21089 (N_21089,N_20135,N_20091);
xor U21090 (N_21090,N_20025,N_20940);
xnor U21091 (N_21091,N_20348,N_20400);
and U21092 (N_21092,N_20963,N_20816);
xor U21093 (N_21093,N_20281,N_20911);
nand U21094 (N_21094,N_20612,N_20142);
xor U21095 (N_21095,N_20618,N_20273);
and U21096 (N_21096,N_20804,N_20277);
and U21097 (N_21097,N_20539,N_20153);
or U21098 (N_21098,N_20788,N_20794);
nor U21099 (N_21099,N_20852,N_20912);
xor U21100 (N_21100,N_20034,N_20060);
or U21101 (N_21101,N_20947,N_20199);
and U21102 (N_21102,N_20132,N_20759);
nand U21103 (N_21103,N_20244,N_20242);
nand U21104 (N_21104,N_20355,N_20349);
xor U21105 (N_21105,N_20458,N_20149);
nor U21106 (N_21106,N_20097,N_20271);
xor U21107 (N_21107,N_20718,N_20874);
or U21108 (N_21108,N_20351,N_20067);
nand U21109 (N_21109,N_20180,N_20510);
and U21110 (N_21110,N_20122,N_20195);
and U21111 (N_21111,N_20059,N_20831);
nand U21112 (N_21112,N_20925,N_20511);
nand U21113 (N_21113,N_20124,N_20566);
or U21114 (N_21114,N_20315,N_20198);
and U21115 (N_21115,N_20688,N_20376);
or U21116 (N_21116,N_20692,N_20693);
nand U21117 (N_21117,N_20906,N_20112);
and U21118 (N_21118,N_20740,N_20404);
or U21119 (N_21119,N_20893,N_20184);
and U21120 (N_21120,N_20208,N_20424);
nand U21121 (N_21121,N_20216,N_20465);
xnor U21122 (N_21122,N_20836,N_20578);
nand U21123 (N_21123,N_20846,N_20460);
nand U21124 (N_21124,N_20885,N_20196);
xnor U21125 (N_21125,N_20997,N_20992);
xor U21126 (N_21126,N_20126,N_20431);
nor U21127 (N_21127,N_20468,N_20061);
or U21128 (N_21128,N_20623,N_20531);
xor U21129 (N_21129,N_20289,N_20801);
nand U21130 (N_21130,N_20686,N_20915);
nor U21131 (N_21131,N_20803,N_20288);
nor U21132 (N_21132,N_20259,N_20634);
nor U21133 (N_21133,N_20350,N_20447);
xnor U21134 (N_21134,N_20600,N_20996);
xnor U21135 (N_21135,N_20868,N_20642);
nand U21136 (N_21136,N_20178,N_20683);
xnor U21137 (N_21137,N_20585,N_20016);
xor U21138 (N_21138,N_20825,N_20783);
or U21139 (N_21139,N_20538,N_20588);
nor U21140 (N_21140,N_20024,N_20989);
nand U21141 (N_21141,N_20525,N_20190);
xor U21142 (N_21142,N_20435,N_20939);
and U21143 (N_21143,N_20367,N_20000);
and U21144 (N_21144,N_20778,N_20187);
or U21145 (N_21145,N_20591,N_20357);
or U21146 (N_21146,N_20448,N_20733);
or U21147 (N_21147,N_20108,N_20728);
nor U21148 (N_21148,N_20859,N_20381);
or U21149 (N_21149,N_20143,N_20631);
nand U21150 (N_21150,N_20865,N_20078);
and U21151 (N_21151,N_20514,N_20856);
nor U21152 (N_21152,N_20870,N_20611);
xnor U21153 (N_21153,N_20532,N_20659);
nand U21154 (N_21154,N_20008,N_20136);
and U21155 (N_21155,N_20524,N_20018);
nor U21156 (N_21156,N_20770,N_20286);
xor U21157 (N_21157,N_20384,N_20904);
and U21158 (N_21158,N_20841,N_20942);
nand U21159 (N_21159,N_20275,N_20308);
nor U21160 (N_21160,N_20369,N_20727);
nor U21161 (N_21161,N_20991,N_20455);
xor U21162 (N_21162,N_20373,N_20994);
nand U21163 (N_21163,N_20100,N_20335);
nor U21164 (N_21164,N_20826,N_20990);
nand U21165 (N_21165,N_20543,N_20529);
and U21166 (N_21166,N_20118,N_20720);
nand U21167 (N_21167,N_20356,N_20470);
or U21168 (N_21168,N_20622,N_20898);
nor U21169 (N_21169,N_20737,N_20383);
nand U21170 (N_21170,N_20170,N_20487);
or U21171 (N_21171,N_20453,N_20207);
or U21172 (N_21172,N_20314,N_20302);
or U21173 (N_21173,N_20233,N_20902);
xor U21174 (N_21174,N_20290,N_20776);
xnor U21175 (N_21175,N_20604,N_20711);
and U21176 (N_21176,N_20797,N_20370);
or U21177 (N_21177,N_20494,N_20316);
or U21178 (N_21178,N_20469,N_20639);
or U21179 (N_21179,N_20918,N_20110);
or U21180 (N_21180,N_20765,N_20704);
or U21181 (N_21181,N_20161,N_20046);
xnor U21182 (N_21182,N_20333,N_20037);
or U21183 (N_21183,N_20105,N_20402);
and U21184 (N_21184,N_20973,N_20405);
nand U21185 (N_21185,N_20806,N_20320);
nor U21186 (N_21186,N_20039,N_20238);
nand U21187 (N_21187,N_20175,N_20030);
and U21188 (N_21188,N_20512,N_20095);
nor U21189 (N_21189,N_20152,N_20975);
and U21190 (N_21190,N_20651,N_20133);
nor U21191 (N_21191,N_20960,N_20624);
nor U21192 (N_21192,N_20932,N_20953);
or U21193 (N_21193,N_20627,N_20478);
xnor U21194 (N_21194,N_20887,N_20466);
and U21195 (N_21195,N_20590,N_20541);
and U21196 (N_21196,N_20658,N_20421);
and U21197 (N_21197,N_20635,N_20959);
or U21198 (N_21198,N_20419,N_20736);
and U21199 (N_21199,N_20891,N_20336);
and U21200 (N_21200,N_20407,N_20970);
nor U21201 (N_21201,N_20422,N_20486);
nand U21202 (N_21202,N_20966,N_20265);
xnor U21203 (N_21203,N_20701,N_20495);
and U21204 (N_21204,N_20020,N_20863);
or U21205 (N_21205,N_20293,N_20483);
and U21206 (N_21206,N_20626,N_20012);
or U21207 (N_21207,N_20176,N_20690);
nor U21208 (N_21208,N_20146,N_20449);
xnor U21209 (N_21209,N_20828,N_20401);
xnor U21210 (N_21210,N_20165,N_20389);
or U21211 (N_21211,N_20123,N_20892);
and U21212 (N_21212,N_20557,N_20148);
or U21213 (N_21213,N_20785,N_20418);
nand U21214 (N_21214,N_20934,N_20650);
or U21215 (N_21215,N_20452,N_20884);
xnor U21216 (N_21216,N_20312,N_20669);
and U21217 (N_21217,N_20266,N_20710);
and U21218 (N_21218,N_20685,N_20766);
or U21219 (N_21219,N_20743,N_20227);
nor U21220 (N_21220,N_20522,N_20450);
nand U21221 (N_21221,N_20089,N_20645);
and U21222 (N_21222,N_20200,N_20417);
or U21223 (N_21223,N_20677,N_20744);
nand U21224 (N_21224,N_20559,N_20049);
xnor U21225 (N_21225,N_20721,N_20819);
nand U21226 (N_21226,N_20144,N_20513);
xor U21227 (N_21227,N_20753,N_20873);
nor U21228 (N_21228,N_20428,N_20949);
nand U21229 (N_21229,N_20235,N_20079);
nor U21230 (N_21230,N_20156,N_20900);
or U21231 (N_21231,N_20223,N_20081);
nor U21232 (N_21232,N_20201,N_20807);
nor U21233 (N_21233,N_20699,N_20496);
nor U21234 (N_21234,N_20391,N_20313);
xor U21235 (N_21235,N_20533,N_20749);
nand U21236 (N_21236,N_20877,N_20246);
nand U21237 (N_21237,N_20725,N_20561);
and U21238 (N_21238,N_20544,N_20680);
or U21239 (N_21239,N_20866,N_20798);
nand U21240 (N_21240,N_20691,N_20687);
nor U21241 (N_21241,N_20547,N_20976);
and U21242 (N_21242,N_20792,N_20026);
xnor U21243 (N_21243,N_20545,N_20412);
or U21244 (N_21244,N_20479,N_20109);
and U21245 (N_21245,N_20998,N_20368);
or U21246 (N_21246,N_20092,N_20416);
and U21247 (N_21247,N_20344,N_20094);
nor U21248 (N_21248,N_20827,N_20166);
xnor U21249 (N_21249,N_20489,N_20193);
nor U21250 (N_21250,N_20064,N_20444);
nor U21251 (N_21251,N_20927,N_20775);
nor U21252 (N_21252,N_20820,N_20957);
or U21253 (N_21253,N_20630,N_20594);
and U21254 (N_21254,N_20476,N_20053);
nor U21255 (N_21255,N_20550,N_20614);
and U21256 (N_21256,N_20474,N_20432);
nand U21257 (N_21257,N_20579,N_20296);
and U21258 (N_21258,N_20096,N_20439);
xor U21259 (N_21259,N_20665,N_20745);
and U21260 (N_21260,N_20502,N_20347);
or U21261 (N_21261,N_20573,N_20613);
xnor U21262 (N_21262,N_20041,N_20058);
and U21263 (N_21263,N_20537,N_20241);
and U21264 (N_21264,N_20280,N_20076);
nand U21265 (N_21265,N_20731,N_20572);
and U21266 (N_21266,N_20086,N_20211);
nor U21267 (N_21267,N_20955,N_20717);
nand U21268 (N_21268,N_20011,N_20871);
or U21269 (N_21269,N_20088,N_20901);
and U21270 (N_21270,N_20908,N_20517);
and U21271 (N_21271,N_20772,N_20986);
or U21272 (N_21272,N_20615,N_20337);
or U21273 (N_21273,N_20042,N_20172);
xor U21274 (N_21274,N_20768,N_20882);
nor U21275 (N_21275,N_20795,N_20243);
or U21276 (N_21276,N_20667,N_20903);
nand U21277 (N_21277,N_20980,N_20371);
nand U21278 (N_21278,N_20234,N_20250);
and U21279 (N_21279,N_20036,N_20386);
or U21280 (N_21280,N_20480,N_20228);
or U21281 (N_21281,N_20551,N_20295);
or U21282 (N_21282,N_20440,N_20782);
and U21283 (N_21283,N_20646,N_20821);
nand U21284 (N_21284,N_20861,N_20771);
nand U21285 (N_21285,N_20451,N_20397);
and U21286 (N_21286,N_20890,N_20212);
nor U21287 (N_21287,N_20328,N_20632);
nand U21288 (N_21288,N_20748,N_20601);
xnor U21289 (N_21289,N_20406,N_20931);
nand U21290 (N_21290,N_20917,N_20179);
xor U21291 (N_21291,N_20331,N_20130);
nor U21292 (N_21292,N_20093,N_20850);
or U21293 (N_21293,N_20506,N_20263);
nand U21294 (N_21294,N_20062,N_20719);
nor U21295 (N_21295,N_20805,N_20977);
or U21296 (N_21296,N_20214,N_20473);
nor U21297 (N_21297,N_20220,N_20379);
nand U21298 (N_21298,N_20299,N_20441);
xor U21299 (N_21299,N_20102,N_20022);
nor U21300 (N_21300,N_20569,N_20520);
and U21301 (N_21301,N_20077,N_20330);
xor U21302 (N_21302,N_20408,N_20461);
and U21303 (N_21303,N_20896,N_20009);
nor U21304 (N_21304,N_20675,N_20830);
nor U21305 (N_21305,N_20763,N_20938);
xnor U21306 (N_21306,N_20051,N_20968);
nand U21307 (N_21307,N_20607,N_20192);
and U21308 (N_21308,N_20399,N_20082);
and U21309 (N_21309,N_20387,N_20305);
xnor U21310 (N_21310,N_20670,N_20779);
and U21311 (N_21311,N_20965,N_20249);
or U21312 (N_21312,N_20070,N_20213);
xor U21313 (N_21313,N_20656,N_20303);
nor U21314 (N_21314,N_20229,N_20188);
or U21315 (N_21315,N_20185,N_20527);
or U21316 (N_21316,N_20799,N_20780);
xnor U21317 (N_21317,N_20015,N_20358);
or U21318 (N_21318,N_20043,N_20443);
nand U21319 (N_21319,N_20065,N_20028);
nor U21320 (N_21320,N_20054,N_20057);
nor U21321 (N_21321,N_20257,N_20519);
or U21322 (N_21322,N_20636,N_20587);
or U21323 (N_21323,N_20702,N_20629);
nand U21324 (N_21324,N_20761,N_20285);
and U21325 (N_21325,N_20549,N_20705);
xor U21326 (N_21326,N_20177,N_20048);
xnor U21327 (N_21327,N_20121,N_20014);
xor U21328 (N_21328,N_20926,N_20274);
xor U21329 (N_21329,N_20583,N_20886);
xor U21330 (N_21330,N_20322,N_20158);
and U21331 (N_21331,N_20365,N_20972);
nor U21332 (N_21332,N_20164,N_20565);
or U21333 (N_21333,N_20159,N_20191);
or U21334 (N_21334,N_20834,N_20954);
xor U21335 (N_21335,N_20226,N_20706);
and U21336 (N_21336,N_20523,N_20426);
xor U21337 (N_21337,N_20385,N_20463);
xor U21338 (N_21338,N_20261,N_20390);
xnor U21339 (N_21339,N_20442,N_20767);
or U21340 (N_21340,N_20948,N_20855);
nor U21341 (N_21341,N_20230,N_20914);
nand U21342 (N_21342,N_20988,N_20935);
nor U21343 (N_21343,N_20916,N_20682);
or U21344 (N_21344,N_20875,N_20215);
nor U21345 (N_21345,N_20562,N_20500);
nor U21346 (N_21346,N_20392,N_20713);
xnor U21347 (N_21347,N_20291,N_20862);
or U21348 (N_21348,N_20167,N_20072);
nand U21349 (N_21349,N_20698,N_20485);
xnor U21350 (N_21350,N_20712,N_20256);
nand U21351 (N_21351,N_20617,N_20396);
and U21352 (N_21352,N_20338,N_20080);
xnor U21353 (N_21353,N_20818,N_20962);
and U21354 (N_21354,N_20427,N_20644);
xnor U21355 (N_21355,N_20592,N_20880);
nand U21356 (N_21356,N_20734,N_20276);
nor U21357 (N_21357,N_20638,N_20173);
xor U21358 (N_21358,N_20003,N_20472);
xnor U21359 (N_21359,N_20842,N_20488);
xor U21360 (N_21360,N_20509,N_20138);
nand U21361 (N_21361,N_20608,N_20751);
xor U21362 (N_21362,N_20781,N_20380);
xnor U21363 (N_21363,N_20808,N_20894);
or U21364 (N_21364,N_20628,N_20324);
and U21365 (N_21365,N_20668,N_20924);
nand U21366 (N_21366,N_20323,N_20878);
or U21367 (N_21367,N_20217,N_20854);
or U21368 (N_21368,N_20021,N_20967);
nand U21369 (N_21369,N_20073,N_20006);
xnor U21370 (N_21370,N_20377,N_20258);
xnor U21371 (N_21371,N_20653,N_20115);
and U21372 (N_21372,N_20742,N_20822);
and U21373 (N_21373,N_20858,N_20662);
nand U21374 (N_21374,N_20602,N_20004);
or U21375 (N_21375,N_20664,N_20596);
and U21376 (N_21376,N_20784,N_20724);
nor U21377 (N_21377,N_20964,N_20354);
xnor U21378 (N_21378,N_20864,N_20031);
nor U21379 (N_21379,N_20910,N_20952);
and U21380 (N_21380,N_20945,N_20125);
nor U21381 (N_21381,N_20075,N_20446);
xnor U21382 (N_21382,N_20203,N_20002);
xor U21383 (N_21383,N_20183,N_20703);
or U21384 (N_21384,N_20599,N_20169);
and U21385 (N_21385,N_20084,N_20867);
nand U21386 (N_21386,N_20554,N_20297);
and U21387 (N_21387,N_20823,N_20264);
xor U21388 (N_21388,N_20503,N_20414);
xor U21389 (N_21389,N_20707,N_20813);
or U21390 (N_21390,N_20437,N_20413);
xnor U21391 (N_21391,N_20433,N_20714);
xor U21392 (N_21392,N_20553,N_20941);
nor U21393 (N_21393,N_20346,N_20311);
nand U21394 (N_21394,N_20849,N_20007);
or U21395 (N_21395,N_20921,N_20374);
and U21396 (N_21396,N_20735,N_20567);
or U21397 (N_21397,N_20260,N_20252);
nor U21398 (N_21398,N_20762,N_20652);
or U21399 (N_21399,N_20113,N_20546);
nor U21400 (N_21400,N_20709,N_20729);
xor U21401 (N_21401,N_20098,N_20774);
and U21402 (N_21402,N_20145,N_20833);
nand U21403 (N_21403,N_20319,N_20099);
or U21404 (N_21404,N_20786,N_20083);
xnor U21405 (N_21405,N_20364,N_20876);
nor U21406 (N_21406,N_20919,N_20210);
xnor U21407 (N_21407,N_20459,N_20464);
xnor U21408 (N_21408,N_20481,N_20694);
nor U21409 (N_21409,N_20928,N_20343);
nand U21410 (N_21410,N_20151,N_20239);
and U21411 (N_21411,N_20283,N_20708);
nand U21412 (N_21412,N_20310,N_20995);
or U21413 (N_21413,N_20467,N_20340);
and U21414 (N_21414,N_20050,N_20526);
nor U21415 (N_21415,N_20857,N_20633);
or U21416 (N_21416,N_20318,N_20548);
nand U21417 (N_21417,N_20570,N_20044);
and U21418 (N_21418,N_20493,N_20796);
nand U21419 (N_21419,N_20817,N_20425);
and U21420 (N_21420,N_20516,N_20209);
xor U21421 (N_21421,N_20897,N_20726);
nand U21422 (N_21422,N_20106,N_20793);
nand U21423 (N_21423,N_20157,N_20279);
nand U21424 (N_21424,N_20394,N_20750);
nand U21425 (N_21425,N_20270,N_20536);
or U21426 (N_21426,N_20267,N_20056);
or U21427 (N_21427,N_20946,N_20141);
and U21428 (N_21428,N_20899,N_20456);
nand U21429 (N_21429,N_20732,N_20087);
nand U21430 (N_21430,N_20951,N_20671);
nor U21431 (N_21431,N_20754,N_20327);
or U21432 (N_21432,N_20150,N_20174);
nand U21433 (N_21433,N_20920,N_20829);
nor U21434 (N_21434,N_20961,N_20298);
xnor U21435 (N_21435,N_20853,N_20838);
or U21436 (N_21436,N_20171,N_20741);
and U21437 (N_21437,N_20162,N_20040);
nor U21438 (N_21438,N_20429,N_20219);
xnor U21439 (N_21439,N_20074,N_20205);
nor U21440 (N_21440,N_20643,N_20462);
or U21441 (N_21441,N_20010,N_20773);
and U21442 (N_21442,N_20508,N_20913);
nor U21443 (N_21443,N_20593,N_20598);
nand U21444 (N_21444,N_20155,N_20556);
nand U21445 (N_21445,N_20905,N_20985);
nand U21446 (N_21446,N_20979,N_20679);
and U21447 (N_21447,N_20610,N_20045);
or U21448 (N_21448,N_20909,N_20747);
nand U21449 (N_21449,N_20225,N_20787);
and U21450 (N_21450,N_20116,N_20815);
or U21451 (N_21451,N_20969,N_20684);
xor U21452 (N_21452,N_20722,N_20247);
or U21453 (N_21453,N_20168,N_20482);
or U21454 (N_21454,N_20660,N_20621);
xnor U21455 (N_21455,N_20202,N_20521);
nor U21456 (N_21456,N_20518,N_20811);
and U21457 (N_21457,N_20542,N_20929);
nand U21458 (N_21458,N_20253,N_20033);
nand U21459 (N_21459,N_20304,N_20649);
nand U21460 (N_21460,N_20129,N_20581);
and U21461 (N_21461,N_20332,N_20971);
nand U21462 (N_21462,N_20309,N_20923);
xnor U21463 (N_21463,N_20362,N_20812);
or U21464 (N_21464,N_20206,N_20204);
nand U21465 (N_21465,N_20388,N_20027);
and U21466 (N_21466,N_20107,N_20255);
nand U21467 (N_21467,N_20282,N_20071);
or U21468 (N_21468,N_20353,N_20119);
nor U21469 (N_21469,N_20576,N_20420);
xor U21470 (N_21470,N_20584,N_20791);
or U21471 (N_21471,N_20637,N_20844);
nand U21472 (N_21472,N_20268,N_20657);
xor U21473 (N_21473,N_20254,N_20715);
nand U21474 (N_21474,N_20922,N_20746);
or U21475 (N_21475,N_20647,N_20888);
xnor U21476 (N_21476,N_20835,N_20982);
nand U21477 (N_21477,N_20411,N_20471);
or U21478 (N_21478,N_20294,N_20492);
nor U21479 (N_21479,N_20403,N_20540);
xnor U21480 (N_21480,N_20457,N_20194);
and U21481 (N_21481,N_20580,N_20907);
and U21482 (N_21482,N_20029,N_20695);
nand U21483 (N_21483,N_20410,N_20606);
nor U21484 (N_21484,N_20958,N_20758);
and U21485 (N_21485,N_20981,N_20114);
and U21486 (N_21486,N_20777,N_20063);
and U21487 (N_21487,N_20438,N_20005);
nand U21488 (N_21488,N_20555,N_20603);
nand U21489 (N_21489,N_20137,N_20983);
xor U21490 (N_21490,N_20052,N_20069);
nor U21491 (N_21491,N_20307,N_20055);
nor U21492 (N_21492,N_20563,N_20697);
xor U21493 (N_21493,N_20360,N_20661);
nand U21494 (N_21494,N_20047,N_20589);
nand U21495 (N_21495,N_20454,N_20363);
xor U21496 (N_21496,N_20575,N_20574);
or U21497 (N_21497,N_20127,N_20950);
or U21498 (N_21498,N_20564,N_20085);
and U21499 (N_21499,N_20240,N_20017);
nand U21500 (N_21500,N_20886,N_20629);
and U21501 (N_21501,N_20448,N_20043);
and U21502 (N_21502,N_20596,N_20635);
and U21503 (N_21503,N_20719,N_20963);
or U21504 (N_21504,N_20420,N_20642);
or U21505 (N_21505,N_20108,N_20155);
or U21506 (N_21506,N_20706,N_20514);
nand U21507 (N_21507,N_20004,N_20266);
nor U21508 (N_21508,N_20061,N_20342);
nand U21509 (N_21509,N_20101,N_20411);
xor U21510 (N_21510,N_20549,N_20230);
and U21511 (N_21511,N_20334,N_20911);
and U21512 (N_21512,N_20753,N_20981);
or U21513 (N_21513,N_20360,N_20396);
or U21514 (N_21514,N_20864,N_20413);
xnor U21515 (N_21515,N_20424,N_20103);
nand U21516 (N_21516,N_20254,N_20209);
nand U21517 (N_21517,N_20228,N_20875);
xnor U21518 (N_21518,N_20946,N_20942);
xor U21519 (N_21519,N_20490,N_20822);
xnor U21520 (N_21520,N_20268,N_20426);
xor U21521 (N_21521,N_20161,N_20728);
or U21522 (N_21522,N_20597,N_20840);
or U21523 (N_21523,N_20677,N_20720);
or U21524 (N_21524,N_20956,N_20201);
xor U21525 (N_21525,N_20235,N_20827);
xnor U21526 (N_21526,N_20922,N_20366);
nor U21527 (N_21527,N_20221,N_20048);
or U21528 (N_21528,N_20300,N_20684);
nor U21529 (N_21529,N_20178,N_20935);
xor U21530 (N_21530,N_20276,N_20335);
and U21531 (N_21531,N_20867,N_20620);
nor U21532 (N_21532,N_20203,N_20105);
nand U21533 (N_21533,N_20519,N_20100);
xnor U21534 (N_21534,N_20811,N_20977);
or U21535 (N_21535,N_20963,N_20796);
or U21536 (N_21536,N_20577,N_20077);
and U21537 (N_21537,N_20162,N_20269);
nand U21538 (N_21538,N_20742,N_20344);
nor U21539 (N_21539,N_20369,N_20489);
nand U21540 (N_21540,N_20248,N_20055);
and U21541 (N_21541,N_20102,N_20925);
nand U21542 (N_21542,N_20988,N_20567);
nand U21543 (N_21543,N_20156,N_20139);
xor U21544 (N_21544,N_20343,N_20669);
nor U21545 (N_21545,N_20927,N_20234);
or U21546 (N_21546,N_20196,N_20882);
nor U21547 (N_21547,N_20181,N_20664);
nor U21548 (N_21548,N_20639,N_20148);
and U21549 (N_21549,N_20594,N_20749);
nand U21550 (N_21550,N_20718,N_20899);
nor U21551 (N_21551,N_20055,N_20448);
nor U21552 (N_21552,N_20499,N_20216);
or U21553 (N_21553,N_20651,N_20644);
xor U21554 (N_21554,N_20376,N_20556);
nand U21555 (N_21555,N_20564,N_20838);
nor U21556 (N_21556,N_20713,N_20789);
or U21557 (N_21557,N_20048,N_20491);
nor U21558 (N_21558,N_20866,N_20684);
and U21559 (N_21559,N_20028,N_20315);
nand U21560 (N_21560,N_20389,N_20066);
or U21561 (N_21561,N_20686,N_20514);
xnor U21562 (N_21562,N_20016,N_20525);
nor U21563 (N_21563,N_20134,N_20099);
and U21564 (N_21564,N_20568,N_20377);
xor U21565 (N_21565,N_20016,N_20262);
nor U21566 (N_21566,N_20483,N_20941);
nor U21567 (N_21567,N_20888,N_20379);
nand U21568 (N_21568,N_20636,N_20852);
or U21569 (N_21569,N_20627,N_20155);
xnor U21570 (N_21570,N_20355,N_20559);
xor U21571 (N_21571,N_20260,N_20846);
xnor U21572 (N_21572,N_20209,N_20136);
or U21573 (N_21573,N_20764,N_20690);
or U21574 (N_21574,N_20950,N_20437);
nand U21575 (N_21575,N_20246,N_20518);
and U21576 (N_21576,N_20926,N_20355);
or U21577 (N_21577,N_20190,N_20478);
nor U21578 (N_21578,N_20701,N_20865);
nor U21579 (N_21579,N_20812,N_20683);
and U21580 (N_21580,N_20398,N_20469);
or U21581 (N_21581,N_20433,N_20718);
xor U21582 (N_21582,N_20681,N_20416);
nor U21583 (N_21583,N_20170,N_20385);
nor U21584 (N_21584,N_20891,N_20788);
or U21585 (N_21585,N_20344,N_20169);
and U21586 (N_21586,N_20598,N_20849);
nand U21587 (N_21587,N_20038,N_20773);
xnor U21588 (N_21588,N_20675,N_20351);
nor U21589 (N_21589,N_20477,N_20933);
or U21590 (N_21590,N_20730,N_20693);
and U21591 (N_21591,N_20635,N_20798);
nor U21592 (N_21592,N_20276,N_20000);
xnor U21593 (N_21593,N_20513,N_20416);
nor U21594 (N_21594,N_20188,N_20020);
or U21595 (N_21595,N_20471,N_20334);
nor U21596 (N_21596,N_20852,N_20662);
nor U21597 (N_21597,N_20704,N_20049);
nor U21598 (N_21598,N_20426,N_20630);
and U21599 (N_21599,N_20205,N_20258);
xnor U21600 (N_21600,N_20358,N_20334);
and U21601 (N_21601,N_20265,N_20388);
xnor U21602 (N_21602,N_20094,N_20512);
xor U21603 (N_21603,N_20024,N_20137);
nand U21604 (N_21604,N_20339,N_20197);
or U21605 (N_21605,N_20664,N_20654);
or U21606 (N_21606,N_20987,N_20849);
nand U21607 (N_21607,N_20114,N_20078);
xnor U21608 (N_21608,N_20093,N_20439);
nand U21609 (N_21609,N_20651,N_20413);
or U21610 (N_21610,N_20617,N_20297);
xnor U21611 (N_21611,N_20831,N_20010);
or U21612 (N_21612,N_20717,N_20550);
and U21613 (N_21613,N_20840,N_20617);
nor U21614 (N_21614,N_20425,N_20607);
and U21615 (N_21615,N_20012,N_20059);
and U21616 (N_21616,N_20451,N_20775);
or U21617 (N_21617,N_20257,N_20778);
nor U21618 (N_21618,N_20818,N_20629);
xnor U21619 (N_21619,N_20753,N_20762);
or U21620 (N_21620,N_20451,N_20798);
or U21621 (N_21621,N_20123,N_20044);
and U21622 (N_21622,N_20413,N_20306);
nor U21623 (N_21623,N_20104,N_20170);
xnor U21624 (N_21624,N_20191,N_20962);
xor U21625 (N_21625,N_20803,N_20336);
and U21626 (N_21626,N_20334,N_20929);
nor U21627 (N_21627,N_20000,N_20931);
or U21628 (N_21628,N_20961,N_20129);
nand U21629 (N_21629,N_20062,N_20680);
or U21630 (N_21630,N_20027,N_20562);
nand U21631 (N_21631,N_20442,N_20537);
nor U21632 (N_21632,N_20986,N_20888);
nor U21633 (N_21633,N_20719,N_20264);
xor U21634 (N_21634,N_20544,N_20839);
nand U21635 (N_21635,N_20403,N_20218);
or U21636 (N_21636,N_20173,N_20737);
nor U21637 (N_21637,N_20454,N_20339);
nand U21638 (N_21638,N_20008,N_20131);
nor U21639 (N_21639,N_20186,N_20760);
xor U21640 (N_21640,N_20364,N_20679);
xor U21641 (N_21641,N_20816,N_20594);
xnor U21642 (N_21642,N_20863,N_20896);
nor U21643 (N_21643,N_20183,N_20972);
and U21644 (N_21644,N_20101,N_20806);
and U21645 (N_21645,N_20074,N_20572);
xnor U21646 (N_21646,N_20519,N_20721);
nand U21647 (N_21647,N_20957,N_20516);
nand U21648 (N_21648,N_20652,N_20812);
xnor U21649 (N_21649,N_20198,N_20558);
and U21650 (N_21650,N_20165,N_20392);
xnor U21651 (N_21651,N_20505,N_20407);
nand U21652 (N_21652,N_20756,N_20543);
nor U21653 (N_21653,N_20703,N_20079);
and U21654 (N_21654,N_20733,N_20237);
or U21655 (N_21655,N_20220,N_20969);
nor U21656 (N_21656,N_20084,N_20254);
nor U21657 (N_21657,N_20240,N_20725);
nand U21658 (N_21658,N_20233,N_20890);
nor U21659 (N_21659,N_20038,N_20091);
or U21660 (N_21660,N_20826,N_20440);
nand U21661 (N_21661,N_20740,N_20199);
and U21662 (N_21662,N_20752,N_20831);
nor U21663 (N_21663,N_20113,N_20808);
and U21664 (N_21664,N_20994,N_20237);
or U21665 (N_21665,N_20927,N_20286);
or U21666 (N_21666,N_20776,N_20613);
nor U21667 (N_21667,N_20610,N_20994);
nand U21668 (N_21668,N_20697,N_20812);
and U21669 (N_21669,N_20470,N_20450);
nand U21670 (N_21670,N_20108,N_20984);
nand U21671 (N_21671,N_20910,N_20247);
xnor U21672 (N_21672,N_20836,N_20964);
nor U21673 (N_21673,N_20519,N_20838);
xor U21674 (N_21674,N_20275,N_20888);
and U21675 (N_21675,N_20592,N_20813);
xnor U21676 (N_21676,N_20534,N_20971);
or U21677 (N_21677,N_20395,N_20659);
and U21678 (N_21678,N_20306,N_20501);
or U21679 (N_21679,N_20282,N_20575);
or U21680 (N_21680,N_20800,N_20137);
or U21681 (N_21681,N_20548,N_20137);
or U21682 (N_21682,N_20643,N_20749);
or U21683 (N_21683,N_20347,N_20849);
and U21684 (N_21684,N_20367,N_20985);
or U21685 (N_21685,N_20122,N_20078);
nand U21686 (N_21686,N_20923,N_20357);
nand U21687 (N_21687,N_20863,N_20412);
and U21688 (N_21688,N_20664,N_20285);
nor U21689 (N_21689,N_20757,N_20077);
nor U21690 (N_21690,N_20666,N_20870);
xnor U21691 (N_21691,N_20093,N_20182);
and U21692 (N_21692,N_20469,N_20084);
or U21693 (N_21693,N_20703,N_20155);
xnor U21694 (N_21694,N_20352,N_20657);
xor U21695 (N_21695,N_20434,N_20981);
nand U21696 (N_21696,N_20775,N_20559);
nor U21697 (N_21697,N_20297,N_20728);
nor U21698 (N_21698,N_20850,N_20886);
and U21699 (N_21699,N_20854,N_20059);
nor U21700 (N_21700,N_20101,N_20543);
nor U21701 (N_21701,N_20260,N_20437);
xor U21702 (N_21702,N_20599,N_20397);
nor U21703 (N_21703,N_20950,N_20595);
nand U21704 (N_21704,N_20717,N_20517);
and U21705 (N_21705,N_20893,N_20117);
nand U21706 (N_21706,N_20040,N_20205);
nor U21707 (N_21707,N_20199,N_20842);
or U21708 (N_21708,N_20577,N_20522);
nand U21709 (N_21709,N_20880,N_20833);
or U21710 (N_21710,N_20629,N_20601);
and U21711 (N_21711,N_20386,N_20975);
xnor U21712 (N_21712,N_20016,N_20473);
nor U21713 (N_21713,N_20312,N_20466);
or U21714 (N_21714,N_20312,N_20793);
or U21715 (N_21715,N_20698,N_20734);
nand U21716 (N_21716,N_20570,N_20941);
xnor U21717 (N_21717,N_20373,N_20042);
and U21718 (N_21718,N_20073,N_20485);
xor U21719 (N_21719,N_20164,N_20634);
and U21720 (N_21720,N_20578,N_20567);
nor U21721 (N_21721,N_20112,N_20367);
and U21722 (N_21722,N_20921,N_20351);
or U21723 (N_21723,N_20812,N_20417);
or U21724 (N_21724,N_20261,N_20196);
nor U21725 (N_21725,N_20405,N_20778);
or U21726 (N_21726,N_20095,N_20870);
nand U21727 (N_21727,N_20048,N_20676);
and U21728 (N_21728,N_20732,N_20270);
xnor U21729 (N_21729,N_20746,N_20182);
nand U21730 (N_21730,N_20542,N_20732);
and U21731 (N_21731,N_20934,N_20507);
and U21732 (N_21732,N_20304,N_20283);
nand U21733 (N_21733,N_20012,N_20202);
xnor U21734 (N_21734,N_20665,N_20960);
xor U21735 (N_21735,N_20285,N_20269);
xor U21736 (N_21736,N_20928,N_20885);
nor U21737 (N_21737,N_20101,N_20634);
xnor U21738 (N_21738,N_20796,N_20103);
xnor U21739 (N_21739,N_20167,N_20439);
nor U21740 (N_21740,N_20721,N_20972);
xor U21741 (N_21741,N_20805,N_20987);
nor U21742 (N_21742,N_20909,N_20011);
nand U21743 (N_21743,N_20348,N_20369);
and U21744 (N_21744,N_20264,N_20403);
xor U21745 (N_21745,N_20703,N_20064);
or U21746 (N_21746,N_20106,N_20297);
and U21747 (N_21747,N_20020,N_20755);
and U21748 (N_21748,N_20776,N_20725);
nor U21749 (N_21749,N_20864,N_20960);
and U21750 (N_21750,N_20317,N_20009);
nand U21751 (N_21751,N_20877,N_20703);
or U21752 (N_21752,N_20411,N_20916);
xor U21753 (N_21753,N_20225,N_20721);
and U21754 (N_21754,N_20031,N_20119);
nand U21755 (N_21755,N_20191,N_20843);
nand U21756 (N_21756,N_20978,N_20354);
xor U21757 (N_21757,N_20035,N_20292);
and U21758 (N_21758,N_20461,N_20697);
nand U21759 (N_21759,N_20708,N_20248);
nand U21760 (N_21760,N_20316,N_20543);
or U21761 (N_21761,N_20391,N_20106);
or U21762 (N_21762,N_20735,N_20667);
and U21763 (N_21763,N_20968,N_20177);
nand U21764 (N_21764,N_20314,N_20679);
nor U21765 (N_21765,N_20351,N_20051);
and U21766 (N_21766,N_20439,N_20917);
nor U21767 (N_21767,N_20472,N_20584);
nand U21768 (N_21768,N_20819,N_20383);
xnor U21769 (N_21769,N_20720,N_20464);
xor U21770 (N_21770,N_20315,N_20487);
xor U21771 (N_21771,N_20548,N_20488);
or U21772 (N_21772,N_20526,N_20809);
nor U21773 (N_21773,N_20489,N_20902);
nand U21774 (N_21774,N_20162,N_20937);
nor U21775 (N_21775,N_20742,N_20435);
and U21776 (N_21776,N_20069,N_20648);
nand U21777 (N_21777,N_20346,N_20923);
or U21778 (N_21778,N_20899,N_20964);
nand U21779 (N_21779,N_20466,N_20944);
xnor U21780 (N_21780,N_20171,N_20864);
and U21781 (N_21781,N_20374,N_20847);
or U21782 (N_21782,N_20560,N_20964);
nand U21783 (N_21783,N_20801,N_20472);
or U21784 (N_21784,N_20225,N_20181);
and U21785 (N_21785,N_20884,N_20791);
or U21786 (N_21786,N_20856,N_20100);
xnor U21787 (N_21787,N_20863,N_20928);
or U21788 (N_21788,N_20581,N_20949);
xor U21789 (N_21789,N_20194,N_20901);
nor U21790 (N_21790,N_20254,N_20464);
xor U21791 (N_21791,N_20397,N_20566);
nor U21792 (N_21792,N_20878,N_20987);
nand U21793 (N_21793,N_20364,N_20142);
nor U21794 (N_21794,N_20043,N_20886);
xnor U21795 (N_21795,N_20479,N_20086);
or U21796 (N_21796,N_20299,N_20258);
nand U21797 (N_21797,N_20816,N_20906);
nor U21798 (N_21798,N_20057,N_20134);
nor U21799 (N_21799,N_20757,N_20727);
nor U21800 (N_21800,N_20000,N_20351);
and U21801 (N_21801,N_20143,N_20970);
nor U21802 (N_21802,N_20542,N_20113);
nand U21803 (N_21803,N_20551,N_20486);
and U21804 (N_21804,N_20635,N_20548);
xnor U21805 (N_21805,N_20472,N_20548);
nor U21806 (N_21806,N_20451,N_20640);
nand U21807 (N_21807,N_20189,N_20453);
nand U21808 (N_21808,N_20673,N_20087);
and U21809 (N_21809,N_20539,N_20064);
nor U21810 (N_21810,N_20528,N_20101);
nor U21811 (N_21811,N_20552,N_20134);
nand U21812 (N_21812,N_20850,N_20622);
nand U21813 (N_21813,N_20020,N_20741);
or U21814 (N_21814,N_20124,N_20796);
nor U21815 (N_21815,N_20281,N_20944);
and U21816 (N_21816,N_20573,N_20528);
nor U21817 (N_21817,N_20556,N_20634);
or U21818 (N_21818,N_20862,N_20000);
nand U21819 (N_21819,N_20072,N_20547);
xnor U21820 (N_21820,N_20100,N_20670);
or U21821 (N_21821,N_20174,N_20226);
nor U21822 (N_21822,N_20646,N_20660);
nand U21823 (N_21823,N_20482,N_20933);
xnor U21824 (N_21824,N_20524,N_20693);
nor U21825 (N_21825,N_20863,N_20659);
or U21826 (N_21826,N_20494,N_20844);
xor U21827 (N_21827,N_20108,N_20934);
nor U21828 (N_21828,N_20635,N_20845);
xor U21829 (N_21829,N_20219,N_20517);
xnor U21830 (N_21830,N_20390,N_20666);
and U21831 (N_21831,N_20170,N_20293);
nand U21832 (N_21832,N_20285,N_20092);
xnor U21833 (N_21833,N_20210,N_20334);
or U21834 (N_21834,N_20580,N_20115);
or U21835 (N_21835,N_20785,N_20125);
xnor U21836 (N_21836,N_20196,N_20569);
xor U21837 (N_21837,N_20622,N_20586);
and U21838 (N_21838,N_20392,N_20374);
xor U21839 (N_21839,N_20168,N_20723);
nor U21840 (N_21840,N_20732,N_20302);
xnor U21841 (N_21841,N_20776,N_20929);
xnor U21842 (N_21842,N_20298,N_20646);
nand U21843 (N_21843,N_20313,N_20450);
and U21844 (N_21844,N_20316,N_20527);
xnor U21845 (N_21845,N_20495,N_20090);
xnor U21846 (N_21846,N_20673,N_20717);
or U21847 (N_21847,N_20474,N_20348);
nor U21848 (N_21848,N_20908,N_20790);
or U21849 (N_21849,N_20568,N_20832);
or U21850 (N_21850,N_20396,N_20145);
xnor U21851 (N_21851,N_20643,N_20690);
nor U21852 (N_21852,N_20104,N_20052);
nor U21853 (N_21853,N_20518,N_20161);
xor U21854 (N_21854,N_20531,N_20921);
nand U21855 (N_21855,N_20137,N_20349);
or U21856 (N_21856,N_20309,N_20540);
nand U21857 (N_21857,N_20009,N_20087);
or U21858 (N_21858,N_20317,N_20094);
nor U21859 (N_21859,N_20281,N_20929);
xor U21860 (N_21860,N_20864,N_20153);
nor U21861 (N_21861,N_20830,N_20511);
nand U21862 (N_21862,N_20866,N_20195);
and U21863 (N_21863,N_20735,N_20271);
nand U21864 (N_21864,N_20679,N_20546);
xnor U21865 (N_21865,N_20621,N_20229);
nor U21866 (N_21866,N_20508,N_20739);
xnor U21867 (N_21867,N_20833,N_20762);
nor U21868 (N_21868,N_20085,N_20463);
xnor U21869 (N_21869,N_20815,N_20240);
xor U21870 (N_21870,N_20577,N_20894);
xnor U21871 (N_21871,N_20867,N_20534);
or U21872 (N_21872,N_20216,N_20326);
and U21873 (N_21873,N_20383,N_20107);
nand U21874 (N_21874,N_20346,N_20455);
or U21875 (N_21875,N_20261,N_20732);
nor U21876 (N_21876,N_20698,N_20765);
nand U21877 (N_21877,N_20240,N_20878);
and U21878 (N_21878,N_20042,N_20747);
or U21879 (N_21879,N_20023,N_20667);
xor U21880 (N_21880,N_20529,N_20535);
xnor U21881 (N_21881,N_20402,N_20285);
xnor U21882 (N_21882,N_20808,N_20622);
nand U21883 (N_21883,N_20928,N_20241);
nor U21884 (N_21884,N_20573,N_20139);
nand U21885 (N_21885,N_20594,N_20807);
or U21886 (N_21886,N_20123,N_20749);
nor U21887 (N_21887,N_20792,N_20368);
nand U21888 (N_21888,N_20091,N_20269);
and U21889 (N_21889,N_20578,N_20278);
xor U21890 (N_21890,N_20924,N_20994);
nand U21891 (N_21891,N_20091,N_20608);
or U21892 (N_21892,N_20969,N_20677);
and U21893 (N_21893,N_20588,N_20445);
or U21894 (N_21894,N_20056,N_20394);
nand U21895 (N_21895,N_20555,N_20284);
and U21896 (N_21896,N_20982,N_20829);
nor U21897 (N_21897,N_20092,N_20508);
nand U21898 (N_21898,N_20827,N_20618);
or U21899 (N_21899,N_20151,N_20320);
nor U21900 (N_21900,N_20389,N_20744);
nor U21901 (N_21901,N_20383,N_20245);
and U21902 (N_21902,N_20120,N_20036);
xor U21903 (N_21903,N_20169,N_20929);
nand U21904 (N_21904,N_20627,N_20575);
xor U21905 (N_21905,N_20699,N_20192);
or U21906 (N_21906,N_20085,N_20483);
or U21907 (N_21907,N_20771,N_20357);
or U21908 (N_21908,N_20480,N_20667);
or U21909 (N_21909,N_20999,N_20971);
or U21910 (N_21910,N_20682,N_20933);
or U21911 (N_21911,N_20202,N_20871);
nor U21912 (N_21912,N_20985,N_20638);
xnor U21913 (N_21913,N_20587,N_20605);
or U21914 (N_21914,N_20017,N_20275);
xnor U21915 (N_21915,N_20405,N_20481);
and U21916 (N_21916,N_20346,N_20282);
or U21917 (N_21917,N_20416,N_20626);
nor U21918 (N_21918,N_20172,N_20591);
nor U21919 (N_21919,N_20755,N_20848);
nor U21920 (N_21920,N_20487,N_20375);
or U21921 (N_21921,N_20794,N_20539);
or U21922 (N_21922,N_20242,N_20468);
xor U21923 (N_21923,N_20760,N_20157);
nor U21924 (N_21924,N_20048,N_20449);
or U21925 (N_21925,N_20274,N_20749);
or U21926 (N_21926,N_20848,N_20503);
and U21927 (N_21927,N_20020,N_20903);
and U21928 (N_21928,N_20305,N_20138);
and U21929 (N_21929,N_20901,N_20379);
xnor U21930 (N_21930,N_20270,N_20208);
and U21931 (N_21931,N_20031,N_20255);
and U21932 (N_21932,N_20614,N_20597);
or U21933 (N_21933,N_20898,N_20411);
xor U21934 (N_21934,N_20579,N_20177);
xor U21935 (N_21935,N_20174,N_20378);
or U21936 (N_21936,N_20102,N_20383);
xor U21937 (N_21937,N_20588,N_20776);
and U21938 (N_21938,N_20080,N_20262);
and U21939 (N_21939,N_20143,N_20048);
or U21940 (N_21940,N_20269,N_20831);
nor U21941 (N_21941,N_20140,N_20078);
or U21942 (N_21942,N_20874,N_20490);
or U21943 (N_21943,N_20234,N_20802);
nand U21944 (N_21944,N_20537,N_20735);
nand U21945 (N_21945,N_20413,N_20462);
or U21946 (N_21946,N_20735,N_20722);
and U21947 (N_21947,N_20490,N_20946);
or U21948 (N_21948,N_20025,N_20099);
nor U21949 (N_21949,N_20337,N_20545);
or U21950 (N_21950,N_20287,N_20392);
nand U21951 (N_21951,N_20036,N_20301);
nand U21952 (N_21952,N_20567,N_20112);
xor U21953 (N_21953,N_20037,N_20845);
xnor U21954 (N_21954,N_20664,N_20712);
nor U21955 (N_21955,N_20668,N_20652);
xnor U21956 (N_21956,N_20163,N_20224);
xnor U21957 (N_21957,N_20010,N_20176);
and U21958 (N_21958,N_20803,N_20448);
and U21959 (N_21959,N_20729,N_20477);
nand U21960 (N_21960,N_20164,N_20439);
nor U21961 (N_21961,N_20699,N_20432);
nor U21962 (N_21962,N_20728,N_20524);
xor U21963 (N_21963,N_20452,N_20501);
or U21964 (N_21964,N_20048,N_20129);
or U21965 (N_21965,N_20849,N_20943);
or U21966 (N_21966,N_20123,N_20220);
nand U21967 (N_21967,N_20039,N_20701);
or U21968 (N_21968,N_20035,N_20436);
nand U21969 (N_21969,N_20580,N_20940);
and U21970 (N_21970,N_20112,N_20141);
xor U21971 (N_21971,N_20105,N_20361);
nor U21972 (N_21972,N_20030,N_20398);
nor U21973 (N_21973,N_20727,N_20111);
xor U21974 (N_21974,N_20340,N_20786);
xor U21975 (N_21975,N_20895,N_20708);
nand U21976 (N_21976,N_20093,N_20927);
nand U21977 (N_21977,N_20636,N_20786);
nor U21978 (N_21978,N_20640,N_20218);
and U21979 (N_21979,N_20058,N_20040);
xor U21980 (N_21980,N_20290,N_20369);
nand U21981 (N_21981,N_20532,N_20174);
and U21982 (N_21982,N_20895,N_20296);
xnor U21983 (N_21983,N_20757,N_20270);
or U21984 (N_21984,N_20896,N_20606);
xnor U21985 (N_21985,N_20103,N_20143);
and U21986 (N_21986,N_20928,N_20359);
and U21987 (N_21987,N_20024,N_20327);
xor U21988 (N_21988,N_20497,N_20191);
nor U21989 (N_21989,N_20969,N_20085);
and U21990 (N_21990,N_20795,N_20706);
and U21991 (N_21991,N_20841,N_20014);
and U21992 (N_21992,N_20069,N_20057);
xnor U21993 (N_21993,N_20362,N_20990);
and U21994 (N_21994,N_20040,N_20122);
and U21995 (N_21995,N_20707,N_20491);
xor U21996 (N_21996,N_20109,N_20864);
xnor U21997 (N_21997,N_20730,N_20688);
and U21998 (N_21998,N_20177,N_20898);
and U21999 (N_21999,N_20741,N_20688);
nor U22000 (N_22000,N_21384,N_21208);
or U22001 (N_22001,N_21137,N_21115);
and U22002 (N_22002,N_21278,N_21023);
nor U22003 (N_22003,N_21445,N_21908);
and U22004 (N_22004,N_21341,N_21449);
or U22005 (N_22005,N_21574,N_21436);
and U22006 (N_22006,N_21031,N_21952);
nor U22007 (N_22007,N_21662,N_21894);
or U22008 (N_22008,N_21372,N_21757);
nand U22009 (N_22009,N_21466,N_21728);
xor U22010 (N_22010,N_21541,N_21104);
xor U22011 (N_22011,N_21802,N_21509);
or U22012 (N_22012,N_21551,N_21114);
xnor U22013 (N_22013,N_21712,N_21156);
xor U22014 (N_22014,N_21258,N_21090);
xnor U22015 (N_22015,N_21781,N_21929);
and U22016 (N_22016,N_21299,N_21048);
and U22017 (N_22017,N_21798,N_21423);
xor U22018 (N_22018,N_21378,N_21331);
and U22019 (N_22019,N_21027,N_21112);
nand U22020 (N_22020,N_21742,N_21022);
and U22021 (N_22021,N_21769,N_21035);
and U22022 (N_22022,N_21191,N_21374);
xnor U22023 (N_22023,N_21032,N_21223);
nand U22024 (N_22024,N_21109,N_21864);
or U22025 (N_22025,N_21256,N_21825);
and U22026 (N_22026,N_21653,N_21316);
or U22027 (N_22027,N_21996,N_21873);
or U22028 (N_22028,N_21155,N_21025);
or U22029 (N_22029,N_21094,N_21508);
or U22030 (N_22030,N_21797,N_21555);
and U22031 (N_22031,N_21790,N_21598);
nor U22032 (N_22032,N_21001,N_21393);
xnor U22033 (N_22033,N_21514,N_21334);
nand U22034 (N_22034,N_21865,N_21992);
or U22035 (N_22035,N_21298,N_21260);
or U22036 (N_22036,N_21990,N_21755);
nor U22037 (N_22037,N_21167,N_21146);
nor U22038 (N_22038,N_21454,N_21077);
and U22039 (N_22039,N_21792,N_21743);
nand U22040 (N_22040,N_21589,N_21178);
or U22041 (N_22041,N_21909,N_21314);
and U22042 (N_22042,N_21738,N_21666);
and U22043 (N_22043,N_21373,N_21296);
or U22044 (N_22044,N_21088,N_21093);
or U22045 (N_22045,N_21692,N_21435);
xor U22046 (N_22046,N_21877,N_21029);
xnor U22047 (N_22047,N_21713,N_21214);
xor U22048 (N_22048,N_21487,N_21740);
or U22049 (N_22049,N_21481,N_21659);
nor U22050 (N_22050,N_21690,N_21678);
and U22051 (N_22051,N_21236,N_21564);
nand U22052 (N_22052,N_21193,N_21335);
or U22053 (N_22053,N_21931,N_21768);
or U22054 (N_22054,N_21679,N_21421);
or U22055 (N_22055,N_21889,N_21732);
and U22056 (N_22056,N_21087,N_21203);
nand U22057 (N_22057,N_21917,N_21745);
nor U22058 (N_22058,N_21180,N_21938);
nor U22059 (N_22059,N_21513,N_21493);
xor U22060 (N_22060,N_21106,N_21630);
nor U22061 (N_22061,N_21361,N_21741);
nand U22062 (N_22062,N_21015,N_21351);
nand U22063 (N_22063,N_21476,N_21561);
nand U22064 (N_22064,N_21726,N_21762);
nand U22065 (N_22065,N_21394,N_21615);
xnor U22066 (N_22066,N_21703,N_21302);
xnor U22067 (N_22067,N_21154,N_21309);
and U22068 (N_22068,N_21707,N_21885);
or U22069 (N_22069,N_21338,N_21357);
or U22070 (N_22070,N_21629,N_21469);
nand U22071 (N_22071,N_21535,N_21572);
nor U22072 (N_22072,N_21641,N_21091);
nor U22073 (N_22073,N_21567,N_21892);
or U22074 (N_22074,N_21654,N_21720);
nor U22075 (N_22075,N_21969,N_21324);
or U22076 (N_22076,N_21689,N_21585);
or U22077 (N_22077,N_21233,N_21044);
or U22078 (N_22078,N_21642,N_21100);
nor U22079 (N_22079,N_21113,N_21472);
xnor U22080 (N_22080,N_21839,N_21490);
nand U22081 (N_22081,N_21295,N_21447);
or U22082 (N_22082,N_21080,N_21446);
nand U22083 (N_22083,N_21681,N_21353);
nand U22084 (N_22084,N_21166,N_21565);
xnor U22085 (N_22085,N_21544,N_21566);
nand U22086 (N_22086,N_21796,N_21748);
and U22087 (N_22087,N_21016,N_21013);
nand U22088 (N_22088,N_21517,N_21063);
nor U22089 (N_22089,N_21542,N_21949);
nand U22090 (N_22090,N_21479,N_21608);
or U22091 (N_22091,N_21684,N_21340);
nand U22092 (N_22092,N_21052,N_21614);
nor U22093 (N_22093,N_21528,N_21623);
and U22094 (N_22094,N_21227,N_21941);
and U22095 (N_22095,N_21511,N_21122);
and U22096 (N_22096,N_21283,N_21304);
xor U22097 (N_22097,N_21640,N_21079);
xor U22098 (N_22098,N_21587,N_21257);
nor U22099 (N_22099,N_21102,N_21682);
nand U22100 (N_22100,N_21414,N_21054);
xnor U22101 (N_22101,N_21377,N_21005);
and U22102 (N_22102,N_21842,N_21368);
nor U22103 (N_22103,N_21664,N_21516);
or U22104 (N_22104,N_21096,N_21006);
nand U22105 (N_22105,N_21793,N_21636);
nand U22106 (N_22106,N_21422,N_21847);
xor U22107 (N_22107,N_21600,N_21785);
and U22108 (N_22108,N_21669,N_21158);
xor U22109 (N_22109,N_21495,N_21882);
nand U22110 (N_22110,N_21134,N_21880);
or U22111 (N_22111,N_21285,N_21951);
or U22112 (N_22112,N_21021,N_21019);
and U22113 (N_22113,N_21083,N_21136);
or U22114 (N_22114,N_21263,N_21914);
and U22115 (N_22115,N_21431,N_21474);
xor U22116 (N_22116,N_21795,N_21000);
or U22117 (N_22117,N_21721,N_21905);
or U22118 (N_22118,N_21903,N_21550);
or U22119 (N_22119,N_21596,N_21456);
nor U22120 (N_22120,N_21074,N_21637);
or U22121 (N_22121,N_21303,N_21014);
nor U22122 (N_22122,N_21343,N_21638);
nor U22123 (N_22123,N_21458,N_21558);
nand U22124 (N_22124,N_21226,N_21066);
xnor U22125 (N_22125,N_21310,N_21046);
and U22126 (N_22126,N_21519,N_21869);
or U22127 (N_22127,N_21776,N_21126);
and U22128 (N_22128,N_21186,N_21264);
or U22129 (N_22129,N_21665,N_21881);
or U22130 (N_22130,N_21277,N_21563);
nand U22131 (N_22131,N_21876,N_21715);
xnor U22132 (N_22132,N_21747,N_21663);
and U22133 (N_22133,N_21603,N_21627);
nand U22134 (N_22134,N_21979,N_21269);
nand U22135 (N_22135,N_21228,N_21694);
xor U22136 (N_22136,N_21968,N_21185);
and U22137 (N_22137,N_21230,N_21024);
and U22138 (N_22138,N_21028,N_21286);
nand U22139 (N_22139,N_21232,N_21358);
nand U22140 (N_22140,N_21330,N_21098);
or U22141 (N_22141,N_21696,N_21271);
xnor U22142 (N_22142,N_21430,N_21287);
or U22143 (N_22143,N_21680,N_21658);
nor U22144 (N_22144,N_21462,N_21464);
nor U22145 (N_22145,N_21457,N_21062);
nand U22146 (N_22146,N_21848,N_21778);
nand U22147 (N_22147,N_21925,N_21655);
nor U22148 (N_22148,N_21497,N_21554);
and U22149 (N_22149,N_21701,N_21010);
nor U22150 (N_22150,N_21860,N_21577);
and U22151 (N_22151,N_21266,N_21238);
and U22152 (N_22152,N_21834,N_21009);
xor U22153 (N_22153,N_21200,N_21926);
xnor U22154 (N_22154,N_21526,N_21759);
and U22155 (N_22155,N_21501,N_21532);
and U22156 (N_22156,N_21400,N_21862);
nor U22157 (N_22157,N_21904,N_21279);
or U22158 (N_22158,N_21007,N_21211);
and U22159 (N_22159,N_21950,N_21116);
nor U22160 (N_22160,N_21945,N_21103);
and U22161 (N_22161,N_21890,N_21254);
or U22162 (N_22162,N_21901,N_21717);
or U22163 (N_22163,N_21282,N_21492);
and U22164 (N_22164,N_21518,N_21830);
nor U22165 (N_22165,N_21716,N_21977);
nand U22166 (N_22166,N_21646,N_21718);
and U22167 (N_22167,N_21455,N_21329);
and U22168 (N_22168,N_21843,N_21504);
nand U22169 (N_22169,N_21594,N_21360);
nor U22170 (N_22170,N_21484,N_21383);
or U22171 (N_22171,N_21042,N_21245);
xnor U22172 (N_22172,N_21810,N_21922);
nor U22173 (N_22173,N_21705,N_21183);
xor U22174 (N_22174,N_21837,N_21610);
xnor U22175 (N_22175,N_21012,N_21473);
or U22176 (N_22176,N_21121,N_21893);
xnor U22177 (N_22177,N_21159,N_21828);
nor U22178 (N_22178,N_21710,N_21783);
and U22179 (N_22179,N_21936,N_21099);
or U22180 (N_22180,N_21339,N_21132);
xor U22181 (N_22181,N_21592,N_21319);
and U22182 (N_22182,N_21415,N_21039);
xor U22183 (N_22183,N_21127,N_21240);
xor U22184 (N_22184,N_21349,N_21390);
xor U22185 (N_22185,N_21043,N_21078);
and U22186 (N_22186,N_21853,N_21426);
xor U22187 (N_22187,N_21725,N_21050);
and U22188 (N_22188,N_21290,N_21300);
xnor U22189 (N_22189,N_21625,N_21736);
nor U22190 (N_22190,N_21459,N_21347);
or U22191 (N_22191,N_21405,N_21182);
or U22192 (N_22192,N_21082,N_21863);
nand U22193 (N_22193,N_21534,N_21986);
nand U22194 (N_22194,N_21386,N_21907);
and U22195 (N_22195,N_21261,N_21190);
nand U22196 (N_22196,N_21766,N_21852);
xor U22197 (N_22197,N_21691,N_21808);
or U22198 (N_22198,N_21089,N_21174);
or U22199 (N_22199,N_21123,N_21581);
and U22200 (N_22200,N_21411,N_21311);
nor U22201 (N_22201,N_21760,N_21620);
or U22202 (N_22202,N_21997,N_21225);
xnor U22203 (N_22203,N_21605,N_21499);
and U22204 (N_22204,N_21609,N_21879);
and U22205 (N_22205,N_21651,N_21438);
and U22206 (N_22206,N_21375,N_21246);
or U22207 (N_22207,N_21677,N_21588);
or U22208 (N_22208,N_21294,N_21595);
nor U22209 (N_22209,N_21590,N_21234);
nor U22210 (N_22210,N_21205,N_21161);
nor U22211 (N_22211,N_21305,N_21222);
nor U22212 (N_22212,N_21409,N_21382);
nor U22213 (N_22213,N_21398,N_21546);
and U22214 (N_22214,N_21788,N_21172);
xor U22215 (N_22215,N_21560,N_21686);
xnor U22216 (N_22216,N_21189,N_21056);
or U22217 (N_22217,N_21631,N_21058);
or U22218 (N_22218,N_21955,N_21536);
xnor U22219 (N_22219,N_21924,N_21671);
nand U22220 (N_22220,N_21841,N_21367);
or U22221 (N_22221,N_21317,N_21521);
xnor U22222 (N_22222,N_21051,N_21346);
or U22223 (N_22223,N_21259,N_21756);
or U22224 (N_22224,N_21318,N_21380);
xor U22225 (N_22225,N_21417,N_21477);
xnor U22226 (N_22226,N_21896,N_21751);
or U22227 (N_22227,N_21849,N_21195);
xor U22228 (N_22228,N_21060,N_21003);
or U22229 (N_22229,N_21342,N_21424);
xor U22230 (N_22230,N_21645,N_21273);
nor U22231 (N_22231,N_21582,N_21068);
xnor U22232 (N_22232,N_21453,N_21500);
xnor U22233 (N_22233,N_21209,N_21819);
nand U22234 (N_22234,N_21761,N_21537);
and U22235 (N_22235,N_21915,N_21789);
xor U22236 (N_22236,N_21130,N_21359);
nand U22237 (N_22237,N_21972,N_21601);
nor U22238 (N_22238,N_21510,N_21800);
xor U22239 (N_22239,N_21957,N_21505);
and U22240 (N_22240,N_21970,N_21391);
nor U22241 (N_22241,N_21782,N_21765);
nor U22242 (N_22242,N_21463,N_21838);
nand U22243 (N_22243,N_21612,N_21496);
nand U22244 (N_22244,N_21727,N_21084);
nand U22245 (N_22245,N_21478,N_21235);
nor U22246 (N_22246,N_21752,N_21937);
nand U22247 (N_22247,N_21061,N_21268);
nand U22248 (N_22248,N_21771,N_21072);
or U22249 (N_22249,N_21606,N_21965);
nand U22250 (N_22250,N_21583,N_21026);
nor U22251 (N_22251,N_21212,N_21939);
xor U22252 (N_22252,N_21219,N_21198);
nor U22253 (N_22253,N_21962,N_21385);
and U22254 (N_22254,N_21213,N_21471);
xnor U22255 (N_22255,N_21777,N_21580);
xor U22256 (N_22256,N_21856,N_21451);
xnor U22257 (N_22257,N_21954,N_21075);
nor U22258 (N_22258,N_21498,N_21163);
nor U22259 (N_22259,N_21365,N_21370);
xor U22260 (N_22260,N_21932,N_21900);
nor U22261 (N_22261,N_21364,N_21241);
xnor U22262 (N_22262,N_21170,N_21111);
or U22263 (N_22263,N_21779,N_21323);
and U22264 (N_22264,N_21832,N_21253);
or U22265 (N_22265,N_21911,N_21450);
and U22266 (N_22266,N_21943,N_21814);
or U22267 (N_22267,N_21753,N_21724);
and U22268 (N_22268,N_21059,N_21995);
nand U22269 (N_22269,N_21468,N_21321);
nand U22270 (N_22270,N_21959,N_21433);
or U22271 (N_22271,N_21619,N_21821);
nand U22272 (N_22272,N_21557,N_21419);
and U22273 (N_22273,N_21846,N_21650);
nand U22274 (N_22274,N_21540,N_21131);
or U22275 (N_22275,N_21206,N_21735);
or U22276 (N_22276,N_21181,N_21151);
nor U22277 (N_22277,N_21201,N_21772);
or U22278 (N_22278,N_21418,N_21221);
and U22279 (N_22279,N_21723,N_21153);
nand U22280 (N_22280,N_21045,N_21661);
or U22281 (N_22281,N_21095,N_21416);
xnor U22282 (N_22282,N_21617,N_21412);
nor U22283 (N_22283,N_21387,N_21754);
xnor U22284 (N_22284,N_21845,N_21086);
and U22285 (N_22285,N_21921,N_21399);
nor U22286 (N_22286,N_21371,N_21998);
nor U22287 (N_22287,N_21410,N_21744);
xnor U22288 (N_22288,N_21624,N_21437);
nand U22289 (N_22289,N_21429,N_21401);
or U22290 (N_22290,N_21488,N_21980);
and U22291 (N_22291,N_21611,N_21327);
xnor U22292 (N_22292,N_21442,N_21971);
nand U22293 (N_22293,N_21657,N_21482);
xnor U22294 (N_22294,N_21250,N_21584);
or U22295 (N_22295,N_21171,N_21483);
or U22296 (N_22296,N_21345,N_21815);
nand U22297 (N_22297,N_21571,N_21942);
or U22298 (N_22298,N_21008,N_21218);
xor U22299 (N_22299,N_21337,N_21820);
and U22300 (N_22300,N_21780,N_21770);
nand U22301 (N_22301,N_21613,N_21593);
or U22302 (N_22302,N_21556,N_21529);
and U22303 (N_22303,N_21674,N_21823);
or U22304 (N_22304,N_21229,N_21366);
or U22305 (N_22305,N_21933,N_21799);
nor U22306 (N_22306,N_21276,N_21160);
and U22307 (N_22307,N_21953,N_21425);
or U22308 (N_22308,N_21210,N_21520);
or U22309 (N_22309,N_21672,N_21836);
nor U22310 (N_22310,N_21961,N_21981);
and U22311 (N_22311,N_21784,N_21177);
xnor U22312 (N_22312,N_21656,N_21649);
or U22313 (N_22313,N_21530,N_21135);
and U22314 (N_22314,N_21702,N_21396);
or U22315 (N_22315,N_21874,N_21002);
xnor U22316 (N_22316,N_21251,N_21987);
and U22317 (N_22317,N_21685,N_21774);
nor U22318 (N_22318,N_21543,N_21963);
and U22319 (N_22319,N_21117,N_21733);
nand U22320 (N_22320,N_21315,N_21176);
nor U22321 (N_22321,N_21737,N_21306);
xor U22322 (N_22322,N_21773,N_21144);
xnor U22323 (N_22323,N_21982,N_21729);
or U22324 (N_22324,N_21055,N_21242);
and U22325 (N_22325,N_21199,N_21579);
nand U22326 (N_22326,N_21110,N_21714);
and U22327 (N_22327,N_21291,N_21886);
or U22328 (N_22328,N_21363,N_21887);
nor U22329 (N_22329,N_21439,N_21859);
nand U22330 (N_22330,N_21602,N_21767);
xnor U22331 (N_22331,N_21325,N_21244);
xnor U22332 (N_22332,N_21197,N_21017);
or U22333 (N_22333,N_21355,N_21041);
xor U22334 (N_22334,N_21960,N_21280);
or U22335 (N_22335,N_21912,N_21352);
and U22336 (N_22336,N_21247,N_21120);
nor U22337 (N_22337,N_21923,N_21578);
and U22338 (N_22338,N_21073,N_21467);
or U22339 (N_22339,N_21576,N_21575);
and U22340 (N_22340,N_21207,N_21739);
nand U22341 (N_22341,N_21693,N_21020);
and U22342 (N_22342,N_21322,N_21307);
and U22343 (N_22343,N_21164,N_21850);
or U22344 (N_22344,N_21857,N_21764);
and U22345 (N_22345,N_21215,N_21272);
and U22346 (N_22346,N_21107,N_21441);
nand U22347 (N_22347,N_21597,N_21673);
or U22348 (N_22348,N_21660,N_21958);
or U22349 (N_22349,N_21652,N_21297);
nor U22350 (N_22350,N_21216,N_21379);
xnor U22351 (N_22351,N_21827,N_21711);
nor U22352 (N_22352,N_21804,N_21806);
and U22353 (N_22353,N_21070,N_21333);
xor U22354 (N_22354,N_21255,N_21947);
nor U22355 (N_22355,N_21906,N_21427);
or U22356 (N_22356,N_21133,N_21867);
or U22357 (N_22357,N_21527,N_21549);
xnor U22358 (N_22358,N_21204,N_21573);
nor U22359 (N_22359,N_21868,N_21591);
xnor U22360 (N_22360,N_21786,N_21069);
nand U22361 (N_22361,N_21854,N_21047);
nor U22362 (N_22362,N_21999,N_21775);
xnor U22363 (N_22363,N_21895,N_21731);
nand U22364 (N_22364,N_21813,N_21168);
xnor U22365 (N_22365,N_21397,N_21750);
and U22366 (N_22366,N_21248,N_21699);
and U22367 (N_22367,N_21097,N_21559);
and U22368 (N_22368,N_21983,N_21452);
nand U22369 (N_22369,N_21175,N_21354);
xnor U22370 (N_22370,N_21067,N_21522);
and U22371 (N_22371,N_21138,N_21267);
and U22372 (N_22372,N_21991,N_21284);
xor U22373 (N_22373,N_21118,N_21293);
nor U22374 (N_22374,N_21988,N_21243);
xor U22375 (N_22375,N_21406,N_21037);
and U22376 (N_22376,N_21192,N_21494);
or U22377 (N_22377,N_21408,N_21404);
nand U22378 (N_22378,N_21794,N_21101);
and U22379 (N_22379,N_21944,N_21875);
nand U22380 (N_22380,N_21440,N_21749);
and U22381 (N_22381,N_21030,N_21697);
or U22382 (N_22382,N_21381,N_21220);
xor U22383 (N_22383,N_21217,N_21108);
and U22384 (N_22384,N_21038,N_21486);
nand U22385 (N_22385,N_21670,N_21237);
xnor U22386 (N_22386,N_21643,N_21460);
and U22387 (N_22387,N_21803,N_21157);
xor U22388 (N_22388,N_21407,N_21928);
nand U22389 (N_22389,N_21872,N_21362);
nand U22390 (N_22390,N_21855,N_21918);
nand U22391 (N_22391,N_21470,N_21622);
and U22392 (N_22392,N_21465,N_21826);
nor U22393 (N_22393,N_21281,N_21179);
nor U22394 (N_22394,N_21369,N_21628);
nor U22395 (N_22395,N_21708,N_21147);
xnor U22396 (N_22396,N_21688,N_21475);
and U22397 (N_22397,N_21833,N_21967);
and U22398 (N_22398,N_21548,N_21523);
nand U22399 (N_22399,N_21706,N_21547);
or U22400 (N_22400,N_21320,N_21392);
or U22401 (N_22401,N_21142,N_21884);
nand U22402 (N_22402,N_21148,N_21934);
nor U22403 (N_22403,N_21966,N_21604);
xor U22404 (N_22404,N_21626,N_21822);
or U22405 (N_22405,N_21011,N_21902);
and U22406 (N_22406,N_21910,N_21719);
xor U22407 (N_22407,N_21344,N_21139);
and U22408 (N_22408,N_21145,N_21162);
nand U22409 (N_22409,N_21644,N_21552);
or U22410 (N_22410,N_21870,N_21840);
nor U22411 (N_22411,N_21916,N_21861);
nor U22412 (N_22412,N_21202,N_21076);
nor U22413 (N_22413,N_21811,N_21913);
nor U22414 (N_22414,N_21668,N_21621);
xor U22415 (N_22415,N_21196,N_21252);
and U22416 (N_22416,N_21975,N_21709);
nor U22417 (N_22417,N_21831,N_21607);
or U22418 (N_22418,N_21239,N_21515);
or U22419 (N_22419,N_21695,N_21676);
xnor U22420 (N_22420,N_21489,N_21851);
nand U22421 (N_22421,N_21432,N_21376);
nor U22422 (N_22422,N_21420,N_21919);
nand U22423 (N_22423,N_21443,N_21946);
xor U22424 (N_22424,N_21149,N_21635);
and U22425 (N_22425,N_21791,N_21336);
nand U22426 (N_22426,N_21978,N_21698);
nand U22427 (N_22427,N_21675,N_21275);
nand U22428 (N_22428,N_21507,N_21289);
nor U22429 (N_22429,N_21812,N_21506);
and U22430 (N_22430,N_21599,N_21816);
or U22431 (N_22431,N_21004,N_21639);
or U22432 (N_22432,N_21502,N_21878);
and U22433 (N_22433,N_21040,N_21265);
nor U22434 (N_22434,N_21143,N_21633);
or U22435 (N_22435,N_21866,N_21491);
and U22436 (N_22436,N_21899,N_21092);
and U22437 (N_22437,N_21533,N_21128);
nand U22438 (N_22438,N_21730,N_21824);
or U22439 (N_22439,N_21231,N_21188);
xnor U22440 (N_22440,N_21187,N_21787);
nand U22441 (N_22441,N_21956,N_21524);
xor U22442 (N_22442,N_21817,N_21033);
nor U22443 (N_22443,N_21964,N_21085);
and U22444 (N_22444,N_21562,N_21891);
or U22445 (N_22445,N_21616,N_21801);
nor U22446 (N_22446,N_21350,N_21683);
nor U22447 (N_22447,N_21184,N_21053);
xnor U22448 (N_22448,N_21935,N_21388);
or U22449 (N_22449,N_21389,N_21525);
nor U22450 (N_22450,N_21129,N_21634);
or U22451 (N_22451,N_21428,N_21888);
nand U22452 (N_22452,N_21413,N_21071);
xor U22453 (N_22453,N_21434,N_21119);
nand U22454 (N_22454,N_21993,N_21332);
and U22455 (N_22455,N_21758,N_21064);
and U22456 (N_22456,N_21539,N_21402);
or U22457 (N_22457,N_21844,N_21348);
nor U22458 (N_22458,N_21057,N_21036);
nor U22459 (N_22459,N_21485,N_21898);
xor U22460 (N_22460,N_21538,N_21569);
nor U22461 (N_22461,N_21545,N_21461);
nand U22462 (N_22462,N_21722,N_21940);
or U22463 (N_22463,N_21152,N_21262);
or U22464 (N_22464,N_21531,N_21125);
and U22465 (N_22465,N_21173,N_21763);
nor U22466 (N_22466,N_21647,N_21700);
nor U22467 (N_22467,N_21480,N_21632);
xor U22468 (N_22468,N_21312,N_21403);
nand U22469 (N_22469,N_21328,N_21807);
xnor U22470 (N_22470,N_21897,N_21667);
xnor U22471 (N_22471,N_21140,N_21989);
and U22472 (N_22472,N_21858,N_21065);
and U22473 (N_22473,N_21274,N_21586);
and U22474 (N_22474,N_21687,N_21034);
nor U22475 (N_22475,N_21270,N_21974);
nand U22476 (N_22476,N_21444,N_21553);
xor U22477 (N_22477,N_21930,N_21920);
xor U22478 (N_22478,N_21984,N_21809);
or U22479 (N_22479,N_21249,N_21292);
or U22480 (N_22480,N_21818,N_21224);
xor U22481 (N_22481,N_21648,N_21150);
nand U22482 (N_22482,N_21448,N_21618);
nand U22483 (N_22483,N_21503,N_21948);
xnor U22484 (N_22484,N_21985,N_21081);
nor U22485 (N_22485,N_21704,N_21973);
xnor U22486 (N_22486,N_21994,N_21124);
nor U22487 (N_22487,N_21194,N_21883);
nor U22488 (N_22488,N_21169,N_21746);
and U22489 (N_22489,N_21805,N_21018);
and U22490 (N_22490,N_21301,N_21326);
nand U22491 (N_22491,N_21568,N_21835);
nand U22492 (N_22492,N_21308,N_21105);
and U22493 (N_22493,N_21141,N_21313);
and U22494 (N_22494,N_21734,N_21512);
or U22495 (N_22495,N_21829,N_21570);
or U22496 (N_22496,N_21049,N_21356);
nand U22497 (N_22497,N_21871,N_21288);
nand U22498 (N_22498,N_21165,N_21927);
nor U22499 (N_22499,N_21976,N_21395);
nand U22500 (N_22500,N_21189,N_21382);
or U22501 (N_22501,N_21513,N_21881);
xnor U22502 (N_22502,N_21484,N_21150);
or U22503 (N_22503,N_21561,N_21037);
nand U22504 (N_22504,N_21455,N_21029);
nor U22505 (N_22505,N_21010,N_21492);
and U22506 (N_22506,N_21988,N_21723);
and U22507 (N_22507,N_21368,N_21520);
nand U22508 (N_22508,N_21090,N_21708);
or U22509 (N_22509,N_21050,N_21310);
and U22510 (N_22510,N_21332,N_21691);
nor U22511 (N_22511,N_21662,N_21882);
nand U22512 (N_22512,N_21660,N_21270);
nor U22513 (N_22513,N_21287,N_21337);
xor U22514 (N_22514,N_21356,N_21680);
nand U22515 (N_22515,N_21397,N_21999);
nand U22516 (N_22516,N_21445,N_21802);
xnor U22517 (N_22517,N_21054,N_21223);
nand U22518 (N_22518,N_21190,N_21427);
nor U22519 (N_22519,N_21476,N_21821);
or U22520 (N_22520,N_21392,N_21775);
and U22521 (N_22521,N_21309,N_21201);
nand U22522 (N_22522,N_21090,N_21351);
nand U22523 (N_22523,N_21865,N_21291);
and U22524 (N_22524,N_21084,N_21961);
nand U22525 (N_22525,N_21236,N_21521);
and U22526 (N_22526,N_21525,N_21725);
nor U22527 (N_22527,N_21926,N_21764);
xor U22528 (N_22528,N_21803,N_21510);
nand U22529 (N_22529,N_21161,N_21329);
xnor U22530 (N_22530,N_21892,N_21770);
nor U22531 (N_22531,N_21989,N_21052);
nand U22532 (N_22532,N_21618,N_21036);
or U22533 (N_22533,N_21511,N_21982);
nor U22534 (N_22534,N_21158,N_21321);
and U22535 (N_22535,N_21723,N_21771);
and U22536 (N_22536,N_21311,N_21518);
nand U22537 (N_22537,N_21113,N_21106);
xor U22538 (N_22538,N_21586,N_21905);
and U22539 (N_22539,N_21549,N_21035);
and U22540 (N_22540,N_21024,N_21983);
nor U22541 (N_22541,N_21353,N_21318);
xor U22542 (N_22542,N_21269,N_21362);
nand U22543 (N_22543,N_21242,N_21207);
xnor U22544 (N_22544,N_21648,N_21205);
or U22545 (N_22545,N_21218,N_21665);
nor U22546 (N_22546,N_21403,N_21818);
nand U22547 (N_22547,N_21988,N_21391);
xor U22548 (N_22548,N_21768,N_21452);
nor U22549 (N_22549,N_21037,N_21229);
nand U22550 (N_22550,N_21994,N_21903);
nor U22551 (N_22551,N_21773,N_21069);
and U22552 (N_22552,N_21282,N_21593);
or U22553 (N_22553,N_21112,N_21902);
or U22554 (N_22554,N_21934,N_21826);
xor U22555 (N_22555,N_21230,N_21626);
xnor U22556 (N_22556,N_21922,N_21767);
xor U22557 (N_22557,N_21556,N_21072);
and U22558 (N_22558,N_21860,N_21630);
nand U22559 (N_22559,N_21483,N_21371);
and U22560 (N_22560,N_21092,N_21772);
or U22561 (N_22561,N_21315,N_21200);
or U22562 (N_22562,N_21485,N_21590);
nor U22563 (N_22563,N_21072,N_21312);
nor U22564 (N_22564,N_21498,N_21207);
nor U22565 (N_22565,N_21862,N_21475);
nor U22566 (N_22566,N_21688,N_21152);
nor U22567 (N_22567,N_21036,N_21415);
and U22568 (N_22568,N_21782,N_21115);
nand U22569 (N_22569,N_21738,N_21745);
or U22570 (N_22570,N_21086,N_21682);
nor U22571 (N_22571,N_21101,N_21633);
or U22572 (N_22572,N_21111,N_21487);
nand U22573 (N_22573,N_21870,N_21773);
xor U22574 (N_22574,N_21169,N_21850);
or U22575 (N_22575,N_21942,N_21318);
nor U22576 (N_22576,N_21086,N_21520);
or U22577 (N_22577,N_21458,N_21721);
and U22578 (N_22578,N_21827,N_21771);
nand U22579 (N_22579,N_21965,N_21604);
or U22580 (N_22580,N_21873,N_21622);
and U22581 (N_22581,N_21411,N_21392);
nor U22582 (N_22582,N_21234,N_21281);
nor U22583 (N_22583,N_21871,N_21827);
or U22584 (N_22584,N_21206,N_21551);
nand U22585 (N_22585,N_21449,N_21171);
nand U22586 (N_22586,N_21486,N_21478);
and U22587 (N_22587,N_21032,N_21419);
nor U22588 (N_22588,N_21339,N_21191);
nand U22589 (N_22589,N_21507,N_21017);
xnor U22590 (N_22590,N_21288,N_21221);
xnor U22591 (N_22591,N_21546,N_21336);
or U22592 (N_22592,N_21596,N_21443);
nor U22593 (N_22593,N_21363,N_21123);
nand U22594 (N_22594,N_21151,N_21493);
nor U22595 (N_22595,N_21659,N_21069);
and U22596 (N_22596,N_21247,N_21940);
and U22597 (N_22597,N_21654,N_21274);
nor U22598 (N_22598,N_21467,N_21043);
xor U22599 (N_22599,N_21174,N_21780);
nand U22600 (N_22600,N_21562,N_21450);
and U22601 (N_22601,N_21890,N_21849);
xor U22602 (N_22602,N_21897,N_21096);
nand U22603 (N_22603,N_21242,N_21452);
or U22604 (N_22604,N_21342,N_21383);
xor U22605 (N_22605,N_21590,N_21091);
xnor U22606 (N_22606,N_21824,N_21281);
xnor U22607 (N_22607,N_21661,N_21948);
nand U22608 (N_22608,N_21762,N_21354);
nand U22609 (N_22609,N_21654,N_21353);
and U22610 (N_22610,N_21805,N_21051);
xor U22611 (N_22611,N_21454,N_21685);
nor U22612 (N_22612,N_21136,N_21651);
xnor U22613 (N_22613,N_21172,N_21091);
nor U22614 (N_22614,N_21110,N_21353);
and U22615 (N_22615,N_21212,N_21004);
nand U22616 (N_22616,N_21669,N_21115);
xnor U22617 (N_22617,N_21825,N_21720);
and U22618 (N_22618,N_21696,N_21976);
xnor U22619 (N_22619,N_21283,N_21926);
nand U22620 (N_22620,N_21406,N_21546);
nor U22621 (N_22621,N_21630,N_21922);
nand U22622 (N_22622,N_21562,N_21604);
or U22623 (N_22623,N_21743,N_21392);
or U22624 (N_22624,N_21334,N_21247);
or U22625 (N_22625,N_21866,N_21009);
and U22626 (N_22626,N_21942,N_21289);
and U22627 (N_22627,N_21309,N_21076);
or U22628 (N_22628,N_21413,N_21313);
or U22629 (N_22629,N_21725,N_21155);
and U22630 (N_22630,N_21583,N_21721);
xnor U22631 (N_22631,N_21769,N_21870);
xnor U22632 (N_22632,N_21778,N_21410);
or U22633 (N_22633,N_21683,N_21399);
nor U22634 (N_22634,N_21921,N_21276);
xor U22635 (N_22635,N_21925,N_21770);
nand U22636 (N_22636,N_21067,N_21465);
nor U22637 (N_22637,N_21659,N_21521);
and U22638 (N_22638,N_21426,N_21830);
and U22639 (N_22639,N_21790,N_21064);
and U22640 (N_22640,N_21928,N_21277);
xor U22641 (N_22641,N_21047,N_21894);
nor U22642 (N_22642,N_21736,N_21219);
xor U22643 (N_22643,N_21356,N_21152);
and U22644 (N_22644,N_21859,N_21982);
nand U22645 (N_22645,N_21843,N_21620);
nand U22646 (N_22646,N_21613,N_21637);
nand U22647 (N_22647,N_21158,N_21141);
or U22648 (N_22648,N_21313,N_21883);
or U22649 (N_22649,N_21291,N_21708);
xor U22650 (N_22650,N_21004,N_21624);
or U22651 (N_22651,N_21284,N_21256);
nand U22652 (N_22652,N_21925,N_21156);
nor U22653 (N_22653,N_21203,N_21079);
nand U22654 (N_22654,N_21251,N_21913);
xnor U22655 (N_22655,N_21804,N_21294);
and U22656 (N_22656,N_21843,N_21084);
nand U22657 (N_22657,N_21543,N_21263);
nand U22658 (N_22658,N_21517,N_21064);
and U22659 (N_22659,N_21975,N_21096);
nor U22660 (N_22660,N_21214,N_21344);
xnor U22661 (N_22661,N_21021,N_21493);
or U22662 (N_22662,N_21263,N_21667);
nor U22663 (N_22663,N_21807,N_21894);
and U22664 (N_22664,N_21852,N_21501);
nand U22665 (N_22665,N_21275,N_21600);
nand U22666 (N_22666,N_21191,N_21224);
and U22667 (N_22667,N_21738,N_21432);
and U22668 (N_22668,N_21515,N_21085);
xnor U22669 (N_22669,N_21025,N_21294);
and U22670 (N_22670,N_21155,N_21118);
nand U22671 (N_22671,N_21576,N_21366);
xor U22672 (N_22672,N_21389,N_21533);
xnor U22673 (N_22673,N_21911,N_21470);
or U22674 (N_22674,N_21739,N_21564);
nand U22675 (N_22675,N_21616,N_21026);
or U22676 (N_22676,N_21791,N_21464);
nor U22677 (N_22677,N_21287,N_21389);
nor U22678 (N_22678,N_21385,N_21422);
xnor U22679 (N_22679,N_21693,N_21541);
xnor U22680 (N_22680,N_21957,N_21434);
nand U22681 (N_22681,N_21200,N_21664);
xnor U22682 (N_22682,N_21624,N_21087);
nor U22683 (N_22683,N_21989,N_21585);
nor U22684 (N_22684,N_21114,N_21550);
nor U22685 (N_22685,N_21972,N_21365);
and U22686 (N_22686,N_21423,N_21286);
nand U22687 (N_22687,N_21254,N_21024);
nor U22688 (N_22688,N_21655,N_21127);
xnor U22689 (N_22689,N_21168,N_21935);
and U22690 (N_22690,N_21549,N_21579);
nand U22691 (N_22691,N_21478,N_21188);
nor U22692 (N_22692,N_21546,N_21161);
xnor U22693 (N_22693,N_21223,N_21076);
and U22694 (N_22694,N_21961,N_21428);
or U22695 (N_22695,N_21848,N_21480);
nor U22696 (N_22696,N_21548,N_21009);
nand U22697 (N_22697,N_21428,N_21177);
and U22698 (N_22698,N_21773,N_21993);
or U22699 (N_22699,N_21223,N_21400);
or U22700 (N_22700,N_21212,N_21243);
or U22701 (N_22701,N_21770,N_21718);
and U22702 (N_22702,N_21304,N_21162);
nor U22703 (N_22703,N_21075,N_21639);
and U22704 (N_22704,N_21328,N_21693);
or U22705 (N_22705,N_21692,N_21615);
nor U22706 (N_22706,N_21829,N_21463);
nor U22707 (N_22707,N_21603,N_21179);
xnor U22708 (N_22708,N_21130,N_21271);
or U22709 (N_22709,N_21939,N_21457);
or U22710 (N_22710,N_21298,N_21064);
xnor U22711 (N_22711,N_21385,N_21053);
nand U22712 (N_22712,N_21597,N_21436);
nand U22713 (N_22713,N_21985,N_21479);
xor U22714 (N_22714,N_21899,N_21764);
nand U22715 (N_22715,N_21106,N_21384);
nand U22716 (N_22716,N_21757,N_21889);
and U22717 (N_22717,N_21532,N_21955);
nand U22718 (N_22718,N_21263,N_21284);
nand U22719 (N_22719,N_21683,N_21823);
xnor U22720 (N_22720,N_21177,N_21298);
xor U22721 (N_22721,N_21406,N_21517);
or U22722 (N_22722,N_21885,N_21577);
xnor U22723 (N_22723,N_21604,N_21823);
xor U22724 (N_22724,N_21732,N_21361);
xor U22725 (N_22725,N_21992,N_21396);
nand U22726 (N_22726,N_21508,N_21276);
nor U22727 (N_22727,N_21020,N_21255);
or U22728 (N_22728,N_21752,N_21254);
nor U22729 (N_22729,N_21761,N_21206);
nor U22730 (N_22730,N_21542,N_21633);
xnor U22731 (N_22731,N_21725,N_21533);
nand U22732 (N_22732,N_21525,N_21532);
or U22733 (N_22733,N_21238,N_21142);
nor U22734 (N_22734,N_21656,N_21091);
xor U22735 (N_22735,N_21997,N_21601);
xor U22736 (N_22736,N_21836,N_21243);
and U22737 (N_22737,N_21056,N_21877);
nand U22738 (N_22738,N_21419,N_21907);
nor U22739 (N_22739,N_21805,N_21483);
nor U22740 (N_22740,N_21585,N_21254);
nor U22741 (N_22741,N_21512,N_21976);
or U22742 (N_22742,N_21432,N_21664);
nor U22743 (N_22743,N_21806,N_21678);
nand U22744 (N_22744,N_21168,N_21387);
nand U22745 (N_22745,N_21889,N_21582);
and U22746 (N_22746,N_21556,N_21273);
or U22747 (N_22747,N_21806,N_21852);
nor U22748 (N_22748,N_21839,N_21531);
nand U22749 (N_22749,N_21387,N_21427);
nand U22750 (N_22750,N_21955,N_21270);
or U22751 (N_22751,N_21625,N_21804);
nand U22752 (N_22752,N_21706,N_21276);
xnor U22753 (N_22753,N_21147,N_21181);
nand U22754 (N_22754,N_21200,N_21668);
nor U22755 (N_22755,N_21785,N_21406);
and U22756 (N_22756,N_21877,N_21405);
nor U22757 (N_22757,N_21364,N_21544);
xor U22758 (N_22758,N_21320,N_21555);
nand U22759 (N_22759,N_21343,N_21717);
xnor U22760 (N_22760,N_21784,N_21994);
and U22761 (N_22761,N_21412,N_21263);
or U22762 (N_22762,N_21061,N_21822);
nand U22763 (N_22763,N_21103,N_21041);
nand U22764 (N_22764,N_21771,N_21274);
or U22765 (N_22765,N_21657,N_21269);
xnor U22766 (N_22766,N_21811,N_21883);
nand U22767 (N_22767,N_21322,N_21804);
nor U22768 (N_22768,N_21829,N_21560);
xor U22769 (N_22769,N_21282,N_21942);
nand U22770 (N_22770,N_21300,N_21432);
nand U22771 (N_22771,N_21985,N_21100);
and U22772 (N_22772,N_21598,N_21766);
and U22773 (N_22773,N_21785,N_21452);
and U22774 (N_22774,N_21860,N_21106);
nand U22775 (N_22775,N_21074,N_21170);
and U22776 (N_22776,N_21613,N_21282);
and U22777 (N_22777,N_21659,N_21453);
or U22778 (N_22778,N_21615,N_21216);
nand U22779 (N_22779,N_21892,N_21912);
or U22780 (N_22780,N_21003,N_21876);
nor U22781 (N_22781,N_21733,N_21915);
nor U22782 (N_22782,N_21631,N_21875);
and U22783 (N_22783,N_21421,N_21886);
or U22784 (N_22784,N_21451,N_21729);
xnor U22785 (N_22785,N_21567,N_21235);
xor U22786 (N_22786,N_21814,N_21624);
or U22787 (N_22787,N_21389,N_21453);
xnor U22788 (N_22788,N_21154,N_21084);
xor U22789 (N_22789,N_21095,N_21008);
and U22790 (N_22790,N_21433,N_21565);
xnor U22791 (N_22791,N_21456,N_21572);
xnor U22792 (N_22792,N_21451,N_21251);
xor U22793 (N_22793,N_21511,N_21203);
nor U22794 (N_22794,N_21524,N_21933);
or U22795 (N_22795,N_21794,N_21392);
nand U22796 (N_22796,N_21344,N_21765);
nand U22797 (N_22797,N_21850,N_21749);
or U22798 (N_22798,N_21834,N_21970);
nand U22799 (N_22799,N_21497,N_21061);
nor U22800 (N_22800,N_21807,N_21404);
xor U22801 (N_22801,N_21433,N_21019);
xor U22802 (N_22802,N_21368,N_21053);
nor U22803 (N_22803,N_21474,N_21211);
nor U22804 (N_22804,N_21441,N_21763);
nand U22805 (N_22805,N_21478,N_21248);
and U22806 (N_22806,N_21771,N_21119);
nor U22807 (N_22807,N_21921,N_21624);
xor U22808 (N_22808,N_21602,N_21889);
or U22809 (N_22809,N_21473,N_21872);
or U22810 (N_22810,N_21390,N_21235);
xnor U22811 (N_22811,N_21630,N_21814);
nor U22812 (N_22812,N_21778,N_21839);
and U22813 (N_22813,N_21158,N_21181);
or U22814 (N_22814,N_21510,N_21749);
nor U22815 (N_22815,N_21694,N_21853);
nor U22816 (N_22816,N_21407,N_21411);
and U22817 (N_22817,N_21430,N_21155);
xor U22818 (N_22818,N_21288,N_21905);
nor U22819 (N_22819,N_21355,N_21819);
nand U22820 (N_22820,N_21098,N_21777);
or U22821 (N_22821,N_21004,N_21777);
nor U22822 (N_22822,N_21331,N_21870);
and U22823 (N_22823,N_21336,N_21870);
or U22824 (N_22824,N_21102,N_21622);
or U22825 (N_22825,N_21791,N_21230);
xnor U22826 (N_22826,N_21969,N_21030);
or U22827 (N_22827,N_21846,N_21446);
or U22828 (N_22828,N_21313,N_21810);
nand U22829 (N_22829,N_21189,N_21712);
nand U22830 (N_22830,N_21209,N_21677);
nor U22831 (N_22831,N_21784,N_21132);
xnor U22832 (N_22832,N_21782,N_21012);
nor U22833 (N_22833,N_21759,N_21710);
nand U22834 (N_22834,N_21823,N_21425);
xor U22835 (N_22835,N_21861,N_21311);
and U22836 (N_22836,N_21736,N_21760);
and U22837 (N_22837,N_21620,N_21517);
xor U22838 (N_22838,N_21677,N_21600);
or U22839 (N_22839,N_21049,N_21843);
and U22840 (N_22840,N_21664,N_21366);
or U22841 (N_22841,N_21965,N_21021);
xnor U22842 (N_22842,N_21491,N_21583);
and U22843 (N_22843,N_21107,N_21522);
xor U22844 (N_22844,N_21550,N_21682);
and U22845 (N_22845,N_21244,N_21144);
nand U22846 (N_22846,N_21139,N_21737);
nor U22847 (N_22847,N_21298,N_21189);
or U22848 (N_22848,N_21228,N_21638);
or U22849 (N_22849,N_21797,N_21554);
and U22850 (N_22850,N_21288,N_21461);
and U22851 (N_22851,N_21691,N_21162);
or U22852 (N_22852,N_21031,N_21576);
and U22853 (N_22853,N_21915,N_21199);
nor U22854 (N_22854,N_21109,N_21882);
nand U22855 (N_22855,N_21361,N_21321);
nor U22856 (N_22856,N_21719,N_21759);
nor U22857 (N_22857,N_21106,N_21079);
or U22858 (N_22858,N_21155,N_21531);
xor U22859 (N_22859,N_21851,N_21528);
and U22860 (N_22860,N_21999,N_21734);
nor U22861 (N_22861,N_21983,N_21149);
nor U22862 (N_22862,N_21126,N_21118);
xnor U22863 (N_22863,N_21312,N_21827);
and U22864 (N_22864,N_21241,N_21186);
nand U22865 (N_22865,N_21286,N_21851);
nor U22866 (N_22866,N_21685,N_21072);
and U22867 (N_22867,N_21812,N_21325);
xor U22868 (N_22868,N_21336,N_21939);
xor U22869 (N_22869,N_21597,N_21076);
and U22870 (N_22870,N_21489,N_21997);
nand U22871 (N_22871,N_21795,N_21666);
nor U22872 (N_22872,N_21783,N_21563);
nor U22873 (N_22873,N_21671,N_21644);
and U22874 (N_22874,N_21457,N_21921);
nand U22875 (N_22875,N_21836,N_21101);
nand U22876 (N_22876,N_21558,N_21983);
nor U22877 (N_22877,N_21510,N_21227);
nor U22878 (N_22878,N_21415,N_21857);
and U22879 (N_22879,N_21966,N_21933);
or U22880 (N_22880,N_21583,N_21770);
nand U22881 (N_22881,N_21598,N_21053);
nand U22882 (N_22882,N_21647,N_21120);
or U22883 (N_22883,N_21201,N_21333);
nor U22884 (N_22884,N_21913,N_21279);
and U22885 (N_22885,N_21903,N_21648);
or U22886 (N_22886,N_21494,N_21789);
nor U22887 (N_22887,N_21059,N_21959);
nor U22888 (N_22888,N_21595,N_21330);
nor U22889 (N_22889,N_21761,N_21917);
xor U22890 (N_22890,N_21728,N_21841);
nor U22891 (N_22891,N_21740,N_21533);
or U22892 (N_22892,N_21624,N_21739);
and U22893 (N_22893,N_21129,N_21579);
nor U22894 (N_22894,N_21631,N_21091);
and U22895 (N_22895,N_21801,N_21622);
or U22896 (N_22896,N_21170,N_21441);
nor U22897 (N_22897,N_21029,N_21892);
and U22898 (N_22898,N_21671,N_21712);
xor U22899 (N_22899,N_21072,N_21530);
and U22900 (N_22900,N_21439,N_21337);
nand U22901 (N_22901,N_21395,N_21537);
or U22902 (N_22902,N_21229,N_21279);
and U22903 (N_22903,N_21687,N_21539);
nand U22904 (N_22904,N_21842,N_21893);
and U22905 (N_22905,N_21784,N_21325);
or U22906 (N_22906,N_21088,N_21936);
nor U22907 (N_22907,N_21174,N_21750);
nand U22908 (N_22908,N_21304,N_21215);
or U22909 (N_22909,N_21493,N_21445);
nand U22910 (N_22910,N_21887,N_21838);
or U22911 (N_22911,N_21763,N_21273);
nand U22912 (N_22912,N_21376,N_21230);
nand U22913 (N_22913,N_21614,N_21942);
or U22914 (N_22914,N_21498,N_21951);
xor U22915 (N_22915,N_21131,N_21645);
or U22916 (N_22916,N_21614,N_21194);
xor U22917 (N_22917,N_21366,N_21228);
nor U22918 (N_22918,N_21190,N_21648);
and U22919 (N_22919,N_21949,N_21197);
xnor U22920 (N_22920,N_21338,N_21075);
and U22921 (N_22921,N_21463,N_21792);
xor U22922 (N_22922,N_21029,N_21986);
xor U22923 (N_22923,N_21621,N_21030);
or U22924 (N_22924,N_21793,N_21106);
nand U22925 (N_22925,N_21940,N_21842);
and U22926 (N_22926,N_21890,N_21087);
and U22927 (N_22927,N_21739,N_21603);
xor U22928 (N_22928,N_21305,N_21708);
or U22929 (N_22929,N_21013,N_21517);
and U22930 (N_22930,N_21254,N_21378);
and U22931 (N_22931,N_21525,N_21047);
xnor U22932 (N_22932,N_21237,N_21780);
nor U22933 (N_22933,N_21039,N_21042);
xor U22934 (N_22934,N_21022,N_21980);
xnor U22935 (N_22935,N_21463,N_21760);
nor U22936 (N_22936,N_21693,N_21261);
or U22937 (N_22937,N_21698,N_21837);
nand U22938 (N_22938,N_21623,N_21632);
nand U22939 (N_22939,N_21922,N_21558);
xnor U22940 (N_22940,N_21462,N_21445);
nand U22941 (N_22941,N_21072,N_21627);
and U22942 (N_22942,N_21589,N_21910);
or U22943 (N_22943,N_21067,N_21832);
xor U22944 (N_22944,N_21326,N_21022);
or U22945 (N_22945,N_21897,N_21316);
or U22946 (N_22946,N_21788,N_21856);
and U22947 (N_22947,N_21136,N_21309);
nand U22948 (N_22948,N_21610,N_21688);
nor U22949 (N_22949,N_21185,N_21695);
and U22950 (N_22950,N_21887,N_21394);
or U22951 (N_22951,N_21251,N_21005);
nor U22952 (N_22952,N_21065,N_21094);
or U22953 (N_22953,N_21678,N_21519);
and U22954 (N_22954,N_21906,N_21264);
nand U22955 (N_22955,N_21788,N_21746);
xnor U22956 (N_22956,N_21382,N_21167);
xor U22957 (N_22957,N_21153,N_21447);
and U22958 (N_22958,N_21923,N_21681);
nand U22959 (N_22959,N_21030,N_21050);
or U22960 (N_22960,N_21630,N_21640);
xor U22961 (N_22961,N_21371,N_21390);
xnor U22962 (N_22962,N_21450,N_21665);
nor U22963 (N_22963,N_21733,N_21983);
xor U22964 (N_22964,N_21413,N_21665);
or U22965 (N_22965,N_21536,N_21120);
xor U22966 (N_22966,N_21297,N_21204);
or U22967 (N_22967,N_21994,N_21471);
nand U22968 (N_22968,N_21081,N_21179);
nor U22969 (N_22969,N_21693,N_21925);
and U22970 (N_22970,N_21058,N_21303);
xor U22971 (N_22971,N_21571,N_21899);
or U22972 (N_22972,N_21335,N_21786);
nor U22973 (N_22973,N_21295,N_21827);
and U22974 (N_22974,N_21851,N_21598);
and U22975 (N_22975,N_21217,N_21014);
or U22976 (N_22976,N_21093,N_21150);
nand U22977 (N_22977,N_21908,N_21688);
nor U22978 (N_22978,N_21807,N_21908);
nor U22979 (N_22979,N_21984,N_21403);
xnor U22980 (N_22980,N_21827,N_21928);
or U22981 (N_22981,N_21464,N_21273);
xnor U22982 (N_22982,N_21028,N_21524);
or U22983 (N_22983,N_21548,N_21866);
and U22984 (N_22984,N_21683,N_21731);
xnor U22985 (N_22985,N_21372,N_21547);
xnor U22986 (N_22986,N_21066,N_21607);
nand U22987 (N_22987,N_21013,N_21322);
nand U22988 (N_22988,N_21713,N_21851);
xor U22989 (N_22989,N_21532,N_21583);
and U22990 (N_22990,N_21611,N_21854);
and U22991 (N_22991,N_21272,N_21869);
nand U22992 (N_22992,N_21468,N_21901);
nor U22993 (N_22993,N_21268,N_21916);
and U22994 (N_22994,N_21816,N_21409);
nor U22995 (N_22995,N_21890,N_21705);
or U22996 (N_22996,N_21389,N_21954);
nor U22997 (N_22997,N_21854,N_21996);
and U22998 (N_22998,N_21250,N_21829);
and U22999 (N_22999,N_21387,N_21290);
or U23000 (N_23000,N_22262,N_22969);
nor U23001 (N_23001,N_22219,N_22248);
or U23002 (N_23002,N_22561,N_22827);
and U23003 (N_23003,N_22281,N_22451);
xor U23004 (N_23004,N_22263,N_22837);
nor U23005 (N_23005,N_22950,N_22095);
and U23006 (N_23006,N_22133,N_22325);
nand U23007 (N_23007,N_22205,N_22454);
and U23008 (N_23008,N_22960,N_22329);
nor U23009 (N_23009,N_22218,N_22925);
nor U23010 (N_23010,N_22384,N_22268);
nor U23011 (N_23011,N_22241,N_22479);
nand U23012 (N_23012,N_22171,N_22440);
nand U23013 (N_23013,N_22422,N_22142);
and U23014 (N_23014,N_22695,N_22784);
nor U23015 (N_23015,N_22944,N_22773);
xnor U23016 (N_23016,N_22506,N_22723);
or U23017 (N_23017,N_22697,N_22802);
or U23018 (N_23018,N_22852,N_22733);
and U23019 (N_23019,N_22487,N_22242);
xnor U23020 (N_23020,N_22126,N_22476);
xor U23021 (N_23021,N_22610,N_22534);
and U23022 (N_23022,N_22257,N_22707);
and U23023 (N_23023,N_22352,N_22047);
and U23024 (N_23024,N_22520,N_22536);
xor U23025 (N_23025,N_22220,N_22799);
or U23026 (N_23026,N_22350,N_22264);
and U23027 (N_23027,N_22307,N_22050);
and U23028 (N_23028,N_22470,N_22651);
nand U23029 (N_23029,N_22767,N_22239);
and U23030 (N_23030,N_22668,N_22083);
or U23031 (N_23031,N_22472,N_22369);
or U23032 (N_23032,N_22914,N_22211);
xnor U23033 (N_23033,N_22190,N_22720);
and U23034 (N_23034,N_22014,N_22062);
and U23035 (N_23035,N_22687,N_22546);
nand U23036 (N_23036,N_22216,N_22521);
nand U23037 (N_23037,N_22669,N_22232);
nor U23038 (N_23038,N_22836,N_22726);
and U23039 (N_23039,N_22866,N_22448);
nand U23040 (N_23040,N_22402,N_22031);
xnor U23041 (N_23041,N_22727,N_22692);
nor U23042 (N_23042,N_22990,N_22786);
nor U23043 (N_23043,N_22735,N_22603);
nor U23044 (N_23044,N_22922,N_22652);
and U23045 (N_23045,N_22309,N_22404);
nand U23046 (N_23046,N_22102,N_22703);
xnor U23047 (N_23047,N_22233,N_22469);
nand U23048 (N_23048,N_22986,N_22206);
or U23049 (N_23049,N_22569,N_22801);
or U23050 (N_23050,N_22516,N_22373);
nand U23051 (N_23051,N_22838,N_22097);
or U23052 (N_23052,N_22478,N_22379);
xor U23053 (N_23053,N_22549,N_22121);
xor U23054 (N_23054,N_22928,N_22975);
xnor U23055 (N_23055,N_22061,N_22533);
and U23056 (N_23056,N_22443,N_22165);
or U23057 (N_23057,N_22435,N_22347);
nand U23058 (N_23058,N_22332,N_22674);
nor U23059 (N_23059,N_22391,N_22452);
or U23060 (N_23060,N_22236,N_22956);
or U23061 (N_23061,N_22084,N_22833);
nor U23062 (N_23062,N_22887,N_22064);
nand U23063 (N_23063,N_22888,N_22306);
nor U23064 (N_23064,N_22428,N_22623);
xnor U23065 (N_23065,N_22125,N_22071);
and U23066 (N_23066,N_22052,N_22834);
nor U23067 (N_23067,N_22434,N_22431);
xnor U23068 (N_23068,N_22529,N_22716);
nor U23069 (N_23069,N_22885,N_22804);
xnor U23070 (N_23070,N_22375,N_22486);
nor U23071 (N_23071,N_22629,N_22365);
nor U23072 (N_23072,N_22730,N_22869);
and U23073 (N_23073,N_22667,N_22895);
or U23074 (N_23074,N_22810,N_22210);
and U23075 (N_23075,N_22924,N_22442);
and U23076 (N_23076,N_22929,N_22049);
or U23077 (N_23077,N_22835,N_22675);
nand U23078 (N_23078,N_22983,N_22967);
nand U23079 (N_23079,N_22096,N_22468);
xor U23080 (N_23080,N_22297,N_22907);
nand U23081 (N_23081,N_22612,N_22955);
or U23082 (N_23082,N_22395,N_22698);
nand U23083 (N_23083,N_22457,N_22387);
or U23084 (N_23084,N_22338,N_22568);
and U23085 (N_23085,N_22854,N_22985);
and U23086 (N_23086,N_22266,N_22381);
nand U23087 (N_23087,N_22278,N_22065);
nor U23088 (N_23088,N_22634,N_22566);
or U23089 (N_23089,N_22656,N_22089);
nor U23090 (N_23090,N_22138,N_22140);
and U23091 (N_23091,N_22092,N_22245);
nand U23092 (N_23092,N_22542,N_22269);
nor U23093 (N_23093,N_22295,N_22413);
nor U23094 (N_23094,N_22234,N_22686);
nand U23095 (N_23095,N_22382,N_22937);
xnor U23096 (N_23096,N_22107,N_22565);
and U23097 (N_23097,N_22167,N_22615);
xnor U23098 (N_23098,N_22864,N_22367);
nor U23099 (N_23099,N_22587,N_22871);
nor U23100 (N_23100,N_22557,N_22886);
xnor U23101 (N_23101,N_22672,N_22409);
and U23102 (N_23102,N_22933,N_22574);
and U23103 (N_23103,N_22324,N_22116);
nor U23104 (N_23104,N_22737,N_22224);
or U23105 (N_23105,N_22830,N_22678);
or U23106 (N_23106,N_22068,N_22017);
nand U23107 (N_23107,N_22355,N_22754);
and U23108 (N_23108,N_22495,N_22082);
xor U23109 (N_23109,N_22340,N_22146);
and U23110 (N_23110,N_22290,N_22471);
and U23111 (N_23111,N_22039,N_22906);
and U23112 (N_23112,N_22770,N_22978);
nor U23113 (N_23113,N_22492,N_22890);
or U23114 (N_23114,N_22825,N_22203);
nand U23115 (N_23115,N_22644,N_22556);
xnor U23116 (N_23116,N_22905,N_22339);
xnor U23117 (N_23117,N_22988,N_22401);
xnor U23118 (N_23118,N_22093,N_22769);
xnor U23119 (N_23119,N_22514,N_22874);
and U23120 (N_23120,N_22625,N_22484);
or U23121 (N_23121,N_22054,N_22385);
xnor U23122 (N_23122,N_22993,N_22323);
nor U23123 (N_23123,N_22882,N_22115);
and U23124 (N_23124,N_22500,N_22821);
xor U23125 (N_23125,N_22035,N_22319);
or U23126 (N_23126,N_22923,N_22376);
or U23127 (N_23127,N_22345,N_22507);
nor U23128 (N_23128,N_22721,N_22671);
nor U23129 (N_23129,N_22392,N_22616);
xor U23130 (N_23130,N_22994,N_22676);
nand U23131 (N_23131,N_22328,N_22129);
nor U23132 (N_23132,N_22072,N_22526);
nor U23133 (N_23133,N_22456,N_22088);
xnor U23134 (N_23134,N_22560,N_22109);
nor U23135 (N_23135,N_22490,N_22460);
nor U23136 (N_23136,N_22894,N_22617);
or U23137 (N_23137,N_22540,N_22377);
and U23138 (N_23138,N_22594,N_22795);
nand U23139 (N_23139,N_22455,N_22078);
xnor U23140 (N_23140,N_22805,N_22518);
nand U23141 (N_23141,N_22026,N_22781);
nand U23142 (N_23142,N_22467,N_22363);
nor U23143 (N_23143,N_22511,N_22333);
and U23144 (N_23144,N_22912,N_22282);
xor U23145 (N_23145,N_22630,N_22627);
and U23146 (N_23146,N_22744,N_22745);
nand U23147 (N_23147,N_22003,N_22680);
nand U23148 (N_23148,N_22194,N_22981);
nand U23149 (N_23149,N_22356,N_22114);
nand U23150 (N_23150,N_22578,N_22868);
xnor U23151 (N_23151,N_22073,N_22284);
xnor U23152 (N_23152,N_22650,N_22762);
nand U23153 (N_23153,N_22554,N_22909);
or U23154 (N_23154,N_22398,N_22150);
nand U23155 (N_23155,N_22177,N_22724);
nor U23156 (N_23156,N_22645,N_22311);
nand U23157 (N_23157,N_22494,N_22664);
xor U23158 (N_23158,N_22601,N_22277);
and U23159 (N_23159,N_22036,N_22091);
nor U23160 (N_23160,N_22934,N_22798);
nor U23161 (N_23161,N_22335,N_22289);
and U23162 (N_23162,N_22648,N_22932);
nand U23163 (N_23163,N_22238,N_22020);
nor U23164 (N_23164,N_22747,N_22876);
nand U23165 (N_23165,N_22947,N_22168);
nor U23166 (N_23166,N_22702,N_22436);
and U23167 (N_23167,N_22719,N_22087);
nor U23168 (N_23168,N_22149,N_22544);
xnor U23169 (N_23169,N_22417,N_22229);
xor U23170 (N_23170,N_22419,N_22538);
xor U23171 (N_23171,N_22599,N_22493);
nor U23172 (N_23172,N_22286,N_22952);
nand U23173 (N_23173,N_22708,N_22600);
nor U23174 (N_23174,N_22447,N_22853);
xnor U23175 (N_23175,N_22408,N_22666);
and U23176 (N_23176,N_22274,N_22689);
nor U23177 (N_23177,N_22649,N_22900);
nand U23178 (N_23178,N_22372,N_22130);
or U23179 (N_23179,N_22972,N_22732);
nand U23180 (N_23180,N_22646,N_22429);
xnor U23181 (N_23181,N_22785,N_22998);
nand U23182 (N_23182,N_22011,N_22684);
or U23183 (N_23183,N_22742,N_22850);
nor U23184 (N_23184,N_22098,N_22197);
nor U23185 (N_23185,N_22973,N_22037);
and U23186 (N_23186,N_22293,N_22714);
and U23187 (N_23187,N_22539,N_22631);
nand U23188 (N_23188,N_22462,N_22639);
and U23189 (N_23189,N_22788,N_22946);
and U23190 (N_23190,N_22287,N_22371);
xor U23191 (N_23191,N_22410,N_22597);
nand U23192 (N_23192,N_22787,N_22915);
nand U23193 (N_23193,N_22080,N_22178);
nand U23194 (N_23194,N_22063,N_22883);
nand U23195 (N_23195,N_22368,N_22240);
and U23196 (N_23196,N_22041,N_22294);
nor U23197 (N_23197,N_22873,N_22193);
or U23198 (N_23198,N_22326,N_22661);
nor U23199 (N_23199,N_22420,N_22814);
nand U23200 (N_23200,N_22212,N_22145);
xor U23201 (N_23201,N_22693,N_22127);
and U23202 (N_23202,N_22132,N_22483);
xnor U23203 (N_23203,N_22665,N_22485);
and U23204 (N_23204,N_22614,N_22094);
nor U23205 (N_23205,N_22341,N_22111);
xnor U23206 (N_23206,N_22179,N_22200);
nor U23207 (N_23207,N_22748,N_22731);
and U23208 (N_23208,N_22655,N_22042);
nand U23209 (N_23209,N_22501,N_22101);
nor U23210 (N_23210,N_22851,N_22161);
nor U23211 (N_23211,N_22766,N_22509);
or U23212 (N_23212,N_22270,N_22060);
and U23213 (N_23213,N_22336,N_22881);
xnor U23214 (N_23214,N_22662,N_22044);
and U23215 (N_23215,N_22989,N_22996);
nor U23216 (N_23216,N_22180,N_22271);
xor U23217 (N_23217,N_22273,N_22824);
and U23218 (N_23218,N_22343,N_22641);
or U23219 (N_23219,N_22131,N_22351);
xor U23220 (N_23220,N_22066,N_22144);
and U23221 (N_23221,N_22337,N_22059);
xor U23222 (N_23222,N_22043,N_22204);
or U23223 (N_23223,N_22941,N_22221);
and U23224 (N_23224,N_22023,N_22891);
or U23225 (N_23225,N_22105,N_22535);
and U23226 (N_23226,N_22753,N_22175);
xnor U23227 (N_23227,N_22342,N_22817);
nor U23228 (N_23228,N_22513,N_22815);
xnor U23229 (N_23229,N_22939,N_22296);
nor U23230 (N_23230,N_22421,N_22688);
xnor U23231 (N_23231,N_22772,N_22550);
nand U23232 (N_23232,N_22260,N_22075);
and U23233 (N_23233,N_22943,N_22449);
nand U23234 (N_23234,N_22581,N_22198);
and U23235 (N_23235,N_22285,N_22250);
and U23236 (N_23236,N_22622,N_22917);
nor U23237 (N_23237,N_22430,N_22357);
xnor U23238 (N_23238,N_22718,N_22991);
nor U23239 (N_23239,N_22104,N_22249);
nor U23240 (N_23240,N_22426,N_22942);
nor U23241 (N_23241,N_22681,N_22532);
or U23242 (N_23242,N_22811,N_22143);
and U23243 (N_23243,N_22605,N_22364);
or U23244 (N_23244,N_22330,N_22067);
nor U23245 (N_23245,N_22828,N_22822);
and U23246 (N_23246,N_22845,N_22734);
or U23247 (N_23247,N_22604,N_22908);
or U23248 (N_23248,N_22418,N_22548);
and U23249 (N_23249,N_22118,N_22207);
nor U23250 (N_23250,N_22005,N_22740);
nand U23251 (N_23251,N_22840,N_22170);
and U23252 (N_23252,N_22862,N_22450);
nor U23253 (N_23253,N_22970,N_22108);
or U23254 (N_23254,N_22778,N_22808);
nor U23255 (N_23255,N_22860,N_22839);
and U23256 (N_23256,N_22164,N_22412);
nor U23257 (N_23257,N_22018,N_22916);
xor U23258 (N_23258,N_22058,N_22761);
nand U23259 (N_23259,N_22793,N_22004);
nor U23260 (N_23260,N_22424,N_22189);
nor U23261 (N_23261,N_22595,N_22706);
nor U23262 (N_23262,N_22659,N_22099);
and U23263 (N_23263,N_22782,N_22582);
xnor U23264 (N_23264,N_22348,N_22910);
nor U23265 (N_23265,N_22028,N_22048);
and U23266 (N_23266,N_22562,N_22209);
xnor U23267 (N_23267,N_22196,N_22002);
and U23268 (N_23268,N_22030,N_22846);
and U23269 (N_23269,N_22812,N_22797);
xor U23270 (N_23270,N_22304,N_22445);
nand U23271 (N_23271,N_22819,N_22559);
or U23272 (N_23272,N_22757,N_22153);
and U23273 (N_23273,N_22855,N_22022);
or U23274 (N_23274,N_22477,N_22244);
nand U23275 (N_23275,N_22032,N_22963);
and U23276 (N_23276,N_22776,N_22522);
or U23277 (N_23277,N_22505,N_22016);
and U23278 (N_23278,N_22015,N_22405);
nor U23279 (N_23279,N_22820,N_22425);
xor U23280 (N_23280,N_22583,N_22038);
nand U23281 (N_23281,N_22729,N_22749);
nand U23282 (N_23282,N_22055,N_22987);
nor U23283 (N_23283,N_22918,N_22272);
and U23284 (N_23284,N_22438,N_22620);
nor U23285 (N_23285,N_22683,N_22354);
and U23286 (N_23286,N_22971,N_22564);
xnor U23287 (N_23287,N_22791,N_22301);
nor U23288 (N_23288,N_22951,N_22593);
and U23289 (N_23289,N_22636,N_22013);
nor U23290 (N_23290,N_22523,N_22525);
and U23291 (N_23291,N_22663,N_22809);
nand U23292 (N_23292,N_22399,N_22106);
xnor U23293 (N_23293,N_22463,N_22166);
or U23294 (N_23294,N_22312,N_22938);
and U23295 (N_23295,N_22353,N_22400);
xnor U23296 (N_23296,N_22654,N_22441);
xnor U23297 (N_23297,N_22465,N_22057);
and U23298 (N_23298,N_22361,N_22849);
and U23299 (N_23299,N_22162,N_22006);
and U23300 (N_23300,N_22247,N_22642);
nor U23301 (N_23301,N_22660,N_22458);
and U23302 (N_23302,N_22034,N_22154);
or U23303 (N_23303,N_22122,N_22638);
nor U23304 (N_23304,N_22545,N_22151);
xor U23305 (N_23305,N_22764,N_22508);
xor U23306 (N_23306,N_22183,N_22892);
nand U23307 (N_23307,N_22024,N_22100);
or U23308 (N_23308,N_22349,N_22589);
or U23309 (N_23309,N_22743,N_22069);
nand U23310 (N_23310,N_22818,N_22459);
or U23311 (N_23311,N_22844,N_22585);
xor U23312 (N_23312,N_22406,N_22159);
or U23313 (N_23313,N_22884,N_22201);
xnor U23314 (N_23314,N_22658,N_22362);
and U23315 (N_23315,N_22292,N_22964);
and U23316 (N_23316,N_22374,N_22911);
xnor U23317 (N_23317,N_22524,N_22552);
and U23318 (N_23318,N_22009,N_22618);
xor U23319 (N_23319,N_22710,N_22267);
and U23320 (N_23320,N_22573,N_22217);
or U23321 (N_23321,N_22752,N_22551);
nor U23322 (N_23322,N_22877,N_22256);
nand U23323 (N_23323,N_22279,N_22921);
or U23324 (N_23324,N_22632,N_22191);
nand U23325 (N_23325,N_22965,N_22813);
nand U23326 (N_23326,N_22314,N_22530);
or U23327 (N_23327,N_22739,N_22579);
xor U23328 (N_23328,N_22711,N_22637);
and U23329 (N_23329,N_22685,N_22537);
and U23330 (N_23330,N_22502,N_22156);
or U23331 (N_23331,N_22000,N_22158);
and U23332 (N_23332,N_22794,N_22543);
and U23333 (N_23333,N_22741,N_22453);
nand U23334 (N_23334,N_22553,N_22588);
xnor U23335 (N_23335,N_22977,N_22859);
nor U23336 (N_23336,N_22673,N_22223);
nand U23337 (N_23337,N_22765,N_22699);
and U23338 (N_23338,N_22021,N_22169);
nand U23339 (N_23339,N_22358,N_22694);
nor U23340 (N_23340,N_22226,N_22128);
nor U23341 (N_23341,N_22222,N_22386);
or U23342 (N_23342,N_22863,N_22275);
nand U23343 (N_23343,N_22019,N_22736);
nor U23344 (N_23344,N_22310,N_22300);
nand U23345 (N_23345,N_22712,N_22299);
nor U23346 (N_23346,N_22070,N_22510);
nand U23347 (N_23347,N_22258,N_22903);
and U23348 (N_23348,N_22136,N_22848);
and U23349 (N_23349,N_22225,N_22790);
nor U23350 (N_23350,N_22705,N_22407);
nand U23351 (N_23351,N_22570,N_22135);
xor U23352 (N_23352,N_22461,N_22653);
or U23353 (N_23353,N_22626,N_22380);
nand U23354 (N_23354,N_22611,N_22842);
or U23355 (N_23355,N_22228,N_22878);
nand U23356 (N_23356,N_22755,N_22246);
xnor U23357 (N_23357,N_22777,N_22081);
xnor U23358 (N_23358,N_22475,N_22051);
nand U23359 (N_23359,N_22331,N_22252);
nand U23360 (N_23360,N_22397,N_22437);
nor U23361 (N_23361,N_22253,N_22870);
and U23362 (N_23362,N_22227,N_22961);
and U23363 (N_23363,N_22930,N_22756);
nor U23364 (N_23364,N_22968,N_22025);
xor U23365 (N_23365,N_22893,N_22677);
nand U23366 (N_23366,N_22856,N_22902);
xor U23367 (N_23367,N_22090,N_22346);
nand U23368 (N_23368,N_22033,N_22433);
nor U23369 (N_23369,N_22255,N_22997);
xnor U23370 (N_23370,N_22633,N_22174);
nor U23371 (N_23371,N_22195,N_22920);
and U23372 (N_23372,N_22959,N_22531);
nand U23373 (N_23373,N_22760,N_22586);
xor U23374 (N_23374,N_22606,N_22491);
or U23375 (N_23375,N_22155,N_22643);
nor U23376 (N_23376,N_22213,N_22889);
and U23377 (N_23377,N_22803,N_22590);
nor U23378 (N_23378,N_22283,N_22919);
or U23379 (N_23379,N_22576,N_22713);
nand U23380 (N_23380,N_22029,N_22215);
xnor U23381 (N_23381,N_22308,N_22120);
or U23382 (N_23382,N_22980,N_22079);
nand U23383 (N_23383,N_22053,N_22528);
and U23384 (N_23384,N_22628,N_22113);
and U23385 (N_23385,N_22110,N_22202);
and U23386 (N_23386,N_22214,N_22624);
xnor U23387 (N_23387,N_22792,N_22112);
nor U23388 (N_23388,N_22366,N_22867);
nor U23389 (N_23389,N_22547,N_22427);
or U23390 (N_23390,N_22935,N_22690);
and U23391 (N_23391,N_22394,N_22187);
nor U23392 (N_23392,N_22841,N_22515);
nand U23393 (N_23393,N_22334,N_22746);
and U23394 (N_23394,N_22446,N_22148);
nor U23395 (N_23395,N_22945,N_22701);
xnor U23396 (N_23396,N_22488,N_22974);
or U23397 (N_23397,N_22503,N_22291);
or U23398 (N_23398,N_22512,N_22592);
and U23399 (N_23399,N_22321,N_22875);
xor U23400 (N_23400,N_22259,N_22415);
or U23401 (N_23401,N_22647,N_22826);
xnor U23402 (N_23402,N_22489,N_22682);
or U23403 (N_23403,N_22995,N_22298);
and U23404 (N_23404,N_22388,N_22439);
xor U23405 (N_23405,N_22498,N_22327);
xnor U23406 (N_23406,N_22575,N_22580);
or U23407 (N_23407,N_22235,N_22482);
nand U23408 (N_23408,N_22184,N_22897);
or U23409 (N_23409,N_22318,N_22619);
xnor U23410 (N_23410,N_22322,N_22176);
or U23411 (N_23411,N_22390,N_22771);
nor U23412 (N_23412,N_22763,N_22123);
or U23413 (N_23413,N_22208,N_22584);
or U23414 (N_23414,N_22497,N_22953);
nor U23415 (N_23415,N_22008,N_22829);
nand U23416 (N_23416,N_22831,N_22962);
nor U23417 (N_23417,N_22779,N_22904);
nand U23418 (N_23418,N_22567,N_22806);
or U23419 (N_23419,N_22403,N_22172);
nand U23420 (N_23420,N_22807,N_22157);
or U23421 (N_23421,N_22393,N_22768);
nor U23422 (N_23422,N_22609,N_22572);
nor U23423 (N_23423,N_22186,N_22519);
nor U23424 (N_23424,N_22185,N_22315);
nand U23425 (N_23425,N_22635,N_22861);
and U23426 (N_23426,N_22173,N_22775);
nand U23427 (N_23427,N_22152,N_22077);
nand U23428 (N_23428,N_22954,N_22280);
and U23429 (N_23429,N_22370,N_22541);
and U23430 (N_23430,N_22007,N_22056);
nand U23431 (N_23431,N_22027,N_22276);
and U23432 (N_23432,N_22999,N_22696);
nand U23433 (N_23433,N_22243,N_22966);
or U23434 (N_23434,N_22416,N_22832);
nand U23435 (N_23435,N_22709,N_22896);
or U23436 (N_23436,N_22378,N_22504);
or U23437 (N_23437,N_22473,N_22948);
or U23438 (N_23438,N_22958,N_22320);
xor U23439 (N_23439,N_22657,N_22192);
nor U23440 (N_23440,N_22237,N_22141);
nor U23441 (N_23441,N_22045,N_22847);
xnor U23442 (N_23442,N_22816,N_22265);
nand U23443 (N_23443,N_22931,N_22957);
and U23444 (N_23444,N_22251,N_22979);
xor U23445 (N_23445,N_22466,N_22139);
xor U23446 (N_23446,N_22432,N_22389);
or U23447 (N_23447,N_22927,N_22517);
nand U23448 (N_23448,N_22317,N_22774);
xnor U23449 (N_23449,N_22360,N_22722);
and U23450 (N_23450,N_22750,N_22001);
and U23451 (N_23451,N_22046,N_22474);
nand U23452 (N_23452,N_22383,N_22872);
and U23453 (N_23453,N_22783,N_22857);
nor U23454 (N_23454,N_22423,N_22704);
xor U23455 (N_23455,N_22313,N_22679);
and U23456 (N_23456,N_22444,N_22899);
nor U23457 (N_23457,N_22181,N_22596);
xnor U23458 (N_23458,N_22598,N_22571);
or U23459 (N_23459,N_22411,N_22738);
xor U23460 (N_23460,N_22396,N_22344);
nor U23461 (N_23461,N_22302,N_22086);
xnor U23462 (N_23462,N_22940,N_22305);
or U23463 (N_23463,N_22481,N_22480);
and U23464 (N_23464,N_22728,N_22759);
or U23465 (N_23465,N_22577,N_22880);
xnor U23466 (N_23466,N_22231,N_22926);
nor U23467 (N_23467,N_22124,N_22188);
nand U23468 (N_23468,N_22117,N_22901);
nand U23469 (N_23469,N_22134,N_22879);
and U23470 (N_23470,N_22984,N_22316);
xnor U23471 (N_23471,N_22607,N_22858);
nand U23472 (N_23472,N_22137,N_22464);
or U23473 (N_23473,N_22602,N_22992);
or U23474 (N_23474,N_22010,N_22163);
nor U23475 (N_23475,N_22254,N_22074);
nor U23476 (N_23476,N_22725,N_22613);
or U23477 (N_23477,N_22796,N_22012);
and U23478 (N_23478,N_22976,N_22949);
or U23479 (N_23479,N_22670,N_22898);
and U23480 (N_23480,N_22563,N_22751);
xor U23481 (N_23481,N_22499,N_22691);
nand U23482 (N_23482,N_22715,N_22608);
and U23483 (N_23483,N_22780,N_22936);
nand U23484 (N_23484,N_22230,N_22700);
xor U23485 (N_23485,N_22982,N_22758);
or U23486 (N_23486,N_22527,N_22800);
nor U23487 (N_23487,N_22591,N_22555);
nand U23488 (N_23488,N_22182,N_22303);
nor U23489 (N_23489,N_22147,N_22823);
nor U23490 (N_23490,N_22119,N_22789);
nand U23491 (N_23491,N_22414,N_22199);
or U23492 (N_23492,N_22843,N_22103);
nor U23493 (N_23493,N_22621,N_22040);
nand U23494 (N_23494,N_22558,N_22717);
nand U23495 (N_23495,N_22865,N_22076);
or U23496 (N_23496,N_22496,N_22261);
and U23497 (N_23497,N_22160,N_22913);
nand U23498 (N_23498,N_22640,N_22085);
or U23499 (N_23499,N_22359,N_22288);
nor U23500 (N_23500,N_22048,N_22162);
nand U23501 (N_23501,N_22287,N_22134);
nand U23502 (N_23502,N_22501,N_22165);
and U23503 (N_23503,N_22393,N_22373);
and U23504 (N_23504,N_22174,N_22884);
or U23505 (N_23505,N_22287,N_22923);
nand U23506 (N_23506,N_22868,N_22553);
nor U23507 (N_23507,N_22355,N_22139);
nand U23508 (N_23508,N_22721,N_22151);
xnor U23509 (N_23509,N_22310,N_22185);
nand U23510 (N_23510,N_22002,N_22997);
and U23511 (N_23511,N_22082,N_22230);
or U23512 (N_23512,N_22966,N_22236);
or U23513 (N_23513,N_22696,N_22737);
or U23514 (N_23514,N_22094,N_22634);
nand U23515 (N_23515,N_22049,N_22502);
or U23516 (N_23516,N_22615,N_22863);
and U23517 (N_23517,N_22595,N_22412);
nor U23518 (N_23518,N_22776,N_22624);
and U23519 (N_23519,N_22453,N_22782);
nand U23520 (N_23520,N_22331,N_22038);
and U23521 (N_23521,N_22946,N_22484);
nand U23522 (N_23522,N_22387,N_22809);
nand U23523 (N_23523,N_22797,N_22576);
and U23524 (N_23524,N_22598,N_22647);
xor U23525 (N_23525,N_22783,N_22488);
and U23526 (N_23526,N_22389,N_22753);
nor U23527 (N_23527,N_22718,N_22153);
or U23528 (N_23528,N_22274,N_22237);
nor U23529 (N_23529,N_22170,N_22278);
nand U23530 (N_23530,N_22312,N_22319);
and U23531 (N_23531,N_22384,N_22230);
and U23532 (N_23532,N_22239,N_22883);
nand U23533 (N_23533,N_22912,N_22991);
nor U23534 (N_23534,N_22224,N_22987);
nand U23535 (N_23535,N_22884,N_22701);
or U23536 (N_23536,N_22458,N_22891);
nor U23537 (N_23537,N_22478,N_22465);
xnor U23538 (N_23538,N_22336,N_22424);
xnor U23539 (N_23539,N_22311,N_22602);
and U23540 (N_23540,N_22436,N_22693);
nand U23541 (N_23541,N_22168,N_22616);
or U23542 (N_23542,N_22495,N_22210);
xor U23543 (N_23543,N_22504,N_22864);
nand U23544 (N_23544,N_22987,N_22875);
xor U23545 (N_23545,N_22870,N_22675);
nand U23546 (N_23546,N_22049,N_22098);
and U23547 (N_23547,N_22869,N_22513);
xnor U23548 (N_23548,N_22510,N_22315);
xor U23549 (N_23549,N_22298,N_22091);
or U23550 (N_23550,N_22019,N_22087);
and U23551 (N_23551,N_22951,N_22809);
and U23552 (N_23552,N_22499,N_22060);
nor U23553 (N_23553,N_22903,N_22496);
nand U23554 (N_23554,N_22392,N_22865);
xor U23555 (N_23555,N_22225,N_22035);
nor U23556 (N_23556,N_22754,N_22171);
or U23557 (N_23557,N_22457,N_22558);
nor U23558 (N_23558,N_22157,N_22574);
nand U23559 (N_23559,N_22211,N_22317);
and U23560 (N_23560,N_22229,N_22512);
and U23561 (N_23561,N_22622,N_22174);
or U23562 (N_23562,N_22680,N_22475);
or U23563 (N_23563,N_22650,N_22003);
nor U23564 (N_23564,N_22221,N_22894);
nand U23565 (N_23565,N_22550,N_22411);
or U23566 (N_23566,N_22371,N_22216);
nand U23567 (N_23567,N_22436,N_22141);
xor U23568 (N_23568,N_22290,N_22753);
xnor U23569 (N_23569,N_22338,N_22113);
xnor U23570 (N_23570,N_22047,N_22858);
or U23571 (N_23571,N_22791,N_22699);
xor U23572 (N_23572,N_22005,N_22045);
xnor U23573 (N_23573,N_22497,N_22745);
or U23574 (N_23574,N_22995,N_22178);
xnor U23575 (N_23575,N_22167,N_22347);
nand U23576 (N_23576,N_22094,N_22957);
xor U23577 (N_23577,N_22825,N_22554);
nand U23578 (N_23578,N_22728,N_22975);
or U23579 (N_23579,N_22774,N_22283);
xor U23580 (N_23580,N_22827,N_22507);
or U23581 (N_23581,N_22866,N_22225);
or U23582 (N_23582,N_22019,N_22316);
nand U23583 (N_23583,N_22989,N_22203);
nand U23584 (N_23584,N_22936,N_22921);
and U23585 (N_23585,N_22715,N_22041);
nor U23586 (N_23586,N_22174,N_22641);
nand U23587 (N_23587,N_22499,N_22686);
nor U23588 (N_23588,N_22484,N_22808);
and U23589 (N_23589,N_22234,N_22076);
nor U23590 (N_23590,N_22454,N_22776);
or U23591 (N_23591,N_22285,N_22692);
nor U23592 (N_23592,N_22827,N_22034);
nor U23593 (N_23593,N_22599,N_22689);
and U23594 (N_23594,N_22658,N_22185);
nand U23595 (N_23595,N_22991,N_22290);
nand U23596 (N_23596,N_22179,N_22486);
xor U23597 (N_23597,N_22606,N_22003);
nor U23598 (N_23598,N_22208,N_22514);
nand U23599 (N_23599,N_22945,N_22743);
and U23600 (N_23600,N_22345,N_22910);
nor U23601 (N_23601,N_22037,N_22944);
xor U23602 (N_23602,N_22322,N_22631);
or U23603 (N_23603,N_22386,N_22401);
xnor U23604 (N_23604,N_22016,N_22919);
xor U23605 (N_23605,N_22732,N_22603);
nand U23606 (N_23606,N_22218,N_22938);
xor U23607 (N_23607,N_22535,N_22459);
or U23608 (N_23608,N_22355,N_22974);
nor U23609 (N_23609,N_22519,N_22310);
nor U23610 (N_23610,N_22168,N_22486);
and U23611 (N_23611,N_22078,N_22358);
nand U23612 (N_23612,N_22657,N_22253);
nand U23613 (N_23613,N_22384,N_22321);
and U23614 (N_23614,N_22334,N_22612);
nor U23615 (N_23615,N_22663,N_22892);
or U23616 (N_23616,N_22542,N_22475);
nor U23617 (N_23617,N_22092,N_22969);
and U23618 (N_23618,N_22983,N_22961);
or U23619 (N_23619,N_22886,N_22607);
xnor U23620 (N_23620,N_22264,N_22848);
nor U23621 (N_23621,N_22758,N_22172);
xnor U23622 (N_23622,N_22867,N_22517);
or U23623 (N_23623,N_22935,N_22305);
xnor U23624 (N_23624,N_22705,N_22002);
or U23625 (N_23625,N_22186,N_22280);
nand U23626 (N_23626,N_22255,N_22094);
xor U23627 (N_23627,N_22859,N_22663);
nand U23628 (N_23628,N_22007,N_22173);
xnor U23629 (N_23629,N_22137,N_22693);
nand U23630 (N_23630,N_22683,N_22321);
xnor U23631 (N_23631,N_22284,N_22890);
nor U23632 (N_23632,N_22601,N_22911);
xor U23633 (N_23633,N_22756,N_22353);
or U23634 (N_23634,N_22671,N_22692);
nand U23635 (N_23635,N_22579,N_22218);
nor U23636 (N_23636,N_22933,N_22141);
and U23637 (N_23637,N_22397,N_22664);
or U23638 (N_23638,N_22222,N_22961);
nand U23639 (N_23639,N_22755,N_22971);
and U23640 (N_23640,N_22906,N_22915);
and U23641 (N_23641,N_22448,N_22086);
nor U23642 (N_23642,N_22591,N_22089);
or U23643 (N_23643,N_22300,N_22609);
nand U23644 (N_23644,N_22988,N_22066);
nor U23645 (N_23645,N_22418,N_22454);
nand U23646 (N_23646,N_22182,N_22916);
or U23647 (N_23647,N_22581,N_22747);
nor U23648 (N_23648,N_22229,N_22343);
and U23649 (N_23649,N_22202,N_22995);
and U23650 (N_23650,N_22933,N_22882);
nor U23651 (N_23651,N_22268,N_22684);
nand U23652 (N_23652,N_22746,N_22974);
nand U23653 (N_23653,N_22250,N_22600);
nand U23654 (N_23654,N_22172,N_22064);
and U23655 (N_23655,N_22194,N_22363);
nand U23656 (N_23656,N_22401,N_22919);
xor U23657 (N_23657,N_22791,N_22384);
and U23658 (N_23658,N_22102,N_22075);
xnor U23659 (N_23659,N_22329,N_22522);
nor U23660 (N_23660,N_22298,N_22424);
or U23661 (N_23661,N_22264,N_22136);
nor U23662 (N_23662,N_22875,N_22609);
nand U23663 (N_23663,N_22908,N_22096);
or U23664 (N_23664,N_22943,N_22243);
and U23665 (N_23665,N_22199,N_22191);
nor U23666 (N_23666,N_22294,N_22622);
or U23667 (N_23667,N_22672,N_22746);
or U23668 (N_23668,N_22136,N_22352);
xor U23669 (N_23669,N_22429,N_22777);
or U23670 (N_23670,N_22812,N_22109);
nor U23671 (N_23671,N_22871,N_22307);
nor U23672 (N_23672,N_22702,N_22373);
or U23673 (N_23673,N_22042,N_22937);
or U23674 (N_23674,N_22764,N_22046);
nand U23675 (N_23675,N_22658,N_22541);
xor U23676 (N_23676,N_22230,N_22678);
and U23677 (N_23677,N_22431,N_22685);
and U23678 (N_23678,N_22329,N_22603);
or U23679 (N_23679,N_22832,N_22432);
nand U23680 (N_23680,N_22111,N_22200);
nand U23681 (N_23681,N_22986,N_22650);
xnor U23682 (N_23682,N_22984,N_22311);
and U23683 (N_23683,N_22675,N_22699);
and U23684 (N_23684,N_22856,N_22493);
nor U23685 (N_23685,N_22148,N_22383);
nand U23686 (N_23686,N_22004,N_22086);
and U23687 (N_23687,N_22738,N_22218);
nor U23688 (N_23688,N_22662,N_22434);
and U23689 (N_23689,N_22054,N_22622);
xor U23690 (N_23690,N_22813,N_22899);
nand U23691 (N_23691,N_22001,N_22517);
nor U23692 (N_23692,N_22921,N_22741);
and U23693 (N_23693,N_22577,N_22223);
or U23694 (N_23694,N_22094,N_22620);
nor U23695 (N_23695,N_22642,N_22981);
or U23696 (N_23696,N_22102,N_22738);
nand U23697 (N_23697,N_22985,N_22662);
nand U23698 (N_23698,N_22076,N_22411);
and U23699 (N_23699,N_22943,N_22009);
or U23700 (N_23700,N_22260,N_22925);
nand U23701 (N_23701,N_22977,N_22193);
nand U23702 (N_23702,N_22712,N_22498);
and U23703 (N_23703,N_22222,N_22428);
or U23704 (N_23704,N_22713,N_22366);
nor U23705 (N_23705,N_22564,N_22490);
and U23706 (N_23706,N_22939,N_22256);
or U23707 (N_23707,N_22298,N_22099);
and U23708 (N_23708,N_22495,N_22613);
or U23709 (N_23709,N_22048,N_22783);
or U23710 (N_23710,N_22635,N_22539);
and U23711 (N_23711,N_22737,N_22214);
nor U23712 (N_23712,N_22003,N_22740);
xor U23713 (N_23713,N_22055,N_22464);
nand U23714 (N_23714,N_22457,N_22416);
xor U23715 (N_23715,N_22428,N_22520);
or U23716 (N_23716,N_22885,N_22869);
nand U23717 (N_23717,N_22123,N_22134);
xor U23718 (N_23718,N_22145,N_22774);
nand U23719 (N_23719,N_22271,N_22607);
or U23720 (N_23720,N_22729,N_22407);
nand U23721 (N_23721,N_22522,N_22960);
xnor U23722 (N_23722,N_22632,N_22988);
xor U23723 (N_23723,N_22925,N_22298);
and U23724 (N_23724,N_22144,N_22534);
nand U23725 (N_23725,N_22934,N_22872);
nand U23726 (N_23726,N_22269,N_22417);
nor U23727 (N_23727,N_22501,N_22665);
xnor U23728 (N_23728,N_22173,N_22461);
nor U23729 (N_23729,N_22495,N_22075);
and U23730 (N_23730,N_22668,N_22119);
and U23731 (N_23731,N_22674,N_22685);
nand U23732 (N_23732,N_22912,N_22249);
or U23733 (N_23733,N_22526,N_22592);
nand U23734 (N_23734,N_22748,N_22151);
or U23735 (N_23735,N_22061,N_22016);
nand U23736 (N_23736,N_22866,N_22813);
xnor U23737 (N_23737,N_22443,N_22303);
or U23738 (N_23738,N_22707,N_22157);
xor U23739 (N_23739,N_22781,N_22149);
or U23740 (N_23740,N_22355,N_22814);
or U23741 (N_23741,N_22669,N_22018);
and U23742 (N_23742,N_22232,N_22179);
nor U23743 (N_23743,N_22122,N_22688);
nor U23744 (N_23744,N_22559,N_22885);
xnor U23745 (N_23745,N_22325,N_22910);
and U23746 (N_23746,N_22215,N_22062);
xnor U23747 (N_23747,N_22494,N_22650);
or U23748 (N_23748,N_22294,N_22631);
xor U23749 (N_23749,N_22910,N_22112);
and U23750 (N_23750,N_22705,N_22970);
nor U23751 (N_23751,N_22022,N_22697);
xnor U23752 (N_23752,N_22558,N_22797);
xnor U23753 (N_23753,N_22197,N_22368);
and U23754 (N_23754,N_22020,N_22414);
nor U23755 (N_23755,N_22595,N_22744);
nand U23756 (N_23756,N_22672,N_22242);
nor U23757 (N_23757,N_22659,N_22527);
and U23758 (N_23758,N_22918,N_22859);
nand U23759 (N_23759,N_22251,N_22688);
nand U23760 (N_23760,N_22527,N_22567);
nor U23761 (N_23761,N_22798,N_22738);
xnor U23762 (N_23762,N_22564,N_22297);
and U23763 (N_23763,N_22909,N_22151);
or U23764 (N_23764,N_22512,N_22812);
nand U23765 (N_23765,N_22805,N_22528);
and U23766 (N_23766,N_22023,N_22765);
xor U23767 (N_23767,N_22445,N_22983);
xnor U23768 (N_23768,N_22131,N_22224);
nor U23769 (N_23769,N_22097,N_22588);
or U23770 (N_23770,N_22731,N_22412);
nor U23771 (N_23771,N_22730,N_22242);
nor U23772 (N_23772,N_22418,N_22926);
nor U23773 (N_23773,N_22757,N_22552);
and U23774 (N_23774,N_22226,N_22905);
or U23775 (N_23775,N_22434,N_22125);
or U23776 (N_23776,N_22587,N_22403);
nor U23777 (N_23777,N_22583,N_22096);
xnor U23778 (N_23778,N_22506,N_22737);
or U23779 (N_23779,N_22431,N_22074);
or U23780 (N_23780,N_22949,N_22848);
nor U23781 (N_23781,N_22116,N_22344);
and U23782 (N_23782,N_22506,N_22077);
or U23783 (N_23783,N_22929,N_22343);
and U23784 (N_23784,N_22119,N_22757);
nor U23785 (N_23785,N_22274,N_22084);
or U23786 (N_23786,N_22335,N_22956);
or U23787 (N_23787,N_22249,N_22819);
and U23788 (N_23788,N_22454,N_22953);
nor U23789 (N_23789,N_22386,N_22103);
nor U23790 (N_23790,N_22914,N_22104);
nor U23791 (N_23791,N_22605,N_22207);
and U23792 (N_23792,N_22626,N_22883);
nand U23793 (N_23793,N_22821,N_22200);
and U23794 (N_23794,N_22717,N_22071);
xnor U23795 (N_23795,N_22704,N_22366);
and U23796 (N_23796,N_22797,N_22111);
nor U23797 (N_23797,N_22782,N_22668);
nand U23798 (N_23798,N_22304,N_22477);
or U23799 (N_23799,N_22792,N_22002);
or U23800 (N_23800,N_22354,N_22820);
xor U23801 (N_23801,N_22744,N_22807);
xnor U23802 (N_23802,N_22687,N_22903);
and U23803 (N_23803,N_22827,N_22428);
and U23804 (N_23804,N_22462,N_22078);
or U23805 (N_23805,N_22796,N_22006);
nor U23806 (N_23806,N_22783,N_22328);
xor U23807 (N_23807,N_22468,N_22895);
nand U23808 (N_23808,N_22379,N_22389);
xor U23809 (N_23809,N_22202,N_22657);
and U23810 (N_23810,N_22030,N_22416);
nor U23811 (N_23811,N_22028,N_22536);
nand U23812 (N_23812,N_22610,N_22882);
nand U23813 (N_23813,N_22642,N_22131);
xor U23814 (N_23814,N_22716,N_22640);
nor U23815 (N_23815,N_22785,N_22896);
xnor U23816 (N_23816,N_22368,N_22927);
nor U23817 (N_23817,N_22341,N_22035);
xor U23818 (N_23818,N_22043,N_22873);
nor U23819 (N_23819,N_22142,N_22839);
nor U23820 (N_23820,N_22776,N_22302);
and U23821 (N_23821,N_22530,N_22989);
or U23822 (N_23822,N_22015,N_22234);
and U23823 (N_23823,N_22688,N_22343);
xor U23824 (N_23824,N_22396,N_22209);
nand U23825 (N_23825,N_22944,N_22353);
or U23826 (N_23826,N_22670,N_22079);
nand U23827 (N_23827,N_22629,N_22057);
xnor U23828 (N_23828,N_22790,N_22274);
or U23829 (N_23829,N_22277,N_22395);
or U23830 (N_23830,N_22513,N_22278);
xor U23831 (N_23831,N_22187,N_22463);
nor U23832 (N_23832,N_22463,N_22749);
xor U23833 (N_23833,N_22451,N_22821);
xor U23834 (N_23834,N_22994,N_22839);
and U23835 (N_23835,N_22790,N_22027);
xor U23836 (N_23836,N_22520,N_22948);
nor U23837 (N_23837,N_22349,N_22973);
xor U23838 (N_23838,N_22341,N_22902);
nand U23839 (N_23839,N_22698,N_22767);
or U23840 (N_23840,N_22544,N_22260);
nand U23841 (N_23841,N_22954,N_22519);
nand U23842 (N_23842,N_22218,N_22897);
nor U23843 (N_23843,N_22664,N_22488);
nand U23844 (N_23844,N_22573,N_22652);
nand U23845 (N_23845,N_22279,N_22888);
nand U23846 (N_23846,N_22700,N_22638);
xor U23847 (N_23847,N_22735,N_22675);
or U23848 (N_23848,N_22973,N_22917);
xor U23849 (N_23849,N_22983,N_22198);
or U23850 (N_23850,N_22372,N_22896);
nor U23851 (N_23851,N_22984,N_22351);
or U23852 (N_23852,N_22793,N_22040);
nor U23853 (N_23853,N_22721,N_22198);
nand U23854 (N_23854,N_22424,N_22121);
nand U23855 (N_23855,N_22114,N_22218);
or U23856 (N_23856,N_22318,N_22425);
nand U23857 (N_23857,N_22951,N_22819);
nand U23858 (N_23858,N_22832,N_22344);
or U23859 (N_23859,N_22110,N_22597);
or U23860 (N_23860,N_22316,N_22113);
and U23861 (N_23861,N_22876,N_22233);
nor U23862 (N_23862,N_22779,N_22331);
or U23863 (N_23863,N_22562,N_22373);
nor U23864 (N_23864,N_22506,N_22216);
nand U23865 (N_23865,N_22215,N_22086);
and U23866 (N_23866,N_22114,N_22683);
or U23867 (N_23867,N_22697,N_22724);
nor U23868 (N_23868,N_22947,N_22792);
xnor U23869 (N_23869,N_22447,N_22543);
nor U23870 (N_23870,N_22597,N_22162);
xnor U23871 (N_23871,N_22988,N_22617);
nand U23872 (N_23872,N_22834,N_22844);
xor U23873 (N_23873,N_22920,N_22390);
nand U23874 (N_23874,N_22383,N_22065);
nor U23875 (N_23875,N_22489,N_22499);
or U23876 (N_23876,N_22409,N_22693);
xor U23877 (N_23877,N_22300,N_22007);
nor U23878 (N_23878,N_22287,N_22483);
nand U23879 (N_23879,N_22313,N_22424);
nand U23880 (N_23880,N_22944,N_22196);
nor U23881 (N_23881,N_22738,N_22348);
and U23882 (N_23882,N_22102,N_22154);
and U23883 (N_23883,N_22402,N_22638);
and U23884 (N_23884,N_22950,N_22378);
nand U23885 (N_23885,N_22071,N_22836);
nor U23886 (N_23886,N_22869,N_22020);
and U23887 (N_23887,N_22490,N_22988);
or U23888 (N_23888,N_22578,N_22335);
or U23889 (N_23889,N_22280,N_22733);
nor U23890 (N_23890,N_22743,N_22191);
nor U23891 (N_23891,N_22655,N_22498);
and U23892 (N_23892,N_22830,N_22618);
or U23893 (N_23893,N_22721,N_22227);
xor U23894 (N_23894,N_22272,N_22336);
nand U23895 (N_23895,N_22193,N_22292);
or U23896 (N_23896,N_22689,N_22050);
nand U23897 (N_23897,N_22611,N_22440);
nand U23898 (N_23898,N_22559,N_22066);
xnor U23899 (N_23899,N_22309,N_22829);
nand U23900 (N_23900,N_22310,N_22030);
and U23901 (N_23901,N_22740,N_22542);
nor U23902 (N_23902,N_22364,N_22609);
or U23903 (N_23903,N_22064,N_22723);
and U23904 (N_23904,N_22069,N_22232);
nor U23905 (N_23905,N_22889,N_22967);
and U23906 (N_23906,N_22631,N_22723);
nand U23907 (N_23907,N_22133,N_22672);
nand U23908 (N_23908,N_22715,N_22345);
nor U23909 (N_23909,N_22735,N_22952);
or U23910 (N_23910,N_22901,N_22899);
or U23911 (N_23911,N_22274,N_22737);
xnor U23912 (N_23912,N_22324,N_22711);
xor U23913 (N_23913,N_22618,N_22801);
and U23914 (N_23914,N_22036,N_22780);
and U23915 (N_23915,N_22157,N_22508);
or U23916 (N_23916,N_22722,N_22682);
xnor U23917 (N_23917,N_22137,N_22323);
or U23918 (N_23918,N_22673,N_22619);
and U23919 (N_23919,N_22377,N_22171);
or U23920 (N_23920,N_22797,N_22215);
xnor U23921 (N_23921,N_22139,N_22866);
or U23922 (N_23922,N_22035,N_22789);
nand U23923 (N_23923,N_22804,N_22642);
nand U23924 (N_23924,N_22522,N_22451);
nand U23925 (N_23925,N_22753,N_22065);
nand U23926 (N_23926,N_22673,N_22211);
xnor U23927 (N_23927,N_22941,N_22893);
xnor U23928 (N_23928,N_22064,N_22001);
or U23929 (N_23929,N_22274,N_22192);
and U23930 (N_23930,N_22515,N_22750);
or U23931 (N_23931,N_22757,N_22787);
nand U23932 (N_23932,N_22145,N_22180);
nor U23933 (N_23933,N_22264,N_22865);
and U23934 (N_23934,N_22211,N_22350);
nand U23935 (N_23935,N_22646,N_22390);
xnor U23936 (N_23936,N_22862,N_22495);
nand U23937 (N_23937,N_22997,N_22592);
nand U23938 (N_23938,N_22971,N_22862);
and U23939 (N_23939,N_22889,N_22227);
or U23940 (N_23940,N_22556,N_22031);
xnor U23941 (N_23941,N_22805,N_22331);
nor U23942 (N_23942,N_22742,N_22888);
or U23943 (N_23943,N_22791,N_22640);
and U23944 (N_23944,N_22367,N_22655);
nor U23945 (N_23945,N_22007,N_22567);
or U23946 (N_23946,N_22449,N_22714);
xnor U23947 (N_23947,N_22298,N_22360);
nor U23948 (N_23948,N_22486,N_22128);
nand U23949 (N_23949,N_22642,N_22639);
nand U23950 (N_23950,N_22516,N_22849);
nand U23951 (N_23951,N_22435,N_22710);
nand U23952 (N_23952,N_22034,N_22635);
nor U23953 (N_23953,N_22171,N_22526);
nand U23954 (N_23954,N_22581,N_22627);
nand U23955 (N_23955,N_22726,N_22432);
xnor U23956 (N_23956,N_22355,N_22605);
nor U23957 (N_23957,N_22074,N_22056);
xnor U23958 (N_23958,N_22136,N_22881);
nor U23959 (N_23959,N_22884,N_22569);
or U23960 (N_23960,N_22207,N_22259);
nor U23961 (N_23961,N_22553,N_22577);
nor U23962 (N_23962,N_22396,N_22177);
or U23963 (N_23963,N_22806,N_22124);
nor U23964 (N_23964,N_22534,N_22327);
xnor U23965 (N_23965,N_22285,N_22630);
nor U23966 (N_23966,N_22033,N_22582);
nor U23967 (N_23967,N_22468,N_22555);
and U23968 (N_23968,N_22746,N_22342);
and U23969 (N_23969,N_22498,N_22335);
and U23970 (N_23970,N_22643,N_22706);
or U23971 (N_23971,N_22093,N_22307);
nor U23972 (N_23972,N_22478,N_22190);
xnor U23973 (N_23973,N_22967,N_22416);
nand U23974 (N_23974,N_22894,N_22543);
nand U23975 (N_23975,N_22648,N_22978);
and U23976 (N_23976,N_22146,N_22626);
nand U23977 (N_23977,N_22659,N_22883);
nor U23978 (N_23978,N_22186,N_22241);
xnor U23979 (N_23979,N_22442,N_22678);
xor U23980 (N_23980,N_22278,N_22413);
or U23981 (N_23981,N_22745,N_22990);
xor U23982 (N_23982,N_22178,N_22143);
xor U23983 (N_23983,N_22533,N_22380);
nand U23984 (N_23984,N_22988,N_22580);
or U23985 (N_23985,N_22232,N_22620);
or U23986 (N_23986,N_22317,N_22653);
and U23987 (N_23987,N_22247,N_22105);
xor U23988 (N_23988,N_22536,N_22905);
nor U23989 (N_23989,N_22175,N_22147);
and U23990 (N_23990,N_22834,N_22195);
xnor U23991 (N_23991,N_22877,N_22913);
or U23992 (N_23992,N_22438,N_22233);
or U23993 (N_23993,N_22791,N_22823);
xor U23994 (N_23994,N_22858,N_22250);
and U23995 (N_23995,N_22743,N_22375);
xor U23996 (N_23996,N_22402,N_22213);
nor U23997 (N_23997,N_22698,N_22131);
and U23998 (N_23998,N_22031,N_22796);
and U23999 (N_23999,N_22393,N_22784);
or U24000 (N_24000,N_23546,N_23469);
nand U24001 (N_24001,N_23760,N_23033);
nor U24002 (N_24002,N_23341,N_23733);
and U24003 (N_24003,N_23648,N_23309);
xnor U24004 (N_24004,N_23856,N_23406);
nor U24005 (N_24005,N_23574,N_23378);
nand U24006 (N_24006,N_23670,N_23553);
xor U24007 (N_24007,N_23799,N_23485);
nand U24008 (N_24008,N_23071,N_23305);
or U24009 (N_24009,N_23468,N_23295);
or U24010 (N_24010,N_23519,N_23885);
nor U24011 (N_24011,N_23112,N_23391);
or U24012 (N_24012,N_23579,N_23690);
or U24013 (N_24013,N_23296,N_23915);
and U24014 (N_24014,N_23820,N_23607);
or U24015 (N_24015,N_23286,N_23601);
or U24016 (N_24016,N_23830,N_23695);
nand U24017 (N_24017,N_23409,N_23746);
xor U24018 (N_24018,N_23421,N_23793);
nand U24019 (N_24019,N_23169,N_23490);
and U24020 (N_24020,N_23496,N_23012);
xor U24021 (N_24021,N_23004,N_23124);
xor U24022 (N_24022,N_23927,N_23275);
or U24023 (N_24023,N_23541,N_23942);
nor U24024 (N_24024,N_23470,N_23527);
nor U24025 (N_24025,N_23375,N_23896);
xnor U24026 (N_24026,N_23214,N_23351);
nand U24027 (N_24027,N_23843,N_23879);
and U24028 (N_24028,N_23552,N_23499);
nand U24029 (N_24029,N_23431,N_23997);
xor U24030 (N_24030,N_23453,N_23903);
or U24031 (N_24031,N_23940,N_23741);
nor U24032 (N_24032,N_23443,N_23430);
xnor U24033 (N_24033,N_23835,N_23037);
or U24034 (N_24034,N_23845,N_23855);
and U24035 (N_24035,N_23818,N_23397);
and U24036 (N_24036,N_23560,N_23795);
and U24037 (N_24037,N_23102,N_23403);
or U24038 (N_24038,N_23866,N_23376);
xnor U24039 (N_24039,N_23256,N_23252);
and U24040 (N_24040,N_23266,N_23123);
xnor U24041 (N_24041,N_23304,N_23639);
nand U24042 (N_24042,N_23128,N_23543);
nor U24043 (N_24043,N_23762,N_23192);
and U24044 (N_24044,N_23901,N_23941);
nand U24045 (N_24045,N_23188,N_23075);
and U24046 (N_24046,N_23987,N_23898);
nor U24047 (N_24047,N_23681,N_23357);
nand U24048 (N_24048,N_23478,N_23775);
or U24049 (N_24049,N_23907,N_23474);
nor U24050 (N_24050,N_23246,N_23205);
nand U24051 (N_24051,N_23161,N_23968);
nand U24052 (N_24052,N_23166,N_23328);
nand U24053 (N_24053,N_23159,N_23819);
nor U24054 (N_24054,N_23668,N_23702);
or U24055 (N_24055,N_23966,N_23571);
and U24056 (N_24056,N_23491,N_23239);
or U24057 (N_24057,N_23976,N_23580);
or U24058 (N_24058,N_23174,N_23081);
nand U24059 (N_24059,N_23720,N_23742);
nand U24060 (N_24060,N_23360,N_23326);
or U24061 (N_24061,N_23404,N_23797);
xor U24062 (N_24062,N_23954,N_23595);
or U24063 (N_24063,N_23999,N_23718);
and U24064 (N_24064,N_23931,N_23025);
nor U24065 (N_24065,N_23938,N_23427);
and U24066 (N_24066,N_23685,N_23583);
nand U24067 (N_24067,N_23255,N_23992);
or U24068 (N_24068,N_23899,N_23343);
nand U24069 (N_24069,N_23748,N_23022);
and U24070 (N_24070,N_23094,N_23612);
and U24071 (N_24071,N_23704,N_23608);
xor U24072 (N_24072,N_23577,N_23238);
nand U24073 (N_24073,N_23644,N_23600);
nor U24074 (N_24074,N_23947,N_23194);
nor U24075 (N_24075,N_23928,N_23952);
or U24076 (N_24076,N_23047,N_23617);
nor U24077 (N_24077,N_23038,N_23509);
or U24078 (N_24078,N_23418,N_23611);
xnor U24079 (N_24079,N_23722,N_23413);
and U24080 (N_24080,N_23806,N_23867);
xor U24081 (N_24081,N_23098,N_23243);
or U24082 (N_24082,N_23209,N_23631);
nand U24083 (N_24083,N_23105,N_23164);
nand U24084 (N_24084,N_23039,N_23851);
nor U24085 (N_24085,N_23183,N_23086);
nor U24086 (N_24086,N_23627,N_23794);
and U24087 (N_24087,N_23125,N_23429);
nor U24088 (N_24088,N_23324,N_23298);
nand U24089 (N_24089,N_23686,N_23828);
or U24090 (N_24090,N_23729,N_23002);
nand U24091 (N_24091,N_23281,N_23291);
and U24092 (N_24092,N_23028,N_23504);
and U24093 (N_24093,N_23700,N_23532);
nor U24094 (N_24094,N_23176,N_23307);
xor U24095 (N_24095,N_23590,N_23861);
nand U24096 (N_24096,N_23833,N_23329);
or U24097 (N_24097,N_23944,N_23754);
or U24098 (N_24098,N_23758,N_23015);
xnor U24099 (N_24099,N_23078,N_23143);
nand U24100 (N_24100,N_23676,N_23278);
or U24101 (N_24101,N_23459,N_23331);
and U24102 (N_24102,N_23454,N_23218);
nor U24103 (N_24103,N_23597,N_23807);
and U24104 (N_24104,N_23419,N_23688);
or U24105 (N_24105,N_23318,N_23005);
nor U24106 (N_24106,N_23585,N_23212);
nand U24107 (N_24107,N_23492,N_23502);
or U24108 (N_24108,N_23813,N_23996);
and U24109 (N_24109,N_23207,N_23522);
and U24110 (N_24110,N_23642,N_23147);
nand U24111 (N_24111,N_23394,N_23562);
nor U24112 (N_24112,N_23353,N_23026);
nor U24113 (N_24113,N_23046,N_23556);
nor U24114 (N_24114,N_23370,N_23500);
and U24115 (N_24115,N_23364,N_23725);
nor U24116 (N_24116,N_23507,N_23961);
or U24117 (N_24117,N_23900,N_23031);
xor U24118 (N_24118,N_23717,N_23823);
xor U24119 (N_24119,N_23067,N_23044);
or U24120 (N_24120,N_23696,N_23203);
nor U24121 (N_24121,N_23584,N_23604);
nor U24122 (N_24122,N_23036,N_23618);
nand U24123 (N_24123,N_23674,N_23144);
or U24124 (N_24124,N_23603,N_23279);
and U24125 (N_24125,N_23913,N_23850);
nor U24126 (N_24126,N_23724,N_23021);
xor U24127 (N_24127,N_23354,N_23313);
and U24128 (N_24128,N_23241,N_23276);
xor U24129 (N_24129,N_23069,N_23133);
xor U24130 (N_24130,N_23934,N_23237);
or U24131 (N_24131,N_23189,N_23323);
and U24132 (N_24132,N_23854,N_23435);
nor U24133 (N_24133,N_23488,N_23626);
nor U24134 (N_24134,N_23625,N_23985);
xnor U24135 (N_24135,N_23653,N_23058);
nand U24136 (N_24136,N_23905,N_23182);
or U24137 (N_24137,N_23637,N_23959);
and U24138 (N_24138,N_23146,N_23735);
nor U24139 (N_24139,N_23489,N_23929);
nor U24140 (N_24140,N_23063,N_23082);
and U24141 (N_24141,N_23220,N_23493);
or U24142 (N_24142,N_23342,N_23388);
nor U24143 (N_24143,N_23930,N_23042);
xor U24144 (N_24144,N_23651,N_23272);
xnor U24145 (N_24145,N_23535,N_23247);
and U24146 (N_24146,N_23020,N_23288);
nor U24147 (N_24147,N_23974,N_23377);
and U24148 (N_24148,N_23529,N_23134);
nor U24149 (N_24149,N_23740,N_23616);
nor U24150 (N_24150,N_23461,N_23614);
nor U24151 (N_24151,N_23344,N_23520);
nor U24152 (N_24152,N_23066,N_23744);
nor U24153 (N_24153,N_23578,N_23154);
nor U24154 (N_24154,N_23780,N_23089);
and U24155 (N_24155,N_23392,N_23713);
nor U24156 (N_24156,N_23184,N_23486);
nand U24157 (N_24157,N_23848,N_23814);
and U24158 (N_24158,N_23263,N_23822);
nand U24159 (N_24159,N_23077,N_23340);
and U24160 (N_24160,N_23727,N_23308);
and U24161 (N_24161,N_23294,N_23691);
and U24162 (N_24162,N_23960,N_23951);
xor U24163 (N_24163,N_23609,N_23737);
nor U24164 (N_24164,N_23709,N_23108);
nand U24165 (N_24165,N_23936,N_23200);
and U24166 (N_24166,N_23372,N_23426);
nor U24167 (N_24167,N_23178,N_23827);
nand U24168 (N_24168,N_23716,N_23043);
xnor U24169 (N_24169,N_23883,N_23208);
nor U24170 (N_24170,N_23945,N_23710);
xor U24171 (N_24171,N_23283,N_23630);
nor U24172 (N_24172,N_23721,N_23761);
nor U24173 (N_24173,N_23569,N_23008);
and U24174 (N_24174,N_23211,N_23389);
or U24175 (N_24175,N_23395,N_23369);
nor U24176 (N_24176,N_23635,N_23027);
nand U24177 (N_24177,N_23346,N_23667);
or U24178 (N_24178,N_23763,N_23085);
and U24179 (N_24179,N_23647,N_23816);
xnor U24180 (N_24180,N_23240,N_23684);
nor U24181 (N_24181,N_23080,N_23092);
nor U24182 (N_24182,N_23692,N_23191);
or U24183 (N_24183,N_23998,N_23223);
and U24184 (N_24184,N_23363,N_23683);
nor U24185 (N_24185,N_23165,N_23712);
and U24186 (N_24186,N_23589,N_23137);
and U24187 (N_24187,N_23407,N_23621);
nand U24188 (N_24188,N_23399,N_23955);
nor U24189 (N_24189,N_23113,N_23593);
nand U24190 (N_24190,N_23510,N_23153);
xnor U24191 (N_24191,N_23887,N_23193);
and U24192 (N_24192,N_23769,N_23707);
or U24193 (N_24193,N_23753,N_23972);
nor U24194 (N_24194,N_23400,N_23187);
or U24195 (N_24195,N_23384,N_23675);
or U24196 (N_24196,N_23456,N_23736);
xor U24197 (N_24197,N_23477,N_23523);
xnor U24198 (N_24198,N_23317,N_23935);
and U24199 (N_24199,N_23497,N_23963);
and U24200 (N_24200,N_23265,N_23356);
or U24201 (N_24201,N_23749,N_23759);
and U24202 (N_24202,N_23594,N_23832);
or U24203 (N_24203,N_23870,N_23424);
and U24204 (N_24204,N_23706,N_23536);
and U24205 (N_24205,N_23895,N_23978);
nor U24206 (N_24206,N_23290,N_23054);
nor U24207 (N_24207,N_23110,N_23267);
and U24208 (N_24208,N_23473,N_23781);
and U24209 (N_24209,N_23206,N_23412);
or U24210 (N_24210,N_23817,N_23554);
or U24211 (N_24211,N_23352,N_23268);
xnor U24212 (N_24212,N_23518,N_23142);
nor U24213 (N_24213,N_23204,N_23844);
xnor U24214 (N_24214,N_23916,N_23437);
and U24215 (N_24215,N_23783,N_23877);
and U24216 (N_24216,N_23049,N_23311);
and U24217 (N_24217,N_23259,N_23697);
nand U24218 (N_24218,N_23083,N_23258);
xnor U24219 (N_24219,N_23777,N_23139);
or U24220 (N_24220,N_23231,N_23751);
nor U24221 (N_24221,N_23250,N_23990);
and U24222 (N_24222,N_23052,N_23784);
nand U24223 (N_24223,N_23458,N_23977);
xnor U24224 (N_24224,N_23414,N_23480);
or U24225 (N_24225,N_23198,N_23116);
and U24226 (N_24226,N_23774,N_23572);
xor U24227 (N_24227,N_23677,N_23649);
xor U24228 (N_24228,N_23251,N_23306);
xor U24229 (N_24229,N_23055,N_23068);
and U24230 (N_24230,N_23533,N_23476);
nor U24231 (N_24231,N_23921,N_23100);
nor U24232 (N_24232,N_23408,N_23048);
nor U24233 (N_24233,N_23076,N_23993);
and U24234 (N_24234,N_23658,N_23396);
and U24235 (N_24235,N_23619,N_23149);
or U24236 (N_24236,N_23967,N_23221);
xnor U24237 (N_24237,N_23024,N_23687);
nand U24238 (N_24238,N_23141,N_23228);
and U24239 (N_24239,N_23906,N_23368);
or U24240 (N_24240,N_23641,N_23757);
nand U24241 (N_24241,N_23715,N_23638);
xnor U24242 (N_24242,N_23890,N_23472);
xnor U24243 (N_24243,N_23528,N_23242);
xor U24244 (N_24244,N_23869,N_23444);
nand U24245 (N_24245,N_23506,N_23160);
nand U24246 (N_24246,N_23103,N_23872);
nor U24247 (N_24247,N_23558,N_23287);
xor U24248 (N_24248,N_23857,N_23514);
and U24249 (N_24249,N_23565,N_23186);
nor U24250 (N_24250,N_23981,N_23766);
xnor U24251 (N_24251,N_23462,N_23765);
xnor U24252 (N_24252,N_23917,N_23138);
nand U24253 (N_24253,N_23876,N_23986);
nor U24254 (N_24254,N_23904,N_23162);
xnor U24255 (N_24255,N_23873,N_23949);
or U24256 (N_24256,N_23132,N_23656);
or U24257 (N_24257,N_23332,N_23150);
and U24258 (N_24258,N_23547,N_23050);
nor U24259 (N_24259,N_23277,N_23016);
or U24260 (N_24260,N_23564,N_23787);
or U24261 (N_24261,N_23312,N_23064);
and U24262 (N_24262,N_23126,N_23932);
xnor U24263 (N_24263,N_23982,N_23320);
nor U24264 (N_24264,N_23484,N_23127);
and U24265 (N_24265,N_23771,N_23338);
and U24266 (N_24266,N_23910,N_23074);
xnor U24267 (N_24267,N_23515,N_23643);
or U24268 (N_24268,N_23274,N_23225);
nand U24269 (N_24269,N_23979,N_23350);
or U24270 (N_24270,N_23227,N_23889);
xnor U24271 (N_24271,N_23262,N_23512);
nor U24272 (N_24272,N_23728,N_23678);
nor U24273 (N_24273,N_23705,N_23975);
nor U24274 (N_24274,N_23269,N_23097);
nand U24275 (N_24275,N_23666,N_23285);
xnor U24276 (N_24276,N_23448,N_23257);
or U24277 (N_24277,N_23301,N_23017);
or U24278 (N_24278,N_23994,N_23390);
or U24279 (N_24279,N_23471,N_23646);
nor U24280 (N_24280,N_23483,N_23339);
xor U24281 (N_24281,N_23282,N_23734);
nor U24282 (N_24282,N_23197,N_23337);
nor U24283 (N_24283,N_23460,N_23411);
and U24284 (N_24284,N_23219,N_23826);
xor U24285 (N_24285,N_23310,N_23316);
and U24286 (N_24286,N_23417,N_23669);
or U24287 (N_24287,N_23701,N_23786);
xnor U24288 (N_24288,N_23442,N_23550);
xnor U24289 (N_24289,N_23096,N_23232);
or U24290 (N_24290,N_23542,N_23933);
nor U24291 (N_24291,N_23420,N_23778);
nor U24292 (N_24292,N_23185,N_23596);
nor U24293 (N_24293,N_23000,N_23964);
xor U24294 (N_24294,N_23950,N_23088);
or U24295 (N_24295,N_23222,N_23289);
or U24296 (N_24296,N_23365,N_23447);
xor U24297 (N_24297,N_23217,N_23040);
and U24298 (N_24298,N_23321,N_23383);
or U24299 (N_24299,N_23567,N_23121);
xnor U24300 (N_24300,N_23682,N_23755);
or U24301 (N_24301,N_23155,N_23802);
nor U24302 (N_24302,N_23436,N_23965);
nand U24303 (N_24303,N_23773,N_23852);
xnor U24304 (N_24304,N_23348,N_23897);
xnor U24305 (N_24305,N_23815,N_23422);
and U24306 (N_24306,N_23776,N_23629);
nand U24307 (N_24307,N_23847,N_23130);
xor U24308 (N_24308,N_23152,N_23136);
and U24309 (N_24309,N_23838,N_23576);
or U24310 (N_24310,N_23464,N_23151);
or U24311 (N_24311,N_23107,N_23561);
and U24312 (N_24312,N_23293,N_23072);
or U24313 (N_24313,N_23371,N_23011);
or U24314 (N_24314,N_23606,N_23505);
nor U24315 (N_24315,N_23382,N_23591);
or U24316 (N_24316,N_23210,N_23292);
or U24317 (N_24317,N_23234,N_23962);
nor U24318 (N_24318,N_23451,N_23498);
nor U24319 (N_24319,N_23559,N_23358);
and U24320 (N_24320,N_23875,N_23622);
xor U24321 (N_24321,N_23248,N_23260);
xor U24322 (N_24322,N_23620,N_23602);
or U24323 (N_24323,N_23236,N_23202);
nor U24324 (N_24324,N_23393,N_23445);
or U24325 (N_24325,N_23860,N_23768);
nand U24326 (N_24326,N_23923,N_23446);
or U24327 (N_24327,N_23273,N_23079);
nor U24328 (N_24328,N_23652,N_23534);
nand U24329 (N_24329,N_23805,N_23432);
xnor U24330 (N_24330,N_23171,N_23937);
or U24331 (N_24331,N_23109,N_23912);
xor U24332 (N_24332,N_23235,N_23789);
and U24333 (N_24333,N_23190,N_23398);
xor U24334 (N_24334,N_23662,N_23172);
nand U24335 (N_24335,N_23009,N_23610);
xor U24336 (N_24336,N_23849,N_23615);
or U24337 (N_24337,N_23730,N_23525);
nand U24338 (N_24338,N_23167,N_23811);
nand U24339 (N_24339,N_23654,N_23117);
nor U24340 (N_24340,N_23441,N_23423);
nor U24341 (N_24341,N_23747,N_23415);
nor U24342 (N_24342,N_23333,N_23573);
and U24343 (N_24343,N_23111,N_23018);
nor U24344 (N_24344,N_23632,N_23664);
xor U24345 (N_24345,N_23672,N_23764);
nand U24346 (N_24346,N_23581,N_23919);
and U24347 (N_24347,N_23800,N_23439);
nand U24348 (N_24348,N_23970,N_23057);
xor U24349 (N_24349,N_23362,N_23201);
nor U24350 (N_24350,N_23327,N_23948);
or U24351 (N_24351,N_23060,N_23156);
and U24352 (N_24352,N_23531,N_23538);
or U24353 (N_24353,N_23373,N_23014);
and U24354 (N_24354,N_23598,N_23482);
and U24355 (N_24355,N_23714,N_23361);
nand U24356 (N_24356,N_23566,N_23582);
and U24357 (N_24357,N_23253,N_23772);
nor U24358 (N_24358,N_23943,N_23264);
and U24359 (N_24359,N_23853,N_23841);
and U24360 (N_24360,N_23041,N_23592);
xor U24361 (N_24361,N_23636,N_23463);
nand U24362 (N_24362,N_23980,N_23886);
xor U24363 (N_24363,N_23455,N_23387);
nor U24364 (N_24364,N_23693,N_23095);
nand U24365 (N_24365,N_23623,N_23158);
nor U24366 (N_24366,N_23719,N_23539);
or U24367 (N_24367,N_23120,N_23003);
nand U24368 (N_24368,N_23325,N_23989);
xor U24369 (N_24369,N_23599,N_23660);
and U24370 (N_24370,N_23628,N_23261);
nor U24371 (N_24371,N_23380,N_23181);
or U24372 (N_24372,N_23892,N_23467);
nor U24373 (N_24373,N_23732,N_23405);
nor U24374 (N_24374,N_23812,N_23891);
nor U24375 (N_24375,N_23330,N_23379);
xnor U24376 (N_24376,N_23481,N_23624);
xor U24377 (N_24377,N_23129,N_23254);
nor U24378 (N_24378,N_23359,N_23971);
xor U24379 (N_24379,N_23694,N_23524);
or U24380 (N_24380,N_23540,N_23902);
and U24381 (N_24381,N_23029,N_23679);
or U24382 (N_24382,N_23946,N_23738);
or U24383 (N_24383,N_23824,N_23177);
nor U24384 (N_24384,N_23884,N_23703);
or U24385 (N_24385,N_23106,N_23297);
nor U24386 (N_24386,N_23557,N_23425);
xor U24387 (N_24387,N_23053,N_23314);
xnor U24388 (N_24388,N_23548,N_23030);
nand U24389 (N_24389,N_23229,N_23645);
nor U24390 (N_24390,N_23871,N_23804);
and U24391 (N_24391,N_23821,N_23745);
and U24392 (N_24392,N_23487,N_23801);
nand U24393 (N_24393,N_23195,N_23726);
or U24394 (N_24394,N_23791,N_23061);
xnor U24395 (N_24395,N_23180,N_23680);
xnor U24396 (N_24396,N_23549,N_23032);
nand U24397 (N_24397,N_23299,N_23792);
and U24398 (N_24398,N_23551,N_23173);
nor U24399 (N_24399,N_23544,N_23019);
nor U24400 (N_24400,N_23410,N_23839);
or U24401 (N_24401,N_23864,N_23034);
and U24402 (N_24402,N_23157,N_23428);
nand U24403 (N_24403,N_23846,N_23374);
or U24404 (N_24404,N_23013,N_23750);
and U24405 (N_24405,N_23059,N_23918);
and U24406 (N_24406,N_23588,N_23213);
or U24407 (N_24407,N_23785,N_23479);
and U24408 (N_24408,N_23516,N_23926);
nor U24409 (N_24409,N_23655,N_23909);
or U24410 (N_24410,N_23659,N_23475);
and U24411 (N_24411,N_23163,N_23663);
xnor U24412 (N_24412,N_23035,N_23452);
nor U24413 (N_24413,N_23334,N_23640);
xor U24414 (N_24414,N_23465,N_23770);
or U24415 (N_24415,N_23501,N_23731);
nand U24416 (N_24416,N_23803,N_23319);
nor U24417 (N_24417,N_23006,N_23115);
xor U24418 (N_24418,N_23335,N_23302);
and U24419 (N_24419,N_23671,N_23526);
xor U24420 (N_24420,N_23010,N_23756);
and U24421 (N_24421,N_23840,N_23494);
and U24422 (N_24422,N_23991,N_23689);
xor U24423 (N_24423,N_23587,N_23914);
or U24424 (N_24424,N_23118,N_23245);
xnor U24425 (N_24425,N_23216,N_23099);
or U24426 (N_24426,N_23056,N_23140);
xnor U24427 (N_24427,N_23810,N_23570);
and U24428 (N_24428,N_23175,N_23226);
or U24429 (N_24429,N_23790,N_23956);
and U24430 (N_24430,N_23233,N_23779);
and U24431 (N_24431,N_23336,N_23752);
and U24432 (N_24432,N_23284,N_23101);
xor U24433 (N_24433,N_23215,N_23087);
nor U24434 (N_24434,N_23673,N_23349);
and U24435 (N_24435,N_23969,N_23434);
xnor U24436 (N_24436,N_23995,N_23825);
or U24437 (N_24437,N_23808,N_23093);
nand U24438 (N_24438,N_23104,N_23315);
xnor U24439 (N_24439,N_23148,N_23657);
nor U24440 (N_24440,N_23347,N_23957);
or U24441 (N_24441,N_23782,N_23894);
xor U24442 (N_24442,N_23586,N_23530);
nor U24443 (N_24443,N_23984,N_23416);
xnor U24444 (N_24444,N_23386,N_23122);
or U24445 (N_24445,N_23605,N_23988);
or U24446 (N_24446,N_23788,N_23874);
and U24447 (N_24447,N_23051,N_23303);
xnor U24448 (N_24448,N_23466,N_23402);
nor U24449 (N_24449,N_23842,N_23537);
nand U24450 (N_24450,N_23135,N_23575);
or U24451 (N_24451,N_23230,N_23723);
xnor U24452 (N_24452,N_23449,N_23563);
xor U24453 (N_24453,N_23070,N_23743);
nand U24454 (N_24454,N_23767,N_23555);
nand U24455 (N_24455,N_23862,N_23834);
nor U24456 (N_24456,N_23859,N_23661);
xnor U24457 (N_24457,N_23045,N_23865);
and U24458 (N_24458,N_23433,N_23922);
nand U24459 (N_24459,N_23888,N_23708);
or U24460 (N_24460,N_23280,N_23073);
or U24461 (N_24461,N_23355,N_23495);
or U24462 (N_24462,N_23863,N_23196);
and U24463 (N_24463,N_23880,N_23119);
nor U24464 (N_24464,N_23367,N_23809);
nor U24465 (N_24465,N_23440,N_23958);
nor U24466 (N_24466,N_23381,N_23168);
and U24467 (N_24467,N_23882,N_23114);
xor U24468 (N_24468,N_23345,N_23001);
or U24469 (N_24469,N_23503,N_23953);
nor U24470 (N_24470,N_23739,N_23322);
nor U24471 (N_24471,N_23270,N_23007);
xor U24472 (N_24472,N_23665,N_23179);
nand U24473 (N_24473,N_23831,N_23796);
nor U24474 (N_24474,N_23521,N_23545);
nor U24475 (N_24475,N_23145,N_23084);
or U24476 (N_24476,N_23911,N_23401);
or U24477 (N_24477,N_23798,N_23517);
and U24478 (N_24478,N_23199,N_23983);
xnor U24479 (N_24479,N_23508,N_23878);
and U24480 (N_24480,N_23908,N_23858);
nor U24481 (N_24481,N_23385,N_23300);
or U24482 (N_24482,N_23893,N_23438);
and U24483 (N_24483,N_23091,N_23711);
xnor U24484 (N_24484,N_23837,N_23249);
or U24485 (N_24485,N_23868,N_23634);
nor U24486 (N_24486,N_23131,N_23633);
or U24487 (N_24487,N_23090,N_23450);
nor U24488 (N_24488,N_23939,N_23925);
nand U24489 (N_24489,N_23170,N_23062);
xor U24490 (N_24490,N_23457,N_23881);
xor U24491 (N_24491,N_23613,N_23650);
xnor U24492 (N_24492,N_23023,N_23271);
and U24493 (N_24493,N_23513,N_23698);
or U24494 (N_24494,N_23065,N_23924);
nand U24495 (N_24495,N_23511,N_23366);
and U24496 (N_24496,N_23920,N_23699);
xnor U24497 (N_24497,N_23973,N_23829);
nor U24498 (N_24498,N_23568,N_23836);
or U24499 (N_24499,N_23224,N_23244);
or U24500 (N_24500,N_23338,N_23041);
xor U24501 (N_24501,N_23857,N_23725);
xor U24502 (N_24502,N_23191,N_23771);
or U24503 (N_24503,N_23786,N_23322);
nand U24504 (N_24504,N_23482,N_23650);
or U24505 (N_24505,N_23085,N_23881);
nor U24506 (N_24506,N_23534,N_23896);
nand U24507 (N_24507,N_23556,N_23105);
xor U24508 (N_24508,N_23231,N_23114);
nor U24509 (N_24509,N_23919,N_23842);
nor U24510 (N_24510,N_23043,N_23943);
or U24511 (N_24511,N_23813,N_23326);
nor U24512 (N_24512,N_23639,N_23917);
nor U24513 (N_24513,N_23323,N_23498);
xor U24514 (N_24514,N_23718,N_23496);
and U24515 (N_24515,N_23244,N_23880);
nor U24516 (N_24516,N_23643,N_23286);
or U24517 (N_24517,N_23282,N_23998);
or U24518 (N_24518,N_23729,N_23100);
nand U24519 (N_24519,N_23803,N_23340);
or U24520 (N_24520,N_23437,N_23014);
and U24521 (N_24521,N_23142,N_23796);
xnor U24522 (N_24522,N_23637,N_23240);
or U24523 (N_24523,N_23560,N_23139);
nand U24524 (N_24524,N_23201,N_23796);
nor U24525 (N_24525,N_23282,N_23001);
nand U24526 (N_24526,N_23987,N_23054);
nand U24527 (N_24527,N_23170,N_23696);
or U24528 (N_24528,N_23526,N_23118);
nor U24529 (N_24529,N_23677,N_23772);
xor U24530 (N_24530,N_23694,N_23119);
and U24531 (N_24531,N_23480,N_23335);
nor U24532 (N_24532,N_23013,N_23578);
nor U24533 (N_24533,N_23475,N_23459);
and U24534 (N_24534,N_23533,N_23066);
nor U24535 (N_24535,N_23615,N_23687);
or U24536 (N_24536,N_23876,N_23882);
or U24537 (N_24537,N_23851,N_23907);
xor U24538 (N_24538,N_23564,N_23985);
and U24539 (N_24539,N_23212,N_23719);
xor U24540 (N_24540,N_23661,N_23666);
and U24541 (N_24541,N_23480,N_23504);
and U24542 (N_24542,N_23798,N_23451);
xor U24543 (N_24543,N_23729,N_23372);
xnor U24544 (N_24544,N_23441,N_23704);
nand U24545 (N_24545,N_23365,N_23841);
xor U24546 (N_24546,N_23863,N_23199);
nor U24547 (N_24547,N_23730,N_23504);
nand U24548 (N_24548,N_23370,N_23896);
and U24549 (N_24549,N_23817,N_23893);
or U24550 (N_24550,N_23166,N_23184);
and U24551 (N_24551,N_23986,N_23128);
nand U24552 (N_24552,N_23429,N_23685);
nand U24553 (N_24553,N_23476,N_23126);
xor U24554 (N_24554,N_23097,N_23999);
nand U24555 (N_24555,N_23034,N_23974);
nor U24556 (N_24556,N_23208,N_23784);
or U24557 (N_24557,N_23198,N_23226);
or U24558 (N_24558,N_23962,N_23836);
xor U24559 (N_24559,N_23412,N_23798);
xor U24560 (N_24560,N_23015,N_23195);
xnor U24561 (N_24561,N_23211,N_23256);
nor U24562 (N_24562,N_23800,N_23960);
or U24563 (N_24563,N_23705,N_23814);
nand U24564 (N_24564,N_23800,N_23823);
nor U24565 (N_24565,N_23371,N_23554);
and U24566 (N_24566,N_23756,N_23181);
xnor U24567 (N_24567,N_23457,N_23412);
and U24568 (N_24568,N_23934,N_23555);
nor U24569 (N_24569,N_23804,N_23230);
or U24570 (N_24570,N_23496,N_23515);
and U24571 (N_24571,N_23825,N_23872);
xnor U24572 (N_24572,N_23151,N_23669);
nor U24573 (N_24573,N_23369,N_23385);
nor U24574 (N_24574,N_23458,N_23869);
and U24575 (N_24575,N_23077,N_23872);
or U24576 (N_24576,N_23233,N_23530);
nor U24577 (N_24577,N_23971,N_23432);
and U24578 (N_24578,N_23722,N_23166);
nand U24579 (N_24579,N_23971,N_23006);
or U24580 (N_24580,N_23497,N_23094);
nand U24581 (N_24581,N_23763,N_23206);
xnor U24582 (N_24582,N_23852,N_23214);
nor U24583 (N_24583,N_23899,N_23835);
nor U24584 (N_24584,N_23937,N_23087);
xor U24585 (N_24585,N_23050,N_23236);
nand U24586 (N_24586,N_23347,N_23372);
nand U24587 (N_24587,N_23585,N_23228);
xor U24588 (N_24588,N_23813,N_23367);
or U24589 (N_24589,N_23028,N_23886);
or U24590 (N_24590,N_23997,N_23766);
nor U24591 (N_24591,N_23432,N_23723);
nand U24592 (N_24592,N_23531,N_23861);
or U24593 (N_24593,N_23873,N_23756);
or U24594 (N_24594,N_23087,N_23468);
xnor U24595 (N_24595,N_23537,N_23897);
or U24596 (N_24596,N_23476,N_23794);
xnor U24597 (N_24597,N_23960,N_23874);
nand U24598 (N_24598,N_23979,N_23124);
nor U24599 (N_24599,N_23861,N_23129);
xor U24600 (N_24600,N_23662,N_23611);
and U24601 (N_24601,N_23930,N_23437);
or U24602 (N_24602,N_23477,N_23677);
or U24603 (N_24603,N_23333,N_23716);
and U24604 (N_24604,N_23325,N_23231);
nor U24605 (N_24605,N_23298,N_23628);
nand U24606 (N_24606,N_23870,N_23846);
or U24607 (N_24607,N_23102,N_23384);
xor U24608 (N_24608,N_23166,N_23021);
or U24609 (N_24609,N_23220,N_23185);
xor U24610 (N_24610,N_23915,N_23209);
nand U24611 (N_24611,N_23213,N_23699);
or U24612 (N_24612,N_23505,N_23717);
and U24613 (N_24613,N_23615,N_23283);
nor U24614 (N_24614,N_23022,N_23169);
nand U24615 (N_24615,N_23587,N_23961);
nor U24616 (N_24616,N_23113,N_23322);
nor U24617 (N_24617,N_23448,N_23814);
nor U24618 (N_24618,N_23897,N_23713);
xnor U24619 (N_24619,N_23089,N_23941);
nor U24620 (N_24620,N_23298,N_23164);
nor U24621 (N_24621,N_23301,N_23053);
or U24622 (N_24622,N_23924,N_23520);
or U24623 (N_24623,N_23737,N_23835);
or U24624 (N_24624,N_23330,N_23820);
xnor U24625 (N_24625,N_23077,N_23342);
nand U24626 (N_24626,N_23493,N_23558);
or U24627 (N_24627,N_23212,N_23686);
xor U24628 (N_24628,N_23014,N_23445);
nor U24629 (N_24629,N_23134,N_23108);
xnor U24630 (N_24630,N_23640,N_23919);
or U24631 (N_24631,N_23327,N_23082);
xor U24632 (N_24632,N_23583,N_23100);
or U24633 (N_24633,N_23100,N_23400);
or U24634 (N_24634,N_23399,N_23766);
nor U24635 (N_24635,N_23419,N_23808);
nor U24636 (N_24636,N_23887,N_23563);
and U24637 (N_24637,N_23798,N_23181);
or U24638 (N_24638,N_23603,N_23091);
nand U24639 (N_24639,N_23911,N_23279);
and U24640 (N_24640,N_23583,N_23804);
and U24641 (N_24641,N_23452,N_23377);
or U24642 (N_24642,N_23743,N_23406);
xnor U24643 (N_24643,N_23639,N_23331);
nand U24644 (N_24644,N_23800,N_23790);
and U24645 (N_24645,N_23047,N_23104);
xnor U24646 (N_24646,N_23242,N_23711);
nand U24647 (N_24647,N_23622,N_23545);
and U24648 (N_24648,N_23533,N_23707);
and U24649 (N_24649,N_23660,N_23032);
nor U24650 (N_24650,N_23201,N_23090);
nor U24651 (N_24651,N_23808,N_23114);
nor U24652 (N_24652,N_23337,N_23489);
nand U24653 (N_24653,N_23091,N_23756);
and U24654 (N_24654,N_23996,N_23567);
nand U24655 (N_24655,N_23025,N_23887);
and U24656 (N_24656,N_23625,N_23348);
or U24657 (N_24657,N_23309,N_23533);
and U24658 (N_24658,N_23538,N_23923);
xnor U24659 (N_24659,N_23445,N_23186);
or U24660 (N_24660,N_23740,N_23720);
or U24661 (N_24661,N_23175,N_23438);
nor U24662 (N_24662,N_23096,N_23106);
nand U24663 (N_24663,N_23920,N_23655);
nor U24664 (N_24664,N_23723,N_23352);
or U24665 (N_24665,N_23343,N_23362);
xor U24666 (N_24666,N_23297,N_23685);
or U24667 (N_24667,N_23832,N_23352);
xnor U24668 (N_24668,N_23637,N_23358);
nand U24669 (N_24669,N_23053,N_23562);
nand U24670 (N_24670,N_23437,N_23226);
nor U24671 (N_24671,N_23298,N_23459);
and U24672 (N_24672,N_23252,N_23545);
nand U24673 (N_24673,N_23155,N_23158);
xnor U24674 (N_24674,N_23718,N_23177);
or U24675 (N_24675,N_23046,N_23102);
nand U24676 (N_24676,N_23342,N_23356);
or U24677 (N_24677,N_23589,N_23145);
or U24678 (N_24678,N_23917,N_23327);
or U24679 (N_24679,N_23607,N_23264);
and U24680 (N_24680,N_23818,N_23278);
nor U24681 (N_24681,N_23170,N_23173);
and U24682 (N_24682,N_23449,N_23713);
or U24683 (N_24683,N_23323,N_23151);
and U24684 (N_24684,N_23138,N_23267);
nand U24685 (N_24685,N_23847,N_23287);
and U24686 (N_24686,N_23427,N_23970);
and U24687 (N_24687,N_23463,N_23008);
and U24688 (N_24688,N_23927,N_23767);
xor U24689 (N_24689,N_23689,N_23248);
or U24690 (N_24690,N_23726,N_23633);
and U24691 (N_24691,N_23365,N_23652);
nand U24692 (N_24692,N_23178,N_23787);
or U24693 (N_24693,N_23321,N_23534);
xor U24694 (N_24694,N_23230,N_23663);
and U24695 (N_24695,N_23365,N_23164);
xnor U24696 (N_24696,N_23007,N_23898);
nor U24697 (N_24697,N_23496,N_23069);
nand U24698 (N_24698,N_23303,N_23975);
xnor U24699 (N_24699,N_23557,N_23606);
xor U24700 (N_24700,N_23998,N_23132);
and U24701 (N_24701,N_23422,N_23292);
nor U24702 (N_24702,N_23998,N_23625);
nand U24703 (N_24703,N_23647,N_23099);
and U24704 (N_24704,N_23857,N_23777);
nor U24705 (N_24705,N_23393,N_23400);
nor U24706 (N_24706,N_23240,N_23772);
xor U24707 (N_24707,N_23950,N_23778);
xor U24708 (N_24708,N_23073,N_23521);
nor U24709 (N_24709,N_23221,N_23622);
and U24710 (N_24710,N_23049,N_23875);
nor U24711 (N_24711,N_23153,N_23543);
nand U24712 (N_24712,N_23677,N_23618);
xnor U24713 (N_24713,N_23688,N_23932);
nand U24714 (N_24714,N_23187,N_23575);
or U24715 (N_24715,N_23306,N_23888);
nor U24716 (N_24716,N_23306,N_23359);
nand U24717 (N_24717,N_23388,N_23131);
or U24718 (N_24718,N_23678,N_23285);
xor U24719 (N_24719,N_23902,N_23159);
nand U24720 (N_24720,N_23697,N_23101);
xnor U24721 (N_24721,N_23758,N_23322);
nand U24722 (N_24722,N_23132,N_23027);
nand U24723 (N_24723,N_23000,N_23054);
nor U24724 (N_24724,N_23306,N_23804);
nor U24725 (N_24725,N_23473,N_23099);
or U24726 (N_24726,N_23621,N_23446);
or U24727 (N_24727,N_23278,N_23531);
or U24728 (N_24728,N_23031,N_23693);
xnor U24729 (N_24729,N_23560,N_23915);
and U24730 (N_24730,N_23792,N_23439);
xor U24731 (N_24731,N_23693,N_23146);
or U24732 (N_24732,N_23517,N_23546);
and U24733 (N_24733,N_23147,N_23256);
or U24734 (N_24734,N_23602,N_23287);
nor U24735 (N_24735,N_23791,N_23743);
or U24736 (N_24736,N_23470,N_23785);
nor U24737 (N_24737,N_23759,N_23698);
or U24738 (N_24738,N_23628,N_23718);
and U24739 (N_24739,N_23633,N_23201);
nor U24740 (N_24740,N_23111,N_23776);
and U24741 (N_24741,N_23088,N_23224);
xnor U24742 (N_24742,N_23103,N_23580);
and U24743 (N_24743,N_23039,N_23728);
and U24744 (N_24744,N_23385,N_23230);
or U24745 (N_24745,N_23934,N_23874);
nor U24746 (N_24746,N_23303,N_23199);
or U24747 (N_24747,N_23198,N_23406);
nand U24748 (N_24748,N_23488,N_23555);
xnor U24749 (N_24749,N_23255,N_23778);
or U24750 (N_24750,N_23280,N_23616);
and U24751 (N_24751,N_23519,N_23212);
or U24752 (N_24752,N_23243,N_23176);
and U24753 (N_24753,N_23457,N_23162);
and U24754 (N_24754,N_23242,N_23523);
and U24755 (N_24755,N_23030,N_23806);
nand U24756 (N_24756,N_23429,N_23980);
xor U24757 (N_24757,N_23349,N_23436);
or U24758 (N_24758,N_23305,N_23663);
nand U24759 (N_24759,N_23049,N_23429);
or U24760 (N_24760,N_23552,N_23125);
and U24761 (N_24761,N_23455,N_23748);
or U24762 (N_24762,N_23244,N_23086);
nor U24763 (N_24763,N_23377,N_23074);
and U24764 (N_24764,N_23658,N_23587);
nor U24765 (N_24765,N_23442,N_23824);
and U24766 (N_24766,N_23648,N_23255);
xnor U24767 (N_24767,N_23728,N_23548);
nand U24768 (N_24768,N_23113,N_23555);
or U24769 (N_24769,N_23978,N_23604);
nand U24770 (N_24770,N_23860,N_23476);
nand U24771 (N_24771,N_23277,N_23110);
and U24772 (N_24772,N_23531,N_23596);
xnor U24773 (N_24773,N_23538,N_23505);
or U24774 (N_24774,N_23557,N_23453);
nand U24775 (N_24775,N_23733,N_23542);
and U24776 (N_24776,N_23945,N_23351);
or U24777 (N_24777,N_23683,N_23577);
xnor U24778 (N_24778,N_23507,N_23790);
and U24779 (N_24779,N_23119,N_23923);
or U24780 (N_24780,N_23665,N_23029);
nor U24781 (N_24781,N_23374,N_23051);
or U24782 (N_24782,N_23574,N_23714);
nand U24783 (N_24783,N_23458,N_23549);
xnor U24784 (N_24784,N_23586,N_23185);
nand U24785 (N_24785,N_23009,N_23434);
or U24786 (N_24786,N_23674,N_23711);
nor U24787 (N_24787,N_23505,N_23806);
and U24788 (N_24788,N_23216,N_23664);
or U24789 (N_24789,N_23411,N_23778);
and U24790 (N_24790,N_23376,N_23668);
and U24791 (N_24791,N_23733,N_23574);
and U24792 (N_24792,N_23797,N_23186);
nand U24793 (N_24793,N_23263,N_23276);
nor U24794 (N_24794,N_23996,N_23001);
nor U24795 (N_24795,N_23186,N_23235);
xor U24796 (N_24796,N_23127,N_23517);
nor U24797 (N_24797,N_23005,N_23362);
xor U24798 (N_24798,N_23601,N_23405);
nand U24799 (N_24799,N_23734,N_23220);
nor U24800 (N_24800,N_23727,N_23762);
or U24801 (N_24801,N_23891,N_23251);
and U24802 (N_24802,N_23330,N_23160);
or U24803 (N_24803,N_23021,N_23114);
or U24804 (N_24804,N_23571,N_23375);
xor U24805 (N_24805,N_23970,N_23707);
xnor U24806 (N_24806,N_23054,N_23063);
nand U24807 (N_24807,N_23397,N_23650);
or U24808 (N_24808,N_23989,N_23821);
nand U24809 (N_24809,N_23627,N_23919);
nand U24810 (N_24810,N_23529,N_23218);
nor U24811 (N_24811,N_23800,N_23028);
xor U24812 (N_24812,N_23598,N_23987);
nor U24813 (N_24813,N_23216,N_23432);
and U24814 (N_24814,N_23222,N_23815);
or U24815 (N_24815,N_23708,N_23376);
nor U24816 (N_24816,N_23646,N_23845);
xnor U24817 (N_24817,N_23320,N_23176);
nand U24818 (N_24818,N_23678,N_23777);
xor U24819 (N_24819,N_23607,N_23711);
nand U24820 (N_24820,N_23085,N_23904);
nor U24821 (N_24821,N_23542,N_23346);
and U24822 (N_24822,N_23850,N_23535);
nand U24823 (N_24823,N_23093,N_23770);
nor U24824 (N_24824,N_23988,N_23878);
nand U24825 (N_24825,N_23433,N_23713);
xor U24826 (N_24826,N_23057,N_23134);
or U24827 (N_24827,N_23534,N_23201);
or U24828 (N_24828,N_23183,N_23133);
nor U24829 (N_24829,N_23199,N_23972);
nand U24830 (N_24830,N_23752,N_23435);
and U24831 (N_24831,N_23735,N_23958);
nand U24832 (N_24832,N_23454,N_23537);
or U24833 (N_24833,N_23122,N_23490);
and U24834 (N_24834,N_23651,N_23204);
and U24835 (N_24835,N_23721,N_23760);
and U24836 (N_24836,N_23072,N_23781);
xor U24837 (N_24837,N_23039,N_23350);
or U24838 (N_24838,N_23295,N_23444);
xnor U24839 (N_24839,N_23425,N_23336);
nand U24840 (N_24840,N_23843,N_23239);
nand U24841 (N_24841,N_23073,N_23973);
and U24842 (N_24842,N_23358,N_23668);
and U24843 (N_24843,N_23653,N_23250);
and U24844 (N_24844,N_23282,N_23987);
xor U24845 (N_24845,N_23336,N_23404);
xnor U24846 (N_24846,N_23243,N_23583);
nand U24847 (N_24847,N_23271,N_23751);
xor U24848 (N_24848,N_23444,N_23561);
nor U24849 (N_24849,N_23095,N_23070);
nand U24850 (N_24850,N_23356,N_23662);
xor U24851 (N_24851,N_23220,N_23290);
xor U24852 (N_24852,N_23952,N_23609);
xor U24853 (N_24853,N_23143,N_23595);
xnor U24854 (N_24854,N_23010,N_23114);
nand U24855 (N_24855,N_23474,N_23547);
or U24856 (N_24856,N_23566,N_23055);
nand U24857 (N_24857,N_23037,N_23569);
nand U24858 (N_24858,N_23298,N_23171);
or U24859 (N_24859,N_23745,N_23581);
and U24860 (N_24860,N_23607,N_23006);
xnor U24861 (N_24861,N_23684,N_23271);
and U24862 (N_24862,N_23209,N_23072);
nand U24863 (N_24863,N_23167,N_23503);
or U24864 (N_24864,N_23953,N_23299);
and U24865 (N_24865,N_23270,N_23848);
or U24866 (N_24866,N_23818,N_23967);
xnor U24867 (N_24867,N_23546,N_23237);
and U24868 (N_24868,N_23263,N_23316);
or U24869 (N_24869,N_23931,N_23381);
nand U24870 (N_24870,N_23613,N_23187);
and U24871 (N_24871,N_23871,N_23426);
nand U24872 (N_24872,N_23782,N_23836);
and U24873 (N_24873,N_23399,N_23690);
nand U24874 (N_24874,N_23646,N_23025);
xor U24875 (N_24875,N_23872,N_23189);
xnor U24876 (N_24876,N_23829,N_23287);
or U24877 (N_24877,N_23998,N_23638);
xor U24878 (N_24878,N_23726,N_23291);
and U24879 (N_24879,N_23885,N_23585);
or U24880 (N_24880,N_23171,N_23650);
xor U24881 (N_24881,N_23379,N_23421);
or U24882 (N_24882,N_23671,N_23066);
nor U24883 (N_24883,N_23963,N_23249);
nand U24884 (N_24884,N_23098,N_23262);
nor U24885 (N_24885,N_23697,N_23170);
nand U24886 (N_24886,N_23919,N_23036);
nand U24887 (N_24887,N_23505,N_23833);
and U24888 (N_24888,N_23917,N_23712);
nand U24889 (N_24889,N_23843,N_23474);
and U24890 (N_24890,N_23906,N_23475);
nand U24891 (N_24891,N_23110,N_23845);
nor U24892 (N_24892,N_23326,N_23380);
and U24893 (N_24893,N_23235,N_23694);
nand U24894 (N_24894,N_23064,N_23652);
nand U24895 (N_24895,N_23002,N_23885);
and U24896 (N_24896,N_23499,N_23683);
nand U24897 (N_24897,N_23355,N_23237);
and U24898 (N_24898,N_23398,N_23233);
and U24899 (N_24899,N_23934,N_23130);
xor U24900 (N_24900,N_23558,N_23665);
nor U24901 (N_24901,N_23407,N_23987);
or U24902 (N_24902,N_23819,N_23956);
or U24903 (N_24903,N_23407,N_23865);
nor U24904 (N_24904,N_23862,N_23586);
and U24905 (N_24905,N_23418,N_23628);
and U24906 (N_24906,N_23497,N_23355);
and U24907 (N_24907,N_23708,N_23990);
and U24908 (N_24908,N_23635,N_23480);
nand U24909 (N_24909,N_23215,N_23088);
xnor U24910 (N_24910,N_23120,N_23229);
and U24911 (N_24911,N_23972,N_23139);
or U24912 (N_24912,N_23435,N_23381);
xnor U24913 (N_24913,N_23774,N_23677);
nand U24914 (N_24914,N_23222,N_23111);
nor U24915 (N_24915,N_23076,N_23310);
and U24916 (N_24916,N_23592,N_23591);
xnor U24917 (N_24917,N_23988,N_23794);
nor U24918 (N_24918,N_23460,N_23088);
nand U24919 (N_24919,N_23429,N_23698);
and U24920 (N_24920,N_23821,N_23488);
xor U24921 (N_24921,N_23307,N_23600);
nor U24922 (N_24922,N_23481,N_23421);
and U24923 (N_24923,N_23928,N_23481);
and U24924 (N_24924,N_23386,N_23285);
xnor U24925 (N_24925,N_23032,N_23553);
nand U24926 (N_24926,N_23875,N_23093);
and U24927 (N_24927,N_23636,N_23557);
nor U24928 (N_24928,N_23601,N_23196);
nor U24929 (N_24929,N_23474,N_23492);
nand U24930 (N_24930,N_23238,N_23163);
or U24931 (N_24931,N_23442,N_23813);
nor U24932 (N_24932,N_23602,N_23809);
nand U24933 (N_24933,N_23595,N_23000);
and U24934 (N_24934,N_23917,N_23112);
or U24935 (N_24935,N_23981,N_23300);
and U24936 (N_24936,N_23480,N_23065);
and U24937 (N_24937,N_23226,N_23321);
or U24938 (N_24938,N_23174,N_23508);
or U24939 (N_24939,N_23243,N_23137);
or U24940 (N_24940,N_23810,N_23514);
and U24941 (N_24941,N_23344,N_23097);
xor U24942 (N_24942,N_23955,N_23974);
or U24943 (N_24943,N_23780,N_23878);
nor U24944 (N_24944,N_23318,N_23845);
nand U24945 (N_24945,N_23897,N_23590);
or U24946 (N_24946,N_23646,N_23126);
xor U24947 (N_24947,N_23352,N_23489);
and U24948 (N_24948,N_23108,N_23275);
xor U24949 (N_24949,N_23997,N_23330);
xor U24950 (N_24950,N_23799,N_23100);
or U24951 (N_24951,N_23121,N_23935);
and U24952 (N_24952,N_23352,N_23503);
or U24953 (N_24953,N_23844,N_23170);
or U24954 (N_24954,N_23814,N_23674);
and U24955 (N_24955,N_23582,N_23602);
and U24956 (N_24956,N_23800,N_23982);
nand U24957 (N_24957,N_23457,N_23479);
nor U24958 (N_24958,N_23325,N_23272);
xnor U24959 (N_24959,N_23843,N_23849);
or U24960 (N_24960,N_23591,N_23005);
nor U24961 (N_24961,N_23615,N_23939);
xor U24962 (N_24962,N_23714,N_23242);
or U24963 (N_24963,N_23539,N_23789);
nor U24964 (N_24964,N_23928,N_23723);
xor U24965 (N_24965,N_23732,N_23016);
xor U24966 (N_24966,N_23073,N_23845);
nand U24967 (N_24967,N_23246,N_23848);
nor U24968 (N_24968,N_23181,N_23567);
and U24969 (N_24969,N_23113,N_23371);
xor U24970 (N_24970,N_23562,N_23875);
and U24971 (N_24971,N_23765,N_23269);
nand U24972 (N_24972,N_23689,N_23238);
nor U24973 (N_24973,N_23279,N_23595);
nand U24974 (N_24974,N_23495,N_23486);
and U24975 (N_24975,N_23103,N_23235);
or U24976 (N_24976,N_23185,N_23527);
and U24977 (N_24977,N_23257,N_23273);
nand U24978 (N_24978,N_23246,N_23402);
xnor U24979 (N_24979,N_23126,N_23787);
or U24980 (N_24980,N_23948,N_23676);
xor U24981 (N_24981,N_23093,N_23651);
nor U24982 (N_24982,N_23345,N_23364);
nor U24983 (N_24983,N_23637,N_23227);
or U24984 (N_24984,N_23341,N_23280);
or U24985 (N_24985,N_23745,N_23411);
xnor U24986 (N_24986,N_23583,N_23408);
or U24987 (N_24987,N_23489,N_23560);
xnor U24988 (N_24988,N_23803,N_23977);
nor U24989 (N_24989,N_23726,N_23469);
xnor U24990 (N_24990,N_23530,N_23017);
or U24991 (N_24991,N_23602,N_23283);
xnor U24992 (N_24992,N_23261,N_23807);
nor U24993 (N_24993,N_23961,N_23040);
nand U24994 (N_24994,N_23542,N_23358);
nor U24995 (N_24995,N_23327,N_23942);
nand U24996 (N_24996,N_23895,N_23267);
nand U24997 (N_24997,N_23227,N_23624);
nor U24998 (N_24998,N_23655,N_23264);
nor U24999 (N_24999,N_23502,N_23900);
nand U25000 (N_25000,N_24582,N_24808);
nand U25001 (N_25001,N_24666,N_24597);
nand U25002 (N_25002,N_24458,N_24440);
and U25003 (N_25003,N_24335,N_24815);
nor U25004 (N_25004,N_24369,N_24384);
nor U25005 (N_25005,N_24093,N_24621);
nor U25006 (N_25006,N_24619,N_24333);
or U25007 (N_25007,N_24761,N_24600);
xnor U25008 (N_25008,N_24089,N_24747);
or U25009 (N_25009,N_24324,N_24095);
or U25010 (N_25010,N_24437,N_24935);
and U25011 (N_25011,N_24628,N_24494);
or U25012 (N_25012,N_24717,N_24834);
xor U25013 (N_25013,N_24595,N_24280);
or U25014 (N_25014,N_24147,N_24273);
nor U25015 (N_25015,N_24455,N_24577);
or U25016 (N_25016,N_24130,N_24141);
nand U25017 (N_25017,N_24902,N_24780);
nor U25018 (N_25018,N_24565,N_24194);
or U25019 (N_25019,N_24844,N_24842);
xnor U25020 (N_25020,N_24905,N_24078);
nand U25021 (N_25021,N_24336,N_24663);
and U25022 (N_25022,N_24830,N_24138);
and U25023 (N_25023,N_24061,N_24643);
and U25024 (N_25024,N_24197,N_24681);
nor U25025 (N_25025,N_24738,N_24325);
nor U25026 (N_25026,N_24735,N_24987);
or U25027 (N_25027,N_24817,N_24288);
nand U25028 (N_25028,N_24835,N_24930);
and U25029 (N_25029,N_24013,N_24563);
or U25030 (N_25030,N_24767,N_24493);
nor U25031 (N_25031,N_24328,N_24202);
nor U25032 (N_25032,N_24166,N_24322);
nor U25033 (N_25033,N_24318,N_24572);
and U25034 (N_25034,N_24467,N_24486);
and U25035 (N_25035,N_24272,N_24199);
or U25036 (N_25036,N_24119,N_24294);
nor U25037 (N_25037,N_24695,N_24693);
nor U25038 (N_25038,N_24488,N_24598);
nor U25039 (N_25039,N_24376,N_24821);
or U25040 (N_25040,N_24886,N_24772);
or U25041 (N_25041,N_24079,N_24476);
and U25042 (N_25042,N_24670,N_24733);
or U25043 (N_25043,N_24776,N_24450);
or U25044 (N_25044,N_24106,N_24029);
nor U25045 (N_25045,N_24893,N_24407);
xnor U25046 (N_25046,N_24216,N_24814);
xnor U25047 (N_25047,N_24775,N_24849);
or U25048 (N_25048,N_24185,N_24825);
nand U25049 (N_25049,N_24262,N_24224);
nor U25050 (N_25050,N_24118,N_24610);
nand U25051 (N_25051,N_24806,N_24230);
nor U25052 (N_25052,N_24510,N_24059);
xor U25053 (N_25053,N_24140,N_24474);
nand U25054 (N_25054,N_24640,N_24154);
nand U25055 (N_25055,N_24323,N_24860);
xor U25056 (N_25056,N_24927,N_24740);
nand U25057 (N_25057,N_24671,N_24536);
xnor U25058 (N_25058,N_24265,N_24951);
or U25059 (N_25059,N_24850,N_24451);
and U25060 (N_25060,N_24659,N_24960);
and U25061 (N_25061,N_24961,N_24848);
xnor U25062 (N_25062,N_24971,N_24604);
xor U25063 (N_25063,N_24491,N_24603);
or U25064 (N_25064,N_24657,N_24487);
or U25065 (N_25065,N_24091,N_24665);
nand U25066 (N_25066,N_24792,N_24897);
and U25067 (N_25067,N_24003,N_24007);
nand U25068 (N_25068,N_24354,N_24006);
nand U25069 (N_25069,N_24633,N_24215);
nor U25070 (N_25070,N_24949,N_24172);
nand U25071 (N_25071,N_24000,N_24084);
and U25072 (N_25072,N_24757,N_24465);
and U25073 (N_25073,N_24749,N_24532);
nand U25074 (N_25074,N_24877,N_24570);
and U25075 (N_25075,N_24947,N_24590);
and U25076 (N_25076,N_24094,N_24307);
nand U25077 (N_25077,N_24857,N_24941);
nand U25078 (N_25078,N_24129,N_24716);
xnor U25079 (N_25079,N_24655,N_24372);
nor U25080 (N_25080,N_24746,N_24405);
nor U25081 (N_25081,N_24074,N_24165);
or U25082 (N_25082,N_24067,N_24589);
nand U25083 (N_25083,N_24542,N_24641);
nor U25084 (N_25084,N_24470,N_24446);
xor U25085 (N_25085,N_24082,N_24368);
xnor U25086 (N_25086,N_24321,N_24448);
xor U25087 (N_25087,N_24876,N_24312);
nand U25088 (N_25088,N_24358,N_24841);
and U25089 (N_25089,N_24192,N_24364);
xor U25090 (N_25090,N_24182,N_24092);
nand U25091 (N_25091,N_24497,N_24462);
xnor U25092 (N_25092,N_24612,N_24001);
nor U25093 (N_25093,N_24791,N_24296);
nor U25094 (N_25094,N_24564,N_24900);
or U25095 (N_25095,N_24469,N_24471);
nand U25096 (N_25096,N_24546,N_24235);
nor U25097 (N_25097,N_24763,N_24466);
nand U25098 (N_25098,N_24204,N_24226);
nor U25099 (N_25099,N_24583,N_24178);
or U25100 (N_25100,N_24188,N_24447);
xor U25101 (N_25101,N_24558,N_24514);
and U25102 (N_25102,N_24480,N_24395);
nor U25103 (N_25103,N_24018,N_24143);
or U25104 (N_25104,N_24501,N_24855);
or U25105 (N_25105,N_24948,N_24708);
xor U25106 (N_25106,N_24828,N_24797);
nor U25107 (N_25107,N_24962,N_24525);
nand U25108 (N_25108,N_24310,N_24910);
and U25109 (N_25109,N_24424,N_24380);
or U25110 (N_25110,N_24909,N_24254);
and U25111 (N_25111,N_24195,N_24113);
nand U25112 (N_25112,N_24517,N_24736);
xnor U25113 (N_25113,N_24631,N_24766);
or U25114 (N_25114,N_24712,N_24915);
nand U25115 (N_25115,N_24452,N_24913);
nand U25116 (N_25116,N_24015,N_24575);
nand U25117 (N_25117,N_24556,N_24073);
nor U25118 (N_25118,N_24731,N_24315);
xnor U25119 (N_25119,N_24174,N_24439);
nor U25120 (N_25120,N_24115,N_24186);
and U25121 (N_25121,N_24365,N_24979);
xor U25122 (N_25122,N_24618,N_24959);
nand U25123 (N_25123,N_24329,N_24387);
or U25124 (N_25124,N_24933,N_24157);
nand U25125 (N_25125,N_24403,N_24754);
xor U25126 (N_25126,N_24730,N_24954);
or U25127 (N_25127,N_24433,N_24654);
nand U25128 (N_25128,N_24786,N_24410);
xor U25129 (N_25129,N_24161,N_24972);
xnor U25130 (N_25130,N_24184,N_24152);
xnor U25131 (N_25131,N_24997,N_24173);
and U25132 (N_25132,N_24225,N_24114);
xor U25133 (N_25133,N_24685,N_24862);
and U25134 (N_25134,N_24503,N_24704);
nand U25135 (N_25135,N_24229,N_24021);
nor U25136 (N_25136,N_24861,N_24127);
nor U25137 (N_25137,N_24158,N_24179);
and U25138 (N_25138,N_24033,N_24858);
and U25139 (N_25139,N_24697,N_24617);
and U25140 (N_25140,N_24903,N_24978);
xor U25141 (N_25141,N_24788,N_24406);
nand U25142 (N_25142,N_24098,N_24946);
nor U25143 (N_25143,N_24944,N_24112);
and U25144 (N_25144,N_24574,N_24313);
xor U25145 (N_25145,N_24551,N_24534);
xor U25146 (N_25146,N_24982,N_24236);
and U25147 (N_25147,N_24203,N_24468);
nand U25148 (N_25148,N_24649,N_24048);
xor U25149 (N_25149,N_24602,N_24969);
and U25150 (N_25150,N_24014,N_24819);
xor U25151 (N_25151,N_24170,N_24461);
nor U25152 (N_25152,N_24484,N_24168);
and U25153 (N_25153,N_24726,N_24499);
and U25154 (N_25154,N_24557,N_24164);
nand U25155 (N_25155,N_24568,N_24481);
and U25156 (N_25156,N_24686,N_24581);
nor U25157 (N_25157,N_24995,N_24263);
or U25158 (N_25158,N_24402,N_24764);
and U25159 (N_25159,N_24989,N_24725);
or U25160 (N_25160,N_24264,N_24327);
and U25161 (N_25161,N_24413,N_24832);
nor U25162 (N_25162,N_24991,N_24269);
nand U25163 (N_25163,N_24076,N_24929);
nand U25164 (N_25164,N_24824,N_24386);
nand U25165 (N_25165,N_24777,N_24679);
or U25166 (N_25166,N_24055,N_24023);
nor U25167 (N_25167,N_24249,N_24240);
or U25168 (N_25168,N_24587,N_24613);
or U25169 (N_25169,N_24529,N_24227);
nor U25170 (N_25170,N_24477,N_24658);
nor U25171 (N_25171,N_24986,N_24316);
or U25172 (N_25172,N_24219,N_24911);
and U25173 (N_25173,N_24317,N_24629);
and U25174 (N_25174,N_24438,N_24734);
nor U25175 (N_25175,N_24647,N_24921);
and U25176 (N_25176,N_24136,N_24637);
nor U25177 (N_25177,N_24258,N_24445);
nand U25178 (N_25178,N_24537,N_24046);
or U25179 (N_25179,N_24099,N_24702);
or U25180 (N_25180,N_24706,N_24159);
xnor U25181 (N_25181,N_24722,N_24282);
nand U25182 (N_25182,N_24081,N_24668);
xor U25183 (N_25183,N_24759,N_24753);
and U25184 (N_25184,N_24632,N_24210);
or U25185 (N_25185,N_24751,N_24482);
xnor U25186 (N_25186,N_24520,N_24802);
or U25187 (N_25187,N_24412,N_24576);
xor U25188 (N_25188,N_24349,N_24701);
and U25189 (N_25189,N_24459,N_24769);
xnor U25190 (N_25190,N_24890,N_24284);
and U25191 (N_25191,N_24765,N_24648);
nand U25192 (N_25192,N_24332,N_24075);
or U25193 (N_25193,N_24398,N_24247);
nand U25194 (N_25194,N_24882,N_24856);
and U25195 (N_25195,N_24360,N_24155);
xor U25196 (N_25196,N_24677,N_24126);
xnor U25197 (N_25197,N_24884,N_24634);
and U25198 (N_25198,N_24418,N_24005);
and U25199 (N_25199,N_24518,N_24024);
nor U25200 (N_25200,N_24383,N_24382);
or U25201 (N_25201,N_24965,N_24901);
nand U25202 (N_25202,N_24371,N_24276);
and U25203 (N_25203,N_24506,N_24153);
xnor U25204 (N_25204,N_24928,N_24943);
xor U25205 (N_25205,N_24885,N_24270);
nor U25206 (N_25206,N_24286,N_24116);
and U25207 (N_25207,N_24580,N_24758);
nor U25208 (N_25208,N_24285,N_24826);
nand U25209 (N_25209,N_24783,N_24220);
and U25210 (N_25210,N_24086,N_24346);
and U25211 (N_25211,N_24243,N_24920);
or U25212 (N_25212,N_24070,N_24588);
xor U25213 (N_25213,N_24069,N_24690);
nand U25214 (N_25214,N_24401,N_24871);
nor U25215 (N_25215,N_24472,N_24801);
xor U25216 (N_25216,N_24895,N_24109);
nor U25217 (N_25217,N_24778,N_24146);
and U25218 (N_25218,N_24297,N_24680);
and U25219 (N_25219,N_24879,N_24837);
nor U25220 (N_25220,N_24111,N_24293);
xnor U25221 (N_25221,N_24718,N_24974);
nor U25222 (N_25222,N_24331,N_24038);
nor U25223 (N_25223,N_24952,N_24274);
nor U25224 (N_25224,N_24653,N_24483);
and U25225 (N_25225,N_24060,N_24275);
nor U25226 (N_25226,N_24966,N_24205);
nand U25227 (N_25227,N_24696,N_24020);
nor U25228 (N_25228,N_24427,N_24611);
and U25229 (N_25229,N_24530,N_24592);
or U25230 (N_25230,N_24102,N_24266);
nand U25231 (N_25231,N_24429,N_24540);
nor U25232 (N_25232,N_24739,N_24362);
nand U25233 (N_25233,N_24430,N_24381);
xnor U25234 (N_25234,N_24566,N_24496);
or U25235 (N_25235,N_24422,N_24077);
and U25236 (N_25236,N_24123,N_24149);
and U25237 (N_25237,N_24756,N_24976);
nand U25238 (N_25238,N_24097,N_24892);
nor U25239 (N_25239,N_24088,N_24200);
nor U25240 (N_25240,N_24498,N_24584);
and U25241 (N_25241,N_24311,N_24635);
nand U25242 (N_25242,N_24132,N_24388);
nand U25243 (N_25243,N_24615,N_24605);
and U25244 (N_25244,N_24507,N_24515);
nor U25245 (N_25245,N_24348,N_24934);
nand U25246 (N_25246,N_24950,N_24586);
or U25247 (N_25247,N_24793,N_24710);
xnor U25248 (N_25248,N_24125,N_24298);
and U25249 (N_25249,N_24223,N_24087);
and U25250 (N_25250,N_24083,N_24139);
nor U25251 (N_25251,N_24538,N_24500);
nor U25252 (N_25252,N_24134,N_24341);
and U25253 (N_25253,N_24443,N_24970);
nor U25254 (N_25254,N_24355,N_24594);
xnor U25255 (N_25255,N_24964,N_24460);
nor U25256 (N_25256,N_24867,N_24217);
or U25257 (N_25257,N_24745,N_24812);
xnor U25258 (N_25258,N_24423,N_24998);
nor U25259 (N_25259,N_24177,N_24539);
xor U25260 (N_25260,N_24441,N_24044);
or U25261 (N_25261,N_24508,N_24531);
nor U25262 (N_25262,N_24868,N_24350);
or U25263 (N_25263,N_24554,N_24727);
nor U25264 (N_25264,N_24790,N_24009);
nor U25265 (N_25265,N_24444,N_24805);
nor U25266 (N_25266,N_24620,N_24207);
nand U25267 (N_25267,N_24804,N_24032);
nand U25268 (N_25268,N_24419,N_24417);
nand U25269 (N_25269,N_24241,N_24063);
nand U25270 (N_25270,N_24148,N_24359);
and U25271 (N_25271,N_24743,N_24373);
xor U25272 (N_25272,N_24031,N_24627);
and U25273 (N_25273,N_24682,N_24011);
nand U25274 (N_25274,N_24672,N_24926);
nand U25275 (N_25275,N_24356,N_24278);
xor U25276 (N_25276,N_24822,N_24002);
and U25277 (N_25277,N_24923,N_24919);
and U25278 (N_25278,N_24408,N_24956);
or U25279 (N_25279,N_24958,N_24521);
or U25280 (N_25280,N_24261,N_24068);
or U25281 (N_25281,N_24435,N_24492);
nand U25282 (N_25282,N_24287,N_24160);
or U25283 (N_25283,N_24700,N_24251);
nor U25284 (N_25284,N_24963,N_24827);
nor U25285 (N_25285,N_24122,N_24357);
and U25286 (N_25286,N_24898,N_24541);
nor U25287 (N_25287,N_24522,N_24809);
nand U25288 (N_25288,N_24870,N_24673);
and U25289 (N_25289,N_24985,N_24295);
xnor U25290 (N_25290,N_24457,N_24117);
or U25291 (N_25291,N_24051,N_24569);
nor U25292 (N_25292,N_24524,N_24544);
nor U25293 (N_25293,N_24973,N_24720);
nand U25294 (N_25294,N_24645,N_24669);
or U25295 (N_25295,N_24085,N_24945);
nand U25296 (N_25296,N_24176,N_24596);
xnor U25297 (N_25297,N_24509,N_24523);
nor U25298 (N_25298,N_24782,N_24957);
nand U25299 (N_25299,N_24370,N_24660);
or U25300 (N_25300,N_24916,N_24794);
xor U25301 (N_25301,N_24400,N_24840);
nor U25302 (N_25302,N_24426,N_24464);
nor U25303 (N_25303,N_24244,N_24454);
nand U25304 (N_25304,N_24415,N_24684);
nor U25305 (N_25305,N_24343,N_24212);
and U25306 (N_25306,N_24428,N_24090);
and U25307 (N_25307,N_24361,N_24337);
and U25308 (N_25308,N_24990,N_24548);
xnor U25309 (N_25309,N_24728,N_24290);
nand U25310 (N_25310,N_24744,N_24260);
xnor U25311 (N_25311,N_24820,N_24624);
or U25312 (N_25312,N_24646,N_24065);
nand U25313 (N_25313,N_24238,N_24340);
or U25314 (N_25314,N_24456,N_24233);
and U25315 (N_25315,N_24560,N_24209);
or U25316 (N_25316,N_24411,N_24888);
xnor U25317 (N_25317,N_24213,N_24246);
nor U25318 (N_25318,N_24232,N_24839);
nor U25319 (N_25319,N_24585,N_24891);
nand U25320 (N_25320,N_24432,N_24028);
xor U25321 (N_25321,N_24664,N_24742);
nand U25322 (N_25322,N_24449,N_24255);
xor U25323 (N_25323,N_24908,N_24342);
nand U25324 (N_25324,N_24931,N_24938);
xor U25325 (N_25325,N_24768,N_24397);
or U25326 (N_25326,N_24818,N_24519);
or U25327 (N_25327,N_24442,N_24306);
and U25328 (N_25328,N_24054,N_24512);
nand U25329 (N_25329,N_24105,N_24936);
nand U25330 (N_25330,N_24683,N_24156);
xnor U25331 (N_25331,N_24463,N_24393);
nor U25332 (N_25332,N_24881,N_24846);
and U25333 (N_25333,N_24390,N_24338);
or U25334 (N_25334,N_24301,N_24131);
xnor U25335 (N_25335,N_24579,N_24345);
xor U25336 (N_25336,N_24218,N_24843);
xor U25337 (N_25337,N_24833,N_24875);
xnor U25338 (N_25338,N_24907,N_24277);
or U25339 (N_25339,N_24072,N_24080);
and U25340 (N_25340,N_24636,N_24019);
and U25341 (N_25341,N_24404,N_24562);
nand U25342 (N_25342,N_24779,N_24661);
nor U25343 (N_25343,N_24353,N_24479);
nand U25344 (N_25344,N_24473,N_24914);
and U25345 (N_25345,N_24351,N_24193);
xor U25346 (N_25346,N_24291,N_24108);
xor U25347 (N_25347,N_24609,N_24511);
nor U25348 (N_25348,N_24513,N_24707);
or U25349 (N_25349,N_24567,N_24721);
and U25350 (N_25350,N_24344,N_24656);
or U25351 (N_25351,N_24939,N_24968);
nand U25352 (N_25352,N_24859,N_24101);
xnor U25353 (N_25353,N_24810,N_24256);
xor U25354 (N_25354,N_24942,N_24169);
nand U25355 (N_25355,N_24593,N_24495);
xnor U25356 (N_25356,N_24851,N_24561);
and U25357 (N_25357,N_24741,N_24042);
nor U25358 (N_25358,N_24289,N_24626);
nor U25359 (N_25359,N_24250,N_24925);
or U25360 (N_25360,N_24550,N_24694);
or U25361 (N_25361,N_24121,N_24729);
xnor U25362 (N_25362,N_24773,N_24993);
and U25363 (N_25363,N_24894,N_24389);
nand U25364 (N_25364,N_24367,N_24922);
and U25365 (N_25365,N_24896,N_24535);
nand U25366 (N_25366,N_24151,N_24279);
xnor U25367 (N_25367,N_24181,N_24874);
nor U25368 (N_25368,N_24008,N_24045);
and U25369 (N_25369,N_24394,N_24110);
xor U25370 (N_25370,N_24676,N_24221);
nand U25371 (N_25371,N_24789,N_24392);
and U25372 (N_25372,N_24211,N_24918);
nor U25373 (N_25373,N_24050,N_24999);
and U25374 (N_25374,N_24552,N_24135);
nand U25375 (N_25375,N_24137,N_24719);
nor U25376 (N_25376,N_24652,N_24391);
nand U25377 (N_25377,N_24052,N_24699);
or U25378 (N_25378,N_24267,N_24591);
xnor U25379 (N_25379,N_24724,N_24889);
xnor U25380 (N_25380,N_24163,N_24614);
nand U25381 (N_25381,N_24813,N_24863);
xnor U25382 (N_25382,N_24883,N_24760);
xor U25383 (N_25383,N_24533,N_24326);
and U25384 (N_25384,N_24198,N_24906);
or U25385 (N_25385,N_24816,N_24162);
nor U25386 (N_25386,N_24796,N_24010);
nor U25387 (N_25387,N_24320,N_24687);
nand U25388 (N_25388,N_24887,N_24303);
nor U25389 (N_25389,N_24300,N_24252);
or U25390 (N_25390,N_24994,N_24057);
nand U25391 (N_25391,N_24691,N_24490);
or U25392 (N_25392,N_24543,N_24606);
xor U25393 (N_25393,N_24049,N_24838);
nand U25394 (N_25394,N_24379,N_24774);
nand U25395 (N_25395,N_24651,N_24416);
xnor U25396 (N_25396,N_24977,N_24257);
nor U25397 (N_25397,N_24107,N_24899);
xor U25398 (N_25398,N_24573,N_24453);
nor U25399 (N_25399,N_24638,N_24191);
or U25400 (N_25400,N_24056,N_24831);
xnor U25401 (N_25401,N_24852,N_24363);
nor U25402 (N_25402,N_24692,N_24022);
xor U25403 (N_25403,N_24854,N_24242);
and U25404 (N_25404,N_24988,N_24281);
or U25405 (N_25405,N_24709,N_24715);
or U25406 (N_25406,N_24502,N_24674);
and U25407 (N_25407,N_24366,N_24066);
xnor U25408 (N_25408,N_24559,N_24528);
and U25409 (N_25409,N_24836,N_24489);
nor U25410 (N_25410,N_24180,N_24555);
or U25411 (N_25411,N_24142,N_24399);
nand U25412 (N_25412,N_24678,N_24795);
and U25413 (N_25413,N_24064,N_24639);
and U25414 (N_25414,N_24431,N_24034);
and U25415 (N_25415,N_24016,N_24516);
or U25416 (N_25416,N_24330,N_24434);
nand U25417 (N_25417,N_24737,N_24864);
xor U25418 (N_25418,N_24425,N_24784);
xor U25419 (N_25419,N_24421,N_24026);
or U25420 (N_25420,N_24845,N_24374);
nor U25421 (N_25421,N_24880,N_24248);
nor U25422 (N_25422,N_24040,N_24984);
nor U25423 (N_25423,N_24750,N_24667);
nand U25424 (N_25424,N_24231,N_24017);
or U25425 (N_25425,N_24062,N_24189);
xnor U25426 (N_25426,N_24770,N_24283);
xor U25427 (N_25427,N_24785,N_24352);
xnor U25428 (N_25428,N_24145,N_24030);
nor U25429 (N_25429,N_24675,N_24711);
nand U25430 (N_25430,N_24043,N_24807);
nor U25431 (N_25431,N_24004,N_24190);
nor U25432 (N_25432,N_24940,N_24622);
and U25433 (N_25433,N_24955,N_24187);
xnor U25434 (N_25434,N_24025,N_24713);
xnor U25435 (N_25435,N_24436,N_24799);
xor U25436 (N_25436,N_24339,N_24904);
nor U25437 (N_25437,N_24698,N_24504);
or U25438 (N_25438,N_24803,N_24748);
xnor U25439 (N_25439,N_24798,N_24314);
xnor U25440 (N_25440,N_24245,N_24917);
and U25441 (N_25441,N_24214,N_24201);
or U25442 (N_25442,N_24228,N_24752);
nor U25443 (N_25443,N_24829,N_24414);
or U25444 (N_25444,N_24037,N_24623);
or U25445 (N_25445,N_24420,N_24128);
nand U25446 (N_25446,N_24865,N_24475);
xor U25447 (N_25447,N_24239,N_24630);
nand U25448 (N_25448,N_24302,N_24378);
nor U25449 (N_25449,N_24571,N_24259);
and U25450 (N_25450,N_24662,N_24309);
or U25451 (N_25451,N_24175,N_24932);
nor U25452 (N_25452,N_24608,N_24409);
nand U25453 (N_25453,N_24047,N_24937);
nand U25454 (N_25454,N_24305,N_24071);
and U25455 (N_25455,N_24319,N_24103);
nand U25456 (N_25456,N_24787,N_24732);
nor U25457 (N_25457,N_24396,N_24992);
or U25458 (N_25458,N_24642,N_24755);
xnor U25459 (N_25459,N_24878,N_24866);
nor U25460 (N_25460,N_24607,N_24375);
nand U25461 (N_25461,N_24762,N_24553);
nand U25462 (N_25462,N_24100,N_24967);
nor U25463 (N_25463,N_24975,N_24253);
xnor U25464 (N_25464,N_24981,N_24616);
or U25465 (N_25465,N_24924,N_24485);
and U25466 (N_25466,N_24912,N_24526);
xor U25467 (N_25467,N_24222,N_24237);
or U25468 (N_25468,N_24206,N_24853);
or U25469 (N_25469,N_24377,N_24234);
xor U25470 (N_25470,N_24053,N_24578);
and U25471 (N_25471,N_24271,N_24847);
nor U25472 (N_25472,N_24800,N_24545);
nor U25473 (N_25473,N_24781,N_24304);
xnor U25474 (N_25474,N_24996,N_24983);
and U25475 (N_25475,N_24549,N_24385);
or U25476 (N_25476,N_24505,N_24027);
and U25477 (N_25477,N_24705,N_24703);
nand U25478 (N_25478,N_24723,N_24334);
or U25479 (N_25479,N_24120,N_24039);
nand U25480 (N_25480,N_24208,N_24689);
or U25481 (N_25481,N_24347,N_24171);
nor U25482 (N_25482,N_24124,N_24299);
nand U25483 (N_25483,N_24823,N_24150);
nand U25484 (N_25484,N_24980,N_24527);
and U25485 (N_25485,N_24714,N_24144);
and U25486 (N_25486,N_24688,N_24104);
and U25487 (N_25487,N_24644,N_24167);
xor U25488 (N_25488,N_24012,N_24035);
nand U25489 (N_25489,N_24292,N_24547);
xor U25490 (N_25490,N_24308,N_24869);
or U25491 (N_25491,N_24096,N_24873);
xnor U25492 (N_25492,N_24771,N_24811);
and U25493 (N_25493,N_24625,N_24599);
xnor U25494 (N_25494,N_24953,N_24041);
nor U25495 (N_25495,N_24650,N_24478);
or U25496 (N_25496,N_24268,N_24601);
and U25497 (N_25497,N_24196,N_24058);
xor U25498 (N_25498,N_24872,N_24036);
or U25499 (N_25499,N_24133,N_24183);
or U25500 (N_25500,N_24231,N_24883);
and U25501 (N_25501,N_24198,N_24938);
and U25502 (N_25502,N_24345,N_24731);
or U25503 (N_25503,N_24638,N_24824);
and U25504 (N_25504,N_24654,N_24803);
xnor U25505 (N_25505,N_24771,N_24386);
and U25506 (N_25506,N_24770,N_24878);
and U25507 (N_25507,N_24262,N_24666);
or U25508 (N_25508,N_24138,N_24755);
and U25509 (N_25509,N_24765,N_24088);
nand U25510 (N_25510,N_24158,N_24418);
or U25511 (N_25511,N_24720,N_24284);
xor U25512 (N_25512,N_24556,N_24185);
nand U25513 (N_25513,N_24802,N_24405);
xor U25514 (N_25514,N_24155,N_24525);
or U25515 (N_25515,N_24477,N_24931);
and U25516 (N_25516,N_24219,N_24567);
or U25517 (N_25517,N_24174,N_24656);
xor U25518 (N_25518,N_24386,N_24818);
and U25519 (N_25519,N_24846,N_24077);
nor U25520 (N_25520,N_24146,N_24722);
and U25521 (N_25521,N_24279,N_24676);
or U25522 (N_25522,N_24767,N_24750);
nor U25523 (N_25523,N_24741,N_24121);
nand U25524 (N_25524,N_24810,N_24918);
xor U25525 (N_25525,N_24045,N_24356);
xor U25526 (N_25526,N_24485,N_24540);
xnor U25527 (N_25527,N_24519,N_24138);
nand U25528 (N_25528,N_24542,N_24890);
or U25529 (N_25529,N_24151,N_24250);
or U25530 (N_25530,N_24407,N_24926);
nand U25531 (N_25531,N_24415,N_24287);
nand U25532 (N_25532,N_24468,N_24335);
and U25533 (N_25533,N_24283,N_24253);
or U25534 (N_25534,N_24572,N_24590);
and U25535 (N_25535,N_24869,N_24123);
nor U25536 (N_25536,N_24179,N_24000);
or U25537 (N_25537,N_24720,N_24968);
and U25538 (N_25538,N_24913,N_24540);
xor U25539 (N_25539,N_24208,N_24501);
and U25540 (N_25540,N_24220,N_24703);
nor U25541 (N_25541,N_24581,N_24299);
nand U25542 (N_25542,N_24760,N_24557);
nor U25543 (N_25543,N_24340,N_24874);
and U25544 (N_25544,N_24695,N_24691);
nor U25545 (N_25545,N_24555,N_24049);
nor U25546 (N_25546,N_24948,N_24620);
or U25547 (N_25547,N_24013,N_24700);
nor U25548 (N_25548,N_24378,N_24247);
or U25549 (N_25549,N_24880,N_24159);
nor U25550 (N_25550,N_24273,N_24868);
or U25551 (N_25551,N_24785,N_24271);
and U25552 (N_25552,N_24512,N_24677);
or U25553 (N_25553,N_24877,N_24373);
or U25554 (N_25554,N_24022,N_24341);
nor U25555 (N_25555,N_24321,N_24396);
nand U25556 (N_25556,N_24095,N_24492);
or U25557 (N_25557,N_24881,N_24315);
nand U25558 (N_25558,N_24562,N_24193);
and U25559 (N_25559,N_24106,N_24028);
xor U25560 (N_25560,N_24089,N_24578);
xnor U25561 (N_25561,N_24433,N_24841);
and U25562 (N_25562,N_24486,N_24805);
nand U25563 (N_25563,N_24233,N_24014);
or U25564 (N_25564,N_24247,N_24317);
nand U25565 (N_25565,N_24880,N_24202);
xor U25566 (N_25566,N_24369,N_24043);
and U25567 (N_25567,N_24048,N_24911);
and U25568 (N_25568,N_24280,N_24150);
nor U25569 (N_25569,N_24067,N_24057);
or U25570 (N_25570,N_24218,N_24528);
nor U25571 (N_25571,N_24726,N_24982);
nand U25572 (N_25572,N_24323,N_24395);
nor U25573 (N_25573,N_24093,N_24001);
xor U25574 (N_25574,N_24500,N_24061);
xor U25575 (N_25575,N_24044,N_24012);
or U25576 (N_25576,N_24583,N_24086);
or U25577 (N_25577,N_24133,N_24820);
nor U25578 (N_25578,N_24599,N_24461);
or U25579 (N_25579,N_24117,N_24467);
nand U25580 (N_25580,N_24549,N_24306);
xor U25581 (N_25581,N_24395,N_24661);
or U25582 (N_25582,N_24773,N_24984);
or U25583 (N_25583,N_24422,N_24737);
nand U25584 (N_25584,N_24696,N_24147);
nand U25585 (N_25585,N_24300,N_24956);
and U25586 (N_25586,N_24427,N_24360);
or U25587 (N_25587,N_24457,N_24887);
nor U25588 (N_25588,N_24506,N_24898);
nor U25589 (N_25589,N_24225,N_24603);
and U25590 (N_25590,N_24863,N_24613);
and U25591 (N_25591,N_24549,N_24429);
xnor U25592 (N_25592,N_24195,N_24197);
or U25593 (N_25593,N_24962,N_24676);
or U25594 (N_25594,N_24124,N_24186);
nor U25595 (N_25595,N_24492,N_24354);
nand U25596 (N_25596,N_24021,N_24594);
xor U25597 (N_25597,N_24037,N_24179);
nor U25598 (N_25598,N_24888,N_24192);
nor U25599 (N_25599,N_24940,N_24910);
and U25600 (N_25600,N_24474,N_24361);
nand U25601 (N_25601,N_24899,N_24509);
and U25602 (N_25602,N_24254,N_24788);
nor U25603 (N_25603,N_24098,N_24895);
nor U25604 (N_25604,N_24705,N_24874);
nor U25605 (N_25605,N_24629,N_24679);
nand U25606 (N_25606,N_24567,N_24944);
and U25607 (N_25607,N_24724,N_24152);
xnor U25608 (N_25608,N_24470,N_24699);
xor U25609 (N_25609,N_24938,N_24374);
and U25610 (N_25610,N_24402,N_24967);
nor U25611 (N_25611,N_24505,N_24538);
nand U25612 (N_25612,N_24379,N_24407);
xnor U25613 (N_25613,N_24610,N_24361);
nor U25614 (N_25614,N_24248,N_24684);
nand U25615 (N_25615,N_24191,N_24821);
and U25616 (N_25616,N_24361,N_24668);
and U25617 (N_25617,N_24971,N_24165);
or U25618 (N_25618,N_24097,N_24295);
and U25619 (N_25619,N_24822,N_24890);
nand U25620 (N_25620,N_24761,N_24770);
nand U25621 (N_25621,N_24134,N_24275);
nor U25622 (N_25622,N_24811,N_24094);
and U25623 (N_25623,N_24063,N_24986);
xnor U25624 (N_25624,N_24420,N_24510);
and U25625 (N_25625,N_24433,N_24777);
nor U25626 (N_25626,N_24287,N_24131);
nand U25627 (N_25627,N_24770,N_24440);
nor U25628 (N_25628,N_24795,N_24829);
nand U25629 (N_25629,N_24243,N_24513);
xor U25630 (N_25630,N_24968,N_24812);
nand U25631 (N_25631,N_24597,N_24218);
or U25632 (N_25632,N_24460,N_24795);
xor U25633 (N_25633,N_24332,N_24623);
and U25634 (N_25634,N_24337,N_24537);
or U25635 (N_25635,N_24694,N_24426);
or U25636 (N_25636,N_24871,N_24909);
nor U25637 (N_25637,N_24454,N_24843);
xor U25638 (N_25638,N_24492,N_24645);
or U25639 (N_25639,N_24373,N_24042);
nand U25640 (N_25640,N_24224,N_24031);
nand U25641 (N_25641,N_24527,N_24509);
or U25642 (N_25642,N_24337,N_24153);
nand U25643 (N_25643,N_24773,N_24713);
nand U25644 (N_25644,N_24643,N_24914);
nor U25645 (N_25645,N_24385,N_24859);
xor U25646 (N_25646,N_24003,N_24989);
nand U25647 (N_25647,N_24750,N_24575);
and U25648 (N_25648,N_24667,N_24021);
nand U25649 (N_25649,N_24156,N_24951);
nor U25650 (N_25650,N_24879,N_24644);
nor U25651 (N_25651,N_24295,N_24660);
or U25652 (N_25652,N_24343,N_24560);
nor U25653 (N_25653,N_24235,N_24933);
nor U25654 (N_25654,N_24606,N_24086);
nor U25655 (N_25655,N_24383,N_24375);
or U25656 (N_25656,N_24898,N_24250);
nor U25657 (N_25657,N_24481,N_24352);
xor U25658 (N_25658,N_24066,N_24311);
nor U25659 (N_25659,N_24908,N_24332);
and U25660 (N_25660,N_24920,N_24531);
nand U25661 (N_25661,N_24184,N_24115);
and U25662 (N_25662,N_24210,N_24387);
and U25663 (N_25663,N_24518,N_24979);
and U25664 (N_25664,N_24341,N_24782);
or U25665 (N_25665,N_24815,N_24035);
nand U25666 (N_25666,N_24981,N_24645);
xor U25667 (N_25667,N_24287,N_24701);
and U25668 (N_25668,N_24227,N_24257);
and U25669 (N_25669,N_24216,N_24018);
nand U25670 (N_25670,N_24471,N_24224);
and U25671 (N_25671,N_24773,N_24170);
nand U25672 (N_25672,N_24870,N_24629);
or U25673 (N_25673,N_24176,N_24895);
nor U25674 (N_25674,N_24452,N_24168);
nor U25675 (N_25675,N_24551,N_24139);
or U25676 (N_25676,N_24068,N_24353);
xor U25677 (N_25677,N_24873,N_24226);
nand U25678 (N_25678,N_24244,N_24431);
or U25679 (N_25679,N_24011,N_24436);
nand U25680 (N_25680,N_24686,N_24477);
nor U25681 (N_25681,N_24789,N_24198);
nor U25682 (N_25682,N_24500,N_24087);
or U25683 (N_25683,N_24304,N_24661);
and U25684 (N_25684,N_24173,N_24522);
or U25685 (N_25685,N_24730,N_24444);
or U25686 (N_25686,N_24541,N_24954);
or U25687 (N_25687,N_24863,N_24759);
or U25688 (N_25688,N_24189,N_24070);
and U25689 (N_25689,N_24817,N_24441);
or U25690 (N_25690,N_24147,N_24656);
or U25691 (N_25691,N_24346,N_24187);
and U25692 (N_25692,N_24154,N_24624);
and U25693 (N_25693,N_24459,N_24205);
and U25694 (N_25694,N_24691,N_24019);
xor U25695 (N_25695,N_24517,N_24107);
nand U25696 (N_25696,N_24506,N_24597);
xnor U25697 (N_25697,N_24343,N_24811);
and U25698 (N_25698,N_24385,N_24251);
nand U25699 (N_25699,N_24932,N_24868);
nor U25700 (N_25700,N_24419,N_24906);
or U25701 (N_25701,N_24190,N_24719);
xor U25702 (N_25702,N_24405,N_24851);
nor U25703 (N_25703,N_24021,N_24135);
nor U25704 (N_25704,N_24275,N_24992);
or U25705 (N_25705,N_24584,N_24384);
and U25706 (N_25706,N_24651,N_24500);
or U25707 (N_25707,N_24261,N_24009);
nand U25708 (N_25708,N_24282,N_24727);
nand U25709 (N_25709,N_24502,N_24185);
nor U25710 (N_25710,N_24095,N_24931);
nor U25711 (N_25711,N_24268,N_24939);
xor U25712 (N_25712,N_24764,N_24208);
and U25713 (N_25713,N_24629,N_24309);
or U25714 (N_25714,N_24242,N_24892);
or U25715 (N_25715,N_24475,N_24368);
or U25716 (N_25716,N_24371,N_24358);
nand U25717 (N_25717,N_24481,N_24686);
nand U25718 (N_25718,N_24047,N_24915);
nor U25719 (N_25719,N_24154,N_24133);
and U25720 (N_25720,N_24253,N_24060);
and U25721 (N_25721,N_24506,N_24312);
xnor U25722 (N_25722,N_24423,N_24487);
nand U25723 (N_25723,N_24648,N_24787);
xor U25724 (N_25724,N_24597,N_24414);
nand U25725 (N_25725,N_24505,N_24556);
xor U25726 (N_25726,N_24809,N_24811);
nand U25727 (N_25727,N_24129,N_24913);
xor U25728 (N_25728,N_24809,N_24833);
or U25729 (N_25729,N_24784,N_24645);
and U25730 (N_25730,N_24458,N_24512);
xnor U25731 (N_25731,N_24856,N_24755);
nand U25732 (N_25732,N_24812,N_24428);
or U25733 (N_25733,N_24155,N_24223);
or U25734 (N_25734,N_24118,N_24744);
nand U25735 (N_25735,N_24869,N_24233);
xor U25736 (N_25736,N_24481,N_24378);
nand U25737 (N_25737,N_24977,N_24246);
xor U25738 (N_25738,N_24870,N_24594);
xor U25739 (N_25739,N_24784,N_24514);
nand U25740 (N_25740,N_24989,N_24909);
and U25741 (N_25741,N_24176,N_24491);
and U25742 (N_25742,N_24237,N_24594);
nand U25743 (N_25743,N_24433,N_24811);
nand U25744 (N_25744,N_24737,N_24709);
nand U25745 (N_25745,N_24986,N_24963);
nor U25746 (N_25746,N_24924,N_24283);
or U25747 (N_25747,N_24649,N_24603);
and U25748 (N_25748,N_24091,N_24511);
nor U25749 (N_25749,N_24241,N_24574);
nand U25750 (N_25750,N_24726,N_24353);
nand U25751 (N_25751,N_24366,N_24069);
and U25752 (N_25752,N_24235,N_24668);
and U25753 (N_25753,N_24647,N_24934);
xnor U25754 (N_25754,N_24638,N_24954);
nand U25755 (N_25755,N_24169,N_24295);
xnor U25756 (N_25756,N_24094,N_24265);
or U25757 (N_25757,N_24698,N_24277);
xnor U25758 (N_25758,N_24651,N_24711);
or U25759 (N_25759,N_24845,N_24220);
nand U25760 (N_25760,N_24408,N_24034);
nand U25761 (N_25761,N_24013,N_24289);
xor U25762 (N_25762,N_24765,N_24353);
or U25763 (N_25763,N_24790,N_24629);
nand U25764 (N_25764,N_24648,N_24930);
or U25765 (N_25765,N_24219,N_24222);
nand U25766 (N_25766,N_24143,N_24211);
and U25767 (N_25767,N_24220,N_24641);
and U25768 (N_25768,N_24535,N_24345);
nor U25769 (N_25769,N_24837,N_24814);
nand U25770 (N_25770,N_24070,N_24693);
nand U25771 (N_25771,N_24432,N_24097);
and U25772 (N_25772,N_24753,N_24796);
nand U25773 (N_25773,N_24787,N_24991);
xor U25774 (N_25774,N_24140,N_24894);
or U25775 (N_25775,N_24903,N_24848);
nor U25776 (N_25776,N_24046,N_24751);
nor U25777 (N_25777,N_24956,N_24754);
nand U25778 (N_25778,N_24076,N_24307);
or U25779 (N_25779,N_24281,N_24594);
and U25780 (N_25780,N_24232,N_24113);
and U25781 (N_25781,N_24632,N_24165);
or U25782 (N_25782,N_24478,N_24356);
nand U25783 (N_25783,N_24588,N_24146);
xnor U25784 (N_25784,N_24028,N_24192);
xnor U25785 (N_25785,N_24287,N_24733);
xor U25786 (N_25786,N_24465,N_24925);
and U25787 (N_25787,N_24097,N_24481);
or U25788 (N_25788,N_24932,N_24538);
xnor U25789 (N_25789,N_24859,N_24004);
nor U25790 (N_25790,N_24276,N_24742);
nor U25791 (N_25791,N_24022,N_24666);
nand U25792 (N_25792,N_24823,N_24807);
xor U25793 (N_25793,N_24974,N_24480);
nor U25794 (N_25794,N_24521,N_24419);
or U25795 (N_25795,N_24952,N_24494);
nor U25796 (N_25796,N_24130,N_24657);
nand U25797 (N_25797,N_24392,N_24015);
nand U25798 (N_25798,N_24846,N_24398);
nand U25799 (N_25799,N_24868,N_24271);
and U25800 (N_25800,N_24569,N_24952);
nor U25801 (N_25801,N_24895,N_24906);
and U25802 (N_25802,N_24975,N_24431);
nor U25803 (N_25803,N_24428,N_24477);
nand U25804 (N_25804,N_24048,N_24900);
nand U25805 (N_25805,N_24713,N_24051);
nand U25806 (N_25806,N_24024,N_24751);
or U25807 (N_25807,N_24150,N_24730);
and U25808 (N_25808,N_24609,N_24556);
xnor U25809 (N_25809,N_24681,N_24057);
or U25810 (N_25810,N_24734,N_24502);
or U25811 (N_25811,N_24153,N_24046);
nor U25812 (N_25812,N_24225,N_24011);
or U25813 (N_25813,N_24375,N_24379);
or U25814 (N_25814,N_24764,N_24822);
xnor U25815 (N_25815,N_24733,N_24251);
nor U25816 (N_25816,N_24622,N_24633);
and U25817 (N_25817,N_24164,N_24644);
or U25818 (N_25818,N_24003,N_24159);
nand U25819 (N_25819,N_24497,N_24505);
nor U25820 (N_25820,N_24785,N_24884);
or U25821 (N_25821,N_24433,N_24839);
or U25822 (N_25822,N_24673,N_24515);
nor U25823 (N_25823,N_24650,N_24177);
xor U25824 (N_25824,N_24846,N_24861);
or U25825 (N_25825,N_24206,N_24987);
xor U25826 (N_25826,N_24762,N_24622);
nand U25827 (N_25827,N_24723,N_24410);
and U25828 (N_25828,N_24778,N_24403);
nor U25829 (N_25829,N_24532,N_24638);
or U25830 (N_25830,N_24693,N_24439);
nor U25831 (N_25831,N_24185,N_24482);
nor U25832 (N_25832,N_24596,N_24872);
nand U25833 (N_25833,N_24331,N_24173);
nand U25834 (N_25834,N_24464,N_24539);
or U25835 (N_25835,N_24042,N_24123);
or U25836 (N_25836,N_24738,N_24015);
or U25837 (N_25837,N_24776,N_24970);
nand U25838 (N_25838,N_24536,N_24846);
or U25839 (N_25839,N_24537,N_24622);
or U25840 (N_25840,N_24976,N_24179);
nand U25841 (N_25841,N_24987,N_24508);
nor U25842 (N_25842,N_24756,N_24571);
nand U25843 (N_25843,N_24991,N_24534);
or U25844 (N_25844,N_24101,N_24861);
and U25845 (N_25845,N_24775,N_24111);
or U25846 (N_25846,N_24169,N_24446);
xor U25847 (N_25847,N_24888,N_24332);
nand U25848 (N_25848,N_24920,N_24225);
and U25849 (N_25849,N_24279,N_24005);
nor U25850 (N_25850,N_24923,N_24465);
xnor U25851 (N_25851,N_24340,N_24781);
nand U25852 (N_25852,N_24240,N_24949);
xor U25853 (N_25853,N_24222,N_24939);
or U25854 (N_25854,N_24022,N_24086);
nor U25855 (N_25855,N_24598,N_24753);
nor U25856 (N_25856,N_24473,N_24604);
nor U25857 (N_25857,N_24361,N_24243);
or U25858 (N_25858,N_24848,N_24745);
nor U25859 (N_25859,N_24000,N_24075);
xnor U25860 (N_25860,N_24940,N_24265);
or U25861 (N_25861,N_24311,N_24852);
xor U25862 (N_25862,N_24662,N_24013);
nor U25863 (N_25863,N_24740,N_24010);
or U25864 (N_25864,N_24815,N_24721);
or U25865 (N_25865,N_24677,N_24900);
nand U25866 (N_25866,N_24033,N_24121);
or U25867 (N_25867,N_24970,N_24676);
and U25868 (N_25868,N_24170,N_24150);
and U25869 (N_25869,N_24667,N_24264);
nand U25870 (N_25870,N_24982,N_24359);
and U25871 (N_25871,N_24532,N_24122);
nor U25872 (N_25872,N_24702,N_24225);
and U25873 (N_25873,N_24397,N_24338);
xnor U25874 (N_25874,N_24463,N_24806);
xor U25875 (N_25875,N_24527,N_24876);
and U25876 (N_25876,N_24152,N_24883);
nand U25877 (N_25877,N_24183,N_24726);
nand U25878 (N_25878,N_24403,N_24087);
nor U25879 (N_25879,N_24484,N_24375);
and U25880 (N_25880,N_24505,N_24946);
xor U25881 (N_25881,N_24062,N_24713);
nor U25882 (N_25882,N_24229,N_24528);
nand U25883 (N_25883,N_24178,N_24833);
xor U25884 (N_25884,N_24129,N_24636);
and U25885 (N_25885,N_24624,N_24360);
and U25886 (N_25886,N_24522,N_24655);
nor U25887 (N_25887,N_24371,N_24873);
or U25888 (N_25888,N_24402,N_24413);
nand U25889 (N_25889,N_24259,N_24509);
nor U25890 (N_25890,N_24987,N_24829);
or U25891 (N_25891,N_24191,N_24145);
and U25892 (N_25892,N_24624,N_24850);
nand U25893 (N_25893,N_24810,N_24007);
nor U25894 (N_25894,N_24308,N_24488);
nand U25895 (N_25895,N_24010,N_24224);
nor U25896 (N_25896,N_24646,N_24167);
and U25897 (N_25897,N_24312,N_24954);
xor U25898 (N_25898,N_24339,N_24816);
and U25899 (N_25899,N_24214,N_24266);
nand U25900 (N_25900,N_24078,N_24161);
nand U25901 (N_25901,N_24678,N_24408);
and U25902 (N_25902,N_24045,N_24661);
xor U25903 (N_25903,N_24754,N_24428);
and U25904 (N_25904,N_24822,N_24768);
nor U25905 (N_25905,N_24689,N_24674);
or U25906 (N_25906,N_24134,N_24533);
xor U25907 (N_25907,N_24312,N_24409);
nand U25908 (N_25908,N_24595,N_24242);
nor U25909 (N_25909,N_24262,N_24163);
or U25910 (N_25910,N_24466,N_24745);
nand U25911 (N_25911,N_24198,N_24411);
and U25912 (N_25912,N_24017,N_24700);
or U25913 (N_25913,N_24883,N_24570);
and U25914 (N_25914,N_24330,N_24798);
xor U25915 (N_25915,N_24849,N_24413);
and U25916 (N_25916,N_24789,N_24847);
xnor U25917 (N_25917,N_24889,N_24349);
xnor U25918 (N_25918,N_24265,N_24113);
or U25919 (N_25919,N_24679,N_24542);
and U25920 (N_25920,N_24956,N_24595);
or U25921 (N_25921,N_24088,N_24300);
and U25922 (N_25922,N_24016,N_24957);
nand U25923 (N_25923,N_24725,N_24850);
nor U25924 (N_25924,N_24849,N_24891);
or U25925 (N_25925,N_24769,N_24187);
and U25926 (N_25926,N_24251,N_24445);
or U25927 (N_25927,N_24785,N_24395);
or U25928 (N_25928,N_24433,N_24992);
xnor U25929 (N_25929,N_24230,N_24738);
xor U25930 (N_25930,N_24208,N_24084);
xor U25931 (N_25931,N_24376,N_24060);
nand U25932 (N_25932,N_24499,N_24663);
and U25933 (N_25933,N_24134,N_24543);
or U25934 (N_25934,N_24521,N_24760);
and U25935 (N_25935,N_24230,N_24716);
nand U25936 (N_25936,N_24044,N_24150);
or U25937 (N_25937,N_24517,N_24609);
nand U25938 (N_25938,N_24884,N_24903);
nand U25939 (N_25939,N_24197,N_24346);
and U25940 (N_25940,N_24229,N_24712);
or U25941 (N_25941,N_24588,N_24528);
nor U25942 (N_25942,N_24488,N_24932);
nand U25943 (N_25943,N_24473,N_24257);
and U25944 (N_25944,N_24639,N_24559);
nand U25945 (N_25945,N_24819,N_24898);
xor U25946 (N_25946,N_24979,N_24895);
and U25947 (N_25947,N_24197,N_24137);
nand U25948 (N_25948,N_24795,N_24307);
xnor U25949 (N_25949,N_24906,N_24095);
or U25950 (N_25950,N_24471,N_24974);
nor U25951 (N_25951,N_24164,N_24667);
nand U25952 (N_25952,N_24487,N_24715);
xnor U25953 (N_25953,N_24846,N_24848);
nor U25954 (N_25954,N_24336,N_24604);
or U25955 (N_25955,N_24703,N_24924);
nand U25956 (N_25956,N_24339,N_24218);
nor U25957 (N_25957,N_24844,N_24606);
xnor U25958 (N_25958,N_24160,N_24633);
or U25959 (N_25959,N_24039,N_24692);
xor U25960 (N_25960,N_24304,N_24749);
nor U25961 (N_25961,N_24000,N_24214);
nand U25962 (N_25962,N_24758,N_24003);
xor U25963 (N_25963,N_24078,N_24609);
nor U25964 (N_25964,N_24215,N_24620);
xnor U25965 (N_25965,N_24051,N_24256);
nor U25966 (N_25966,N_24267,N_24118);
or U25967 (N_25967,N_24677,N_24198);
and U25968 (N_25968,N_24555,N_24237);
nor U25969 (N_25969,N_24867,N_24625);
and U25970 (N_25970,N_24278,N_24627);
xnor U25971 (N_25971,N_24556,N_24975);
xnor U25972 (N_25972,N_24491,N_24943);
or U25973 (N_25973,N_24775,N_24797);
nand U25974 (N_25974,N_24164,N_24697);
nand U25975 (N_25975,N_24523,N_24116);
or U25976 (N_25976,N_24566,N_24061);
or U25977 (N_25977,N_24479,N_24416);
or U25978 (N_25978,N_24286,N_24205);
and U25979 (N_25979,N_24455,N_24335);
xnor U25980 (N_25980,N_24766,N_24557);
and U25981 (N_25981,N_24731,N_24486);
and U25982 (N_25982,N_24057,N_24592);
nand U25983 (N_25983,N_24745,N_24681);
and U25984 (N_25984,N_24417,N_24185);
or U25985 (N_25985,N_24442,N_24985);
and U25986 (N_25986,N_24328,N_24719);
xnor U25987 (N_25987,N_24716,N_24145);
xor U25988 (N_25988,N_24000,N_24840);
or U25989 (N_25989,N_24883,N_24415);
nor U25990 (N_25990,N_24567,N_24669);
nor U25991 (N_25991,N_24703,N_24142);
nor U25992 (N_25992,N_24196,N_24733);
nand U25993 (N_25993,N_24331,N_24623);
xor U25994 (N_25994,N_24505,N_24975);
or U25995 (N_25995,N_24727,N_24156);
xor U25996 (N_25996,N_24833,N_24647);
xnor U25997 (N_25997,N_24826,N_24744);
nor U25998 (N_25998,N_24211,N_24345);
and U25999 (N_25999,N_24130,N_24587);
xnor U26000 (N_26000,N_25049,N_25296);
nor U26001 (N_26001,N_25860,N_25289);
xnor U26002 (N_26002,N_25500,N_25398);
xor U26003 (N_26003,N_25630,N_25275);
and U26004 (N_26004,N_25664,N_25827);
nor U26005 (N_26005,N_25897,N_25667);
nor U26006 (N_26006,N_25358,N_25681);
nor U26007 (N_26007,N_25817,N_25937);
and U26008 (N_26008,N_25163,N_25910);
nor U26009 (N_26009,N_25976,N_25766);
xnor U26010 (N_26010,N_25890,N_25438);
and U26011 (N_26011,N_25613,N_25226);
and U26012 (N_26012,N_25521,N_25487);
or U26013 (N_26013,N_25559,N_25673);
or U26014 (N_26014,N_25599,N_25370);
or U26015 (N_26015,N_25765,N_25182);
xor U26016 (N_26016,N_25381,N_25669);
nor U26017 (N_26017,N_25116,N_25084);
and U26018 (N_26018,N_25379,N_25479);
nand U26019 (N_26019,N_25456,N_25792);
nand U26020 (N_26020,N_25421,N_25045);
nand U26021 (N_26021,N_25187,N_25899);
nor U26022 (N_26022,N_25790,N_25248);
and U26023 (N_26023,N_25231,N_25811);
nor U26024 (N_26024,N_25822,N_25861);
and U26025 (N_26025,N_25682,N_25198);
or U26026 (N_26026,N_25623,N_25193);
nor U26027 (N_26027,N_25697,N_25680);
and U26028 (N_26028,N_25570,N_25507);
and U26029 (N_26029,N_25747,N_25905);
or U26030 (N_26030,N_25262,N_25945);
nor U26031 (N_26031,N_25484,N_25033);
nand U26032 (N_26032,N_25843,N_25459);
and U26033 (N_26033,N_25314,N_25646);
and U26034 (N_26034,N_25213,N_25183);
nor U26035 (N_26035,N_25549,N_25395);
nand U26036 (N_26036,N_25350,N_25263);
nor U26037 (N_26037,N_25956,N_25810);
xnor U26038 (N_26038,N_25533,N_25875);
nor U26039 (N_26039,N_25424,N_25752);
nand U26040 (N_26040,N_25774,N_25031);
or U26041 (N_26041,N_25057,N_25287);
nand U26042 (N_26042,N_25058,N_25399);
or U26043 (N_26043,N_25684,N_25706);
xor U26044 (N_26044,N_25809,N_25329);
or U26045 (N_26045,N_25118,N_25064);
or U26046 (N_26046,N_25857,N_25082);
or U26047 (N_26047,N_25908,N_25126);
xor U26048 (N_26048,N_25659,N_25631);
xor U26049 (N_26049,N_25292,N_25089);
xor U26050 (N_26050,N_25010,N_25526);
xnor U26051 (N_26051,N_25284,N_25462);
xnor U26052 (N_26052,N_25216,N_25018);
nor U26053 (N_26053,N_25728,N_25607);
nor U26054 (N_26054,N_25083,N_25217);
and U26055 (N_26055,N_25471,N_25420);
or U26056 (N_26056,N_25334,N_25678);
nand U26057 (N_26057,N_25628,N_25553);
nor U26058 (N_26058,N_25565,N_25230);
nor U26059 (N_26059,N_25796,N_25577);
nand U26060 (N_26060,N_25436,N_25944);
xnor U26061 (N_26061,N_25994,N_25611);
and U26062 (N_26062,N_25940,N_25692);
nor U26063 (N_26063,N_25693,N_25404);
nand U26064 (N_26064,N_25191,N_25483);
nand U26065 (N_26065,N_25541,N_25992);
nand U26066 (N_26066,N_25584,N_25236);
and U26067 (N_26067,N_25000,N_25759);
xnor U26068 (N_26068,N_25786,N_25925);
xor U26069 (N_26069,N_25167,N_25982);
or U26070 (N_26070,N_25297,N_25390);
nand U26071 (N_26071,N_25281,N_25699);
nor U26072 (N_26072,N_25952,N_25301);
nand U26073 (N_26073,N_25209,N_25917);
xor U26074 (N_26074,N_25290,N_25141);
xor U26075 (N_26075,N_25671,N_25594);
nor U26076 (N_26076,N_25862,N_25489);
xnor U26077 (N_26077,N_25722,N_25869);
and U26078 (N_26078,N_25199,N_25896);
nand U26079 (N_26079,N_25685,N_25174);
nand U26080 (N_26080,N_25146,N_25353);
nor U26081 (N_26081,N_25439,N_25845);
nand U26082 (N_26082,N_25733,N_25098);
nor U26083 (N_26083,N_25271,N_25557);
nor U26084 (N_26084,N_25008,N_25641);
xor U26085 (N_26085,N_25007,N_25046);
or U26086 (N_26086,N_25232,N_25957);
nor U26087 (N_26087,N_25151,N_25465);
nand U26088 (N_26088,N_25509,N_25502);
nand U26089 (N_26089,N_25918,N_25269);
and U26090 (N_26090,N_25019,N_25804);
nand U26091 (N_26091,N_25514,N_25388);
nand U26092 (N_26092,N_25719,N_25361);
nand U26093 (N_26093,N_25989,N_25214);
nand U26094 (N_26094,N_25556,N_25336);
or U26095 (N_26095,N_25322,N_25755);
nand U26096 (N_26096,N_25690,N_25879);
nand U26097 (N_26097,N_25863,N_25453);
nand U26098 (N_26098,N_25285,N_25427);
and U26099 (N_26099,N_25177,N_25704);
or U26100 (N_26100,N_25805,N_25367);
or U26101 (N_26101,N_25318,N_25121);
nand U26102 (N_26102,N_25197,N_25405);
and U26103 (N_26103,N_25619,N_25640);
or U26104 (N_26104,N_25195,N_25142);
nor U26105 (N_26105,N_25482,N_25294);
nor U26106 (N_26106,N_25349,N_25180);
or U26107 (N_26107,N_25407,N_25328);
xor U26108 (N_26108,N_25799,N_25305);
nand U26109 (N_26109,N_25620,N_25803);
nor U26110 (N_26110,N_25635,N_25555);
xor U26111 (N_26111,N_25877,N_25586);
xnor U26112 (N_26112,N_25868,N_25758);
or U26113 (N_26113,N_25380,N_25069);
and U26114 (N_26114,N_25593,N_25658);
nor U26115 (N_26115,N_25872,N_25249);
nand U26116 (N_26116,N_25830,N_25475);
and U26117 (N_26117,N_25060,N_25833);
nand U26118 (N_26118,N_25892,N_25189);
or U26119 (N_26119,N_25639,N_25698);
xor U26120 (N_26120,N_25653,N_25445);
nor U26121 (N_26121,N_25298,N_25392);
nand U26122 (N_26122,N_25288,N_25539);
xor U26123 (N_26123,N_25815,N_25677);
and U26124 (N_26124,N_25369,N_25510);
or U26125 (N_26125,N_25092,N_25423);
and U26126 (N_26126,N_25601,N_25859);
nor U26127 (N_26127,N_25964,N_25742);
xor U26128 (N_26128,N_25788,N_25903);
and U26129 (N_26129,N_25666,N_25731);
nand U26130 (N_26130,N_25154,N_25178);
xor U26131 (N_26131,N_25039,N_25355);
or U26132 (N_26132,N_25716,N_25464);
xor U26133 (N_26133,N_25820,N_25321);
xnor U26134 (N_26134,N_25534,N_25256);
xnor U26135 (N_26135,N_25186,N_25603);
and U26136 (N_26136,N_25540,N_25980);
xor U26137 (N_26137,N_25764,N_25695);
or U26138 (N_26138,N_25968,N_25855);
xnor U26139 (N_26139,N_25338,N_25274);
nand U26140 (N_26140,N_25023,N_25821);
xor U26141 (N_26141,N_25396,N_25739);
nand U26142 (N_26142,N_25309,N_25165);
xnor U26143 (N_26143,N_25444,N_25532);
nand U26144 (N_26144,N_25105,N_25201);
nor U26145 (N_26145,N_25419,N_25250);
nor U26146 (N_26146,N_25068,N_25975);
or U26147 (N_26147,N_25783,N_25576);
and U26148 (N_26148,N_25273,N_25055);
nor U26149 (N_26149,N_25223,N_25266);
and U26150 (N_26150,N_25853,N_25703);
xor U26151 (N_26151,N_25346,N_25938);
nand U26152 (N_26152,N_25589,N_25147);
xor U26153 (N_26153,N_25629,N_25725);
nand U26154 (N_26154,N_25286,N_25743);
xnor U26155 (N_26155,N_25348,N_25161);
nand U26156 (N_26156,N_25047,N_25354);
nand U26157 (N_26157,N_25034,N_25365);
nand U26158 (N_26158,N_25442,N_25441);
nand U26159 (N_26159,N_25867,N_25610);
nand U26160 (N_26160,N_25070,N_25575);
xnor U26161 (N_26161,N_25564,N_25443);
or U26162 (N_26162,N_25627,N_25962);
nor U26163 (N_26163,N_25683,N_25079);
xor U26164 (N_26164,N_25384,N_25950);
and U26165 (N_26165,N_25362,N_25544);
and U26166 (N_26166,N_25686,N_25970);
xnor U26167 (N_26167,N_25915,N_25429);
or U26168 (N_26168,N_25492,N_25066);
and U26169 (N_26169,N_25538,N_25470);
and U26170 (N_26170,N_25319,N_25818);
and U26171 (N_26171,N_25573,N_25866);
nand U26172 (N_26172,N_25158,N_25268);
xnor U26173 (N_26173,N_25308,N_25014);
and U26174 (N_26174,N_25622,N_25661);
nand U26175 (N_26175,N_25073,N_25837);
or U26176 (N_26176,N_25779,N_25410);
and U26177 (N_26177,N_25648,N_25519);
xor U26178 (N_26178,N_25824,N_25654);
nand U26179 (N_26179,N_25130,N_25676);
nand U26180 (N_26180,N_25205,N_25839);
or U26181 (N_26181,N_25780,N_25708);
xnor U26182 (N_26182,N_25485,N_25922);
nand U26183 (N_26183,N_25711,N_25785);
or U26184 (N_26184,N_25996,N_25048);
nand U26185 (N_26185,N_25668,N_25689);
nand U26186 (N_26186,N_25156,N_25965);
or U26187 (N_26187,N_25215,N_25551);
and U26188 (N_26188,N_25826,N_25042);
and U26189 (N_26189,N_25734,N_25452);
xor U26190 (N_26190,N_25457,N_25440);
nor U26191 (N_26191,N_25360,N_25920);
xor U26192 (N_26192,N_25501,N_25961);
and U26193 (N_26193,N_25303,N_25313);
nor U26194 (N_26194,N_25679,N_25935);
or U26195 (N_26195,N_25015,N_25582);
nand U26196 (N_26196,N_25227,N_25075);
nor U26197 (N_26197,N_25037,N_25200);
and U26198 (N_26198,N_25907,N_25772);
nor U26199 (N_26199,N_25478,N_25889);
xor U26200 (N_26200,N_25431,N_25649);
xor U26201 (N_26201,N_25850,N_25590);
nand U26202 (N_26202,N_25041,N_25123);
xnor U26203 (N_26203,N_25254,N_25221);
nor U26204 (N_26204,N_25953,N_25966);
nand U26205 (N_26205,N_25763,N_25408);
nand U26206 (N_26206,N_25311,N_25312);
nand U26207 (N_26207,N_25846,N_25991);
nor U26208 (N_26208,N_25481,N_25325);
nor U26209 (N_26209,N_25097,N_25170);
or U26210 (N_26210,N_25304,N_25542);
or U26211 (N_26211,N_25135,N_25212);
and U26212 (N_26212,N_25310,N_25473);
nand U26213 (N_26213,N_25545,N_25691);
and U26214 (N_26214,N_25062,N_25616);
xor U26215 (N_26215,N_25736,N_25086);
or U26216 (N_26216,N_25029,N_25138);
or U26217 (N_26217,N_25076,N_25351);
nand U26218 (N_26218,N_25751,N_25854);
or U26219 (N_26219,N_25418,N_25633);
xnor U26220 (N_26220,N_25235,N_25552);
and U26221 (N_26221,N_25798,N_25881);
and U26222 (N_26222,N_25270,N_25497);
nand U26223 (N_26223,N_25537,N_25302);
and U26224 (N_26224,N_25761,N_25460);
or U26225 (N_26225,N_25625,N_25694);
and U26226 (N_26226,N_25749,N_25243);
xnor U26227 (N_26227,N_25016,N_25277);
nor U26228 (N_26228,N_25021,N_25080);
nand U26229 (N_26229,N_25754,N_25709);
nand U26230 (N_26230,N_25928,N_25762);
nor U26231 (N_26231,N_25276,N_25508);
nor U26232 (N_26232,N_25035,N_25995);
nand U26233 (N_26233,N_25449,N_25687);
nor U26234 (N_26234,N_25612,N_25265);
or U26235 (N_26235,N_25579,N_25280);
nand U26236 (N_26236,N_25373,N_25784);
and U26237 (N_26237,N_25376,N_25063);
nor U26238 (N_26238,N_25518,N_25983);
or U26239 (N_26239,N_25463,N_25374);
nor U26240 (N_26240,N_25997,N_25224);
or U26241 (N_26241,N_25315,N_25588);
and U26242 (N_26242,N_25776,N_25283);
xor U26243 (N_26243,N_25657,N_25595);
or U26244 (N_26244,N_25852,N_25025);
nand U26245 (N_26245,N_25825,N_25834);
xor U26246 (N_26246,N_25366,N_25413);
nor U26247 (N_26247,N_25958,N_25411);
nand U26248 (N_26248,N_25307,N_25166);
or U26249 (N_26249,N_25674,N_25530);
nand U26250 (N_26250,N_25753,N_25732);
nor U26251 (N_26251,N_25909,N_25737);
nor U26252 (N_26252,N_25746,N_25233);
nor U26253 (N_26253,N_25394,N_25878);
and U26254 (N_26254,N_25368,N_25503);
nand U26255 (N_26255,N_25255,N_25517);
nor U26256 (N_26256,N_25644,N_25583);
or U26257 (N_26257,N_25490,N_25655);
xnor U26258 (N_26258,N_25652,N_25451);
xnor U26259 (N_26259,N_25819,N_25119);
xnor U26260 (N_26260,N_25572,N_25851);
or U26261 (N_26261,N_25088,N_25051);
and U26262 (N_26262,N_25257,N_25750);
nand U26263 (N_26263,N_25880,N_25560);
or U26264 (N_26264,N_25172,N_25115);
or U26265 (N_26265,N_25054,N_25173);
and U26266 (N_26266,N_25009,N_25777);
nor U26267 (N_26267,N_25986,N_25972);
nand U26268 (N_26268,N_25768,N_25162);
xnor U26269 (N_26269,N_25901,N_25637);
and U26270 (N_26270,N_25617,N_25122);
and U26271 (N_26271,N_25888,N_25546);
nand U26272 (N_26272,N_25238,N_25211);
nor U26273 (N_26273,N_25943,N_25320);
and U26274 (N_26274,N_25941,N_25642);
and U26275 (N_26275,N_25383,N_25352);
xnor U26276 (N_26276,N_25259,N_25760);
nand U26277 (N_26277,N_25293,N_25488);
nand U26278 (N_26278,N_25038,N_25192);
or U26279 (N_26279,N_25515,N_25933);
and U26280 (N_26280,N_25117,N_25359);
or U26281 (N_26281,N_25978,N_25397);
or U26282 (N_26282,N_25948,N_25587);
and U26283 (N_26283,N_25306,N_25596);
nand U26284 (N_26284,N_25131,N_25446);
and U26285 (N_26285,N_25900,N_25067);
xor U26286 (N_26286,N_25378,N_25636);
nand U26287 (N_26287,N_25428,N_25331);
and U26288 (N_26288,N_25513,N_25251);
and U26289 (N_26289,N_25977,N_25455);
and U26290 (N_26290,N_25894,N_25100);
xnor U26291 (N_26291,N_25876,N_25099);
xnor U26292 (N_26292,N_25159,N_25108);
xnor U26293 (N_26293,N_25904,N_25973);
xnor U26294 (N_26294,N_25494,N_25971);
and U26295 (N_26295,N_25787,N_25245);
and U26296 (N_26296,N_25364,N_25112);
nand U26297 (N_26297,N_25210,N_25239);
and U26298 (N_26298,N_25344,N_25554);
or U26299 (N_26299,N_25149,N_25795);
xor U26300 (N_26300,N_25713,N_25527);
nand U26301 (N_26301,N_25342,N_25581);
or U26302 (N_26302,N_25279,N_25234);
nand U26303 (N_26303,N_25433,N_25114);
or U26304 (N_26304,N_25730,N_25461);
nand U26305 (N_26305,N_25006,N_25144);
or U26306 (N_26306,N_25912,N_25044);
nand U26307 (N_26307,N_25528,N_25767);
and U26308 (N_26308,N_25794,N_25206);
nand U26309 (N_26309,N_25065,N_25832);
and U26310 (N_26310,N_25955,N_25916);
nand U26311 (N_26311,N_25887,N_25203);
xor U26312 (N_26312,N_25190,N_25153);
nor U26313 (N_26313,N_25715,N_25061);
nor U26314 (N_26314,N_25476,N_25477);
nand U26315 (N_26315,N_25504,N_25873);
or U26316 (N_26316,N_25700,N_25134);
nand U26317 (N_26317,N_25024,N_25624);
nand U26318 (N_26318,N_25536,N_25299);
and U26319 (N_26319,N_25152,N_25241);
nand U26320 (N_26320,N_25393,N_25095);
xnor U26321 (N_26321,N_25505,N_25343);
nor U26322 (N_26322,N_25775,N_25591);
and U26323 (N_26323,N_25643,N_25771);
nand U26324 (N_26324,N_25005,N_25726);
nor U26325 (N_26325,N_25415,N_25979);
or U26326 (N_26326,N_25335,N_25931);
nand U26327 (N_26327,N_25333,N_25729);
or U26328 (N_26328,N_25562,N_25988);
xor U26329 (N_26329,N_25807,N_25264);
nor U26330 (N_26330,N_25326,N_25074);
nand U26331 (N_26331,N_25244,N_25672);
nor U26332 (N_26332,N_25101,N_25797);
or U26333 (N_26333,N_25574,N_25078);
and U26334 (N_26334,N_25437,N_25634);
or U26335 (N_26335,N_25157,N_25842);
nor U26336 (N_26336,N_25128,N_25168);
or U26337 (N_26337,N_25535,N_25847);
or U26338 (N_26338,N_25204,N_25498);
and U26339 (N_26339,N_25874,N_25735);
nor U26340 (N_26340,N_25710,N_25930);
nor U26341 (N_26341,N_25895,N_25090);
nand U26342 (N_26342,N_25053,N_25469);
nand U26343 (N_26343,N_25228,N_25295);
nor U26344 (N_26344,N_25645,N_25432);
or U26345 (N_26345,N_25939,N_25430);
xor U26346 (N_26346,N_25357,N_25647);
nor U26347 (N_26347,N_25416,N_25592);
nor U26348 (N_26348,N_25696,N_25614);
xnor U26349 (N_26349,N_25011,N_25145);
and U26350 (N_26350,N_25838,N_25450);
nand U26351 (N_26351,N_25727,N_25323);
and U26352 (N_26352,N_25985,N_25017);
and U26353 (N_26353,N_25447,N_25942);
xor U26354 (N_26354,N_25841,N_25417);
nand U26355 (N_26355,N_25884,N_25181);
nand U26356 (N_26356,N_25618,N_25929);
and U26357 (N_26357,N_25769,N_25782);
nand U26358 (N_26358,N_25998,N_25836);
or U26359 (N_26359,N_25885,N_25139);
or U26360 (N_26360,N_25106,N_25778);
or U26361 (N_26361,N_25414,N_25604);
xnor U26362 (N_26362,N_25954,N_25113);
nand U26363 (N_26363,N_25184,N_25125);
xor U26364 (N_26364,N_25026,N_25401);
and U26365 (N_26365,N_25040,N_25791);
nand U26366 (N_26366,N_25372,N_25813);
and U26367 (N_26367,N_25531,N_25237);
nor U26368 (N_26368,N_25656,N_25651);
xor U26369 (N_26369,N_25247,N_25701);
nand U26370 (N_26370,N_25013,N_25104);
xor U26371 (N_26371,N_25844,N_25835);
or U26372 (N_26372,N_25402,N_25984);
nor U26373 (N_26373,N_25914,N_25773);
and U26374 (N_26374,N_25558,N_25300);
or U26375 (N_26375,N_25665,N_25548);
nor U26376 (N_26376,N_25330,N_25512);
and U26377 (N_26377,N_25721,N_25022);
and U26378 (N_26378,N_25148,N_25282);
xnor U26379 (N_26379,N_25882,N_25688);
xor U26380 (N_26380,N_25160,N_25218);
nand U26381 (N_26381,N_25403,N_25609);
and U26382 (N_26382,N_25120,N_25185);
or U26383 (N_26383,N_25102,N_25525);
and U26384 (N_26384,N_25003,N_25317);
and U26385 (N_26385,N_25563,N_25176);
nor U26386 (N_26386,N_25466,N_25906);
or U26387 (N_26387,N_25856,N_25770);
nor U26388 (N_26388,N_25004,N_25756);
xnor U26389 (N_26389,N_25606,N_25883);
xor U26390 (N_26390,N_25175,N_25926);
xnor U26391 (N_26391,N_25981,N_25087);
and U26392 (N_26392,N_25150,N_25849);
xor U26393 (N_26393,N_25071,N_25801);
and U26394 (N_26394,N_25164,N_25332);
nor U26395 (N_26395,N_25155,N_25571);
or U26396 (N_26396,N_25027,N_25043);
or U26397 (N_26397,N_25602,N_25702);
nand U26398 (N_26398,N_25638,N_25272);
nor U26399 (N_26399,N_25600,N_25871);
xor U26400 (N_26400,N_25523,N_25387);
nor U26401 (N_26401,N_25435,N_25094);
nor U26402 (N_26402,N_25188,N_25036);
or U26403 (N_26403,N_25608,N_25002);
nor U26404 (N_26404,N_25949,N_25426);
xor U26405 (N_26405,N_25806,N_25663);
or U26406 (N_26406,N_25793,N_25382);
or U26407 (N_26407,N_25816,N_25127);
xnor U26408 (N_26408,N_25111,N_25963);
nand U26409 (N_26409,N_25936,N_25550);
xnor U26410 (N_26410,N_25179,N_25136);
and U26411 (N_26411,N_25828,N_25969);
or U26412 (N_26412,N_25567,N_25093);
xnor U26413 (N_26413,N_25347,N_25720);
nor U26414 (N_26414,N_25605,N_25670);
xor U26415 (N_26415,N_25748,N_25240);
or U26416 (N_26416,N_25050,N_25495);
and U26417 (N_26417,N_25356,N_25621);
nand U26418 (N_26418,N_25516,N_25220);
and U26419 (N_26419,N_25434,N_25171);
nand U26420 (N_26420,N_25529,N_25202);
and U26421 (N_26421,N_25454,N_25072);
or U26422 (N_26422,N_25511,N_25278);
and U26423 (N_26423,N_25091,N_25675);
nand U26424 (N_26424,N_25267,N_25143);
xnor U26425 (N_26425,N_25831,N_25705);
nor U26426 (N_26426,N_25707,N_25615);
or U26427 (N_26427,N_25923,N_25260);
nand U26428 (N_26428,N_25001,N_25110);
nand U26429 (N_26429,N_25840,N_25823);
xnor U26430 (N_26430,N_25789,N_25020);
nor U26431 (N_26431,N_25327,N_25493);
nand U26432 (N_26432,N_25626,N_25052);
or U26433 (N_26433,N_25967,N_25800);
or U26434 (N_26434,N_25472,N_25246);
or U26435 (N_26435,N_25081,N_25946);
or U26436 (N_26436,N_25391,N_25561);
and U26437 (N_26437,N_25345,N_25520);
xor U26438 (N_26438,N_25261,N_25898);
nor U26439 (N_26439,N_25341,N_25085);
or U26440 (N_26440,N_25316,N_25253);
xnor U26441 (N_26441,N_25096,N_25886);
and U26442 (N_26442,N_25580,N_25802);
xnor U26443 (N_26443,N_25717,N_25566);
or U26444 (N_26444,N_25389,N_25012);
nand U26445 (N_26445,N_25578,N_25448);
or U26446 (N_26446,N_25137,N_25714);
or U26447 (N_26447,N_25660,N_25340);
nor U26448 (N_26448,N_25409,N_25524);
and U26449 (N_26449,N_25568,N_25543);
nand U26450 (N_26450,N_25425,N_25377);
and U26451 (N_26451,N_25960,N_25107);
or U26452 (N_26452,N_25597,N_25406);
xnor U26453 (N_26453,N_25412,N_25077);
or U26454 (N_26454,N_25324,N_25891);
xnor U26455 (N_26455,N_25662,N_25650);
nor U26456 (N_26456,N_25757,N_25339);
and U26457 (N_26457,N_25194,N_25129);
xor U26458 (N_26458,N_25169,N_25207);
and U26459 (N_26459,N_25723,N_25934);
and U26460 (N_26460,N_25208,N_25400);
xor U26461 (N_26461,N_25913,N_25506);
nand U26462 (N_26462,N_25987,N_25893);
xnor U26463 (N_26463,N_25724,N_25196);
xnor U26464 (N_26464,N_25829,N_25858);
or U26465 (N_26465,N_25109,N_25993);
nand U26466 (N_26466,N_25291,N_25814);
xor U26467 (N_26467,N_25974,N_25219);
nor U26468 (N_26468,N_25028,N_25865);
nor U26469 (N_26469,N_25458,N_25921);
xor U26470 (N_26470,N_25864,N_25059);
and U26471 (N_26471,N_25499,N_25598);
nor U26472 (N_26472,N_25547,N_25927);
nor U26473 (N_26473,N_25386,N_25712);
nand U26474 (N_26474,N_25140,N_25569);
nor U26475 (N_26475,N_25467,N_25902);
nand U26476 (N_26476,N_25225,N_25474);
xor U26477 (N_26477,N_25812,N_25999);
and U26478 (N_26478,N_25258,N_25229);
nor U26479 (N_26479,N_25103,N_25371);
and U26480 (N_26480,N_25924,N_25133);
nor U26481 (N_26481,N_25242,N_25947);
nand U26482 (N_26482,N_25363,N_25480);
nand U26483 (N_26483,N_25632,N_25468);
nor U26484 (N_26484,N_25486,N_25744);
or U26485 (N_26485,N_25496,N_25056);
or U26486 (N_26486,N_25491,N_25252);
or U26487 (N_26487,N_25919,N_25848);
and U26488 (N_26488,N_25422,N_25932);
xnor U26489 (N_26489,N_25375,N_25030);
xnor U26490 (N_26490,N_25741,N_25718);
and U26491 (N_26491,N_25222,N_25990);
and U26492 (N_26492,N_25385,N_25781);
xnor U26493 (N_26493,N_25337,N_25132);
nand U26494 (N_26494,N_25808,N_25738);
nor U26495 (N_26495,N_25740,N_25585);
and U26496 (N_26496,N_25745,N_25959);
or U26497 (N_26497,N_25951,N_25911);
nand U26498 (N_26498,N_25032,N_25870);
and U26499 (N_26499,N_25522,N_25124);
xnor U26500 (N_26500,N_25108,N_25205);
xnor U26501 (N_26501,N_25309,N_25582);
or U26502 (N_26502,N_25773,N_25338);
nand U26503 (N_26503,N_25616,N_25345);
nor U26504 (N_26504,N_25086,N_25091);
xnor U26505 (N_26505,N_25774,N_25367);
xor U26506 (N_26506,N_25531,N_25924);
xor U26507 (N_26507,N_25737,N_25178);
nor U26508 (N_26508,N_25525,N_25338);
and U26509 (N_26509,N_25592,N_25997);
nand U26510 (N_26510,N_25950,N_25199);
or U26511 (N_26511,N_25864,N_25706);
nor U26512 (N_26512,N_25481,N_25276);
xnor U26513 (N_26513,N_25746,N_25639);
and U26514 (N_26514,N_25043,N_25616);
xnor U26515 (N_26515,N_25481,N_25468);
nand U26516 (N_26516,N_25203,N_25691);
or U26517 (N_26517,N_25235,N_25070);
nand U26518 (N_26518,N_25556,N_25983);
or U26519 (N_26519,N_25418,N_25635);
and U26520 (N_26520,N_25466,N_25822);
or U26521 (N_26521,N_25136,N_25937);
and U26522 (N_26522,N_25531,N_25516);
and U26523 (N_26523,N_25691,N_25749);
and U26524 (N_26524,N_25438,N_25558);
or U26525 (N_26525,N_25792,N_25097);
and U26526 (N_26526,N_25373,N_25121);
nor U26527 (N_26527,N_25379,N_25892);
nand U26528 (N_26528,N_25172,N_25603);
nor U26529 (N_26529,N_25933,N_25380);
xor U26530 (N_26530,N_25205,N_25487);
nor U26531 (N_26531,N_25198,N_25699);
nand U26532 (N_26532,N_25121,N_25092);
xnor U26533 (N_26533,N_25952,N_25483);
nand U26534 (N_26534,N_25264,N_25995);
xnor U26535 (N_26535,N_25956,N_25190);
or U26536 (N_26536,N_25655,N_25374);
and U26537 (N_26537,N_25912,N_25808);
nand U26538 (N_26538,N_25365,N_25585);
xor U26539 (N_26539,N_25108,N_25565);
and U26540 (N_26540,N_25017,N_25812);
nand U26541 (N_26541,N_25466,N_25350);
or U26542 (N_26542,N_25189,N_25290);
or U26543 (N_26543,N_25845,N_25020);
xnor U26544 (N_26544,N_25485,N_25441);
nor U26545 (N_26545,N_25535,N_25848);
or U26546 (N_26546,N_25251,N_25008);
xor U26547 (N_26547,N_25925,N_25697);
or U26548 (N_26548,N_25953,N_25629);
nor U26549 (N_26549,N_25058,N_25507);
nand U26550 (N_26550,N_25898,N_25987);
nand U26551 (N_26551,N_25047,N_25211);
xor U26552 (N_26552,N_25770,N_25231);
and U26553 (N_26553,N_25788,N_25728);
xor U26554 (N_26554,N_25433,N_25813);
nor U26555 (N_26555,N_25065,N_25442);
xnor U26556 (N_26556,N_25141,N_25945);
xor U26557 (N_26557,N_25824,N_25738);
xor U26558 (N_26558,N_25340,N_25405);
nand U26559 (N_26559,N_25669,N_25102);
nor U26560 (N_26560,N_25462,N_25086);
or U26561 (N_26561,N_25759,N_25017);
xnor U26562 (N_26562,N_25989,N_25418);
nand U26563 (N_26563,N_25763,N_25359);
nand U26564 (N_26564,N_25122,N_25007);
or U26565 (N_26565,N_25282,N_25550);
and U26566 (N_26566,N_25155,N_25201);
nor U26567 (N_26567,N_25480,N_25725);
or U26568 (N_26568,N_25607,N_25649);
nor U26569 (N_26569,N_25034,N_25330);
or U26570 (N_26570,N_25008,N_25720);
and U26571 (N_26571,N_25035,N_25276);
or U26572 (N_26572,N_25720,N_25299);
xnor U26573 (N_26573,N_25420,N_25316);
and U26574 (N_26574,N_25852,N_25530);
nor U26575 (N_26575,N_25499,N_25934);
and U26576 (N_26576,N_25264,N_25876);
and U26577 (N_26577,N_25837,N_25962);
or U26578 (N_26578,N_25811,N_25316);
and U26579 (N_26579,N_25763,N_25735);
nand U26580 (N_26580,N_25814,N_25213);
and U26581 (N_26581,N_25179,N_25605);
xor U26582 (N_26582,N_25495,N_25768);
and U26583 (N_26583,N_25504,N_25092);
and U26584 (N_26584,N_25045,N_25546);
or U26585 (N_26585,N_25906,N_25313);
nand U26586 (N_26586,N_25862,N_25632);
nand U26587 (N_26587,N_25091,N_25915);
xor U26588 (N_26588,N_25353,N_25707);
xnor U26589 (N_26589,N_25804,N_25623);
xnor U26590 (N_26590,N_25013,N_25048);
or U26591 (N_26591,N_25278,N_25251);
nand U26592 (N_26592,N_25416,N_25343);
and U26593 (N_26593,N_25615,N_25328);
or U26594 (N_26594,N_25356,N_25216);
nand U26595 (N_26595,N_25808,N_25242);
nor U26596 (N_26596,N_25689,N_25313);
and U26597 (N_26597,N_25157,N_25928);
and U26598 (N_26598,N_25307,N_25897);
or U26599 (N_26599,N_25461,N_25071);
or U26600 (N_26600,N_25075,N_25471);
nor U26601 (N_26601,N_25015,N_25604);
xnor U26602 (N_26602,N_25017,N_25442);
xor U26603 (N_26603,N_25358,N_25566);
xor U26604 (N_26604,N_25407,N_25269);
xor U26605 (N_26605,N_25946,N_25321);
nor U26606 (N_26606,N_25348,N_25551);
nor U26607 (N_26607,N_25169,N_25960);
or U26608 (N_26608,N_25633,N_25085);
nor U26609 (N_26609,N_25011,N_25549);
nand U26610 (N_26610,N_25319,N_25789);
and U26611 (N_26611,N_25625,N_25987);
nor U26612 (N_26612,N_25467,N_25898);
nand U26613 (N_26613,N_25891,N_25018);
nor U26614 (N_26614,N_25701,N_25616);
xor U26615 (N_26615,N_25379,N_25795);
nand U26616 (N_26616,N_25344,N_25280);
and U26617 (N_26617,N_25462,N_25857);
or U26618 (N_26618,N_25306,N_25741);
nand U26619 (N_26619,N_25685,N_25810);
xor U26620 (N_26620,N_25143,N_25649);
nand U26621 (N_26621,N_25120,N_25440);
nand U26622 (N_26622,N_25697,N_25981);
nor U26623 (N_26623,N_25967,N_25602);
or U26624 (N_26624,N_25112,N_25866);
or U26625 (N_26625,N_25183,N_25927);
or U26626 (N_26626,N_25420,N_25583);
nor U26627 (N_26627,N_25938,N_25480);
nand U26628 (N_26628,N_25553,N_25666);
or U26629 (N_26629,N_25754,N_25962);
and U26630 (N_26630,N_25041,N_25796);
xor U26631 (N_26631,N_25727,N_25866);
or U26632 (N_26632,N_25307,N_25450);
nand U26633 (N_26633,N_25145,N_25236);
nor U26634 (N_26634,N_25401,N_25435);
xor U26635 (N_26635,N_25851,N_25943);
nor U26636 (N_26636,N_25268,N_25733);
or U26637 (N_26637,N_25245,N_25340);
xor U26638 (N_26638,N_25234,N_25340);
xnor U26639 (N_26639,N_25782,N_25125);
nor U26640 (N_26640,N_25599,N_25203);
xnor U26641 (N_26641,N_25392,N_25249);
nor U26642 (N_26642,N_25280,N_25399);
and U26643 (N_26643,N_25265,N_25530);
and U26644 (N_26644,N_25730,N_25989);
nand U26645 (N_26645,N_25491,N_25284);
or U26646 (N_26646,N_25424,N_25385);
or U26647 (N_26647,N_25478,N_25825);
or U26648 (N_26648,N_25453,N_25866);
nor U26649 (N_26649,N_25624,N_25622);
and U26650 (N_26650,N_25004,N_25053);
or U26651 (N_26651,N_25609,N_25751);
xnor U26652 (N_26652,N_25288,N_25351);
or U26653 (N_26653,N_25780,N_25932);
xor U26654 (N_26654,N_25803,N_25448);
nand U26655 (N_26655,N_25142,N_25356);
nor U26656 (N_26656,N_25932,N_25743);
xor U26657 (N_26657,N_25324,N_25322);
or U26658 (N_26658,N_25600,N_25361);
xnor U26659 (N_26659,N_25974,N_25680);
or U26660 (N_26660,N_25200,N_25045);
or U26661 (N_26661,N_25941,N_25872);
xnor U26662 (N_26662,N_25256,N_25658);
nand U26663 (N_26663,N_25923,N_25659);
or U26664 (N_26664,N_25265,N_25165);
xnor U26665 (N_26665,N_25573,N_25672);
and U26666 (N_26666,N_25646,N_25503);
xnor U26667 (N_26667,N_25567,N_25517);
nand U26668 (N_26668,N_25811,N_25491);
nor U26669 (N_26669,N_25431,N_25742);
or U26670 (N_26670,N_25538,N_25634);
xnor U26671 (N_26671,N_25319,N_25843);
or U26672 (N_26672,N_25204,N_25021);
xnor U26673 (N_26673,N_25517,N_25983);
nor U26674 (N_26674,N_25779,N_25307);
and U26675 (N_26675,N_25184,N_25027);
and U26676 (N_26676,N_25691,N_25181);
xnor U26677 (N_26677,N_25670,N_25894);
xnor U26678 (N_26678,N_25211,N_25184);
xor U26679 (N_26679,N_25519,N_25439);
or U26680 (N_26680,N_25775,N_25643);
nor U26681 (N_26681,N_25966,N_25503);
nor U26682 (N_26682,N_25656,N_25839);
xor U26683 (N_26683,N_25669,N_25095);
xnor U26684 (N_26684,N_25566,N_25965);
xor U26685 (N_26685,N_25275,N_25794);
xnor U26686 (N_26686,N_25871,N_25060);
nand U26687 (N_26687,N_25980,N_25314);
or U26688 (N_26688,N_25418,N_25123);
or U26689 (N_26689,N_25483,N_25233);
and U26690 (N_26690,N_25132,N_25937);
xor U26691 (N_26691,N_25732,N_25842);
nand U26692 (N_26692,N_25884,N_25798);
nand U26693 (N_26693,N_25586,N_25064);
and U26694 (N_26694,N_25673,N_25252);
and U26695 (N_26695,N_25975,N_25313);
or U26696 (N_26696,N_25582,N_25048);
xnor U26697 (N_26697,N_25341,N_25785);
nand U26698 (N_26698,N_25273,N_25391);
and U26699 (N_26699,N_25505,N_25657);
xnor U26700 (N_26700,N_25984,N_25252);
nor U26701 (N_26701,N_25954,N_25502);
and U26702 (N_26702,N_25193,N_25566);
and U26703 (N_26703,N_25348,N_25256);
nand U26704 (N_26704,N_25555,N_25736);
or U26705 (N_26705,N_25233,N_25080);
nand U26706 (N_26706,N_25949,N_25546);
nor U26707 (N_26707,N_25520,N_25689);
nor U26708 (N_26708,N_25033,N_25364);
xor U26709 (N_26709,N_25900,N_25673);
nand U26710 (N_26710,N_25756,N_25342);
nand U26711 (N_26711,N_25714,N_25332);
nor U26712 (N_26712,N_25524,N_25478);
nor U26713 (N_26713,N_25171,N_25608);
nor U26714 (N_26714,N_25543,N_25910);
or U26715 (N_26715,N_25802,N_25096);
or U26716 (N_26716,N_25210,N_25464);
nor U26717 (N_26717,N_25116,N_25279);
or U26718 (N_26718,N_25017,N_25600);
nand U26719 (N_26719,N_25088,N_25816);
or U26720 (N_26720,N_25414,N_25519);
nor U26721 (N_26721,N_25487,N_25175);
nand U26722 (N_26722,N_25071,N_25636);
nand U26723 (N_26723,N_25614,N_25805);
nor U26724 (N_26724,N_25272,N_25936);
nand U26725 (N_26725,N_25237,N_25477);
nor U26726 (N_26726,N_25984,N_25327);
and U26727 (N_26727,N_25554,N_25539);
and U26728 (N_26728,N_25705,N_25740);
and U26729 (N_26729,N_25250,N_25457);
xnor U26730 (N_26730,N_25748,N_25214);
nand U26731 (N_26731,N_25170,N_25190);
nand U26732 (N_26732,N_25107,N_25942);
and U26733 (N_26733,N_25592,N_25835);
and U26734 (N_26734,N_25380,N_25301);
or U26735 (N_26735,N_25326,N_25574);
nor U26736 (N_26736,N_25047,N_25605);
nand U26737 (N_26737,N_25339,N_25737);
nor U26738 (N_26738,N_25210,N_25875);
nand U26739 (N_26739,N_25115,N_25801);
nand U26740 (N_26740,N_25477,N_25422);
nor U26741 (N_26741,N_25545,N_25634);
nand U26742 (N_26742,N_25584,N_25954);
and U26743 (N_26743,N_25647,N_25557);
xnor U26744 (N_26744,N_25864,N_25876);
or U26745 (N_26745,N_25865,N_25701);
nor U26746 (N_26746,N_25193,N_25408);
or U26747 (N_26747,N_25237,N_25017);
nand U26748 (N_26748,N_25128,N_25702);
nand U26749 (N_26749,N_25295,N_25779);
or U26750 (N_26750,N_25488,N_25671);
nor U26751 (N_26751,N_25034,N_25842);
xor U26752 (N_26752,N_25001,N_25342);
nand U26753 (N_26753,N_25466,N_25361);
and U26754 (N_26754,N_25677,N_25958);
and U26755 (N_26755,N_25094,N_25905);
xnor U26756 (N_26756,N_25437,N_25610);
and U26757 (N_26757,N_25641,N_25629);
or U26758 (N_26758,N_25693,N_25444);
xor U26759 (N_26759,N_25955,N_25872);
and U26760 (N_26760,N_25821,N_25618);
nand U26761 (N_26761,N_25455,N_25562);
nand U26762 (N_26762,N_25997,N_25857);
nand U26763 (N_26763,N_25855,N_25691);
nor U26764 (N_26764,N_25389,N_25040);
nand U26765 (N_26765,N_25267,N_25989);
and U26766 (N_26766,N_25474,N_25092);
and U26767 (N_26767,N_25347,N_25112);
or U26768 (N_26768,N_25688,N_25167);
nor U26769 (N_26769,N_25902,N_25291);
nand U26770 (N_26770,N_25751,N_25397);
and U26771 (N_26771,N_25160,N_25308);
nor U26772 (N_26772,N_25582,N_25612);
xor U26773 (N_26773,N_25251,N_25320);
nor U26774 (N_26774,N_25519,N_25814);
or U26775 (N_26775,N_25347,N_25527);
xnor U26776 (N_26776,N_25117,N_25734);
nor U26777 (N_26777,N_25992,N_25285);
xor U26778 (N_26778,N_25644,N_25754);
xor U26779 (N_26779,N_25399,N_25613);
nor U26780 (N_26780,N_25878,N_25679);
or U26781 (N_26781,N_25670,N_25484);
or U26782 (N_26782,N_25523,N_25456);
nand U26783 (N_26783,N_25873,N_25091);
nor U26784 (N_26784,N_25059,N_25751);
nand U26785 (N_26785,N_25903,N_25387);
nor U26786 (N_26786,N_25789,N_25599);
nand U26787 (N_26787,N_25444,N_25309);
and U26788 (N_26788,N_25185,N_25769);
nand U26789 (N_26789,N_25296,N_25630);
nor U26790 (N_26790,N_25085,N_25588);
nand U26791 (N_26791,N_25198,N_25519);
nand U26792 (N_26792,N_25910,N_25787);
xnor U26793 (N_26793,N_25999,N_25218);
nand U26794 (N_26794,N_25007,N_25601);
and U26795 (N_26795,N_25656,N_25544);
or U26796 (N_26796,N_25831,N_25924);
nor U26797 (N_26797,N_25082,N_25198);
nand U26798 (N_26798,N_25367,N_25141);
xnor U26799 (N_26799,N_25990,N_25885);
nor U26800 (N_26800,N_25963,N_25953);
xor U26801 (N_26801,N_25298,N_25879);
and U26802 (N_26802,N_25070,N_25326);
xnor U26803 (N_26803,N_25321,N_25934);
and U26804 (N_26804,N_25167,N_25597);
nand U26805 (N_26805,N_25766,N_25605);
nand U26806 (N_26806,N_25676,N_25175);
nand U26807 (N_26807,N_25763,N_25478);
xnor U26808 (N_26808,N_25475,N_25698);
nand U26809 (N_26809,N_25603,N_25979);
nand U26810 (N_26810,N_25911,N_25389);
and U26811 (N_26811,N_25844,N_25968);
and U26812 (N_26812,N_25397,N_25261);
and U26813 (N_26813,N_25404,N_25170);
or U26814 (N_26814,N_25134,N_25849);
or U26815 (N_26815,N_25340,N_25495);
and U26816 (N_26816,N_25395,N_25123);
nor U26817 (N_26817,N_25187,N_25573);
nor U26818 (N_26818,N_25558,N_25410);
nand U26819 (N_26819,N_25209,N_25609);
xnor U26820 (N_26820,N_25083,N_25290);
xnor U26821 (N_26821,N_25934,N_25822);
or U26822 (N_26822,N_25855,N_25354);
xnor U26823 (N_26823,N_25086,N_25082);
nor U26824 (N_26824,N_25209,N_25890);
nand U26825 (N_26825,N_25048,N_25152);
and U26826 (N_26826,N_25473,N_25487);
or U26827 (N_26827,N_25099,N_25638);
nor U26828 (N_26828,N_25867,N_25417);
xnor U26829 (N_26829,N_25235,N_25561);
nor U26830 (N_26830,N_25934,N_25842);
nand U26831 (N_26831,N_25123,N_25523);
nor U26832 (N_26832,N_25352,N_25269);
and U26833 (N_26833,N_25618,N_25545);
and U26834 (N_26834,N_25997,N_25435);
or U26835 (N_26835,N_25244,N_25163);
or U26836 (N_26836,N_25778,N_25266);
and U26837 (N_26837,N_25013,N_25747);
xnor U26838 (N_26838,N_25939,N_25257);
nor U26839 (N_26839,N_25470,N_25889);
nor U26840 (N_26840,N_25189,N_25433);
nor U26841 (N_26841,N_25693,N_25200);
nand U26842 (N_26842,N_25356,N_25130);
nand U26843 (N_26843,N_25523,N_25360);
nand U26844 (N_26844,N_25072,N_25308);
nand U26845 (N_26845,N_25528,N_25812);
or U26846 (N_26846,N_25263,N_25536);
and U26847 (N_26847,N_25226,N_25510);
nor U26848 (N_26848,N_25536,N_25191);
and U26849 (N_26849,N_25387,N_25676);
nor U26850 (N_26850,N_25064,N_25471);
xnor U26851 (N_26851,N_25578,N_25545);
nand U26852 (N_26852,N_25297,N_25298);
and U26853 (N_26853,N_25357,N_25592);
and U26854 (N_26854,N_25649,N_25159);
or U26855 (N_26855,N_25692,N_25089);
nor U26856 (N_26856,N_25090,N_25017);
and U26857 (N_26857,N_25357,N_25917);
or U26858 (N_26858,N_25519,N_25501);
nand U26859 (N_26859,N_25446,N_25051);
xor U26860 (N_26860,N_25823,N_25717);
xor U26861 (N_26861,N_25393,N_25926);
xnor U26862 (N_26862,N_25507,N_25920);
nor U26863 (N_26863,N_25760,N_25162);
nor U26864 (N_26864,N_25614,N_25933);
nor U26865 (N_26865,N_25582,N_25104);
or U26866 (N_26866,N_25554,N_25931);
or U26867 (N_26867,N_25476,N_25155);
nor U26868 (N_26868,N_25898,N_25365);
nor U26869 (N_26869,N_25212,N_25649);
xnor U26870 (N_26870,N_25839,N_25054);
nor U26871 (N_26871,N_25901,N_25728);
nand U26872 (N_26872,N_25301,N_25579);
nor U26873 (N_26873,N_25126,N_25100);
xnor U26874 (N_26874,N_25084,N_25473);
nand U26875 (N_26875,N_25943,N_25986);
nand U26876 (N_26876,N_25606,N_25422);
or U26877 (N_26877,N_25395,N_25746);
and U26878 (N_26878,N_25017,N_25431);
or U26879 (N_26879,N_25259,N_25041);
and U26880 (N_26880,N_25595,N_25326);
and U26881 (N_26881,N_25190,N_25163);
nor U26882 (N_26882,N_25635,N_25517);
nor U26883 (N_26883,N_25147,N_25734);
nand U26884 (N_26884,N_25051,N_25079);
and U26885 (N_26885,N_25863,N_25019);
or U26886 (N_26886,N_25801,N_25484);
nor U26887 (N_26887,N_25694,N_25381);
xor U26888 (N_26888,N_25406,N_25416);
xor U26889 (N_26889,N_25703,N_25110);
or U26890 (N_26890,N_25514,N_25373);
and U26891 (N_26891,N_25686,N_25028);
nand U26892 (N_26892,N_25051,N_25582);
xnor U26893 (N_26893,N_25176,N_25721);
nand U26894 (N_26894,N_25056,N_25862);
or U26895 (N_26895,N_25977,N_25110);
nor U26896 (N_26896,N_25623,N_25238);
nor U26897 (N_26897,N_25512,N_25351);
and U26898 (N_26898,N_25731,N_25418);
nor U26899 (N_26899,N_25666,N_25794);
or U26900 (N_26900,N_25252,N_25828);
or U26901 (N_26901,N_25187,N_25362);
or U26902 (N_26902,N_25545,N_25270);
nor U26903 (N_26903,N_25031,N_25849);
and U26904 (N_26904,N_25190,N_25910);
and U26905 (N_26905,N_25546,N_25432);
nand U26906 (N_26906,N_25006,N_25745);
xor U26907 (N_26907,N_25589,N_25242);
xor U26908 (N_26908,N_25088,N_25849);
or U26909 (N_26909,N_25484,N_25278);
nand U26910 (N_26910,N_25934,N_25719);
nand U26911 (N_26911,N_25801,N_25998);
and U26912 (N_26912,N_25813,N_25034);
nand U26913 (N_26913,N_25540,N_25113);
nor U26914 (N_26914,N_25296,N_25568);
xor U26915 (N_26915,N_25602,N_25147);
and U26916 (N_26916,N_25585,N_25648);
nor U26917 (N_26917,N_25546,N_25683);
nor U26918 (N_26918,N_25903,N_25345);
nor U26919 (N_26919,N_25160,N_25681);
xnor U26920 (N_26920,N_25739,N_25387);
and U26921 (N_26921,N_25322,N_25230);
and U26922 (N_26922,N_25014,N_25675);
nand U26923 (N_26923,N_25584,N_25151);
and U26924 (N_26924,N_25994,N_25849);
nand U26925 (N_26925,N_25489,N_25948);
nand U26926 (N_26926,N_25509,N_25607);
xor U26927 (N_26927,N_25009,N_25668);
or U26928 (N_26928,N_25245,N_25896);
and U26929 (N_26929,N_25060,N_25861);
xnor U26930 (N_26930,N_25196,N_25121);
nand U26931 (N_26931,N_25662,N_25897);
or U26932 (N_26932,N_25961,N_25379);
nand U26933 (N_26933,N_25085,N_25981);
nand U26934 (N_26934,N_25724,N_25232);
nor U26935 (N_26935,N_25201,N_25361);
xor U26936 (N_26936,N_25348,N_25132);
and U26937 (N_26937,N_25930,N_25392);
nor U26938 (N_26938,N_25491,N_25323);
and U26939 (N_26939,N_25752,N_25337);
nand U26940 (N_26940,N_25395,N_25896);
nand U26941 (N_26941,N_25527,N_25122);
xnor U26942 (N_26942,N_25862,N_25491);
or U26943 (N_26943,N_25666,N_25188);
nand U26944 (N_26944,N_25903,N_25811);
nand U26945 (N_26945,N_25932,N_25545);
and U26946 (N_26946,N_25110,N_25800);
xnor U26947 (N_26947,N_25529,N_25047);
xor U26948 (N_26948,N_25541,N_25097);
nand U26949 (N_26949,N_25803,N_25876);
and U26950 (N_26950,N_25449,N_25130);
and U26951 (N_26951,N_25637,N_25974);
nand U26952 (N_26952,N_25728,N_25386);
nand U26953 (N_26953,N_25311,N_25381);
xnor U26954 (N_26954,N_25874,N_25994);
xnor U26955 (N_26955,N_25994,N_25190);
nor U26956 (N_26956,N_25981,N_25917);
nor U26957 (N_26957,N_25263,N_25175);
nor U26958 (N_26958,N_25176,N_25667);
xor U26959 (N_26959,N_25323,N_25459);
xnor U26960 (N_26960,N_25645,N_25104);
and U26961 (N_26961,N_25118,N_25878);
nand U26962 (N_26962,N_25951,N_25422);
xnor U26963 (N_26963,N_25185,N_25861);
nor U26964 (N_26964,N_25216,N_25024);
xor U26965 (N_26965,N_25386,N_25517);
xnor U26966 (N_26966,N_25538,N_25316);
or U26967 (N_26967,N_25063,N_25311);
nand U26968 (N_26968,N_25573,N_25836);
or U26969 (N_26969,N_25729,N_25616);
nand U26970 (N_26970,N_25033,N_25163);
and U26971 (N_26971,N_25352,N_25595);
or U26972 (N_26972,N_25927,N_25586);
or U26973 (N_26973,N_25110,N_25903);
xor U26974 (N_26974,N_25863,N_25941);
and U26975 (N_26975,N_25186,N_25670);
and U26976 (N_26976,N_25458,N_25274);
or U26977 (N_26977,N_25954,N_25982);
or U26978 (N_26978,N_25561,N_25281);
xor U26979 (N_26979,N_25480,N_25373);
and U26980 (N_26980,N_25465,N_25357);
or U26981 (N_26981,N_25150,N_25310);
xnor U26982 (N_26982,N_25647,N_25289);
or U26983 (N_26983,N_25951,N_25274);
and U26984 (N_26984,N_25917,N_25402);
nand U26985 (N_26985,N_25489,N_25193);
nor U26986 (N_26986,N_25339,N_25271);
and U26987 (N_26987,N_25794,N_25940);
nor U26988 (N_26988,N_25748,N_25180);
or U26989 (N_26989,N_25933,N_25286);
and U26990 (N_26990,N_25109,N_25659);
or U26991 (N_26991,N_25615,N_25219);
and U26992 (N_26992,N_25740,N_25842);
xor U26993 (N_26993,N_25528,N_25702);
and U26994 (N_26994,N_25571,N_25880);
nor U26995 (N_26995,N_25934,N_25506);
and U26996 (N_26996,N_25439,N_25266);
nor U26997 (N_26997,N_25185,N_25521);
nand U26998 (N_26998,N_25640,N_25681);
or U26999 (N_26999,N_25913,N_25772);
or U27000 (N_27000,N_26045,N_26462);
or U27001 (N_27001,N_26257,N_26439);
or U27002 (N_27002,N_26375,N_26816);
xnor U27003 (N_27003,N_26326,N_26145);
and U27004 (N_27004,N_26229,N_26446);
and U27005 (N_27005,N_26417,N_26719);
nand U27006 (N_27006,N_26562,N_26563);
nor U27007 (N_27007,N_26499,N_26502);
nor U27008 (N_27008,N_26634,N_26508);
xor U27009 (N_27009,N_26636,N_26961);
nor U27010 (N_27010,N_26349,N_26359);
nand U27011 (N_27011,N_26791,N_26975);
or U27012 (N_27012,N_26560,N_26172);
nor U27013 (N_27013,N_26146,N_26454);
nor U27014 (N_27014,N_26773,N_26472);
and U27015 (N_27015,N_26666,N_26277);
and U27016 (N_27016,N_26201,N_26280);
nand U27017 (N_27017,N_26995,N_26405);
xnor U27018 (N_27018,N_26874,N_26970);
and U27019 (N_27019,N_26735,N_26497);
and U27020 (N_27020,N_26677,N_26569);
nor U27021 (N_27021,N_26253,N_26701);
or U27022 (N_27022,N_26565,N_26682);
nor U27023 (N_27023,N_26904,N_26096);
or U27024 (N_27024,N_26684,N_26415);
or U27025 (N_27025,N_26534,N_26265);
xor U27026 (N_27026,N_26383,N_26004);
or U27027 (N_27027,N_26269,N_26545);
and U27028 (N_27028,N_26721,N_26709);
nand U27029 (N_27029,N_26268,N_26079);
and U27030 (N_27030,N_26912,N_26817);
xor U27031 (N_27031,N_26109,N_26780);
nand U27032 (N_27032,N_26604,N_26959);
and U27033 (N_27033,N_26142,N_26498);
xnor U27034 (N_27034,N_26882,N_26585);
or U27035 (N_27035,N_26270,N_26188);
or U27036 (N_27036,N_26619,N_26749);
or U27037 (N_27037,N_26181,N_26612);
xor U27038 (N_27038,N_26302,N_26789);
nor U27039 (N_27039,N_26605,N_26595);
or U27040 (N_27040,N_26191,N_26160);
nand U27041 (N_27041,N_26189,N_26070);
xor U27042 (N_27042,N_26111,N_26695);
nand U27043 (N_27043,N_26430,N_26121);
and U27044 (N_27044,N_26019,N_26960);
nor U27045 (N_27045,N_26292,N_26517);
xor U27046 (N_27046,N_26140,N_26209);
and U27047 (N_27047,N_26575,N_26566);
xor U27048 (N_27048,N_26944,N_26414);
xnor U27049 (N_27049,N_26710,N_26673);
nor U27050 (N_27050,N_26224,N_26821);
and U27051 (N_27051,N_26119,N_26078);
nand U27052 (N_27052,N_26842,N_26781);
nand U27053 (N_27053,N_26514,N_26969);
nor U27054 (N_27054,N_26819,N_26449);
and U27055 (N_27055,N_26543,N_26425);
xor U27056 (N_27056,N_26128,N_26927);
nor U27057 (N_27057,N_26579,N_26473);
and U27058 (N_27058,N_26977,N_26031);
nand U27059 (N_27059,N_26014,N_26306);
and U27060 (N_27060,N_26437,N_26830);
and U27061 (N_27061,N_26086,N_26590);
and U27062 (N_27062,N_26054,N_26312);
and U27063 (N_27063,N_26914,N_26748);
nand U27064 (N_27064,N_26124,N_26782);
xor U27065 (N_27065,N_26422,N_26840);
and U27066 (N_27066,N_26831,N_26993);
and U27067 (N_27067,N_26456,N_26942);
or U27068 (N_27068,N_26835,N_26335);
xnor U27069 (N_27069,N_26548,N_26101);
xnor U27070 (N_27070,N_26934,N_26374);
nand U27071 (N_27071,N_26857,N_26899);
nor U27072 (N_27072,N_26123,N_26032);
xor U27073 (N_27073,N_26327,N_26216);
or U27074 (N_27074,N_26600,N_26175);
nor U27075 (N_27075,N_26855,N_26587);
and U27076 (N_27076,N_26367,N_26561);
xor U27077 (N_27077,N_26853,N_26578);
and U27078 (N_27078,N_26668,N_26826);
nor U27079 (N_27079,N_26594,N_26930);
and U27080 (N_27080,N_26152,N_26949);
and U27081 (N_27081,N_26137,N_26156);
or U27082 (N_27082,N_26161,N_26809);
or U27083 (N_27083,N_26402,N_26676);
nor U27084 (N_27084,N_26282,N_26073);
or U27085 (N_27085,N_26737,N_26495);
nor U27086 (N_27086,N_26386,N_26599);
and U27087 (N_27087,N_26505,N_26445);
nand U27088 (N_27088,N_26886,N_26767);
xnor U27089 (N_27089,N_26255,N_26916);
nor U27090 (N_27090,N_26616,N_26915);
or U27091 (N_27091,N_26174,N_26378);
nor U27092 (N_27092,N_26082,N_26479);
and U27093 (N_27093,N_26071,N_26918);
and U27094 (N_27094,N_26114,N_26510);
or U27095 (N_27095,N_26968,N_26401);
xnor U27096 (N_27096,N_26868,N_26810);
and U27097 (N_27097,N_26557,N_26556);
and U27098 (N_27098,N_26528,N_26048);
nor U27099 (N_27099,N_26435,N_26500);
or U27100 (N_27100,N_26696,N_26751);
nand U27101 (N_27101,N_26615,N_26726);
nand U27102 (N_27102,N_26559,N_26159);
nor U27103 (N_27103,N_26226,N_26803);
or U27104 (N_27104,N_26281,N_26586);
nand U27105 (N_27105,N_26740,N_26741);
nand U27106 (N_27106,N_26978,N_26602);
and U27107 (N_27107,N_26406,N_26653);
nand U27108 (N_27108,N_26471,N_26897);
and U27109 (N_27109,N_26639,N_26481);
xor U27110 (N_27110,N_26347,N_26834);
and U27111 (N_27111,N_26240,N_26824);
and U27112 (N_27112,N_26245,N_26275);
nand U27113 (N_27113,N_26911,N_26228);
xnor U27114 (N_27114,N_26584,N_26311);
nand U27115 (N_27115,N_26660,N_26232);
or U27116 (N_27116,N_26689,N_26363);
xnor U27117 (N_27117,N_26458,N_26766);
nand U27118 (N_27118,N_26443,N_26203);
or U27119 (N_27119,N_26488,N_26962);
xor U27120 (N_27120,N_26610,N_26008);
and U27121 (N_27121,N_26067,N_26618);
nor U27122 (N_27122,N_26890,N_26597);
and U27123 (N_27123,N_26625,N_26219);
xor U27124 (N_27124,N_26340,N_26080);
xor U27125 (N_27125,N_26711,N_26720);
or U27126 (N_27126,N_26672,N_26820);
nor U27127 (N_27127,N_26316,N_26016);
nor U27128 (N_27128,N_26410,N_26272);
or U27129 (N_27129,N_26674,N_26376);
nor U27130 (N_27130,N_26023,N_26509);
nand U27131 (N_27131,N_26923,N_26681);
nand U27132 (N_27132,N_26800,N_26461);
and U27133 (N_27133,N_26036,N_26870);
nor U27134 (N_27134,N_26427,N_26309);
xor U27135 (N_27135,N_26167,N_26515);
or U27136 (N_27136,N_26837,N_26012);
or U27137 (N_27137,N_26558,N_26343);
nor U27138 (N_27138,N_26654,N_26254);
nor U27139 (N_27139,N_26250,N_26704);
xor U27140 (N_27140,N_26732,N_26865);
xor U27141 (N_27141,N_26757,N_26394);
nand U27142 (N_27142,N_26039,N_26733);
and U27143 (N_27143,N_26208,N_26413);
and U27144 (N_27144,N_26771,N_26999);
or U27145 (N_27145,N_26516,N_26945);
or U27146 (N_27146,N_26804,N_26907);
nand U27147 (N_27147,N_26843,N_26005);
or U27148 (N_27148,N_26205,N_26656);
nor U27149 (N_27149,N_26527,N_26183);
xnor U27150 (N_27150,N_26341,N_26832);
nand U27151 (N_27151,N_26379,N_26165);
nor U27152 (N_27152,N_26358,N_26954);
or U27153 (N_27153,N_26365,N_26103);
xor U27154 (N_27154,N_26357,N_26623);
nand U27155 (N_27155,N_26348,N_26200);
nand U27156 (N_27156,N_26997,N_26238);
nor U27157 (N_27157,N_26779,N_26922);
or U27158 (N_27158,N_26469,N_26428);
and U27159 (N_27159,N_26755,N_26396);
nor U27160 (N_27160,N_26025,N_26910);
or U27161 (N_27161,N_26763,N_26806);
and U27162 (N_27162,N_26212,N_26686);
and U27163 (N_27163,N_26220,N_26705);
and U27164 (N_27164,N_26210,N_26889);
nand U27165 (N_27165,N_26490,N_26313);
and U27166 (N_27166,N_26017,N_26679);
nor U27167 (N_27167,N_26187,N_26083);
xnor U27168 (N_27168,N_26027,N_26215);
nor U27169 (N_27169,N_26862,N_26539);
nor U27170 (N_27170,N_26092,N_26029);
and U27171 (N_27171,N_26589,N_26131);
or U27172 (N_27172,N_26972,N_26278);
or U27173 (N_27173,N_26568,N_26787);
nor U27174 (N_27174,N_26049,N_26033);
xor U27175 (N_27175,N_26052,N_26451);
and U27176 (N_27176,N_26518,N_26043);
nand U27177 (N_27177,N_26521,N_26796);
nand U27178 (N_27178,N_26056,N_26106);
nor U27179 (N_27179,N_26544,N_26845);
nor U27180 (N_27180,N_26013,N_26062);
or U27181 (N_27181,N_26424,N_26760);
nand U27182 (N_27182,N_26284,N_26380);
nand U27183 (N_27183,N_26593,N_26613);
or U27184 (N_27184,N_26580,N_26433);
and U27185 (N_27185,N_26503,N_26724);
or U27186 (N_27186,N_26667,N_26838);
and U27187 (N_27187,N_26141,N_26324);
and U27188 (N_27188,N_26592,N_26876);
and U27189 (N_27189,N_26117,N_26021);
nand U27190 (N_27190,N_26801,N_26251);
or U27191 (N_27191,N_26296,N_26474);
and U27192 (N_27192,N_26011,N_26744);
nor U27193 (N_27193,N_26227,N_26345);
or U27194 (N_27194,N_26990,N_26567);
xnor U27195 (N_27195,N_26289,N_26196);
or U27196 (N_27196,N_26798,N_26797);
nor U27197 (N_27197,N_26941,N_26397);
nand U27198 (N_27198,N_26986,N_26342);
xnor U27199 (N_27199,N_26179,N_26053);
nand U27200 (N_27200,N_26426,N_26850);
and U27201 (N_27201,N_26463,N_26659);
nand U27202 (N_27202,N_26290,N_26601);
nor U27203 (N_27203,N_26887,N_26967);
and U27204 (N_27204,N_26630,N_26871);
nor U27205 (N_27205,N_26136,N_26132);
nand U27206 (N_27206,N_26328,N_26574);
xor U27207 (N_27207,N_26901,N_26678);
or U27208 (N_27208,N_26632,N_26157);
nor U27209 (N_27209,N_26943,N_26948);
nand U27210 (N_27210,N_26947,N_26264);
or U27211 (N_27211,N_26906,N_26088);
nor U27212 (N_27212,N_26535,N_26493);
nor U27213 (N_27213,N_26143,N_26135);
nor U27214 (N_27214,N_26223,N_26989);
nor U27215 (N_27215,N_26467,N_26926);
xnor U27216 (N_27216,N_26211,N_26649);
xnor U27217 (N_27217,N_26304,N_26982);
nand U27218 (N_27218,N_26504,N_26195);
xnor U27219 (N_27219,N_26511,N_26412);
nand U27220 (N_27220,N_26310,N_26362);
or U27221 (N_27221,N_26716,N_26194);
and U27222 (N_27222,N_26643,N_26841);
or U27223 (N_27223,N_26645,N_26102);
nand U27224 (N_27224,N_26846,N_26294);
xnor U27225 (N_27225,N_26644,N_26973);
or U27226 (N_27226,N_26526,N_26369);
or U27227 (N_27227,N_26880,N_26308);
nor U27228 (N_27228,N_26670,N_26647);
and U27229 (N_27229,N_26317,N_26182);
xnor U27230 (N_27230,N_26884,N_26747);
nand U27231 (N_27231,N_26069,N_26758);
and U27232 (N_27232,N_26350,N_26093);
and U27233 (N_27233,N_26790,N_26337);
xor U27234 (N_27234,N_26026,N_26745);
nand U27235 (N_27235,N_26553,N_26598);
or U27236 (N_27236,N_26450,N_26494);
or U27237 (N_27237,N_26844,N_26496);
xor U27238 (N_27238,N_26418,N_26665);
and U27239 (N_27239,N_26084,N_26966);
or U27240 (N_27240,N_26828,N_26155);
and U27241 (N_27241,N_26356,N_26723);
and U27242 (N_27242,N_26629,N_26662);
and U27243 (N_27243,N_26697,N_26808);
and U27244 (N_27244,N_26464,N_26655);
nor U27245 (N_27245,N_26734,N_26525);
and U27246 (N_27246,N_26385,N_26120);
and U27247 (N_27247,N_26717,N_26089);
xor U27248 (N_27248,N_26138,N_26468);
nor U27249 (N_27249,N_26607,N_26110);
nor U27250 (N_27250,N_26244,N_26176);
and U27251 (N_27251,N_26105,N_26455);
and U27252 (N_27252,N_26407,N_26115);
nor U27253 (N_27253,N_26772,N_26778);
nor U27254 (N_27254,N_26318,N_26933);
and U27255 (N_27255,N_26133,N_26177);
and U27256 (N_27256,N_26230,N_26072);
xnor U27257 (N_27257,N_26044,N_26202);
nand U27258 (N_27258,N_26929,N_26752);
nand U27259 (N_27259,N_26388,N_26241);
nor U27260 (N_27260,N_26074,N_26785);
or U27261 (N_27261,N_26010,N_26366);
xnor U27262 (N_27262,N_26419,N_26344);
xnor U27263 (N_27263,N_26743,N_26242);
nand U27264 (N_27264,N_26829,N_26063);
or U27265 (N_27265,N_26932,N_26707);
and U27266 (N_27266,N_26153,N_26742);
or U27267 (N_27267,N_26532,N_26739);
xor U27268 (N_27268,N_26002,N_26207);
and U27269 (N_27269,N_26163,N_26154);
and U27270 (N_27270,N_26442,N_26576);
and U27271 (N_27271,N_26998,N_26786);
nor U27272 (N_27272,N_26950,N_26395);
or U27273 (N_27273,N_26620,N_26288);
nor U27274 (N_27274,N_26368,N_26409);
or U27275 (N_27275,N_26979,N_26325);
nand U27276 (N_27276,N_26487,N_26299);
nor U27277 (N_27277,N_26094,N_26713);
nand U27278 (N_27278,N_26529,N_26485);
nor U27279 (N_27279,N_26403,N_26400);
and U27280 (N_27280,N_26551,N_26387);
nor U27281 (N_27281,N_26691,N_26323);
and U27282 (N_27282,N_26814,N_26606);
or U27283 (N_27283,N_26762,N_26564);
or U27284 (N_27284,N_26098,N_26399);
nand U27285 (N_27285,N_26003,N_26041);
and U27286 (N_27286,N_26746,N_26883);
or U27287 (N_27287,N_26293,N_26935);
xor U27288 (N_27288,N_26951,N_26770);
xor U27289 (N_27289,N_26756,N_26730);
or U27290 (N_27290,N_26637,N_26596);
nor U27291 (N_27291,N_26222,N_26908);
or U27292 (N_27292,N_26271,N_26928);
nand U27293 (N_27293,N_26283,N_26192);
nand U27294 (N_27294,N_26300,N_26940);
nand U27295 (N_27295,N_26204,N_26895);
and U27296 (N_27296,N_26221,N_26675);
nand U27297 (N_27297,N_26197,N_26411);
xor U27298 (N_27298,N_26823,N_26583);
and U27299 (N_27299,N_26231,N_26650);
xnor U27300 (N_27300,N_26286,N_26122);
nor U27301 (N_27301,N_26171,N_26432);
nor U27302 (N_27302,N_26050,N_26902);
and U27303 (N_27303,N_26812,N_26046);
or U27304 (N_27304,N_26247,N_26169);
nand U27305 (N_27305,N_26118,N_26956);
or U27306 (N_27306,N_26009,N_26813);
and U27307 (N_27307,N_26507,N_26992);
or U27308 (N_27308,N_26307,N_26875);
nor U27309 (N_27309,N_26055,N_26075);
or U27310 (N_27310,N_26994,N_26663);
nor U27311 (N_27311,N_26646,N_26833);
or U27312 (N_27312,N_26692,N_26060);
nand U27313 (N_27313,N_26051,N_26444);
and U27314 (N_27314,N_26164,N_26759);
xnor U27315 (N_27315,N_26001,N_26694);
or U27316 (N_27316,N_26953,N_26470);
xnor U27317 (N_27317,N_26699,N_26037);
and U27318 (N_27318,N_26851,N_26000);
and U27319 (N_27319,N_26218,N_26658);
xnor U27320 (N_27320,N_26788,N_26848);
xnor U27321 (N_27321,N_26130,N_26669);
or U27322 (N_27322,N_26638,N_26693);
xnor U27323 (N_27323,N_26769,N_26522);
nand U27324 (N_27324,N_26081,N_26248);
nor U27325 (N_27325,N_26775,N_26621);
or U27326 (N_27326,N_26541,N_26492);
nand U27327 (N_27327,N_26239,N_26536);
nor U27328 (N_27328,N_26761,N_26382);
xnor U27329 (N_27329,N_26753,N_26184);
nand U27330 (N_27330,N_26090,N_26898);
xor U27331 (N_27331,N_26793,N_26477);
nor U27332 (N_27332,N_26429,N_26107);
nand U27333 (N_27333,N_26420,N_26506);
and U27334 (N_27334,N_26134,N_26917);
or U27335 (N_27335,N_26077,N_26991);
or U27336 (N_27336,N_26909,N_26519);
nor U27337 (N_27337,N_26199,N_26664);
nor U27338 (N_27338,N_26768,N_26162);
nor U27339 (N_27339,N_26214,N_26708);
xor U27340 (N_27340,N_26466,N_26034);
and U27341 (N_27341,N_26524,N_26577);
nand U27342 (N_27342,N_26501,N_26698);
and U27343 (N_27343,N_26364,N_26206);
or U27344 (N_27344,N_26291,N_26836);
and U27345 (N_27345,N_26729,N_26641);
and U27346 (N_27346,N_26869,N_26261);
and U27347 (N_27347,N_26878,N_26893);
nor U27348 (N_27348,N_26249,N_26104);
or U27349 (N_27349,N_26546,N_26166);
nor U27350 (N_27350,N_26173,N_26258);
nand U27351 (N_27351,N_26059,N_26398);
nand U27352 (N_27352,N_26794,N_26217);
nand U27353 (N_27353,N_26351,N_26888);
nor U27354 (N_27354,N_26040,N_26702);
xor U27355 (N_27355,N_26852,N_26421);
and U27356 (N_27356,N_26322,N_26651);
nor U27357 (N_27357,N_26393,N_26885);
and U27358 (N_27358,N_26712,N_26984);
nand U27359 (N_27359,N_26158,N_26811);
nor U27360 (N_27360,N_26611,N_26151);
or U27361 (N_27361,N_26937,N_26097);
nor U27362 (N_27362,N_26225,N_26360);
nand U27363 (N_27363,N_26572,N_26854);
or U27364 (N_27364,N_26859,N_26457);
nand U27365 (N_27365,N_26996,N_26981);
xor U27366 (N_27366,N_26864,N_26703);
or U27367 (N_27367,N_26861,N_26028);
xor U27368 (N_27368,N_26180,N_26314);
or U27369 (N_27369,N_26475,N_26648);
or U27370 (N_27370,N_26147,N_26279);
and U27371 (N_27371,N_26346,N_26127);
or U27372 (N_27372,N_26185,N_26671);
nor U27373 (N_27373,N_26974,N_26603);
and U27374 (N_27374,N_26148,N_26390);
nor U27375 (N_27375,N_26866,N_26391);
nand U27376 (N_27376,N_26964,N_26822);
nor U27377 (N_27377,N_26987,N_26236);
or U27378 (N_27378,N_26267,N_26246);
nor U27379 (N_27379,N_26125,N_26020);
or U27380 (N_27380,N_26571,N_26447);
nand U27381 (N_27381,N_26983,N_26448);
nand U27382 (N_27382,N_26038,N_26873);
or U27383 (N_27383,N_26022,N_26608);
nand U27384 (N_27384,N_26617,N_26139);
xor U27385 (N_27385,N_26867,N_26263);
xor U27386 (N_27386,N_26233,N_26657);
or U27387 (N_27387,N_26714,N_26352);
nor U27388 (N_27388,N_26178,N_26980);
nor U27389 (N_27389,N_26483,N_26774);
nand U27390 (N_27390,N_26065,N_26058);
and U27391 (N_27391,N_26087,N_26491);
or U27392 (N_27392,N_26795,N_26554);
or U27393 (N_27393,N_26389,N_26642);
and U27394 (N_27394,N_26727,N_26334);
and U27395 (N_27395,N_26530,N_26513);
nand U27396 (N_27396,N_26355,N_26095);
and U27397 (N_27397,N_26321,N_26331);
xnor U27398 (N_27398,N_26903,N_26298);
or U27399 (N_27399,N_26581,N_26482);
nand U27400 (N_27400,N_26377,N_26715);
or U27401 (N_27401,N_26476,N_26408);
and U27402 (N_27402,N_26573,N_26700);
xnor U27403 (N_27403,N_26879,N_26858);
xor U27404 (N_27404,N_26988,N_26894);
or U27405 (N_27405,N_26633,N_26434);
nor U27406 (N_27406,N_26295,N_26061);
or U27407 (N_27407,N_26030,N_26068);
nand U27408 (N_27408,N_26736,N_26144);
and U27409 (N_27409,N_26416,N_26549);
or U27410 (N_27410,N_26237,N_26750);
xnor U27411 (N_27411,N_26392,N_26531);
nand U27412 (N_27412,N_26591,N_26100);
xnor U27413 (N_27413,N_26900,N_26542);
nor U27414 (N_27414,N_26338,N_26116);
nand U27415 (N_27415,N_26685,N_26799);
nor U27416 (N_27416,N_26877,N_26582);
and U27417 (N_27417,N_26537,N_26486);
nand U27418 (N_27418,N_26881,N_26423);
or U27419 (N_27419,N_26431,N_26688);
or U27420 (N_27420,N_26807,N_26330);
or U27421 (N_27421,N_26628,N_26336);
xor U27422 (N_27422,N_26818,N_26126);
nand U27423 (N_27423,N_26622,N_26384);
nand U27424 (N_27424,N_26627,N_26404);
or U27425 (N_27425,N_26066,N_26333);
nand U27426 (N_27426,N_26035,N_26460);
nand U27427 (N_27427,N_26776,N_26452);
or U27428 (N_27428,N_26971,N_26985);
and U27429 (N_27429,N_26856,N_26170);
nand U27430 (N_27430,N_26064,N_26440);
and U27431 (N_27431,N_26640,N_26287);
nor U27432 (N_27432,N_26276,N_26213);
xor U27433 (N_27433,N_26976,N_26849);
xor U27434 (N_27434,N_26936,N_26896);
nand U27435 (N_27435,N_26243,N_26520);
nor U27436 (N_27436,N_26301,N_26738);
xnor U27437 (N_27437,N_26453,N_26805);
or U27438 (N_27438,N_26371,N_26149);
and U27439 (N_27439,N_26792,N_26722);
and U27440 (N_27440,N_26765,N_26108);
nand U27441 (N_27441,N_26234,N_26783);
and U27442 (N_27442,N_26085,N_26007);
nand U27443 (N_27443,N_26905,N_26252);
nand U27444 (N_27444,N_26373,N_26319);
and U27445 (N_27445,N_26547,N_26274);
and U27446 (N_27446,N_26754,N_26706);
or U27447 (N_27447,N_26847,N_26683);
nor U27448 (N_27448,N_26190,N_26614);
xor U27449 (N_27449,N_26361,N_26168);
or U27450 (N_27450,N_26259,N_26047);
nand U27451 (N_27451,N_26921,N_26939);
nor U27452 (N_27452,N_26764,N_26480);
nor U27453 (N_27453,N_26198,N_26262);
xnor U27454 (N_27454,N_26459,N_26112);
nand U27455 (N_27455,N_26297,N_26353);
xnor U27456 (N_27456,N_26091,N_26784);
xnor U27457 (N_27457,N_26725,N_26320);
xor U27458 (N_27458,N_26913,N_26303);
nor U27459 (N_27459,N_26478,N_26436);
nand U27460 (N_27460,N_26015,N_26777);
nor U27461 (N_27461,N_26931,N_26260);
xor U27462 (N_27462,N_26687,N_26919);
xor U27463 (N_27463,N_26113,N_26533);
and U27464 (N_27464,N_26938,N_26256);
or U27465 (N_27465,N_26955,N_26489);
xor U27466 (N_27466,N_26285,N_26690);
or U27467 (N_27467,N_26925,N_26370);
and U27468 (N_27468,N_26129,N_26957);
and U27469 (N_27469,N_26273,N_26839);
xnor U27470 (N_27470,N_26963,N_26266);
xnor U27471 (N_27471,N_26728,N_26441);
xor U27472 (N_27472,N_26652,N_26661);
xor U27473 (N_27473,N_26718,N_26891);
nand U27474 (N_27474,N_26484,N_26635);
nor U27475 (N_27475,N_26609,N_26825);
and U27476 (N_27476,N_26680,N_26550);
nand U27477 (N_27477,N_26827,N_26193);
nor U27478 (N_27478,N_26626,N_26523);
nor U27479 (N_27479,N_26965,N_26860);
and U27480 (N_27480,N_26555,N_26372);
or U27481 (N_27481,N_26438,N_26958);
xnor U27482 (N_27482,N_26018,N_26024);
and U27483 (N_27483,N_26538,N_26186);
nor U27484 (N_27484,N_26329,N_26339);
or U27485 (N_27485,N_26512,N_26946);
and U27486 (N_27486,N_26588,N_26315);
and U27487 (N_27487,N_26802,N_26332);
xnor U27488 (N_27488,N_26624,N_26305);
xor U27489 (N_27489,N_26924,N_26863);
nor U27490 (N_27490,N_26099,N_26076);
or U27491 (N_27491,N_26235,N_26150);
nor U27492 (N_27492,N_26892,N_26354);
nor U27493 (N_27493,N_26952,N_26381);
xor U27494 (N_27494,N_26815,N_26042);
nor U27495 (N_27495,N_26872,N_26540);
and U27496 (N_27496,N_26006,N_26570);
and U27497 (N_27497,N_26731,N_26920);
nand U27498 (N_27498,N_26552,N_26057);
and U27499 (N_27499,N_26465,N_26631);
nand U27500 (N_27500,N_26843,N_26891);
or U27501 (N_27501,N_26425,N_26092);
and U27502 (N_27502,N_26090,N_26161);
or U27503 (N_27503,N_26872,N_26376);
nor U27504 (N_27504,N_26809,N_26773);
or U27505 (N_27505,N_26875,N_26268);
and U27506 (N_27506,N_26578,N_26918);
nand U27507 (N_27507,N_26031,N_26787);
nor U27508 (N_27508,N_26850,N_26270);
xor U27509 (N_27509,N_26999,N_26757);
nor U27510 (N_27510,N_26283,N_26476);
xor U27511 (N_27511,N_26239,N_26297);
and U27512 (N_27512,N_26629,N_26327);
or U27513 (N_27513,N_26822,N_26588);
or U27514 (N_27514,N_26683,N_26109);
or U27515 (N_27515,N_26834,N_26653);
and U27516 (N_27516,N_26272,N_26612);
and U27517 (N_27517,N_26456,N_26552);
nand U27518 (N_27518,N_26729,N_26812);
or U27519 (N_27519,N_26123,N_26013);
nor U27520 (N_27520,N_26042,N_26802);
xnor U27521 (N_27521,N_26812,N_26147);
and U27522 (N_27522,N_26708,N_26351);
nor U27523 (N_27523,N_26860,N_26865);
or U27524 (N_27524,N_26662,N_26970);
and U27525 (N_27525,N_26504,N_26835);
and U27526 (N_27526,N_26175,N_26332);
nand U27527 (N_27527,N_26308,N_26159);
nor U27528 (N_27528,N_26443,N_26809);
xnor U27529 (N_27529,N_26131,N_26039);
nand U27530 (N_27530,N_26897,N_26661);
nand U27531 (N_27531,N_26998,N_26004);
and U27532 (N_27532,N_26650,N_26099);
or U27533 (N_27533,N_26606,N_26829);
nand U27534 (N_27534,N_26483,N_26392);
nor U27535 (N_27535,N_26039,N_26260);
or U27536 (N_27536,N_26197,N_26302);
xnor U27537 (N_27537,N_26246,N_26629);
or U27538 (N_27538,N_26068,N_26647);
or U27539 (N_27539,N_26929,N_26539);
nor U27540 (N_27540,N_26861,N_26653);
xor U27541 (N_27541,N_26690,N_26185);
nand U27542 (N_27542,N_26719,N_26065);
xor U27543 (N_27543,N_26855,N_26046);
nor U27544 (N_27544,N_26552,N_26250);
nor U27545 (N_27545,N_26195,N_26245);
xnor U27546 (N_27546,N_26109,N_26445);
or U27547 (N_27547,N_26343,N_26889);
xnor U27548 (N_27548,N_26099,N_26955);
or U27549 (N_27549,N_26338,N_26436);
or U27550 (N_27550,N_26231,N_26965);
xnor U27551 (N_27551,N_26918,N_26633);
nor U27552 (N_27552,N_26020,N_26279);
and U27553 (N_27553,N_26664,N_26029);
nand U27554 (N_27554,N_26326,N_26084);
or U27555 (N_27555,N_26273,N_26133);
xor U27556 (N_27556,N_26189,N_26477);
nand U27557 (N_27557,N_26444,N_26609);
nand U27558 (N_27558,N_26232,N_26976);
and U27559 (N_27559,N_26151,N_26906);
or U27560 (N_27560,N_26793,N_26610);
nor U27561 (N_27561,N_26876,N_26995);
nor U27562 (N_27562,N_26486,N_26529);
xor U27563 (N_27563,N_26505,N_26774);
nor U27564 (N_27564,N_26402,N_26235);
nand U27565 (N_27565,N_26751,N_26680);
or U27566 (N_27566,N_26571,N_26490);
xnor U27567 (N_27567,N_26373,N_26404);
and U27568 (N_27568,N_26797,N_26104);
xor U27569 (N_27569,N_26554,N_26081);
or U27570 (N_27570,N_26465,N_26374);
xor U27571 (N_27571,N_26658,N_26001);
or U27572 (N_27572,N_26223,N_26788);
or U27573 (N_27573,N_26779,N_26184);
nor U27574 (N_27574,N_26890,N_26925);
or U27575 (N_27575,N_26462,N_26548);
or U27576 (N_27576,N_26381,N_26342);
nand U27577 (N_27577,N_26194,N_26871);
nor U27578 (N_27578,N_26237,N_26497);
nor U27579 (N_27579,N_26143,N_26985);
nand U27580 (N_27580,N_26869,N_26274);
or U27581 (N_27581,N_26106,N_26526);
xnor U27582 (N_27582,N_26642,N_26238);
xor U27583 (N_27583,N_26772,N_26802);
or U27584 (N_27584,N_26016,N_26972);
xor U27585 (N_27585,N_26314,N_26890);
and U27586 (N_27586,N_26381,N_26143);
nor U27587 (N_27587,N_26906,N_26036);
nor U27588 (N_27588,N_26532,N_26668);
or U27589 (N_27589,N_26798,N_26674);
and U27590 (N_27590,N_26760,N_26832);
nor U27591 (N_27591,N_26688,N_26174);
xnor U27592 (N_27592,N_26081,N_26630);
nor U27593 (N_27593,N_26013,N_26282);
xnor U27594 (N_27594,N_26860,N_26479);
or U27595 (N_27595,N_26796,N_26358);
nand U27596 (N_27596,N_26377,N_26563);
nand U27597 (N_27597,N_26990,N_26371);
xor U27598 (N_27598,N_26032,N_26146);
nor U27599 (N_27599,N_26854,N_26344);
or U27600 (N_27600,N_26943,N_26432);
nand U27601 (N_27601,N_26784,N_26136);
nor U27602 (N_27602,N_26169,N_26957);
nand U27603 (N_27603,N_26010,N_26870);
nor U27604 (N_27604,N_26584,N_26229);
or U27605 (N_27605,N_26488,N_26868);
nor U27606 (N_27606,N_26806,N_26001);
nand U27607 (N_27607,N_26882,N_26863);
nand U27608 (N_27608,N_26082,N_26151);
xor U27609 (N_27609,N_26897,N_26358);
xnor U27610 (N_27610,N_26604,N_26687);
nor U27611 (N_27611,N_26215,N_26002);
and U27612 (N_27612,N_26989,N_26732);
nand U27613 (N_27613,N_26573,N_26156);
nand U27614 (N_27614,N_26443,N_26247);
nor U27615 (N_27615,N_26474,N_26627);
xnor U27616 (N_27616,N_26415,N_26134);
and U27617 (N_27617,N_26632,N_26020);
or U27618 (N_27618,N_26236,N_26758);
nand U27619 (N_27619,N_26402,N_26478);
xnor U27620 (N_27620,N_26380,N_26831);
nor U27621 (N_27621,N_26745,N_26576);
nand U27622 (N_27622,N_26407,N_26645);
nand U27623 (N_27623,N_26014,N_26790);
xor U27624 (N_27624,N_26110,N_26559);
and U27625 (N_27625,N_26190,N_26156);
nand U27626 (N_27626,N_26775,N_26671);
or U27627 (N_27627,N_26747,N_26659);
or U27628 (N_27628,N_26971,N_26925);
and U27629 (N_27629,N_26599,N_26843);
or U27630 (N_27630,N_26828,N_26592);
nor U27631 (N_27631,N_26478,N_26062);
and U27632 (N_27632,N_26892,N_26288);
and U27633 (N_27633,N_26667,N_26013);
or U27634 (N_27634,N_26715,N_26141);
and U27635 (N_27635,N_26927,N_26502);
nand U27636 (N_27636,N_26141,N_26875);
nor U27637 (N_27637,N_26991,N_26032);
xnor U27638 (N_27638,N_26912,N_26844);
xnor U27639 (N_27639,N_26559,N_26208);
and U27640 (N_27640,N_26838,N_26918);
or U27641 (N_27641,N_26159,N_26833);
nor U27642 (N_27642,N_26222,N_26355);
or U27643 (N_27643,N_26418,N_26097);
nor U27644 (N_27644,N_26818,N_26025);
nor U27645 (N_27645,N_26151,N_26859);
xor U27646 (N_27646,N_26564,N_26691);
nor U27647 (N_27647,N_26368,N_26899);
nand U27648 (N_27648,N_26872,N_26100);
or U27649 (N_27649,N_26250,N_26784);
xor U27650 (N_27650,N_26891,N_26937);
xor U27651 (N_27651,N_26213,N_26062);
nand U27652 (N_27652,N_26854,N_26117);
or U27653 (N_27653,N_26018,N_26431);
nor U27654 (N_27654,N_26180,N_26761);
and U27655 (N_27655,N_26981,N_26555);
xnor U27656 (N_27656,N_26646,N_26533);
nand U27657 (N_27657,N_26293,N_26791);
or U27658 (N_27658,N_26036,N_26094);
xor U27659 (N_27659,N_26620,N_26054);
nand U27660 (N_27660,N_26585,N_26998);
or U27661 (N_27661,N_26740,N_26784);
or U27662 (N_27662,N_26950,N_26772);
nor U27663 (N_27663,N_26945,N_26683);
nand U27664 (N_27664,N_26093,N_26263);
nand U27665 (N_27665,N_26051,N_26583);
and U27666 (N_27666,N_26531,N_26556);
nand U27667 (N_27667,N_26405,N_26755);
xor U27668 (N_27668,N_26906,N_26755);
nor U27669 (N_27669,N_26918,N_26749);
nor U27670 (N_27670,N_26230,N_26067);
nor U27671 (N_27671,N_26866,N_26206);
nand U27672 (N_27672,N_26561,N_26173);
or U27673 (N_27673,N_26505,N_26297);
xnor U27674 (N_27674,N_26585,N_26697);
and U27675 (N_27675,N_26880,N_26892);
or U27676 (N_27676,N_26128,N_26561);
or U27677 (N_27677,N_26147,N_26187);
nor U27678 (N_27678,N_26035,N_26420);
nor U27679 (N_27679,N_26307,N_26789);
nor U27680 (N_27680,N_26459,N_26665);
and U27681 (N_27681,N_26371,N_26262);
or U27682 (N_27682,N_26504,N_26143);
nor U27683 (N_27683,N_26676,N_26519);
xnor U27684 (N_27684,N_26849,N_26402);
and U27685 (N_27685,N_26728,N_26965);
or U27686 (N_27686,N_26304,N_26574);
and U27687 (N_27687,N_26599,N_26887);
nand U27688 (N_27688,N_26693,N_26408);
xnor U27689 (N_27689,N_26828,N_26563);
xnor U27690 (N_27690,N_26194,N_26005);
nand U27691 (N_27691,N_26133,N_26617);
nor U27692 (N_27692,N_26364,N_26299);
nand U27693 (N_27693,N_26923,N_26993);
xnor U27694 (N_27694,N_26815,N_26032);
nor U27695 (N_27695,N_26855,N_26498);
nand U27696 (N_27696,N_26523,N_26943);
xnor U27697 (N_27697,N_26649,N_26272);
nand U27698 (N_27698,N_26331,N_26058);
and U27699 (N_27699,N_26613,N_26963);
or U27700 (N_27700,N_26051,N_26957);
nor U27701 (N_27701,N_26862,N_26721);
nor U27702 (N_27702,N_26633,N_26540);
or U27703 (N_27703,N_26064,N_26071);
and U27704 (N_27704,N_26773,N_26846);
nand U27705 (N_27705,N_26883,N_26361);
or U27706 (N_27706,N_26278,N_26094);
nor U27707 (N_27707,N_26985,N_26205);
and U27708 (N_27708,N_26953,N_26578);
nor U27709 (N_27709,N_26750,N_26726);
nor U27710 (N_27710,N_26267,N_26397);
nand U27711 (N_27711,N_26634,N_26998);
and U27712 (N_27712,N_26971,N_26710);
and U27713 (N_27713,N_26628,N_26580);
and U27714 (N_27714,N_26533,N_26240);
nand U27715 (N_27715,N_26610,N_26625);
nor U27716 (N_27716,N_26925,N_26102);
or U27717 (N_27717,N_26162,N_26454);
or U27718 (N_27718,N_26798,N_26080);
and U27719 (N_27719,N_26641,N_26786);
nand U27720 (N_27720,N_26609,N_26110);
or U27721 (N_27721,N_26786,N_26293);
and U27722 (N_27722,N_26760,N_26599);
and U27723 (N_27723,N_26317,N_26380);
xnor U27724 (N_27724,N_26974,N_26944);
nand U27725 (N_27725,N_26713,N_26930);
nor U27726 (N_27726,N_26971,N_26009);
or U27727 (N_27727,N_26546,N_26368);
xnor U27728 (N_27728,N_26005,N_26957);
nor U27729 (N_27729,N_26969,N_26313);
nor U27730 (N_27730,N_26956,N_26392);
nor U27731 (N_27731,N_26479,N_26233);
or U27732 (N_27732,N_26614,N_26111);
and U27733 (N_27733,N_26496,N_26124);
xor U27734 (N_27734,N_26607,N_26074);
xnor U27735 (N_27735,N_26905,N_26982);
or U27736 (N_27736,N_26402,N_26214);
nand U27737 (N_27737,N_26039,N_26842);
or U27738 (N_27738,N_26338,N_26604);
nand U27739 (N_27739,N_26369,N_26398);
and U27740 (N_27740,N_26304,N_26406);
or U27741 (N_27741,N_26712,N_26129);
and U27742 (N_27742,N_26953,N_26027);
and U27743 (N_27743,N_26733,N_26204);
xor U27744 (N_27744,N_26427,N_26803);
and U27745 (N_27745,N_26426,N_26781);
nand U27746 (N_27746,N_26563,N_26050);
xor U27747 (N_27747,N_26152,N_26512);
and U27748 (N_27748,N_26427,N_26062);
and U27749 (N_27749,N_26762,N_26821);
xor U27750 (N_27750,N_26440,N_26642);
or U27751 (N_27751,N_26383,N_26785);
and U27752 (N_27752,N_26219,N_26110);
nor U27753 (N_27753,N_26034,N_26839);
and U27754 (N_27754,N_26980,N_26117);
or U27755 (N_27755,N_26055,N_26445);
nor U27756 (N_27756,N_26734,N_26967);
or U27757 (N_27757,N_26942,N_26909);
and U27758 (N_27758,N_26632,N_26346);
or U27759 (N_27759,N_26244,N_26205);
nand U27760 (N_27760,N_26563,N_26898);
or U27761 (N_27761,N_26887,N_26546);
nand U27762 (N_27762,N_26117,N_26984);
xor U27763 (N_27763,N_26504,N_26467);
or U27764 (N_27764,N_26177,N_26041);
xor U27765 (N_27765,N_26006,N_26875);
xnor U27766 (N_27766,N_26271,N_26277);
xor U27767 (N_27767,N_26511,N_26246);
or U27768 (N_27768,N_26183,N_26863);
or U27769 (N_27769,N_26722,N_26988);
xnor U27770 (N_27770,N_26804,N_26979);
nand U27771 (N_27771,N_26524,N_26558);
nand U27772 (N_27772,N_26972,N_26917);
nand U27773 (N_27773,N_26829,N_26518);
nor U27774 (N_27774,N_26915,N_26376);
nand U27775 (N_27775,N_26100,N_26088);
xnor U27776 (N_27776,N_26252,N_26561);
nand U27777 (N_27777,N_26830,N_26628);
or U27778 (N_27778,N_26783,N_26354);
nor U27779 (N_27779,N_26868,N_26064);
xor U27780 (N_27780,N_26887,N_26016);
and U27781 (N_27781,N_26586,N_26888);
or U27782 (N_27782,N_26003,N_26375);
and U27783 (N_27783,N_26161,N_26740);
nor U27784 (N_27784,N_26617,N_26925);
nand U27785 (N_27785,N_26012,N_26144);
or U27786 (N_27786,N_26723,N_26859);
xnor U27787 (N_27787,N_26266,N_26228);
or U27788 (N_27788,N_26296,N_26936);
xor U27789 (N_27789,N_26398,N_26876);
nand U27790 (N_27790,N_26584,N_26390);
and U27791 (N_27791,N_26620,N_26606);
and U27792 (N_27792,N_26869,N_26041);
and U27793 (N_27793,N_26325,N_26051);
xor U27794 (N_27794,N_26225,N_26737);
nor U27795 (N_27795,N_26167,N_26895);
xor U27796 (N_27796,N_26175,N_26176);
nor U27797 (N_27797,N_26949,N_26880);
and U27798 (N_27798,N_26438,N_26704);
nand U27799 (N_27799,N_26226,N_26436);
nor U27800 (N_27800,N_26943,N_26828);
nor U27801 (N_27801,N_26466,N_26626);
and U27802 (N_27802,N_26128,N_26824);
nor U27803 (N_27803,N_26255,N_26663);
xor U27804 (N_27804,N_26968,N_26733);
nand U27805 (N_27805,N_26960,N_26828);
xor U27806 (N_27806,N_26058,N_26041);
and U27807 (N_27807,N_26824,N_26291);
xnor U27808 (N_27808,N_26010,N_26712);
or U27809 (N_27809,N_26967,N_26854);
nor U27810 (N_27810,N_26636,N_26750);
nand U27811 (N_27811,N_26302,N_26138);
or U27812 (N_27812,N_26125,N_26699);
nor U27813 (N_27813,N_26361,N_26314);
or U27814 (N_27814,N_26217,N_26308);
or U27815 (N_27815,N_26671,N_26990);
or U27816 (N_27816,N_26615,N_26560);
nand U27817 (N_27817,N_26906,N_26183);
nor U27818 (N_27818,N_26052,N_26001);
xor U27819 (N_27819,N_26513,N_26902);
nor U27820 (N_27820,N_26512,N_26994);
nor U27821 (N_27821,N_26294,N_26795);
xnor U27822 (N_27822,N_26713,N_26995);
nor U27823 (N_27823,N_26281,N_26196);
nand U27824 (N_27824,N_26460,N_26304);
xnor U27825 (N_27825,N_26651,N_26940);
nand U27826 (N_27826,N_26913,N_26601);
xnor U27827 (N_27827,N_26200,N_26035);
nand U27828 (N_27828,N_26939,N_26197);
nor U27829 (N_27829,N_26525,N_26480);
and U27830 (N_27830,N_26790,N_26110);
and U27831 (N_27831,N_26347,N_26175);
nand U27832 (N_27832,N_26844,N_26579);
and U27833 (N_27833,N_26193,N_26749);
xnor U27834 (N_27834,N_26751,N_26104);
xnor U27835 (N_27835,N_26877,N_26931);
nor U27836 (N_27836,N_26976,N_26952);
nand U27837 (N_27837,N_26584,N_26210);
xor U27838 (N_27838,N_26297,N_26260);
nor U27839 (N_27839,N_26518,N_26791);
nand U27840 (N_27840,N_26718,N_26593);
xor U27841 (N_27841,N_26445,N_26680);
nor U27842 (N_27842,N_26717,N_26401);
xnor U27843 (N_27843,N_26784,N_26604);
xnor U27844 (N_27844,N_26028,N_26740);
nor U27845 (N_27845,N_26921,N_26167);
xor U27846 (N_27846,N_26987,N_26853);
and U27847 (N_27847,N_26640,N_26917);
nor U27848 (N_27848,N_26237,N_26478);
xnor U27849 (N_27849,N_26910,N_26236);
or U27850 (N_27850,N_26503,N_26983);
nor U27851 (N_27851,N_26740,N_26513);
and U27852 (N_27852,N_26236,N_26964);
nor U27853 (N_27853,N_26756,N_26422);
or U27854 (N_27854,N_26317,N_26191);
xor U27855 (N_27855,N_26971,N_26923);
nand U27856 (N_27856,N_26039,N_26373);
and U27857 (N_27857,N_26028,N_26285);
and U27858 (N_27858,N_26119,N_26560);
and U27859 (N_27859,N_26856,N_26068);
and U27860 (N_27860,N_26791,N_26743);
xnor U27861 (N_27861,N_26772,N_26924);
nand U27862 (N_27862,N_26677,N_26184);
and U27863 (N_27863,N_26592,N_26184);
nand U27864 (N_27864,N_26319,N_26242);
xnor U27865 (N_27865,N_26624,N_26343);
nand U27866 (N_27866,N_26295,N_26741);
or U27867 (N_27867,N_26335,N_26757);
and U27868 (N_27868,N_26125,N_26061);
nand U27869 (N_27869,N_26883,N_26378);
and U27870 (N_27870,N_26960,N_26741);
or U27871 (N_27871,N_26313,N_26866);
xor U27872 (N_27872,N_26904,N_26760);
and U27873 (N_27873,N_26245,N_26580);
and U27874 (N_27874,N_26836,N_26195);
and U27875 (N_27875,N_26847,N_26017);
or U27876 (N_27876,N_26940,N_26595);
and U27877 (N_27877,N_26496,N_26685);
and U27878 (N_27878,N_26002,N_26116);
xor U27879 (N_27879,N_26596,N_26902);
nor U27880 (N_27880,N_26008,N_26207);
nand U27881 (N_27881,N_26406,N_26411);
nand U27882 (N_27882,N_26768,N_26538);
nor U27883 (N_27883,N_26731,N_26381);
or U27884 (N_27884,N_26598,N_26986);
nor U27885 (N_27885,N_26804,N_26389);
nand U27886 (N_27886,N_26292,N_26241);
or U27887 (N_27887,N_26804,N_26960);
nor U27888 (N_27888,N_26933,N_26835);
nor U27889 (N_27889,N_26713,N_26659);
and U27890 (N_27890,N_26226,N_26405);
nand U27891 (N_27891,N_26142,N_26126);
or U27892 (N_27892,N_26956,N_26709);
xor U27893 (N_27893,N_26749,N_26272);
nand U27894 (N_27894,N_26101,N_26553);
xor U27895 (N_27895,N_26048,N_26621);
xnor U27896 (N_27896,N_26445,N_26571);
xor U27897 (N_27897,N_26908,N_26932);
and U27898 (N_27898,N_26718,N_26723);
nand U27899 (N_27899,N_26842,N_26511);
xor U27900 (N_27900,N_26272,N_26192);
xor U27901 (N_27901,N_26012,N_26745);
nor U27902 (N_27902,N_26940,N_26694);
and U27903 (N_27903,N_26862,N_26640);
and U27904 (N_27904,N_26777,N_26464);
nand U27905 (N_27905,N_26448,N_26176);
nor U27906 (N_27906,N_26138,N_26522);
nand U27907 (N_27907,N_26879,N_26188);
nand U27908 (N_27908,N_26522,N_26529);
or U27909 (N_27909,N_26953,N_26216);
or U27910 (N_27910,N_26359,N_26720);
and U27911 (N_27911,N_26012,N_26334);
or U27912 (N_27912,N_26067,N_26524);
or U27913 (N_27913,N_26909,N_26963);
or U27914 (N_27914,N_26671,N_26238);
or U27915 (N_27915,N_26924,N_26560);
or U27916 (N_27916,N_26820,N_26754);
nand U27917 (N_27917,N_26739,N_26289);
xnor U27918 (N_27918,N_26583,N_26748);
or U27919 (N_27919,N_26250,N_26646);
nor U27920 (N_27920,N_26588,N_26383);
nor U27921 (N_27921,N_26955,N_26409);
nand U27922 (N_27922,N_26678,N_26329);
xnor U27923 (N_27923,N_26934,N_26724);
and U27924 (N_27924,N_26526,N_26291);
and U27925 (N_27925,N_26654,N_26899);
and U27926 (N_27926,N_26723,N_26572);
nor U27927 (N_27927,N_26579,N_26330);
nand U27928 (N_27928,N_26668,N_26699);
nand U27929 (N_27929,N_26905,N_26664);
or U27930 (N_27930,N_26706,N_26381);
nand U27931 (N_27931,N_26772,N_26818);
xor U27932 (N_27932,N_26731,N_26227);
nor U27933 (N_27933,N_26906,N_26152);
nor U27934 (N_27934,N_26709,N_26103);
nor U27935 (N_27935,N_26289,N_26279);
xor U27936 (N_27936,N_26417,N_26889);
nand U27937 (N_27937,N_26307,N_26447);
xnor U27938 (N_27938,N_26439,N_26893);
xor U27939 (N_27939,N_26254,N_26919);
and U27940 (N_27940,N_26232,N_26930);
nor U27941 (N_27941,N_26254,N_26448);
nor U27942 (N_27942,N_26414,N_26397);
or U27943 (N_27943,N_26182,N_26483);
xnor U27944 (N_27944,N_26480,N_26768);
nor U27945 (N_27945,N_26980,N_26402);
nor U27946 (N_27946,N_26438,N_26168);
nand U27947 (N_27947,N_26454,N_26506);
and U27948 (N_27948,N_26823,N_26912);
or U27949 (N_27949,N_26155,N_26638);
nor U27950 (N_27950,N_26596,N_26678);
and U27951 (N_27951,N_26575,N_26176);
nand U27952 (N_27952,N_26762,N_26693);
nor U27953 (N_27953,N_26312,N_26848);
nor U27954 (N_27954,N_26138,N_26110);
nand U27955 (N_27955,N_26477,N_26698);
xnor U27956 (N_27956,N_26728,N_26480);
nand U27957 (N_27957,N_26327,N_26586);
nand U27958 (N_27958,N_26627,N_26581);
and U27959 (N_27959,N_26454,N_26895);
xnor U27960 (N_27960,N_26674,N_26950);
nor U27961 (N_27961,N_26579,N_26919);
nand U27962 (N_27962,N_26332,N_26746);
xnor U27963 (N_27963,N_26238,N_26388);
or U27964 (N_27964,N_26070,N_26553);
or U27965 (N_27965,N_26257,N_26804);
nor U27966 (N_27966,N_26115,N_26060);
nand U27967 (N_27967,N_26134,N_26591);
nor U27968 (N_27968,N_26910,N_26961);
nand U27969 (N_27969,N_26365,N_26635);
xor U27970 (N_27970,N_26666,N_26646);
xnor U27971 (N_27971,N_26396,N_26102);
nor U27972 (N_27972,N_26554,N_26899);
nor U27973 (N_27973,N_26107,N_26505);
xor U27974 (N_27974,N_26888,N_26080);
nor U27975 (N_27975,N_26835,N_26347);
and U27976 (N_27976,N_26505,N_26298);
or U27977 (N_27977,N_26859,N_26233);
and U27978 (N_27978,N_26900,N_26895);
and U27979 (N_27979,N_26872,N_26724);
nor U27980 (N_27980,N_26216,N_26240);
or U27981 (N_27981,N_26412,N_26602);
nor U27982 (N_27982,N_26007,N_26986);
nand U27983 (N_27983,N_26366,N_26421);
or U27984 (N_27984,N_26398,N_26368);
and U27985 (N_27985,N_26854,N_26769);
nor U27986 (N_27986,N_26356,N_26322);
nand U27987 (N_27987,N_26995,N_26469);
xor U27988 (N_27988,N_26508,N_26525);
or U27989 (N_27989,N_26606,N_26330);
nand U27990 (N_27990,N_26790,N_26567);
nand U27991 (N_27991,N_26898,N_26684);
nand U27992 (N_27992,N_26422,N_26132);
and U27993 (N_27993,N_26177,N_26619);
or U27994 (N_27994,N_26341,N_26308);
nand U27995 (N_27995,N_26060,N_26722);
and U27996 (N_27996,N_26808,N_26599);
nor U27997 (N_27997,N_26376,N_26195);
or U27998 (N_27998,N_26850,N_26347);
and U27999 (N_27999,N_26760,N_26087);
xor U28000 (N_28000,N_27253,N_27394);
xor U28001 (N_28001,N_27134,N_27649);
xnor U28002 (N_28002,N_27207,N_27668);
nand U28003 (N_28003,N_27202,N_27659);
nor U28004 (N_28004,N_27320,N_27452);
nor U28005 (N_28005,N_27525,N_27030);
or U28006 (N_28006,N_27069,N_27203);
and U28007 (N_28007,N_27157,N_27606);
or U28008 (N_28008,N_27964,N_27699);
and U28009 (N_28009,N_27067,N_27095);
xor U28010 (N_28010,N_27573,N_27513);
or U28011 (N_28011,N_27379,N_27053);
xor U28012 (N_28012,N_27881,N_27289);
nor U28013 (N_28013,N_27671,N_27152);
nand U28014 (N_28014,N_27988,N_27776);
nand U28015 (N_28015,N_27862,N_27024);
xnor U28016 (N_28016,N_27901,N_27723);
nor U28017 (N_28017,N_27799,N_27651);
or U28018 (N_28018,N_27204,N_27883);
xnor U28019 (N_28019,N_27488,N_27623);
and U28020 (N_28020,N_27822,N_27821);
nand U28021 (N_28021,N_27762,N_27811);
nor U28022 (N_28022,N_27629,N_27419);
nor U28023 (N_28023,N_27866,N_27459);
or U28024 (N_28024,N_27630,N_27820);
or U28025 (N_28025,N_27354,N_27605);
xor U28026 (N_28026,N_27201,N_27208);
or U28027 (N_28027,N_27945,N_27491);
and U28028 (N_28028,N_27250,N_27195);
xnor U28029 (N_28029,N_27585,N_27843);
xnor U28030 (N_28030,N_27947,N_27802);
or U28031 (N_28031,N_27738,N_27443);
nand U28032 (N_28032,N_27865,N_27123);
nand U28033 (N_28033,N_27806,N_27353);
xor U28034 (N_28034,N_27080,N_27679);
and U28035 (N_28035,N_27010,N_27023);
xnor U28036 (N_28036,N_27984,N_27189);
nor U28037 (N_28037,N_27756,N_27277);
or U28038 (N_28038,N_27692,N_27700);
nor U28039 (N_28039,N_27054,N_27797);
or U28040 (N_28040,N_27689,N_27227);
nor U28041 (N_28041,N_27589,N_27507);
nor U28042 (N_28042,N_27008,N_27991);
nor U28043 (N_28043,N_27100,N_27621);
nand U28044 (N_28044,N_27117,N_27166);
and U28045 (N_28045,N_27757,N_27778);
xnor U28046 (N_28046,N_27955,N_27261);
or U28047 (N_28047,N_27766,N_27849);
nand U28048 (N_28048,N_27707,N_27193);
nor U28049 (N_28049,N_27462,N_27345);
and U28050 (N_28050,N_27058,N_27230);
or U28051 (N_28051,N_27887,N_27504);
and U28052 (N_28052,N_27118,N_27744);
or U28053 (N_28053,N_27436,N_27851);
and U28054 (N_28054,N_27015,N_27678);
nor U28055 (N_28055,N_27724,N_27056);
or U28056 (N_28056,N_27251,N_27470);
and U28057 (N_28057,N_27433,N_27200);
or U28058 (N_28058,N_27855,N_27021);
nor U28059 (N_28059,N_27347,N_27047);
nand U28060 (N_28060,N_27911,N_27194);
xor U28061 (N_28061,N_27524,N_27558);
xor U28062 (N_28062,N_27860,N_27636);
nor U28063 (N_28063,N_27934,N_27405);
nand U28064 (N_28064,N_27870,N_27378);
xnor U28065 (N_28065,N_27141,N_27545);
nand U28066 (N_28066,N_27046,N_27076);
and U28067 (N_28067,N_27281,N_27027);
nand U28068 (N_28068,N_27654,N_27174);
and U28069 (N_28069,N_27420,N_27803);
and U28070 (N_28070,N_27771,N_27265);
or U28071 (N_28071,N_27686,N_27539);
xnor U28072 (N_28072,N_27341,N_27428);
nor U28073 (N_28073,N_27472,N_27617);
or U28074 (N_28074,N_27940,N_27455);
xor U28075 (N_28075,N_27665,N_27684);
and U28076 (N_28076,N_27244,N_27492);
xor U28077 (N_28077,N_27161,N_27995);
nand U28078 (N_28078,N_27041,N_27872);
nor U28079 (N_28079,N_27561,N_27963);
nand U28080 (N_28080,N_27368,N_27165);
or U28081 (N_28081,N_27482,N_27550);
nand U28082 (N_28082,N_27135,N_27309);
or U28083 (N_28083,N_27681,N_27078);
nand U28084 (N_28084,N_27541,N_27217);
and U28085 (N_28085,N_27187,N_27535);
nand U28086 (N_28086,N_27526,N_27685);
nand U28087 (N_28087,N_27645,N_27993);
or U28088 (N_28088,N_27418,N_27599);
xor U28089 (N_28089,N_27424,N_27314);
nand U28090 (N_28090,N_27241,N_27846);
or U28091 (N_28091,N_27119,N_27716);
or U28092 (N_28092,N_27228,N_27596);
nor U28093 (N_28093,N_27381,N_27626);
nor U28094 (N_28094,N_27761,N_27310);
and U28095 (N_28095,N_27348,N_27708);
and U28096 (N_28096,N_27094,N_27976);
nor U28097 (N_28097,N_27680,N_27185);
or U28098 (N_28098,N_27276,N_27885);
nand U28099 (N_28099,N_27956,N_27594);
xnor U28100 (N_28100,N_27703,N_27129);
nand U28101 (N_28101,N_27385,N_27019);
nor U28102 (N_28102,N_27569,N_27350);
nand U28103 (N_28103,N_27907,N_27831);
or U28104 (N_28104,N_27549,N_27718);
nand U28105 (N_28105,N_27877,N_27474);
nor U28106 (N_28106,N_27715,N_27790);
nand U28107 (N_28107,N_27900,N_27985);
nor U28108 (N_28108,N_27987,N_27393);
nor U28109 (N_28109,N_27970,N_27879);
xnor U28110 (N_28110,N_27301,N_27223);
and U28111 (N_28111,N_27231,N_27952);
and U28112 (N_28112,N_27236,N_27827);
xor U28113 (N_28113,N_27868,N_27465);
nor U28114 (N_28114,N_27858,N_27034);
or U28115 (N_28115,N_27302,N_27112);
and U28116 (N_28116,N_27212,N_27631);
xnor U28117 (N_28117,N_27180,N_27701);
or U28118 (N_28118,N_27475,N_27562);
and U28119 (N_28119,N_27752,N_27528);
or U28120 (N_28120,N_27552,N_27782);
nor U28121 (N_28121,N_27640,N_27974);
nor U28122 (N_28122,N_27902,N_27237);
and U28123 (N_28123,N_27601,N_27068);
nand U28124 (N_28124,N_27374,N_27113);
xor U28125 (N_28125,N_27464,N_27499);
or U28126 (N_28126,N_27255,N_27800);
or U28127 (N_28127,N_27088,N_27727);
nand U28128 (N_28128,N_27845,N_27136);
or U28129 (N_28129,N_27346,N_27614);
xor U28130 (N_28130,N_27677,N_27178);
nand U28131 (N_28131,N_27229,N_27017);
nand U28132 (N_28132,N_27226,N_27839);
xnor U28133 (N_28133,N_27825,N_27456);
and U28134 (N_28134,N_27090,N_27401);
xor U28135 (N_28135,N_27085,N_27089);
nor U28136 (N_28136,N_27399,N_27918);
or U28137 (N_28137,N_27422,N_27026);
nand U28138 (N_28138,N_27408,N_27184);
and U28139 (N_28139,N_27303,N_27780);
nand U28140 (N_28140,N_27737,N_27337);
or U28141 (N_28141,N_27505,N_27763);
and U28142 (N_28142,N_27548,N_27938);
and U28143 (N_28143,N_27613,N_27814);
nor U28144 (N_28144,N_27833,N_27662);
nor U28145 (N_28145,N_27300,N_27619);
xor U28146 (N_28146,N_27876,N_27240);
and U28147 (N_28147,N_27116,N_27308);
nor U28148 (N_28148,N_27795,N_27823);
and U28149 (N_28149,N_27743,N_27275);
nand U28150 (N_28150,N_27830,N_27765);
or U28151 (N_28151,N_27576,N_27914);
nand U28152 (N_28152,N_27247,N_27642);
nor U28153 (N_28153,N_27990,N_27086);
xor U28154 (N_28154,N_27572,N_27392);
or U28155 (N_28155,N_27367,N_27177);
xor U28156 (N_28156,N_27656,N_27785);
or U28157 (N_28157,N_27294,N_27442);
nor U28158 (N_28158,N_27547,N_27018);
or U28159 (N_28159,N_27371,N_27182);
and U28160 (N_28160,N_27480,N_27339);
xor U28161 (N_28161,N_27647,N_27867);
nand U28162 (N_28162,N_27485,N_27687);
nor U28163 (N_28163,N_27953,N_27931);
nand U28164 (N_28164,N_27039,N_27676);
and U28165 (N_28165,N_27511,N_27733);
or U28166 (N_28166,N_27978,N_27832);
nand U28167 (N_28167,N_27893,N_27835);
nor U28168 (N_28168,N_27643,N_27622);
xnor U28169 (N_28169,N_27211,N_27001);
xor U28170 (N_28170,N_27603,N_27891);
xor U28171 (N_28171,N_27804,N_27777);
nor U28172 (N_28172,N_27179,N_27035);
and U28173 (N_28173,N_27454,N_27736);
or U28174 (N_28174,N_27000,N_27981);
nand U28175 (N_28175,N_27221,N_27755);
nand U28176 (N_28176,N_27527,N_27633);
or U28177 (N_28177,N_27591,N_27259);
xor U28178 (N_28178,N_27509,N_27888);
nand U28179 (N_28179,N_27579,N_27741);
or U28180 (N_28180,N_27126,N_27077);
or U28181 (N_28181,N_27127,N_27897);
nor U28182 (N_28182,N_27714,N_27999);
or U28183 (N_28183,N_27372,N_27045);
and U28184 (N_28184,N_27789,N_27463);
nand U28185 (N_28185,N_27245,N_27163);
and U28186 (N_28186,N_27406,N_27798);
nand U28187 (N_28187,N_27224,N_27666);
and U28188 (N_28188,N_27147,N_27412);
nand U28189 (N_28189,N_27239,N_27951);
xor U28190 (N_28190,N_27105,N_27404);
and U28191 (N_28191,N_27458,N_27554);
or U28192 (N_28192,N_27817,N_27739);
xor U28193 (N_28193,N_27397,N_27775);
and U28194 (N_28194,N_27523,N_27989);
and U28195 (N_28195,N_27567,N_27175);
or U28196 (N_28196,N_27824,N_27975);
nand U28197 (N_28197,N_27198,N_27444);
nand U28198 (N_28198,N_27972,N_27711);
or U28199 (N_28199,N_27819,N_27531);
xnor U28200 (N_28200,N_27220,N_27501);
nor U28201 (N_28201,N_27906,N_27516);
or U28202 (N_28202,N_27384,N_27323);
and U28203 (N_28203,N_27287,N_27847);
and U28204 (N_28204,N_27690,N_27369);
nand U28205 (N_28205,N_27751,N_27828);
or U28206 (N_28206,N_27587,N_27653);
xnor U28207 (N_28207,N_27884,N_27913);
xor U28208 (N_28208,N_27584,N_27486);
and U28209 (N_28209,N_27453,N_27959);
and U28210 (N_28210,N_27878,N_27279);
nor U28211 (N_28211,N_27604,N_27417);
nand U28212 (N_28212,N_27783,N_27097);
nor U28213 (N_28213,N_27293,N_27917);
xor U28214 (N_28214,N_27764,N_27387);
nand U28215 (N_28215,N_27364,N_27439);
xor U28216 (N_28216,N_27115,N_27402);
and U28217 (N_28217,N_27489,N_27908);
xor U28218 (N_28218,N_27807,N_27950);
nor U28219 (N_28219,N_27563,N_27361);
or U28220 (N_28220,N_27683,N_27837);
nand U28221 (N_28221,N_27894,N_27156);
xor U28222 (N_28222,N_27256,N_27383);
or U28223 (N_28223,N_27553,N_27682);
or U28224 (N_28224,N_27267,N_27377);
nand U28225 (N_28225,N_27375,N_27466);
nand U28226 (N_28226,N_27618,N_27467);
nor U28227 (N_28227,N_27538,N_27784);
or U28228 (N_28228,N_27358,N_27121);
and U28229 (N_28229,N_27895,N_27205);
xor U28230 (N_28230,N_27996,N_27400);
or U28231 (N_28231,N_27122,N_27600);
and U28232 (N_28232,N_27431,N_27081);
or U28233 (N_28233,N_27328,N_27304);
or U28234 (N_28234,N_27274,N_27434);
nor U28235 (N_28235,N_27336,N_27712);
xnor U28236 (N_28236,N_27874,N_27927);
xor U28237 (N_28237,N_27268,N_27044);
and U28238 (N_28238,N_27694,N_27490);
xnor U28239 (N_28239,N_27871,N_27215);
or U28240 (N_28240,N_27886,N_27889);
nor U28241 (N_28241,N_27355,N_27427);
nand U28242 (N_28242,N_27448,N_27731);
and U28243 (N_28243,N_27264,N_27786);
and U28244 (N_28244,N_27188,N_27219);
or U28245 (N_28245,N_27298,N_27183);
xor U28246 (N_28246,N_27471,N_27052);
and U28247 (N_28247,N_27297,N_27810);
and U28248 (N_28248,N_27049,N_27106);
xor U28249 (N_28249,N_27065,N_27093);
nand U28250 (N_28250,N_27331,N_27740);
xnor U28251 (N_28251,N_27840,N_27329);
or U28252 (N_28252,N_27536,N_27948);
xor U28253 (N_28253,N_27382,N_27270);
xor U28254 (N_28254,N_27403,N_27079);
nand U28255 (N_28255,N_27349,N_27838);
xnor U28256 (N_28256,N_27937,N_27648);
nand U28257 (N_28257,N_27338,N_27057);
or U28258 (N_28258,N_27064,N_27091);
nor U28259 (N_28259,N_27222,N_27238);
nand U28260 (N_28260,N_27941,N_27932);
and U28261 (N_28261,N_27266,N_27770);
xnor U28262 (N_28262,N_27675,N_27853);
and U28263 (N_28263,N_27627,N_27670);
and U28264 (N_28264,N_27646,N_27657);
or U28265 (N_28265,N_27609,N_27059);
xnor U28266 (N_28266,N_27199,N_27450);
nor U28267 (N_28267,N_27131,N_27153);
nor U28268 (N_28268,N_27791,N_27011);
or U28269 (N_28269,N_27801,N_27330);
or U28270 (N_28270,N_27650,N_27357);
nand U28271 (N_28271,N_27468,N_27447);
or U28272 (N_28272,N_27446,N_27432);
and U28273 (N_28273,N_27016,N_27578);
and U28274 (N_28274,N_27242,N_27143);
or U28275 (N_28275,N_27588,N_27216);
nand U28276 (N_28276,N_27570,N_27958);
or U28277 (N_28277,N_27598,N_27597);
nor U28278 (N_28278,N_27313,N_27248);
nand U28279 (N_28279,N_27842,N_27409);
nand U28280 (N_28280,N_27568,N_27171);
nand U28281 (N_28281,N_27391,N_27898);
and U28282 (N_28282,N_27667,N_27542);
nand U28283 (N_28283,N_27658,N_27863);
or U28284 (N_28284,N_27344,N_27299);
and U28285 (N_28285,N_27788,N_27998);
nor U28286 (N_28286,N_27191,N_27904);
and U28287 (N_28287,N_27546,N_27518);
and U28288 (N_28288,N_27413,N_27559);
nor U28289 (N_28289,N_27580,N_27673);
or U28290 (N_28290,N_27957,N_27534);
nand U28291 (N_28291,N_27396,N_27721);
nor U28292 (N_28292,N_27278,N_27768);
and U28293 (N_28293,N_27243,N_27343);
xor U28294 (N_28294,N_27273,N_27162);
xnor U28295 (N_28295,N_27457,N_27048);
and U28296 (N_28296,N_27730,N_27942);
xnor U28297 (N_28297,N_27004,N_27484);
and U28298 (N_28298,N_27669,N_27813);
and U28299 (N_28299,N_27632,N_27290);
nor U28300 (N_28300,N_27875,N_27258);
or U28301 (N_28301,N_27398,N_27774);
nor U28302 (N_28302,N_27386,N_27373);
xor U28303 (N_28303,N_27082,N_27103);
nand U28304 (N_28304,N_27960,N_27710);
and U28305 (N_28305,N_27944,N_27109);
nand U28306 (N_28306,N_27286,N_27172);
and U28307 (N_28307,N_27038,N_27232);
xnor U28308 (N_28308,N_27962,N_27148);
and U28309 (N_28309,N_27025,N_27029);
xnor U28310 (N_28310,N_27850,N_27728);
nor U28311 (N_28311,N_27968,N_27495);
nor U28312 (N_28312,N_27426,N_27512);
and U28313 (N_28313,N_27796,N_27181);
xor U28314 (N_28314,N_27214,N_27794);
or U28315 (N_28315,N_27316,N_27007);
or U28316 (N_28316,N_27410,N_27478);
xnor U28317 (N_28317,N_27916,N_27028);
xor U28318 (N_28318,N_27022,N_27869);
or U28319 (N_28319,N_27042,N_27133);
and U28320 (N_28320,N_27691,N_27779);
or U28321 (N_28321,N_27571,N_27149);
nand U28322 (N_28322,N_27359,N_27529);
and U28323 (N_28323,N_27315,N_27360);
and U28324 (N_28324,N_27164,N_27652);
xnor U28325 (N_28325,N_27257,N_27928);
xnor U28326 (N_28326,N_27722,N_27726);
nand U28327 (N_28327,N_27407,N_27812);
and U28328 (N_28328,N_27625,N_27150);
nand U28329 (N_28329,N_27415,N_27051);
and U28330 (N_28330,N_27753,N_27695);
nor U28331 (N_28331,N_27271,N_27370);
xnor U28332 (N_28332,N_27066,N_27429);
xnor U28333 (N_28333,N_27324,N_27688);
nand U28334 (N_28334,N_27834,N_27729);
nor U28335 (N_28335,N_27732,N_27983);
nand U28336 (N_28336,N_27734,N_27020);
xnor U28337 (N_28337,N_27923,N_27033);
and U28338 (N_28338,N_27356,N_27252);
and U28339 (N_28339,N_27235,N_27709);
nor U28340 (N_28340,N_27943,N_27969);
nor U28341 (N_28341,N_27595,N_27905);
nor U28342 (N_28342,N_27145,N_27748);
nand U28343 (N_28343,N_27861,N_27074);
nand U28344 (N_28344,N_27269,N_27698);
nor U28345 (N_28345,N_27713,N_27295);
xor U28346 (N_28346,N_27479,N_27787);
and U28347 (N_28347,N_27130,N_27036);
nand U28348 (N_28348,N_27880,N_27635);
nor U28349 (N_28349,N_27760,N_27890);
nor U28350 (N_28350,N_27859,N_27986);
nand U28351 (N_28351,N_27793,N_27146);
xnor U28352 (N_28352,N_27532,N_27071);
and U28353 (N_28353,N_27735,N_27994);
nor U28354 (N_28354,N_27624,N_27611);
and U28355 (N_28355,N_27909,N_27352);
or U28356 (N_28356,N_27169,N_27674);
nand U28357 (N_28357,N_27967,N_27892);
nor U28358 (N_28358,N_27754,N_27725);
xnor U28359 (N_28359,N_27206,N_27530);
nand U28360 (N_28360,N_27717,N_27210);
or U28361 (N_28361,N_27586,N_27128);
and U28362 (N_28362,N_27696,N_27769);
nor U28363 (N_28363,N_27560,N_27857);
or U28364 (N_28364,N_27749,N_27070);
nand U28365 (N_28365,N_27848,N_27140);
nor U28366 (N_28366,N_27852,N_27213);
or U28367 (N_28367,N_27098,N_27351);
and U28368 (N_28368,N_27414,N_27977);
xor U28369 (N_28369,N_27321,N_27487);
nand U28370 (N_28370,N_27672,N_27961);
nand U28371 (N_28371,N_27389,N_27190);
nor U28372 (N_28372,N_27151,N_27610);
or U28373 (N_28373,N_27005,N_27288);
nor U28374 (N_28374,N_27154,N_27919);
or U28375 (N_28375,N_27903,N_27395);
nand U28376 (N_28376,N_27540,N_27805);
nand U28377 (N_28377,N_27110,N_27639);
nand U28378 (N_28378,N_27582,N_27272);
or U28379 (N_28379,N_27544,N_27296);
nor U28380 (N_28380,N_27421,N_27697);
xor U28381 (N_28381,N_27254,N_27234);
and U28382 (N_28382,N_27380,N_27196);
nand U28383 (N_28383,N_27158,N_27508);
nor U28384 (N_28384,N_27921,N_27925);
or U28385 (N_28385,N_27844,N_27750);
and U28386 (N_28386,N_27073,N_27481);
and U28387 (N_28387,N_27664,N_27808);
or U28388 (N_28388,N_27451,N_27575);
nor U28389 (N_28389,N_27144,N_27411);
nor U28390 (N_28390,N_27390,N_27280);
nor U28391 (N_28391,N_27494,N_27638);
nor U28392 (N_28392,N_27543,N_27930);
and U28393 (N_28393,N_27445,N_27013);
nand U28394 (N_28394,N_27818,N_27767);
and U28395 (N_28395,N_27517,N_27882);
and U28396 (N_28396,N_27602,N_27461);
and U28397 (N_28397,N_27062,N_27920);
nor U28398 (N_28398,N_27641,N_27155);
nor U28399 (N_28399,N_27173,N_27661);
nand U28400 (N_28400,N_27792,N_27327);
or U28401 (N_28401,N_27965,N_27759);
nor U28402 (N_28402,N_27705,N_27002);
nor U28403 (N_28403,N_27137,N_27291);
and U28404 (N_28404,N_27745,N_27773);
or U28405 (N_28405,N_27120,N_27829);
xor U28406 (N_28406,N_27933,N_27037);
xor U28407 (N_28407,N_27111,N_27922);
and U28408 (N_28408,N_27325,N_27520);
or U28409 (N_28409,N_27043,N_27132);
xor U28410 (N_28410,N_27282,N_27809);
and U28411 (N_28411,N_27644,N_27284);
nand U28412 (N_28412,N_27108,N_27781);
and U28413 (N_28413,N_27092,N_27170);
nand U28414 (N_28414,N_27873,N_27425);
nor U28415 (N_28415,N_27620,N_27896);
xnor U28416 (N_28416,N_27365,N_27772);
and U28417 (N_28417,N_27612,N_27075);
nand U28418 (N_28418,N_27363,N_27102);
xor U28419 (N_28419,N_27939,N_27583);
nand U28420 (N_28420,N_27225,N_27719);
xnor U28421 (N_28421,N_27114,N_27311);
xnor U28422 (N_28422,N_27929,N_27469);
and U28423 (N_28423,N_27519,N_27263);
nand U28424 (N_28424,N_27979,N_27936);
nor U28425 (N_28425,N_27565,N_27285);
xnor U28426 (N_28426,N_27388,N_27521);
or U28427 (N_28427,N_27483,N_27006);
nor U28428 (N_28428,N_27924,N_27593);
and U28429 (N_28429,N_27317,N_27440);
and U28430 (N_28430,N_27012,N_27176);
nor U28431 (N_28431,N_27502,N_27634);
nor U28432 (N_28432,N_27514,N_27854);
nand U28433 (N_28433,N_27342,N_27306);
or U28434 (N_28434,N_27305,N_27555);
and U28435 (N_28435,N_27720,N_27966);
nor U28436 (N_28436,N_27926,N_27477);
and U28437 (N_28437,N_27233,N_27340);
or U28438 (N_28438,N_27096,N_27910);
or U28439 (N_28439,N_27607,N_27441);
and U28440 (N_28440,N_27437,N_27551);
or U28441 (N_28441,N_27083,N_27564);
and U28442 (N_28442,N_27856,N_27581);
or U28443 (N_28443,N_27435,N_27982);
nor U28444 (N_28444,N_27496,N_27826);
nand U28445 (N_28445,N_27031,N_27072);
and U28446 (N_28446,N_27515,N_27099);
nand U28447 (N_28447,N_27160,N_27706);
nand U28448 (N_28448,N_27124,N_27125);
xnor U28449 (N_28449,N_27742,N_27104);
nor U28450 (N_28450,N_27326,N_27592);
nor U28451 (N_28451,N_27138,N_27040);
or U28452 (N_28452,N_27493,N_27935);
nand U28453 (N_28453,N_27335,N_27510);
xnor U28454 (N_28454,N_27032,N_27616);
xor U28455 (N_28455,N_27556,N_27973);
and U28456 (N_28456,N_27946,N_27262);
and U28457 (N_28457,N_27615,N_27577);
and U28458 (N_28458,N_27473,N_27061);
nand U28459 (N_28459,N_27899,N_27319);
xor U28460 (N_28460,N_27009,N_27246);
nor U28461 (N_28461,N_27980,N_27628);
xnor U28462 (N_28462,N_27334,N_27167);
or U28463 (N_28463,N_27283,N_27660);
or U28464 (N_28464,N_27912,N_27333);
and U28465 (N_28465,N_27142,N_27366);
or U28466 (N_28466,N_27590,N_27758);
nor U28467 (N_28467,N_27704,N_27312);
xor U28468 (N_28468,N_27971,N_27815);
or U28469 (N_28469,N_27003,N_27702);
nand U28470 (N_28470,N_27503,N_27836);
or U28471 (N_28471,N_27566,N_27500);
nand U28472 (N_28472,N_27460,N_27438);
xnor U28473 (N_28473,N_27537,N_27816);
nand U28474 (N_28474,N_27746,N_27307);
or U28475 (N_28475,N_27533,N_27522);
and U28476 (N_28476,N_27498,N_27655);
nor U28477 (N_28477,N_27430,N_27476);
and U28478 (N_28478,N_27055,N_27218);
nand U28479 (N_28479,N_27693,N_27260);
and U28480 (N_28480,N_27159,N_27292);
or U28481 (N_28481,N_27864,N_27637);
and U28482 (N_28482,N_27997,N_27168);
xor U28483 (N_28483,N_27084,N_27992);
nand U28484 (N_28484,N_27318,N_27747);
or U28485 (N_28485,N_27841,N_27107);
nand U28486 (N_28486,N_27087,N_27423);
nand U28487 (N_28487,N_27557,N_27506);
and U28488 (N_28488,N_27322,N_27574);
nand U28489 (N_28489,N_27050,N_27608);
nor U28490 (N_28490,N_27139,N_27497);
nor U28491 (N_28491,N_27663,N_27376);
nand U28492 (N_28492,N_27332,N_27915);
and U28493 (N_28493,N_27063,N_27209);
nor U28494 (N_28494,N_27101,N_27186);
xnor U28495 (N_28495,N_27192,N_27060);
and U28496 (N_28496,N_27014,N_27954);
nor U28497 (N_28497,N_27449,N_27197);
nor U28498 (N_28498,N_27249,N_27362);
xnor U28499 (N_28499,N_27416,N_27949);
nor U28500 (N_28500,N_27148,N_27039);
xor U28501 (N_28501,N_27152,N_27983);
nor U28502 (N_28502,N_27466,N_27239);
nand U28503 (N_28503,N_27443,N_27828);
xnor U28504 (N_28504,N_27885,N_27043);
and U28505 (N_28505,N_27476,N_27914);
or U28506 (N_28506,N_27474,N_27493);
xnor U28507 (N_28507,N_27028,N_27486);
xor U28508 (N_28508,N_27857,N_27739);
or U28509 (N_28509,N_27394,N_27717);
xnor U28510 (N_28510,N_27119,N_27250);
and U28511 (N_28511,N_27247,N_27918);
nand U28512 (N_28512,N_27937,N_27078);
or U28513 (N_28513,N_27373,N_27665);
and U28514 (N_28514,N_27757,N_27245);
and U28515 (N_28515,N_27870,N_27646);
xnor U28516 (N_28516,N_27227,N_27237);
or U28517 (N_28517,N_27192,N_27456);
nor U28518 (N_28518,N_27531,N_27855);
or U28519 (N_28519,N_27003,N_27135);
or U28520 (N_28520,N_27107,N_27914);
nor U28521 (N_28521,N_27073,N_27029);
nor U28522 (N_28522,N_27083,N_27920);
nand U28523 (N_28523,N_27353,N_27944);
nand U28524 (N_28524,N_27463,N_27601);
and U28525 (N_28525,N_27749,N_27023);
nor U28526 (N_28526,N_27363,N_27854);
and U28527 (N_28527,N_27265,N_27282);
nand U28528 (N_28528,N_27166,N_27263);
xor U28529 (N_28529,N_27095,N_27148);
nor U28530 (N_28530,N_27675,N_27547);
nand U28531 (N_28531,N_27832,N_27543);
or U28532 (N_28532,N_27946,N_27524);
and U28533 (N_28533,N_27543,N_27163);
or U28534 (N_28534,N_27717,N_27815);
xor U28535 (N_28535,N_27606,N_27138);
xor U28536 (N_28536,N_27673,N_27117);
nor U28537 (N_28537,N_27797,N_27135);
or U28538 (N_28538,N_27407,N_27144);
and U28539 (N_28539,N_27395,N_27941);
and U28540 (N_28540,N_27763,N_27136);
nor U28541 (N_28541,N_27024,N_27339);
or U28542 (N_28542,N_27317,N_27627);
nor U28543 (N_28543,N_27678,N_27696);
xnor U28544 (N_28544,N_27086,N_27709);
and U28545 (N_28545,N_27001,N_27828);
and U28546 (N_28546,N_27020,N_27810);
nor U28547 (N_28547,N_27597,N_27939);
nand U28548 (N_28548,N_27177,N_27461);
xnor U28549 (N_28549,N_27070,N_27454);
nand U28550 (N_28550,N_27132,N_27514);
xnor U28551 (N_28551,N_27354,N_27830);
or U28552 (N_28552,N_27331,N_27075);
xor U28553 (N_28553,N_27296,N_27136);
nor U28554 (N_28554,N_27148,N_27697);
xnor U28555 (N_28555,N_27091,N_27243);
nand U28556 (N_28556,N_27052,N_27224);
nor U28557 (N_28557,N_27571,N_27909);
nand U28558 (N_28558,N_27205,N_27169);
or U28559 (N_28559,N_27794,N_27980);
and U28560 (N_28560,N_27646,N_27228);
or U28561 (N_28561,N_27315,N_27215);
or U28562 (N_28562,N_27565,N_27596);
nand U28563 (N_28563,N_27888,N_27281);
nor U28564 (N_28564,N_27314,N_27845);
nor U28565 (N_28565,N_27012,N_27760);
and U28566 (N_28566,N_27784,N_27640);
and U28567 (N_28567,N_27052,N_27685);
nor U28568 (N_28568,N_27183,N_27968);
nor U28569 (N_28569,N_27258,N_27829);
xnor U28570 (N_28570,N_27728,N_27195);
nand U28571 (N_28571,N_27540,N_27915);
nand U28572 (N_28572,N_27775,N_27804);
xor U28573 (N_28573,N_27699,N_27451);
and U28574 (N_28574,N_27688,N_27831);
nand U28575 (N_28575,N_27972,N_27849);
xnor U28576 (N_28576,N_27034,N_27097);
xor U28577 (N_28577,N_27781,N_27176);
and U28578 (N_28578,N_27382,N_27429);
or U28579 (N_28579,N_27185,N_27119);
nand U28580 (N_28580,N_27644,N_27968);
nor U28581 (N_28581,N_27569,N_27942);
or U28582 (N_28582,N_27190,N_27315);
or U28583 (N_28583,N_27625,N_27819);
nor U28584 (N_28584,N_27855,N_27442);
and U28585 (N_28585,N_27164,N_27192);
nand U28586 (N_28586,N_27451,N_27168);
nor U28587 (N_28587,N_27090,N_27381);
nor U28588 (N_28588,N_27919,N_27732);
and U28589 (N_28589,N_27464,N_27171);
nor U28590 (N_28590,N_27762,N_27785);
nand U28591 (N_28591,N_27167,N_27241);
xor U28592 (N_28592,N_27237,N_27331);
nor U28593 (N_28593,N_27601,N_27492);
and U28594 (N_28594,N_27989,N_27057);
and U28595 (N_28595,N_27622,N_27773);
and U28596 (N_28596,N_27595,N_27377);
or U28597 (N_28597,N_27760,N_27577);
and U28598 (N_28598,N_27740,N_27221);
nor U28599 (N_28599,N_27943,N_27970);
and U28600 (N_28600,N_27680,N_27950);
nor U28601 (N_28601,N_27937,N_27957);
xor U28602 (N_28602,N_27814,N_27747);
xor U28603 (N_28603,N_27167,N_27501);
nor U28604 (N_28604,N_27581,N_27981);
nor U28605 (N_28605,N_27488,N_27927);
and U28606 (N_28606,N_27872,N_27328);
or U28607 (N_28607,N_27599,N_27806);
nor U28608 (N_28608,N_27915,N_27495);
or U28609 (N_28609,N_27091,N_27036);
and U28610 (N_28610,N_27991,N_27876);
or U28611 (N_28611,N_27398,N_27134);
xor U28612 (N_28612,N_27392,N_27272);
nor U28613 (N_28613,N_27312,N_27363);
or U28614 (N_28614,N_27635,N_27567);
and U28615 (N_28615,N_27312,N_27246);
nand U28616 (N_28616,N_27120,N_27964);
and U28617 (N_28617,N_27995,N_27901);
xnor U28618 (N_28618,N_27281,N_27126);
nand U28619 (N_28619,N_27829,N_27621);
xnor U28620 (N_28620,N_27939,N_27051);
or U28621 (N_28621,N_27427,N_27089);
nand U28622 (N_28622,N_27516,N_27315);
nand U28623 (N_28623,N_27041,N_27575);
and U28624 (N_28624,N_27257,N_27091);
nand U28625 (N_28625,N_27108,N_27790);
nor U28626 (N_28626,N_27021,N_27322);
nor U28627 (N_28627,N_27997,N_27438);
xor U28628 (N_28628,N_27013,N_27923);
and U28629 (N_28629,N_27328,N_27543);
xor U28630 (N_28630,N_27520,N_27497);
nor U28631 (N_28631,N_27026,N_27508);
nand U28632 (N_28632,N_27911,N_27311);
xnor U28633 (N_28633,N_27580,N_27507);
nand U28634 (N_28634,N_27507,N_27287);
or U28635 (N_28635,N_27494,N_27848);
nor U28636 (N_28636,N_27414,N_27212);
xnor U28637 (N_28637,N_27780,N_27448);
nand U28638 (N_28638,N_27971,N_27337);
xnor U28639 (N_28639,N_27957,N_27098);
xor U28640 (N_28640,N_27037,N_27959);
or U28641 (N_28641,N_27741,N_27002);
and U28642 (N_28642,N_27481,N_27952);
and U28643 (N_28643,N_27719,N_27985);
xor U28644 (N_28644,N_27872,N_27977);
nand U28645 (N_28645,N_27986,N_27171);
nand U28646 (N_28646,N_27188,N_27926);
and U28647 (N_28647,N_27396,N_27057);
or U28648 (N_28648,N_27661,N_27646);
xnor U28649 (N_28649,N_27745,N_27098);
and U28650 (N_28650,N_27808,N_27564);
nor U28651 (N_28651,N_27238,N_27508);
nor U28652 (N_28652,N_27717,N_27502);
nor U28653 (N_28653,N_27463,N_27556);
or U28654 (N_28654,N_27396,N_27316);
or U28655 (N_28655,N_27400,N_27257);
xor U28656 (N_28656,N_27466,N_27402);
nand U28657 (N_28657,N_27046,N_27054);
and U28658 (N_28658,N_27234,N_27135);
or U28659 (N_28659,N_27861,N_27041);
xor U28660 (N_28660,N_27213,N_27621);
xnor U28661 (N_28661,N_27567,N_27524);
xor U28662 (N_28662,N_27520,N_27635);
nand U28663 (N_28663,N_27418,N_27200);
or U28664 (N_28664,N_27913,N_27074);
xor U28665 (N_28665,N_27534,N_27535);
or U28666 (N_28666,N_27832,N_27130);
nand U28667 (N_28667,N_27753,N_27629);
and U28668 (N_28668,N_27014,N_27639);
nand U28669 (N_28669,N_27972,N_27449);
and U28670 (N_28670,N_27726,N_27369);
xnor U28671 (N_28671,N_27531,N_27089);
and U28672 (N_28672,N_27356,N_27395);
nand U28673 (N_28673,N_27294,N_27125);
nand U28674 (N_28674,N_27671,N_27095);
or U28675 (N_28675,N_27040,N_27069);
xnor U28676 (N_28676,N_27577,N_27738);
xor U28677 (N_28677,N_27780,N_27318);
or U28678 (N_28678,N_27726,N_27623);
or U28679 (N_28679,N_27171,N_27733);
xor U28680 (N_28680,N_27898,N_27559);
nor U28681 (N_28681,N_27968,N_27732);
xor U28682 (N_28682,N_27830,N_27529);
or U28683 (N_28683,N_27576,N_27438);
nor U28684 (N_28684,N_27233,N_27420);
nor U28685 (N_28685,N_27545,N_27867);
xnor U28686 (N_28686,N_27047,N_27776);
or U28687 (N_28687,N_27896,N_27482);
or U28688 (N_28688,N_27044,N_27496);
nor U28689 (N_28689,N_27424,N_27931);
or U28690 (N_28690,N_27200,N_27821);
nor U28691 (N_28691,N_27415,N_27003);
and U28692 (N_28692,N_27724,N_27087);
nand U28693 (N_28693,N_27162,N_27838);
xnor U28694 (N_28694,N_27783,N_27818);
or U28695 (N_28695,N_27637,N_27920);
or U28696 (N_28696,N_27811,N_27953);
or U28697 (N_28697,N_27475,N_27066);
nand U28698 (N_28698,N_27183,N_27599);
or U28699 (N_28699,N_27773,N_27528);
nand U28700 (N_28700,N_27022,N_27858);
and U28701 (N_28701,N_27426,N_27341);
nor U28702 (N_28702,N_27061,N_27717);
xor U28703 (N_28703,N_27415,N_27323);
or U28704 (N_28704,N_27111,N_27273);
or U28705 (N_28705,N_27838,N_27809);
xor U28706 (N_28706,N_27808,N_27370);
or U28707 (N_28707,N_27666,N_27781);
xnor U28708 (N_28708,N_27729,N_27004);
nand U28709 (N_28709,N_27564,N_27659);
nand U28710 (N_28710,N_27545,N_27916);
and U28711 (N_28711,N_27159,N_27107);
nor U28712 (N_28712,N_27350,N_27015);
nand U28713 (N_28713,N_27322,N_27588);
xor U28714 (N_28714,N_27654,N_27961);
and U28715 (N_28715,N_27088,N_27782);
or U28716 (N_28716,N_27450,N_27971);
and U28717 (N_28717,N_27768,N_27513);
and U28718 (N_28718,N_27079,N_27671);
or U28719 (N_28719,N_27133,N_27624);
xor U28720 (N_28720,N_27858,N_27213);
or U28721 (N_28721,N_27410,N_27025);
xnor U28722 (N_28722,N_27386,N_27886);
nand U28723 (N_28723,N_27515,N_27891);
or U28724 (N_28724,N_27478,N_27466);
nand U28725 (N_28725,N_27852,N_27159);
and U28726 (N_28726,N_27658,N_27706);
and U28727 (N_28727,N_27198,N_27169);
xor U28728 (N_28728,N_27698,N_27197);
or U28729 (N_28729,N_27364,N_27310);
nor U28730 (N_28730,N_27595,N_27676);
nand U28731 (N_28731,N_27249,N_27301);
xor U28732 (N_28732,N_27704,N_27622);
and U28733 (N_28733,N_27137,N_27456);
or U28734 (N_28734,N_27101,N_27555);
nor U28735 (N_28735,N_27078,N_27102);
xor U28736 (N_28736,N_27220,N_27337);
and U28737 (N_28737,N_27860,N_27237);
or U28738 (N_28738,N_27179,N_27765);
nand U28739 (N_28739,N_27352,N_27106);
nand U28740 (N_28740,N_27614,N_27046);
nand U28741 (N_28741,N_27389,N_27536);
or U28742 (N_28742,N_27189,N_27723);
xnor U28743 (N_28743,N_27505,N_27834);
nor U28744 (N_28744,N_27262,N_27117);
nor U28745 (N_28745,N_27152,N_27009);
xnor U28746 (N_28746,N_27027,N_27394);
nand U28747 (N_28747,N_27594,N_27319);
or U28748 (N_28748,N_27296,N_27736);
nand U28749 (N_28749,N_27561,N_27321);
xnor U28750 (N_28750,N_27693,N_27118);
xor U28751 (N_28751,N_27480,N_27590);
xnor U28752 (N_28752,N_27031,N_27218);
and U28753 (N_28753,N_27355,N_27512);
and U28754 (N_28754,N_27498,N_27643);
nand U28755 (N_28755,N_27799,N_27284);
xor U28756 (N_28756,N_27529,N_27901);
and U28757 (N_28757,N_27422,N_27727);
nand U28758 (N_28758,N_27053,N_27274);
xnor U28759 (N_28759,N_27479,N_27594);
or U28760 (N_28760,N_27620,N_27062);
and U28761 (N_28761,N_27325,N_27664);
xor U28762 (N_28762,N_27862,N_27737);
nand U28763 (N_28763,N_27014,N_27114);
and U28764 (N_28764,N_27767,N_27334);
and U28765 (N_28765,N_27968,N_27355);
and U28766 (N_28766,N_27118,N_27723);
nand U28767 (N_28767,N_27592,N_27516);
and U28768 (N_28768,N_27886,N_27491);
nor U28769 (N_28769,N_27875,N_27375);
nand U28770 (N_28770,N_27242,N_27190);
and U28771 (N_28771,N_27094,N_27846);
and U28772 (N_28772,N_27808,N_27605);
and U28773 (N_28773,N_27831,N_27336);
or U28774 (N_28774,N_27097,N_27954);
nand U28775 (N_28775,N_27113,N_27182);
or U28776 (N_28776,N_27056,N_27829);
xnor U28777 (N_28777,N_27386,N_27875);
nor U28778 (N_28778,N_27350,N_27731);
or U28779 (N_28779,N_27173,N_27171);
xor U28780 (N_28780,N_27724,N_27216);
and U28781 (N_28781,N_27754,N_27282);
nand U28782 (N_28782,N_27927,N_27897);
xor U28783 (N_28783,N_27998,N_27284);
nor U28784 (N_28784,N_27002,N_27389);
nor U28785 (N_28785,N_27738,N_27150);
nor U28786 (N_28786,N_27533,N_27792);
nor U28787 (N_28787,N_27276,N_27147);
nor U28788 (N_28788,N_27659,N_27371);
nand U28789 (N_28789,N_27846,N_27975);
nor U28790 (N_28790,N_27297,N_27558);
or U28791 (N_28791,N_27505,N_27617);
and U28792 (N_28792,N_27831,N_27990);
xor U28793 (N_28793,N_27969,N_27654);
and U28794 (N_28794,N_27988,N_27186);
or U28795 (N_28795,N_27378,N_27801);
or U28796 (N_28796,N_27259,N_27310);
nand U28797 (N_28797,N_27664,N_27190);
nand U28798 (N_28798,N_27125,N_27856);
nand U28799 (N_28799,N_27146,N_27081);
or U28800 (N_28800,N_27537,N_27336);
nand U28801 (N_28801,N_27351,N_27533);
and U28802 (N_28802,N_27074,N_27352);
nor U28803 (N_28803,N_27423,N_27888);
xor U28804 (N_28804,N_27127,N_27738);
nor U28805 (N_28805,N_27610,N_27527);
nand U28806 (N_28806,N_27855,N_27478);
and U28807 (N_28807,N_27762,N_27886);
or U28808 (N_28808,N_27926,N_27048);
or U28809 (N_28809,N_27274,N_27017);
xnor U28810 (N_28810,N_27162,N_27463);
nand U28811 (N_28811,N_27435,N_27319);
and U28812 (N_28812,N_27477,N_27675);
and U28813 (N_28813,N_27700,N_27629);
and U28814 (N_28814,N_27149,N_27807);
xnor U28815 (N_28815,N_27287,N_27273);
nand U28816 (N_28816,N_27807,N_27960);
and U28817 (N_28817,N_27777,N_27563);
nand U28818 (N_28818,N_27960,N_27990);
and U28819 (N_28819,N_27065,N_27676);
or U28820 (N_28820,N_27194,N_27612);
xor U28821 (N_28821,N_27038,N_27034);
nand U28822 (N_28822,N_27067,N_27794);
nand U28823 (N_28823,N_27576,N_27691);
and U28824 (N_28824,N_27565,N_27777);
or U28825 (N_28825,N_27264,N_27867);
nand U28826 (N_28826,N_27739,N_27541);
and U28827 (N_28827,N_27913,N_27512);
nor U28828 (N_28828,N_27953,N_27702);
and U28829 (N_28829,N_27143,N_27462);
and U28830 (N_28830,N_27696,N_27576);
xnor U28831 (N_28831,N_27755,N_27965);
xnor U28832 (N_28832,N_27045,N_27352);
nand U28833 (N_28833,N_27073,N_27686);
and U28834 (N_28834,N_27381,N_27681);
and U28835 (N_28835,N_27574,N_27265);
and U28836 (N_28836,N_27331,N_27609);
xor U28837 (N_28837,N_27821,N_27644);
and U28838 (N_28838,N_27223,N_27870);
and U28839 (N_28839,N_27700,N_27822);
and U28840 (N_28840,N_27833,N_27744);
or U28841 (N_28841,N_27860,N_27320);
xnor U28842 (N_28842,N_27283,N_27613);
or U28843 (N_28843,N_27316,N_27779);
xor U28844 (N_28844,N_27831,N_27519);
nand U28845 (N_28845,N_27537,N_27000);
nor U28846 (N_28846,N_27495,N_27591);
or U28847 (N_28847,N_27166,N_27412);
nand U28848 (N_28848,N_27557,N_27284);
and U28849 (N_28849,N_27446,N_27714);
nand U28850 (N_28850,N_27087,N_27864);
nor U28851 (N_28851,N_27267,N_27578);
nand U28852 (N_28852,N_27815,N_27368);
xnor U28853 (N_28853,N_27507,N_27062);
or U28854 (N_28854,N_27905,N_27545);
nand U28855 (N_28855,N_27956,N_27635);
nor U28856 (N_28856,N_27754,N_27239);
nand U28857 (N_28857,N_27843,N_27112);
and U28858 (N_28858,N_27409,N_27385);
and U28859 (N_28859,N_27144,N_27742);
nand U28860 (N_28860,N_27689,N_27369);
xor U28861 (N_28861,N_27055,N_27729);
and U28862 (N_28862,N_27301,N_27934);
nand U28863 (N_28863,N_27508,N_27744);
nand U28864 (N_28864,N_27971,N_27584);
and U28865 (N_28865,N_27340,N_27991);
nand U28866 (N_28866,N_27506,N_27697);
nor U28867 (N_28867,N_27882,N_27426);
nand U28868 (N_28868,N_27735,N_27504);
nand U28869 (N_28869,N_27922,N_27839);
nor U28870 (N_28870,N_27868,N_27088);
nand U28871 (N_28871,N_27933,N_27510);
and U28872 (N_28872,N_27083,N_27982);
xnor U28873 (N_28873,N_27058,N_27479);
nor U28874 (N_28874,N_27209,N_27092);
nor U28875 (N_28875,N_27194,N_27881);
xor U28876 (N_28876,N_27114,N_27105);
nor U28877 (N_28877,N_27160,N_27304);
or U28878 (N_28878,N_27814,N_27534);
or U28879 (N_28879,N_27616,N_27563);
nor U28880 (N_28880,N_27506,N_27997);
nor U28881 (N_28881,N_27634,N_27820);
and U28882 (N_28882,N_27105,N_27919);
xor U28883 (N_28883,N_27636,N_27173);
nor U28884 (N_28884,N_27310,N_27655);
nand U28885 (N_28885,N_27629,N_27262);
nand U28886 (N_28886,N_27587,N_27107);
or U28887 (N_28887,N_27993,N_27152);
nand U28888 (N_28888,N_27023,N_27073);
or U28889 (N_28889,N_27543,N_27156);
nor U28890 (N_28890,N_27773,N_27710);
xor U28891 (N_28891,N_27003,N_27493);
or U28892 (N_28892,N_27091,N_27568);
or U28893 (N_28893,N_27275,N_27263);
nand U28894 (N_28894,N_27783,N_27722);
or U28895 (N_28895,N_27085,N_27623);
nand U28896 (N_28896,N_27902,N_27077);
or U28897 (N_28897,N_27848,N_27929);
and U28898 (N_28898,N_27594,N_27634);
xnor U28899 (N_28899,N_27059,N_27533);
and U28900 (N_28900,N_27182,N_27348);
and U28901 (N_28901,N_27140,N_27814);
xor U28902 (N_28902,N_27343,N_27713);
nand U28903 (N_28903,N_27027,N_27552);
and U28904 (N_28904,N_27194,N_27058);
nand U28905 (N_28905,N_27978,N_27760);
nand U28906 (N_28906,N_27901,N_27097);
and U28907 (N_28907,N_27981,N_27283);
or U28908 (N_28908,N_27324,N_27481);
nand U28909 (N_28909,N_27807,N_27842);
nand U28910 (N_28910,N_27011,N_27198);
nor U28911 (N_28911,N_27660,N_27313);
xor U28912 (N_28912,N_27308,N_27480);
nand U28913 (N_28913,N_27910,N_27448);
or U28914 (N_28914,N_27412,N_27874);
or U28915 (N_28915,N_27516,N_27777);
xor U28916 (N_28916,N_27963,N_27910);
nand U28917 (N_28917,N_27057,N_27956);
or U28918 (N_28918,N_27962,N_27440);
or U28919 (N_28919,N_27152,N_27267);
nand U28920 (N_28920,N_27664,N_27171);
nand U28921 (N_28921,N_27265,N_27047);
nor U28922 (N_28922,N_27817,N_27569);
or U28923 (N_28923,N_27145,N_27015);
or U28924 (N_28924,N_27249,N_27389);
nor U28925 (N_28925,N_27945,N_27470);
or U28926 (N_28926,N_27646,N_27530);
or U28927 (N_28927,N_27337,N_27197);
or U28928 (N_28928,N_27545,N_27534);
nand U28929 (N_28929,N_27383,N_27853);
nor U28930 (N_28930,N_27913,N_27473);
and U28931 (N_28931,N_27674,N_27227);
nand U28932 (N_28932,N_27062,N_27438);
or U28933 (N_28933,N_27022,N_27152);
or U28934 (N_28934,N_27326,N_27662);
and U28935 (N_28935,N_27441,N_27343);
nor U28936 (N_28936,N_27092,N_27936);
xnor U28937 (N_28937,N_27245,N_27413);
and U28938 (N_28938,N_27223,N_27737);
nand U28939 (N_28939,N_27645,N_27308);
or U28940 (N_28940,N_27943,N_27507);
nor U28941 (N_28941,N_27689,N_27160);
and U28942 (N_28942,N_27010,N_27661);
and U28943 (N_28943,N_27205,N_27135);
nor U28944 (N_28944,N_27032,N_27930);
or U28945 (N_28945,N_27501,N_27212);
or U28946 (N_28946,N_27436,N_27784);
xor U28947 (N_28947,N_27928,N_27791);
or U28948 (N_28948,N_27273,N_27959);
xnor U28949 (N_28949,N_27296,N_27126);
nor U28950 (N_28950,N_27947,N_27149);
nor U28951 (N_28951,N_27288,N_27912);
nor U28952 (N_28952,N_27542,N_27995);
xnor U28953 (N_28953,N_27082,N_27515);
xor U28954 (N_28954,N_27197,N_27383);
or U28955 (N_28955,N_27268,N_27716);
nor U28956 (N_28956,N_27200,N_27053);
nor U28957 (N_28957,N_27803,N_27260);
nand U28958 (N_28958,N_27009,N_27800);
or U28959 (N_28959,N_27071,N_27840);
nand U28960 (N_28960,N_27365,N_27526);
nor U28961 (N_28961,N_27572,N_27542);
and U28962 (N_28962,N_27249,N_27006);
or U28963 (N_28963,N_27464,N_27281);
nor U28964 (N_28964,N_27472,N_27869);
nand U28965 (N_28965,N_27198,N_27835);
nor U28966 (N_28966,N_27004,N_27720);
xnor U28967 (N_28967,N_27450,N_27780);
or U28968 (N_28968,N_27721,N_27630);
and U28969 (N_28969,N_27957,N_27407);
xnor U28970 (N_28970,N_27856,N_27481);
or U28971 (N_28971,N_27571,N_27646);
and U28972 (N_28972,N_27135,N_27470);
and U28973 (N_28973,N_27687,N_27902);
xor U28974 (N_28974,N_27895,N_27590);
xor U28975 (N_28975,N_27591,N_27172);
and U28976 (N_28976,N_27588,N_27256);
xor U28977 (N_28977,N_27143,N_27042);
xor U28978 (N_28978,N_27271,N_27296);
or U28979 (N_28979,N_27174,N_27918);
or U28980 (N_28980,N_27878,N_27678);
nand U28981 (N_28981,N_27915,N_27776);
and U28982 (N_28982,N_27182,N_27419);
or U28983 (N_28983,N_27750,N_27154);
nor U28984 (N_28984,N_27505,N_27271);
and U28985 (N_28985,N_27415,N_27691);
nor U28986 (N_28986,N_27781,N_27135);
and U28987 (N_28987,N_27850,N_27428);
and U28988 (N_28988,N_27220,N_27795);
or U28989 (N_28989,N_27837,N_27753);
nand U28990 (N_28990,N_27578,N_27598);
and U28991 (N_28991,N_27734,N_27335);
nand U28992 (N_28992,N_27114,N_27834);
and U28993 (N_28993,N_27182,N_27737);
xor U28994 (N_28994,N_27742,N_27870);
nor U28995 (N_28995,N_27447,N_27757);
or U28996 (N_28996,N_27626,N_27849);
nor U28997 (N_28997,N_27120,N_27908);
nor U28998 (N_28998,N_27227,N_27707);
and U28999 (N_28999,N_27788,N_27451);
nor U29000 (N_29000,N_28435,N_28711);
xnor U29001 (N_29001,N_28847,N_28628);
xor U29002 (N_29002,N_28565,N_28553);
xor U29003 (N_29003,N_28930,N_28000);
xnor U29004 (N_29004,N_28952,N_28589);
or U29005 (N_29005,N_28498,N_28597);
nand U29006 (N_29006,N_28983,N_28904);
xnor U29007 (N_29007,N_28801,N_28095);
nand U29008 (N_29008,N_28272,N_28499);
nor U29009 (N_29009,N_28738,N_28773);
nor U29010 (N_29010,N_28433,N_28366);
and U29011 (N_29011,N_28003,N_28261);
or U29012 (N_29012,N_28294,N_28408);
and U29013 (N_29013,N_28196,N_28211);
nand U29014 (N_29014,N_28315,N_28251);
nor U29015 (N_29015,N_28919,N_28461);
and U29016 (N_29016,N_28041,N_28091);
nor U29017 (N_29017,N_28682,N_28683);
nand U29018 (N_29018,N_28198,N_28364);
nor U29019 (N_29019,N_28720,N_28101);
xnor U29020 (N_29020,N_28723,N_28579);
nor U29021 (N_29021,N_28910,N_28824);
nor U29022 (N_29022,N_28523,N_28921);
nand U29023 (N_29023,N_28977,N_28304);
or U29024 (N_29024,N_28854,N_28155);
nand U29025 (N_29025,N_28106,N_28451);
xor U29026 (N_29026,N_28354,N_28283);
nor U29027 (N_29027,N_28744,N_28885);
xor U29028 (N_29028,N_28163,N_28993);
nor U29029 (N_29029,N_28672,N_28244);
nor U29030 (N_29030,N_28607,N_28633);
nand U29031 (N_29031,N_28061,N_28753);
nor U29032 (N_29032,N_28317,N_28994);
xnor U29033 (N_29033,N_28956,N_28049);
nand U29034 (N_29034,N_28563,N_28782);
xor U29035 (N_29035,N_28120,N_28249);
nand U29036 (N_29036,N_28265,N_28800);
nand U29037 (N_29037,N_28180,N_28043);
or U29038 (N_29038,N_28159,N_28025);
or U29039 (N_29039,N_28403,N_28205);
nand U29040 (N_29040,N_28342,N_28743);
or U29041 (N_29041,N_28142,N_28503);
nand U29042 (N_29042,N_28221,N_28873);
nor U29043 (N_29043,N_28083,N_28989);
nor U29044 (N_29044,N_28543,N_28395);
nand U29045 (N_29045,N_28511,N_28680);
nand U29046 (N_29046,N_28588,N_28644);
or U29047 (N_29047,N_28538,N_28183);
or U29048 (N_29048,N_28526,N_28337);
or U29049 (N_29049,N_28259,N_28689);
xor U29050 (N_29050,N_28105,N_28379);
nor U29051 (N_29051,N_28604,N_28121);
xor U29052 (N_29052,N_28730,N_28102);
nor U29053 (N_29053,N_28750,N_28975);
and U29054 (N_29054,N_28030,N_28849);
nor U29055 (N_29055,N_28623,N_28314);
xnor U29056 (N_29056,N_28216,N_28243);
or U29057 (N_29057,N_28973,N_28616);
nand U29058 (N_29058,N_28137,N_28358);
nor U29059 (N_29059,N_28129,N_28088);
xor U29060 (N_29060,N_28039,N_28201);
nand U29061 (N_29061,N_28718,N_28475);
xor U29062 (N_29062,N_28762,N_28518);
nor U29063 (N_29063,N_28349,N_28869);
or U29064 (N_29064,N_28562,N_28751);
and U29065 (N_29065,N_28386,N_28681);
nand U29066 (N_29066,N_28587,N_28465);
and U29067 (N_29067,N_28996,N_28979);
xor U29068 (N_29068,N_28040,N_28027);
nand U29069 (N_29069,N_28731,N_28799);
and U29070 (N_29070,N_28146,N_28638);
or U29071 (N_29071,N_28482,N_28065);
xor U29072 (N_29072,N_28233,N_28104);
and U29073 (N_29073,N_28299,N_28405);
nand U29074 (N_29074,N_28640,N_28370);
and U29075 (N_29075,N_28365,N_28241);
nor U29076 (N_29076,N_28350,N_28019);
xor U29077 (N_29077,N_28046,N_28937);
xnor U29078 (N_29078,N_28504,N_28110);
or U29079 (N_29079,N_28319,N_28341);
or U29080 (N_29080,N_28207,N_28546);
xor U29081 (N_29081,N_28316,N_28918);
xnor U29082 (N_29082,N_28313,N_28428);
nor U29083 (N_29083,N_28085,N_28507);
nand U29084 (N_29084,N_28480,N_28577);
and U29085 (N_29085,N_28463,N_28974);
nand U29086 (N_29086,N_28410,N_28450);
nor U29087 (N_29087,N_28008,N_28360);
nor U29088 (N_29088,N_28510,N_28048);
xor U29089 (N_29089,N_28236,N_28182);
nor U29090 (N_29090,N_28111,N_28266);
and U29091 (N_29091,N_28339,N_28031);
xor U29092 (N_29092,N_28772,N_28479);
nor U29093 (N_29093,N_28281,N_28929);
nor U29094 (N_29094,N_28520,N_28760);
and U29095 (N_29095,N_28652,N_28914);
xnor U29096 (N_29096,N_28456,N_28462);
xor U29097 (N_29097,N_28164,N_28044);
xor U29098 (N_29098,N_28592,N_28246);
nand U29099 (N_29099,N_28225,N_28162);
xor U29100 (N_29100,N_28070,N_28492);
or U29101 (N_29101,N_28792,N_28861);
or U29102 (N_29102,N_28306,N_28122);
and U29103 (N_29103,N_28412,N_28785);
and U29104 (N_29104,N_28945,N_28856);
nor U29105 (N_29105,N_28813,N_28367);
xor U29106 (N_29106,N_28470,N_28627);
or U29107 (N_29107,N_28965,N_28344);
xnor U29108 (N_29108,N_28212,N_28896);
nor U29109 (N_29109,N_28015,N_28356);
or U29110 (N_29110,N_28431,N_28348);
nand U29111 (N_29111,N_28234,N_28999);
nor U29112 (N_29112,N_28312,N_28472);
or U29113 (N_29113,N_28735,N_28248);
or U29114 (N_29114,N_28815,N_28415);
nor U29115 (N_29115,N_28630,N_28264);
and U29116 (N_29116,N_28050,N_28571);
xnor U29117 (N_29117,N_28485,N_28136);
and U29118 (N_29118,N_28273,N_28926);
nand U29119 (N_29119,N_28399,N_28833);
nand U29120 (N_29120,N_28277,N_28798);
and U29121 (N_29121,N_28636,N_28330);
or U29122 (N_29122,N_28335,N_28508);
nor U29123 (N_29123,N_28840,N_28559);
xnor U29124 (N_29124,N_28852,N_28355);
and U29125 (N_29125,N_28222,N_28948);
nand U29126 (N_29126,N_28987,N_28900);
nor U29127 (N_29127,N_28867,N_28779);
and U29128 (N_29128,N_28497,N_28255);
or U29129 (N_29129,N_28823,N_28026);
xnor U29130 (N_29130,N_28758,N_28880);
nand U29131 (N_29131,N_28516,N_28686);
xnor U29132 (N_29132,N_28581,N_28804);
or U29133 (N_29133,N_28858,N_28641);
or U29134 (N_29134,N_28373,N_28915);
nand U29135 (N_29135,N_28547,N_28887);
xor U29136 (N_29136,N_28086,N_28401);
nor U29137 (N_29137,N_28906,N_28834);
or U29138 (N_29138,N_28156,N_28647);
and U29139 (N_29139,N_28981,N_28296);
xnor U29140 (N_29140,N_28634,N_28694);
and U29141 (N_29141,N_28862,N_28676);
nor U29142 (N_29142,N_28545,N_28580);
or U29143 (N_29143,N_28009,N_28584);
xor U29144 (N_29144,N_28097,N_28032);
nand U29145 (N_29145,N_28074,N_28194);
and U29146 (N_29146,N_28447,N_28883);
xor U29147 (N_29147,N_28971,N_28382);
nand U29148 (N_29148,N_28611,N_28837);
or U29149 (N_29149,N_28033,N_28420);
xnor U29150 (N_29150,N_28622,N_28899);
and U29151 (N_29151,N_28958,N_28171);
xor U29152 (N_29152,N_28615,N_28922);
and U29153 (N_29153,N_28489,N_28748);
nor U29154 (N_29154,N_28522,N_28071);
nor U29155 (N_29155,N_28712,N_28793);
nor U29156 (N_29156,N_28028,N_28903);
and U29157 (N_29157,N_28034,N_28671);
and U29158 (N_29158,N_28536,N_28181);
nand U29159 (N_29159,N_28960,N_28340);
or U29160 (N_29160,N_28232,N_28529);
and U29161 (N_29161,N_28651,N_28632);
nand U29162 (N_29162,N_28675,N_28307);
nor U29163 (N_29163,N_28590,N_28566);
nor U29164 (N_29164,N_28179,N_28139);
and U29165 (N_29165,N_28884,N_28116);
and U29166 (N_29166,N_28274,N_28667);
nor U29167 (N_29167,N_28016,N_28795);
nand U29168 (N_29168,N_28124,N_28661);
and U29169 (N_29169,N_28568,N_28911);
or U29170 (N_29170,N_28093,N_28333);
or U29171 (N_29171,N_28501,N_28717);
or U29172 (N_29172,N_28708,N_28542);
and U29173 (N_29173,N_28902,N_28662);
or U29174 (N_29174,N_28995,N_28178);
nand U29175 (N_29175,N_28893,N_28006);
nand U29176 (N_29176,N_28879,N_28453);
xnor U29177 (N_29177,N_28202,N_28610);
xor U29178 (N_29178,N_28092,N_28154);
and U29179 (N_29179,N_28690,N_28020);
nand U29180 (N_29180,N_28493,N_28371);
and U29181 (N_29181,N_28619,N_28505);
and U29182 (N_29182,N_28811,N_28514);
nand U29183 (N_29183,N_28646,N_28115);
nor U29184 (N_29184,N_28052,N_28208);
or U29185 (N_29185,N_28250,N_28305);
nand U29186 (N_29186,N_28318,N_28957);
and U29187 (N_29187,N_28186,N_28649);
and U29188 (N_29188,N_28368,N_28291);
and U29189 (N_29189,N_28013,N_28332);
and U29190 (N_29190,N_28007,N_28214);
xnor U29191 (N_29191,N_28416,N_28969);
nor U29192 (N_29192,N_28459,N_28362);
xnor U29193 (N_29193,N_28603,N_28444);
nand U29194 (N_29194,N_28912,N_28474);
xor U29195 (N_29195,N_28572,N_28099);
and U29196 (N_29196,N_28806,N_28369);
or U29197 (N_29197,N_28113,N_28190);
and U29198 (N_29198,N_28817,N_28696);
xnor U29199 (N_29199,N_28875,N_28509);
and U29200 (N_29200,N_28396,N_28173);
nor U29201 (N_29201,N_28169,N_28907);
xor U29202 (N_29202,N_28471,N_28068);
xor U29203 (N_29203,N_28483,N_28725);
and U29204 (N_29204,N_28950,N_28695);
and U29205 (N_29205,N_28557,N_28199);
nand U29206 (N_29206,N_28077,N_28160);
and U29207 (N_29207,N_28022,N_28004);
nand U29208 (N_29208,N_28018,N_28506);
nand U29209 (N_29209,N_28287,N_28716);
nand U29210 (N_29210,N_28601,N_28347);
nand U29211 (N_29211,N_28944,N_28011);
nand U29212 (N_29212,N_28949,N_28765);
xnor U29213 (N_29213,N_28147,N_28351);
or U29214 (N_29214,N_28037,N_28658);
and U29215 (N_29215,N_28374,N_28700);
xnor U29216 (N_29216,N_28998,N_28564);
and U29217 (N_29217,N_28103,N_28639);
nand U29218 (N_29218,N_28166,N_28413);
or U29219 (N_29219,N_28768,N_28901);
or U29220 (N_29220,N_28621,N_28593);
nand U29221 (N_29221,N_28684,N_28826);
nand U29222 (N_29222,N_28353,N_28531);
nor U29223 (N_29223,N_28786,N_28361);
or U29224 (N_29224,N_28802,N_28150);
nand U29225 (N_29225,N_28596,N_28814);
or U29226 (N_29226,N_28109,N_28775);
and U29227 (N_29227,N_28612,N_28528);
nand U29228 (N_29228,N_28059,N_28794);
nand U29229 (N_29229,N_28767,N_28189);
xor U29230 (N_29230,N_28582,N_28846);
nor U29231 (N_29231,N_28326,N_28323);
or U29232 (N_29232,N_28406,N_28737);
or U29233 (N_29233,N_28527,N_28674);
nor U29234 (N_29234,N_28935,N_28759);
xnor U29235 (N_29235,N_28943,N_28185);
nand U29236 (N_29236,N_28585,N_28325);
xor U29237 (N_29237,N_28739,N_28012);
and U29238 (N_29238,N_28978,N_28699);
nor U29239 (N_29239,N_28445,N_28336);
nand U29240 (N_29240,N_28439,N_28418);
nor U29241 (N_29241,N_28964,N_28057);
or U29242 (N_29242,N_28938,N_28787);
and U29243 (N_29243,N_28486,N_28831);
and U29244 (N_29244,N_28845,N_28388);
nor U29245 (N_29245,N_28732,N_28223);
xnor U29246 (N_29246,N_28567,N_28148);
xor U29247 (N_29247,N_28855,N_28275);
nand U29248 (N_29248,N_28532,N_28886);
nand U29249 (N_29249,N_28238,N_28770);
nand U29250 (N_29250,N_28829,N_28144);
or U29251 (N_29251,N_28835,N_28704);
nand U29252 (N_29252,N_28123,N_28311);
nand U29253 (N_29253,N_28158,N_28345);
nor U29254 (N_29254,N_28449,N_28766);
nor U29255 (N_29255,N_28905,N_28478);
nand U29256 (N_29256,N_28024,N_28613);
xnor U29257 (N_29257,N_28067,N_28942);
nand U29258 (N_29258,N_28962,N_28473);
nor U29259 (N_29259,N_28894,N_28108);
and U29260 (N_29260,N_28558,N_28090);
and U29261 (N_29261,N_28890,N_28087);
xor U29262 (N_29262,N_28437,N_28138);
or U29263 (N_29263,N_28828,N_28295);
nand U29264 (N_29264,N_28414,N_28728);
or U29265 (N_29265,N_28864,N_28913);
nand U29266 (N_29266,N_28170,N_28600);
and U29267 (N_29267,N_28502,N_28126);
or U29268 (N_29268,N_28286,N_28256);
nor U29269 (N_29269,N_28530,N_28062);
nand U29270 (N_29270,N_28594,N_28187);
and U29271 (N_29271,N_28084,N_28496);
and U29272 (N_29272,N_28177,N_28380);
nand U29273 (N_29273,N_28426,N_28320);
xnor U29274 (N_29274,N_28328,N_28818);
nand U29275 (N_29275,N_28288,N_28297);
nor U29276 (N_29276,N_28383,N_28719);
nor U29277 (N_29277,N_28573,N_28656);
nand U29278 (N_29278,N_28460,N_28733);
nor U29279 (N_29279,N_28740,N_28051);
or U29280 (N_29280,N_28678,N_28143);
nor U29281 (N_29281,N_28165,N_28014);
nor U29282 (N_29282,N_28219,N_28721);
and U29283 (N_29283,N_28617,N_28079);
nor U29284 (N_29284,N_28359,N_28583);
xnor U29285 (N_29285,N_28140,N_28534);
xnor U29286 (N_29286,N_28860,N_28832);
nand U29287 (N_29287,N_28591,N_28191);
nand U29288 (N_29288,N_28857,N_28430);
or U29289 (N_29289,N_28608,N_28218);
nand U29290 (N_29290,N_28217,N_28161);
and U29291 (N_29291,N_28643,N_28988);
xor U29292 (N_29292,N_28642,N_28245);
and U29293 (N_29293,N_28467,N_28931);
nor U29294 (N_29294,N_28796,N_28133);
nor U29295 (N_29295,N_28853,N_28363);
nand U29296 (N_29296,N_28434,N_28253);
and U29297 (N_29297,N_28544,N_28967);
nand U29298 (N_29298,N_28227,N_28820);
nor U29299 (N_29299,N_28292,N_28727);
or U29300 (N_29300,N_28394,N_28635);
nand U29301 (N_29301,N_28549,N_28803);
nor U29302 (N_29302,N_28118,N_28659);
nand U29303 (N_29303,N_28955,N_28290);
nand U29304 (N_29304,N_28512,N_28812);
and U29305 (N_29305,N_28454,N_28117);
nor U29306 (N_29306,N_28517,N_28045);
or U29307 (N_29307,N_28168,N_28329);
or U29308 (N_29308,N_28047,N_28539);
nor U29309 (N_29309,N_28665,N_28076);
nor U29310 (N_29310,N_28469,N_28660);
xor U29311 (N_29311,N_28747,N_28231);
or U29312 (N_29312,N_28822,N_28419);
nand U29313 (N_29313,N_28343,N_28936);
xnor U29314 (N_29314,N_28877,N_28764);
or U29315 (N_29315,N_28576,N_28677);
xnor U29316 (N_29316,N_28197,N_28407);
nor U29317 (N_29317,N_28586,N_28693);
nor U29318 (N_29318,N_28427,N_28188);
nand U29319 (N_29319,N_28980,N_28513);
nand U29320 (N_29320,N_28448,N_28392);
and U29321 (N_29321,N_28920,N_28230);
and U29322 (N_29322,N_28209,N_28494);
and U29323 (N_29323,N_28324,N_28540);
xnor U29324 (N_29324,N_28821,N_28081);
or U29325 (N_29325,N_28771,N_28206);
nor U29326 (N_29326,N_28002,N_28736);
nor U29327 (N_29327,N_28908,N_28954);
nand U29328 (N_29328,N_28114,N_28391);
or U29329 (N_29329,N_28816,N_28927);
nand U29330 (N_29330,N_28841,N_28058);
nand U29331 (N_29331,N_28490,N_28992);
xnor U29332 (N_29332,N_28038,N_28262);
nor U29333 (N_29333,N_28021,N_28859);
and U29334 (N_29334,N_28481,N_28986);
nor U29335 (N_29335,N_28226,N_28707);
or U29336 (N_29336,N_28664,N_28637);
xnor U29337 (N_29337,N_28280,N_28094);
nand U29338 (N_29338,N_28300,N_28703);
nor U29339 (N_29339,N_28174,N_28882);
nand U29340 (N_29340,N_28928,N_28881);
or U29341 (N_29341,N_28064,N_28655);
and U29342 (N_29342,N_28258,N_28670);
or U29343 (N_29343,N_28754,N_28001);
nor U29344 (N_29344,N_28135,N_28519);
and U29345 (N_29345,N_28521,N_28119);
and U29346 (N_29346,N_28863,N_28278);
nand U29347 (N_29347,N_28100,N_28741);
or U29348 (N_29348,N_28263,N_28790);
and U29349 (N_29349,N_28533,N_28152);
nand U29350 (N_29350,N_28443,N_28215);
nand U29351 (N_29351,N_28868,N_28078);
nand U29352 (N_29352,N_28252,N_28404);
nor U29353 (N_29353,N_28897,N_28606);
or U29354 (N_29354,N_28555,N_28130);
nand U29355 (N_29355,N_28247,N_28836);
nor U29356 (N_29356,N_28387,N_28458);
or U29357 (N_29357,N_28271,N_28784);
nand U29358 (N_29358,N_28609,N_28301);
nor U29359 (N_29359,N_28865,N_28982);
xnor U29360 (N_29360,N_28346,N_28552);
nor U29361 (N_29361,N_28310,N_28334);
nand U29362 (N_29362,N_28734,N_28213);
or U29363 (N_29363,N_28618,N_28438);
nand U29364 (N_29364,N_28060,N_28710);
xor U29365 (N_29365,N_28035,N_28331);
or U29366 (N_29366,N_28745,N_28551);
xnor U29367 (N_29367,N_28424,N_28228);
nand U29368 (N_29368,N_28172,N_28303);
xor U29369 (N_29369,N_28848,N_28535);
and U29370 (N_29370,N_28941,N_28688);
and U29371 (N_29371,N_28440,N_28276);
nand U29372 (N_29372,N_28267,N_28560);
xor U29373 (N_29373,N_28153,N_28279);
xor U29374 (N_29374,N_28200,N_28176);
nand U29375 (N_29375,N_28780,N_28805);
xnor U29376 (N_29376,N_28080,N_28175);
xnor U29377 (N_29377,N_28484,N_28570);
or U29378 (N_29378,N_28569,N_28763);
nand U29379 (N_29379,N_28878,N_28838);
nand U29380 (N_29380,N_28605,N_28556);
and U29381 (N_29381,N_28839,N_28891);
nand U29382 (N_29382,N_28237,N_28774);
and U29383 (N_29383,N_28352,N_28970);
xor U29384 (N_29384,N_28706,N_28697);
nand U29385 (N_29385,N_28436,N_28010);
nor U29386 (N_29386,N_28691,N_28871);
and U29387 (N_29387,N_28224,N_28575);
nor U29388 (N_29388,N_28284,N_28916);
and U29389 (N_29389,N_28749,N_28476);
or U29390 (N_29390,N_28089,N_28017);
and U29391 (N_29391,N_28417,N_28468);
and U29392 (N_29392,N_28631,N_28477);
or U29393 (N_29393,N_28289,N_28705);
xnor U29394 (N_29394,N_28654,N_28141);
nor U29395 (N_29395,N_28425,N_28423);
xnor U29396 (N_29396,N_28066,N_28429);
or U29397 (N_29397,N_28193,N_28385);
nor U29398 (N_29398,N_28776,N_28872);
nor U29399 (N_29399,N_28554,N_28726);
nand U29400 (N_29400,N_28843,N_28112);
xnor U29401 (N_29401,N_28242,N_28714);
nand U29402 (N_29402,N_28309,N_28491);
and U29403 (N_29403,N_28338,N_28807);
and U29404 (N_29404,N_28679,N_28107);
or U29405 (N_29405,N_28537,N_28073);
xnor U29406 (N_29406,N_28402,N_28939);
or U29407 (N_29407,N_28932,N_28808);
nand U29408 (N_29408,N_28599,N_28151);
nand U29409 (N_29409,N_28614,N_28783);
nor U29410 (N_29410,N_28398,N_28825);
and U29411 (N_29411,N_28844,N_28327);
or U29412 (N_29412,N_28809,N_28777);
nor U29413 (N_29413,N_28963,N_28550);
nand U29414 (N_29414,N_28072,N_28874);
or U29415 (N_29415,N_28457,N_28959);
nor U29416 (N_29416,N_28561,N_28991);
and U29417 (N_29417,N_28372,N_28663);
and U29418 (N_29418,N_28953,N_28668);
xor U29419 (N_29419,N_28257,N_28895);
nand U29420 (N_29420,N_28990,N_28381);
nor U29421 (N_29421,N_28761,N_28357);
nor U29422 (N_29422,N_28029,N_28925);
or U29423 (N_29423,N_28966,N_28254);
and U29424 (N_29424,N_28446,N_28645);
and U29425 (N_29425,N_28204,N_28673);
and U29426 (N_29426,N_28778,N_28149);
xor U29427 (N_29427,N_28713,N_28466);
nor U29428 (N_29428,N_28791,N_28432);
nand U29429 (N_29429,N_28023,N_28192);
nor U29430 (N_29430,N_28229,N_28270);
nand U29431 (N_29431,N_28653,N_28602);
xnor U29432 (N_29432,N_28898,N_28082);
xnor U29433 (N_29433,N_28648,N_28715);
and U29434 (N_29434,N_28260,N_28390);
or U29435 (N_29435,N_28240,N_28378);
or U29436 (N_29436,N_28524,N_28629);
or U29437 (N_29437,N_28157,N_28709);
nand U29438 (N_29438,N_28195,N_28298);
or U29439 (N_29439,N_28624,N_28598);
nor U29440 (N_29440,N_28220,N_28293);
nor U29441 (N_29441,N_28620,N_28042);
and U29442 (N_29442,N_28452,N_28495);
nor U29443 (N_29443,N_28742,N_28375);
or U29444 (N_29444,N_28282,N_28924);
nor U29445 (N_29445,N_28757,N_28909);
xor U29446 (N_29446,N_28203,N_28525);
nor U29447 (N_29447,N_28053,N_28923);
or U29448 (N_29448,N_28578,N_28827);
nor U29449 (N_29449,N_28400,N_28934);
and U29450 (N_29450,N_28626,N_28917);
xnor U29451 (N_29451,N_28167,N_28698);
xor U29452 (N_29452,N_28892,N_28666);
and U29453 (N_29453,N_28889,N_28746);
or U29454 (N_29454,N_28384,N_28876);
or U29455 (N_29455,N_28131,N_28830);
xor U29456 (N_29456,N_28625,N_28036);
nor U29457 (N_29457,N_28850,N_28132);
and U29458 (N_29458,N_28724,N_28984);
nand U29459 (N_29459,N_28968,N_28797);
or U29460 (N_29460,N_28184,N_28393);
nand U29461 (N_29461,N_28075,N_28389);
nand U29462 (N_29462,N_28268,N_28756);
nand U29463 (N_29463,N_28722,N_28870);
xnor U29464 (N_29464,N_28054,N_28789);
nand U29465 (N_29465,N_28541,N_28692);
nand U29466 (N_29466,N_28210,N_28657);
nor U29467 (N_29467,N_28976,N_28866);
nor U29468 (N_29468,N_28500,N_28302);
and U29469 (N_29469,N_28933,N_28888);
nor U29470 (N_29470,N_28687,N_28422);
or U29471 (N_29471,N_28997,N_28755);
nand U29472 (N_29472,N_28810,N_28377);
xor U29473 (N_29473,N_28441,N_28285);
and U29474 (N_29474,N_28701,N_28239);
nand U29475 (N_29475,N_28972,N_28411);
nand U29476 (N_29476,N_28488,N_28851);
or U29477 (N_29477,N_28769,N_28781);
nand U29478 (N_29478,N_28421,N_28397);
nor U29479 (N_29479,N_28134,N_28145);
and U29480 (N_29480,N_28055,N_28702);
xnor U29481 (N_29481,N_28788,N_28961);
nand U29482 (N_29482,N_28985,N_28752);
and U29483 (N_29483,N_28128,N_28063);
or U29484 (N_29484,N_28269,N_28308);
nand U29485 (N_29485,N_28515,N_28951);
nand U29486 (N_29486,N_28056,N_28322);
xor U29487 (N_29487,N_28574,N_28005);
nor U29488 (N_29488,N_28487,N_28455);
and U29489 (N_29489,N_28685,N_28096);
xor U29490 (N_29490,N_28442,N_28947);
or U29491 (N_29491,N_28098,N_28595);
and U29492 (N_29492,N_28376,N_28464);
nor U29493 (N_29493,N_28940,N_28548);
xnor U29494 (N_29494,N_28669,N_28235);
nor U29495 (N_29495,N_28729,N_28819);
or U29496 (N_29496,N_28650,N_28125);
xnor U29497 (N_29497,N_28321,N_28069);
and U29498 (N_29498,N_28946,N_28842);
or U29499 (N_29499,N_28409,N_28127);
or U29500 (N_29500,N_28214,N_28188);
or U29501 (N_29501,N_28996,N_28127);
xor U29502 (N_29502,N_28112,N_28690);
and U29503 (N_29503,N_28622,N_28426);
or U29504 (N_29504,N_28498,N_28249);
xor U29505 (N_29505,N_28883,N_28607);
xor U29506 (N_29506,N_28012,N_28349);
and U29507 (N_29507,N_28548,N_28920);
nor U29508 (N_29508,N_28711,N_28215);
or U29509 (N_29509,N_28068,N_28679);
nor U29510 (N_29510,N_28933,N_28447);
nand U29511 (N_29511,N_28569,N_28297);
or U29512 (N_29512,N_28317,N_28086);
nor U29513 (N_29513,N_28827,N_28258);
or U29514 (N_29514,N_28332,N_28507);
nand U29515 (N_29515,N_28315,N_28407);
nor U29516 (N_29516,N_28533,N_28782);
nand U29517 (N_29517,N_28668,N_28859);
nand U29518 (N_29518,N_28044,N_28863);
nor U29519 (N_29519,N_28079,N_28625);
xor U29520 (N_29520,N_28148,N_28144);
or U29521 (N_29521,N_28477,N_28481);
xnor U29522 (N_29522,N_28120,N_28924);
and U29523 (N_29523,N_28480,N_28429);
nand U29524 (N_29524,N_28110,N_28727);
nand U29525 (N_29525,N_28802,N_28643);
xor U29526 (N_29526,N_28587,N_28898);
nor U29527 (N_29527,N_28530,N_28884);
and U29528 (N_29528,N_28191,N_28711);
nor U29529 (N_29529,N_28575,N_28056);
or U29530 (N_29530,N_28169,N_28816);
or U29531 (N_29531,N_28244,N_28134);
nor U29532 (N_29532,N_28477,N_28031);
nor U29533 (N_29533,N_28695,N_28353);
nand U29534 (N_29534,N_28247,N_28977);
nor U29535 (N_29535,N_28236,N_28942);
xnor U29536 (N_29536,N_28131,N_28342);
nor U29537 (N_29537,N_28477,N_28286);
xor U29538 (N_29538,N_28679,N_28735);
or U29539 (N_29539,N_28177,N_28383);
nor U29540 (N_29540,N_28773,N_28178);
nand U29541 (N_29541,N_28643,N_28602);
or U29542 (N_29542,N_28229,N_28520);
or U29543 (N_29543,N_28952,N_28625);
and U29544 (N_29544,N_28867,N_28398);
and U29545 (N_29545,N_28112,N_28376);
xor U29546 (N_29546,N_28565,N_28571);
nor U29547 (N_29547,N_28522,N_28730);
nand U29548 (N_29548,N_28134,N_28296);
or U29549 (N_29549,N_28867,N_28085);
nand U29550 (N_29550,N_28401,N_28303);
xnor U29551 (N_29551,N_28841,N_28859);
nor U29552 (N_29552,N_28994,N_28458);
nor U29553 (N_29553,N_28908,N_28387);
and U29554 (N_29554,N_28598,N_28428);
and U29555 (N_29555,N_28153,N_28689);
nand U29556 (N_29556,N_28445,N_28586);
nor U29557 (N_29557,N_28915,N_28103);
xor U29558 (N_29558,N_28227,N_28752);
nand U29559 (N_29559,N_28839,N_28732);
or U29560 (N_29560,N_28890,N_28612);
nor U29561 (N_29561,N_28773,N_28673);
and U29562 (N_29562,N_28824,N_28772);
nand U29563 (N_29563,N_28952,N_28671);
xor U29564 (N_29564,N_28375,N_28729);
nor U29565 (N_29565,N_28395,N_28514);
nor U29566 (N_29566,N_28004,N_28629);
or U29567 (N_29567,N_28168,N_28791);
nand U29568 (N_29568,N_28366,N_28377);
nand U29569 (N_29569,N_28104,N_28323);
or U29570 (N_29570,N_28646,N_28360);
or U29571 (N_29571,N_28702,N_28865);
or U29572 (N_29572,N_28247,N_28551);
xor U29573 (N_29573,N_28309,N_28163);
and U29574 (N_29574,N_28939,N_28526);
and U29575 (N_29575,N_28265,N_28728);
nand U29576 (N_29576,N_28505,N_28325);
nand U29577 (N_29577,N_28695,N_28731);
nor U29578 (N_29578,N_28495,N_28089);
xor U29579 (N_29579,N_28090,N_28452);
nor U29580 (N_29580,N_28376,N_28737);
and U29581 (N_29581,N_28285,N_28658);
xnor U29582 (N_29582,N_28379,N_28867);
and U29583 (N_29583,N_28409,N_28744);
xor U29584 (N_29584,N_28568,N_28887);
nor U29585 (N_29585,N_28988,N_28420);
or U29586 (N_29586,N_28620,N_28219);
nand U29587 (N_29587,N_28971,N_28385);
nand U29588 (N_29588,N_28421,N_28616);
and U29589 (N_29589,N_28776,N_28157);
and U29590 (N_29590,N_28546,N_28344);
or U29591 (N_29591,N_28361,N_28992);
xor U29592 (N_29592,N_28038,N_28256);
or U29593 (N_29593,N_28440,N_28442);
or U29594 (N_29594,N_28437,N_28638);
or U29595 (N_29595,N_28794,N_28374);
or U29596 (N_29596,N_28121,N_28782);
or U29597 (N_29597,N_28467,N_28299);
nand U29598 (N_29598,N_28110,N_28799);
or U29599 (N_29599,N_28573,N_28363);
or U29600 (N_29600,N_28872,N_28711);
or U29601 (N_29601,N_28211,N_28233);
xor U29602 (N_29602,N_28807,N_28576);
and U29603 (N_29603,N_28386,N_28630);
nor U29604 (N_29604,N_28518,N_28340);
or U29605 (N_29605,N_28427,N_28877);
nor U29606 (N_29606,N_28822,N_28844);
or U29607 (N_29607,N_28475,N_28627);
xnor U29608 (N_29608,N_28243,N_28183);
and U29609 (N_29609,N_28538,N_28280);
nor U29610 (N_29610,N_28488,N_28908);
and U29611 (N_29611,N_28447,N_28100);
nor U29612 (N_29612,N_28911,N_28313);
or U29613 (N_29613,N_28119,N_28692);
and U29614 (N_29614,N_28835,N_28877);
xnor U29615 (N_29615,N_28599,N_28851);
xor U29616 (N_29616,N_28495,N_28868);
nor U29617 (N_29617,N_28578,N_28975);
nand U29618 (N_29618,N_28044,N_28107);
and U29619 (N_29619,N_28940,N_28606);
or U29620 (N_29620,N_28628,N_28719);
or U29621 (N_29621,N_28941,N_28008);
nand U29622 (N_29622,N_28198,N_28107);
nand U29623 (N_29623,N_28466,N_28749);
nor U29624 (N_29624,N_28317,N_28478);
nor U29625 (N_29625,N_28018,N_28631);
nand U29626 (N_29626,N_28676,N_28967);
xnor U29627 (N_29627,N_28375,N_28886);
nor U29628 (N_29628,N_28882,N_28775);
or U29629 (N_29629,N_28514,N_28163);
nor U29630 (N_29630,N_28693,N_28345);
or U29631 (N_29631,N_28055,N_28042);
or U29632 (N_29632,N_28883,N_28660);
xnor U29633 (N_29633,N_28167,N_28549);
xor U29634 (N_29634,N_28433,N_28739);
and U29635 (N_29635,N_28107,N_28573);
or U29636 (N_29636,N_28467,N_28759);
nor U29637 (N_29637,N_28369,N_28993);
nor U29638 (N_29638,N_28856,N_28160);
and U29639 (N_29639,N_28431,N_28284);
and U29640 (N_29640,N_28559,N_28573);
nor U29641 (N_29641,N_28742,N_28886);
xnor U29642 (N_29642,N_28435,N_28696);
or U29643 (N_29643,N_28601,N_28961);
and U29644 (N_29644,N_28176,N_28704);
and U29645 (N_29645,N_28034,N_28265);
nand U29646 (N_29646,N_28812,N_28312);
nand U29647 (N_29647,N_28352,N_28188);
nand U29648 (N_29648,N_28955,N_28447);
nand U29649 (N_29649,N_28400,N_28220);
or U29650 (N_29650,N_28825,N_28507);
xor U29651 (N_29651,N_28019,N_28516);
xnor U29652 (N_29652,N_28295,N_28379);
or U29653 (N_29653,N_28894,N_28408);
and U29654 (N_29654,N_28714,N_28423);
or U29655 (N_29655,N_28697,N_28329);
xor U29656 (N_29656,N_28039,N_28474);
xnor U29657 (N_29657,N_28989,N_28011);
and U29658 (N_29658,N_28331,N_28773);
nor U29659 (N_29659,N_28572,N_28513);
and U29660 (N_29660,N_28054,N_28002);
xor U29661 (N_29661,N_28249,N_28199);
nor U29662 (N_29662,N_28271,N_28436);
nor U29663 (N_29663,N_28463,N_28488);
nor U29664 (N_29664,N_28963,N_28450);
nor U29665 (N_29665,N_28281,N_28963);
or U29666 (N_29666,N_28578,N_28708);
xor U29667 (N_29667,N_28540,N_28386);
nor U29668 (N_29668,N_28038,N_28260);
nor U29669 (N_29669,N_28045,N_28241);
and U29670 (N_29670,N_28953,N_28868);
nor U29671 (N_29671,N_28975,N_28462);
xor U29672 (N_29672,N_28028,N_28775);
and U29673 (N_29673,N_28415,N_28368);
xor U29674 (N_29674,N_28685,N_28524);
nor U29675 (N_29675,N_28423,N_28661);
nand U29676 (N_29676,N_28727,N_28378);
or U29677 (N_29677,N_28452,N_28379);
nand U29678 (N_29678,N_28004,N_28933);
nor U29679 (N_29679,N_28423,N_28820);
or U29680 (N_29680,N_28391,N_28498);
xor U29681 (N_29681,N_28375,N_28515);
or U29682 (N_29682,N_28432,N_28225);
and U29683 (N_29683,N_28450,N_28353);
or U29684 (N_29684,N_28506,N_28640);
or U29685 (N_29685,N_28085,N_28989);
nor U29686 (N_29686,N_28760,N_28826);
nor U29687 (N_29687,N_28041,N_28721);
or U29688 (N_29688,N_28189,N_28259);
xor U29689 (N_29689,N_28801,N_28400);
nand U29690 (N_29690,N_28010,N_28251);
or U29691 (N_29691,N_28839,N_28818);
nand U29692 (N_29692,N_28424,N_28427);
xor U29693 (N_29693,N_28146,N_28002);
nor U29694 (N_29694,N_28502,N_28799);
nand U29695 (N_29695,N_28094,N_28197);
or U29696 (N_29696,N_28218,N_28263);
and U29697 (N_29697,N_28571,N_28457);
nand U29698 (N_29698,N_28293,N_28077);
or U29699 (N_29699,N_28316,N_28350);
nor U29700 (N_29700,N_28231,N_28003);
nor U29701 (N_29701,N_28096,N_28456);
xnor U29702 (N_29702,N_28954,N_28309);
or U29703 (N_29703,N_28105,N_28486);
and U29704 (N_29704,N_28628,N_28210);
nor U29705 (N_29705,N_28602,N_28576);
or U29706 (N_29706,N_28316,N_28539);
nand U29707 (N_29707,N_28908,N_28898);
nor U29708 (N_29708,N_28421,N_28623);
xnor U29709 (N_29709,N_28447,N_28079);
and U29710 (N_29710,N_28031,N_28809);
or U29711 (N_29711,N_28318,N_28902);
and U29712 (N_29712,N_28737,N_28853);
nand U29713 (N_29713,N_28869,N_28389);
nor U29714 (N_29714,N_28241,N_28523);
xor U29715 (N_29715,N_28799,N_28181);
or U29716 (N_29716,N_28524,N_28681);
nand U29717 (N_29717,N_28913,N_28515);
nor U29718 (N_29718,N_28060,N_28769);
nand U29719 (N_29719,N_28586,N_28107);
or U29720 (N_29720,N_28260,N_28981);
xor U29721 (N_29721,N_28026,N_28492);
or U29722 (N_29722,N_28148,N_28849);
xor U29723 (N_29723,N_28310,N_28331);
nor U29724 (N_29724,N_28608,N_28164);
xnor U29725 (N_29725,N_28047,N_28715);
nor U29726 (N_29726,N_28726,N_28928);
xnor U29727 (N_29727,N_28691,N_28788);
xnor U29728 (N_29728,N_28649,N_28938);
or U29729 (N_29729,N_28827,N_28086);
or U29730 (N_29730,N_28235,N_28302);
and U29731 (N_29731,N_28518,N_28746);
xor U29732 (N_29732,N_28683,N_28081);
or U29733 (N_29733,N_28233,N_28829);
nor U29734 (N_29734,N_28911,N_28760);
xnor U29735 (N_29735,N_28234,N_28534);
nand U29736 (N_29736,N_28426,N_28179);
xor U29737 (N_29737,N_28219,N_28363);
nand U29738 (N_29738,N_28958,N_28866);
xor U29739 (N_29739,N_28000,N_28672);
nor U29740 (N_29740,N_28112,N_28629);
or U29741 (N_29741,N_28460,N_28493);
and U29742 (N_29742,N_28407,N_28735);
nand U29743 (N_29743,N_28500,N_28962);
nor U29744 (N_29744,N_28904,N_28238);
nor U29745 (N_29745,N_28531,N_28049);
and U29746 (N_29746,N_28707,N_28138);
and U29747 (N_29747,N_28581,N_28419);
and U29748 (N_29748,N_28310,N_28963);
or U29749 (N_29749,N_28258,N_28671);
nor U29750 (N_29750,N_28404,N_28495);
xor U29751 (N_29751,N_28934,N_28779);
and U29752 (N_29752,N_28291,N_28466);
and U29753 (N_29753,N_28195,N_28153);
nor U29754 (N_29754,N_28749,N_28619);
or U29755 (N_29755,N_28174,N_28899);
nand U29756 (N_29756,N_28058,N_28724);
xor U29757 (N_29757,N_28780,N_28071);
nor U29758 (N_29758,N_28794,N_28259);
and U29759 (N_29759,N_28650,N_28784);
and U29760 (N_29760,N_28767,N_28291);
nand U29761 (N_29761,N_28779,N_28572);
or U29762 (N_29762,N_28059,N_28180);
and U29763 (N_29763,N_28898,N_28087);
nand U29764 (N_29764,N_28217,N_28184);
nor U29765 (N_29765,N_28493,N_28147);
or U29766 (N_29766,N_28735,N_28503);
or U29767 (N_29767,N_28011,N_28898);
xor U29768 (N_29768,N_28324,N_28482);
nand U29769 (N_29769,N_28035,N_28509);
or U29770 (N_29770,N_28874,N_28014);
nand U29771 (N_29771,N_28123,N_28818);
xnor U29772 (N_29772,N_28215,N_28823);
or U29773 (N_29773,N_28658,N_28409);
nand U29774 (N_29774,N_28228,N_28788);
nor U29775 (N_29775,N_28045,N_28668);
nand U29776 (N_29776,N_28153,N_28489);
nor U29777 (N_29777,N_28589,N_28311);
nand U29778 (N_29778,N_28395,N_28735);
nand U29779 (N_29779,N_28407,N_28089);
nand U29780 (N_29780,N_28260,N_28655);
or U29781 (N_29781,N_28782,N_28546);
xnor U29782 (N_29782,N_28547,N_28002);
nor U29783 (N_29783,N_28099,N_28063);
xnor U29784 (N_29784,N_28013,N_28420);
or U29785 (N_29785,N_28430,N_28498);
nand U29786 (N_29786,N_28537,N_28387);
nand U29787 (N_29787,N_28767,N_28356);
xor U29788 (N_29788,N_28652,N_28556);
nand U29789 (N_29789,N_28510,N_28406);
or U29790 (N_29790,N_28599,N_28030);
xor U29791 (N_29791,N_28607,N_28558);
nand U29792 (N_29792,N_28997,N_28285);
or U29793 (N_29793,N_28749,N_28623);
or U29794 (N_29794,N_28004,N_28875);
and U29795 (N_29795,N_28915,N_28925);
and U29796 (N_29796,N_28375,N_28290);
or U29797 (N_29797,N_28164,N_28315);
nand U29798 (N_29798,N_28242,N_28289);
nand U29799 (N_29799,N_28319,N_28634);
or U29800 (N_29800,N_28228,N_28993);
and U29801 (N_29801,N_28612,N_28095);
nor U29802 (N_29802,N_28663,N_28692);
xnor U29803 (N_29803,N_28741,N_28657);
and U29804 (N_29804,N_28886,N_28798);
nor U29805 (N_29805,N_28489,N_28006);
nand U29806 (N_29806,N_28689,N_28101);
nand U29807 (N_29807,N_28014,N_28830);
xor U29808 (N_29808,N_28302,N_28551);
xnor U29809 (N_29809,N_28743,N_28788);
or U29810 (N_29810,N_28876,N_28345);
nand U29811 (N_29811,N_28749,N_28126);
or U29812 (N_29812,N_28531,N_28945);
and U29813 (N_29813,N_28364,N_28072);
nand U29814 (N_29814,N_28682,N_28066);
or U29815 (N_29815,N_28566,N_28932);
nor U29816 (N_29816,N_28845,N_28140);
nand U29817 (N_29817,N_28115,N_28754);
nand U29818 (N_29818,N_28763,N_28481);
and U29819 (N_29819,N_28325,N_28983);
xnor U29820 (N_29820,N_28517,N_28660);
or U29821 (N_29821,N_28698,N_28101);
xnor U29822 (N_29822,N_28894,N_28483);
nand U29823 (N_29823,N_28965,N_28030);
nand U29824 (N_29824,N_28443,N_28921);
nand U29825 (N_29825,N_28533,N_28109);
nor U29826 (N_29826,N_28015,N_28228);
nor U29827 (N_29827,N_28757,N_28237);
xnor U29828 (N_29828,N_28024,N_28228);
or U29829 (N_29829,N_28878,N_28432);
nor U29830 (N_29830,N_28683,N_28744);
and U29831 (N_29831,N_28858,N_28077);
nand U29832 (N_29832,N_28952,N_28493);
nor U29833 (N_29833,N_28783,N_28957);
nor U29834 (N_29834,N_28949,N_28561);
and U29835 (N_29835,N_28144,N_28577);
or U29836 (N_29836,N_28462,N_28823);
and U29837 (N_29837,N_28091,N_28836);
or U29838 (N_29838,N_28121,N_28624);
nor U29839 (N_29839,N_28484,N_28930);
xor U29840 (N_29840,N_28827,N_28526);
nor U29841 (N_29841,N_28717,N_28411);
xnor U29842 (N_29842,N_28487,N_28880);
nand U29843 (N_29843,N_28073,N_28195);
and U29844 (N_29844,N_28988,N_28782);
nor U29845 (N_29845,N_28350,N_28407);
xor U29846 (N_29846,N_28364,N_28058);
nand U29847 (N_29847,N_28571,N_28746);
xnor U29848 (N_29848,N_28730,N_28700);
xor U29849 (N_29849,N_28441,N_28421);
or U29850 (N_29850,N_28231,N_28098);
and U29851 (N_29851,N_28462,N_28030);
or U29852 (N_29852,N_28758,N_28735);
nor U29853 (N_29853,N_28038,N_28379);
nand U29854 (N_29854,N_28951,N_28720);
or U29855 (N_29855,N_28888,N_28294);
or U29856 (N_29856,N_28492,N_28675);
or U29857 (N_29857,N_28386,N_28733);
and U29858 (N_29858,N_28674,N_28683);
xor U29859 (N_29859,N_28379,N_28787);
and U29860 (N_29860,N_28309,N_28132);
nor U29861 (N_29861,N_28244,N_28421);
or U29862 (N_29862,N_28519,N_28242);
nor U29863 (N_29863,N_28966,N_28006);
and U29864 (N_29864,N_28253,N_28587);
xnor U29865 (N_29865,N_28613,N_28247);
nor U29866 (N_29866,N_28173,N_28052);
xnor U29867 (N_29867,N_28143,N_28822);
or U29868 (N_29868,N_28623,N_28722);
and U29869 (N_29869,N_28904,N_28780);
and U29870 (N_29870,N_28590,N_28797);
xnor U29871 (N_29871,N_28687,N_28743);
xnor U29872 (N_29872,N_28383,N_28404);
nand U29873 (N_29873,N_28728,N_28568);
or U29874 (N_29874,N_28766,N_28303);
xor U29875 (N_29875,N_28906,N_28038);
xor U29876 (N_29876,N_28707,N_28112);
or U29877 (N_29877,N_28626,N_28391);
and U29878 (N_29878,N_28533,N_28610);
and U29879 (N_29879,N_28280,N_28474);
and U29880 (N_29880,N_28209,N_28730);
nor U29881 (N_29881,N_28609,N_28045);
xor U29882 (N_29882,N_28904,N_28525);
xor U29883 (N_29883,N_28073,N_28062);
or U29884 (N_29884,N_28096,N_28637);
xnor U29885 (N_29885,N_28187,N_28022);
nand U29886 (N_29886,N_28371,N_28159);
or U29887 (N_29887,N_28743,N_28496);
xnor U29888 (N_29888,N_28470,N_28509);
nand U29889 (N_29889,N_28118,N_28393);
or U29890 (N_29890,N_28305,N_28550);
nor U29891 (N_29891,N_28428,N_28559);
and U29892 (N_29892,N_28339,N_28102);
nor U29893 (N_29893,N_28601,N_28864);
or U29894 (N_29894,N_28529,N_28302);
xnor U29895 (N_29895,N_28458,N_28091);
nand U29896 (N_29896,N_28441,N_28813);
and U29897 (N_29897,N_28546,N_28192);
and U29898 (N_29898,N_28608,N_28040);
nand U29899 (N_29899,N_28246,N_28660);
or U29900 (N_29900,N_28245,N_28857);
and U29901 (N_29901,N_28329,N_28274);
and U29902 (N_29902,N_28669,N_28716);
or U29903 (N_29903,N_28216,N_28045);
nand U29904 (N_29904,N_28756,N_28567);
nor U29905 (N_29905,N_28564,N_28213);
xor U29906 (N_29906,N_28025,N_28240);
nor U29907 (N_29907,N_28207,N_28810);
nor U29908 (N_29908,N_28176,N_28901);
nor U29909 (N_29909,N_28623,N_28269);
nand U29910 (N_29910,N_28918,N_28024);
nor U29911 (N_29911,N_28842,N_28994);
xnor U29912 (N_29912,N_28909,N_28556);
nand U29913 (N_29913,N_28470,N_28354);
nand U29914 (N_29914,N_28808,N_28788);
or U29915 (N_29915,N_28202,N_28562);
nand U29916 (N_29916,N_28968,N_28911);
nor U29917 (N_29917,N_28200,N_28724);
xor U29918 (N_29918,N_28873,N_28643);
or U29919 (N_29919,N_28930,N_28540);
and U29920 (N_29920,N_28563,N_28841);
nor U29921 (N_29921,N_28601,N_28351);
nand U29922 (N_29922,N_28464,N_28941);
or U29923 (N_29923,N_28695,N_28668);
nand U29924 (N_29924,N_28093,N_28941);
xor U29925 (N_29925,N_28533,N_28015);
nor U29926 (N_29926,N_28752,N_28255);
xor U29927 (N_29927,N_28074,N_28980);
nor U29928 (N_29928,N_28895,N_28897);
nand U29929 (N_29929,N_28232,N_28591);
nand U29930 (N_29930,N_28739,N_28797);
and U29931 (N_29931,N_28285,N_28303);
nand U29932 (N_29932,N_28528,N_28954);
xor U29933 (N_29933,N_28266,N_28759);
xnor U29934 (N_29934,N_28900,N_28623);
xor U29935 (N_29935,N_28754,N_28396);
nand U29936 (N_29936,N_28577,N_28599);
nand U29937 (N_29937,N_28095,N_28595);
or U29938 (N_29938,N_28394,N_28940);
and U29939 (N_29939,N_28932,N_28262);
nor U29940 (N_29940,N_28255,N_28872);
nand U29941 (N_29941,N_28526,N_28026);
or U29942 (N_29942,N_28090,N_28158);
xnor U29943 (N_29943,N_28433,N_28196);
xor U29944 (N_29944,N_28352,N_28914);
xor U29945 (N_29945,N_28077,N_28053);
nor U29946 (N_29946,N_28866,N_28722);
nand U29947 (N_29947,N_28504,N_28012);
nand U29948 (N_29948,N_28842,N_28893);
nand U29949 (N_29949,N_28211,N_28682);
and U29950 (N_29950,N_28256,N_28394);
and U29951 (N_29951,N_28156,N_28736);
nor U29952 (N_29952,N_28291,N_28685);
and U29953 (N_29953,N_28859,N_28907);
or U29954 (N_29954,N_28381,N_28615);
and U29955 (N_29955,N_28205,N_28249);
or U29956 (N_29956,N_28678,N_28145);
or U29957 (N_29957,N_28451,N_28243);
and U29958 (N_29958,N_28981,N_28274);
and U29959 (N_29959,N_28928,N_28763);
nor U29960 (N_29960,N_28396,N_28410);
or U29961 (N_29961,N_28395,N_28068);
and U29962 (N_29962,N_28377,N_28334);
nand U29963 (N_29963,N_28592,N_28052);
or U29964 (N_29964,N_28598,N_28994);
and U29965 (N_29965,N_28812,N_28216);
and U29966 (N_29966,N_28581,N_28757);
nor U29967 (N_29967,N_28674,N_28481);
nand U29968 (N_29968,N_28047,N_28554);
nor U29969 (N_29969,N_28643,N_28818);
xor U29970 (N_29970,N_28560,N_28093);
xnor U29971 (N_29971,N_28000,N_28938);
nand U29972 (N_29972,N_28556,N_28323);
or U29973 (N_29973,N_28034,N_28470);
or U29974 (N_29974,N_28597,N_28662);
nand U29975 (N_29975,N_28231,N_28640);
or U29976 (N_29976,N_28828,N_28260);
and U29977 (N_29977,N_28579,N_28220);
xnor U29978 (N_29978,N_28207,N_28491);
nand U29979 (N_29979,N_28079,N_28255);
nand U29980 (N_29980,N_28771,N_28070);
xnor U29981 (N_29981,N_28252,N_28363);
or U29982 (N_29982,N_28519,N_28493);
xor U29983 (N_29983,N_28364,N_28587);
and U29984 (N_29984,N_28805,N_28542);
xor U29985 (N_29985,N_28657,N_28347);
xor U29986 (N_29986,N_28006,N_28639);
and U29987 (N_29987,N_28311,N_28849);
or U29988 (N_29988,N_28264,N_28888);
nor U29989 (N_29989,N_28627,N_28076);
nand U29990 (N_29990,N_28503,N_28456);
xnor U29991 (N_29991,N_28913,N_28373);
and U29992 (N_29992,N_28791,N_28559);
and U29993 (N_29993,N_28646,N_28031);
or U29994 (N_29994,N_28793,N_28356);
nand U29995 (N_29995,N_28494,N_28459);
and U29996 (N_29996,N_28931,N_28601);
nand U29997 (N_29997,N_28278,N_28572);
nor U29998 (N_29998,N_28312,N_28923);
xor U29999 (N_29999,N_28023,N_28746);
nand U30000 (N_30000,N_29200,N_29549);
xnor U30001 (N_30001,N_29864,N_29280);
or U30002 (N_30002,N_29868,N_29900);
nand U30003 (N_30003,N_29847,N_29578);
nand U30004 (N_30004,N_29247,N_29621);
and U30005 (N_30005,N_29938,N_29834);
xnor U30006 (N_30006,N_29403,N_29624);
and U30007 (N_30007,N_29581,N_29614);
nand U30008 (N_30008,N_29756,N_29151);
or U30009 (N_30009,N_29187,N_29147);
nor U30010 (N_30010,N_29750,N_29226);
or U30011 (N_30011,N_29925,N_29110);
nand U30012 (N_30012,N_29466,N_29958);
or U30013 (N_30013,N_29781,N_29746);
and U30014 (N_30014,N_29485,N_29617);
nand U30015 (N_30015,N_29168,N_29783);
nand U30016 (N_30016,N_29074,N_29348);
or U30017 (N_30017,N_29383,N_29113);
or U30018 (N_30018,N_29358,N_29611);
nor U30019 (N_30019,N_29917,N_29133);
and U30020 (N_30020,N_29607,N_29608);
nor U30021 (N_30021,N_29311,N_29196);
or U30022 (N_30022,N_29648,N_29653);
nand U30023 (N_30023,N_29237,N_29981);
nor U30024 (N_30024,N_29256,N_29012);
and U30025 (N_30025,N_29803,N_29404);
or U30026 (N_30026,N_29000,N_29270);
xnor U30027 (N_30027,N_29625,N_29907);
nand U30028 (N_30028,N_29165,N_29380);
or U30029 (N_30029,N_29203,N_29456);
nand U30030 (N_30030,N_29856,N_29206);
nor U30031 (N_30031,N_29512,N_29181);
or U30032 (N_30032,N_29792,N_29088);
nand U30033 (N_30033,N_29221,N_29804);
nand U30034 (N_30034,N_29109,N_29100);
nor U30035 (N_30035,N_29170,N_29274);
or U30036 (N_30036,N_29492,N_29169);
xor U30037 (N_30037,N_29889,N_29341);
xor U30038 (N_30038,N_29263,N_29338);
xor U30039 (N_30039,N_29066,N_29812);
and U30040 (N_30040,N_29150,N_29697);
nor U30041 (N_30041,N_29399,N_29437);
nand U30042 (N_30042,N_29733,N_29503);
nor U30043 (N_30043,N_29535,N_29392);
and U30044 (N_30044,N_29236,N_29445);
or U30045 (N_30045,N_29959,N_29789);
nor U30046 (N_30046,N_29896,N_29830);
nor U30047 (N_30047,N_29031,N_29068);
or U30048 (N_30048,N_29590,N_29273);
xor U30049 (N_30049,N_29575,N_29062);
or U30050 (N_30050,N_29351,N_29742);
or U30051 (N_30051,N_29396,N_29817);
nand U30052 (N_30052,N_29172,N_29701);
and U30053 (N_30053,N_29965,N_29442);
xor U30054 (N_30054,N_29252,N_29258);
and U30055 (N_30055,N_29257,N_29866);
xor U30056 (N_30056,N_29239,N_29486);
nand U30057 (N_30057,N_29585,N_29367);
nor U30058 (N_30058,N_29279,N_29217);
or U30059 (N_30059,N_29353,N_29527);
or U30060 (N_30060,N_29121,N_29618);
xnor U30061 (N_30061,N_29390,N_29568);
or U30062 (N_30062,N_29644,N_29725);
and U30063 (N_30063,N_29683,N_29797);
nand U30064 (N_30064,N_29534,N_29550);
or U30065 (N_30065,N_29054,N_29796);
and U30066 (N_30066,N_29173,N_29325);
and U30067 (N_30067,N_29337,N_29028);
or U30068 (N_30068,N_29251,N_29452);
nand U30069 (N_30069,N_29366,N_29061);
nor U30070 (N_30070,N_29176,N_29122);
and U30071 (N_30071,N_29316,N_29954);
or U30072 (N_30072,N_29080,N_29519);
xnor U30073 (N_30073,N_29021,N_29870);
or U30074 (N_30074,N_29881,N_29933);
and U30075 (N_30075,N_29778,N_29670);
and U30076 (N_30076,N_29971,N_29805);
xnor U30077 (N_30077,N_29384,N_29106);
nor U30078 (N_30078,N_29344,N_29587);
or U30079 (N_30079,N_29042,N_29432);
nand U30080 (N_30080,N_29077,N_29631);
and U30081 (N_30081,N_29360,N_29349);
nor U30082 (N_30082,N_29298,N_29598);
nand U30083 (N_30083,N_29167,N_29643);
or U30084 (N_30084,N_29674,N_29924);
nor U30085 (N_30085,N_29030,N_29779);
nor U30086 (N_30086,N_29788,N_29595);
nor U30087 (N_30087,N_29634,N_29820);
or U30088 (N_30088,N_29078,N_29973);
nand U30089 (N_30089,N_29374,N_29695);
or U30090 (N_30090,N_29798,N_29627);
nand U30091 (N_30091,N_29131,N_29141);
xnor U30092 (N_30092,N_29703,N_29580);
nor U30093 (N_30093,N_29806,N_29937);
and U30094 (N_30094,N_29418,N_29497);
nor U30095 (N_30095,N_29057,N_29069);
nand U30096 (N_30096,N_29949,N_29397);
or U30097 (N_30097,N_29424,N_29545);
nor U30098 (N_30098,N_29563,N_29034);
xor U30099 (N_30099,N_29751,N_29458);
xor U30100 (N_30100,N_29795,N_29964);
nand U30101 (N_30101,N_29860,N_29713);
and U30102 (N_30102,N_29556,N_29542);
nand U30103 (N_30103,N_29320,N_29435);
and U30104 (N_30104,N_29330,N_29079);
or U30105 (N_30105,N_29183,N_29092);
nor U30106 (N_30106,N_29350,N_29939);
nand U30107 (N_30107,N_29044,N_29376);
nor U30108 (N_30108,N_29696,N_29738);
xor U30109 (N_30109,N_29036,N_29210);
and U30110 (N_30110,N_29577,N_29240);
xnor U30111 (N_30111,N_29089,N_29479);
or U30112 (N_30112,N_29177,N_29522);
nand U30113 (N_30113,N_29749,N_29554);
or U30114 (N_30114,N_29639,N_29935);
or U30115 (N_30115,N_29129,N_29065);
xnor U30116 (N_30116,N_29365,N_29983);
nand U30117 (N_30117,N_29623,N_29967);
nor U30118 (N_30118,N_29026,N_29205);
nor U30119 (N_30119,N_29553,N_29056);
xnor U30120 (N_30120,N_29543,N_29293);
nand U30121 (N_30121,N_29513,N_29771);
nand U30122 (N_30122,N_29510,N_29102);
xor U30123 (N_30123,N_29120,N_29855);
xnor U30124 (N_30124,N_29601,N_29858);
or U30125 (N_30125,N_29946,N_29451);
nand U30126 (N_30126,N_29304,N_29559);
xor U30127 (N_30127,N_29364,N_29333);
or U30128 (N_30128,N_29869,N_29775);
or U30129 (N_30129,N_29572,N_29963);
nand U30130 (N_30130,N_29667,N_29790);
xor U30131 (N_30131,N_29666,N_29928);
nand U30132 (N_30132,N_29526,N_29671);
nor U30133 (N_30133,N_29905,N_29574);
and U30134 (N_30134,N_29851,N_29888);
nand U30135 (N_30135,N_29076,N_29936);
nor U30136 (N_30136,N_29159,N_29107);
nand U30137 (N_30137,N_29827,N_29516);
and U30138 (N_30138,N_29476,N_29306);
nor U30139 (N_30139,N_29214,N_29943);
nor U30140 (N_30140,N_29053,N_29158);
and U30141 (N_30141,N_29677,N_29768);
nand U30142 (N_30142,N_29986,N_29882);
and U30143 (N_30143,N_29395,N_29067);
nand U30144 (N_30144,N_29430,N_29090);
xor U30145 (N_30145,N_29022,N_29006);
nand U30146 (N_30146,N_29588,N_29813);
xor U30147 (N_30147,N_29539,N_29862);
nor U30148 (N_30148,N_29013,N_29225);
and U30149 (N_30149,N_29615,N_29009);
nor U30150 (N_30150,N_29191,N_29734);
and U30151 (N_30151,N_29676,N_29879);
xnor U30152 (N_30152,N_29363,N_29091);
xnor U30153 (N_30153,N_29582,N_29266);
or U30154 (N_30154,N_29184,N_29331);
nor U30155 (N_30155,N_29471,N_29824);
xor U30156 (N_30156,N_29586,N_29705);
nand U30157 (N_30157,N_29930,N_29199);
nor U30158 (N_30158,N_29767,N_29345);
nor U30159 (N_30159,N_29914,N_29887);
xor U30160 (N_30160,N_29763,N_29468);
or U30161 (N_30161,N_29753,N_29926);
or U30162 (N_30162,N_29413,N_29385);
xor U30163 (N_30163,N_29632,N_29599);
or U30164 (N_30164,N_29499,N_29050);
or U30165 (N_30165,N_29098,N_29823);
xnor U30166 (N_30166,N_29689,N_29748);
xor U30167 (N_30167,N_29142,N_29886);
and U30168 (N_30168,N_29537,N_29831);
nand U30169 (N_30169,N_29224,N_29629);
xnor U30170 (N_30170,N_29319,N_29443);
and U30171 (N_30171,N_29517,N_29362);
nand U30172 (N_30172,N_29058,N_29863);
nor U30173 (N_30173,N_29455,N_29420);
or U30174 (N_30174,N_29276,N_29112);
xnor U30175 (N_30175,N_29460,N_29202);
nor U30176 (N_30176,N_29139,N_29436);
nor U30177 (N_30177,N_29470,N_29988);
nor U30178 (N_30178,N_29248,N_29439);
xnor U30179 (N_30179,N_29229,N_29425);
nand U30180 (N_30180,N_29950,N_29394);
xnor U30181 (N_30181,N_29897,N_29381);
nor U30182 (N_30182,N_29194,N_29682);
xor U30183 (N_30183,N_29149,N_29814);
and U30184 (N_30184,N_29464,N_29228);
nor U30185 (N_30185,N_29271,N_29246);
xor U30186 (N_30186,N_29315,N_29844);
or U30187 (N_30187,N_29650,N_29669);
xnor U30188 (N_30188,N_29387,N_29945);
nor U30189 (N_30189,N_29509,N_29893);
or U30190 (N_30190,N_29832,N_29357);
nand U30191 (N_30191,N_29125,N_29429);
nand U30192 (N_30192,N_29233,N_29745);
nand U30193 (N_30193,N_29114,N_29651);
xor U30194 (N_30194,N_29604,N_29083);
nor U30195 (N_30195,N_29547,N_29462);
or U30196 (N_30196,N_29828,N_29721);
nand U30197 (N_30197,N_29340,N_29772);
nand U30198 (N_30198,N_29454,N_29402);
or U30199 (N_30199,N_29810,N_29219);
nand U30200 (N_30200,N_29448,N_29087);
and U30201 (N_30201,N_29691,N_29504);
or U30202 (N_30202,N_29453,N_29017);
nor U30203 (N_30203,N_29447,N_29567);
or U30204 (N_30204,N_29037,N_29528);
and U30205 (N_30205,N_29638,N_29867);
nand U30206 (N_30206,N_29175,N_29536);
nand U30207 (N_30207,N_29794,N_29999);
nor U30208 (N_30208,N_29530,N_29377);
nand U30209 (N_30209,N_29154,N_29010);
xor U30210 (N_30210,N_29081,N_29564);
or U30211 (N_30211,N_29446,N_29487);
xnor U30212 (N_30212,N_29693,N_29164);
nor U30213 (N_30213,N_29819,N_29603);
nand U30214 (N_30214,N_29871,N_29473);
and U30215 (N_30215,N_29300,N_29321);
xor U30216 (N_30216,N_29195,N_29941);
nand U30217 (N_30217,N_29305,N_29412);
xor U30218 (N_30218,N_29663,N_29123);
or U30219 (N_30219,N_29033,N_29301);
xnor U30220 (N_30220,N_29619,N_29722);
nand U30221 (N_30221,N_29138,N_29609);
xor U30222 (N_30222,N_29576,N_29329);
and U30223 (N_30223,N_29208,N_29494);
nor U30224 (N_30224,N_29808,N_29980);
nand U30225 (N_30225,N_29726,N_29754);
and U30226 (N_30226,N_29524,N_29207);
xnor U30227 (N_30227,N_29014,N_29414);
or U30228 (N_30228,N_29288,N_29681);
xor U30229 (N_30229,N_29264,N_29096);
nor U30230 (N_30230,N_29500,N_29707);
nor U30231 (N_30231,N_29143,N_29406);
xnor U30232 (N_30232,N_29440,N_29277);
and U30233 (N_30233,N_29923,N_29729);
nand U30234 (N_30234,N_29839,N_29188);
nand U30235 (N_30235,N_29531,N_29894);
or U30236 (N_30236,N_29211,N_29773);
nor U30237 (N_30237,N_29525,N_29444);
nand U30238 (N_30238,N_29148,N_29920);
nand U30239 (N_30239,N_29190,N_29613);
nor U30240 (N_30240,N_29163,N_29557);
or U30241 (N_30241,N_29498,N_29902);
or U30242 (N_30242,N_29060,N_29269);
xor U30243 (N_30243,N_29708,N_29180);
xnor U30244 (N_30244,N_29714,N_29511);
xnor U30245 (N_30245,N_29242,N_29835);
or U30246 (N_30246,N_29178,N_29032);
and U30247 (N_30247,N_29640,N_29731);
or U30248 (N_30248,N_29339,N_29898);
nor U30249 (N_30249,N_29047,N_29658);
nand U30250 (N_30250,N_29777,N_29343);
or U30251 (N_30251,N_29649,N_29704);
and U30252 (N_30252,N_29244,N_29475);
nor U30253 (N_30253,N_29019,N_29997);
and U30254 (N_30254,N_29850,N_29282);
xnor U30255 (N_30255,N_29405,N_29326);
nor U30256 (N_30256,N_29063,N_29185);
or U30257 (N_30257,N_29502,N_29630);
xnor U30258 (N_30258,N_29477,N_29840);
and U30259 (N_30259,N_29985,N_29160);
nor U30260 (N_30260,N_29720,N_29884);
nor U30261 (N_30261,N_29490,N_29463);
nand U30262 (N_30262,N_29822,N_29931);
nand U30263 (N_30263,N_29117,N_29426);
or U30264 (N_30264,N_29375,N_29140);
and U30265 (N_30265,N_29904,N_29097);
nor U30266 (N_30266,N_29153,N_29489);
or U30267 (N_30267,N_29419,N_29807);
nand U30268 (N_30268,N_29307,N_29231);
nor U30269 (N_30269,N_29015,N_29232);
and U30270 (N_30270,N_29961,N_29126);
and U30271 (N_30271,N_29571,N_29346);
or U30272 (N_30272,N_29286,N_29059);
and U30273 (N_30273,N_29791,N_29438);
xor U30274 (N_30274,N_29927,N_29987);
xnor U30275 (N_30275,N_29921,N_29001);
nor U30276 (N_30276,N_29467,N_29314);
or U30277 (N_30277,N_29686,N_29801);
and U30278 (N_30278,N_29323,N_29417);
xnor U30279 (N_30279,N_29991,N_29659);
and U30280 (N_30280,N_29312,N_29996);
nand U30281 (N_30281,N_29873,N_29260);
or U30282 (N_30282,N_29755,N_29786);
or U30283 (N_30283,N_29739,N_29952);
and U30284 (N_30284,N_29508,N_29876);
nand U30285 (N_30285,N_29837,N_29968);
or U30286 (N_30286,N_29825,N_29573);
nand U30287 (N_30287,N_29128,N_29660);
nand U30288 (N_30288,N_29171,N_29646);
nor U30289 (N_30289,N_29597,N_29398);
xnor U30290 (N_30290,N_29035,N_29235);
nand U30291 (N_30291,N_29433,N_29787);
xor U30292 (N_30292,N_29241,N_29785);
and U30293 (N_30293,N_29506,N_29386);
nor U30294 (N_30294,N_29647,N_29685);
nor U30295 (N_30295,N_29024,N_29197);
nor U30296 (N_30296,N_29723,N_29025);
or U30297 (N_30297,N_29043,N_29268);
and U30298 (N_30298,N_29626,N_29027);
nand U30299 (N_30299,N_29679,N_29583);
and U30300 (N_30300,N_29372,N_29724);
xnor U30301 (N_30301,N_29474,N_29029);
nand U30302 (N_30302,N_29654,N_29193);
nor U30303 (N_30303,N_29491,N_29267);
or U30304 (N_30304,N_29551,N_29234);
or U30305 (N_30305,N_29570,N_29003);
xor U30306 (N_30306,N_29422,N_29322);
and U30307 (N_30307,N_29799,N_29673);
xnor U30308 (N_30308,N_29484,N_29774);
nor U30309 (N_30309,N_29605,N_29152);
and U30310 (N_30310,N_29505,N_29145);
nor U30311 (N_30311,N_29101,N_29428);
or U30312 (N_30312,N_29073,N_29070);
and U30313 (N_30313,N_29262,N_29736);
and U30314 (N_30314,N_29094,N_29566);
and U30315 (N_30315,N_29974,N_29932);
nand U30316 (N_30316,N_29633,N_29761);
nand U30317 (N_30317,N_29480,N_29045);
or U30318 (N_30318,N_29493,N_29661);
or U30319 (N_30319,N_29995,N_29481);
and U30320 (N_30320,N_29303,N_29916);
nor U30321 (N_30321,N_29055,N_29238);
xor U30322 (N_30322,N_29912,N_29104);
or U30323 (N_30323,N_29132,N_29410);
xnor U30324 (N_30324,N_29600,N_29878);
and U30325 (N_30325,N_29711,N_29023);
xor U30326 (N_30326,N_29816,N_29018);
or U30327 (N_30327,N_29728,N_29833);
nand U30328 (N_30328,N_29741,N_29488);
and U30329 (N_30329,N_29483,N_29215);
xor U30330 (N_30330,N_29213,N_29334);
or U30331 (N_30331,N_29953,N_29982);
or U30332 (N_30332,N_29540,N_29296);
and U30333 (N_30333,N_29718,N_29877);
or U30334 (N_30334,N_29450,N_29085);
nand U30335 (N_30335,N_29423,N_29890);
nor U30336 (N_30336,N_29622,N_29415);
or U30337 (N_30337,N_29901,N_29845);
nand U30338 (N_30338,N_29284,N_29292);
and U30339 (N_30339,N_29811,N_29218);
or U30340 (N_30340,N_29944,N_29969);
xnor U30341 (N_30341,N_29727,N_29616);
nor U30342 (N_30342,N_29368,N_29291);
nor U30343 (N_30343,N_29780,N_29678);
nand U30344 (N_30344,N_29116,N_29389);
or U30345 (N_30345,N_29465,N_29198);
nor U30346 (N_30346,N_29099,N_29883);
nor U30347 (N_30347,N_29735,N_29544);
xor U30348 (N_30348,N_29161,N_29408);
nand U30349 (N_30349,N_29716,N_29702);
nand U30350 (N_30350,N_29523,N_29836);
nand U30351 (N_30351,N_29308,N_29719);
nor U30352 (N_30352,N_29243,N_29744);
and U30353 (N_30353,N_29361,N_29230);
or U30354 (N_30354,N_29495,N_29310);
and U30355 (N_30355,N_29960,N_29119);
and U30356 (N_30356,N_29457,N_29355);
nand U30357 (N_30357,N_29684,N_29594);
nand U30358 (N_30358,N_29335,N_29918);
and U30359 (N_30359,N_29086,N_29776);
nand U30360 (N_30360,N_29265,N_29136);
nor U30361 (N_30361,N_29212,N_29668);
or U30362 (N_30362,N_29715,N_29815);
or U30363 (N_30363,N_29977,N_29400);
and U30364 (N_30364,N_29124,N_29910);
or U30365 (N_30365,N_29108,N_29848);
nand U30366 (N_30366,N_29514,N_29911);
or U30367 (N_30367,N_29710,N_29990);
xnor U30368 (N_30368,N_29072,N_29765);
or U30369 (N_30369,N_29093,N_29838);
nand U30370 (N_30370,N_29302,N_29318);
xnor U30371 (N_30371,N_29299,N_29294);
nand U30372 (N_30372,N_29008,N_29421);
or U30373 (N_30373,N_29039,N_29747);
or U30374 (N_30374,N_29717,N_29692);
xor U30375 (N_30375,N_29352,N_29758);
and U30376 (N_30376,N_29743,N_29347);
and U30377 (N_30377,N_29324,N_29281);
nand U30378 (N_30378,N_29841,N_29254);
xnor U30379 (N_30379,N_29144,N_29818);
nor U30380 (N_30380,N_29706,N_29223);
or U30381 (N_30381,N_29642,N_29111);
and U30382 (N_30382,N_29427,N_29441);
xor U30383 (N_30383,N_29853,N_29259);
and U30384 (N_30384,N_29913,N_29994);
xor U30385 (N_30385,N_29051,N_29700);
or U30386 (N_30386,N_29075,N_29955);
or U30387 (N_30387,N_29843,N_29411);
nor U30388 (N_30388,N_29662,N_29478);
or U30389 (N_30389,N_29992,N_29784);
xor U30390 (N_30390,N_29407,N_29846);
nand U30391 (N_30391,N_29041,N_29665);
or U30392 (N_30392,N_29285,N_29645);
xor U30393 (N_30393,N_29589,N_29993);
nand U30394 (N_30394,N_29250,N_29546);
or U30395 (N_30395,N_29975,N_29371);
nor U30396 (N_30396,N_29602,N_29095);
and U30397 (N_30397,N_29103,N_29760);
or U30398 (N_30398,N_29998,N_29929);
xnor U30399 (N_30399,N_29687,N_29127);
or U30400 (N_30400,N_29875,N_29675);
xor U30401 (N_30401,N_29762,N_29272);
nand U30402 (N_30402,N_29852,N_29857);
nor U30403 (N_30403,N_29354,N_29680);
and U30404 (N_30404,N_29874,N_29189);
nor U30405 (N_30405,N_29956,N_29222);
and U30406 (N_30406,N_29652,N_29628);
xor U30407 (N_30407,N_29606,N_29694);
and U30408 (N_30408,N_29209,N_29934);
or U30409 (N_30409,N_29737,N_29664);
nor U30410 (N_30410,N_29962,N_29501);
nor U30411 (N_30411,N_29712,N_29290);
or U30412 (N_30412,N_29038,N_29431);
xnor U30413 (N_30413,N_29885,N_29002);
or U30414 (N_30414,N_29186,N_29984);
and U30415 (N_30415,N_29472,N_29569);
xor U30416 (N_30416,N_29393,N_29596);
xnor U30417 (N_30417,N_29249,N_29891);
nor U30418 (N_30418,N_29579,N_29793);
and U30419 (N_30419,N_29192,N_29922);
nand U30420 (N_30420,N_29007,N_29555);
nor U30421 (N_30421,N_29903,N_29016);
or U30422 (N_30422,N_29561,N_29872);
nor U30423 (N_30423,N_29182,N_29156);
nand U30424 (N_30424,N_29533,N_29227);
xnor U30425 (N_30425,N_29204,N_29565);
or U30426 (N_30426,N_29854,N_29434);
and U30427 (N_30427,N_29507,N_29809);
nand U30428 (N_30428,N_29688,N_29255);
xnor U30429 (N_30429,N_29261,N_29620);
and U30430 (N_30430,N_29155,N_29105);
nor U30431 (N_30431,N_29342,N_29558);
nand U30432 (N_30432,N_29461,N_29880);
nor U30433 (N_30433,N_29378,N_29842);
and U30434 (N_30434,N_29637,N_29730);
xnor U30435 (N_30435,N_29040,N_29915);
xnor U30436 (N_30436,N_29297,N_29005);
xnor U30437 (N_30437,N_29740,N_29782);
nand U30438 (N_30438,N_29336,N_29826);
xnor U30439 (N_30439,N_29541,N_29942);
and U30440 (N_30440,N_29560,N_29048);
and U30441 (N_30441,N_29115,N_29940);
and U30442 (N_30442,N_29289,N_29989);
and U30443 (N_30443,N_29657,N_29591);
and U30444 (N_30444,N_29859,N_29947);
and U30445 (N_30445,N_29592,N_29449);
nor U30446 (N_30446,N_29179,N_29709);
xor U30447 (N_30447,N_29909,N_29220);
nand U30448 (N_30448,N_29908,N_29895);
and U30449 (N_30449,N_29166,N_29593);
or U30450 (N_30450,N_29972,N_29532);
nor U30451 (N_30451,N_29146,N_29802);
or U30452 (N_30452,N_29275,N_29071);
xnor U30453 (N_30453,N_29979,N_29957);
and U30454 (N_30454,N_29732,N_29636);
and U30455 (N_30455,N_29518,N_29548);
and U30456 (N_30456,N_29552,N_29004);
xnor U30457 (N_30457,N_29201,N_29174);
nand U30458 (N_30458,N_29356,N_29137);
or U30459 (N_30459,N_29052,N_29295);
nor U30460 (N_30460,N_29388,N_29082);
or U30461 (N_30461,N_29157,N_29752);
or U30462 (N_30462,N_29401,N_29278);
xor U30463 (N_30463,N_29892,N_29562);
and U30464 (N_30464,N_29245,N_29757);
nand U30465 (N_30465,N_29970,N_29369);
or U30466 (N_30466,N_29469,N_29359);
nor U30467 (N_30467,N_29821,N_29635);
nand U30468 (N_30468,N_29610,N_29865);
and U30469 (N_30469,N_29416,N_29655);
xnor U30470 (N_30470,N_29515,N_29584);
nor U30471 (N_30471,N_29049,N_29978);
xor U30472 (N_30472,N_29287,N_29118);
and U30473 (N_30473,N_29084,N_29672);
or U30474 (N_30474,N_29134,N_29332);
nor U30475 (N_30475,N_29011,N_29759);
nor U30476 (N_30476,N_29764,N_29919);
nor U30477 (N_30477,N_29313,N_29861);
and U30478 (N_30478,N_29064,N_29328);
or U30479 (N_30479,N_29976,N_29899);
or U30480 (N_30480,N_29130,N_29496);
nor U30481 (N_30481,N_29046,N_29379);
nor U30482 (N_30482,N_29690,N_29391);
xnor U30483 (N_30483,N_29253,N_29766);
or U30484 (N_30484,N_29906,N_29459);
or U30485 (N_30485,N_29309,N_29966);
or U30486 (N_30486,N_29162,N_29656);
xor U30487 (N_30487,N_29382,N_29698);
xor U30488 (N_30488,N_29699,N_29135);
or U30489 (N_30489,N_29770,N_29849);
and U30490 (N_30490,N_29216,N_29521);
xor U30491 (N_30491,N_29529,N_29373);
or U30492 (N_30492,N_29948,N_29538);
nand U30493 (N_30493,N_29520,N_29020);
and U30494 (N_30494,N_29800,N_29283);
xnor U30495 (N_30495,N_29370,N_29409);
or U30496 (N_30496,N_29641,N_29829);
and U30497 (N_30497,N_29482,N_29612);
nand U30498 (N_30498,N_29317,N_29951);
nand U30499 (N_30499,N_29327,N_29769);
and U30500 (N_30500,N_29483,N_29092);
nor U30501 (N_30501,N_29168,N_29488);
nor U30502 (N_30502,N_29566,N_29125);
or U30503 (N_30503,N_29262,N_29743);
nand U30504 (N_30504,N_29010,N_29030);
or U30505 (N_30505,N_29346,N_29932);
xnor U30506 (N_30506,N_29340,N_29567);
and U30507 (N_30507,N_29771,N_29222);
nand U30508 (N_30508,N_29322,N_29516);
and U30509 (N_30509,N_29992,N_29859);
and U30510 (N_30510,N_29470,N_29823);
nor U30511 (N_30511,N_29306,N_29104);
or U30512 (N_30512,N_29674,N_29271);
nor U30513 (N_30513,N_29565,N_29558);
nor U30514 (N_30514,N_29060,N_29251);
or U30515 (N_30515,N_29304,N_29663);
or U30516 (N_30516,N_29104,N_29363);
nand U30517 (N_30517,N_29766,N_29014);
and U30518 (N_30518,N_29045,N_29293);
and U30519 (N_30519,N_29076,N_29456);
nor U30520 (N_30520,N_29444,N_29114);
nand U30521 (N_30521,N_29156,N_29967);
nor U30522 (N_30522,N_29154,N_29529);
xor U30523 (N_30523,N_29272,N_29202);
nor U30524 (N_30524,N_29708,N_29363);
or U30525 (N_30525,N_29680,N_29002);
and U30526 (N_30526,N_29063,N_29652);
nor U30527 (N_30527,N_29537,N_29826);
or U30528 (N_30528,N_29683,N_29721);
nor U30529 (N_30529,N_29180,N_29114);
or U30530 (N_30530,N_29723,N_29130);
xor U30531 (N_30531,N_29631,N_29023);
nor U30532 (N_30532,N_29130,N_29465);
and U30533 (N_30533,N_29495,N_29359);
or U30534 (N_30534,N_29467,N_29685);
nor U30535 (N_30535,N_29147,N_29750);
xnor U30536 (N_30536,N_29652,N_29617);
nand U30537 (N_30537,N_29091,N_29241);
or U30538 (N_30538,N_29202,N_29967);
nor U30539 (N_30539,N_29992,N_29915);
nor U30540 (N_30540,N_29315,N_29656);
and U30541 (N_30541,N_29479,N_29388);
and U30542 (N_30542,N_29727,N_29136);
xor U30543 (N_30543,N_29089,N_29881);
or U30544 (N_30544,N_29745,N_29285);
or U30545 (N_30545,N_29089,N_29700);
nand U30546 (N_30546,N_29687,N_29505);
xor U30547 (N_30547,N_29470,N_29615);
nand U30548 (N_30548,N_29552,N_29587);
xor U30549 (N_30549,N_29647,N_29691);
nand U30550 (N_30550,N_29863,N_29251);
and U30551 (N_30551,N_29352,N_29785);
xnor U30552 (N_30552,N_29715,N_29939);
or U30553 (N_30553,N_29614,N_29999);
nor U30554 (N_30554,N_29782,N_29242);
nor U30555 (N_30555,N_29797,N_29082);
nor U30556 (N_30556,N_29942,N_29892);
nor U30557 (N_30557,N_29237,N_29085);
xnor U30558 (N_30558,N_29784,N_29361);
and U30559 (N_30559,N_29378,N_29535);
nand U30560 (N_30560,N_29664,N_29103);
nor U30561 (N_30561,N_29354,N_29558);
nand U30562 (N_30562,N_29691,N_29417);
xor U30563 (N_30563,N_29808,N_29736);
nor U30564 (N_30564,N_29140,N_29986);
and U30565 (N_30565,N_29670,N_29285);
nor U30566 (N_30566,N_29964,N_29511);
nand U30567 (N_30567,N_29070,N_29092);
nand U30568 (N_30568,N_29600,N_29862);
nand U30569 (N_30569,N_29231,N_29561);
and U30570 (N_30570,N_29645,N_29196);
nor U30571 (N_30571,N_29017,N_29623);
or U30572 (N_30572,N_29545,N_29681);
nand U30573 (N_30573,N_29074,N_29207);
xor U30574 (N_30574,N_29364,N_29888);
nand U30575 (N_30575,N_29396,N_29154);
xor U30576 (N_30576,N_29652,N_29479);
nand U30577 (N_30577,N_29597,N_29977);
nor U30578 (N_30578,N_29620,N_29099);
nand U30579 (N_30579,N_29118,N_29336);
or U30580 (N_30580,N_29683,N_29604);
xor U30581 (N_30581,N_29058,N_29100);
xnor U30582 (N_30582,N_29258,N_29949);
or U30583 (N_30583,N_29252,N_29617);
nor U30584 (N_30584,N_29389,N_29266);
nand U30585 (N_30585,N_29824,N_29680);
or U30586 (N_30586,N_29722,N_29100);
xor U30587 (N_30587,N_29174,N_29415);
nor U30588 (N_30588,N_29999,N_29492);
and U30589 (N_30589,N_29754,N_29257);
xor U30590 (N_30590,N_29203,N_29586);
and U30591 (N_30591,N_29551,N_29970);
nor U30592 (N_30592,N_29337,N_29022);
or U30593 (N_30593,N_29333,N_29780);
xor U30594 (N_30594,N_29107,N_29992);
nand U30595 (N_30595,N_29588,N_29966);
nand U30596 (N_30596,N_29730,N_29409);
nor U30597 (N_30597,N_29360,N_29845);
and U30598 (N_30598,N_29801,N_29544);
xor U30599 (N_30599,N_29172,N_29489);
xnor U30600 (N_30600,N_29753,N_29316);
or U30601 (N_30601,N_29342,N_29545);
xnor U30602 (N_30602,N_29699,N_29140);
xnor U30603 (N_30603,N_29565,N_29574);
or U30604 (N_30604,N_29454,N_29437);
or U30605 (N_30605,N_29512,N_29432);
or U30606 (N_30606,N_29571,N_29990);
or U30607 (N_30607,N_29533,N_29342);
nor U30608 (N_30608,N_29382,N_29681);
or U30609 (N_30609,N_29714,N_29113);
nand U30610 (N_30610,N_29412,N_29775);
nor U30611 (N_30611,N_29198,N_29985);
or U30612 (N_30612,N_29379,N_29761);
and U30613 (N_30613,N_29437,N_29894);
nor U30614 (N_30614,N_29793,N_29741);
or U30615 (N_30615,N_29936,N_29345);
and U30616 (N_30616,N_29195,N_29762);
nand U30617 (N_30617,N_29505,N_29246);
nand U30618 (N_30618,N_29592,N_29350);
nand U30619 (N_30619,N_29423,N_29789);
or U30620 (N_30620,N_29594,N_29295);
and U30621 (N_30621,N_29044,N_29251);
nand U30622 (N_30622,N_29859,N_29789);
nand U30623 (N_30623,N_29930,N_29047);
nor U30624 (N_30624,N_29529,N_29073);
nand U30625 (N_30625,N_29095,N_29824);
nand U30626 (N_30626,N_29742,N_29382);
nand U30627 (N_30627,N_29745,N_29848);
nor U30628 (N_30628,N_29601,N_29467);
xor U30629 (N_30629,N_29293,N_29624);
nand U30630 (N_30630,N_29647,N_29018);
and U30631 (N_30631,N_29518,N_29294);
nand U30632 (N_30632,N_29735,N_29409);
or U30633 (N_30633,N_29512,N_29963);
nand U30634 (N_30634,N_29333,N_29313);
xor U30635 (N_30635,N_29559,N_29780);
nand U30636 (N_30636,N_29117,N_29554);
or U30637 (N_30637,N_29913,N_29583);
or U30638 (N_30638,N_29423,N_29576);
nand U30639 (N_30639,N_29939,N_29447);
and U30640 (N_30640,N_29490,N_29749);
xnor U30641 (N_30641,N_29033,N_29724);
xnor U30642 (N_30642,N_29483,N_29054);
or U30643 (N_30643,N_29331,N_29840);
xor U30644 (N_30644,N_29867,N_29903);
and U30645 (N_30645,N_29559,N_29775);
or U30646 (N_30646,N_29085,N_29781);
nand U30647 (N_30647,N_29446,N_29330);
nand U30648 (N_30648,N_29897,N_29811);
xor U30649 (N_30649,N_29219,N_29001);
nand U30650 (N_30650,N_29292,N_29286);
xnor U30651 (N_30651,N_29797,N_29580);
nor U30652 (N_30652,N_29751,N_29677);
xor U30653 (N_30653,N_29747,N_29559);
xor U30654 (N_30654,N_29099,N_29019);
and U30655 (N_30655,N_29712,N_29730);
xnor U30656 (N_30656,N_29247,N_29948);
and U30657 (N_30657,N_29143,N_29820);
nand U30658 (N_30658,N_29058,N_29536);
or U30659 (N_30659,N_29515,N_29765);
nor U30660 (N_30660,N_29104,N_29399);
or U30661 (N_30661,N_29607,N_29480);
or U30662 (N_30662,N_29157,N_29102);
xor U30663 (N_30663,N_29008,N_29844);
or U30664 (N_30664,N_29098,N_29721);
nor U30665 (N_30665,N_29774,N_29216);
xor U30666 (N_30666,N_29104,N_29461);
nor U30667 (N_30667,N_29583,N_29093);
nor U30668 (N_30668,N_29793,N_29035);
nand U30669 (N_30669,N_29779,N_29941);
or U30670 (N_30670,N_29130,N_29266);
nor U30671 (N_30671,N_29770,N_29476);
and U30672 (N_30672,N_29888,N_29713);
or U30673 (N_30673,N_29150,N_29005);
or U30674 (N_30674,N_29174,N_29336);
nor U30675 (N_30675,N_29541,N_29787);
or U30676 (N_30676,N_29348,N_29772);
and U30677 (N_30677,N_29647,N_29851);
and U30678 (N_30678,N_29054,N_29662);
and U30679 (N_30679,N_29444,N_29766);
nor U30680 (N_30680,N_29001,N_29316);
nor U30681 (N_30681,N_29324,N_29949);
and U30682 (N_30682,N_29102,N_29350);
nand U30683 (N_30683,N_29288,N_29262);
nand U30684 (N_30684,N_29513,N_29070);
nor U30685 (N_30685,N_29380,N_29512);
nor U30686 (N_30686,N_29153,N_29313);
and U30687 (N_30687,N_29770,N_29653);
and U30688 (N_30688,N_29245,N_29917);
nand U30689 (N_30689,N_29506,N_29990);
xor U30690 (N_30690,N_29083,N_29090);
xor U30691 (N_30691,N_29474,N_29228);
nor U30692 (N_30692,N_29040,N_29324);
and U30693 (N_30693,N_29054,N_29500);
or U30694 (N_30694,N_29582,N_29866);
or U30695 (N_30695,N_29968,N_29657);
or U30696 (N_30696,N_29007,N_29692);
and U30697 (N_30697,N_29090,N_29477);
nor U30698 (N_30698,N_29556,N_29951);
and U30699 (N_30699,N_29872,N_29869);
xnor U30700 (N_30700,N_29966,N_29094);
nor U30701 (N_30701,N_29162,N_29181);
and U30702 (N_30702,N_29384,N_29881);
and U30703 (N_30703,N_29700,N_29837);
or U30704 (N_30704,N_29091,N_29320);
or U30705 (N_30705,N_29313,N_29890);
and U30706 (N_30706,N_29948,N_29041);
nor U30707 (N_30707,N_29957,N_29442);
or U30708 (N_30708,N_29120,N_29797);
xor U30709 (N_30709,N_29195,N_29444);
or U30710 (N_30710,N_29561,N_29269);
nand U30711 (N_30711,N_29009,N_29397);
nand U30712 (N_30712,N_29236,N_29428);
and U30713 (N_30713,N_29375,N_29931);
xor U30714 (N_30714,N_29635,N_29005);
xnor U30715 (N_30715,N_29575,N_29167);
or U30716 (N_30716,N_29384,N_29267);
nand U30717 (N_30717,N_29238,N_29278);
or U30718 (N_30718,N_29091,N_29235);
and U30719 (N_30719,N_29455,N_29654);
and U30720 (N_30720,N_29521,N_29898);
or U30721 (N_30721,N_29602,N_29003);
or U30722 (N_30722,N_29846,N_29275);
or U30723 (N_30723,N_29509,N_29857);
xnor U30724 (N_30724,N_29022,N_29490);
or U30725 (N_30725,N_29509,N_29412);
xnor U30726 (N_30726,N_29917,N_29593);
xnor U30727 (N_30727,N_29979,N_29755);
or U30728 (N_30728,N_29590,N_29419);
and U30729 (N_30729,N_29502,N_29147);
or U30730 (N_30730,N_29439,N_29010);
or U30731 (N_30731,N_29499,N_29092);
nand U30732 (N_30732,N_29483,N_29912);
nor U30733 (N_30733,N_29173,N_29780);
nor U30734 (N_30734,N_29650,N_29617);
nand U30735 (N_30735,N_29592,N_29830);
or U30736 (N_30736,N_29147,N_29703);
and U30737 (N_30737,N_29486,N_29359);
and U30738 (N_30738,N_29708,N_29512);
nor U30739 (N_30739,N_29553,N_29937);
xnor U30740 (N_30740,N_29658,N_29746);
nor U30741 (N_30741,N_29962,N_29640);
nand U30742 (N_30742,N_29746,N_29935);
or U30743 (N_30743,N_29836,N_29387);
xnor U30744 (N_30744,N_29898,N_29824);
and U30745 (N_30745,N_29600,N_29340);
and U30746 (N_30746,N_29714,N_29003);
xor U30747 (N_30747,N_29169,N_29637);
nand U30748 (N_30748,N_29751,N_29933);
nand U30749 (N_30749,N_29560,N_29106);
xor U30750 (N_30750,N_29428,N_29811);
xnor U30751 (N_30751,N_29668,N_29333);
and U30752 (N_30752,N_29030,N_29948);
nor U30753 (N_30753,N_29932,N_29830);
nand U30754 (N_30754,N_29538,N_29779);
and U30755 (N_30755,N_29621,N_29003);
xnor U30756 (N_30756,N_29844,N_29098);
and U30757 (N_30757,N_29410,N_29175);
nand U30758 (N_30758,N_29767,N_29144);
nor U30759 (N_30759,N_29633,N_29965);
or U30760 (N_30760,N_29612,N_29585);
nor U30761 (N_30761,N_29058,N_29213);
nand U30762 (N_30762,N_29322,N_29597);
xor U30763 (N_30763,N_29578,N_29905);
nand U30764 (N_30764,N_29099,N_29578);
xnor U30765 (N_30765,N_29469,N_29763);
nand U30766 (N_30766,N_29600,N_29341);
nor U30767 (N_30767,N_29645,N_29272);
nand U30768 (N_30768,N_29411,N_29522);
nor U30769 (N_30769,N_29985,N_29015);
xnor U30770 (N_30770,N_29702,N_29288);
nor U30771 (N_30771,N_29216,N_29058);
or U30772 (N_30772,N_29667,N_29976);
xnor U30773 (N_30773,N_29810,N_29639);
xor U30774 (N_30774,N_29870,N_29845);
or U30775 (N_30775,N_29026,N_29946);
nand U30776 (N_30776,N_29578,N_29171);
and U30777 (N_30777,N_29080,N_29760);
and U30778 (N_30778,N_29561,N_29556);
or U30779 (N_30779,N_29994,N_29103);
nor U30780 (N_30780,N_29980,N_29527);
or U30781 (N_30781,N_29884,N_29219);
or U30782 (N_30782,N_29838,N_29027);
nand U30783 (N_30783,N_29026,N_29255);
nor U30784 (N_30784,N_29977,N_29386);
nor U30785 (N_30785,N_29686,N_29984);
and U30786 (N_30786,N_29600,N_29779);
or U30787 (N_30787,N_29171,N_29148);
nor U30788 (N_30788,N_29856,N_29547);
or U30789 (N_30789,N_29869,N_29603);
and U30790 (N_30790,N_29935,N_29420);
xnor U30791 (N_30791,N_29729,N_29465);
or U30792 (N_30792,N_29753,N_29632);
xor U30793 (N_30793,N_29128,N_29775);
or U30794 (N_30794,N_29364,N_29938);
nand U30795 (N_30795,N_29210,N_29193);
xnor U30796 (N_30796,N_29933,N_29662);
or U30797 (N_30797,N_29511,N_29853);
nand U30798 (N_30798,N_29514,N_29402);
nor U30799 (N_30799,N_29261,N_29636);
and U30800 (N_30800,N_29134,N_29718);
nand U30801 (N_30801,N_29265,N_29976);
nor U30802 (N_30802,N_29618,N_29683);
and U30803 (N_30803,N_29560,N_29097);
xor U30804 (N_30804,N_29855,N_29898);
or U30805 (N_30805,N_29241,N_29781);
nand U30806 (N_30806,N_29482,N_29886);
and U30807 (N_30807,N_29512,N_29937);
or U30808 (N_30808,N_29857,N_29314);
nor U30809 (N_30809,N_29967,N_29764);
and U30810 (N_30810,N_29883,N_29125);
nor U30811 (N_30811,N_29323,N_29120);
and U30812 (N_30812,N_29744,N_29469);
nor U30813 (N_30813,N_29465,N_29479);
and U30814 (N_30814,N_29954,N_29646);
and U30815 (N_30815,N_29624,N_29743);
nor U30816 (N_30816,N_29857,N_29883);
xnor U30817 (N_30817,N_29575,N_29550);
nand U30818 (N_30818,N_29848,N_29385);
xor U30819 (N_30819,N_29730,N_29771);
nor U30820 (N_30820,N_29237,N_29141);
nor U30821 (N_30821,N_29421,N_29884);
nor U30822 (N_30822,N_29277,N_29725);
and U30823 (N_30823,N_29987,N_29235);
xor U30824 (N_30824,N_29080,N_29280);
and U30825 (N_30825,N_29979,N_29678);
or U30826 (N_30826,N_29883,N_29426);
nor U30827 (N_30827,N_29247,N_29039);
and U30828 (N_30828,N_29111,N_29837);
and U30829 (N_30829,N_29768,N_29354);
nor U30830 (N_30830,N_29838,N_29090);
or U30831 (N_30831,N_29502,N_29871);
nand U30832 (N_30832,N_29573,N_29810);
or U30833 (N_30833,N_29608,N_29528);
nand U30834 (N_30834,N_29033,N_29266);
and U30835 (N_30835,N_29104,N_29706);
nand U30836 (N_30836,N_29398,N_29567);
nor U30837 (N_30837,N_29988,N_29208);
xor U30838 (N_30838,N_29378,N_29271);
and U30839 (N_30839,N_29825,N_29941);
or U30840 (N_30840,N_29073,N_29105);
xnor U30841 (N_30841,N_29329,N_29347);
nor U30842 (N_30842,N_29666,N_29844);
xor U30843 (N_30843,N_29551,N_29788);
nand U30844 (N_30844,N_29943,N_29099);
and U30845 (N_30845,N_29960,N_29537);
xor U30846 (N_30846,N_29626,N_29741);
xnor U30847 (N_30847,N_29637,N_29093);
xor U30848 (N_30848,N_29836,N_29493);
xnor U30849 (N_30849,N_29317,N_29205);
nand U30850 (N_30850,N_29152,N_29398);
or U30851 (N_30851,N_29120,N_29960);
and U30852 (N_30852,N_29351,N_29913);
and U30853 (N_30853,N_29466,N_29054);
nand U30854 (N_30854,N_29744,N_29623);
nor U30855 (N_30855,N_29285,N_29153);
and U30856 (N_30856,N_29244,N_29424);
nor U30857 (N_30857,N_29851,N_29587);
nor U30858 (N_30858,N_29999,N_29233);
nor U30859 (N_30859,N_29700,N_29605);
nor U30860 (N_30860,N_29839,N_29636);
or U30861 (N_30861,N_29395,N_29091);
xor U30862 (N_30862,N_29449,N_29498);
or U30863 (N_30863,N_29741,N_29777);
xor U30864 (N_30864,N_29923,N_29080);
nor U30865 (N_30865,N_29078,N_29412);
xnor U30866 (N_30866,N_29327,N_29669);
nor U30867 (N_30867,N_29295,N_29514);
nor U30868 (N_30868,N_29477,N_29921);
nand U30869 (N_30869,N_29142,N_29610);
and U30870 (N_30870,N_29727,N_29052);
and U30871 (N_30871,N_29123,N_29155);
and U30872 (N_30872,N_29905,N_29173);
and U30873 (N_30873,N_29724,N_29943);
nand U30874 (N_30874,N_29175,N_29225);
nor U30875 (N_30875,N_29398,N_29211);
or U30876 (N_30876,N_29886,N_29153);
xnor U30877 (N_30877,N_29446,N_29509);
or U30878 (N_30878,N_29449,N_29369);
xnor U30879 (N_30879,N_29071,N_29659);
nor U30880 (N_30880,N_29222,N_29068);
xor U30881 (N_30881,N_29333,N_29611);
and U30882 (N_30882,N_29529,N_29653);
and U30883 (N_30883,N_29240,N_29212);
nand U30884 (N_30884,N_29438,N_29934);
or U30885 (N_30885,N_29349,N_29862);
xnor U30886 (N_30886,N_29541,N_29946);
or U30887 (N_30887,N_29652,N_29788);
xor U30888 (N_30888,N_29916,N_29020);
xor U30889 (N_30889,N_29741,N_29322);
and U30890 (N_30890,N_29474,N_29807);
and U30891 (N_30891,N_29591,N_29281);
xnor U30892 (N_30892,N_29680,N_29226);
nand U30893 (N_30893,N_29314,N_29391);
xor U30894 (N_30894,N_29876,N_29063);
or U30895 (N_30895,N_29687,N_29677);
and U30896 (N_30896,N_29789,N_29820);
and U30897 (N_30897,N_29451,N_29730);
nor U30898 (N_30898,N_29737,N_29775);
and U30899 (N_30899,N_29162,N_29555);
nand U30900 (N_30900,N_29635,N_29699);
nor U30901 (N_30901,N_29203,N_29305);
nand U30902 (N_30902,N_29089,N_29128);
or U30903 (N_30903,N_29092,N_29318);
or U30904 (N_30904,N_29573,N_29711);
nand U30905 (N_30905,N_29835,N_29265);
xnor U30906 (N_30906,N_29242,N_29068);
and U30907 (N_30907,N_29280,N_29999);
nand U30908 (N_30908,N_29825,N_29465);
nand U30909 (N_30909,N_29091,N_29116);
nand U30910 (N_30910,N_29597,N_29490);
or U30911 (N_30911,N_29844,N_29637);
or U30912 (N_30912,N_29851,N_29478);
and U30913 (N_30913,N_29946,N_29990);
nor U30914 (N_30914,N_29797,N_29868);
nor U30915 (N_30915,N_29495,N_29854);
and U30916 (N_30916,N_29879,N_29507);
nand U30917 (N_30917,N_29632,N_29989);
and U30918 (N_30918,N_29926,N_29166);
xor U30919 (N_30919,N_29421,N_29493);
nor U30920 (N_30920,N_29834,N_29534);
xor U30921 (N_30921,N_29788,N_29622);
and U30922 (N_30922,N_29001,N_29883);
or U30923 (N_30923,N_29788,N_29521);
nand U30924 (N_30924,N_29466,N_29759);
xor U30925 (N_30925,N_29531,N_29888);
and U30926 (N_30926,N_29071,N_29465);
xor U30927 (N_30927,N_29089,N_29278);
nor U30928 (N_30928,N_29998,N_29264);
or U30929 (N_30929,N_29772,N_29032);
and U30930 (N_30930,N_29723,N_29456);
xnor U30931 (N_30931,N_29558,N_29360);
xnor U30932 (N_30932,N_29879,N_29284);
nand U30933 (N_30933,N_29244,N_29932);
nor U30934 (N_30934,N_29714,N_29502);
nor U30935 (N_30935,N_29511,N_29494);
nor U30936 (N_30936,N_29490,N_29278);
nand U30937 (N_30937,N_29165,N_29760);
nand U30938 (N_30938,N_29572,N_29176);
and U30939 (N_30939,N_29380,N_29265);
nor U30940 (N_30940,N_29490,N_29141);
nor U30941 (N_30941,N_29869,N_29311);
nor U30942 (N_30942,N_29604,N_29455);
and U30943 (N_30943,N_29750,N_29195);
and U30944 (N_30944,N_29367,N_29192);
and U30945 (N_30945,N_29984,N_29727);
and U30946 (N_30946,N_29502,N_29300);
or U30947 (N_30947,N_29755,N_29224);
or U30948 (N_30948,N_29055,N_29498);
xnor U30949 (N_30949,N_29888,N_29740);
xnor U30950 (N_30950,N_29539,N_29251);
nor U30951 (N_30951,N_29939,N_29075);
and U30952 (N_30952,N_29195,N_29461);
and U30953 (N_30953,N_29214,N_29905);
nand U30954 (N_30954,N_29795,N_29122);
and U30955 (N_30955,N_29467,N_29592);
xnor U30956 (N_30956,N_29763,N_29030);
or U30957 (N_30957,N_29375,N_29504);
xor U30958 (N_30958,N_29822,N_29389);
or U30959 (N_30959,N_29996,N_29038);
nand U30960 (N_30960,N_29159,N_29101);
or U30961 (N_30961,N_29986,N_29862);
xnor U30962 (N_30962,N_29367,N_29202);
and U30963 (N_30963,N_29848,N_29949);
nor U30964 (N_30964,N_29794,N_29243);
and U30965 (N_30965,N_29288,N_29415);
and U30966 (N_30966,N_29698,N_29883);
xor U30967 (N_30967,N_29648,N_29300);
xor U30968 (N_30968,N_29562,N_29508);
or U30969 (N_30969,N_29020,N_29279);
or U30970 (N_30970,N_29029,N_29921);
xor U30971 (N_30971,N_29640,N_29605);
or U30972 (N_30972,N_29191,N_29127);
and U30973 (N_30973,N_29385,N_29631);
nand U30974 (N_30974,N_29404,N_29892);
and U30975 (N_30975,N_29774,N_29687);
or U30976 (N_30976,N_29806,N_29195);
and U30977 (N_30977,N_29328,N_29019);
xnor U30978 (N_30978,N_29420,N_29802);
xor U30979 (N_30979,N_29569,N_29533);
nor U30980 (N_30980,N_29272,N_29674);
or U30981 (N_30981,N_29016,N_29902);
and U30982 (N_30982,N_29370,N_29301);
nand U30983 (N_30983,N_29069,N_29973);
or U30984 (N_30984,N_29630,N_29565);
and U30985 (N_30985,N_29656,N_29529);
nor U30986 (N_30986,N_29961,N_29612);
xnor U30987 (N_30987,N_29130,N_29165);
and U30988 (N_30988,N_29801,N_29730);
or U30989 (N_30989,N_29442,N_29303);
and U30990 (N_30990,N_29427,N_29209);
or U30991 (N_30991,N_29591,N_29406);
nand U30992 (N_30992,N_29567,N_29921);
xor U30993 (N_30993,N_29396,N_29349);
nor U30994 (N_30994,N_29322,N_29303);
and U30995 (N_30995,N_29571,N_29705);
nand U30996 (N_30996,N_29063,N_29926);
and U30997 (N_30997,N_29903,N_29240);
or U30998 (N_30998,N_29231,N_29562);
nor U30999 (N_30999,N_29971,N_29324);
nand U31000 (N_31000,N_30677,N_30641);
and U31001 (N_31001,N_30497,N_30123);
xnor U31002 (N_31002,N_30605,N_30846);
nor U31003 (N_31003,N_30749,N_30137);
or U31004 (N_31004,N_30107,N_30191);
or U31005 (N_31005,N_30366,N_30817);
xor U31006 (N_31006,N_30401,N_30766);
nor U31007 (N_31007,N_30144,N_30014);
xor U31008 (N_31008,N_30593,N_30073);
or U31009 (N_31009,N_30718,N_30692);
and U31010 (N_31010,N_30238,N_30503);
or U31011 (N_31011,N_30303,N_30312);
nor U31012 (N_31012,N_30765,N_30147);
nor U31013 (N_31013,N_30720,N_30042);
or U31014 (N_31014,N_30878,N_30842);
or U31015 (N_31015,N_30127,N_30086);
nor U31016 (N_31016,N_30635,N_30654);
or U31017 (N_31017,N_30645,N_30828);
nand U31018 (N_31018,N_30166,N_30811);
and U31019 (N_31019,N_30214,N_30262);
or U31020 (N_31020,N_30923,N_30355);
and U31021 (N_31021,N_30689,N_30728);
nand U31022 (N_31022,N_30610,N_30442);
nand U31023 (N_31023,N_30016,N_30311);
nand U31024 (N_31024,N_30545,N_30911);
nor U31025 (N_31025,N_30320,N_30054);
xnor U31026 (N_31026,N_30393,N_30854);
and U31027 (N_31027,N_30939,N_30348);
xor U31028 (N_31028,N_30023,N_30776);
nand U31029 (N_31029,N_30027,N_30213);
and U31030 (N_31030,N_30268,N_30211);
nor U31031 (N_31031,N_30972,N_30255);
or U31032 (N_31032,N_30101,N_30921);
and U31033 (N_31033,N_30087,N_30660);
xor U31034 (N_31034,N_30987,N_30613);
nand U31035 (N_31035,N_30914,N_30050);
and U31036 (N_31036,N_30427,N_30192);
and U31037 (N_31037,N_30063,N_30864);
nor U31038 (N_31038,N_30411,N_30479);
and U31039 (N_31039,N_30335,N_30448);
nand U31040 (N_31040,N_30602,N_30406);
nor U31041 (N_31041,N_30536,N_30104);
nor U31042 (N_31042,N_30953,N_30224);
and U31043 (N_31043,N_30724,N_30621);
or U31044 (N_31044,N_30652,N_30866);
and U31045 (N_31045,N_30746,N_30186);
and U31046 (N_31046,N_30528,N_30785);
nor U31047 (N_31047,N_30417,N_30970);
or U31048 (N_31048,N_30252,N_30465);
nand U31049 (N_31049,N_30793,N_30871);
xor U31050 (N_31050,N_30258,N_30695);
xnor U31051 (N_31051,N_30004,N_30136);
and U31052 (N_31052,N_30261,N_30259);
nand U31053 (N_31053,N_30555,N_30346);
xnor U31054 (N_31054,N_30881,N_30969);
xor U31055 (N_31055,N_30336,N_30025);
and U31056 (N_31056,N_30468,N_30499);
nor U31057 (N_31057,N_30351,N_30625);
or U31058 (N_31058,N_30330,N_30365);
nor U31059 (N_31059,N_30474,N_30640);
nand U31060 (N_31060,N_30813,N_30362);
and U31061 (N_31061,N_30354,N_30217);
xor U31062 (N_31062,N_30380,N_30590);
xnor U31063 (N_31063,N_30582,N_30600);
and U31064 (N_31064,N_30648,N_30575);
nand U31065 (N_31065,N_30650,N_30810);
xor U31066 (N_31066,N_30830,N_30250);
or U31067 (N_31067,N_30378,N_30559);
or U31068 (N_31068,N_30247,N_30463);
or U31069 (N_31069,N_30055,N_30288);
nor U31070 (N_31070,N_30690,N_30790);
and U31071 (N_31071,N_30398,N_30077);
nor U31072 (N_31072,N_30457,N_30342);
xnor U31073 (N_31073,N_30620,N_30289);
nor U31074 (N_31074,N_30230,N_30048);
nand U31075 (N_31075,N_30198,N_30879);
or U31076 (N_31076,N_30476,N_30160);
xor U31077 (N_31077,N_30979,N_30059);
nand U31078 (N_31078,N_30928,N_30314);
nor U31079 (N_31079,N_30840,N_30132);
or U31080 (N_31080,N_30484,N_30642);
or U31081 (N_31081,N_30345,N_30761);
and U31082 (N_31082,N_30157,N_30112);
xor U31083 (N_31083,N_30331,N_30172);
nand U31084 (N_31084,N_30433,N_30013);
nand U31085 (N_31085,N_30540,N_30882);
xnor U31086 (N_31086,N_30002,N_30412);
nand U31087 (N_31087,N_30246,N_30535);
or U31088 (N_31088,N_30341,N_30232);
and U31089 (N_31089,N_30619,N_30973);
nor U31090 (N_31090,N_30103,N_30370);
nand U31091 (N_31091,N_30944,N_30279);
nand U31092 (N_31092,N_30174,N_30824);
xnor U31093 (N_31093,N_30594,N_30332);
nor U31094 (N_31094,N_30905,N_30421);
or U31095 (N_31095,N_30321,N_30437);
xor U31096 (N_31096,N_30357,N_30673);
or U31097 (N_31097,N_30694,N_30361);
xnor U31098 (N_31098,N_30521,N_30805);
xnor U31099 (N_31099,N_30797,N_30825);
or U31100 (N_31100,N_30651,N_30902);
xor U31101 (N_31101,N_30963,N_30742);
and U31102 (N_31102,N_30243,N_30447);
and U31103 (N_31103,N_30129,N_30067);
xor U31104 (N_31104,N_30566,N_30032);
nor U31105 (N_31105,N_30177,N_30164);
xnor U31106 (N_31106,N_30522,N_30773);
and U31107 (N_31107,N_30359,N_30111);
xor U31108 (N_31108,N_30889,N_30748);
and U31109 (N_31109,N_30135,N_30181);
and U31110 (N_31110,N_30723,N_30576);
and U31111 (N_31111,N_30852,N_30041);
or U31112 (N_31112,N_30883,N_30705);
and U31113 (N_31113,N_30900,N_30110);
nand U31114 (N_31114,N_30441,N_30204);
nor U31115 (N_31115,N_30685,N_30633);
nor U31116 (N_31116,N_30139,N_30940);
nand U31117 (N_31117,N_30407,N_30193);
or U31118 (N_31118,N_30901,N_30119);
nor U31119 (N_31119,N_30024,N_30151);
xnor U31120 (N_31120,N_30012,N_30225);
nand U31121 (N_31121,N_30470,N_30502);
and U31122 (N_31122,N_30071,N_30865);
xnor U31123 (N_31123,N_30131,N_30957);
xor U31124 (N_31124,N_30236,N_30426);
nor U31125 (N_31125,N_30924,N_30931);
xnor U31126 (N_31126,N_30767,N_30126);
and U31127 (N_31127,N_30971,N_30892);
and U31128 (N_31128,N_30780,N_30507);
nand U31129 (N_31129,N_30814,N_30933);
and U31130 (N_31130,N_30631,N_30226);
or U31131 (N_31131,N_30095,N_30333);
nand U31132 (N_31132,N_30880,N_30170);
nand U31133 (N_31133,N_30372,N_30493);
nor U31134 (N_31134,N_30294,N_30591);
or U31135 (N_31135,N_30644,N_30952);
and U31136 (N_31136,N_30490,N_30932);
nor U31137 (N_31137,N_30097,N_30158);
xnor U31138 (N_31138,N_30980,N_30809);
or U31139 (N_31139,N_30698,N_30179);
nor U31140 (N_31140,N_30395,N_30385);
or U31141 (N_31141,N_30877,N_30205);
xnor U31142 (N_31142,N_30701,N_30115);
nor U31143 (N_31143,N_30770,N_30783);
and U31144 (N_31144,N_30089,N_30483);
xnor U31145 (N_31145,N_30208,N_30322);
and U31146 (N_31146,N_30315,N_30628);
xor U31147 (N_31147,N_30974,N_30791);
or U31148 (N_31148,N_30683,N_30563);
and U31149 (N_31149,N_30121,N_30416);
or U31150 (N_31150,N_30659,N_30189);
nand U31151 (N_31151,N_30099,N_30612);
nor U31152 (N_31152,N_30287,N_30964);
and U31153 (N_31153,N_30556,N_30245);
xor U31154 (N_31154,N_30904,N_30046);
nand U31155 (N_31155,N_30410,N_30446);
and U31156 (N_31156,N_30327,N_30992);
or U31157 (N_31157,N_30985,N_30532);
or U31158 (N_31158,N_30888,N_30364);
nand U31159 (N_31159,N_30848,N_30508);
or U31160 (N_31160,N_30623,N_30229);
nand U31161 (N_31161,N_30068,N_30168);
xnor U31162 (N_31162,N_30664,N_30235);
xor U31163 (N_31163,N_30898,N_30758);
nor U31164 (N_31164,N_30759,N_30833);
nor U31165 (N_31165,N_30053,N_30845);
nor U31166 (N_31166,N_30832,N_30313);
xor U31167 (N_31167,N_30571,N_30757);
nand U31168 (N_31168,N_30975,N_30965);
xor U31169 (N_31169,N_30386,N_30344);
xor U31170 (N_31170,N_30423,N_30998);
nor U31171 (N_31171,N_30609,N_30498);
and U31172 (N_31172,N_30091,N_30078);
nand U31173 (N_31173,N_30988,N_30171);
xnor U31174 (N_31174,N_30523,N_30873);
or U31175 (N_31175,N_30300,N_30368);
nand U31176 (N_31176,N_30917,N_30572);
or U31177 (N_31177,N_30936,N_30281);
and U31178 (N_31178,N_30719,N_30422);
nor U31179 (N_31179,N_30352,N_30267);
and U31180 (N_31180,N_30968,N_30227);
and U31181 (N_31181,N_30907,N_30467);
nand U31182 (N_31182,N_30496,N_30298);
nor U31183 (N_31183,N_30280,N_30614);
xnor U31184 (N_31184,N_30316,N_30649);
xnor U31185 (N_31185,N_30146,N_30989);
and U31186 (N_31186,N_30360,N_30234);
and U31187 (N_31187,N_30517,N_30000);
or U31188 (N_31188,N_30215,N_30634);
nor U31189 (N_31189,N_30834,N_30688);
nor U31190 (N_31190,N_30925,N_30596);
nand U31191 (N_31191,N_30358,N_30977);
xnor U31192 (N_31192,N_30859,N_30529);
nor U31193 (N_31193,N_30935,N_30734);
and U31194 (N_31194,N_30049,N_30755);
xnor U31195 (N_31195,N_30425,N_30047);
nor U31196 (N_31196,N_30062,N_30339);
nor U31197 (N_31197,N_30663,N_30283);
nand U31198 (N_31198,N_30820,N_30815);
and U31199 (N_31199,N_30819,N_30870);
and U31200 (N_31200,N_30549,N_30491);
or U31201 (N_31201,N_30022,N_30367);
xnor U31202 (N_31202,N_30868,N_30837);
or U31203 (N_31203,N_30750,N_30180);
nor U31204 (N_31204,N_30408,N_30272);
nand U31205 (N_31205,N_30253,N_30927);
nand U31206 (N_31206,N_30741,N_30730);
nand U31207 (N_31207,N_30343,N_30057);
nand U31208 (N_31208,N_30938,N_30578);
xnor U31209 (N_31209,N_30184,N_30960);
or U31210 (N_31210,N_30100,N_30244);
nor U31211 (N_31211,N_30028,N_30849);
or U31212 (N_31212,N_30429,N_30116);
xnor U31213 (N_31213,N_30504,N_30188);
or U31214 (N_31214,N_30264,N_30066);
or U31215 (N_31215,N_30472,N_30093);
nand U31216 (N_31216,N_30375,N_30396);
nor U31217 (N_31217,N_30804,N_30274);
or U31218 (N_31218,N_30376,N_30646);
and U31219 (N_31219,N_30223,N_30318);
nor U31220 (N_31220,N_30550,N_30285);
nor U31221 (N_31221,N_30994,N_30141);
nand U31222 (N_31222,N_30182,N_30976);
xnor U31223 (N_31223,N_30413,N_30800);
or U31224 (N_31224,N_30913,N_30807);
nor U31225 (N_31225,N_30494,N_30886);
nand U31226 (N_31226,N_30282,N_30531);
nand U31227 (N_31227,N_30478,N_30109);
or U31228 (N_31228,N_30430,N_30469);
nand U31229 (N_31229,N_30505,N_30548);
and U31230 (N_31230,N_30302,N_30947);
nor U31231 (N_31231,N_30890,N_30768);
nor U31232 (N_31232,N_30954,N_30639);
or U31233 (N_31233,N_30090,N_30756);
and U31234 (N_31234,N_30251,N_30260);
or U31235 (N_31235,N_30568,N_30176);
nand U31236 (N_31236,N_30473,N_30702);
xnor U31237 (N_31237,N_30542,N_30044);
nor U31238 (N_31238,N_30618,N_30557);
nor U31239 (N_31239,N_30753,N_30875);
nand U31240 (N_31240,N_30220,N_30165);
and U31241 (N_31241,N_30424,N_30801);
or U31242 (N_31242,N_30452,N_30707);
nand U31243 (N_31243,N_30597,N_30029);
xor U31244 (N_31244,N_30169,N_30850);
or U31245 (N_31245,N_30622,N_30291);
nor U31246 (N_31246,N_30983,N_30482);
or U31247 (N_31247,N_30667,N_30661);
nor U31248 (N_31248,N_30299,N_30951);
nand U31249 (N_31249,N_30212,N_30629);
and U31250 (N_31250,N_30604,N_30038);
or U31251 (N_31251,N_30671,N_30037);
and U31252 (N_31252,N_30295,N_30304);
and U31253 (N_31253,N_30996,N_30516);
nor U31254 (N_31254,N_30506,N_30838);
nor U31255 (N_31255,N_30580,N_30802);
nor U31256 (N_31256,N_30069,N_30872);
or U31257 (N_31257,N_30374,N_30058);
or U31258 (N_31258,N_30019,N_30818);
xnor U31259 (N_31259,N_30265,N_30601);
and U31260 (N_31260,N_30567,N_30538);
nor U31261 (N_31261,N_30487,N_30409);
nand U31262 (N_31262,N_30684,N_30812);
and U31263 (N_31263,N_30347,N_30586);
and U31264 (N_31264,N_30606,N_30450);
nand U31265 (N_31265,N_30079,N_30390);
or U31266 (N_31266,N_30981,N_30527);
or U31267 (N_31267,N_30439,N_30826);
xor U31268 (N_31268,N_30240,N_30190);
nand U31269 (N_31269,N_30511,N_30383);
nor U31270 (N_31270,N_30726,N_30569);
nand U31271 (N_31271,N_30562,N_30142);
nand U31272 (N_31272,N_30530,N_30431);
and U31273 (N_31273,N_30449,N_30096);
or U31274 (N_31274,N_30999,N_30993);
and U31275 (N_31275,N_30150,N_30163);
nor U31276 (N_31276,N_30061,N_30722);
or U31277 (N_31277,N_30896,N_30159);
nor U31278 (N_31278,N_30679,N_30662);
xnor U31279 (N_31279,N_30105,N_30754);
nor U31280 (N_31280,N_30821,N_30534);
or U31281 (N_31281,N_30006,N_30435);
or U31282 (N_31282,N_30709,N_30948);
xor U31283 (N_31283,N_30519,N_30309);
xnor U31284 (N_31284,N_30488,N_30518);
xor U31285 (N_31285,N_30665,N_30120);
nand U31286 (N_31286,N_30305,N_30329);
xor U31287 (N_31287,N_30387,N_30277);
nand U31288 (N_31288,N_30772,N_30391);
and U31289 (N_31289,N_30353,N_30585);
and U31290 (N_31290,N_30788,N_30481);
or U31291 (N_31291,N_30843,N_30455);
or U31292 (N_31292,N_30658,N_30686);
xnor U31293 (N_31293,N_30501,N_30611);
nand U31294 (N_31294,N_30145,N_30573);
nand U31295 (N_31295,N_30489,N_30007);
xor U31296 (N_31296,N_30543,N_30713);
or U31297 (N_31297,N_30148,N_30607);
nor U31298 (N_31298,N_30737,N_30194);
and U31299 (N_31299,N_30377,N_30588);
and U31300 (N_31300,N_30434,N_30349);
and U31301 (N_31301,N_30691,N_30231);
or U31302 (N_31302,N_30738,N_30237);
xnor U31303 (N_31303,N_30781,N_30798);
nand U31304 (N_31304,N_30248,N_30031);
or U31305 (N_31305,N_30676,N_30117);
and U31306 (N_31306,N_30862,N_30356);
or U31307 (N_31307,N_30775,N_30161);
nor U31308 (N_31308,N_30884,N_30088);
or U31309 (N_31309,N_30495,N_30554);
nor U31310 (N_31310,N_30143,N_30399);
nand U31311 (N_31311,N_30510,N_30711);
nand U31312 (N_31312,N_30920,N_30477);
or U31313 (N_31313,N_30712,N_30687);
nor U31314 (N_31314,N_30369,N_30937);
nand U31315 (N_31315,N_30466,N_30891);
xnor U31316 (N_31316,N_30736,N_30887);
or U31317 (N_31317,N_30187,N_30419);
xor U31318 (N_31318,N_30906,N_30453);
and U31319 (N_31319,N_30706,N_30856);
and U31320 (N_31320,N_30990,N_30777);
nor U31321 (N_31321,N_30286,N_30106);
xor U31322 (N_31322,N_30978,N_30092);
and U31323 (N_31323,N_30325,N_30789);
xor U31324 (N_31324,N_30492,N_30727);
and U31325 (N_31325,N_30363,N_30130);
nand U31326 (N_31326,N_30853,N_30546);
or U31327 (N_31327,N_30307,N_30949);
and U31328 (N_31328,N_30052,N_30680);
and U31329 (N_31329,N_30216,N_30670);
nand U31330 (N_31330,N_30509,N_30404);
and U31331 (N_31331,N_30729,N_30637);
nand U31332 (N_31332,N_30786,N_30595);
or U31333 (N_31333,N_30196,N_30666);
nand U31334 (N_31334,N_30926,N_30657);
or U31335 (N_31335,N_30486,N_30001);
xnor U31336 (N_31336,N_30323,N_30869);
xnor U31337 (N_31337,N_30743,N_30721);
and U31338 (N_31338,N_30855,N_30570);
nor U31339 (N_31339,N_30133,N_30122);
xor U31340 (N_31340,N_30074,N_30301);
and U31341 (N_31341,N_30459,N_30806);
xor U31342 (N_31342,N_30045,N_30337);
nand U31343 (N_31343,N_30524,N_30156);
xnor U31344 (N_31344,N_30792,N_30056);
xor U31345 (N_31345,N_30039,N_30072);
or U31346 (N_31346,N_30270,N_30296);
or U31347 (N_31347,N_30708,N_30839);
nand U31348 (N_31348,N_30384,N_30577);
nor U31349 (N_31349,N_30273,N_30956);
nor U31350 (N_31350,N_30603,N_30153);
nand U31351 (N_31351,N_30995,N_30615);
or U31352 (N_31352,N_30822,N_30836);
and U31353 (N_31353,N_30460,N_30451);
nor U31354 (N_31354,N_30827,N_30249);
and U31355 (N_31355,N_30740,N_30874);
and U31356 (N_31356,N_30991,N_30829);
or U31357 (N_31357,N_30185,N_30015);
xnor U31358 (N_31358,N_30867,N_30541);
nor U31359 (N_31359,N_30202,N_30796);
nand U31360 (N_31360,N_30895,N_30152);
xnor U31361 (N_31361,N_30831,N_30515);
nand U31362 (N_31362,N_30579,N_30266);
or U31363 (N_31363,N_30725,N_30310);
or U31364 (N_31364,N_30394,N_30254);
nand U31365 (N_31365,N_30292,N_30138);
xnor U31366 (N_31366,N_30700,N_30581);
xor U31367 (N_31367,N_30400,N_30564);
xor U31368 (N_31368,N_30584,N_30678);
and U31369 (N_31369,N_30297,N_30373);
and U31370 (N_31370,N_30608,N_30958);
xnor U31371 (N_31371,N_30520,N_30835);
xnor U31372 (N_31372,N_30514,N_30210);
or U31373 (N_31373,N_30636,N_30922);
and U31374 (N_31374,N_30402,N_30544);
nor U31375 (N_31375,N_30241,N_30233);
nor U31376 (N_31376,N_30128,N_30060);
nor U31377 (N_31377,N_30945,N_30910);
or U31378 (N_31378,N_30456,N_30893);
and U31379 (N_31379,N_30464,N_30065);
or U31380 (N_31380,N_30043,N_30592);
or U31381 (N_31381,N_30269,N_30275);
or U31382 (N_31382,N_30026,N_30080);
or U31383 (N_31383,N_30918,N_30731);
nor U31384 (N_31384,N_30710,N_30219);
or U31385 (N_31385,N_30263,N_30693);
nand U31386 (N_31386,N_30885,N_30714);
nand U31387 (N_31387,N_30512,N_30102);
nor U31388 (N_31388,N_30454,N_30668);
nand U31389 (N_31389,N_30943,N_30716);
nor U31390 (N_31390,N_30076,N_30876);
and U31391 (N_31391,N_30787,N_30445);
nor U31392 (N_31392,N_30183,N_30929);
and U31393 (N_31393,N_30256,N_30010);
xor U31394 (N_31394,N_30715,N_30317);
and U31395 (N_31395,N_30070,N_30500);
nor U31396 (N_31396,N_30035,N_30334);
nor U31397 (N_31397,N_30338,N_30643);
nand U31398 (N_31398,N_30082,N_30203);
and U31399 (N_31399,N_30934,N_30290);
nor U31400 (N_31400,N_30703,N_30271);
or U31401 (N_31401,N_30149,N_30560);
xnor U31402 (N_31402,N_30485,N_30583);
or U31403 (N_31403,N_30098,N_30764);
xnor U31404 (N_31404,N_30199,N_30222);
and U31405 (N_31405,N_30306,N_30967);
xor U31406 (N_31406,N_30392,N_30242);
or U31407 (N_31407,N_30784,N_30340);
or U31408 (N_31408,N_30547,N_30036);
xnor U31409 (N_31409,N_30195,N_30653);
nor U31410 (N_31410,N_30655,N_30950);
nor U31411 (N_31411,N_30844,N_30656);
nand U31412 (N_31412,N_30113,N_30647);
or U31413 (N_31413,N_30760,N_30778);
or U31414 (N_31414,N_30420,N_30173);
nor U31415 (N_31415,N_30388,N_30382);
and U31416 (N_31416,N_30574,N_30284);
and U31417 (N_31417,N_30218,N_30552);
or U31418 (N_31418,N_30669,N_30475);
nor U31419 (N_31419,N_30672,N_30841);
and U31420 (N_31420,N_30403,N_30206);
nor U31421 (N_31421,N_30438,N_30782);
or U31422 (N_31422,N_30397,N_30436);
or U31423 (N_31423,N_30955,N_30860);
xor U31424 (N_31424,N_30379,N_30178);
and U31425 (N_31425,N_30005,N_30617);
nor U31426 (N_31426,N_30897,N_30941);
or U31427 (N_31427,N_30966,N_30732);
nor U31428 (N_31428,N_30697,N_30616);
and U31429 (N_31429,N_30040,N_30744);
or U31430 (N_31430,N_30207,N_30908);
nand U31431 (N_31431,N_30350,N_30751);
or U31432 (N_31432,N_30696,N_30916);
nand U31433 (N_31433,N_30114,N_30735);
or U31434 (N_31434,N_30471,N_30816);
nand U31435 (N_31435,N_30221,N_30175);
nor U31436 (N_31436,N_30167,N_30717);
xor U31437 (N_31437,N_30539,N_30480);
nor U31438 (N_31438,N_30084,N_30381);
xnor U31439 (N_31439,N_30526,N_30458);
nor U31440 (N_31440,N_30986,N_30962);
nand U31441 (N_31441,N_30861,N_30324);
nand U31442 (N_31442,N_30632,N_30795);
nand U31443 (N_31443,N_30771,N_30598);
xnor U31444 (N_31444,N_30011,N_30930);
or U31445 (N_31445,N_30326,N_30699);
nor U31446 (N_31446,N_30553,N_30774);
and U31447 (N_31447,N_30551,N_30857);
nor U31448 (N_31448,N_30858,N_30462);
nand U31449 (N_31449,N_30899,N_30209);
nand U31450 (N_31450,N_30030,N_30108);
or U31451 (N_31451,N_30681,N_30624);
nand U31452 (N_31452,N_30201,N_30682);
nor U31453 (N_31453,N_30009,N_30565);
xnor U31454 (N_31454,N_30440,N_30017);
nor U31455 (N_31455,N_30328,N_30094);
nand U31456 (N_31456,N_30081,N_30984);
and U31457 (N_31457,N_30803,N_30739);
and U31458 (N_31458,N_30154,N_30162);
and U31459 (N_31459,N_30525,N_30308);
and U31460 (N_31460,N_30200,N_30747);
and U31461 (N_31461,N_30414,N_30432);
and U31462 (N_31462,N_30064,N_30704);
nand U31463 (N_31463,N_30239,N_30118);
or U31464 (N_31464,N_30083,N_30942);
nor U31465 (N_31465,N_30033,N_30919);
xor U31466 (N_31466,N_30982,N_30794);
and U31467 (N_31467,N_30799,N_30599);
nand U31468 (N_31468,N_30808,N_30155);
xor U31469 (N_31469,N_30561,N_30959);
nor U31470 (N_31470,N_30863,N_30674);
nor U31471 (N_31471,N_30894,N_30319);
or U31472 (N_31472,N_30779,N_30533);
and U31473 (N_31473,N_30461,N_30587);
or U31474 (N_31474,N_30003,N_30293);
and U31475 (N_31475,N_30444,N_30020);
nand U31476 (N_31476,N_30558,N_30389);
nand U31477 (N_31477,N_30034,N_30075);
nor U31478 (N_31478,N_30769,N_30847);
and U31479 (N_31479,N_30627,N_30745);
nor U31480 (N_31480,N_30630,N_30638);
xnor U31481 (N_31481,N_30903,N_30018);
nor U31482 (N_31482,N_30537,N_30051);
nand U31483 (N_31483,N_30371,N_30946);
nor U31484 (N_31484,N_30675,N_30909);
nor U31485 (N_31485,N_30626,N_30851);
nor U31486 (N_31486,N_30763,N_30140);
xnor U31487 (N_31487,N_30197,N_30134);
nor U31488 (N_31488,N_30823,N_30589);
xor U31489 (N_31489,N_30415,N_30228);
or U31490 (N_31490,N_30021,N_30085);
xor U31491 (N_31491,N_30752,N_30915);
nand U31492 (N_31492,N_30278,N_30008);
xor U31493 (N_31493,N_30428,N_30257);
and U31494 (N_31494,N_30762,N_30513);
nand U31495 (N_31495,N_30997,N_30276);
or U31496 (N_31496,N_30961,N_30418);
or U31497 (N_31497,N_30125,N_30443);
nand U31498 (N_31498,N_30124,N_30912);
or U31499 (N_31499,N_30733,N_30405);
xor U31500 (N_31500,N_30998,N_30583);
nor U31501 (N_31501,N_30552,N_30254);
nor U31502 (N_31502,N_30521,N_30147);
or U31503 (N_31503,N_30700,N_30616);
or U31504 (N_31504,N_30606,N_30946);
and U31505 (N_31505,N_30963,N_30331);
nor U31506 (N_31506,N_30605,N_30924);
nand U31507 (N_31507,N_30382,N_30259);
nor U31508 (N_31508,N_30054,N_30602);
nor U31509 (N_31509,N_30999,N_30236);
xnor U31510 (N_31510,N_30816,N_30425);
nor U31511 (N_31511,N_30993,N_30920);
xor U31512 (N_31512,N_30289,N_30362);
and U31513 (N_31513,N_30043,N_30271);
xor U31514 (N_31514,N_30236,N_30903);
or U31515 (N_31515,N_30901,N_30312);
nor U31516 (N_31516,N_30075,N_30827);
and U31517 (N_31517,N_30943,N_30836);
or U31518 (N_31518,N_30796,N_30722);
or U31519 (N_31519,N_30944,N_30475);
and U31520 (N_31520,N_30069,N_30369);
nor U31521 (N_31521,N_30070,N_30756);
and U31522 (N_31522,N_30220,N_30651);
nor U31523 (N_31523,N_30878,N_30760);
nand U31524 (N_31524,N_30093,N_30851);
nor U31525 (N_31525,N_30380,N_30623);
and U31526 (N_31526,N_30182,N_30158);
and U31527 (N_31527,N_30199,N_30539);
nand U31528 (N_31528,N_30312,N_30252);
and U31529 (N_31529,N_30280,N_30021);
or U31530 (N_31530,N_30080,N_30993);
nor U31531 (N_31531,N_30038,N_30373);
or U31532 (N_31532,N_30404,N_30000);
and U31533 (N_31533,N_30512,N_30333);
nand U31534 (N_31534,N_30032,N_30574);
or U31535 (N_31535,N_30284,N_30783);
nor U31536 (N_31536,N_30269,N_30425);
or U31537 (N_31537,N_30443,N_30220);
or U31538 (N_31538,N_30410,N_30314);
or U31539 (N_31539,N_30489,N_30896);
xnor U31540 (N_31540,N_30226,N_30324);
nor U31541 (N_31541,N_30194,N_30417);
xnor U31542 (N_31542,N_30682,N_30122);
and U31543 (N_31543,N_30490,N_30613);
and U31544 (N_31544,N_30437,N_30042);
and U31545 (N_31545,N_30639,N_30717);
nand U31546 (N_31546,N_30131,N_30898);
nor U31547 (N_31547,N_30547,N_30790);
nand U31548 (N_31548,N_30490,N_30491);
nand U31549 (N_31549,N_30762,N_30751);
nor U31550 (N_31550,N_30590,N_30035);
nand U31551 (N_31551,N_30567,N_30171);
nor U31552 (N_31552,N_30863,N_30902);
nor U31553 (N_31553,N_30382,N_30644);
xnor U31554 (N_31554,N_30892,N_30518);
nor U31555 (N_31555,N_30653,N_30962);
and U31556 (N_31556,N_30064,N_30889);
xnor U31557 (N_31557,N_30153,N_30639);
nand U31558 (N_31558,N_30032,N_30348);
nor U31559 (N_31559,N_30832,N_30819);
nor U31560 (N_31560,N_30471,N_30297);
xor U31561 (N_31561,N_30720,N_30832);
nand U31562 (N_31562,N_30977,N_30275);
and U31563 (N_31563,N_30899,N_30883);
nand U31564 (N_31564,N_30312,N_30172);
and U31565 (N_31565,N_30384,N_30138);
or U31566 (N_31566,N_30696,N_30092);
nand U31567 (N_31567,N_30519,N_30047);
or U31568 (N_31568,N_30622,N_30989);
xnor U31569 (N_31569,N_30881,N_30246);
nor U31570 (N_31570,N_30437,N_30848);
nor U31571 (N_31571,N_30569,N_30678);
nand U31572 (N_31572,N_30363,N_30656);
xnor U31573 (N_31573,N_30597,N_30098);
and U31574 (N_31574,N_30055,N_30899);
or U31575 (N_31575,N_30645,N_30695);
or U31576 (N_31576,N_30865,N_30005);
nor U31577 (N_31577,N_30772,N_30510);
nand U31578 (N_31578,N_30074,N_30410);
nor U31579 (N_31579,N_30161,N_30556);
xor U31580 (N_31580,N_30146,N_30446);
nor U31581 (N_31581,N_30806,N_30203);
xor U31582 (N_31582,N_30449,N_30358);
xor U31583 (N_31583,N_30049,N_30068);
or U31584 (N_31584,N_30614,N_30527);
nand U31585 (N_31585,N_30961,N_30782);
xnor U31586 (N_31586,N_30488,N_30976);
and U31587 (N_31587,N_30690,N_30947);
or U31588 (N_31588,N_30015,N_30048);
and U31589 (N_31589,N_30266,N_30864);
nand U31590 (N_31590,N_30826,N_30982);
nand U31591 (N_31591,N_30926,N_30078);
or U31592 (N_31592,N_30321,N_30766);
xor U31593 (N_31593,N_30925,N_30315);
nand U31594 (N_31594,N_30744,N_30203);
nand U31595 (N_31595,N_30153,N_30664);
nor U31596 (N_31596,N_30330,N_30200);
nor U31597 (N_31597,N_30655,N_30996);
xor U31598 (N_31598,N_30060,N_30272);
xnor U31599 (N_31599,N_30158,N_30364);
xnor U31600 (N_31600,N_30417,N_30092);
nand U31601 (N_31601,N_30643,N_30554);
or U31602 (N_31602,N_30928,N_30838);
nand U31603 (N_31603,N_30695,N_30138);
and U31604 (N_31604,N_30125,N_30168);
nand U31605 (N_31605,N_30426,N_30214);
nor U31606 (N_31606,N_30889,N_30232);
xnor U31607 (N_31607,N_30683,N_30535);
nand U31608 (N_31608,N_30826,N_30814);
xor U31609 (N_31609,N_30173,N_30312);
or U31610 (N_31610,N_30037,N_30840);
or U31611 (N_31611,N_30592,N_30599);
nor U31612 (N_31612,N_30082,N_30989);
and U31613 (N_31613,N_30346,N_30599);
and U31614 (N_31614,N_30294,N_30892);
nand U31615 (N_31615,N_30141,N_30638);
nand U31616 (N_31616,N_30009,N_30524);
or U31617 (N_31617,N_30296,N_30287);
and U31618 (N_31618,N_30344,N_30791);
nand U31619 (N_31619,N_30447,N_30133);
nand U31620 (N_31620,N_30053,N_30708);
and U31621 (N_31621,N_30216,N_30983);
nand U31622 (N_31622,N_30621,N_30099);
nand U31623 (N_31623,N_30353,N_30442);
nand U31624 (N_31624,N_30405,N_30096);
and U31625 (N_31625,N_30016,N_30203);
xor U31626 (N_31626,N_30319,N_30021);
or U31627 (N_31627,N_30952,N_30638);
and U31628 (N_31628,N_30848,N_30035);
and U31629 (N_31629,N_30258,N_30811);
xor U31630 (N_31630,N_30612,N_30993);
nor U31631 (N_31631,N_30488,N_30481);
xnor U31632 (N_31632,N_30331,N_30069);
xnor U31633 (N_31633,N_30999,N_30119);
xor U31634 (N_31634,N_30558,N_30759);
nand U31635 (N_31635,N_30796,N_30322);
nor U31636 (N_31636,N_30980,N_30476);
xor U31637 (N_31637,N_30420,N_30083);
nand U31638 (N_31638,N_30213,N_30153);
and U31639 (N_31639,N_30216,N_30893);
or U31640 (N_31640,N_30255,N_30999);
and U31641 (N_31641,N_30585,N_30062);
nor U31642 (N_31642,N_30751,N_30524);
and U31643 (N_31643,N_30347,N_30665);
and U31644 (N_31644,N_30477,N_30756);
or U31645 (N_31645,N_30628,N_30140);
nand U31646 (N_31646,N_30896,N_30323);
or U31647 (N_31647,N_30099,N_30035);
and U31648 (N_31648,N_30341,N_30718);
xor U31649 (N_31649,N_30038,N_30473);
xor U31650 (N_31650,N_30935,N_30836);
nand U31651 (N_31651,N_30762,N_30904);
nand U31652 (N_31652,N_30592,N_30820);
or U31653 (N_31653,N_30227,N_30850);
nand U31654 (N_31654,N_30873,N_30681);
nor U31655 (N_31655,N_30522,N_30386);
and U31656 (N_31656,N_30920,N_30996);
nand U31657 (N_31657,N_30158,N_30242);
and U31658 (N_31658,N_30934,N_30026);
nor U31659 (N_31659,N_30513,N_30344);
and U31660 (N_31660,N_30981,N_30071);
nor U31661 (N_31661,N_30862,N_30160);
nand U31662 (N_31662,N_30684,N_30309);
and U31663 (N_31663,N_30604,N_30175);
nor U31664 (N_31664,N_30583,N_30481);
and U31665 (N_31665,N_30832,N_30137);
or U31666 (N_31666,N_30559,N_30931);
xor U31667 (N_31667,N_30940,N_30619);
xnor U31668 (N_31668,N_30790,N_30419);
nor U31669 (N_31669,N_30593,N_30953);
and U31670 (N_31670,N_30174,N_30288);
xor U31671 (N_31671,N_30857,N_30012);
xor U31672 (N_31672,N_30353,N_30077);
and U31673 (N_31673,N_30301,N_30230);
xor U31674 (N_31674,N_30053,N_30212);
and U31675 (N_31675,N_30454,N_30466);
xor U31676 (N_31676,N_30477,N_30084);
or U31677 (N_31677,N_30894,N_30918);
nor U31678 (N_31678,N_30101,N_30264);
nor U31679 (N_31679,N_30172,N_30534);
xnor U31680 (N_31680,N_30641,N_30199);
xor U31681 (N_31681,N_30004,N_30793);
or U31682 (N_31682,N_30415,N_30871);
or U31683 (N_31683,N_30387,N_30176);
nand U31684 (N_31684,N_30366,N_30368);
or U31685 (N_31685,N_30471,N_30563);
nor U31686 (N_31686,N_30101,N_30185);
and U31687 (N_31687,N_30660,N_30117);
and U31688 (N_31688,N_30390,N_30771);
or U31689 (N_31689,N_30676,N_30160);
and U31690 (N_31690,N_30014,N_30059);
nand U31691 (N_31691,N_30495,N_30683);
nand U31692 (N_31692,N_30767,N_30457);
xnor U31693 (N_31693,N_30683,N_30608);
and U31694 (N_31694,N_30032,N_30770);
nor U31695 (N_31695,N_30305,N_30011);
or U31696 (N_31696,N_30543,N_30099);
or U31697 (N_31697,N_30541,N_30725);
xnor U31698 (N_31698,N_30845,N_30262);
and U31699 (N_31699,N_30332,N_30641);
nand U31700 (N_31700,N_30468,N_30640);
nor U31701 (N_31701,N_30031,N_30677);
nand U31702 (N_31702,N_30737,N_30873);
xnor U31703 (N_31703,N_30171,N_30773);
nand U31704 (N_31704,N_30527,N_30515);
nand U31705 (N_31705,N_30655,N_30994);
xnor U31706 (N_31706,N_30902,N_30898);
or U31707 (N_31707,N_30638,N_30100);
or U31708 (N_31708,N_30126,N_30335);
and U31709 (N_31709,N_30542,N_30597);
and U31710 (N_31710,N_30519,N_30620);
nand U31711 (N_31711,N_30744,N_30828);
and U31712 (N_31712,N_30528,N_30583);
nand U31713 (N_31713,N_30468,N_30341);
or U31714 (N_31714,N_30798,N_30676);
xnor U31715 (N_31715,N_30468,N_30087);
nand U31716 (N_31716,N_30290,N_30249);
nor U31717 (N_31717,N_30019,N_30205);
or U31718 (N_31718,N_30772,N_30721);
xor U31719 (N_31719,N_30265,N_30980);
or U31720 (N_31720,N_30534,N_30837);
xnor U31721 (N_31721,N_30483,N_30233);
nand U31722 (N_31722,N_30226,N_30207);
and U31723 (N_31723,N_30955,N_30493);
and U31724 (N_31724,N_30115,N_30895);
or U31725 (N_31725,N_30888,N_30988);
nor U31726 (N_31726,N_30164,N_30521);
xor U31727 (N_31727,N_30376,N_30067);
nor U31728 (N_31728,N_30190,N_30858);
nand U31729 (N_31729,N_30255,N_30758);
nor U31730 (N_31730,N_30142,N_30480);
and U31731 (N_31731,N_30102,N_30664);
nand U31732 (N_31732,N_30461,N_30977);
and U31733 (N_31733,N_30425,N_30806);
nor U31734 (N_31734,N_30401,N_30225);
and U31735 (N_31735,N_30777,N_30974);
nand U31736 (N_31736,N_30240,N_30447);
or U31737 (N_31737,N_30094,N_30795);
and U31738 (N_31738,N_30658,N_30435);
xnor U31739 (N_31739,N_30066,N_30969);
nor U31740 (N_31740,N_30992,N_30852);
nand U31741 (N_31741,N_30566,N_30532);
nor U31742 (N_31742,N_30523,N_30234);
or U31743 (N_31743,N_30677,N_30279);
nor U31744 (N_31744,N_30193,N_30474);
nor U31745 (N_31745,N_30703,N_30574);
xor U31746 (N_31746,N_30555,N_30839);
nand U31747 (N_31747,N_30653,N_30891);
nand U31748 (N_31748,N_30352,N_30602);
and U31749 (N_31749,N_30066,N_30350);
and U31750 (N_31750,N_30527,N_30083);
xnor U31751 (N_31751,N_30075,N_30562);
and U31752 (N_31752,N_30709,N_30692);
nor U31753 (N_31753,N_30964,N_30343);
or U31754 (N_31754,N_30976,N_30893);
and U31755 (N_31755,N_30250,N_30314);
nor U31756 (N_31756,N_30645,N_30011);
and U31757 (N_31757,N_30146,N_30040);
nand U31758 (N_31758,N_30102,N_30500);
nand U31759 (N_31759,N_30077,N_30573);
or U31760 (N_31760,N_30894,N_30293);
or U31761 (N_31761,N_30871,N_30515);
and U31762 (N_31762,N_30965,N_30691);
nand U31763 (N_31763,N_30135,N_30253);
and U31764 (N_31764,N_30371,N_30549);
nor U31765 (N_31765,N_30690,N_30162);
or U31766 (N_31766,N_30722,N_30784);
nor U31767 (N_31767,N_30164,N_30891);
nor U31768 (N_31768,N_30794,N_30662);
nand U31769 (N_31769,N_30169,N_30761);
and U31770 (N_31770,N_30492,N_30201);
and U31771 (N_31771,N_30282,N_30963);
xnor U31772 (N_31772,N_30774,N_30850);
nand U31773 (N_31773,N_30240,N_30307);
nor U31774 (N_31774,N_30330,N_30724);
nand U31775 (N_31775,N_30467,N_30690);
nor U31776 (N_31776,N_30393,N_30993);
or U31777 (N_31777,N_30374,N_30996);
nand U31778 (N_31778,N_30787,N_30772);
nand U31779 (N_31779,N_30581,N_30967);
and U31780 (N_31780,N_30900,N_30581);
xnor U31781 (N_31781,N_30658,N_30588);
nand U31782 (N_31782,N_30270,N_30926);
or U31783 (N_31783,N_30062,N_30066);
xnor U31784 (N_31784,N_30878,N_30237);
nand U31785 (N_31785,N_30346,N_30813);
xor U31786 (N_31786,N_30054,N_30299);
and U31787 (N_31787,N_30085,N_30055);
nor U31788 (N_31788,N_30123,N_30811);
xor U31789 (N_31789,N_30991,N_30610);
and U31790 (N_31790,N_30216,N_30392);
nor U31791 (N_31791,N_30785,N_30673);
nand U31792 (N_31792,N_30527,N_30847);
or U31793 (N_31793,N_30040,N_30724);
and U31794 (N_31794,N_30196,N_30638);
nor U31795 (N_31795,N_30491,N_30297);
nor U31796 (N_31796,N_30657,N_30379);
and U31797 (N_31797,N_30694,N_30347);
nor U31798 (N_31798,N_30812,N_30280);
nor U31799 (N_31799,N_30194,N_30751);
nor U31800 (N_31800,N_30076,N_30658);
nand U31801 (N_31801,N_30680,N_30926);
nand U31802 (N_31802,N_30359,N_30175);
and U31803 (N_31803,N_30536,N_30223);
nand U31804 (N_31804,N_30363,N_30344);
nor U31805 (N_31805,N_30483,N_30958);
and U31806 (N_31806,N_30185,N_30514);
and U31807 (N_31807,N_30409,N_30665);
xor U31808 (N_31808,N_30959,N_30249);
nand U31809 (N_31809,N_30856,N_30281);
and U31810 (N_31810,N_30401,N_30325);
xor U31811 (N_31811,N_30821,N_30632);
nor U31812 (N_31812,N_30934,N_30109);
xor U31813 (N_31813,N_30404,N_30087);
nor U31814 (N_31814,N_30519,N_30432);
xor U31815 (N_31815,N_30724,N_30969);
nor U31816 (N_31816,N_30205,N_30207);
or U31817 (N_31817,N_30759,N_30235);
nand U31818 (N_31818,N_30283,N_30959);
xnor U31819 (N_31819,N_30180,N_30019);
xor U31820 (N_31820,N_30069,N_30573);
and U31821 (N_31821,N_30449,N_30719);
or U31822 (N_31822,N_30412,N_30034);
xnor U31823 (N_31823,N_30395,N_30192);
xor U31824 (N_31824,N_30107,N_30261);
or U31825 (N_31825,N_30143,N_30400);
nor U31826 (N_31826,N_30346,N_30515);
nand U31827 (N_31827,N_30708,N_30943);
xor U31828 (N_31828,N_30752,N_30333);
or U31829 (N_31829,N_30354,N_30521);
nand U31830 (N_31830,N_30536,N_30216);
nand U31831 (N_31831,N_30251,N_30026);
nand U31832 (N_31832,N_30869,N_30476);
xnor U31833 (N_31833,N_30405,N_30715);
xor U31834 (N_31834,N_30447,N_30564);
and U31835 (N_31835,N_30299,N_30443);
and U31836 (N_31836,N_30282,N_30693);
and U31837 (N_31837,N_30471,N_30346);
nand U31838 (N_31838,N_30754,N_30435);
nor U31839 (N_31839,N_30393,N_30805);
xor U31840 (N_31840,N_30544,N_30965);
xor U31841 (N_31841,N_30916,N_30244);
and U31842 (N_31842,N_30774,N_30822);
xnor U31843 (N_31843,N_30151,N_30174);
xor U31844 (N_31844,N_30313,N_30910);
or U31845 (N_31845,N_30150,N_30181);
nor U31846 (N_31846,N_30705,N_30582);
xor U31847 (N_31847,N_30575,N_30515);
and U31848 (N_31848,N_30273,N_30636);
or U31849 (N_31849,N_30542,N_30166);
nor U31850 (N_31850,N_30269,N_30291);
and U31851 (N_31851,N_30268,N_30025);
and U31852 (N_31852,N_30318,N_30072);
or U31853 (N_31853,N_30820,N_30142);
or U31854 (N_31854,N_30202,N_30788);
xnor U31855 (N_31855,N_30093,N_30998);
nand U31856 (N_31856,N_30490,N_30248);
nor U31857 (N_31857,N_30286,N_30040);
or U31858 (N_31858,N_30499,N_30237);
and U31859 (N_31859,N_30332,N_30101);
or U31860 (N_31860,N_30165,N_30898);
xor U31861 (N_31861,N_30217,N_30575);
nand U31862 (N_31862,N_30567,N_30280);
and U31863 (N_31863,N_30898,N_30535);
and U31864 (N_31864,N_30705,N_30497);
xnor U31865 (N_31865,N_30655,N_30147);
or U31866 (N_31866,N_30368,N_30659);
and U31867 (N_31867,N_30181,N_30076);
nor U31868 (N_31868,N_30571,N_30398);
xnor U31869 (N_31869,N_30451,N_30329);
and U31870 (N_31870,N_30801,N_30213);
nor U31871 (N_31871,N_30380,N_30683);
or U31872 (N_31872,N_30454,N_30040);
and U31873 (N_31873,N_30302,N_30223);
or U31874 (N_31874,N_30401,N_30177);
nand U31875 (N_31875,N_30120,N_30807);
xnor U31876 (N_31876,N_30172,N_30345);
xor U31877 (N_31877,N_30432,N_30504);
xor U31878 (N_31878,N_30401,N_30550);
or U31879 (N_31879,N_30631,N_30328);
nand U31880 (N_31880,N_30330,N_30782);
nand U31881 (N_31881,N_30206,N_30251);
nand U31882 (N_31882,N_30319,N_30368);
and U31883 (N_31883,N_30495,N_30031);
xor U31884 (N_31884,N_30150,N_30063);
and U31885 (N_31885,N_30546,N_30157);
nand U31886 (N_31886,N_30978,N_30001);
nor U31887 (N_31887,N_30586,N_30041);
xor U31888 (N_31888,N_30535,N_30410);
nand U31889 (N_31889,N_30039,N_30749);
nand U31890 (N_31890,N_30839,N_30424);
xor U31891 (N_31891,N_30038,N_30170);
or U31892 (N_31892,N_30196,N_30683);
nor U31893 (N_31893,N_30576,N_30388);
nand U31894 (N_31894,N_30120,N_30575);
nor U31895 (N_31895,N_30657,N_30237);
nor U31896 (N_31896,N_30704,N_30563);
or U31897 (N_31897,N_30493,N_30887);
nand U31898 (N_31898,N_30870,N_30629);
nand U31899 (N_31899,N_30225,N_30254);
and U31900 (N_31900,N_30440,N_30814);
or U31901 (N_31901,N_30364,N_30106);
nand U31902 (N_31902,N_30780,N_30810);
nor U31903 (N_31903,N_30903,N_30078);
or U31904 (N_31904,N_30195,N_30144);
or U31905 (N_31905,N_30573,N_30425);
and U31906 (N_31906,N_30056,N_30573);
xor U31907 (N_31907,N_30995,N_30778);
nor U31908 (N_31908,N_30060,N_30995);
nand U31909 (N_31909,N_30046,N_30606);
nor U31910 (N_31910,N_30275,N_30203);
xnor U31911 (N_31911,N_30571,N_30640);
xnor U31912 (N_31912,N_30137,N_30583);
or U31913 (N_31913,N_30909,N_30971);
nor U31914 (N_31914,N_30361,N_30762);
and U31915 (N_31915,N_30917,N_30906);
nand U31916 (N_31916,N_30696,N_30172);
xnor U31917 (N_31917,N_30612,N_30547);
or U31918 (N_31918,N_30791,N_30380);
xor U31919 (N_31919,N_30568,N_30016);
xor U31920 (N_31920,N_30431,N_30389);
nor U31921 (N_31921,N_30075,N_30162);
xor U31922 (N_31922,N_30089,N_30577);
nand U31923 (N_31923,N_30790,N_30060);
xnor U31924 (N_31924,N_30375,N_30643);
nand U31925 (N_31925,N_30118,N_30942);
xnor U31926 (N_31926,N_30286,N_30589);
nand U31927 (N_31927,N_30447,N_30856);
nor U31928 (N_31928,N_30093,N_30558);
or U31929 (N_31929,N_30612,N_30673);
xor U31930 (N_31930,N_30153,N_30194);
nand U31931 (N_31931,N_30170,N_30888);
nor U31932 (N_31932,N_30361,N_30501);
and U31933 (N_31933,N_30142,N_30160);
nor U31934 (N_31934,N_30054,N_30303);
or U31935 (N_31935,N_30613,N_30375);
nand U31936 (N_31936,N_30460,N_30430);
and U31937 (N_31937,N_30659,N_30685);
and U31938 (N_31938,N_30885,N_30810);
and U31939 (N_31939,N_30669,N_30847);
xnor U31940 (N_31940,N_30699,N_30337);
or U31941 (N_31941,N_30442,N_30666);
or U31942 (N_31942,N_30718,N_30404);
nor U31943 (N_31943,N_30443,N_30033);
nand U31944 (N_31944,N_30877,N_30374);
nand U31945 (N_31945,N_30397,N_30269);
nand U31946 (N_31946,N_30134,N_30884);
nand U31947 (N_31947,N_30264,N_30407);
nor U31948 (N_31948,N_30732,N_30269);
nor U31949 (N_31949,N_30356,N_30651);
and U31950 (N_31950,N_30539,N_30926);
nand U31951 (N_31951,N_30276,N_30447);
nor U31952 (N_31952,N_30983,N_30328);
or U31953 (N_31953,N_30633,N_30624);
nor U31954 (N_31954,N_30589,N_30751);
xnor U31955 (N_31955,N_30603,N_30755);
and U31956 (N_31956,N_30380,N_30039);
xor U31957 (N_31957,N_30547,N_30209);
or U31958 (N_31958,N_30823,N_30724);
or U31959 (N_31959,N_30502,N_30680);
and U31960 (N_31960,N_30984,N_30401);
xor U31961 (N_31961,N_30529,N_30836);
nor U31962 (N_31962,N_30212,N_30282);
and U31963 (N_31963,N_30719,N_30967);
or U31964 (N_31964,N_30696,N_30689);
nand U31965 (N_31965,N_30312,N_30958);
and U31966 (N_31966,N_30192,N_30900);
xnor U31967 (N_31967,N_30452,N_30198);
xor U31968 (N_31968,N_30241,N_30585);
nand U31969 (N_31969,N_30261,N_30302);
nor U31970 (N_31970,N_30061,N_30917);
nand U31971 (N_31971,N_30706,N_30116);
xnor U31972 (N_31972,N_30667,N_30697);
nor U31973 (N_31973,N_30957,N_30777);
or U31974 (N_31974,N_30536,N_30400);
and U31975 (N_31975,N_30807,N_30461);
nand U31976 (N_31976,N_30145,N_30419);
and U31977 (N_31977,N_30147,N_30411);
or U31978 (N_31978,N_30690,N_30991);
and U31979 (N_31979,N_30277,N_30570);
xnor U31980 (N_31980,N_30298,N_30860);
nand U31981 (N_31981,N_30807,N_30921);
or U31982 (N_31982,N_30587,N_30726);
or U31983 (N_31983,N_30042,N_30242);
and U31984 (N_31984,N_30207,N_30640);
xor U31985 (N_31985,N_30461,N_30374);
xnor U31986 (N_31986,N_30514,N_30542);
or U31987 (N_31987,N_30417,N_30269);
or U31988 (N_31988,N_30593,N_30201);
nor U31989 (N_31989,N_30955,N_30928);
nor U31990 (N_31990,N_30572,N_30182);
nand U31991 (N_31991,N_30172,N_30455);
nand U31992 (N_31992,N_30403,N_30636);
or U31993 (N_31993,N_30537,N_30018);
nor U31994 (N_31994,N_30258,N_30359);
xnor U31995 (N_31995,N_30124,N_30217);
nor U31996 (N_31996,N_30840,N_30185);
or U31997 (N_31997,N_30639,N_30391);
nand U31998 (N_31998,N_30538,N_30849);
xnor U31999 (N_31999,N_30513,N_30349);
xnor U32000 (N_32000,N_31409,N_31501);
and U32001 (N_32001,N_31292,N_31059);
nand U32002 (N_32002,N_31421,N_31634);
or U32003 (N_32003,N_31946,N_31106);
nor U32004 (N_32004,N_31325,N_31701);
and U32005 (N_32005,N_31670,N_31854);
nor U32006 (N_32006,N_31636,N_31151);
and U32007 (N_32007,N_31852,N_31224);
xor U32008 (N_32008,N_31276,N_31211);
nand U32009 (N_32009,N_31690,N_31268);
or U32010 (N_32010,N_31872,N_31991);
or U32011 (N_32011,N_31291,N_31715);
and U32012 (N_32012,N_31627,N_31047);
xor U32013 (N_32013,N_31078,N_31924);
nor U32014 (N_32014,N_31046,N_31316);
xnor U32015 (N_32015,N_31411,N_31708);
xor U32016 (N_32016,N_31179,N_31040);
and U32017 (N_32017,N_31109,N_31076);
nor U32018 (N_32018,N_31776,N_31940);
and U32019 (N_32019,N_31504,N_31485);
xnor U32020 (N_32020,N_31720,N_31650);
and U32021 (N_32021,N_31741,N_31279);
or U32022 (N_32022,N_31365,N_31738);
and U32023 (N_32023,N_31370,N_31631);
or U32024 (N_32024,N_31261,N_31937);
nand U32025 (N_32025,N_31867,N_31577);
or U32026 (N_32026,N_31336,N_31287);
and U32027 (N_32027,N_31153,N_31586);
xor U32028 (N_32028,N_31055,N_31834);
or U32029 (N_32029,N_31551,N_31380);
and U32030 (N_32030,N_31263,N_31548);
or U32031 (N_32031,N_31319,N_31123);
or U32032 (N_32032,N_31964,N_31234);
nor U32033 (N_32033,N_31328,N_31420);
nor U32034 (N_32034,N_31172,N_31133);
xnor U32035 (N_32035,N_31379,N_31466);
and U32036 (N_32036,N_31502,N_31803);
nand U32037 (N_32037,N_31677,N_31347);
and U32038 (N_32038,N_31828,N_31041);
nand U32039 (N_32039,N_31663,N_31910);
or U32040 (N_32040,N_31148,N_31248);
and U32041 (N_32041,N_31724,N_31626);
nand U32042 (N_32042,N_31657,N_31290);
or U32043 (N_32043,N_31825,N_31064);
or U32044 (N_32044,N_31275,N_31077);
or U32045 (N_32045,N_31968,N_31700);
nor U32046 (N_32046,N_31898,N_31798);
nor U32047 (N_32047,N_31402,N_31001);
or U32048 (N_32048,N_31090,N_31449);
or U32049 (N_32049,N_31437,N_31547);
nor U32050 (N_32050,N_31945,N_31288);
or U32051 (N_32051,N_31418,N_31923);
nor U32052 (N_32052,N_31166,N_31095);
and U32053 (N_32053,N_31598,N_31373);
and U32054 (N_32054,N_31213,N_31374);
and U32055 (N_32055,N_31596,N_31870);
nand U32056 (N_32056,N_31809,N_31761);
xnor U32057 (N_32057,N_31416,N_31031);
nand U32058 (N_32058,N_31085,N_31399);
nand U32059 (N_32059,N_31160,N_31388);
nand U32060 (N_32060,N_31578,N_31882);
and U32061 (N_32061,N_31887,N_31120);
xor U32062 (N_32062,N_31661,N_31891);
nor U32063 (N_32063,N_31537,N_31030);
nand U32064 (N_32064,N_31916,N_31067);
and U32065 (N_32065,N_31450,N_31550);
nor U32066 (N_32066,N_31920,N_31839);
nor U32067 (N_32067,N_31136,N_31233);
nor U32068 (N_32068,N_31855,N_31110);
or U32069 (N_32069,N_31829,N_31199);
nand U32070 (N_32070,N_31338,N_31235);
and U32071 (N_32071,N_31405,N_31403);
or U32072 (N_32072,N_31036,N_31394);
and U32073 (N_32073,N_31823,N_31592);
xor U32074 (N_32074,N_31771,N_31125);
xnor U32075 (N_32075,N_31264,N_31396);
nor U32076 (N_32076,N_31746,N_31518);
nor U32077 (N_32077,N_31245,N_31714);
and U32078 (N_32078,N_31807,N_31535);
and U32079 (N_32079,N_31323,N_31764);
and U32080 (N_32080,N_31591,N_31623);
nand U32081 (N_32081,N_31539,N_31000);
or U32082 (N_32082,N_31060,N_31772);
xnor U32083 (N_32083,N_31976,N_31143);
nor U32084 (N_32084,N_31800,N_31680);
nand U32085 (N_32085,N_31894,N_31579);
nand U32086 (N_32086,N_31628,N_31508);
nand U32087 (N_32087,N_31928,N_31258);
nand U32088 (N_32088,N_31020,N_31918);
nor U32089 (N_32089,N_31538,N_31357);
nor U32090 (N_32090,N_31666,N_31273);
nand U32091 (N_32091,N_31806,N_31557);
or U32092 (N_32092,N_31500,N_31297);
nor U32093 (N_32093,N_31671,N_31662);
nor U32094 (N_32094,N_31008,N_31640);
xor U32095 (N_32095,N_31089,N_31312);
nor U32096 (N_32096,N_31072,N_31289);
and U32097 (N_32097,N_31451,N_31257);
xor U32098 (N_32098,N_31564,N_31683);
xnor U32099 (N_32099,N_31185,N_31952);
and U32100 (N_32100,N_31102,N_31146);
nor U32101 (N_32101,N_31897,N_31641);
nand U32102 (N_32102,N_31304,N_31607);
nor U32103 (N_32103,N_31124,N_31006);
xnor U32104 (N_32104,N_31423,N_31506);
nand U32105 (N_32105,N_31818,N_31408);
nor U32106 (N_32106,N_31785,N_31345);
and U32107 (N_32107,N_31997,N_31027);
xor U32108 (N_32108,N_31175,N_31050);
or U32109 (N_32109,N_31063,N_31226);
and U32110 (N_32110,N_31303,N_31676);
and U32111 (N_32111,N_31011,N_31082);
xnor U32112 (N_32112,N_31385,N_31620);
or U32113 (N_32113,N_31361,N_31053);
and U32114 (N_32114,N_31138,N_31885);
and U32115 (N_32115,N_31673,N_31232);
nand U32116 (N_32116,N_31843,N_31019);
nand U32117 (N_32117,N_31993,N_31957);
nor U32118 (N_32118,N_31757,N_31206);
nand U32119 (N_32119,N_31313,N_31498);
and U32120 (N_32120,N_31962,N_31567);
xnor U32121 (N_32121,N_31249,N_31824);
nand U32122 (N_32122,N_31811,N_31490);
nor U32123 (N_32123,N_31941,N_31225);
or U32124 (N_32124,N_31159,N_31516);
or U32125 (N_32125,N_31194,N_31695);
or U32126 (N_32126,N_31719,N_31472);
nand U32127 (N_32127,N_31187,N_31271);
and U32128 (N_32128,N_31530,N_31058);
xnor U32129 (N_32129,N_31049,N_31333);
nand U32130 (N_32130,N_31010,N_31381);
or U32131 (N_32131,N_31349,N_31474);
nand U32132 (N_32132,N_31461,N_31477);
nand U32133 (N_32133,N_31644,N_31096);
and U32134 (N_32134,N_31180,N_31559);
nor U32135 (N_32135,N_31802,N_31355);
nand U32136 (N_32136,N_31066,N_31992);
and U32137 (N_32137,N_31728,N_31025);
and U32138 (N_32138,N_31083,N_31286);
nor U32139 (N_32139,N_31014,N_31996);
or U32140 (N_32140,N_31699,N_31778);
nor U32141 (N_32141,N_31201,N_31116);
xor U32142 (N_32142,N_31588,N_31927);
xor U32143 (N_32143,N_31848,N_31751);
nor U32144 (N_32144,N_31652,N_31979);
or U32145 (N_32145,N_31520,N_31269);
and U32146 (N_32146,N_31955,N_31471);
xnor U32147 (N_32147,N_31963,N_31605);
and U32148 (N_32148,N_31200,N_31004);
and U32149 (N_32149,N_31118,N_31780);
nand U32150 (N_32150,N_31513,N_31075);
and U32151 (N_32151,N_31722,N_31071);
or U32152 (N_32152,N_31913,N_31415);
or U32153 (N_32153,N_31054,N_31481);
nand U32154 (N_32154,N_31158,N_31429);
nand U32155 (N_32155,N_31658,N_31308);
xor U32156 (N_32156,N_31984,N_31922);
nor U32157 (N_32157,N_31101,N_31509);
nand U32158 (N_32158,N_31721,N_31822);
and U32159 (N_32159,N_31087,N_31540);
xnor U32160 (N_32160,N_31468,N_31853);
or U32161 (N_32161,N_31703,N_31723);
and U32162 (N_32162,N_31487,N_31895);
nand U32163 (N_32163,N_31545,N_31947);
xor U32164 (N_32164,N_31122,N_31599);
or U32165 (N_32165,N_31743,N_31042);
nor U32166 (N_32166,N_31524,N_31901);
nand U32167 (N_32167,N_31759,N_31917);
xor U32168 (N_32168,N_31285,N_31262);
and U32169 (N_32169,N_31103,N_31305);
and U32170 (N_32170,N_31007,N_31278);
nor U32171 (N_32171,N_31189,N_31549);
nand U32172 (N_32172,N_31028,N_31121);
nor U32173 (N_32173,N_31961,N_31478);
or U32174 (N_32174,N_31888,N_31018);
nor U32175 (N_32175,N_31654,N_31284);
xnor U32176 (N_32176,N_31614,N_31243);
and U32177 (N_32177,N_31616,N_31817);
nand U32178 (N_32178,N_31613,N_31919);
nand U32179 (N_32179,N_31390,N_31130);
nand U32180 (N_32180,N_31162,N_31622);
or U32181 (N_32181,N_31765,N_31184);
or U32182 (N_32182,N_31340,N_31583);
nor U32183 (N_32183,N_31003,N_31251);
and U32184 (N_32184,N_31117,N_31978);
and U32185 (N_32185,N_31088,N_31600);
or U32186 (N_32186,N_31793,N_31283);
nand U32187 (N_32187,N_31427,N_31845);
nor U32188 (N_32188,N_31821,N_31711);
and U32189 (N_32189,N_31507,N_31925);
nor U32190 (N_32190,N_31202,N_31188);
xnor U32191 (N_32191,N_31590,N_31197);
nand U32192 (N_32192,N_31755,N_31575);
nand U32193 (N_32193,N_31309,N_31944);
xor U32194 (N_32194,N_31029,N_31618);
nor U32195 (N_32195,N_31371,N_31942);
xor U32196 (N_32196,N_31983,N_31352);
or U32197 (N_32197,N_31782,N_31306);
nand U32198 (N_32198,N_31543,N_31051);
nand U32199 (N_32199,N_31182,N_31424);
xor U32200 (N_32200,N_31856,N_31367);
xnor U32201 (N_32201,N_31002,N_31015);
nor U32202 (N_32202,N_31445,N_31168);
nor U32203 (N_32203,N_31070,N_31198);
xor U32204 (N_32204,N_31154,N_31229);
nand U32205 (N_32205,N_31685,N_31382);
xnor U32206 (N_32206,N_31369,N_31769);
or U32207 (N_32207,N_31998,N_31387);
nor U32208 (N_32208,N_31649,N_31929);
xnor U32209 (N_32209,N_31630,N_31960);
or U32210 (N_32210,N_31497,N_31208);
and U32211 (N_32211,N_31482,N_31861);
nor U32212 (N_32212,N_31838,N_31938);
and U32213 (N_32213,N_31820,N_31740);
nand U32214 (N_32214,N_31805,N_31858);
or U32215 (N_32215,N_31165,N_31943);
nand U32216 (N_32216,N_31274,N_31260);
nand U32217 (N_32217,N_31163,N_31692);
xor U32218 (N_32218,N_31904,N_31791);
xor U32219 (N_32219,N_31204,N_31989);
nand U32220 (N_32220,N_31486,N_31433);
or U32221 (N_32221,N_31693,N_31127);
or U32222 (N_32222,N_31637,N_31364);
xor U32223 (N_32223,N_31859,N_31376);
xnor U32224 (N_32224,N_31344,N_31439);
or U32225 (N_32225,N_31298,N_31032);
xor U32226 (N_32226,N_31866,N_31568);
nor U32227 (N_32227,N_31391,N_31026);
nand U32228 (N_32228,N_31280,N_31679);
xnor U32229 (N_32229,N_31813,N_31748);
nor U32230 (N_32230,N_31282,N_31569);
or U32231 (N_32231,N_31021,N_31558);
xor U32232 (N_32232,N_31531,N_31745);
nand U32233 (N_32233,N_31664,N_31300);
nor U32234 (N_32234,N_31544,N_31571);
nand U32235 (N_32235,N_31022,N_31868);
or U32236 (N_32236,N_31436,N_31880);
and U32237 (N_32237,N_31886,N_31762);
nand U32238 (N_32238,N_31536,N_31012);
nand U32239 (N_32239,N_31476,N_31737);
xnor U32240 (N_32240,N_31645,N_31959);
nand U32241 (N_32241,N_31212,N_31646);
nand U32242 (N_32242,N_31191,N_31656);
nand U32243 (N_32243,N_31327,N_31384);
nand U32244 (N_32244,N_31086,N_31389);
and U32245 (N_32245,N_31203,N_31563);
nand U32246 (N_32246,N_31758,N_31024);
or U32247 (N_32247,N_31410,N_31255);
nor U32248 (N_32248,N_31186,N_31768);
nand U32249 (N_32249,N_31417,N_31176);
and U32250 (N_32250,N_31625,N_31013);
nor U32251 (N_32251,N_31438,N_31747);
nor U32252 (N_32252,N_31425,N_31183);
and U32253 (N_32253,N_31844,N_31266);
xnor U32254 (N_32254,N_31665,N_31602);
nand U32255 (N_32255,N_31157,N_31145);
nand U32256 (N_32256,N_31794,N_31035);
nand U32257 (N_32257,N_31840,N_31799);
and U32258 (N_32258,N_31753,N_31893);
or U32259 (N_32259,N_31210,N_31643);
and U32260 (N_32260,N_31359,N_31113);
nand U32261 (N_32261,N_31763,N_31911);
nand U32262 (N_32262,N_31244,N_31601);
and U32263 (N_32263,N_31585,N_31068);
or U32264 (N_32264,N_31847,N_31986);
nand U32265 (N_32265,N_31104,N_31447);
or U32266 (N_32266,N_31883,N_31108);
and U32267 (N_32267,N_31881,N_31404);
nand U32268 (N_32268,N_31038,N_31463);
nand U32269 (N_32269,N_31242,N_31589);
and U32270 (N_32270,N_31267,N_31080);
and U32271 (N_32271,N_31149,N_31494);
xnor U32272 (N_32272,N_31915,N_31775);
xnor U32273 (N_32273,N_31732,N_31256);
and U32274 (N_32274,N_31808,N_31231);
nor U32275 (N_32275,N_31749,N_31648);
or U32276 (N_32276,N_31353,N_31796);
nor U32277 (N_32277,N_31496,N_31810);
nor U32278 (N_32278,N_31057,N_31062);
and U32279 (N_32279,N_31238,N_31519);
nor U32280 (N_32280,N_31045,N_31801);
nand U32281 (N_32281,N_31152,N_31326);
nand U32282 (N_32282,N_31977,N_31773);
nor U32283 (N_32283,N_31668,N_31522);
and U32284 (N_32284,N_31639,N_31691);
xnor U32285 (N_32285,N_31346,N_31573);
xnor U32286 (N_32286,N_31005,N_31223);
nand U32287 (N_32287,N_31967,N_31039);
or U32288 (N_32288,N_31546,N_31167);
nand U32289 (N_32289,N_31097,N_31294);
xor U32290 (N_32290,N_31147,N_31383);
or U32291 (N_32291,N_31735,N_31609);
or U32292 (N_32292,N_31674,N_31056);
nand U32293 (N_32293,N_31980,N_31324);
and U32294 (N_32294,N_31532,N_31492);
nor U32295 (N_32295,N_31552,N_31726);
and U32296 (N_32296,N_31851,N_31190);
or U32297 (N_32297,N_31119,N_31457);
or U32298 (N_32298,N_31788,N_31841);
or U32299 (N_32299,N_31037,N_31017);
xor U32300 (N_32300,N_31862,N_31156);
nand U32301 (N_32301,N_31315,N_31831);
or U32302 (N_32302,N_31906,N_31554);
nor U32303 (N_32303,N_31687,N_31842);
nor U32304 (N_32304,N_31595,N_31479);
xnor U32305 (N_32305,N_31608,N_31395);
nand U32306 (N_32306,N_31678,N_31016);
nor U32307 (N_32307,N_31277,N_31815);
and U32308 (N_32308,N_31227,N_31217);
xnor U32309 (N_32309,N_31562,N_31716);
nand U32310 (N_32310,N_31533,N_31576);
nand U32311 (N_32311,N_31816,N_31455);
nor U32312 (N_32312,N_31733,N_31896);
nand U32313 (N_32313,N_31555,N_31128);
nor U32314 (N_32314,N_31849,N_31434);
and U32315 (N_32315,N_31704,N_31393);
and U32316 (N_32316,N_31511,N_31754);
and U32317 (N_32317,N_31875,N_31871);
or U32318 (N_32318,N_31480,N_31675);
nand U32319 (N_32319,N_31440,N_31899);
nand U32320 (N_32320,N_31081,N_31990);
or U32321 (N_32321,N_31459,N_31632);
xnor U32322 (N_32322,N_31339,N_31669);
nand U32323 (N_32323,N_31193,N_31368);
and U32324 (N_32324,N_31079,N_31987);
xor U32325 (N_32325,N_31099,N_31933);
nor U32326 (N_32326,N_31322,N_31350);
and U32327 (N_32327,N_31836,N_31837);
nor U32328 (N_32328,N_31702,N_31334);
nor U32329 (N_32329,N_31651,N_31584);
nor U32330 (N_32330,N_31241,N_31023);
nand U32331 (N_32331,N_31752,N_31301);
nand U32332 (N_32332,N_31903,N_31401);
or U32333 (N_32333,N_31307,N_31454);
nand U32334 (N_32334,N_31570,N_31377);
or U32335 (N_32335,N_31864,N_31460);
xnor U32336 (N_32336,N_31797,N_31950);
nor U32337 (N_32337,N_31132,N_31850);
or U32338 (N_32338,N_31667,N_31706);
nand U32339 (N_32339,N_31239,N_31642);
or U32340 (N_32340,N_31553,N_31912);
or U32341 (N_32341,N_31982,N_31826);
nand U32342 (N_32342,N_31617,N_31879);
nor U32343 (N_32343,N_31698,N_31766);
and U32344 (N_32344,N_31452,N_31760);
xor U32345 (N_32345,N_31653,N_31742);
nand U32346 (N_32346,N_31150,N_31247);
and U32347 (N_32347,N_31342,N_31526);
nand U32348 (N_32348,N_31783,N_31510);
and U32349 (N_32349,N_31835,N_31320);
and U32350 (N_32350,N_31317,N_31865);
xor U32351 (N_32351,N_31140,N_31448);
xor U32352 (N_32352,N_31318,N_31932);
xor U32353 (N_32353,N_31216,N_31981);
and U32354 (N_32354,N_31612,N_31729);
xor U32355 (N_32355,N_31921,N_31604);
xor U32356 (N_32356,N_31362,N_31712);
nor U32357 (N_32357,N_31196,N_31270);
nand U32358 (N_32358,N_31954,N_31832);
or U32359 (N_32359,N_31787,N_31907);
nor U32360 (N_32360,N_31131,N_31970);
nor U32361 (N_32361,N_31694,N_31792);
or U32362 (N_32362,N_31725,N_31343);
and U32363 (N_32363,N_31582,N_31354);
nand U32364 (N_32364,N_31091,N_31112);
or U32365 (N_32365,N_31512,N_31375);
or U32366 (N_32366,N_31126,N_31739);
nor U32367 (N_32367,N_31556,N_31386);
and U32368 (N_32368,N_31443,N_31293);
nand U32369 (N_32369,N_31331,N_31100);
xnor U32370 (N_32370,N_31398,N_31734);
or U32371 (N_32371,N_31142,N_31515);
xor U32372 (N_32372,N_31422,N_31655);
nor U32373 (N_32373,N_31948,N_31250);
nand U32374 (N_32374,N_31905,N_31697);
nand U32375 (N_32375,N_31139,N_31804);
or U32376 (N_32376,N_31220,N_31337);
and U32377 (N_32377,N_31406,N_31169);
nand U32378 (N_32378,N_31135,N_31560);
and U32379 (N_32379,N_31467,N_31819);
xnor U32380 (N_32380,N_31988,N_31696);
or U32381 (N_32381,N_31884,N_31930);
nand U32382 (N_32382,N_31442,N_31446);
and U32383 (N_32383,N_31789,N_31428);
or U32384 (N_32384,N_31629,N_31876);
or U32385 (N_32385,N_31972,N_31470);
nand U32386 (N_32386,N_31974,N_31400);
nor U32387 (N_32387,N_31332,N_31624);
nand U32388 (N_32388,N_31495,N_31969);
or U32389 (N_32389,N_31936,N_31830);
nand U32390 (N_32390,N_31846,N_31814);
or U32391 (N_32391,N_31727,N_31863);
nor U32392 (N_32392,N_31253,N_31134);
and U32393 (N_32393,N_31709,N_31874);
or U32394 (N_32394,N_31052,N_31705);
nor U32395 (N_32395,N_31593,N_31195);
nor U32396 (N_32396,N_31061,N_31441);
and U32397 (N_32397,N_31392,N_31048);
or U32398 (N_32398,N_31218,N_31619);
nor U32399 (N_32399,N_31660,N_31574);
xnor U32400 (N_32400,N_31335,N_31431);
nand U32401 (N_32401,N_31141,N_31958);
or U32402 (N_32402,N_31935,N_31681);
nand U32403 (N_32403,N_31009,N_31784);
xor U32404 (N_32404,N_31397,N_31458);
xor U32405 (N_32405,N_31603,N_31860);
and U32406 (N_32406,N_31484,N_31228);
nor U32407 (N_32407,N_31222,N_31310);
xnor U32408 (N_32408,N_31908,N_31774);
nor U32409 (N_32409,N_31173,N_31372);
nand U32410 (N_32410,N_31833,N_31033);
and U32411 (N_32411,N_31174,N_31296);
xnor U32412 (N_32412,N_31230,N_31710);
and U32413 (N_32413,N_31951,N_31931);
xor U32414 (N_32414,N_31044,N_31523);
and U32415 (N_32415,N_31069,N_31580);
and U32416 (N_32416,N_31164,N_31985);
xor U32417 (N_32417,N_31129,N_31221);
xnor U32418 (N_32418,N_31462,N_31192);
xnor U32419 (N_32419,N_31246,N_31105);
xnor U32420 (N_32420,N_31566,N_31171);
xor U32421 (N_32421,N_31214,N_31178);
nor U32422 (N_32422,N_31857,N_31779);
xnor U32423 (N_32423,N_31065,N_31525);
or U32424 (N_32424,N_31426,N_31272);
and U32425 (N_32425,N_31956,N_31219);
or U32426 (N_32426,N_31366,N_31215);
nand U32427 (N_32427,N_31236,N_31561);
xnor U32428 (N_32428,N_31412,N_31529);
nor U32429 (N_32429,N_31254,N_31111);
xnor U32430 (N_32430,N_31647,N_31407);
nand U32431 (N_32431,N_31889,N_31786);
nor U32432 (N_32432,N_31378,N_31252);
or U32433 (N_32433,N_31517,N_31456);
nand U32434 (N_32434,N_31767,N_31541);
or U32435 (N_32435,N_31348,N_31311);
or U32436 (N_32436,N_31170,N_31464);
xor U32437 (N_32437,N_31689,N_31034);
and U32438 (N_32438,N_31430,N_31092);
nand U32439 (N_32439,N_31939,N_31707);
nor U32440 (N_32440,N_31900,N_31084);
or U32441 (N_32441,N_31812,N_31505);
nand U32442 (N_32442,N_31621,N_31491);
and U32443 (N_32443,N_31902,N_31414);
nand U32444 (N_32444,N_31949,N_31750);
xnor U32445 (N_32445,N_31790,N_31107);
or U32446 (N_32446,N_31483,N_31493);
and U32447 (N_32447,N_31177,N_31299);
nand U32448 (N_32448,N_31975,N_31730);
or U32449 (N_32449,N_31144,N_31205);
nand U32450 (N_32450,N_31265,N_31360);
xnor U32451 (N_32451,N_31684,N_31594);
and U32452 (N_32452,N_31744,N_31314);
nand U32453 (N_32453,N_31419,N_31994);
or U32454 (N_32454,N_31686,N_31435);
nand U32455 (N_32455,N_31965,N_31770);
nor U32456 (N_32456,N_31953,N_31718);
and U32457 (N_32457,N_31971,N_31514);
nand U32458 (N_32458,N_31973,N_31873);
and U32459 (N_32459,N_31358,N_31475);
xnor U32460 (N_32460,N_31926,N_31713);
nor U32461 (N_32461,N_31638,N_31093);
and U32462 (N_32462,N_31363,N_31351);
nor U32463 (N_32463,N_31717,N_31503);
xor U32464 (N_32464,N_31521,N_31756);
xnor U32465 (N_32465,N_31469,N_31488);
and U32466 (N_32466,N_31413,N_31473);
or U32467 (N_32467,N_31073,N_31114);
xor U32468 (N_32468,N_31688,N_31682);
nor U32469 (N_32469,N_31909,N_31281);
nand U32470 (N_32470,N_31499,N_31736);
nand U32471 (N_32471,N_31161,N_31209);
xnor U32472 (N_32472,N_31934,N_31995);
and U32473 (N_32473,N_31615,N_31572);
nor U32474 (N_32474,N_31542,N_31356);
and U32475 (N_32475,N_31207,N_31259);
and U32476 (N_32476,N_31074,N_31043);
xnor U32477 (N_32477,N_31877,N_31295);
and U32478 (N_32478,N_31237,N_31528);
or U32479 (N_32479,N_31098,N_31890);
nand U32480 (N_32480,N_31330,N_31321);
nand U32481 (N_32481,N_31869,N_31795);
nor U32482 (N_32482,N_31606,N_31489);
and U32483 (N_32483,N_31094,N_31115);
xnor U32484 (N_32484,N_31155,N_31827);
or U32485 (N_32485,N_31181,N_31329);
or U32486 (N_32486,N_31611,N_31341);
and U32487 (N_32487,N_31777,N_31534);
or U32488 (N_32488,N_31781,N_31966);
and U32489 (N_32489,N_31610,N_31302);
xnor U32490 (N_32490,N_31565,N_31527);
and U32491 (N_32491,N_31914,N_31453);
and U32492 (N_32492,N_31465,N_31587);
nor U32493 (N_32493,N_31444,N_31581);
and U32494 (N_32494,N_31878,N_31240);
and U32495 (N_32495,N_31432,N_31659);
nor U32496 (N_32496,N_31597,N_31892);
xor U32497 (N_32497,N_31731,N_31999);
nand U32498 (N_32498,N_31672,N_31633);
and U32499 (N_32499,N_31137,N_31635);
or U32500 (N_32500,N_31752,N_31263);
nand U32501 (N_32501,N_31425,N_31923);
xor U32502 (N_32502,N_31704,N_31870);
xor U32503 (N_32503,N_31738,N_31338);
and U32504 (N_32504,N_31217,N_31900);
nor U32505 (N_32505,N_31571,N_31051);
and U32506 (N_32506,N_31464,N_31573);
and U32507 (N_32507,N_31074,N_31206);
nor U32508 (N_32508,N_31918,N_31946);
nor U32509 (N_32509,N_31366,N_31598);
nand U32510 (N_32510,N_31337,N_31140);
nand U32511 (N_32511,N_31737,N_31444);
or U32512 (N_32512,N_31103,N_31727);
nor U32513 (N_32513,N_31401,N_31620);
and U32514 (N_32514,N_31413,N_31394);
and U32515 (N_32515,N_31108,N_31474);
and U32516 (N_32516,N_31709,N_31339);
xnor U32517 (N_32517,N_31719,N_31676);
or U32518 (N_32518,N_31186,N_31221);
nand U32519 (N_32519,N_31933,N_31079);
nor U32520 (N_32520,N_31248,N_31507);
xnor U32521 (N_32521,N_31594,N_31211);
or U32522 (N_32522,N_31795,N_31683);
or U32523 (N_32523,N_31407,N_31978);
nor U32524 (N_32524,N_31872,N_31190);
nor U32525 (N_32525,N_31986,N_31206);
xor U32526 (N_32526,N_31870,N_31720);
nor U32527 (N_32527,N_31367,N_31673);
xor U32528 (N_32528,N_31395,N_31331);
nand U32529 (N_32529,N_31051,N_31276);
nand U32530 (N_32530,N_31391,N_31181);
or U32531 (N_32531,N_31993,N_31497);
or U32532 (N_32532,N_31941,N_31794);
xor U32533 (N_32533,N_31846,N_31331);
nand U32534 (N_32534,N_31722,N_31135);
or U32535 (N_32535,N_31703,N_31762);
and U32536 (N_32536,N_31341,N_31948);
nand U32537 (N_32537,N_31168,N_31764);
and U32538 (N_32538,N_31323,N_31528);
xnor U32539 (N_32539,N_31289,N_31871);
and U32540 (N_32540,N_31166,N_31820);
xnor U32541 (N_32541,N_31848,N_31786);
and U32542 (N_32542,N_31319,N_31717);
nand U32543 (N_32543,N_31984,N_31328);
or U32544 (N_32544,N_31369,N_31692);
nand U32545 (N_32545,N_31522,N_31361);
and U32546 (N_32546,N_31715,N_31295);
nor U32547 (N_32547,N_31556,N_31137);
xor U32548 (N_32548,N_31551,N_31646);
and U32549 (N_32549,N_31818,N_31810);
nor U32550 (N_32550,N_31496,N_31867);
nor U32551 (N_32551,N_31278,N_31747);
nand U32552 (N_32552,N_31596,N_31334);
nand U32553 (N_32553,N_31043,N_31167);
and U32554 (N_32554,N_31948,N_31860);
and U32555 (N_32555,N_31158,N_31085);
xnor U32556 (N_32556,N_31253,N_31956);
or U32557 (N_32557,N_31943,N_31679);
nand U32558 (N_32558,N_31586,N_31147);
nand U32559 (N_32559,N_31337,N_31445);
nor U32560 (N_32560,N_31710,N_31273);
or U32561 (N_32561,N_31705,N_31256);
nor U32562 (N_32562,N_31076,N_31968);
nor U32563 (N_32563,N_31076,N_31241);
nor U32564 (N_32564,N_31297,N_31752);
nand U32565 (N_32565,N_31294,N_31987);
and U32566 (N_32566,N_31904,N_31289);
and U32567 (N_32567,N_31138,N_31359);
nand U32568 (N_32568,N_31108,N_31093);
nand U32569 (N_32569,N_31606,N_31027);
nor U32570 (N_32570,N_31829,N_31444);
nor U32571 (N_32571,N_31317,N_31854);
or U32572 (N_32572,N_31098,N_31892);
nor U32573 (N_32573,N_31436,N_31628);
nor U32574 (N_32574,N_31323,N_31767);
nand U32575 (N_32575,N_31601,N_31617);
nand U32576 (N_32576,N_31319,N_31674);
nor U32577 (N_32577,N_31138,N_31179);
xor U32578 (N_32578,N_31728,N_31988);
and U32579 (N_32579,N_31598,N_31678);
nand U32580 (N_32580,N_31893,N_31143);
xor U32581 (N_32581,N_31897,N_31723);
nor U32582 (N_32582,N_31322,N_31442);
nand U32583 (N_32583,N_31282,N_31096);
xnor U32584 (N_32584,N_31178,N_31222);
or U32585 (N_32585,N_31253,N_31498);
or U32586 (N_32586,N_31697,N_31551);
nand U32587 (N_32587,N_31074,N_31675);
nand U32588 (N_32588,N_31839,N_31024);
nor U32589 (N_32589,N_31470,N_31885);
xor U32590 (N_32590,N_31509,N_31387);
nand U32591 (N_32591,N_31058,N_31390);
and U32592 (N_32592,N_31045,N_31526);
xnor U32593 (N_32593,N_31208,N_31005);
and U32594 (N_32594,N_31360,N_31326);
nand U32595 (N_32595,N_31004,N_31769);
nand U32596 (N_32596,N_31715,N_31033);
and U32597 (N_32597,N_31048,N_31617);
nand U32598 (N_32598,N_31364,N_31981);
nor U32599 (N_32599,N_31484,N_31001);
nor U32600 (N_32600,N_31255,N_31546);
nor U32601 (N_32601,N_31729,N_31682);
nand U32602 (N_32602,N_31151,N_31114);
or U32603 (N_32603,N_31774,N_31514);
and U32604 (N_32604,N_31116,N_31866);
and U32605 (N_32605,N_31640,N_31802);
nand U32606 (N_32606,N_31008,N_31617);
and U32607 (N_32607,N_31141,N_31539);
nor U32608 (N_32608,N_31285,N_31539);
nor U32609 (N_32609,N_31789,N_31015);
nor U32610 (N_32610,N_31646,N_31074);
nor U32611 (N_32611,N_31802,N_31346);
and U32612 (N_32612,N_31666,N_31588);
or U32613 (N_32613,N_31223,N_31831);
nand U32614 (N_32614,N_31245,N_31112);
or U32615 (N_32615,N_31815,N_31667);
nor U32616 (N_32616,N_31709,N_31516);
nor U32617 (N_32617,N_31381,N_31528);
and U32618 (N_32618,N_31521,N_31137);
xor U32619 (N_32619,N_31277,N_31190);
and U32620 (N_32620,N_31484,N_31501);
nand U32621 (N_32621,N_31045,N_31590);
nor U32622 (N_32622,N_31049,N_31119);
nor U32623 (N_32623,N_31781,N_31525);
or U32624 (N_32624,N_31627,N_31106);
nand U32625 (N_32625,N_31497,N_31032);
nor U32626 (N_32626,N_31585,N_31807);
or U32627 (N_32627,N_31905,N_31544);
nand U32628 (N_32628,N_31577,N_31151);
or U32629 (N_32629,N_31304,N_31513);
or U32630 (N_32630,N_31547,N_31369);
and U32631 (N_32631,N_31190,N_31311);
or U32632 (N_32632,N_31067,N_31790);
or U32633 (N_32633,N_31984,N_31754);
or U32634 (N_32634,N_31449,N_31331);
nor U32635 (N_32635,N_31864,N_31372);
or U32636 (N_32636,N_31739,N_31956);
nor U32637 (N_32637,N_31619,N_31497);
nand U32638 (N_32638,N_31399,N_31890);
and U32639 (N_32639,N_31968,N_31850);
or U32640 (N_32640,N_31939,N_31909);
nor U32641 (N_32641,N_31558,N_31720);
or U32642 (N_32642,N_31227,N_31249);
nor U32643 (N_32643,N_31469,N_31498);
nor U32644 (N_32644,N_31854,N_31787);
or U32645 (N_32645,N_31170,N_31980);
nor U32646 (N_32646,N_31667,N_31198);
and U32647 (N_32647,N_31823,N_31466);
and U32648 (N_32648,N_31883,N_31583);
and U32649 (N_32649,N_31226,N_31464);
or U32650 (N_32650,N_31071,N_31198);
nand U32651 (N_32651,N_31831,N_31065);
xor U32652 (N_32652,N_31989,N_31947);
nor U32653 (N_32653,N_31911,N_31591);
or U32654 (N_32654,N_31621,N_31252);
nand U32655 (N_32655,N_31083,N_31260);
xnor U32656 (N_32656,N_31333,N_31384);
and U32657 (N_32657,N_31451,N_31389);
or U32658 (N_32658,N_31868,N_31061);
nand U32659 (N_32659,N_31840,N_31290);
or U32660 (N_32660,N_31349,N_31394);
or U32661 (N_32661,N_31045,N_31349);
xor U32662 (N_32662,N_31481,N_31628);
xor U32663 (N_32663,N_31515,N_31986);
and U32664 (N_32664,N_31697,N_31386);
and U32665 (N_32665,N_31495,N_31330);
xor U32666 (N_32666,N_31800,N_31561);
and U32667 (N_32667,N_31322,N_31206);
or U32668 (N_32668,N_31806,N_31050);
xnor U32669 (N_32669,N_31310,N_31978);
and U32670 (N_32670,N_31651,N_31094);
xor U32671 (N_32671,N_31612,N_31289);
nor U32672 (N_32672,N_31395,N_31521);
xnor U32673 (N_32673,N_31193,N_31161);
nand U32674 (N_32674,N_31474,N_31639);
xnor U32675 (N_32675,N_31882,N_31171);
nor U32676 (N_32676,N_31946,N_31786);
xor U32677 (N_32677,N_31570,N_31644);
nor U32678 (N_32678,N_31708,N_31630);
and U32679 (N_32679,N_31987,N_31124);
xnor U32680 (N_32680,N_31800,N_31056);
nand U32681 (N_32681,N_31679,N_31941);
xor U32682 (N_32682,N_31479,N_31693);
or U32683 (N_32683,N_31877,N_31856);
nand U32684 (N_32684,N_31820,N_31890);
nand U32685 (N_32685,N_31482,N_31765);
nand U32686 (N_32686,N_31587,N_31373);
or U32687 (N_32687,N_31125,N_31116);
or U32688 (N_32688,N_31477,N_31382);
xor U32689 (N_32689,N_31911,N_31513);
nor U32690 (N_32690,N_31366,N_31570);
or U32691 (N_32691,N_31250,N_31740);
and U32692 (N_32692,N_31582,N_31797);
nand U32693 (N_32693,N_31881,N_31297);
nand U32694 (N_32694,N_31118,N_31957);
nand U32695 (N_32695,N_31479,N_31916);
or U32696 (N_32696,N_31726,N_31088);
xnor U32697 (N_32697,N_31801,N_31872);
nor U32698 (N_32698,N_31965,N_31519);
nand U32699 (N_32699,N_31891,N_31199);
or U32700 (N_32700,N_31663,N_31307);
nor U32701 (N_32701,N_31884,N_31813);
xnor U32702 (N_32702,N_31882,N_31246);
nand U32703 (N_32703,N_31763,N_31772);
or U32704 (N_32704,N_31158,N_31020);
nor U32705 (N_32705,N_31526,N_31175);
xor U32706 (N_32706,N_31527,N_31168);
or U32707 (N_32707,N_31391,N_31790);
nand U32708 (N_32708,N_31221,N_31500);
nor U32709 (N_32709,N_31670,N_31047);
and U32710 (N_32710,N_31340,N_31379);
xor U32711 (N_32711,N_31983,N_31724);
and U32712 (N_32712,N_31095,N_31543);
nand U32713 (N_32713,N_31528,N_31836);
and U32714 (N_32714,N_31920,N_31996);
nor U32715 (N_32715,N_31670,N_31691);
and U32716 (N_32716,N_31151,N_31099);
or U32717 (N_32717,N_31132,N_31406);
nor U32718 (N_32718,N_31118,N_31817);
nand U32719 (N_32719,N_31915,N_31097);
nor U32720 (N_32720,N_31894,N_31782);
xor U32721 (N_32721,N_31779,N_31728);
or U32722 (N_32722,N_31060,N_31022);
or U32723 (N_32723,N_31833,N_31370);
and U32724 (N_32724,N_31233,N_31670);
or U32725 (N_32725,N_31824,N_31667);
nor U32726 (N_32726,N_31654,N_31269);
xnor U32727 (N_32727,N_31586,N_31095);
and U32728 (N_32728,N_31558,N_31354);
or U32729 (N_32729,N_31733,N_31035);
nand U32730 (N_32730,N_31305,N_31733);
xor U32731 (N_32731,N_31974,N_31010);
xor U32732 (N_32732,N_31288,N_31478);
xnor U32733 (N_32733,N_31940,N_31168);
xor U32734 (N_32734,N_31444,N_31471);
or U32735 (N_32735,N_31890,N_31781);
nor U32736 (N_32736,N_31324,N_31018);
nor U32737 (N_32737,N_31068,N_31623);
and U32738 (N_32738,N_31859,N_31348);
nand U32739 (N_32739,N_31863,N_31474);
xor U32740 (N_32740,N_31621,N_31000);
nand U32741 (N_32741,N_31189,N_31964);
and U32742 (N_32742,N_31738,N_31768);
nor U32743 (N_32743,N_31636,N_31010);
and U32744 (N_32744,N_31553,N_31762);
or U32745 (N_32745,N_31717,N_31462);
xor U32746 (N_32746,N_31174,N_31843);
nor U32747 (N_32747,N_31365,N_31772);
xor U32748 (N_32748,N_31128,N_31325);
nand U32749 (N_32749,N_31649,N_31751);
xor U32750 (N_32750,N_31809,N_31996);
or U32751 (N_32751,N_31877,N_31309);
nor U32752 (N_32752,N_31438,N_31288);
nand U32753 (N_32753,N_31610,N_31776);
and U32754 (N_32754,N_31473,N_31634);
and U32755 (N_32755,N_31756,N_31255);
nand U32756 (N_32756,N_31714,N_31738);
nor U32757 (N_32757,N_31105,N_31307);
or U32758 (N_32758,N_31021,N_31749);
or U32759 (N_32759,N_31131,N_31972);
and U32760 (N_32760,N_31969,N_31636);
xnor U32761 (N_32761,N_31481,N_31585);
nor U32762 (N_32762,N_31218,N_31417);
xor U32763 (N_32763,N_31358,N_31071);
xor U32764 (N_32764,N_31821,N_31478);
nand U32765 (N_32765,N_31365,N_31931);
or U32766 (N_32766,N_31113,N_31622);
and U32767 (N_32767,N_31150,N_31007);
and U32768 (N_32768,N_31304,N_31565);
nand U32769 (N_32769,N_31634,N_31295);
xor U32770 (N_32770,N_31109,N_31333);
xor U32771 (N_32771,N_31440,N_31461);
or U32772 (N_32772,N_31331,N_31324);
nand U32773 (N_32773,N_31009,N_31249);
and U32774 (N_32774,N_31212,N_31008);
or U32775 (N_32775,N_31118,N_31664);
nor U32776 (N_32776,N_31728,N_31406);
nand U32777 (N_32777,N_31464,N_31049);
nand U32778 (N_32778,N_31613,N_31525);
nand U32779 (N_32779,N_31703,N_31579);
nor U32780 (N_32780,N_31491,N_31603);
or U32781 (N_32781,N_31242,N_31132);
xnor U32782 (N_32782,N_31139,N_31305);
or U32783 (N_32783,N_31446,N_31545);
xor U32784 (N_32784,N_31848,N_31477);
or U32785 (N_32785,N_31202,N_31869);
nand U32786 (N_32786,N_31366,N_31563);
nand U32787 (N_32787,N_31610,N_31130);
nand U32788 (N_32788,N_31562,N_31816);
nor U32789 (N_32789,N_31458,N_31948);
or U32790 (N_32790,N_31676,N_31540);
nand U32791 (N_32791,N_31687,N_31120);
and U32792 (N_32792,N_31218,N_31492);
xor U32793 (N_32793,N_31309,N_31448);
or U32794 (N_32794,N_31188,N_31982);
nor U32795 (N_32795,N_31669,N_31488);
nor U32796 (N_32796,N_31551,N_31740);
xnor U32797 (N_32797,N_31967,N_31633);
nand U32798 (N_32798,N_31854,N_31819);
xor U32799 (N_32799,N_31887,N_31603);
or U32800 (N_32800,N_31115,N_31299);
nor U32801 (N_32801,N_31249,N_31286);
nor U32802 (N_32802,N_31792,N_31788);
nand U32803 (N_32803,N_31333,N_31140);
xnor U32804 (N_32804,N_31127,N_31541);
xnor U32805 (N_32805,N_31377,N_31023);
nor U32806 (N_32806,N_31397,N_31824);
and U32807 (N_32807,N_31360,N_31519);
xor U32808 (N_32808,N_31674,N_31120);
or U32809 (N_32809,N_31135,N_31048);
and U32810 (N_32810,N_31602,N_31254);
nand U32811 (N_32811,N_31224,N_31489);
or U32812 (N_32812,N_31587,N_31046);
and U32813 (N_32813,N_31066,N_31857);
nor U32814 (N_32814,N_31898,N_31502);
nor U32815 (N_32815,N_31756,N_31047);
and U32816 (N_32816,N_31395,N_31886);
or U32817 (N_32817,N_31180,N_31720);
or U32818 (N_32818,N_31705,N_31650);
nand U32819 (N_32819,N_31102,N_31860);
xnor U32820 (N_32820,N_31184,N_31923);
and U32821 (N_32821,N_31314,N_31972);
and U32822 (N_32822,N_31876,N_31697);
xor U32823 (N_32823,N_31801,N_31967);
xor U32824 (N_32824,N_31877,N_31698);
xnor U32825 (N_32825,N_31380,N_31750);
or U32826 (N_32826,N_31515,N_31327);
or U32827 (N_32827,N_31266,N_31905);
nand U32828 (N_32828,N_31111,N_31766);
or U32829 (N_32829,N_31326,N_31657);
xor U32830 (N_32830,N_31767,N_31364);
and U32831 (N_32831,N_31050,N_31311);
and U32832 (N_32832,N_31577,N_31349);
xor U32833 (N_32833,N_31335,N_31687);
nand U32834 (N_32834,N_31711,N_31314);
and U32835 (N_32835,N_31295,N_31110);
or U32836 (N_32836,N_31714,N_31152);
xor U32837 (N_32837,N_31084,N_31582);
nand U32838 (N_32838,N_31084,N_31168);
xor U32839 (N_32839,N_31630,N_31223);
or U32840 (N_32840,N_31678,N_31121);
nand U32841 (N_32841,N_31641,N_31720);
and U32842 (N_32842,N_31953,N_31615);
nor U32843 (N_32843,N_31218,N_31689);
and U32844 (N_32844,N_31934,N_31013);
nor U32845 (N_32845,N_31996,N_31204);
nand U32846 (N_32846,N_31176,N_31653);
and U32847 (N_32847,N_31646,N_31316);
xor U32848 (N_32848,N_31420,N_31362);
or U32849 (N_32849,N_31011,N_31017);
nand U32850 (N_32850,N_31471,N_31658);
nor U32851 (N_32851,N_31852,N_31893);
nand U32852 (N_32852,N_31507,N_31156);
and U32853 (N_32853,N_31837,N_31220);
and U32854 (N_32854,N_31850,N_31613);
nor U32855 (N_32855,N_31124,N_31506);
and U32856 (N_32856,N_31546,N_31497);
nor U32857 (N_32857,N_31780,N_31270);
or U32858 (N_32858,N_31902,N_31352);
nor U32859 (N_32859,N_31084,N_31394);
nand U32860 (N_32860,N_31388,N_31325);
or U32861 (N_32861,N_31138,N_31074);
or U32862 (N_32862,N_31878,N_31630);
xor U32863 (N_32863,N_31400,N_31297);
nand U32864 (N_32864,N_31366,N_31904);
xnor U32865 (N_32865,N_31107,N_31376);
xor U32866 (N_32866,N_31903,N_31426);
and U32867 (N_32867,N_31759,N_31744);
nand U32868 (N_32868,N_31826,N_31736);
and U32869 (N_32869,N_31036,N_31839);
or U32870 (N_32870,N_31329,N_31348);
and U32871 (N_32871,N_31092,N_31566);
nand U32872 (N_32872,N_31696,N_31251);
and U32873 (N_32873,N_31578,N_31989);
and U32874 (N_32874,N_31737,N_31230);
and U32875 (N_32875,N_31266,N_31719);
and U32876 (N_32876,N_31100,N_31361);
or U32877 (N_32877,N_31325,N_31151);
or U32878 (N_32878,N_31550,N_31387);
or U32879 (N_32879,N_31639,N_31526);
xor U32880 (N_32880,N_31177,N_31901);
and U32881 (N_32881,N_31491,N_31176);
and U32882 (N_32882,N_31555,N_31778);
xor U32883 (N_32883,N_31292,N_31827);
and U32884 (N_32884,N_31737,N_31225);
or U32885 (N_32885,N_31039,N_31493);
or U32886 (N_32886,N_31148,N_31371);
and U32887 (N_32887,N_31949,N_31135);
nor U32888 (N_32888,N_31832,N_31527);
and U32889 (N_32889,N_31564,N_31014);
nor U32890 (N_32890,N_31729,N_31396);
nand U32891 (N_32891,N_31045,N_31659);
or U32892 (N_32892,N_31603,N_31912);
nand U32893 (N_32893,N_31649,N_31529);
nor U32894 (N_32894,N_31370,N_31555);
nand U32895 (N_32895,N_31757,N_31325);
nand U32896 (N_32896,N_31309,N_31896);
xnor U32897 (N_32897,N_31711,N_31180);
nor U32898 (N_32898,N_31157,N_31864);
and U32899 (N_32899,N_31315,N_31492);
or U32900 (N_32900,N_31969,N_31097);
or U32901 (N_32901,N_31635,N_31271);
nor U32902 (N_32902,N_31559,N_31817);
nand U32903 (N_32903,N_31641,N_31340);
nor U32904 (N_32904,N_31675,N_31867);
nand U32905 (N_32905,N_31917,N_31424);
and U32906 (N_32906,N_31847,N_31880);
or U32907 (N_32907,N_31613,N_31596);
xnor U32908 (N_32908,N_31192,N_31028);
xor U32909 (N_32909,N_31853,N_31260);
or U32910 (N_32910,N_31589,N_31954);
xnor U32911 (N_32911,N_31373,N_31246);
nand U32912 (N_32912,N_31210,N_31510);
and U32913 (N_32913,N_31060,N_31827);
nand U32914 (N_32914,N_31109,N_31220);
nor U32915 (N_32915,N_31846,N_31159);
nor U32916 (N_32916,N_31382,N_31151);
nand U32917 (N_32917,N_31358,N_31394);
or U32918 (N_32918,N_31243,N_31546);
xnor U32919 (N_32919,N_31032,N_31248);
nor U32920 (N_32920,N_31965,N_31780);
or U32921 (N_32921,N_31033,N_31809);
xnor U32922 (N_32922,N_31738,N_31943);
or U32923 (N_32923,N_31507,N_31447);
or U32924 (N_32924,N_31998,N_31500);
and U32925 (N_32925,N_31282,N_31522);
xor U32926 (N_32926,N_31158,N_31493);
nand U32927 (N_32927,N_31997,N_31633);
xor U32928 (N_32928,N_31733,N_31940);
or U32929 (N_32929,N_31034,N_31035);
nand U32930 (N_32930,N_31461,N_31048);
xor U32931 (N_32931,N_31960,N_31985);
xnor U32932 (N_32932,N_31834,N_31929);
or U32933 (N_32933,N_31565,N_31139);
nor U32934 (N_32934,N_31912,N_31575);
and U32935 (N_32935,N_31359,N_31157);
or U32936 (N_32936,N_31905,N_31951);
or U32937 (N_32937,N_31535,N_31580);
nor U32938 (N_32938,N_31601,N_31147);
xor U32939 (N_32939,N_31889,N_31980);
xor U32940 (N_32940,N_31114,N_31149);
nor U32941 (N_32941,N_31356,N_31249);
nand U32942 (N_32942,N_31311,N_31768);
or U32943 (N_32943,N_31515,N_31107);
xnor U32944 (N_32944,N_31515,N_31122);
nand U32945 (N_32945,N_31513,N_31967);
nand U32946 (N_32946,N_31113,N_31234);
nor U32947 (N_32947,N_31741,N_31009);
or U32948 (N_32948,N_31567,N_31056);
or U32949 (N_32949,N_31594,N_31468);
nor U32950 (N_32950,N_31605,N_31933);
or U32951 (N_32951,N_31288,N_31472);
nand U32952 (N_32952,N_31717,N_31779);
and U32953 (N_32953,N_31880,N_31229);
nand U32954 (N_32954,N_31200,N_31746);
and U32955 (N_32955,N_31209,N_31477);
or U32956 (N_32956,N_31374,N_31910);
nor U32957 (N_32957,N_31881,N_31188);
nor U32958 (N_32958,N_31877,N_31071);
nor U32959 (N_32959,N_31615,N_31562);
or U32960 (N_32960,N_31617,N_31782);
nand U32961 (N_32961,N_31670,N_31595);
and U32962 (N_32962,N_31375,N_31069);
xnor U32963 (N_32963,N_31283,N_31499);
or U32964 (N_32964,N_31382,N_31927);
and U32965 (N_32965,N_31424,N_31302);
nor U32966 (N_32966,N_31155,N_31377);
nor U32967 (N_32967,N_31714,N_31203);
or U32968 (N_32968,N_31577,N_31120);
and U32969 (N_32969,N_31376,N_31349);
nor U32970 (N_32970,N_31413,N_31124);
nor U32971 (N_32971,N_31520,N_31379);
and U32972 (N_32972,N_31343,N_31754);
or U32973 (N_32973,N_31722,N_31073);
nor U32974 (N_32974,N_31442,N_31764);
xnor U32975 (N_32975,N_31136,N_31268);
xor U32976 (N_32976,N_31581,N_31831);
xor U32977 (N_32977,N_31506,N_31023);
and U32978 (N_32978,N_31853,N_31363);
nor U32979 (N_32979,N_31308,N_31635);
and U32980 (N_32980,N_31421,N_31066);
and U32981 (N_32981,N_31464,N_31984);
or U32982 (N_32982,N_31809,N_31739);
nand U32983 (N_32983,N_31139,N_31780);
and U32984 (N_32984,N_31257,N_31976);
nand U32985 (N_32985,N_31108,N_31388);
nand U32986 (N_32986,N_31622,N_31992);
or U32987 (N_32987,N_31218,N_31406);
xor U32988 (N_32988,N_31147,N_31984);
and U32989 (N_32989,N_31787,N_31598);
nand U32990 (N_32990,N_31119,N_31527);
nor U32991 (N_32991,N_31525,N_31850);
and U32992 (N_32992,N_31450,N_31761);
and U32993 (N_32993,N_31962,N_31213);
nand U32994 (N_32994,N_31217,N_31739);
or U32995 (N_32995,N_31297,N_31293);
nor U32996 (N_32996,N_31758,N_31046);
xnor U32997 (N_32997,N_31410,N_31180);
nor U32998 (N_32998,N_31142,N_31717);
nor U32999 (N_32999,N_31948,N_31515);
or U33000 (N_33000,N_32171,N_32956);
or U33001 (N_33001,N_32652,N_32976);
nand U33002 (N_33002,N_32418,N_32483);
nand U33003 (N_33003,N_32008,N_32580);
xor U33004 (N_33004,N_32472,N_32497);
nand U33005 (N_33005,N_32195,N_32366);
nand U33006 (N_33006,N_32522,N_32688);
nand U33007 (N_33007,N_32491,N_32760);
nand U33008 (N_33008,N_32124,N_32056);
or U33009 (N_33009,N_32602,N_32591);
or U33010 (N_33010,N_32889,N_32631);
nor U33011 (N_33011,N_32630,N_32009);
or U33012 (N_33012,N_32605,N_32334);
nor U33013 (N_33013,N_32044,N_32080);
xor U33014 (N_33014,N_32150,N_32979);
xnor U33015 (N_33015,N_32994,N_32802);
nand U33016 (N_33016,N_32675,N_32494);
nand U33017 (N_33017,N_32348,N_32679);
xor U33018 (N_33018,N_32232,N_32389);
nand U33019 (N_33019,N_32623,N_32779);
xor U33020 (N_33020,N_32249,N_32747);
and U33021 (N_33021,N_32162,N_32419);
and U33022 (N_33022,N_32699,N_32570);
nand U33023 (N_33023,N_32634,N_32545);
nand U33024 (N_33024,N_32191,N_32664);
nand U33025 (N_33025,N_32706,N_32731);
xnor U33026 (N_33026,N_32978,N_32531);
xnor U33027 (N_33027,N_32735,N_32135);
and U33028 (N_33028,N_32017,N_32678);
xnor U33029 (N_33029,N_32544,N_32982);
or U33030 (N_33030,N_32586,N_32256);
nor U33031 (N_33031,N_32159,N_32559);
or U33032 (N_33032,N_32416,N_32999);
xor U33033 (N_33033,N_32324,N_32733);
xor U33034 (N_33034,N_32556,N_32729);
or U33035 (N_33035,N_32975,N_32299);
xor U33036 (N_33036,N_32801,N_32661);
or U33037 (N_33037,N_32386,N_32702);
or U33038 (N_33038,N_32082,N_32873);
and U33039 (N_33039,N_32566,N_32629);
xnor U33040 (N_33040,N_32106,N_32149);
nor U33041 (N_33041,N_32202,N_32266);
nor U33042 (N_33042,N_32551,N_32073);
or U33043 (N_33043,N_32052,N_32216);
nor U33044 (N_33044,N_32786,N_32182);
and U33045 (N_33045,N_32144,N_32924);
and U33046 (N_33046,N_32697,N_32896);
or U33047 (N_33047,N_32774,N_32243);
nand U33048 (N_33048,N_32103,N_32504);
xor U33049 (N_33049,N_32248,N_32743);
nor U33050 (N_33050,N_32154,N_32604);
or U33051 (N_33051,N_32614,N_32961);
xor U33052 (N_33052,N_32196,N_32615);
or U33053 (N_33053,N_32356,N_32708);
or U33054 (N_33054,N_32572,N_32429);
nor U33055 (N_33055,N_32885,N_32881);
nand U33056 (N_33056,N_32111,N_32463);
nand U33057 (N_33057,N_32186,N_32428);
or U33058 (N_33058,N_32293,N_32374);
nand U33059 (N_33059,N_32007,N_32797);
and U33060 (N_33060,N_32573,N_32211);
or U33061 (N_33061,N_32146,N_32684);
xor U33062 (N_33062,N_32446,N_32611);
nor U33063 (N_33063,N_32600,N_32230);
and U33064 (N_33064,N_32244,N_32582);
nand U33065 (N_33065,N_32927,N_32160);
and U33066 (N_33066,N_32270,N_32325);
or U33067 (N_33067,N_32347,N_32808);
xnor U33068 (N_33068,N_32264,N_32798);
nand U33069 (N_33069,N_32425,N_32273);
nand U33070 (N_33070,N_32690,N_32761);
xnor U33071 (N_33071,N_32550,N_32935);
and U33072 (N_33072,N_32110,N_32517);
nor U33073 (N_33073,N_32598,N_32502);
xor U33074 (N_33074,N_32564,N_32886);
xor U33075 (N_33075,N_32465,N_32740);
nand U33076 (N_33076,N_32197,N_32077);
nor U33077 (N_33077,N_32540,N_32910);
and U33078 (N_33078,N_32555,N_32148);
nor U33079 (N_33079,N_32379,N_32867);
or U33080 (N_33080,N_32640,N_32292);
nand U33081 (N_33081,N_32038,N_32753);
xnor U33082 (N_33082,N_32501,N_32345);
or U33083 (N_33083,N_32626,N_32285);
and U33084 (N_33084,N_32701,N_32001);
or U33085 (N_33085,N_32260,N_32468);
nor U33086 (N_33086,N_32721,N_32745);
nand U33087 (N_33087,N_32320,N_32723);
nand U33088 (N_33088,N_32002,N_32929);
xnor U33089 (N_33089,N_32349,N_32547);
or U33090 (N_33090,N_32658,N_32985);
nor U33091 (N_33091,N_32302,N_32856);
xnor U33092 (N_33092,N_32381,N_32968);
nor U33093 (N_33093,N_32335,N_32228);
nor U33094 (N_33094,N_32878,N_32533);
or U33095 (N_33095,N_32754,N_32770);
nor U33096 (N_33096,N_32304,N_32401);
nor U33097 (N_33097,N_32383,N_32673);
and U33098 (N_33098,N_32909,N_32609);
or U33099 (N_33099,N_32827,N_32724);
nor U33100 (N_33100,N_32578,N_32716);
xor U33101 (N_33101,N_32122,N_32902);
nand U33102 (N_33102,N_32950,N_32484);
xor U33103 (N_33103,N_32768,N_32882);
xor U33104 (N_33104,N_32762,N_32460);
xnor U33105 (N_33105,N_32799,N_32834);
or U33106 (N_33106,N_32181,N_32114);
or U33107 (N_33107,N_32445,N_32455);
nor U33108 (N_33108,N_32340,N_32430);
nand U33109 (N_33109,N_32362,N_32554);
or U33110 (N_33110,N_32434,N_32973);
nor U33111 (N_33111,N_32393,N_32964);
nor U33112 (N_33112,N_32793,N_32537);
nor U33113 (N_33113,N_32953,N_32888);
xor U33114 (N_33114,N_32897,N_32986);
and U33115 (N_33115,N_32527,N_32977);
and U33116 (N_33116,N_32033,N_32139);
and U33117 (N_33117,N_32892,N_32601);
and U33118 (N_33118,N_32890,N_32163);
or U33119 (N_33119,N_32342,N_32954);
or U33120 (N_33120,N_32100,N_32289);
or U33121 (N_33121,N_32765,N_32509);
or U33122 (N_33122,N_32741,N_32060);
xor U33123 (N_33123,N_32997,N_32807);
nor U33124 (N_33124,N_32205,N_32200);
and U33125 (N_33125,N_32715,N_32101);
and U33126 (N_33126,N_32086,N_32921);
and U33127 (N_33127,N_32840,N_32507);
or U33128 (N_33128,N_32454,N_32042);
xnor U33129 (N_33129,N_32088,N_32951);
or U33130 (N_33130,N_32041,N_32094);
or U33131 (N_33131,N_32668,N_32229);
or U33132 (N_33132,N_32996,N_32595);
nand U33133 (N_33133,N_32616,N_32378);
xor U33134 (N_33134,N_32129,N_32109);
nor U33135 (N_33135,N_32870,N_32405);
xnor U33136 (N_33136,N_32490,N_32838);
xnor U33137 (N_33137,N_32180,N_32479);
and U33138 (N_33138,N_32521,N_32928);
and U33139 (N_33139,N_32055,N_32506);
and U33140 (N_33140,N_32444,N_32271);
xor U33141 (N_33141,N_32836,N_32584);
or U33142 (N_33142,N_32300,N_32344);
nand U33143 (N_33143,N_32655,N_32792);
nor U33144 (N_33144,N_32981,N_32541);
and U33145 (N_33145,N_32043,N_32680);
nand U33146 (N_33146,N_32423,N_32795);
or U33147 (N_33147,N_32967,N_32470);
nor U33148 (N_33148,N_32955,N_32653);
nor U33149 (N_33149,N_32443,N_32004);
and U33150 (N_33150,N_32843,N_32118);
xnor U33151 (N_33151,N_32394,N_32432);
or U33152 (N_33152,N_32686,N_32860);
xnor U33153 (N_33153,N_32750,N_32102);
and U33154 (N_33154,N_32806,N_32931);
or U33155 (N_33155,N_32717,N_32677);
or U33156 (N_33156,N_32766,N_32865);
nor U33157 (N_33157,N_32089,N_32894);
or U33158 (N_33158,N_32235,N_32764);
xor U33159 (N_33159,N_32995,N_32568);
nand U33160 (N_33160,N_32749,N_32920);
and U33161 (N_33161,N_32046,N_32730);
xnor U33162 (N_33162,N_32301,N_32276);
xor U33163 (N_33163,N_32824,N_32915);
and U33164 (N_33164,N_32656,N_32087);
nand U33165 (N_33165,N_32133,N_32453);
nand U33166 (N_33166,N_32138,N_32567);
or U33167 (N_33167,N_32462,N_32769);
nand U33168 (N_33168,N_32489,N_32830);
nand U33169 (N_33169,N_32755,N_32333);
nor U33170 (N_33170,N_32030,N_32669);
or U33171 (N_33171,N_32923,N_32869);
and U33172 (N_33172,N_32505,N_32189);
xnor U33173 (N_33173,N_32687,N_32746);
nand U33174 (N_33174,N_32647,N_32905);
xnor U33175 (N_33175,N_32571,N_32308);
and U33176 (N_33176,N_32137,N_32670);
nor U33177 (N_33177,N_32406,N_32152);
nand U33178 (N_33178,N_32108,N_32529);
nor U33179 (N_33179,N_32321,N_32650);
nor U33180 (N_33180,N_32855,N_32091);
or U33181 (N_33181,N_32848,N_32663);
or U33182 (N_33182,N_32780,N_32872);
xor U33183 (N_33183,N_32831,N_32127);
xor U33184 (N_33184,N_32667,N_32078);
and U33185 (N_33185,N_32115,N_32599);
and U33186 (N_33186,N_32081,N_32058);
xnor U33187 (N_33187,N_32469,N_32941);
nand U33188 (N_33188,N_32240,N_32261);
or U33189 (N_33189,N_32027,N_32771);
or U33190 (N_33190,N_32164,N_32212);
and U33191 (N_33191,N_32279,N_32158);
nand U33192 (N_33192,N_32391,N_32070);
nor U33193 (N_33193,N_32408,N_32998);
nand U33194 (N_33194,N_32410,N_32364);
xor U33195 (N_33195,N_32777,N_32548);
nand U33196 (N_33196,N_32187,N_32104);
nor U33197 (N_33197,N_32415,N_32911);
xnor U33198 (N_33198,N_32336,N_32738);
or U33199 (N_33199,N_32250,N_32402);
and U33200 (N_33200,N_32718,N_32066);
and U33201 (N_33201,N_32907,N_32709);
nand U33202 (N_33202,N_32280,N_32441);
or U33203 (N_33203,N_32119,N_32492);
and U33204 (N_33204,N_32874,N_32457);
nor U33205 (N_33205,N_32090,N_32560);
and U33206 (N_33206,N_32403,N_32412);
nor U33207 (N_33207,N_32852,N_32859);
and U33208 (N_33208,N_32901,N_32037);
xor U33209 (N_33209,N_32404,N_32606);
xor U33210 (N_33210,N_32047,N_32012);
and U33211 (N_33211,N_32759,N_32612);
nor U33212 (N_33212,N_32858,N_32284);
xnor U33213 (N_33213,N_32096,N_32789);
xnor U33214 (N_33214,N_32553,N_32543);
xnor U33215 (N_33215,N_32665,N_32179);
and U33216 (N_33216,N_32908,N_32832);
xor U33217 (N_33217,N_32711,N_32959);
nand U33218 (N_33218,N_32452,N_32477);
xor U33219 (N_33219,N_32227,N_32355);
xor U33220 (N_33220,N_32372,N_32945);
and U33221 (N_33221,N_32449,N_32318);
and U33222 (N_33222,N_32536,N_32635);
or U33223 (N_33223,N_32918,N_32710);
xor U33224 (N_33224,N_32239,N_32947);
xor U33225 (N_33225,N_32847,N_32512);
nand U33226 (N_33226,N_32175,N_32725);
xor U33227 (N_33227,N_32642,N_32224);
nand U33228 (N_33228,N_32313,N_32949);
nor U33229 (N_33229,N_32628,N_32705);
nand U33230 (N_33230,N_32963,N_32190);
nor U33231 (N_33231,N_32447,N_32513);
and U33232 (N_33232,N_32145,N_32503);
nor U33233 (N_33233,N_32782,N_32552);
xor U33234 (N_33234,N_32074,N_32409);
and U33235 (N_33235,N_32201,N_32322);
nor U33236 (N_33236,N_32514,N_32157);
and U33237 (N_33237,N_32382,N_32011);
and U33238 (N_33238,N_32021,N_32338);
and U33239 (N_33239,N_32204,N_32622);
and U33240 (N_33240,N_32625,N_32295);
nand U33241 (N_33241,N_32944,N_32734);
and U33242 (N_33242,N_32704,N_32035);
nor U33243 (N_33243,N_32937,N_32588);
xnor U33244 (N_33244,N_32407,N_32557);
nand U33245 (N_33245,N_32203,N_32645);
nand U33246 (N_33246,N_32562,N_32987);
and U33247 (N_33247,N_32714,N_32952);
xor U33248 (N_33248,N_32420,N_32194);
nand U33249 (N_33249,N_32330,N_32845);
nor U33250 (N_33250,N_32298,N_32499);
or U33251 (N_33251,N_32072,N_32617);
nand U33252 (N_33252,N_32737,N_32360);
nand U33253 (N_33253,N_32026,N_32130);
and U33254 (N_33254,N_32676,N_32638);
nor U33255 (N_33255,N_32003,N_32960);
or U33256 (N_33256,N_32659,N_32713);
or U33257 (N_33257,N_32822,N_32593);
and U33258 (N_33258,N_32589,N_32359);
or U33259 (N_33259,N_32183,N_32467);
or U33260 (N_33260,N_32172,N_32265);
xnor U33261 (N_33261,N_32871,N_32036);
or U33262 (N_33262,N_32861,N_32833);
nor U33263 (N_33263,N_32828,N_32776);
or U33264 (N_33264,N_32165,N_32850);
xor U33265 (N_33265,N_32636,N_32565);
nand U33266 (N_33266,N_32672,N_32474);
or U33267 (N_33267,N_32475,N_32231);
xor U33268 (N_33268,N_32396,N_32358);
nor U33269 (N_33269,N_32296,N_32252);
and U33270 (N_33270,N_32092,N_32618);
or U33271 (N_33271,N_32728,N_32563);
nand U33272 (N_33272,N_32983,N_32574);
or U33273 (N_33273,N_32019,N_32257);
xnor U33274 (N_33274,N_32694,N_32569);
or U33275 (N_33275,N_32259,N_32117);
nand U33276 (N_33276,N_32587,N_32286);
and U33277 (N_33277,N_32914,N_32222);
xor U33278 (N_33278,N_32121,N_32255);
or U33279 (N_33279,N_32519,N_32083);
xnor U33280 (N_33280,N_32310,N_32226);
nand U33281 (N_33281,N_32691,N_32796);
nor U33282 (N_33282,N_32542,N_32373);
or U33283 (N_33283,N_32040,N_32632);
nor U33284 (N_33284,N_32241,N_32916);
and U33285 (N_33285,N_32829,N_32620);
and U33286 (N_33286,N_32208,N_32974);
nand U33287 (N_33287,N_32895,N_32561);
nor U33288 (N_33288,N_32032,N_32900);
nor U33289 (N_33289,N_32323,N_32245);
and U33290 (N_33290,N_32603,N_32893);
nor U33291 (N_33291,N_32161,N_32290);
nor U33292 (N_33292,N_32919,N_32884);
xor U33293 (N_33293,N_32167,N_32262);
nand U33294 (N_33294,N_32438,N_32525);
nand U33295 (N_33295,N_32681,N_32388);
xnor U33296 (N_33296,N_32868,N_32785);
and U33297 (N_33297,N_32608,N_32069);
xor U33298 (N_33298,N_32597,N_32254);
xnor U33299 (N_33299,N_32498,N_32306);
and U33300 (N_33300,N_32846,N_32267);
nand U33301 (N_33301,N_32633,N_32147);
and U33302 (N_33302,N_32610,N_32530);
xor U33303 (N_33303,N_32247,N_32482);
or U33304 (N_33304,N_32339,N_32098);
xnor U33305 (N_33305,N_32712,N_32524);
or U33306 (N_33306,N_32692,N_32791);
or U33307 (N_33307,N_32596,N_32075);
and U33308 (N_33308,N_32674,N_32079);
or U33309 (N_33309,N_32093,N_32120);
or U33310 (N_33310,N_32948,N_32456);
nand U33311 (N_33311,N_32192,N_32450);
xnor U33312 (N_33312,N_32585,N_32825);
xnor U33313 (N_33313,N_32508,N_32478);
and U33314 (N_33314,N_32486,N_32575);
nand U33315 (N_33315,N_32990,N_32049);
nand U33316 (N_33316,N_32051,N_32215);
or U33317 (N_33317,N_32283,N_32274);
and U33318 (N_33318,N_32485,N_32375);
xnor U33319 (N_33319,N_32234,N_32275);
and U33320 (N_33320,N_32526,N_32437);
xor U33321 (N_33321,N_32875,N_32925);
or U33322 (N_33322,N_32071,N_32969);
nand U33323 (N_33323,N_32461,N_32095);
nand U33324 (N_33324,N_32178,N_32837);
and U33325 (N_33325,N_32696,N_32442);
and U33326 (N_33326,N_32581,N_32065);
nor U33327 (N_33327,N_32938,N_32464);
and U33328 (N_33328,N_32170,N_32748);
and U33329 (N_33329,N_32787,N_32297);
nand U33330 (N_33330,N_32757,N_32131);
nand U33331 (N_33331,N_32500,N_32013);
xnor U33332 (N_33332,N_32218,N_32809);
nor U33333 (N_33333,N_32084,N_32387);
nand U33334 (N_33334,N_32862,N_32365);
and U33335 (N_33335,N_32288,N_32466);
nand U33336 (N_33336,N_32031,N_32991);
nor U33337 (N_33337,N_32337,N_32132);
or U33338 (N_33338,N_32068,N_32767);
and U33339 (N_33339,N_32061,N_32932);
and U33340 (N_33340,N_32353,N_32142);
or U33341 (N_33341,N_32343,N_32854);
nand U33342 (N_33342,N_32989,N_32097);
nor U33343 (N_33343,N_32005,N_32417);
nand U33344 (N_33344,N_32660,N_32305);
nor U33345 (N_33345,N_32763,N_32392);
nor U33346 (N_33346,N_32015,N_32341);
xnor U33347 (N_33347,N_32361,N_32328);
and U33348 (N_33348,N_32592,N_32816);
and U33349 (N_33349,N_32707,N_32815);
and U33350 (N_33350,N_32934,N_32842);
xor U33351 (N_33351,N_32487,N_32010);
and U33352 (N_33352,N_32821,N_32367);
nand U33353 (N_33353,N_32050,N_32168);
nand U33354 (N_33354,N_32930,N_32926);
or U33355 (N_33355,N_32414,N_32957);
xnor U33356 (N_33356,N_32794,N_32644);
xnor U33357 (N_33357,N_32511,N_32020);
and U33358 (N_33358,N_32057,N_32583);
and U33359 (N_33359,N_32188,N_32141);
nor U33360 (N_33360,N_32958,N_32136);
nand U33361 (N_33361,N_32440,N_32458);
nor U33362 (N_33362,N_32326,N_32819);
nor U33363 (N_33363,N_32426,N_32184);
and U33364 (N_33364,N_32804,N_32613);
and U33365 (N_33365,N_32193,N_32346);
nand U33366 (N_33366,N_32853,N_32480);
nor U33367 (N_33367,N_32107,N_32350);
xnor U33368 (N_33368,N_32311,N_32332);
or U33369 (N_33369,N_32277,N_32422);
or U33370 (N_33370,N_32913,N_32282);
nand U33371 (N_33371,N_32922,N_32857);
and U33372 (N_33372,N_32980,N_32233);
and U33373 (N_33373,N_32648,N_32803);
xnor U33374 (N_33374,N_32143,N_32024);
nor U33375 (N_33375,N_32898,N_32451);
and U33376 (N_33376,N_32029,N_32942);
nand U33377 (N_33377,N_32329,N_32214);
nor U33378 (N_33378,N_32048,N_32805);
xor U33379 (N_33379,N_32331,N_32817);
and U33380 (N_33380,N_32539,N_32624);
nor U33381 (N_33381,N_32783,N_32219);
or U33382 (N_33382,N_32646,N_32722);
and U33383 (N_33383,N_32278,N_32876);
nor U33384 (N_33384,N_32291,N_32719);
xnor U33385 (N_33385,N_32221,N_32076);
nand U33386 (N_33386,N_32421,N_32756);
and U33387 (N_33387,N_32621,N_32727);
and U33388 (N_33388,N_32844,N_32811);
or U33389 (N_33389,N_32839,N_32518);
xor U33390 (N_33390,N_32022,N_32814);
and U33391 (N_33391,N_32198,N_32067);
nor U33392 (N_33392,N_32906,N_32695);
or U33393 (N_33393,N_32970,N_32390);
or U33394 (N_33394,N_32384,N_32576);
nor U33395 (N_33395,N_32436,N_32851);
and U33396 (N_33396,N_32546,N_32023);
or U33397 (N_33397,N_32496,N_32818);
xor U33398 (N_33398,N_32377,N_32433);
xor U33399 (N_33399,N_32899,N_32863);
nor U33400 (N_33400,N_32739,N_32395);
and U33401 (N_33401,N_32352,N_32220);
nand U33402 (N_33402,N_32113,N_32354);
nand U33403 (N_33403,N_32813,N_32662);
or U33404 (N_33404,N_32849,N_32820);
nand U33405 (N_33405,N_32363,N_32912);
nor U33406 (N_33406,N_32281,N_32312);
nand U33407 (N_33407,N_32720,N_32128);
or U33408 (N_33408,N_32400,N_32751);
and U33409 (N_33409,N_32357,N_32242);
and U33410 (N_33410,N_32351,N_32726);
nand U33411 (N_33411,N_32772,N_32657);
nor U33412 (N_33412,N_32411,N_32471);
and U33413 (N_33413,N_32327,N_32397);
xor U33414 (N_33414,N_32016,N_32594);
xor U33415 (N_33415,N_32431,N_32493);
nor U33416 (N_33416,N_32287,N_32034);
nor U33417 (N_33417,N_32864,N_32877);
or U33418 (N_33418,N_32316,N_32532);
nor U33419 (N_33419,N_32641,N_32000);
and U33420 (N_33420,N_32213,N_32217);
nand U33421 (N_33421,N_32054,N_32549);
or U33422 (N_33422,N_32018,N_32841);
nor U33423 (N_33423,N_32269,N_32577);
xor U33424 (N_33424,N_32558,N_32778);
or U33425 (N_33425,N_32176,N_32125);
xor U33426 (N_33426,N_32123,N_32099);
nand U33427 (N_33427,N_32314,N_32473);
and U33428 (N_33428,N_32134,N_32253);
xnor U33429 (N_33429,N_32209,N_32904);
xor U33430 (N_33430,N_32053,N_32169);
and U33431 (N_33431,N_32887,N_32966);
nand U33432 (N_33432,N_32237,N_32781);
or U33433 (N_33433,N_32649,N_32510);
nor U33434 (N_33434,N_32736,N_32810);
xnor U33435 (N_33435,N_32579,N_32317);
or U33436 (N_33436,N_32732,N_32946);
nand U33437 (N_33437,N_32972,N_32199);
or U33438 (N_33438,N_32826,N_32627);
or U33439 (N_33439,N_32788,N_32643);
nor U33440 (N_33440,N_32689,N_32105);
xor U33441 (N_33441,N_32126,N_32385);
and U33442 (N_33442,N_32315,N_32059);
xor U33443 (N_33443,N_32427,N_32917);
nor U33444 (N_33444,N_32682,N_32742);
xnor U33445 (N_33445,N_32223,N_32376);
and U33446 (N_33446,N_32654,N_32398);
nor U33447 (N_33447,N_32238,N_32683);
and U33448 (N_33448,N_32940,N_32174);
nor U33449 (N_33449,N_32085,N_32251);
nor U33450 (N_33450,N_32965,N_32319);
or U33451 (N_33451,N_32439,N_32294);
xor U33452 (N_33452,N_32448,N_32272);
nand U33453 (N_33453,N_32784,N_32140);
and U33454 (N_33454,N_32155,N_32619);
xnor U33455 (N_33455,N_32590,N_32516);
and U33456 (N_33456,N_32936,N_32823);
and U33457 (N_33457,N_32062,N_32380);
or U33458 (N_33458,N_32151,N_32303);
nor U33459 (N_33459,N_32800,N_32028);
or U33460 (N_33460,N_32206,N_32639);
nor U33461 (N_33461,N_32435,N_32006);
nand U33462 (N_33462,N_32039,N_32210);
or U33463 (N_33463,N_32459,N_32520);
and U33464 (N_33464,N_32773,N_32225);
or U33465 (N_33465,N_32962,N_32488);
nand U33466 (N_33466,N_32116,N_32971);
or U33467 (N_33467,N_32637,N_32153);
or U33468 (N_33468,N_32263,N_32424);
and U33469 (N_33469,N_32063,N_32258);
nor U33470 (N_33470,N_32515,N_32185);
and U33471 (N_33471,N_32939,N_32866);
nand U33472 (N_33472,N_32984,N_32177);
and U33473 (N_33473,N_32993,N_32476);
nor U33474 (N_33474,N_32307,N_32744);
or U33475 (N_33475,N_32528,N_32369);
nand U33476 (N_33476,N_32534,N_32173);
and U33477 (N_33477,N_32045,N_32790);
nor U33478 (N_33478,N_32064,N_32693);
or U33479 (N_33479,N_32014,N_32671);
xor U33480 (N_33480,N_32698,N_32236);
or U33481 (N_33481,N_32933,N_32883);
or U33482 (N_33482,N_32371,N_32992);
or U33483 (N_33483,N_32651,N_32268);
nand U33484 (N_33484,N_32812,N_32368);
xor U33485 (N_33485,N_32835,N_32891);
nand U33486 (N_33486,N_32523,N_32495);
nand U33487 (N_33487,N_32988,N_32370);
or U33488 (N_33488,N_32880,N_32752);
nor U33489 (N_33489,N_32538,N_32246);
or U33490 (N_33490,N_32309,N_32607);
xor U33491 (N_33491,N_32399,N_32685);
xor U33492 (N_33492,N_32166,N_32207);
nor U33493 (N_33493,N_32156,N_32703);
nor U33494 (N_33494,N_32025,N_32758);
and U33495 (N_33495,N_32481,N_32775);
nand U33496 (N_33496,N_32879,N_32666);
xor U33497 (N_33497,N_32112,N_32943);
nor U33498 (N_33498,N_32413,N_32535);
or U33499 (N_33499,N_32903,N_32700);
or U33500 (N_33500,N_32331,N_32146);
nor U33501 (N_33501,N_32861,N_32852);
and U33502 (N_33502,N_32589,N_32850);
or U33503 (N_33503,N_32234,N_32661);
xnor U33504 (N_33504,N_32558,N_32310);
xnor U33505 (N_33505,N_32674,N_32217);
and U33506 (N_33506,N_32420,N_32259);
xnor U33507 (N_33507,N_32988,N_32015);
nor U33508 (N_33508,N_32546,N_32334);
nand U33509 (N_33509,N_32746,N_32884);
nand U33510 (N_33510,N_32493,N_32112);
or U33511 (N_33511,N_32531,N_32305);
or U33512 (N_33512,N_32788,N_32241);
nand U33513 (N_33513,N_32716,N_32043);
or U33514 (N_33514,N_32318,N_32343);
or U33515 (N_33515,N_32967,N_32482);
or U33516 (N_33516,N_32898,N_32746);
or U33517 (N_33517,N_32685,N_32850);
nand U33518 (N_33518,N_32084,N_32891);
or U33519 (N_33519,N_32089,N_32492);
xnor U33520 (N_33520,N_32785,N_32529);
or U33521 (N_33521,N_32326,N_32119);
nor U33522 (N_33522,N_32812,N_32716);
or U33523 (N_33523,N_32879,N_32428);
nand U33524 (N_33524,N_32879,N_32009);
nor U33525 (N_33525,N_32374,N_32907);
nand U33526 (N_33526,N_32244,N_32347);
nand U33527 (N_33527,N_32707,N_32935);
or U33528 (N_33528,N_32071,N_32450);
xnor U33529 (N_33529,N_32552,N_32642);
nor U33530 (N_33530,N_32669,N_32549);
and U33531 (N_33531,N_32460,N_32026);
xnor U33532 (N_33532,N_32769,N_32055);
and U33533 (N_33533,N_32740,N_32105);
nand U33534 (N_33534,N_32705,N_32384);
nor U33535 (N_33535,N_32163,N_32722);
nand U33536 (N_33536,N_32434,N_32023);
xnor U33537 (N_33537,N_32454,N_32975);
nor U33538 (N_33538,N_32983,N_32919);
or U33539 (N_33539,N_32880,N_32330);
or U33540 (N_33540,N_32215,N_32477);
nor U33541 (N_33541,N_32689,N_32209);
or U33542 (N_33542,N_32927,N_32391);
xor U33543 (N_33543,N_32903,N_32600);
nor U33544 (N_33544,N_32634,N_32410);
nand U33545 (N_33545,N_32234,N_32773);
or U33546 (N_33546,N_32158,N_32591);
or U33547 (N_33547,N_32612,N_32072);
xor U33548 (N_33548,N_32255,N_32757);
xor U33549 (N_33549,N_32455,N_32138);
or U33550 (N_33550,N_32967,N_32259);
and U33551 (N_33551,N_32729,N_32813);
nand U33552 (N_33552,N_32141,N_32391);
nor U33553 (N_33553,N_32241,N_32680);
nor U33554 (N_33554,N_32497,N_32838);
or U33555 (N_33555,N_32912,N_32431);
nor U33556 (N_33556,N_32014,N_32730);
xor U33557 (N_33557,N_32563,N_32330);
xnor U33558 (N_33558,N_32689,N_32115);
xor U33559 (N_33559,N_32726,N_32868);
nor U33560 (N_33560,N_32229,N_32653);
nor U33561 (N_33561,N_32215,N_32424);
xor U33562 (N_33562,N_32673,N_32332);
nand U33563 (N_33563,N_32927,N_32114);
nand U33564 (N_33564,N_32828,N_32234);
and U33565 (N_33565,N_32934,N_32557);
or U33566 (N_33566,N_32071,N_32800);
or U33567 (N_33567,N_32686,N_32024);
nor U33568 (N_33568,N_32379,N_32412);
or U33569 (N_33569,N_32785,N_32748);
nor U33570 (N_33570,N_32837,N_32441);
nor U33571 (N_33571,N_32870,N_32949);
and U33572 (N_33572,N_32779,N_32588);
or U33573 (N_33573,N_32607,N_32328);
nor U33574 (N_33574,N_32482,N_32913);
or U33575 (N_33575,N_32236,N_32682);
and U33576 (N_33576,N_32172,N_32045);
xor U33577 (N_33577,N_32984,N_32289);
nor U33578 (N_33578,N_32484,N_32867);
nand U33579 (N_33579,N_32009,N_32088);
and U33580 (N_33580,N_32646,N_32433);
nor U33581 (N_33581,N_32537,N_32643);
xnor U33582 (N_33582,N_32425,N_32649);
nor U33583 (N_33583,N_32528,N_32377);
and U33584 (N_33584,N_32376,N_32316);
and U33585 (N_33585,N_32019,N_32203);
nand U33586 (N_33586,N_32602,N_32789);
or U33587 (N_33587,N_32108,N_32513);
and U33588 (N_33588,N_32159,N_32920);
nand U33589 (N_33589,N_32039,N_32696);
nor U33590 (N_33590,N_32222,N_32934);
nor U33591 (N_33591,N_32434,N_32853);
xor U33592 (N_33592,N_32877,N_32155);
nor U33593 (N_33593,N_32606,N_32765);
nor U33594 (N_33594,N_32626,N_32070);
or U33595 (N_33595,N_32485,N_32830);
and U33596 (N_33596,N_32562,N_32839);
nand U33597 (N_33597,N_32288,N_32094);
or U33598 (N_33598,N_32077,N_32617);
xnor U33599 (N_33599,N_32655,N_32030);
and U33600 (N_33600,N_32618,N_32270);
nor U33601 (N_33601,N_32524,N_32421);
and U33602 (N_33602,N_32079,N_32475);
nor U33603 (N_33603,N_32052,N_32599);
and U33604 (N_33604,N_32829,N_32483);
nor U33605 (N_33605,N_32117,N_32838);
and U33606 (N_33606,N_32108,N_32637);
and U33607 (N_33607,N_32951,N_32819);
and U33608 (N_33608,N_32240,N_32402);
or U33609 (N_33609,N_32492,N_32145);
xor U33610 (N_33610,N_32628,N_32908);
nor U33611 (N_33611,N_32456,N_32305);
xor U33612 (N_33612,N_32835,N_32630);
nor U33613 (N_33613,N_32280,N_32821);
or U33614 (N_33614,N_32778,N_32834);
nand U33615 (N_33615,N_32406,N_32313);
xor U33616 (N_33616,N_32705,N_32629);
nor U33617 (N_33617,N_32059,N_32844);
nand U33618 (N_33618,N_32280,N_32945);
xor U33619 (N_33619,N_32372,N_32623);
nor U33620 (N_33620,N_32215,N_32574);
or U33621 (N_33621,N_32004,N_32088);
or U33622 (N_33622,N_32069,N_32060);
xnor U33623 (N_33623,N_32343,N_32655);
nand U33624 (N_33624,N_32838,N_32735);
or U33625 (N_33625,N_32499,N_32428);
and U33626 (N_33626,N_32355,N_32977);
nor U33627 (N_33627,N_32998,N_32267);
nand U33628 (N_33628,N_32386,N_32638);
xor U33629 (N_33629,N_32051,N_32992);
or U33630 (N_33630,N_32095,N_32318);
xor U33631 (N_33631,N_32117,N_32817);
and U33632 (N_33632,N_32703,N_32205);
or U33633 (N_33633,N_32112,N_32598);
or U33634 (N_33634,N_32143,N_32028);
and U33635 (N_33635,N_32984,N_32861);
nor U33636 (N_33636,N_32302,N_32740);
xor U33637 (N_33637,N_32974,N_32287);
and U33638 (N_33638,N_32092,N_32827);
and U33639 (N_33639,N_32238,N_32941);
and U33640 (N_33640,N_32743,N_32755);
xor U33641 (N_33641,N_32541,N_32509);
nand U33642 (N_33642,N_32238,N_32567);
and U33643 (N_33643,N_32403,N_32703);
or U33644 (N_33644,N_32367,N_32264);
or U33645 (N_33645,N_32519,N_32106);
or U33646 (N_33646,N_32425,N_32044);
xnor U33647 (N_33647,N_32191,N_32373);
nor U33648 (N_33648,N_32853,N_32633);
and U33649 (N_33649,N_32131,N_32515);
nand U33650 (N_33650,N_32528,N_32447);
nand U33651 (N_33651,N_32812,N_32673);
and U33652 (N_33652,N_32224,N_32958);
or U33653 (N_33653,N_32271,N_32466);
xnor U33654 (N_33654,N_32701,N_32885);
and U33655 (N_33655,N_32449,N_32176);
and U33656 (N_33656,N_32000,N_32218);
nor U33657 (N_33657,N_32499,N_32768);
nor U33658 (N_33658,N_32661,N_32798);
and U33659 (N_33659,N_32060,N_32661);
xnor U33660 (N_33660,N_32274,N_32795);
xor U33661 (N_33661,N_32786,N_32056);
and U33662 (N_33662,N_32696,N_32676);
or U33663 (N_33663,N_32432,N_32533);
and U33664 (N_33664,N_32762,N_32599);
or U33665 (N_33665,N_32242,N_32743);
xor U33666 (N_33666,N_32669,N_32665);
and U33667 (N_33667,N_32963,N_32625);
xor U33668 (N_33668,N_32657,N_32920);
and U33669 (N_33669,N_32277,N_32506);
nor U33670 (N_33670,N_32795,N_32669);
nand U33671 (N_33671,N_32037,N_32424);
or U33672 (N_33672,N_32763,N_32691);
or U33673 (N_33673,N_32026,N_32175);
and U33674 (N_33674,N_32478,N_32311);
nor U33675 (N_33675,N_32013,N_32113);
xnor U33676 (N_33676,N_32937,N_32627);
nor U33677 (N_33677,N_32964,N_32330);
xnor U33678 (N_33678,N_32242,N_32217);
nand U33679 (N_33679,N_32369,N_32691);
xnor U33680 (N_33680,N_32132,N_32752);
and U33681 (N_33681,N_32013,N_32456);
nor U33682 (N_33682,N_32526,N_32584);
xor U33683 (N_33683,N_32805,N_32903);
or U33684 (N_33684,N_32099,N_32889);
or U33685 (N_33685,N_32313,N_32089);
nand U33686 (N_33686,N_32724,N_32118);
or U33687 (N_33687,N_32657,N_32613);
xor U33688 (N_33688,N_32803,N_32488);
and U33689 (N_33689,N_32376,N_32210);
nor U33690 (N_33690,N_32179,N_32952);
or U33691 (N_33691,N_32933,N_32759);
xor U33692 (N_33692,N_32320,N_32138);
and U33693 (N_33693,N_32294,N_32889);
and U33694 (N_33694,N_32262,N_32194);
or U33695 (N_33695,N_32429,N_32871);
nor U33696 (N_33696,N_32068,N_32210);
and U33697 (N_33697,N_32068,N_32239);
nor U33698 (N_33698,N_32116,N_32541);
nand U33699 (N_33699,N_32824,N_32992);
nor U33700 (N_33700,N_32130,N_32428);
or U33701 (N_33701,N_32793,N_32425);
xnor U33702 (N_33702,N_32747,N_32367);
and U33703 (N_33703,N_32750,N_32708);
xnor U33704 (N_33704,N_32980,N_32686);
nor U33705 (N_33705,N_32931,N_32065);
and U33706 (N_33706,N_32872,N_32650);
xor U33707 (N_33707,N_32888,N_32312);
and U33708 (N_33708,N_32764,N_32934);
and U33709 (N_33709,N_32585,N_32558);
nand U33710 (N_33710,N_32013,N_32080);
xor U33711 (N_33711,N_32249,N_32691);
nor U33712 (N_33712,N_32317,N_32974);
nor U33713 (N_33713,N_32611,N_32214);
or U33714 (N_33714,N_32660,N_32517);
nand U33715 (N_33715,N_32798,N_32458);
or U33716 (N_33716,N_32596,N_32128);
xor U33717 (N_33717,N_32576,N_32470);
nand U33718 (N_33718,N_32811,N_32493);
xor U33719 (N_33719,N_32731,N_32085);
and U33720 (N_33720,N_32823,N_32607);
nor U33721 (N_33721,N_32856,N_32976);
or U33722 (N_33722,N_32860,N_32790);
or U33723 (N_33723,N_32122,N_32362);
and U33724 (N_33724,N_32398,N_32401);
or U33725 (N_33725,N_32888,N_32401);
and U33726 (N_33726,N_32262,N_32128);
nand U33727 (N_33727,N_32412,N_32978);
nand U33728 (N_33728,N_32233,N_32176);
nand U33729 (N_33729,N_32207,N_32366);
and U33730 (N_33730,N_32270,N_32396);
and U33731 (N_33731,N_32764,N_32393);
or U33732 (N_33732,N_32490,N_32979);
xnor U33733 (N_33733,N_32421,N_32122);
nor U33734 (N_33734,N_32500,N_32384);
or U33735 (N_33735,N_32980,N_32373);
and U33736 (N_33736,N_32112,N_32121);
or U33737 (N_33737,N_32885,N_32554);
xnor U33738 (N_33738,N_32525,N_32770);
or U33739 (N_33739,N_32213,N_32898);
nor U33740 (N_33740,N_32036,N_32644);
nand U33741 (N_33741,N_32392,N_32554);
and U33742 (N_33742,N_32917,N_32097);
or U33743 (N_33743,N_32428,N_32589);
xor U33744 (N_33744,N_32440,N_32848);
or U33745 (N_33745,N_32526,N_32264);
nor U33746 (N_33746,N_32879,N_32188);
xnor U33747 (N_33747,N_32437,N_32047);
nor U33748 (N_33748,N_32063,N_32394);
xnor U33749 (N_33749,N_32539,N_32227);
xor U33750 (N_33750,N_32020,N_32399);
nand U33751 (N_33751,N_32259,N_32932);
nor U33752 (N_33752,N_32537,N_32041);
and U33753 (N_33753,N_32700,N_32662);
or U33754 (N_33754,N_32455,N_32261);
xor U33755 (N_33755,N_32871,N_32832);
nand U33756 (N_33756,N_32441,N_32543);
nor U33757 (N_33757,N_32004,N_32128);
or U33758 (N_33758,N_32516,N_32354);
nand U33759 (N_33759,N_32603,N_32264);
nor U33760 (N_33760,N_32403,N_32058);
and U33761 (N_33761,N_32219,N_32057);
xor U33762 (N_33762,N_32824,N_32440);
and U33763 (N_33763,N_32953,N_32778);
and U33764 (N_33764,N_32221,N_32453);
nor U33765 (N_33765,N_32759,N_32593);
nor U33766 (N_33766,N_32830,N_32261);
or U33767 (N_33767,N_32704,N_32653);
nor U33768 (N_33768,N_32584,N_32115);
and U33769 (N_33769,N_32978,N_32086);
xnor U33770 (N_33770,N_32998,N_32712);
or U33771 (N_33771,N_32266,N_32743);
nor U33772 (N_33772,N_32172,N_32202);
nor U33773 (N_33773,N_32385,N_32798);
nor U33774 (N_33774,N_32761,N_32514);
xor U33775 (N_33775,N_32354,N_32845);
nor U33776 (N_33776,N_32891,N_32620);
nor U33777 (N_33777,N_32686,N_32815);
and U33778 (N_33778,N_32497,N_32655);
xnor U33779 (N_33779,N_32754,N_32449);
and U33780 (N_33780,N_32767,N_32074);
nor U33781 (N_33781,N_32271,N_32118);
nand U33782 (N_33782,N_32065,N_32493);
or U33783 (N_33783,N_32271,N_32747);
nand U33784 (N_33784,N_32453,N_32136);
nor U33785 (N_33785,N_32517,N_32474);
nor U33786 (N_33786,N_32080,N_32786);
or U33787 (N_33787,N_32782,N_32829);
nor U33788 (N_33788,N_32606,N_32852);
and U33789 (N_33789,N_32336,N_32921);
or U33790 (N_33790,N_32072,N_32959);
nand U33791 (N_33791,N_32208,N_32618);
xor U33792 (N_33792,N_32258,N_32207);
and U33793 (N_33793,N_32932,N_32398);
and U33794 (N_33794,N_32689,N_32496);
nor U33795 (N_33795,N_32591,N_32187);
or U33796 (N_33796,N_32913,N_32357);
and U33797 (N_33797,N_32700,N_32484);
nand U33798 (N_33798,N_32121,N_32895);
xor U33799 (N_33799,N_32046,N_32218);
nor U33800 (N_33800,N_32308,N_32370);
nor U33801 (N_33801,N_32438,N_32100);
and U33802 (N_33802,N_32942,N_32603);
or U33803 (N_33803,N_32683,N_32699);
and U33804 (N_33804,N_32185,N_32076);
nand U33805 (N_33805,N_32242,N_32108);
or U33806 (N_33806,N_32179,N_32320);
and U33807 (N_33807,N_32949,N_32481);
or U33808 (N_33808,N_32511,N_32711);
and U33809 (N_33809,N_32671,N_32786);
and U33810 (N_33810,N_32165,N_32918);
nand U33811 (N_33811,N_32494,N_32371);
and U33812 (N_33812,N_32973,N_32881);
xnor U33813 (N_33813,N_32444,N_32049);
xor U33814 (N_33814,N_32756,N_32514);
or U33815 (N_33815,N_32305,N_32432);
nand U33816 (N_33816,N_32097,N_32767);
xor U33817 (N_33817,N_32720,N_32532);
nor U33818 (N_33818,N_32406,N_32440);
nor U33819 (N_33819,N_32726,N_32700);
or U33820 (N_33820,N_32882,N_32197);
nor U33821 (N_33821,N_32330,N_32194);
xnor U33822 (N_33822,N_32921,N_32171);
or U33823 (N_33823,N_32296,N_32676);
or U33824 (N_33824,N_32959,N_32750);
nand U33825 (N_33825,N_32846,N_32800);
nand U33826 (N_33826,N_32006,N_32921);
or U33827 (N_33827,N_32910,N_32811);
or U33828 (N_33828,N_32722,N_32511);
xnor U33829 (N_33829,N_32507,N_32526);
nand U33830 (N_33830,N_32298,N_32990);
nor U33831 (N_33831,N_32989,N_32954);
and U33832 (N_33832,N_32409,N_32838);
and U33833 (N_33833,N_32000,N_32393);
nand U33834 (N_33834,N_32008,N_32715);
nand U33835 (N_33835,N_32270,N_32977);
xor U33836 (N_33836,N_32119,N_32743);
and U33837 (N_33837,N_32418,N_32186);
xnor U33838 (N_33838,N_32167,N_32825);
nand U33839 (N_33839,N_32036,N_32541);
nor U33840 (N_33840,N_32428,N_32724);
and U33841 (N_33841,N_32152,N_32461);
and U33842 (N_33842,N_32427,N_32464);
or U33843 (N_33843,N_32841,N_32223);
and U33844 (N_33844,N_32105,N_32887);
or U33845 (N_33845,N_32924,N_32392);
nor U33846 (N_33846,N_32415,N_32397);
nor U33847 (N_33847,N_32223,N_32953);
or U33848 (N_33848,N_32141,N_32014);
and U33849 (N_33849,N_32990,N_32236);
or U33850 (N_33850,N_32354,N_32724);
xor U33851 (N_33851,N_32802,N_32391);
nor U33852 (N_33852,N_32878,N_32860);
nor U33853 (N_33853,N_32890,N_32087);
and U33854 (N_33854,N_32078,N_32278);
nor U33855 (N_33855,N_32875,N_32465);
and U33856 (N_33856,N_32133,N_32509);
nor U33857 (N_33857,N_32636,N_32825);
xor U33858 (N_33858,N_32982,N_32965);
and U33859 (N_33859,N_32271,N_32218);
or U33860 (N_33860,N_32702,N_32612);
nand U33861 (N_33861,N_32696,N_32581);
nand U33862 (N_33862,N_32380,N_32093);
or U33863 (N_33863,N_32833,N_32666);
or U33864 (N_33864,N_32961,N_32437);
xor U33865 (N_33865,N_32336,N_32469);
nand U33866 (N_33866,N_32208,N_32251);
and U33867 (N_33867,N_32739,N_32359);
and U33868 (N_33868,N_32026,N_32853);
nand U33869 (N_33869,N_32488,N_32969);
and U33870 (N_33870,N_32176,N_32473);
nor U33871 (N_33871,N_32642,N_32870);
xor U33872 (N_33872,N_32001,N_32576);
nand U33873 (N_33873,N_32252,N_32279);
and U33874 (N_33874,N_32927,N_32787);
and U33875 (N_33875,N_32591,N_32814);
xnor U33876 (N_33876,N_32163,N_32812);
or U33877 (N_33877,N_32396,N_32551);
or U33878 (N_33878,N_32624,N_32553);
or U33879 (N_33879,N_32824,N_32449);
and U33880 (N_33880,N_32516,N_32799);
nand U33881 (N_33881,N_32135,N_32395);
or U33882 (N_33882,N_32017,N_32648);
nor U33883 (N_33883,N_32957,N_32263);
and U33884 (N_33884,N_32253,N_32586);
nor U33885 (N_33885,N_32648,N_32117);
and U33886 (N_33886,N_32307,N_32900);
and U33887 (N_33887,N_32477,N_32686);
nand U33888 (N_33888,N_32965,N_32936);
nand U33889 (N_33889,N_32710,N_32028);
nor U33890 (N_33890,N_32015,N_32171);
or U33891 (N_33891,N_32790,N_32188);
and U33892 (N_33892,N_32414,N_32468);
and U33893 (N_33893,N_32440,N_32018);
and U33894 (N_33894,N_32677,N_32749);
or U33895 (N_33895,N_32149,N_32516);
or U33896 (N_33896,N_32369,N_32563);
xor U33897 (N_33897,N_32316,N_32343);
nor U33898 (N_33898,N_32037,N_32659);
nor U33899 (N_33899,N_32995,N_32010);
xnor U33900 (N_33900,N_32612,N_32784);
or U33901 (N_33901,N_32164,N_32999);
xor U33902 (N_33902,N_32542,N_32374);
nand U33903 (N_33903,N_32745,N_32221);
nor U33904 (N_33904,N_32679,N_32172);
xor U33905 (N_33905,N_32316,N_32111);
xor U33906 (N_33906,N_32734,N_32311);
xor U33907 (N_33907,N_32866,N_32243);
or U33908 (N_33908,N_32057,N_32241);
or U33909 (N_33909,N_32481,N_32388);
xor U33910 (N_33910,N_32948,N_32812);
nand U33911 (N_33911,N_32625,N_32802);
nor U33912 (N_33912,N_32817,N_32886);
and U33913 (N_33913,N_32485,N_32932);
and U33914 (N_33914,N_32408,N_32560);
and U33915 (N_33915,N_32779,N_32680);
xor U33916 (N_33916,N_32692,N_32385);
or U33917 (N_33917,N_32701,N_32164);
xnor U33918 (N_33918,N_32197,N_32713);
or U33919 (N_33919,N_32477,N_32559);
xor U33920 (N_33920,N_32940,N_32733);
and U33921 (N_33921,N_32015,N_32011);
nor U33922 (N_33922,N_32695,N_32646);
xnor U33923 (N_33923,N_32775,N_32899);
xor U33924 (N_33924,N_32880,N_32495);
nor U33925 (N_33925,N_32076,N_32569);
xor U33926 (N_33926,N_32327,N_32086);
or U33927 (N_33927,N_32758,N_32126);
nor U33928 (N_33928,N_32270,N_32464);
nand U33929 (N_33929,N_32824,N_32601);
and U33930 (N_33930,N_32071,N_32470);
xnor U33931 (N_33931,N_32247,N_32634);
or U33932 (N_33932,N_32702,N_32735);
nor U33933 (N_33933,N_32209,N_32380);
nor U33934 (N_33934,N_32248,N_32014);
and U33935 (N_33935,N_32078,N_32619);
xnor U33936 (N_33936,N_32059,N_32236);
nor U33937 (N_33937,N_32880,N_32356);
and U33938 (N_33938,N_32413,N_32487);
and U33939 (N_33939,N_32224,N_32344);
or U33940 (N_33940,N_32473,N_32123);
or U33941 (N_33941,N_32692,N_32536);
nand U33942 (N_33942,N_32125,N_32159);
or U33943 (N_33943,N_32627,N_32322);
or U33944 (N_33944,N_32852,N_32735);
or U33945 (N_33945,N_32406,N_32443);
xnor U33946 (N_33946,N_32104,N_32746);
xnor U33947 (N_33947,N_32350,N_32252);
xor U33948 (N_33948,N_32707,N_32756);
xor U33949 (N_33949,N_32801,N_32060);
or U33950 (N_33950,N_32493,N_32421);
xnor U33951 (N_33951,N_32515,N_32844);
xor U33952 (N_33952,N_32127,N_32978);
nor U33953 (N_33953,N_32586,N_32545);
nor U33954 (N_33954,N_32288,N_32765);
nor U33955 (N_33955,N_32072,N_32004);
xor U33956 (N_33956,N_32920,N_32725);
nor U33957 (N_33957,N_32157,N_32094);
or U33958 (N_33958,N_32307,N_32850);
nor U33959 (N_33959,N_32482,N_32191);
nor U33960 (N_33960,N_32883,N_32113);
and U33961 (N_33961,N_32952,N_32332);
or U33962 (N_33962,N_32892,N_32866);
nand U33963 (N_33963,N_32421,N_32758);
and U33964 (N_33964,N_32921,N_32262);
xor U33965 (N_33965,N_32984,N_32704);
or U33966 (N_33966,N_32632,N_32024);
xnor U33967 (N_33967,N_32059,N_32653);
or U33968 (N_33968,N_32433,N_32266);
nand U33969 (N_33969,N_32716,N_32908);
and U33970 (N_33970,N_32275,N_32313);
and U33971 (N_33971,N_32545,N_32879);
nor U33972 (N_33972,N_32155,N_32273);
xor U33973 (N_33973,N_32103,N_32532);
nand U33974 (N_33974,N_32912,N_32931);
nand U33975 (N_33975,N_32203,N_32524);
nor U33976 (N_33976,N_32831,N_32355);
nor U33977 (N_33977,N_32146,N_32703);
nand U33978 (N_33978,N_32747,N_32328);
or U33979 (N_33979,N_32482,N_32592);
nand U33980 (N_33980,N_32886,N_32556);
and U33981 (N_33981,N_32764,N_32508);
and U33982 (N_33982,N_32183,N_32504);
or U33983 (N_33983,N_32184,N_32789);
and U33984 (N_33984,N_32340,N_32427);
or U33985 (N_33985,N_32904,N_32074);
or U33986 (N_33986,N_32199,N_32216);
nor U33987 (N_33987,N_32285,N_32288);
nand U33988 (N_33988,N_32227,N_32710);
and U33989 (N_33989,N_32915,N_32274);
xor U33990 (N_33990,N_32444,N_32439);
xor U33991 (N_33991,N_32086,N_32443);
nor U33992 (N_33992,N_32010,N_32707);
xor U33993 (N_33993,N_32305,N_32597);
nor U33994 (N_33994,N_32683,N_32106);
xor U33995 (N_33995,N_32861,N_32313);
nand U33996 (N_33996,N_32267,N_32792);
or U33997 (N_33997,N_32983,N_32070);
xor U33998 (N_33998,N_32989,N_32017);
xnor U33999 (N_33999,N_32697,N_32929);
xnor U34000 (N_34000,N_33366,N_33657);
or U34001 (N_34001,N_33481,N_33304);
nand U34002 (N_34002,N_33084,N_33718);
nand U34003 (N_34003,N_33556,N_33261);
nand U34004 (N_34004,N_33981,N_33736);
xor U34005 (N_34005,N_33761,N_33226);
or U34006 (N_34006,N_33547,N_33373);
or U34007 (N_34007,N_33571,N_33318);
or U34008 (N_34008,N_33309,N_33335);
or U34009 (N_34009,N_33884,N_33573);
or U34010 (N_34010,N_33900,N_33579);
or U34011 (N_34011,N_33704,N_33178);
nand U34012 (N_34012,N_33349,N_33281);
nand U34013 (N_34013,N_33805,N_33440);
xor U34014 (N_34014,N_33662,N_33024);
nor U34015 (N_34015,N_33765,N_33705);
xnor U34016 (N_34016,N_33406,N_33750);
nand U34017 (N_34017,N_33343,N_33688);
nor U34018 (N_34018,N_33937,N_33523);
nor U34019 (N_34019,N_33040,N_33910);
nor U34020 (N_34020,N_33693,N_33253);
xnor U34021 (N_34021,N_33001,N_33301);
nor U34022 (N_34022,N_33798,N_33310);
xor U34023 (N_34023,N_33103,N_33127);
or U34024 (N_34024,N_33889,N_33743);
xor U34025 (N_34025,N_33933,N_33460);
xor U34026 (N_34026,N_33307,N_33434);
nor U34027 (N_34027,N_33374,N_33558);
and U34028 (N_34028,N_33104,N_33585);
nor U34029 (N_34029,N_33652,N_33152);
xor U34030 (N_34030,N_33522,N_33569);
or U34031 (N_34031,N_33753,N_33022);
nand U34032 (N_34032,N_33436,N_33991);
and U34033 (N_34033,N_33729,N_33714);
nor U34034 (N_34034,N_33251,N_33636);
and U34035 (N_34035,N_33552,N_33696);
xnor U34036 (N_34036,N_33888,N_33962);
nand U34037 (N_34037,N_33972,N_33027);
and U34038 (N_34038,N_33527,N_33215);
nand U34039 (N_34039,N_33727,N_33297);
xnor U34040 (N_34040,N_33970,N_33295);
xor U34041 (N_34041,N_33268,N_33429);
nand U34042 (N_34042,N_33323,N_33923);
and U34043 (N_34043,N_33288,N_33813);
nand U34044 (N_34044,N_33210,N_33612);
and U34045 (N_34045,N_33786,N_33830);
nand U34046 (N_34046,N_33633,N_33413);
nor U34047 (N_34047,N_33713,N_33875);
xnor U34048 (N_34048,N_33627,N_33728);
and U34049 (N_34049,N_33099,N_33218);
or U34050 (N_34050,N_33255,N_33016);
nand U34051 (N_34051,N_33490,N_33073);
and U34052 (N_34052,N_33299,N_33030);
or U34053 (N_34053,N_33576,N_33128);
nand U34054 (N_34054,N_33326,N_33650);
xnor U34055 (N_34055,N_33467,N_33694);
xor U34056 (N_34056,N_33709,N_33492);
nand U34057 (N_34057,N_33480,N_33118);
and U34058 (N_34058,N_33388,N_33620);
xor U34059 (N_34059,N_33855,N_33140);
nor U34060 (N_34060,N_33354,N_33234);
xnor U34061 (N_34061,N_33363,N_33950);
nand U34062 (N_34062,N_33605,N_33998);
xor U34063 (N_34063,N_33738,N_33046);
nor U34064 (N_34064,N_33320,N_33946);
or U34065 (N_34065,N_33050,N_33428);
nor U34066 (N_34066,N_33154,N_33274);
and U34067 (N_34067,N_33822,N_33465);
nand U34068 (N_34068,N_33616,N_33280);
nor U34069 (N_34069,N_33110,N_33723);
xor U34070 (N_34070,N_33665,N_33034);
or U34071 (N_34071,N_33570,N_33105);
xor U34072 (N_34072,N_33638,N_33092);
xnor U34073 (N_34073,N_33070,N_33425);
and U34074 (N_34074,N_33208,N_33940);
xor U34075 (N_34075,N_33449,N_33083);
and U34076 (N_34076,N_33080,N_33992);
xor U34077 (N_34077,N_33157,N_33634);
nor U34078 (N_34078,N_33063,N_33195);
nor U34079 (N_34079,N_33491,N_33142);
and U34080 (N_34080,N_33895,N_33787);
nand U34081 (N_34081,N_33922,N_33849);
and U34082 (N_34082,N_33200,N_33698);
xnor U34083 (N_34083,N_33516,N_33934);
xnor U34084 (N_34084,N_33305,N_33661);
nand U34085 (N_34085,N_33597,N_33517);
or U34086 (N_34086,N_33609,N_33451);
and U34087 (N_34087,N_33463,N_33566);
xnor U34088 (N_34088,N_33416,N_33872);
nand U34089 (N_34089,N_33230,N_33237);
or U34090 (N_34090,N_33509,N_33414);
nor U34091 (N_34091,N_33062,N_33398);
xnor U34092 (N_34092,N_33859,N_33035);
xor U34093 (N_34093,N_33931,N_33377);
or U34094 (N_34094,N_33702,N_33624);
or U34095 (N_34095,N_33640,N_33801);
nor U34096 (N_34096,N_33550,N_33865);
nor U34097 (N_34097,N_33381,N_33932);
nor U34098 (N_34098,N_33722,N_33328);
nand U34099 (N_34099,N_33468,N_33275);
nand U34100 (N_34100,N_33773,N_33028);
and U34101 (N_34101,N_33114,N_33680);
nand U34102 (N_34102,N_33447,N_33706);
or U34103 (N_34103,N_33220,N_33583);
nand U34104 (N_34104,N_33470,N_33474);
nand U34105 (N_34105,N_33511,N_33975);
and U34106 (N_34106,N_33188,N_33559);
and U34107 (N_34107,N_33689,N_33059);
or U34108 (N_34108,N_33581,N_33068);
nand U34109 (N_34109,N_33951,N_33967);
and U34110 (N_34110,N_33444,N_33047);
nand U34111 (N_34111,N_33256,N_33497);
xor U34112 (N_34112,N_33258,N_33685);
or U34113 (N_34113,N_33867,N_33052);
xnor U34114 (N_34114,N_33580,N_33339);
and U34115 (N_34115,N_33303,N_33541);
nor U34116 (N_34116,N_33401,N_33015);
nor U34117 (N_34117,N_33355,N_33686);
xnor U34118 (N_34118,N_33471,N_33213);
nand U34119 (N_34119,N_33143,N_33648);
xor U34120 (N_34120,N_33877,N_33148);
or U34121 (N_34121,N_33603,N_33365);
and U34122 (N_34122,N_33521,N_33458);
and U34123 (N_34123,N_33639,N_33163);
or U34124 (N_34124,N_33312,N_33908);
nand U34125 (N_34125,N_33893,N_33966);
nor U34126 (N_34126,N_33599,N_33101);
and U34127 (N_34127,N_33668,N_33249);
and U34128 (N_34128,N_33300,N_33431);
xor U34129 (N_34129,N_33645,N_33672);
and U34130 (N_34130,N_33655,N_33594);
nor U34131 (N_34131,N_33803,N_33006);
xnor U34132 (N_34132,N_33044,N_33811);
or U34133 (N_34133,N_33766,N_33131);
and U34134 (N_34134,N_33663,N_33942);
and U34135 (N_34135,N_33741,N_33973);
nor U34136 (N_34136,N_33746,N_33219);
and U34137 (N_34137,N_33825,N_33164);
or U34138 (N_34138,N_33284,N_33224);
nand U34139 (N_34139,N_33710,N_33671);
nand U34140 (N_34140,N_33776,N_33771);
nand U34141 (N_34141,N_33731,N_33774);
nor U34142 (N_34142,N_33149,N_33642);
or U34143 (N_34143,N_33898,N_33415);
nand U34144 (N_34144,N_33278,N_33329);
or U34145 (N_34145,N_33854,N_33069);
nor U34146 (N_34146,N_33504,N_33202);
and U34147 (N_34147,N_33435,N_33364);
or U34148 (N_34148,N_33924,N_33989);
xor U34149 (N_34149,N_33876,N_33051);
or U34150 (N_34150,N_33711,N_33109);
or U34151 (N_34151,N_33315,N_33631);
xnor U34152 (N_34152,N_33170,N_33394);
and U34153 (N_34153,N_33720,N_33197);
or U34154 (N_34154,N_33590,N_33337);
or U34155 (N_34155,N_33955,N_33448);
xor U34156 (N_34156,N_33041,N_33145);
xor U34157 (N_34157,N_33112,N_33411);
nand U34158 (N_34158,N_33681,N_33209);
and U34159 (N_34159,N_33977,N_33461);
and U34160 (N_34160,N_33078,N_33317);
or U34161 (N_34161,N_33782,N_33551);
xnor U34162 (N_34162,N_33454,N_33985);
xor U34163 (N_34163,N_33254,N_33917);
nor U34164 (N_34164,N_33997,N_33919);
nor U34165 (N_34165,N_33762,N_33916);
or U34166 (N_34166,N_33726,N_33863);
or U34167 (N_34167,N_33536,N_33690);
xnor U34168 (N_34168,N_33198,N_33183);
nor U34169 (N_34169,N_33539,N_33821);
and U34170 (N_34170,N_33628,N_33061);
nor U34171 (N_34171,N_33294,N_33348);
and U34172 (N_34172,N_33098,N_33752);
or U34173 (N_34173,N_33405,N_33379);
or U34174 (N_34174,N_33371,N_33217);
nand U34175 (N_34175,N_33546,N_33453);
or U34176 (N_34176,N_33948,N_33356);
and U34177 (N_34177,N_33506,N_33032);
nand U34178 (N_34178,N_33840,N_33831);
or U34179 (N_34179,N_33250,N_33850);
and U34180 (N_34180,N_33980,N_33269);
xnor U34181 (N_34181,N_33277,N_33591);
nand U34182 (N_34182,N_33974,N_33141);
and U34183 (N_34183,N_33735,N_33065);
and U34184 (N_34184,N_33238,N_33928);
and U34185 (N_34185,N_33882,N_33235);
nor U34186 (N_34186,N_33904,N_33144);
or U34187 (N_34187,N_33802,N_33654);
or U34188 (N_34188,N_33563,N_33602);
nand U34189 (N_34189,N_33264,N_33136);
nor U34190 (N_34190,N_33800,N_33700);
nor U34191 (N_34191,N_33717,N_33232);
xor U34192 (N_34192,N_33344,N_33990);
nor U34193 (N_34193,N_33091,N_33995);
xnor U34194 (N_34194,N_33669,N_33938);
xor U34195 (N_34195,N_33246,N_33156);
and U34196 (N_34196,N_33483,N_33804);
and U34197 (N_34197,N_33074,N_33513);
and U34198 (N_34198,N_33093,N_33554);
and U34199 (N_34199,N_33031,N_33896);
xor U34200 (N_34200,N_33675,N_33259);
nand U34201 (N_34201,N_33017,N_33173);
nor U34202 (N_34202,N_33560,N_33376);
nor U34203 (N_34203,N_33572,N_33820);
or U34204 (N_34204,N_33999,N_33336);
and U34205 (N_34205,N_33187,N_33116);
nor U34206 (N_34206,N_33806,N_33687);
nor U34207 (N_34207,N_33996,N_33502);
or U34208 (N_34208,N_33360,N_33222);
nand U34209 (N_34209,N_33902,N_33792);
nand U34210 (N_34210,N_33351,N_33026);
nor U34211 (N_34211,N_33846,N_33290);
nand U34212 (N_34212,N_33166,N_33350);
nand U34213 (N_34213,N_33549,N_33887);
or U34214 (N_34214,N_33677,N_33598);
nor U34215 (N_34215,N_33075,N_33167);
nor U34216 (N_34216,N_33961,N_33361);
nand U34217 (N_34217,N_33538,N_33486);
and U34218 (N_34218,N_33362,N_33482);
and U34219 (N_34219,N_33562,N_33403);
xnor U34220 (N_34220,N_33969,N_33901);
and U34221 (N_34221,N_33287,N_33588);
xnor U34222 (N_34222,N_33760,N_33890);
or U34223 (N_34223,N_33544,N_33879);
and U34224 (N_34224,N_33169,N_33013);
xnor U34225 (N_34225,N_33123,N_33174);
nand U34226 (N_34226,N_33719,N_33132);
or U34227 (N_34227,N_33703,N_33535);
or U34228 (N_34228,N_33834,N_33100);
nand U34229 (N_34229,N_33810,N_33953);
xnor U34230 (N_34230,N_33866,N_33987);
or U34231 (N_34231,N_33676,N_33122);
and U34232 (N_34232,N_33954,N_33370);
and U34233 (N_34233,N_33247,N_33430);
nand U34234 (N_34234,N_33553,N_33759);
nor U34235 (N_34235,N_33777,N_33788);
nand U34236 (N_34236,N_33227,N_33862);
nor U34237 (N_34237,N_33853,N_33039);
and U34238 (N_34238,N_33457,N_33057);
and U34239 (N_34239,N_33125,N_33949);
nor U34240 (N_34240,N_33393,N_33734);
nor U34241 (N_34241,N_33575,N_33493);
and U34242 (N_34242,N_33646,N_33071);
and U34243 (N_34243,N_33387,N_33313);
xnor U34244 (N_34244,N_33503,N_33121);
nor U34245 (N_34245,N_33960,N_33756);
or U34246 (N_34246,N_33469,N_33443);
xor U34247 (N_34247,N_33111,N_33139);
nand U34248 (N_34248,N_33340,N_33871);
nand U34249 (N_34249,N_33367,N_33789);
nor U34250 (N_34250,N_33965,N_33757);
xnor U34251 (N_34251,N_33651,N_33944);
nand U34252 (N_34252,N_33712,N_33930);
xnor U34253 (N_34253,N_33848,N_33011);
or U34254 (N_34254,N_33045,N_33479);
or U34255 (N_34255,N_33240,N_33926);
and U34256 (N_34256,N_33445,N_33883);
nor U34257 (N_34257,N_33799,N_33833);
nor U34258 (N_34258,N_33391,N_33674);
xnor U34259 (N_34259,N_33622,N_33390);
nor U34260 (N_34260,N_33921,N_33494);
or U34261 (N_34261,N_33214,N_33733);
and U34262 (N_34262,N_33090,N_33667);
nor U34263 (N_34263,N_33204,N_33196);
and U34264 (N_34264,N_33126,N_33316);
xnor U34265 (N_34265,N_33697,N_33621);
or U34266 (N_34266,N_33330,N_33437);
nor U34267 (N_34267,N_33333,N_33064);
or U34268 (N_34268,N_33134,N_33137);
xor U34269 (N_34269,N_33984,N_33790);
or U34270 (N_34270,N_33207,N_33791);
nor U34271 (N_34271,N_33283,N_33014);
and U34272 (N_34272,N_33537,N_33577);
nor U34273 (N_34273,N_33557,N_33783);
xor U34274 (N_34274,N_33119,N_33241);
nor U34275 (N_34275,N_33778,N_33262);
nand U34276 (N_34276,N_33421,N_33913);
or U34277 (N_34277,N_33067,N_33858);
nand U34278 (N_34278,N_33909,N_33683);
xor U34279 (N_34279,N_33824,N_33809);
or U34280 (N_34280,N_33678,N_33619);
or U34281 (N_34281,N_33082,N_33918);
xor U34282 (N_34282,N_33927,N_33767);
or U34283 (N_34283,N_33146,N_33427);
nand U34284 (N_34284,N_33113,N_33094);
nor U34285 (N_34285,N_33912,N_33568);
and U34286 (N_34286,N_33565,N_33814);
xnor U34287 (N_34287,N_33357,N_33334);
and U34288 (N_34288,N_33272,N_33520);
and U34289 (N_34289,N_33108,N_33701);
or U34290 (N_34290,N_33632,N_33135);
and U34291 (N_34291,N_33857,N_33542);
xor U34292 (N_34292,N_33656,N_33864);
nand U34293 (N_34293,N_33764,N_33409);
and U34294 (N_34294,N_33420,N_33897);
xor U34295 (N_34295,N_33920,N_33495);
or U34296 (N_34296,N_33225,N_33500);
or U34297 (N_34297,N_33066,N_33817);
nor U34298 (N_34298,N_33604,N_33534);
and U34299 (N_34299,N_33400,N_33768);
nor U34300 (N_34300,N_33012,N_33043);
nor U34301 (N_34301,N_33660,N_33815);
or U34302 (N_34302,N_33891,N_33488);
and U34303 (N_34303,N_33772,N_33223);
xor U34304 (N_34304,N_33679,N_33286);
nand U34305 (N_34305,N_33159,N_33321);
xnor U34306 (N_34306,N_33837,N_33120);
and U34307 (N_34307,N_33666,N_33185);
nand U34308 (N_34308,N_33038,N_33749);
nand U34309 (N_34309,N_33019,N_33839);
xor U34310 (N_34310,N_33976,N_33243);
xnor U34311 (N_34311,N_33658,N_33608);
nor U34312 (N_34312,N_33880,N_33484);
nand U34313 (N_34313,N_33291,N_33115);
xnor U34314 (N_34314,N_33885,N_33939);
nor U34315 (N_34315,N_33221,N_33707);
nor U34316 (N_34316,N_33161,N_33378);
and U34317 (N_34317,N_33724,N_33561);
nand U34318 (N_34318,N_33229,N_33260);
or U34319 (N_34319,N_33832,N_33181);
nand U34320 (N_34320,N_33780,N_33489);
and U34321 (N_34321,N_33625,N_33925);
or U34322 (N_34322,N_33836,N_33129);
nor U34323 (N_34323,N_33641,N_33319);
nor U34324 (N_34324,N_33352,N_33325);
and U34325 (N_34325,N_33342,N_33929);
or U34326 (N_34326,N_33740,N_33056);
nand U34327 (N_34327,N_33308,N_33353);
nor U34328 (N_34328,N_33852,N_33670);
xnor U34329 (N_34329,N_33869,N_33433);
nor U34330 (N_34330,N_33564,N_33004);
nand U34331 (N_34331,N_33359,N_33018);
xnor U34332 (N_34332,N_33311,N_33797);
nand U34333 (N_34333,N_33781,N_33155);
and U34334 (N_34334,N_33838,N_33914);
nand U34335 (N_34335,N_33055,N_33623);
xor U34336 (N_34336,N_33009,N_33054);
nor U34337 (N_34337,N_33058,N_33515);
and U34338 (N_34338,N_33189,N_33314);
xnor U34339 (N_34339,N_33793,N_33191);
nand U34340 (N_34340,N_33410,N_33947);
and U34341 (N_34341,N_33095,N_33555);
xor U34342 (N_34342,N_33124,N_33438);
and U34343 (N_34343,N_33595,N_33160);
nand U34344 (N_34344,N_33533,N_33519);
xor U34345 (N_34345,N_33744,N_33418);
nor U34346 (N_34346,N_33003,N_33397);
xor U34347 (N_34347,N_33886,N_33808);
or U34348 (N_34348,N_33402,N_33881);
or U34349 (N_34349,N_33036,N_33993);
nand U34350 (N_34350,N_33102,N_33372);
or U34351 (N_34351,N_33153,N_33751);
nor U34352 (N_34352,N_33524,N_33239);
nor U34353 (N_34353,N_33994,N_33002);
and U34354 (N_34354,N_33755,N_33190);
or U34355 (N_34355,N_33184,N_33737);
xor U34356 (N_34356,N_33404,N_33456);
nand U34357 (N_34357,N_33589,N_33978);
or U34358 (N_34358,N_33086,N_33945);
and U34359 (N_34359,N_33607,N_33175);
nor U34360 (N_34360,N_33158,N_33338);
nand U34361 (N_34361,N_33276,N_33510);
or U34362 (N_34362,N_33818,N_33851);
nor U34363 (N_34363,N_33423,N_33076);
or U34364 (N_34364,N_33203,N_33029);
nand U34365 (N_34365,N_33835,N_33844);
or U34366 (N_34366,N_33042,N_33206);
or U34367 (N_34367,N_33963,N_33841);
and U34368 (N_34368,N_33567,N_33601);
nand U34369 (N_34369,N_33138,N_33785);
or U34370 (N_34370,N_33265,N_33033);
and U34371 (N_34371,N_33389,N_33165);
nand U34372 (N_34372,N_33081,N_33531);
and U34373 (N_34373,N_33957,N_33692);
and U34374 (N_34374,N_33273,N_33826);
and U34375 (N_34375,N_33770,N_33176);
xnor U34376 (N_34376,N_33244,N_33653);
and U34377 (N_34377,N_33472,N_33475);
and U34378 (N_34378,N_33060,N_33010);
nand U34379 (N_34379,N_33231,N_33545);
nor U34380 (N_34380,N_33828,N_33037);
or U34381 (N_34381,N_33450,N_33508);
nor U34382 (N_34382,N_33899,N_33477);
and U34383 (N_34383,N_33647,N_33201);
and U34384 (N_34384,N_33843,N_33526);
xnor U34385 (N_34385,N_33827,N_33596);
or U34386 (N_34386,N_33708,N_33384);
nand U34387 (N_34387,N_33285,N_33150);
or U34388 (N_34388,N_33530,N_33592);
or U34389 (N_34389,N_33532,N_33085);
xnor U34390 (N_34390,N_33266,N_33496);
xor U34391 (N_34391,N_33979,N_33332);
or U34392 (N_34392,N_33578,N_33079);
nor U34393 (N_34393,N_33845,N_33868);
nand U34394 (N_34394,N_33257,N_33179);
xor U34395 (N_34395,N_33192,N_33915);
and U34396 (N_34396,N_33087,N_33695);
xor U34397 (N_34397,N_33005,N_33691);
nand U34398 (N_34398,N_33498,N_33617);
and U34399 (N_34399,N_33346,N_33341);
and U34400 (N_34400,N_33582,N_33186);
nor U34401 (N_34401,N_33279,N_33892);
xor U34402 (N_34402,N_33873,N_33673);
nand U34403 (N_34403,N_33907,N_33664);
or U34404 (N_34404,N_33459,N_33574);
nand U34405 (N_34405,N_33053,N_33964);
xor U34406 (N_34406,N_33505,N_33807);
nand U34407 (N_34407,N_33630,N_33248);
nand U34408 (N_34408,N_33382,N_33419);
and U34409 (N_34409,N_33263,N_33162);
or U34410 (N_34410,N_33233,N_33107);
nand U34411 (N_34411,N_33172,N_33748);
xor U34412 (N_34412,N_33587,N_33439);
and U34413 (N_34413,N_33613,N_33306);
and U34414 (N_34414,N_33048,N_33614);
nand U34415 (N_34415,N_33441,N_33584);
or U34416 (N_34416,N_33958,N_33327);
xnor U34417 (N_34417,N_33716,N_33117);
nor U34418 (N_34418,N_33518,N_33199);
nor U34419 (N_34419,N_33874,N_33548);
nor U34420 (N_34420,N_33870,N_33725);
or U34421 (N_34421,N_33212,N_33446);
or U34422 (N_34422,N_33543,N_33072);
xor U34423 (N_34423,N_33021,N_33911);
nor U34424 (N_34424,N_33988,N_33369);
xnor U34425 (N_34425,N_33424,N_33182);
nor U34426 (N_34426,N_33715,N_33487);
xor U34427 (N_34427,N_33637,N_33252);
or U34428 (N_34428,N_33245,N_33324);
or U34429 (N_34429,N_33754,N_33228);
or U34430 (N_34430,N_33982,N_33302);
nor U34431 (N_34431,N_33412,N_33747);
nor U34432 (N_34432,N_33968,N_33784);
nand U34433 (N_34433,N_33903,N_33629);
and U34434 (N_34434,N_33860,N_33971);
and U34435 (N_34435,N_33077,N_33742);
or U34436 (N_34436,N_33659,N_33408);
xnor U34437 (N_34437,N_33298,N_33106);
and U34438 (N_34438,N_33133,N_33023);
nand U34439 (N_34439,N_33682,N_33296);
and U34440 (N_34440,N_33829,N_33347);
or U34441 (N_34441,N_33847,N_33606);
or U34442 (N_34442,N_33464,N_33271);
and U34443 (N_34443,N_33422,N_33478);
nor U34444 (N_34444,N_33941,N_33205);
and U34445 (N_34445,N_33194,N_33267);
nor U34446 (N_34446,N_33242,N_33442);
and U34447 (N_34447,N_33611,N_33600);
nand U34448 (N_34448,N_33769,N_33025);
xor U34449 (N_34449,N_33236,N_33699);
xor U34450 (N_34450,N_33745,N_33618);
nand U34451 (N_34451,N_33507,N_33020);
and U34452 (N_34452,N_33452,N_33358);
nand U34453 (N_34453,N_33292,N_33177);
xor U34454 (N_34454,N_33396,N_33097);
nand U34455 (N_34455,N_33345,N_33485);
nor U34456 (N_34456,N_33375,N_33130);
nand U34457 (N_34457,N_33586,N_33935);
and U34458 (N_34458,N_33936,N_33089);
xnor U34459 (N_34459,N_33644,N_33383);
nor U34460 (N_34460,N_33943,N_33499);
or U34461 (N_34461,N_33796,N_33380);
or U34462 (N_34462,N_33861,N_33455);
nand U34463 (N_34463,N_33795,N_33983);
nand U34464 (N_34464,N_33758,N_33615);
or U34465 (N_34465,N_33610,N_33000);
nand U34466 (N_34466,N_33626,N_33501);
or U34467 (N_34467,N_33794,N_33322);
or U34468 (N_34468,N_33151,N_33007);
and U34469 (N_34469,N_33432,N_33171);
nor U34470 (N_34470,N_33407,N_33168);
and U34471 (N_34471,N_33512,N_33635);
and U34472 (N_34472,N_33008,N_33593);
xnor U34473 (N_34473,N_33514,N_33905);
xor U34474 (N_34474,N_33270,N_33816);
xor U34475 (N_34475,N_33473,N_33293);
nand U34476 (N_34476,N_33395,N_33289);
and U34477 (N_34477,N_33878,N_33417);
and U34478 (N_34478,N_33528,N_33466);
xnor U34479 (N_34479,N_33386,N_33732);
or U34480 (N_34480,N_33392,N_33779);
nor U34481 (N_34481,N_33540,N_33643);
nor U34482 (N_34482,N_33216,N_33823);
and U34483 (N_34483,N_33952,N_33812);
nor U34484 (N_34484,N_33147,N_33986);
nor U34485 (N_34485,N_33049,N_33088);
nand U34486 (N_34486,N_33399,N_33959);
nand U34487 (N_34487,N_33529,N_33763);
or U34488 (N_34488,N_33906,N_33842);
and U34489 (N_34489,N_33096,N_33476);
xnor U34490 (N_34490,N_33525,N_33739);
nor U34491 (N_34491,N_33856,N_33730);
or U34492 (N_34492,N_33331,N_33721);
or U34493 (N_34493,N_33426,N_33819);
nor U34494 (N_34494,N_33368,N_33649);
or U34495 (N_34495,N_33211,N_33282);
and U34496 (N_34496,N_33956,N_33684);
or U34497 (N_34497,N_33193,N_33385);
nand U34498 (N_34498,N_33775,N_33894);
and U34499 (N_34499,N_33462,N_33180);
nand U34500 (N_34500,N_33977,N_33725);
xnor U34501 (N_34501,N_33383,N_33806);
or U34502 (N_34502,N_33248,N_33710);
xor U34503 (N_34503,N_33809,N_33947);
and U34504 (N_34504,N_33052,N_33025);
and U34505 (N_34505,N_33604,N_33478);
and U34506 (N_34506,N_33950,N_33185);
nand U34507 (N_34507,N_33899,N_33853);
nand U34508 (N_34508,N_33368,N_33699);
and U34509 (N_34509,N_33923,N_33660);
xnor U34510 (N_34510,N_33915,N_33291);
or U34511 (N_34511,N_33845,N_33976);
nor U34512 (N_34512,N_33525,N_33675);
and U34513 (N_34513,N_33109,N_33101);
or U34514 (N_34514,N_33311,N_33232);
nor U34515 (N_34515,N_33503,N_33575);
nor U34516 (N_34516,N_33901,N_33238);
nand U34517 (N_34517,N_33033,N_33417);
xnor U34518 (N_34518,N_33631,N_33978);
or U34519 (N_34519,N_33417,N_33412);
nand U34520 (N_34520,N_33650,N_33397);
xnor U34521 (N_34521,N_33603,N_33452);
or U34522 (N_34522,N_33531,N_33215);
nor U34523 (N_34523,N_33255,N_33454);
nand U34524 (N_34524,N_33101,N_33583);
xor U34525 (N_34525,N_33536,N_33941);
or U34526 (N_34526,N_33973,N_33143);
and U34527 (N_34527,N_33129,N_33286);
or U34528 (N_34528,N_33018,N_33799);
xor U34529 (N_34529,N_33529,N_33141);
and U34530 (N_34530,N_33916,N_33595);
nand U34531 (N_34531,N_33398,N_33245);
nor U34532 (N_34532,N_33866,N_33373);
and U34533 (N_34533,N_33519,N_33500);
nand U34534 (N_34534,N_33401,N_33918);
nor U34535 (N_34535,N_33066,N_33735);
xnor U34536 (N_34536,N_33041,N_33868);
xnor U34537 (N_34537,N_33254,N_33104);
xnor U34538 (N_34538,N_33193,N_33816);
and U34539 (N_34539,N_33365,N_33119);
nand U34540 (N_34540,N_33049,N_33066);
xor U34541 (N_34541,N_33534,N_33944);
nor U34542 (N_34542,N_33887,N_33066);
xnor U34543 (N_34543,N_33826,N_33869);
or U34544 (N_34544,N_33680,N_33062);
nor U34545 (N_34545,N_33363,N_33842);
xor U34546 (N_34546,N_33646,N_33170);
or U34547 (N_34547,N_33142,N_33792);
xnor U34548 (N_34548,N_33992,N_33175);
nor U34549 (N_34549,N_33990,N_33060);
nand U34550 (N_34550,N_33051,N_33492);
nand U34551 (N_34551,N_33410,N_33569);
or U34552 (N_34552,N_33409,N_33430);
and U34553 (N_34553,N_33036,N_33558);
or U34554 (N_34554,N_33703,N_33644);
xnor U34555 (N_34555,N_33806,N_33140);
xor U34556 (N_34556,N_33582,N_33598);
and U34557 (N_34557,N_33942,N_33384);
and U34558 (N_34558,N_33412,N_33099);
xor U34559 (N_34559,N_33525,N_33536);
xnor U34560 (N_34560,N_33938,N_33029);
xor U34561 (N_34561,N_33997,N_33516);
or U34562 (N_34562,N_33699,N_33614);
nand U34563 (N_34563,N_33371,N_33518);
nor U34564 (N_34564,N_33796,N_33314);
or U34565 (N_34565,N_33767,N_33344);
xor U34566 (N_34566,N_33094,N_33032);
nor U34567 (N_34567,N_33791,N_33568);
nor U34568 (N_34568,N_33195,N_33391);
and U34569 (N_34569,N_33041,N_33112);
xnor U34570 (N_34570,N_33168,N_33795);
or U34571 (N_34571,N_33334,N_33172);
and U34572 (N_34572,N_33957,N_33909);
xor U34573 (N_34573,N_33682,N_33303);
nand U34574 (N_34574,N_33770,N_33386);
nor U34575 (N_34575,N_33411,N_33332);
and U34576 (N_34576,N_33459,N_33086);
or U34577 (N_34577,N_33799,N_33045);
nand U34578 (N_34578,N_33073,N_33111);
and U34579 (N_34579,N_33962,N_33846);
xor U34580 (N_34580,N_33223,N_33015);
xnor U34581 (N_34581,N_33992,N_33553);
and U34582 (N_34582,N_33309,N_33204);
or U34583 (N_34583,N_33931,N_33253);
xor U34584 (N_34584,N_33220,N_33532);
nor U34585 (N_34585,N_33341,N_33945);
and U34586 (N_34586,N_33199,N_33250);
and U34587 (N_34587,N_33753,N_33870);
nand U34588 (N_34588,N_33848,N_33306);
nand U34589 (N_34589,N_33865,N_33907);
and U34590 (N_34590,N_33870,N_33215);
and U34591 (N_34591,N_33042,N_33967);
nand U34592 (N_34592,N_33721,N_33616);
and U34593 (N_34593,N_33596,N_33590);
or U34594 (N_34594,N_33226,N_33687);
or U34595 (N_34595,N_33192,N_33252);
xor U34596 (N_34596,N_33614,N_33330);
and U34597 (N_34597,N_33692,N_33672);
nor U34598 (N_34598,N_33027,N_33172);
xnor U34599 (N_34599,N_33859,N_33813);
xor U34600 (N_34600,N_33325,N_33436);
xor U34601 (N_34601,N_33340,N_33878);
or U34602 (N_34602,N_33433,N_33206);
nand U34603 (N_34603,N_33099,N_33696);
and U34604 (N_34604,N_33211,N_33304);
or U34605 (N_34605,N_33929,N_33777);
and U34606 (N_34606,N_33659,N_33231);
nor U34607 (N_34607,N_33922,N_33288);
and U34608 (N_34608,N_33018,N_33738);
nor U34609 (N_34609,N_33698,N_33281);
and U34610 (N_34610,N_33275,N_33554);
xnor U34611 (N_34611,N_33225,N_33663);
nand U34612 (N_34612,N_33822,N_33712);
nand U34613 (N_34613,N_33174,N_33254);
or U34614 (N_34614,N_33312,N_33426);
and U34615 (N_34615,N_33899,N_33327);
xor U34616 (N_34616,N_33502,N_33715);
or U34617 (N_34617,N_33079,N_33889);
xor U34618 (N_34618,N_33592,N_33366);
nor U34619 (N_34619,N_33109,N_33219);
nand U34620 (N_34620,N_33851,N_33261);
nand U34621 (N_34621,N_33708,N_33064);
nor U34622 (N_34622,N_33295,N_33190);
xnor U34623 (N_34623,N_33693,N_33323);
nor U34624 (N_34624,N_33510,N_33002);
nand U34625 (N_34625,N_33983,N_33259);
nand U34626 (N_34626,N_33496,N_33408);
and U34627 (N_34627,N_33820,N_33183);
and U34628 (N_34628,N_33094,N_33557);
or U34629 (N_34629,N_33383,N_33833);
or U34630 (N_34630,N_33983,N_33135);
or U34631 (N_34631,N_33661,N_33391);
xor U34632 (N_34632,N_33284,N_33014);
nor U34633 (N_34633,N_33965,N_33001);
nand U34634 (N_34634,N_33347,N_33334);
xor U34635 (N_34635,N_33759,N_33472);
nand U34636 (N_34636,N_33098,N_33271);
or U34637 (N_34637,N_33119,N_33303);
or U34638 (N_34638,N_33963,N_33965);
nand U34639 (N_34639,N_33120,N_33623);
or U34640 (N_34640,N_33360,N_33661);
or U34641 (N_34641,N_33918,N_33359);
nand U34642 (N_34642,N_33698,N_33018);
nor U34643 (N_34643,N_33958,N_33889);
and U34644 (N_34644,N_33177,N_33775);
nor U34645 (N_34645,N_33312,N_33406);
and U34646 (N_34646,N_33448,N_33515);
or U34647 (N_34647,N_33497,N_33795);
nor U34648 (N_34648,N_33958,N_33045);
nor U34649 (N_34649,N_33215,N_33838);
or U34650 (N_34650,N_33220,N_33827);
nand U34651 (N_34651,N_33456,N_33869);
nand U34652 (N_34652,N_33229,N_33700);
and U34653 (N_34653,N_33408,N_33449);
and U34654 (N_34654,N_33240,N_33261);
nor U34655 (N_34655,N_33117,N_33595);
and U34656 (N_34656,N_33815,N_33035);
nor U34657 (N_34657,N_33276,N_33788);
and U34658 (N_34658,N_33067,N_33314);
and U34659 (N_34659,N_33660,N_33233);
nor U34660 (N_34660,N_33014,N_33458);
or U34661 (N_34661,N_33287,N_33109);
nor U34662 (N_34662,N_33212,N_33014);
nand U34663 (N_34663,N_33273,N_33170);
or U34664 (N_34664,N_33359,N_33130);
or U34665 (N_34665,N_33315,N_33558);
nand U34666 (N_34666,N_33736,N_33337);
nand U34667 (N_34667,N_33983,N_33286);
nor U34668 (N_34668,N_33389,N_33476);
xor U34669 (N_34669,N_33367,N_33491);
or U34670 (N_34670,N_33007,N_33519);
xor U34671 (N_34671,N_33738,N_33118);
and U34672 (N_34672,N_33522,N_33777);
and U34673 (N_34673,N_33720,N_33838);
or U34674 (N_34674,N_33198,N_33956);
nand U34675 (N_34675,N_33678,N_33381);
or U34676 (N_34676,N_33601,N_33266);
nor U34677 (N_34677,N_33107,N_33797);
or U34678 (N_34678,N_33710,N_33975);
nor U34679 (N_34679,N_33076,N_33999);
nor U34680 (N_34680,N_33292,N_33349);
nor U34681 (N_34681,N_33702,N_33057);
and U34682 (N_34682,N_33115,N_33820);
nor U34683 (N_34683,N_33900,N_33903);
or U34684 (N_34684,N_33719,N_33574);
xor U34685 (N_34685,N_33600,N_33882);
nor U34686 (N_34686,N_33199,N_33630);
or U34687 (N_34687,N_33166,N_33046);
or U34688 (N_34688,N_33746,N_33266);
or U34689 (N_34689,N_33849,N_33533);
nor U34690 (N_34690,N_33890,N_33652);
or U34691 (N_34691,N_33018,N_33037);
or U34692 (N_34692,N_33430,N_33677);
and U34693 (N_34693,N_33983,N_33394);
nand U34694 (N_34694,N_33625,N_33263);
xnor U34695 (N_34695,N_33071,N_33716);
xnor U34696 (N_34696,N_33528,N_33585);
nand U34697 (N_34697,N_33976,N_33953);
nand U34698 (N_34698,N_33318,N_33754);
and U34699 (N_34699,N_33218,N_33937);
nor U34700 (N_34700,N_33979,N_33432);
nand U34701 (N_34701,N_33884,N_33438);
nor U34702 (N_34702,N_33977,N_33805);
xor U34703 (N_34703,N_33317,N_33961);
nor U34704 (N_34704,N_33308,N_33163);
or U34705 (N_34705,N_33862,N_33030);
and U34706 (N_34706,N_33717,N_33951);
xnor U34707 (N_34707,N_33899,N_33919);
and U34708 (N_34708,N_33863,N_33777);
or U34709 (N_34709,N_33621,N_33138);
and U34710 (N_34710,N_33476,N_33876);
and U34711 (N_34711,N_33660,N_33320);
and U34712 (N_34712,N_33771,N_33793);
and U34713 (N_34713,N_33718,N_33663);
or U34714 (N_34714,N_33934,N_33080);
nand U34715 (N_34715,N_33495,N_33134);
or U34716 (N_34716,N_33927,N_33292);
or U34717 (N_34717,N_33659,N_33671);
nor U34718 (N_34718,N_33571,N_33141);
xor U34719 (N_34719,N_33809,N_33141);
or U34720 (N_34720,N_33196,N_33531);
xnor U34721 (N_34721,N_33408,N_33841);
or U34722 (N_34722,N_33492,N_33183);
xnor U34723 (N_34723,N_33300,N_33956);
and U34724 (N_34724,N_33571,N_33909);
nor U34725 (N_34725,N_33886,N_33166);
nor U34726 (N_34726,N_33364,N_33069);
nor U34727 (N_34727,N_33500,N_33865);
or U34728 (N_34728,N_33312,N_33113);
nand U34729 (N_34729,N_33952,N_33287);
nand U34730 (N_34730,N_33224,N_33688);
and U34731 (N_34731,N_33200,N_33385);
nor U34732 (N_34732,N_33012,N_33746);
and U34733 (N_34733,N_33467,N_33952);
xnor U34734 (N_34734,N_33224,N_33993);
or U34735 (N_34735,N_33751,N_33591);
nand U34736 (N_34736,N_33075,N_33579);
xnor U34737 (N_34737,N_33144,N_33083);
or U34738 (N_34738,N_33584,N_33445);
or U34739 (N_34739,N_33932,N_33002);
nor U34740 (N_34740,N_33409,N_33703);
xnor U34741 (N_34741,N_33640,N_33098);
nand U34742 (N_34742,N_33688,N_33271);
and U34743 (N_34743,N_33804,N_33780);
nor U34744 (N_34744,N_33178,N_33127);
xnor U34745 (N_34745,N_33962,N_33730);
and U34746 (N_34746,N_33837,N_33131);
nor U34747 (N_34747,N_33937,N_33087);
xnor U34748 (N_34748,N_33780,N_33210);
and U34749 (N_34749,N_33459,N_33717);
and U34750 (N_34750,N_33885,N_33446);
and U34751 (N_34751,N_33722,N_33455);
nand U34752 (N_34752,N_33198,N_33934);
nand U34753 (N_34753,N_33015,N_33074);
xnor U34754 (N_34754,N_33788,N_33106);
nand U34755 (N_34755,N_33564,N_33068);
or U34756 (N_34756,N_33803,N_33149);
or U34757 (N_34757,N_33298,N_33439);
nand U34758 (N_34758,N_33260,N_33855);
nand U34759 (N_34759,N_33476,N_33517);
nand U34760 (N_34760,N_33315,N_33367);
nand U34761 (N_34761,N_33993,N_33886);
and U34762 (N_34762,N_33142,N_33307);
xor U34763 (N_34763,N_33490,N_33222);
and U34764 (N_34764,N_33248,N_33879);
or U34765 (N_34765,N_33329,N_33472);
nand U34766 (N_34766,N_33196,N_33275);
and U34767 (N_34767,N_33782,N_33260);
nor U34768 (N_34768,N_33923,N_33313);
or U34769 (N_34769,N_33854,N_33733);
or U34770 (N_34770,N_33999,N_33288);
or U34771 (N_34771,N_33709,N_33573);
or U34772 (N_34772,N_33066,N_33162);
and U34773 (N_34773,N_33541,N_33257);
or U34774 (N_34774,N_33823,N_33166);
or U34775 (N_34775,N_33788,N_33954);
and U34776 (N_34776,N_33222,N_33581);
or U34777 (N_34777,N_33292,N_33612);
nand U34778 (N_34778,N_33182,N_33585);
nor U34779 (N_34779,N_33648,N_33176);
or U34780 (N_34780,N_33797,N_33548);
xnor U34781 (N_34781,N_33266,N_33994);
and U34782 (N_34782,N_33135,N_33107);
and U34783 (N_34783,N_33583,N_33669);
xor U34784 (N_34784,N_33842,N_33146);
nor U34785 (N_34785,N_33918,N_33814);
nand U34786 (N_34786,N_33660,N_33540);
nand U34787 (N_34787,N_33014,N_33895);
nor U34788 (N_34788,N_33535,N_33577);
nand U34789 (N_34789,N_33276,N_33265);
xnor U34790 (N_34790,N_33338,N_33396);
nor U34791 (N_34791,N_33920,N_33205);
nand U34792 (N_34792,N_33622,N_33420);
xnor U34793 (N_34793,N_33531,N_33471);
nor U34794 (N_34794,N_33193,N_33685);
xor U34795 (N_34795,N_33960,N_33323);
or U34796 (N_34796,N_33648,N_33959);
nor U34797 (N_34797,N_33015,N_33732);
xor U34798 (N_34798,N_33233,N_33374);
nor U34799 (N_34799,N_33996,N_33336);
and U34800 (N_34800,N_33109,N_33402);
xor U34801 (N_34801,N_33727,N_33587);
or U34802 (N_34802,N_33505,N_33267);
nor U34803 (N_34803,N_33777,N_33508);
or U34804 (N_34804,N_33174,N_33427);
nand U34805 (N_34805,N_33868,N_33619);
or U34806 (N_34806,N_33666,N_33838);
or U34807 (N_34807,N_33865,N_33878);
and U34808 (N_34808,N_33846,N_33277);
or U34809 (N_34809,N_33738,N_33331);
nor U34810 (N_34810,N_33868,N_33568);
or U34811 (N_34811,N_33359,N_33916);
and U34812 (N_34812,N_33138,N_33400);
nand U34813 (N_34813,N_33965,N_33181);
nor U34814 (N_34814,N_33359,N_33161);
xor U34815 (N_34815,N_33363,N_33343);
nand U34816 (N_34816,N_33330,N_33300);
nor U34817 (N_34817,N_33388,N_33044);
nor U34818 (N_34818,N_33275,N_33514);
or U34819 (N_34819,N_33073,N_33541);
nand U34820 (N_34820,N_33947,N_33908);
nor U34821 (N_34821,N_33193,N_33549);
nand U34822 (N_34822,N_33582,N_33853);
xor U34823 (N_34823,N_33941,N_33800);
nand U34824 (N_34824,N_33350,N_33921);
and U34825 (N_34825,N_33828,N_33857);
xor U34826 (N_34826,N_33727,N_33816);
nor U34827 (N_34827,N_33840,N_33737);
nor U34828 (N_34828,N_33666,N_33268);
or U34829 (N_34829,N_33823,N_33042);
nor U34830 (N_34830,N_33617,N_33454);
nor U34831 (N_34831,N_33637,N_33522);
nand U34832 (N_34832,N_33560,N_33710);
xor U34833 (N_34833,N_33018,N_33012);
and U34834 (N_34834,N_33776,N_33823);
nor U34835 (N_34835,N_33405,N_33958);
nand U34836 (N_34836,N_33900,N_33866);
xor U34837 (N_34837,N_33084,N_33175);
nor U34838 (N_34838,N_33329,N_33208);
and U34839 (N_34839,N_33895,N_33823);
nor U34840 (N_34840,N_33691,N_33187);
and U34841 (N_34841,N_33368,N_33983);
or U34842 (N_34842,N_33307,N_33077);
nor U34843 (N_34843,N_33222,N_33242);
xor U34844 (N_34844,N_33252,N_33829);
nand U34845 (N_34845,N_33928,N_33213);
nand U34846 (N_34846,N_33375,N_33752);
nor U34847 (N_34847,N_33412,N_33224);
nand U34848 (N_34848,N_33465,N_33252);
and U34849 (N_34849,N_33873,N_33715);
xnor U34850 (N_34850,N_33527,N_33087);
and U34851 (N_34851,N_33343,N_33639);
nor U34852 (N_34852,N_33630,N_33903);
or U34853 (N_34853,N_33680,N_33561);
nand U34854 (N_34854,N_33567,N_33261);
nand U34855 (N_34855,N_33354,N_33972);
nand U34856 (N_34856,N_33031,N_33630);
nand U34857 (N_34857,N_33895,N_33148);
nand U34858 (N_34858,N_33022,N_33073);
or U34859 (N_34859,N_33456,N_33736);
or U34860 (N_34860,N_33711,N_33885);
xor U34861 (N_34861,N_33170,N_33830);
nor U34862 (N_34862,N_33320,N_33782);
or U34863 (N_34863,N_33913,N_33670);
nor U34864 (N_34864,N_33757,N_33234);
nor U34865 (N_34865,N_33363,N_33176);
and U34866 (N_34866,N_33385,N_33630);
or U34867 (N_34867,N_33533,N_33336);
nand U34868 (N_34868,N_33248,N_33401);
nor U34869 (N_34869,N_33664,N_33278);
nor U34870 (N_34870,N_33551,N_33285);
and U34871 (N_34871,N_33072,N_33538);
and U34872 (N_34872,N_33611,N_33268);
nor U34873 (N_34873,N_33448,N_33283);
or U34874 (N_34874,N_33719,N_33457);
nand U34875 (N_34875,N_33804,N_33424);
and U34876 (N_34876,N_33255,N_33092);
or U34877 (N_34877,N_33611,N_33403);
nand U34878 (N_34878,N_33287,N_33281);
nand U34879 (N_34879,N_33237,N_33324);
and U34880 (N_34880,N_33761,N_33227);
nor U34881 (N_34881,N_33737,N_33899);
or U34882 (N_34882,N_33661,N_33878);
or U34883 (N_34883,N_33741,N_33937);
xnor U34884 (N_34884,N_33184,N_33577);
nand U34885 (N_34885,N_33567,N_33326);
or U34886 (N_34886,N_33028,N_33157);
and U34887 (N_34887,N_33243,N_33066);
and U34888 (N_34888,N_33178,N_33407);
nor U34889 (N_34889,N_33816,N_33648);
and U34890 (N_34890,N_33593,N_33647);
and U34891 (N_34891,N_33594,N_33132);
xor U34892 (N_34892,N_33622,N_33563);
xnor U34893 (N_34893,N_33714,N_33762);
or U34894 (N_34894,N_33423,N_33992);
or U34895 (N_34895,N_33382,N_33664);
and U34896 (N_34896,N_33932,N_33185);
xnor U34897 (N_34897,N_33526,N_33463);
nand U34898 (N_34898,N_33501,N_33377);
and U34899 (N_34899,N_33898,N_33874);
nor U34900 (N_34900,N_33876,N_33881);
xor U34901 (N_34901,N_33028,N_33420);
xnor U34902 (N_34902,N_33647,N_33783);
nand U34903 (N_34903,N_33141,N_33599);
xor U34904 (N_34904,N_33570,N_33758);
xor U34905 (N_34905,N_33560,N_33343);
or U34906 (N_34906,N_33539,N_33149);
and U34907 (N_34907,N_33927,N_33010);
xor U34908 (N_34908,N_33131,N_33913);
xnor U34909 (N_34909,N_33784,N_33311);
and U34910 (N_34910,N_33034,N_33813);
and U34911 (N_34911,N_33793,N_33224);
nor U34912 (N_34912,N_33865,N_33312);
and U34913 (N_34913,N_33808,N_33927);
or U34914 (N_34914,N_33013,N_33737);
or U34915 (N_34915,N_33872,N_33078);
xor U34916 (N_34916,N_33957,N_33501);
xor U34917 (N_34917,N_33560,N_33030);
xnor U34918 (N_34918,N_33179,N_33562);
xor U34919 (N_34919,N_33000,N_33238);
and U34920 (N_34920,N_33814,N_33297);
or U34921 (N_34921,N_33312,N_33784);
and U34922 (N_34922,N_33020,N_33953);
nand U34923 (N_34923,N_33238,N_33132);
or U34924 (N_34924,N_33662,N_33294);
xor U34925 (N_34925,N_33157,N_33462);
nand U34926 (N_34926,N_33132,N_33511);
or U34927 (N_34927,N_33600,N_33403);
xnor U34928 (N_34928,N_33770,N_33329);
or U34929 (N_34929,N_33430,N_33641);
xnor U34930 (N_34930,N_33696,N_33388);
and U34931 (N_34931,N_33608,N_33350);
and U34932 (N_34932,N_33488,N_33345);
nor U34933 (N_34933,N_33020,N_33116);
or U34934 (N_34934,N_33282,N_33705);
nor U34935 (N_34935,N_33006,N_33632);
nand U34936 (N_34936,N_33719,N_33184);
xor U34937 (N_34937,N_33364,N_33395);
nor U34938 (N_34938,N_33598,N_33508);
nand U34939 (N_34939,N_33801,N_33035);
or U34940 (N_34940,N_33018,N_33821);
nand U34941 (N_34941,N_33119,N_33215);
nand U34942 (N_34942,N_33819,N_33701);
nand U34943 (N_34943,N_33965,N_33533);
xnor U34944 (N_34944,N_33958,N_33858);
xor U34945 (N_34945,N_33220,N_33282);
nand U34946 (N_34946,N_33429,N_33243);
or U34947 (N_34947,N_33264,N_33004);
nand U34948 (N_34948,N_33171,N_33465);
xnor U34949 (N_34949,N_33836,N_33705);
or U34950 (N_34950,N_33429,N_33911);
or U34951 (N_34951,N_33840,N_33236);
or U34952 (N_34952,N_33055,N_33264);
or U34953 (N_34953,N_33346,N_33977);
nor U34954 (N_34954,N_33232,N_33790);
nand U34955 (N_34955,N_33120,N_33660);
or U34956 (N_34956,N_33429,N_33117);
and U34957 (N_34957,N_33403,N_33048);
nand U34958 (N_34958,N_33749,N_33049);
and U34959 (N_34959,N_33066,N_33187);
nand U34960 (N_34960,N_33542,N_33379);
or U34961 (N_34961,N_33405,N_33047);
nand U34962 (N_34962,N_33646,N_33173);
xnor U34963 (N_34963,N_33251,N_33484);
xnor U34964 (N_34964,N_33951,N_33973);
nand U34965 (N_34965,N_33170,N_33454);
and U34966 (N_34966,N_33535,N_33851);
nor U34967 (N_34967,N_33437,N_33238);
xnor U34968 (N_34968,N_33935,N_33361);
or U34969 (N_34969,N_33263,N_33564);
or U34970 (N_34970,N_33472,N_33992);
or U34971 (N_34971,N_33746,N_33813);
or U34972 (N_34972,N_33772,N_33528);
or U34973 (N_34973,N_33313,N_33113);
nand U34974 (N_34974,N_33259,N_33366);
nand U34975 (N_34975,N_33612,N_33635);
and U34976 (N_34976,N_33802,N_33506);
or U34977 (N_34977,N_33254,N_33555);
xor U34978 (N_34978,N_33179,N_33857);
nor U34979 (N_34979,N_33422,N_33634);
nand U34980 (N_34980,N_33623,N_33810);
xor U34981 (N_34981,N_33676,N_33702);
nand U34982 (N_34982,N_33353,N_33377);
or U34983 (N_34983,N_33103,N_33276);
xnor U34984 (N_34984,N_33534,N_33277);
nand U34985 (N_34985,N_33193,N_33903);
nand U34986 (N_34986,N_33572,N_33992);
xnor U34987 (N_34987,N_33442,N_33643);
or U34988 (N_34988,N_33551,N_33381);
xnor U34989 (N_34989,N_33322,N_33911);
or U34990 (N_34990,N_33291,N_33484);
nand U34991 (N_34991,N_33022,N_33313);
xnor U34992 (N_34992,N_33903,N_33633);
or U34993 (N_34993,N_33231,N_33828);
xnor U34994 (N_34994,N_33967,N_33631);
xnor U34995 (N_34995,N_33212,N_33177);
nand U34996 (N_34996,N_33439,N_33421);
xor U34997 (N_34997,N_33594,N_33090);
nand U34998 (N_34998,N_33004,N_33495);
and U34999 (N_34999,N_33140,N_33053);
nor U35000 (N_35000,N_34266,N_34991);
nand U35001 (N_35001,N_34234,N_34721);
xor U35002 (N_35002,N_34667,N_34072);
nor U35003 (N_35003,N_34785,N_34094);
nand U35004 (N_35004,N_34863,N_34604);
or U35005 (N_35005,N_34570,N_34079);
or U35006 (N_35006,N_34673,N_34484);
or U35007 (N_35007,N_34766,N_34846);
or U35008 (N_35008,N_34284,N_34262);
or U35009 (N_35009,N_34440,N_34985);
xor U35010 (N_35010,N_34021,N_34066);
xnor U35011 (N_35011,N_34706,N_34314);
or U35012 (N_35012,N_34018,N_34779);
and U35013 (N_35013,N_34416,N_34456);
xnor U35014 (N_35014,N_34660,N_34315);
nand U35015 (N_35015,N_34595,N_34814);
or U35016 (N_35016,N_34940,N_34950);
nor U35017 (N_35017,N_34609,N_34992);
nor U35018 (N_35018,N_34014,N_34689);
and U35019 (N_35019,N_34652,N_34904);
or U35020 (N_35020,N_34822,N_34053);
nand U35021 (N_35021,N_34541,N_34327);
nand U35022 (N_35022,N_34168,N_34463);
xnor U35023 (N_35023,N_34600,N_34573);
or U35024 (N_35024,N_34834,N_34624);
and U35025 (N_35025,N_34441,N_34287);
and U35026 (N_35026,N_34843,N_34974);
xor U35027 (N_35027,N_34251,N_34102);
and U35028 (N_35028,N_34181,N_34349);
or U35029 (N_35029,N_34000,N_34444);
or U35030 (N_35030,N_34049,N_34828);
xor U35031 (N_35031,N_34061,N_34111);
xor U35032 (N_35032,N_34684,N_34083);
xnor U35033 (N_35033,N_34330,N_34382);
xor U35034 (N_35034,N_34644,N_34119);
nor U35035 (N_35035,N_34558,N_34362);
xnor U35036 (N_35036,N_34656,N_34242);
and U35037 (N_35037,N_34140,N_34035);
nor U35038 (N_35038,N_34756,N_34258);
and U35039 (N_35039,N_34998,N_34492);
or U35040 (N_35040,N_34338,N_34618);
xor U35041 (N_35041,N_34322,N_34961);
or U35042 (N_35042,N_34312,N_34276);
nor U35043 (N_35043,N_34143,N_34890);
and U35044 (N_35044,N_34177,N_34336);
and U35045 (N_35045,N_34156,N_34980);
and U35046 (N_35046,N_34979,N_34566);
and U35047 (N_35047,N_34506,N_34200);
and U35048 (N_35048,N_34291,N_34400);
or U35049 (N_35049,N_34132,N_34932);
xor U35050 (N_35050,N_34725,N_34575);
nand U35051 (N_35051,N_34678,N_34305);
or U35052 (N_35052,N_34759,N_34659);
and U35053 (N_35053,N_34183,N_34879);
or U35054 (N_35054,N_34058,N_34044);
and U35055 (N_35055,N_34942,N_34220);
and U35056 (N_35056,N_34219,N_34641);
nor U35057 (N_35057,N_34157,N_34477);
nand U35058 (N_35058,N_34211,N_34135);
or U35059 (N_35059,N_34374,N_34643);
or U35060 (N_35060,N_34622,N_34454);
nand U35061 (N_35061,N_34605,N_34743);
nor U35062 (N_35062,N_34951,N_34538);
and U35063 (N_35063,N_34277,N_34013);
xor U35064 (N_35064,N_34639,N_34474);
xnor U35065 (N_35065,N_34771,N_34246);
nor U35066 (N_35066,N_34762,N_34303);
xnor U35067 (N_35067,N_34707,N_34532);
and U35068 (N_35068,N_34155,N_34994);
xnor U35069 (N_35069,N_34468,N_34414);
and U35070 (N_35070,N_34597,N_34579);
nand U35071 (N_35071,N_34626,N_34473);
xnor U35072 (N_35072,N_34813,N_34872);
or U35073 (N_35073,N_34955,N_34439);
and U35074 (N_35074,N_34380,N_34623);
xnor U35075 (N_35075,N_34628,N_34098);
or U35076 (N_35076,N_34017,N_34563);
and U35077 (N_35077,N_34934,N_34911);
nor U35078 (N_35078,N_34744,N_34255);
xnor U35079 (N_35079,N_34244,N_34329);
or U35080 (N_35080,N_34290,N_34052);
nand U35081 (N_35081,N_34534,N_34669);
nand U35082 (N_35082,N_34580,N_34043);
nor U35083 (N_35083,N_34077,N_34675);
xor U35084 (N_35084,N_34587,N_34524);
xnor U35085 (N_35085,N_34420,N_34801);
and U35086 (N_35086,N_34431,N_34897);
nor U35087 (N_35087,N_34523,N_34106);
nor U35088 (N_35088,N_34100,N_34685);
or U35089 (N_35089,N_34428,N_34032);
nand U35090 (N_35090,N_34356,N_34769);
and U35091 (N_35091,N_34105,N_34496);
nor U35092 (N_35092,N_34245,N_34621);
nor U35093 (N_35093,N_34114,N_34283);
or U35094 (N_35094,N_34778,N_34693);
or U35095 (N_35095,N_34179,N_34003);
nand U35096 (N_35096,N_34895,N_34426);
xor U35097 (N_35097,N_34434,N_34185);
and U35098 (N_35098,N_34295,N_34548);
or U35099 (N_35099,N_34121,N_34436);
and U35100 (N_35100,N_34317,N_34487);
nor U35101 (N_35101,N_34438,N_34661);
and U35102 (N_35102,N_34964,N_34261);
nor U35103 (N_35103,N_34729,N_34529);
and U35104 (N_35104,N_34237,N_34599);
or U35105 (N_35105,N_34823,N_34008);
xnor U35106 (N_35106,N_34511,N_34326);
and U35107 (N_35107,N_34544,N_34345);
nand U35108 (N_35108,N_34218,N_34984);
xor U35109 (N_35109,N_34560,N_34230);
xnor U35110 (N_35110,N_34858,N_34593);
and U35111 (N_35111,N_34210,N_34990);
xor U35112 (N_35112,N_34996,N_34147);
and U35113 (N_35113,N_34582,N_34126);
or U35114 (N_35114,N_34136,N_34686);
and U35115 (N_35115,N_34606,N_34392);
nor U35116 (N_35116,N_34900,N_34227);
or U35117 (N_35117,N_34190,N_34878);
and U35118 (N_35118,N_34848,N_34551);
nand U35119 (N_35119,N_34509,N_34170);
xnor U35120 (N_35120,N_34607,N_34633);
nor U35121 (N_35121,N_34446,N_34804);
nand U35122 (N_35122,N_34835,N_34602);
and U35123 (N_35123,N_34012,N_34125);
or U35124 (N_35124,N_34703,N_34292);
xnor U35125 (N_35125,N_34182,N_34139);
and U35126 (N_35126,N_34152,N_34853);
and U35127 (N_35127,N_34164,N_34186);
xnor U35128 (N_35128,N_34857,N_34727);
or U35129 (N_35129,N_34004,N_34954);
and U35130 (N_35130,N_34921,N_34448);
xnor U35131 (N_35131,N_34761,N_34750);
and U35132 (N_35132,N_34958,N_34923);
xor U35133 (N_35133,N_34452,N_34798);
nand U35134 (N_35134,N_34180,N_34764);
or U35135 (N_35135,N_34719,N_34907);
xor U35136 (N_35136,N_34735,N_34516);
xnor U35137 (N_35137,N_34341,N_34997);
xnor U35138 (N_35138,N_34553,N_34007);
xnor U35139 (N_35139,N_34662,N_34941);
or U35140 (N_35140,N_34343,N_34050);
xor U35141 (N_35141,N_34654,N_34328);
xor U35142 (N_35142,N_34948,N_34819);
nand U35143 (N_35143,N_34867,N_34070);
nand U35144 (N_35144,N_34483,N_34107);
and U35145 (N_35145,N_34700,N_34395);
or U35146 (N_35146,N_34215,N_34298);
nor U35147 (N_35147,N_34161,N_34831);
or U35148 (N_35148,N_34518,N_34581);
or U35149 (N_35149,N_34836,N_34898);
nand U35150 (N_35150,N_34406,N_34281);
nand U35151 (N_35151,N_34883,N_34957);
xnor U35152 (N_35152,N_34115,N_34415);
nor U35153 (N_35153,N_34203,N_34953);
xor U35154 (N_35154,N_34922,N_34398);
or U35155 (N_35155,N_34927,N_34229);
nand U35156 (N_35156,N_34433,N_34977);
xor U35157 (N_35157,N_34788,N_34198);
nand U35158 (N_35158,N_34011,N_34616);
and U35159 (N_35159,N_34821,N_34931);
nor U35160 (N_35160,N_34981,N_34763);
and U35161 (N_35161,N_34559,N_34776);
or U35162 (N_35162,N_34162,N_34758);
nor U35163 (N_35163,N_34240,N_34584);
nand U35164 (N_35164,N_34006,N_34704);
or U35165 (N_35165,N_34130,N_34680);
nor U35166 (N_35166,N_34993,N_34543);
or U35167 (N_35167,N_34630,N_34847);
nor U35168 (N_35168,N_34956,N_34429);
or U35169 (N_35169,N_34339,N_34065);
nand U35170 (N_35170,N_34033,N_34109);
nor U35171 (N_35171,N_34040,N_34588);
or U35172 (N_35172,N_34146,N_34432);
or U35173 (N_35173,N_34540,N_34409);
and U35174 (N_35174,N_34222,N_34316);
nand U35175 (N_35175,N_34672,N_34120);
nand U35176 (N_35176,N_34453,N_34401);
or U35177 (N_35177,N_34894,N_34019);
xnor U35178 (N_35178,N_34731,N_34257);
nor U35179 (N_35179,N_34787,N_34199);
nor U35180 (N_35180,N_34864,N_34490);
nand U35181 (N_35181,N_34090,N_34383);
xor U35182 (N_35182,N_34250,N_34698);
and U35183 (N_35183,N_34590,N_34786);
or U35184 (N_35184,N_34705,N_34679);
and U35185 (N_35185,N_34191,N_34387);
nand U35186 (N_35186,N_34086,N_34873);
and U35187 (N_35187,N_34457,N_34657);
nand U35188 (N_35188,N_34906,N_34507);
or U35189 (N_35189,N_34080,N_34445);
nor U35190 (N_35190,N_34270,N_34057);
nor U35191 (N_35191,N_34555,N_34514);
or U35192 (N_35192,N_34781,N_34394);
or U35193 (N_35193,N_34982,N_34755);
nand U35194 (N_35194,N_34408,N_34084);
and U35195 (N_35195,N_34363,N_34364);
and U35196 (N_35196,N_34187,N_34715);
or U35197 (N_35197,N_34112,N_34466);
nor U35198 (N_35198,N_34866,N_34739);
xnor U35199 (N_35199,N_34877,N_34967);
or U35200 (N_35200,N_34189,N_34784);
xnor U35201 (N_35201,N_34520,N_34567);
xnor U35202 (N_35202,N_34970,N_34213);
nor U35203 (N_35203,N_34082,N_34598);
xor U35204 (N_35204,N_34009,N_34793);
xnor U35205 (N_35205,N_34462,N_34172);
and U35206 (N_35206,N_34351,N_34732);
or U35207 (N_35207,N_34841,N_34375);
or U35208 (N_35208,N_34983,N_34138);
nand U35209 (N_35209,N_34443,N_34508);
and U35210 (N_35210,N_34613,N_34650);
or U35211 (N_35211,N_34876,N_34512);
nor U35212 (N_35212,N_34223,N_34925);
or U35213 (N_35213,N_34175,N_34471);
xnor U35214 (N_35214,N_34891,N_34871);
and U35215 (N_35215,N_34352,N_34074);
and U35216 (N_35216,N_34513,N_34427);
nand U35217 (N_35217,N_34024,N_34472);
nand U35218 (N_35218,N_34748,N_34826);
nor U35219 (N_35219,N_34938,N_34528);
nand U35220 (N_35220,N_34221,N_34617);
and U35221 (N_35221,N_34539,N_34357);
nand U35222 (N_35222,N_34206,N_34493);
xor U35223 (N_35223,N_34965,N_34459);
and U35224 (N_35224,N_34469,N_34235);
and U35225 (N_35225,N_34488,N_34188);
xor U35226 (N_35226,N_34987,N_34212);
nor U35227 (N_35227,N_34248,N_34167);
xnor U35228 (N_35228,N_34173,N_34418);
nand U35229 (N_35229,N_34228,N_34638);
and U35230 (N_35230,N_34367,N_34562);
xnor U35231 (N_35231,N_34461,N_34865);
nand U35232 (N_35232,N_34153,N_34694);
xnor U35233 (N_35233,N_34986,N_34629);
and U35234 (N_35234,N_34391,N_34422);
nor U35235 (N_35235,N_34905,N_34424);
and U35236 (N_35236,N_34738,N_34664);
nor U35237 (N_35237,N_34101,N_34491);
or U35238 (N_35238,N_34952,N_34051);
nor U35239 (N_35239,N_34752,N_34526);
and U35240 (N_35240,N_34184,N_34919);
xnor U35241 (N_35241,N_34464,N_34881);
nor U35242 (N_35242,N_34577,N_34578);
xnor U35243 (N_35243,N_34381,N_34868);
nor U35244 (N_35244,N_34064,N_34709);
and U35245 (N_35245,N_34226,N_34753);
nand U35246 (N_35246,N_34108,N_34099);
nor U35247 (N_35247,N_34712,N_34313);
nand U35248 (N_35248,N_34169,N_34320);
or U35249 (N_35249,N_34144,N_34193);
nand U35250 (N_35250,N_34097,N_34505);
or U35251 (N_35251,N_34133,N_34202);
nand U35252 (N_35252,N_34160,N_34495);
or U35253 (N_35253,N_34574,N_34856);
nor U35254 (N_35254,N_34839,N_34369);
and U35255 (N_35255,N_34999,N_34413);
and U35256 (N_35256,N_34348,N_34696);
and U35257 (N_35257,N_34201,N_34832);
and U35258 (N_35258,N_34500,N_34455);
nand U35259 (N_35259,N_34859,N_34141);
nand U35260 (N_35260,N_34412,N_34936);
xor U35261 (N_35261,N_34384,N_34792);
or U35262 (N_35262,N_34817,N_34365);
xor U35263 (N_35263,N_34159,N_34123);
and U35264 (N_35264,N_34502,N_34377);
or U35265 (N_35265,N_34482,N_34874);
nand U35266 (N_35266,N_34960,N_34335);
or U35267 (N_35267,N_34820,N_34480);
nor U35268 (N_35268,N_34615,N_34734);
nand U35269 (N_35269,N_34194,N_34855);
nor U35270 (N_35270,N_34410,N_34746);
xnor U35271 (N_35271,N_34885,N_34271);
xnor U35272 (N_35272,N_34176,N_34718);
nor U35273 (N_35273,N_34178,N_34378);
nor U35274 (N_35274,N_34665,N_34149);
and U35275 (N_35275,N_34812,N_34803);
and U35276 (N_35276,N_34417,N_34232);
and U35277 (N_35277,N_34002,N_34723);
xor U35278 (N_35278,N_34047,N_34971);
and U35279 (N_35279,N_34419,N_34396);
or U35280 (N_35280,N_34085,N_34347);
nor U35281 (N_35281,N_34275,N_34503);
or U35282 (N_35282,N_34073,N_34056);
xor U35283 (N_35283,N_34268,N_34995);
nand U35284 (N_35284,N_34850,N_34023);
and U35285 (N_35285,N_34451,N_34498);
nor U35286 (N_35286,N_34113,N_34116);
or U35287 (N_35287,N_34854,N_34430);
nand U35288 (N_35288,N_34280,N_34849);
or U35289 (N_35289,N_34465,N_34949);
nand U35290 (N_35290,N_34586,N_34742);
nor U35291 (N_35291,N_34288,N_34810);
or U35292 (N_35292,N_34045,N_34875);
xor U35293 (N_35293,N_34247,N_34637);
nor U35294 (N_35294,N_34241,N_34346);
xnor U35295 (N_35295,N_34279,N_34148);
nor U35296 (N_35296,N_34737,N_34833);
nand U35297 (N_35297,N_34533,N_34069);
nand U35298 (N_35298,N_34360,N_34404);
xnor U35299 (N_35299,N_34745,N_34627);
xor U35300 (N_35300,N_34421,N_34926);
and U35301 (N_35301,N_34930,N_34059);
xnor U35302 (N_35302,N_34265,N_34767);
and U35303 (N_35303,N_34959,N_34751);
nor U35304 (N_35304,N_34063,N_34407);
nand U35305 (N_35305,N_34802,N_34651);
nor U35306 (N_35306,N_34805,N_34988);
and U35307 (N_35307,N_34411,N_34711);
nand U35308 (N_35308,N_34568,N_34368);
and U35309 (N_35309,N_34646,N_34861);
or U35310 (N_35310,N_34425,N_34174);
xnor U35311 (N_35311,N_34882,N_34549);
nand U35312 (N_35312,N_34103,N_34158);
or U35313 (N_35313,N_34478,N_34552);
nor U35314 (N_35314,N_34370,N_34837);
nand U35315 (N_35315,N_34022,N_34209);
or U35316 (N_35316,N_34840,N_34944);
or U35317 (N_35317,N_34799,N_34231);
or U35318 (N_35318,N_34972,N_34358);
xor U35319 (N_35319,N_34852,N_34458);
xor U35320 (N_35320,N_34249,N_34830);
nand U35321 (N_35321,N_34131,N_34196);
and U35322 (N_35322,N_34736,N_34945);
or U35323 (N_35323,N_34321,N_34256);
nor U35324 (N_35324,N_34460,N_34760);
nor U35325 (N_35325,N_34397,N_34104);
nand U35326 (N_35326,N_34713,N_34238);
and U35327 (N_35327,N_34851,N_34844);
or U35328 (N_35328,N_34806,N_34264);
or U35329 (N_35329,N_34968,N_34475);
and U35330 (N_35330,N_34869,N_34681);
nor U35331 (N_35331,N_34355,N_34937);
nor U35332 (N_35332,N_34311,N_34388);
or U35333 (N_35333,N_34901,N_34550);
xnor U35334 (N_35334,N_34260,N_34110);
xor U35335 (N_35335,N_34122,N_34239);
nand U35336 (N_35336,N_34310,N_34128);
and U35337 (N_35337,N_34325,N_34612);
xor U35338 (N_35338,N_34880,N_34499);
nand U35339 (N_35339,N_34794,N_34504);
nand U35340 (N_35340,N_34088,N_34217);
and U35341 (N_35341,N_34888,N_34038);
xor U35342 (N_35342,N_34818,N_34728);
and U35343 (N_35343,N_34710,N_34373);
and U35344 (N_35344,N_34724,N_34037);
or U35345 (N_35345,N_34450,N_34576);
nand U35346 (N_35346,N_34797,N_34842);
nor U35347 (N_35347,N_34583,N_34749);
and U35348 (N_35348,N_34376,N_34337);
or U35349 (N_35349,N_34714,N_34666);
or U35350 (N_35350,N_34677,N_34296);
nand U35351 (N_35351,N_34531,N_34334);
nand U35352 (N_35352,N_34447,N_34253);
or U35353 (N_35353,N_34282,N_34089);
or U35354 (N_35354,N_34301,N_34535);
and U35355 (N_35355,N_34067,N_34670);
or U35356 (N_35356,N_34278,N_34682);
nand U35357 (N_35357,N_34010,N_34909);
nor U35358 (N_35358,N_34323,N_34005);
nor U35359 (N_35359,N_34790,N_34591);
and U35360 (N_35360,N_34163,N_34653);
or U35361 (N_35361,N_34989,N_34078);
xor U35362 (N_35362,N_34494,N_34151);
and U35363 (N_35363,N_34001,N_34655);
xor U35364 (N_35364,N_34770,N_34340);
or U35365 (N_35365,N_34124,N_34807);
and U35366 (N_35366,N_34389,N_34145);
and U35367 (N_35367,N_34716,N_34978);
xnor U35368 (N_35368,N_34062,N_34585);
and U35369 (N_35369,N_34642,N_34071);
or U35370 (N_35370,N_34697,N_34611);
or U35371 (N_35371,N_34306,N_34592);
xnor U35372 (N_35372,N_34034,N_34933);
and U35373 (N_35373,N_34517,N_34829);
or U35374 (N_35374,N_34610,N_34294);
or U35375 (N_35375,N_34402,N_34026);
or U35376 (N_35376,N_34827,N_34556);
nor U35377 (N_35377,N_34485,N_34025);
and U35378 (N_35378,N_34233,N_34297);
and U35379 (N_35379,N_34648,N_34385);
nand U35380 (N_35380,N_34449,N_34920);
xnor U35381 (N_35381,N_34087,N_34525);
nor U35382 (N_35382,N_34683,N_34795);
xor U35383 (N_35383,N_34331,N_34208);
or U35384 (N_35384,N_34963,N_34740);
nor U35385 (N_35385,N_34730,N_34129);
xor U35386 (N_35386,N_34649,N_34809);
xor U35387 (N_35387,N_34060,N_34815);
nor U35388 (N_35388,N_34860,N_34470);
and U35389 (N_35389,N_34091,N_34390);
and U35390 (N_35390,N_34608,N_34372);
and U35391 (N_35391,N_34899,N_34545);
or U35392 (N_35392,N_34783,N_34722);
nand U35393 (N_35393,N_34486,N_34510);
xor U35394 (N_35394,N_34929,N_34635);
nor U35395 (N_35395,N_34537,N_34699);
and U35396 (N_35396,N_34708,N_34913);
nand U35397 (N_35397,N_34489,N_34154);
xor U35398 (N_35398,N_34031,N_34435);
nor U35399 (N_35399,N_34371,N_34224);
and U35400 (N_35400,N_34476,N_34733);
nand U35401 (N_35401,N_34800,N_34572);
or U35402 (N_35402,N_34547,N_34300);
or U35403 (N_35403,N_34893,N_34028);
nor U35404 (N_35404,N_34589,N_34344);
nand U35405 (N_35405,N_34192,N_34824);
nor U35406 (N_35406,N_34142,N_34254);
xnor U35407 (N_35407,N_34691,N_34353);
nor U35408 (N_35408,N_34048,N_34530);
xnor U35409 (N_35409,N_34137,N_34811);
nor U35410 (N_35410,N_34197,N_34695);
or U35411 (N_35411,N_34935,N_34561);
nor U35412 (N_35412,N_34717,N_34274);
xor U35413 (N_35413,N_34442,N_34171);
nand U35414 (N_35414,N_34243,N_34437);
or U35415 (N_35415,N_34565,N_34757);
and U35416 (N_35416,N_34285,N_34319);
nor U35417 (N_35417,N_34908,N_34204);
or U35418 (N_35418,N_34671,N_34501);
nand U35419 (N_35419,N_34216,N_34702);
nor U35420 (N_35420,N_34423,N_34887);
xor U35421 (N_35421,N_34557,N_34366);
nand U35422 (N_35422,N_34289,N_34399);
or U35423 (N_35423,N_34554,N_34636);
or U35424 (N_35424,N_34307,N_34668);
nor U35425 (N_35425,N_34768,N_34594);
and U35426 (N_35426,N_34150,N_34332);
nand U35427 (N_35427,N_34773,N_34886);
or U35428 (N_35428,N_34166,N_34205);
or U35429 (N_35429,N_34947,N_34324);
and U35430 (N_35430,N_34342,N_34273);
xor U35431 (N_35431,N_34701,N_34796);
or U35432 (N_35432,N_34687,N_34569);
and U35433 (N_35433,N_34046,N_34515);
nor U35434 (N_35434,N_34039,N_34903);
nand U35435 (N_35435,N_34962,N_34884);
xnor U35436 (N_35436,N_34915,N_34747);
or U35437 (N_35437,N_34946,N_34674);
nand U35438 (N_35438,N_34772,N_34350);
or U35439 (N_35439,N_34308,N_34015);
or U35440 (N_35440,N_34774,N_34030);
and U35441 (N_35441,N_34092,N_34838);
or U35442 (N_35442,N_34910,N_34892);
xor U35443 (N_35443,N_34127,N_34973);
nand U35444 (N_35444,N_34546,N_34041);
or U35445 (N_35445,N_34386,N_34902);
or U35446 (N_35446,N_34207,N_34658);
or U35447 (N_35447,N_34467,N_34016);
or U35448 (N_35448,N_34522,N_34536);
nand U35449 (N_35449,N_34625,N_34976);
or U35450 (N_35450,N_34521,N_34917);
xor U35451 (N_35451,N_34379,N_34293);
nor U35452 (N_35452,N_34862,N_34081);
nor U35453 (N_35453,N_34225,N_34620);
nor U35454 (N_35454,N_34614,N_34076);
xor U35455 (N_35455,N_34036,N_34870);
or U35456 (N_35456,N_34309,N_34304);
nor U35457 (N_35457,N_34165,N_34808);
or U35458 (N_35458,N_34943,N_34055);
nor U35459 (N_35459,N_34754,N_34095);
nand U35460 (N_35460,N_34791,N_34020);
xnor U35461 (N_35461,N_34564,N_34896);
xnor U35462 (N_35462,N_34916,N_34068);
xor U35463 (N_35463,N_34272,N_34924);
xor U35464 (N_35464,N_34318,N_34780);
or U35465 (N_35465,N_34601,N_34479);
and U35466 (N_35466,N_34688,N_34027);
nand U35467 (N_35467,N_34359,N_34042);
and U35468 (N_35468,N_34789,N_34631);
nand U35469 (N_35469,N_34542,N_34029);
or U35470 (N_35470,N_34720,N_34647);
nor U35471 (N_35471,N_34690,N_34632);
xnor U35472 (N_35472,N_34405,N_34286);
or U35473 (N_35473,N_34741,N_34966);
nand U35474 (N_35474,N_34252,N_34118);
or U35475 (N_35475,N_34975,N_34726);
nor U35476 (N_35476,N_34497,N_34816);
nand U35477 (N_35477,N_34054,N_34333);
and U35478 (N_35478,N_34527,N_34481);
nand U35479 (N_35479,N_34889,N_34603);
xnor U35480 (N_35480,N_34969,N_34093);
nor U35481 (N_35481,N_34361,N_34134);
nand U35482 (N_35482,N_34299,N_34195);
and U35483 (N_35483,N_34096,N_34267);
xor U35484 (N_35484,N_34214,N_34259);
nor U35485 (N_35485,N_34236,N_34263);
nor U35486 (N_35486,N_34075,N_34663);
or U35487 (N_35487,N_34939,N_34640);
nand U35488 (N_35488,N_34775,N_34912);
xnor U35489 (N_35489,N_34825,N_34302);
and U35490 (N_35490,N_34928,N_34782);
and U35491 (N_35491,N_34634,N_34777);
xor U35492 (N_35492,N_34269,N_34393);
nand U35493 (N_35493,N_34692,N_34645);
and U35494 (N_35494,N_34596,N_34676);
and U35495 (N_35495,N_34914,N_34918);
nor U35496 (N_35496,N_34571,N_34117);
or U35497 (N_35497,N_34845,N_34765);
nor U35498 (N_35498,N_34403,N_34619);
and U35499 (N_35499,N_34354,N_34519);
and U35500 (N_35500,N_34132,N_34331);
and U35501 (N_35501,N_34033,N_34376);
and U35502 (N_35502,N_34506,N_34267);
xnor U35503 (N_35503,N_34168,N_34948);
or U35504 (N_35504,N_34898,N_34715);
and U35505 (N_35505,N_34818,N_34299);
nand U35506 (N_35506,N_34894,N_34679);
or U35507 (N_35507,N_34283,N_34718);
xor U35508 (N_35508,N_34768,N_34506);
nor U35509 (N_35509,N_34889,N_34869);
nor U35510 (N_35510,N_34972,N_34201);
and U35511 (N_35511,N_34376,N_34240);
xor U35512 (N_35512,N_34728,N_34088);
xor U35513 (N_35513,N_34650,N_34004);
nand U35514 (N_35514,N_34878,N_34265);
nor U35515 (N_35515,N_34807,N_34447);
or U35516 (N_35516,N_34992,N_34282);
nor U35517 (N_35517,N_34156,N_34639);
nand U35518 (N_35518,N_34438,N_34601);
and U35519 (N_35519,N_34753,N_34100);
and U35520 (N_35520,N_34826,N_34308);
and U35521 (N_35521,N_34220,N_34208);
xor U35522 (N_35522,N_34908,N_34093);
nand U35523 (N_35523,N_34981,N_34515);
and U35524 (N_35524,N_34605,N_34027);
and U35525 (N_35525,N_34002,N_34100);
and U35526 (N_35526,N_34139,N_34317);
and U35527 (N_35527,N_34767,N_34948);
and U35528 (N_35528,N_34748,N_34078);
and U35529 (N_35529,N_34378,N_34358);
xnor U35530 (N_35530,N_34823,N_34929);
or U35531 (N_35531,N_34665,N_34921);
and U35532 (N_35532,N_34868,N_34321);
and U35533 (N_35533,N_34131,N_34736);
and U35534 (N_35534,N_34300,N_34638);
or U35535 (N_35535,N_34327,N_34370);
xnor U35536 (N_35536,N_34874,N_34630);
or U35537 (N_35537,N_34225,N_34887);
nor U35538 (N_35538,N_34070,N_34956);
nand U35539 (N_35539,N_34028,N_34859);
nor U35540 (N_35540,N_34886,N_34751);
nor U35541 (N_35541,N_34765,N_34668);
nor U35542 (N_35542,N_34024,N_34997);
nor U35543 (N_35543,N_34297,N_34173);
nand U35544 (N_35544,N_34269,N_34348);
or U35545 (N_35545,N_34742,N_34556);
nand U35546 (N_35546,N_34788,N_34327);
nor U35547 (N_35547,N_34982,N_34275);
xor U35548 (N_35548,N_34674,N_34555);
or U35549 (N_35549,N_34209,N_34219);
or U35550 (N_35550,N_34235,N_34835);
nor U35551 (N_35551,N_34174,N_34841);
and U35552 (N_35552,N_34628,N_34666);
and U35553 (N_35553,N_34280,N_34916);
and U35554 (N_35554,N_34675,N_34293);
and U35555 (N_35555,N_34889,N_34453);
xnor U35556 (N_35556,N_34942,N_34544);
xor U35557 (N_35557,N_34080,N_34665);
nand U35558 (N_35558,N_34291,N_34000);
nand U35559 (N_35559,N_34901,N_34696);
and U35560 (N_35560,N_34184,N_34897);
xnor U35561 (N_35561,N_34811,N_34319);
and U35562 (N_35562,N_34833,N_34624);
nand U35563 (N_35563,N_34859,N_34046);
or U35564 (N_35564,N_34535,N_34580);
nand U35565 (N_35565,N_34930,N_34239);
and U35566 (N_35566,N_34923,N_34075);
nand U35567 (N_35567,N_34351,N_34157);
xnor U35568 (N_35568,N_34558,N_34101);
nand U35569 (N_35569,N_34144,N_34476);
and U35570 (N_35570,N_34799,N_34528);
and U35571 (N_35571,N_34510,N_34780);
and U35572 (N_35572,N_34091,N_34016);
nand U35573 (N_35573,N_34782,N_34767);
xor U35574 (N_35574,N_34487,N_34986);
xor U35575 (N_35575,N_34624,N_34487);
and U35576 (N_35576,N_34102,N_34010);
xnor U35577 (N_35577,N_34792,N_34582);
nand U35578 (N_35578,N_34038,N_34348);
nor U35579 (N_35579,N_34412,N_34470);
xnor U35580 (N_35580,N_34920,N_34608);
or U35581 (N_35581,N_34547,N_34454);
or U35582 (N_35582,N_34015,N_34209);
and U35583 (N_35583,N_34418,N_34986);
nor U35584 (N_35584,N_34723,N_34090);
nand U35585 (N_35585,N_34075,N_34464);
nor U35586 (N_35586,N_34232,N_34152);
nor U35587 (N_35587,N_34708,N_34982);
or U35588 (N_35588,N_34947,N_34945);
nand U35589 (N_35589,N_34061,N_34016);
nor U35590 (N_35590,N_34532,N_34309);
xor U35591 (N_35591,N_34425,N_34251);
nand U35592 (N_35592,N_34273,N_34762);
nor U35593 (N_35593,N_34743,N_34768);
xor U35594 (N_35594,N_34801,N_34392);
or U35595 (N_35595,N_34904,N_34105);
and U35596 (N_35596,N_34261,N_34905);
xor U35597 (N_35597,N_34529,N_34220);
or U35598 (N_35598,N_34582,N_34046);
nand U35599 (N_35599,N_34184,N_34304);
nor U35600 (N_35600,N_34720,N_34033);
or U35601 (N_35601,N_34003,N_34792);
and U35602 (N_35602,N_34507,N_34014);
nor U35603 (N_35603,N_34230,N_34121);
and U35604 (N_35604,N_34396,N_34977);
nor U35605 (N_35605,N_34326,N_34831);
nor U35606 (N_35606,N_34996,N_34365);
xor U35607 (N_35607,N_34355,N_34643);
xnor U35608 (N_35608,N_34701,N_34436);
and U35609 (N_35609,N_34246,N_34488);
nand U35610 (N_35610,N_34455,N_34689);
nand U35611 (N_35611,N_34608,N_34147);
nor U35612 (N_35612,N_34073,N_34458);
xnor U35613 (N_35613,N_34619,N_34050);
xor U35614 (N_35614,N_34861,N_34737);
nand U35615 (N_35615,N_34537,N_34226);
nor U35616 (N_35616,N_34603,N_34472);
xnor U35617 (N_35617,N_34446,N_34117);
or U35618 (N_35618,N_34447,N_34259);
xor U35619 (N_35619,N_34680,N_34121);
nand U35620 (N_35620,N_34738,N_34253);
nand U35621 (N_35621,N_34910,N_34783);
and U35622 (N_35622,N_34530,N_34527);
or U35623 (N_35623,N_34468,N_34586);
or U35624 (N_35624,N_34130,N_34580);
or U35625 (N_35625,N_34883,N_34813);
and U35626 (N_35626,N_34702,N_34864);
or U35627 (N_35627,N_34315,N_34549);
xor U35628 (N_35628,N_34564,N_34330);
nand U35629 (N_35629,N_34412,N_34853);
nand U35630 (N_35630,N_34750,N_34279);
xnor U35631 (N_35631,N_34451,N_34874);
nand U35632 (N_35632,N_34166,N_34436);
nor U35633 (N_35633,N_34093,N_34471);
nor U35634 (N_35634,N_34474,N_34173);
nand U35635 (N_35635,N_34960,N_34962);
xor U35636 (N_35636,N_34963,N_34075);
nor U35637 (N_35637,N_34796,N_34438);
or U35638 (N_35638,N_34157,N_34668);
or U35639 (N_35639,N_34858,N_34417);
or U35640 (N_35640,N_34384,N_34480);
or U35641 (N_35641,N_34189,N_34328);
nand U35642 (N_35642,N_34040,N_34598);
nor U35643 (N_35643,N_34011,N_34735);
or U35644 (N_35644,N_34938,N_34470);
and U35645 (N_35645,N_34583,N_34746);
and U35646 (N_35646,N_34877,N_34217);
xnor U35647 (N_35647,N_34056,N_34664);
xnor U35648 (N_35648,N_34055,N_34733);
nor U35649 (N_35649,N_34500,N_34383);
nand U35650 (N_35650,N_34073,N_34961);
xnor U35651 (N_35651,N_34133,N_34517);
nand U35652 (N_35652,N_34566,N_34395);
or U35653 (N_35653,N_34534,N_34536);
nand U35654 (N_35654,N_34475,N_34413);
or U35655 (N_35655,N_34612,N_34373);
or U35656 (N_35656,N_34503,N_34862);
and U35657 (N_35657,N_34136,N_34881);
nor U35658 (N_35658,N_34394,N_34277);
and U35659 (N_35659,N_34322,N_34850);
nand U35660 (N_35660,N_34273,N_34098);
and U35661 (N_35661,N_34148,N_34779);
and U35662 (N_35662,N_34427,N_34869);
xnor U35663 (N_35663,N_34947,N_34750);
xnor U35664 (N_35664,N_34118,N_34749);
nand U35665 (N_35665,N_34555,N_34654);
nand U35666 (N_35666,N_34318,N_34252);
nor U35667 (N_35667,N_34116,N_34593);
and U35668 (N_35668,N_34170,N_34672);
nand U35669 (N_35669,N_34034,N_34813);
xnor U35670 (N_35670,N_34691,N_34248);
xor U35671 (N_35671,N_34020,N_34901);
nand U35672 (N_35672,N_34763,N_34780);
nor U35673 (N_35673,N_34376,N_34047);
and U35674 (N_35674,N_34747,N_34813);
or U35675 (N_35675,N_34827,N_34446);
xnor U35676 (N_35676,N_34559,N_34424);
nor U35677 (N_35677,N_34856,N_34050);
nor U35678 (N_35678,N_34100,N_34011);
nor U35679 (N_35679,N_34604,N_34025);
nand U35680 (N_35680,N_34592,N_34421);
xnor U35681 (N_35681,N_34961,N_34082);
nor U35682 (N_35682,N_34613,N_34645);
xnor U35683 (N_35683,N_34484,N_34282);
xor U35684 (N_35684,N_34868,N_34556);
or U35685 (N_35685,N_34917,N_34609);
xor U35686 (N_35686,N_34907,N_34585);
xor U35687 (N_35687,N_34159,N_34788);
nand U35688 (N_35688,N_34585,N_34360);
xnor U35689 (N_35689,N_34024,N_34887);
nor U35690 (N_35690,N_34242,N_34011);
nor U35691 (N_35691,N_34520,N_34817);
or U35692 (N_35692,N_34151,N_34167);
xnor U35693 (N_35693,N_34464,N_34756);
and U35694 (N_35694,N_34964,N_34267);
or U35695 (N_35695,N_34786,N_34264);
nor U35696 (N_35696,N_34732,N_34982);
xnor U35697 (N_35697,N_34363,N_34843);
xnor U35698 (N_35698,N_34586,N_34949);
nor U35699 (N_35699,N_34576,N_34084);
nor U35700 (N_35700,N_34129,N_34652);
nand U35701 (N_35701,N_34251,N_34169);
xnor U35702 (N_35702,N_34152,N_34566);
nand U35703 (N_35703,N_34215,N_34032);
nor U35704 (N_35704,N_34658,N_34857);
nor U35705 (N_35705,N_34381,N_34893);
nor U35706 (N_35706,N_34196,N_34638);
nor U35707 (N_35707,N_34173,N_34743);
or U35708 (N_35708,N_34300,N_34830);
or U35709 (N_35709,N_34863,N_34004);
nand U35710 (N_35710,N_34331,N_34195);
and U35711 (N_35711,N_34329,N_34635);
or U35712 (N_35712,N_34886,N_34526);
and U35713 (N_35713,N_34495,N_34121);
or U35714 (N_35714,N_34167,N_34736);
nand U35715 (N_35715,N_34905,N_34382);
nor U35716 (N_35716,N_34936,N_34560);
nor U35717 (N_35717,N_34397,N_34584);
or U35718 (N_35718,N_34651,N_34921);
and U35719 (N_35719,N_34973,N_34948);
nand U35720 (N_35720,N_34800,N_34406);
and U35721 (N_35721,N_34640,N_34891);
nand U35722 (N_35722,N_34763,N_34793);
nand U35723 (N_35723,N_34760,N_34389);
or U35724 (N_35724,N_34567,N_34989);
or U35725 (N_35725,N_34384,N_34291);
xnor U35726 (N_35726,N_34196,N_34465);
and U35727 (N_35727,N_34610,N_34634);
and U35728 (N_35728,N_34499,N_34961);
nand U35729 (N_35729,N_34238,N_34979);
nand U35730 (N_35730,N_34548,N_34273);
and U35731 (N_35731,N_34952,N_34738);
nor U35732 (N_35732,N_34293,N_34650);
and U35733 (N_35733,N_34376,N_34489);
xor U35734 (N_35734,N_34406,N_34111);
nor U35735 (N_35735,N_34845,N_34508);
xor U35736 (N_35736,N_34260,N_34579);
and U35737 (N_35737,N_34120,N_34030);
nand U35738 (N_35738,N_34067,N_34127);
xnor U35739 (N_35739,N_34888,N_34067);
nand U35740 (N_35740,N_34204,N_34191);
and U35741 (N_35741,N_34199,N_34950);
nor U35742 (N_35742,N_34764,N_34943);
xor U35743 (N_35743,N_34099,N_34395);
nor U35744 (N_35744,N_34387,N_34039);
or U35745 (N_35745,N_34431,N_34403);
or U35746 (N_35746,N_34164,N_34902);
or U35747 (N_35747,N_34423,N_34188);
or U35748 (N_35748,N_34881,N_34828);
and U35749 (N_35749,N_34071,N_34219);
nor U35750 (N_35750,N_34116,N_34059);
nor U35751 (N_35751,N_34590,N_34524);
xnor U35752 (N_35752,N_34629,N_34400);
and U35753 (N_35753,N_34787,N_34586);
or U35754 (N_35754,N_34554,N_34155);
and U35755 (N_35755,N_34722,N_34163);
and U35756 (N_35756,N_34382,N_34043);
nor U35757 (N_35757,N_34277,N_34987);
nor U35758 (N_35758,N_34518,N_34955);
xor U35759 (N_35759,N_34830,N_34906);
xnor U35760 (N_35760,N_34841,N_34098);
nor U35761 (N_35761,N_34162,N_34414);
xor U35762 (N_35762,N_34512,N_34131);
or U35763 (N_35763,N_34985,N_34299);
xor U35764 (N_35764,N_34976,N_34943);
nor U35765 (N_35765,N_34451,N_34844);
nor U35766 (N_35766,N_34057,N_34217);
and U35767 (N_35767,N_34454,N_34081);
or U35768 (N_35768,N_34941,N_34705);
nor U35769 (N_35769,N_34126,N_34159);
nor U35770 (N_35770,N_34073,N_34002);
or U35771 (N_35771,N_34086,N_34123);
nand U35772 (N_35772,N_34645,N_34917);
nor U35773 (N_35773,N_34659,N_34617);
or U35774 (N_35774,N_34343,N_34683);
xor U35775 (N_35775,N_34540,N_34521);
nor U35776 (N_35776,N_34680,N_34588);
nor U35777 (N_35777,N_34071,N_34070);
nand U35778 (N_35778,N_34226,N_34827);
nand U35779 (N_35779,N_34005,N_34472);
or U35780 (N_35780,N_34504,N_34431);
and U35781 (N_35781,N_34152,N_34691);
and U35782 (N_35782,N_34320,N_34292);
nand U35783 (N_35783,N_34242,N_34543);
nand U35784 (N_35784,N_34632,N_34209);
nor U35785 (N_35785,N_34816,N_34118);
and U35786 (N_35786,N_34245,N_34766);
or U35787 (N_35787,N_34851,N_34192);
or U35788 (N_35788,N_34674,N_34692);
xnor U35789 (N_35789,N_34582,N_34930);
or U35790 (N_35790,N_34139,N_34051);
nand U35791 (N_35791,N_34136,N_34657);
nand U35792 (N_35792,N_34421,N_34928);
nand U35793 (N_35793,N_34140,N_34761);
nand U35794 (N_35794,N_34531,N_34030);
and U35795 (N_35795,N_34349,N_34905);
xor U35796 (N_35796,N_34857,N_34580);
and U35797 (N_35797,N_34099,N_34274);
nor U35798 (N_35798,N_34980,N_34328);
and U35799 (N_35799,N_34879,N_34987);
nand U35800 (N_35800,N_34629,N_34064);
nand U35801 (N_35801,N_34833,N_34575);
and U35802 (N_35802,N_34504,N_34341);
nand U35803 (N_35803,N_34052,N_34352);
nor U35804 (N_35804,N_34307,N_34498);
nor U35805 (N_35805,N_34142,N_34455);
and U35806 (N_35806,N_34954,N_34234);
xor U35807 (N_35807,N_34631,N_34063);
nand U35808 (N_35808,N_34760,N_34411);
nor U35809 (N_35809,N_34167,N_34681);
nand U35810 (N_35810,N_34763,N_34551);
xor U35811 (N_35811,N_34531,N_34927);
and U35812 (N_35812,N_34590,N_34037);
nand U35813 (N_35813,N_34577,N_34257);
xor U35814 (N_35814,N_34085,N_34703);
or U35815 (N_35815,N_34494,N_34946);
nor U35816 (N_35816,N_34975,N_34211);
xor U35817 (N_35817,N_34360,N_34918);
nor U35818 (N_35818,N_34971,N_34700);
nand U35819 (N_35819,N_34853,N_34964);
nand U35820 (N_35820,N_34286,N_34371);
nand U35821 (N_35821,N_34518,N_34411);
and U35822 (N_35822,N_34638,N_34854);
nand U35823 (N_35823,N_34741,N_34412);
xnor U35824 (N_35824,N_34183,N_34390);
xor U35825 (N_35825,N_34813,N_34874);
nand U35826 (N_35826,N_34202,N_34694);
or U35827 (N_35827,N_34341,N_34939);
and U35828 (N_35828,N_34518,N_34841);
or U35829 (N_35829,N_34035,N_34625);
nor U35830 (N_35830,N_34828,N_34511);
and U35831 (N_35831,N_34024,N_34386);
nor U35832 (N_35832,N_34675,N_34203);
nor U35833 (N_35833,N_34161,N_34083);
nand U35834 (N_35834,N_34182,N_34644);
xor U35835 (N_35835,N_34686,N_34363);
and U35836 (N_35836,N_34981,N_34219);
or U35837 (N_35837,N_34286,N_34150);
nor U35838 (N_35838,N_34799,N_34174);
and U35839 (N_35839,N_34406,N_34923);
nand U35840 (N_35840,N_34898,N_34609);
and U35841 (N_35841,N_34937,N_34549);
nand U35842 (N_35842,N_34914,N_34141);
or U35843 (N_35843,N_34784,N_34138);
xnor U35844 (N_35844,N_34401,N_34238);
nand U35845 (N_35845,N_34545,N_34257);
and U35846 (N_35846,N_34438,N_34746);
xor U35847 (N_35847,N_34068,N_34803);
and U35848 (N_35848,N_34689,N_34010);
xnor U35849 (N_35849,N_34071,N_34347);
nand U35850 (N_35850,N_34949,N_34955);
nor U35851 (N_35851,N_34660,N_34380);
nor U35852 (N_35852,N_34482,N_34553);
and U35853 (N_35853,N_34620,N_34426);
or U35854 (N_35854,N_34766,N_34374);
xor U35855 (N_35855,N_34454,N_34269);
nand U35856 (N_35856,N_34154,N_34854);
nand U35857 (N_35857,N_34155,N_34506);
nor U35858 (N_35858,N_34805,N_34993);
and U35859 (N_35859,N_34860,N_34106);
nand U35860 (N_35860,N_34011,N_34077);
nor U35861 (N_35861,N_34934,N_34877);
nor U35862 (N_35862,N_34781,N_34742);
and U35863 (N_35863,N_34584,N_34489);
nor U35864 (N_35864,N_34188,N_34688);
nand U35865 (N_35865,N_34954,N_34867);
and U35866 (N_35866,N_34476,N_34041);
nor U35867 (N_35867,N_34840,N_34866);
xor U35868 (N_35868,N_34338,N_34854);
nand U35869 (N_35869,N_34725,N_34201);
or U35870 (N_35870,N_34686,N_34493);
and U35871 (N_35871,N_34114,N_34666);
nand U35872 (N_35872,N_34247,N_34275);
or U35873 (N_35873,N_34525,N_34553);
nand U35874 (N_35874,N_34544,N_34279);
or U35875 (N_35875,N_34795,N_34656);
xor U35876 (N_35876,N_34167,N_34919);
xnor U35877 (N_35877,N_34454,N_34966);
nor U35878 (N_35878,N_34779,N_34060);
nor U35879 (N_35879,N_34659,N_34379);
xor U35880 (N_35880,N_34051,N_34821);
and U35881 (N_35881,N_34190,N_34643);
xor U35882 (N_35882,N_34387,N_34944);
and U35883 (N_35883,N_34293,N_34406);
or U35884 (N_35884,N_34353,N_34196);
nand U35885 (N_35885,N_34157,N_34407);
or U35886 (N_35886,N_34726,N_34024);
xnor U35887 (N_35887,N_34356,N_34424);
nand U35888 (N_35888,N_34780,N_34206);
or U35889 (N_35889,N_34284,N_34366);
or U35890 (N_35890,N_34497,N_34544);
nor U35891 (N_35891,N_34055,N_34014);
and U35892 (N_35892,N_34019,N_34468);
nand U35893 (N_35893,N_34390,N_34382);
or U35894 (N_35894,N_34399,N_34059);
and U35895 (N_35895,N_34353,N_34450);
nor U35896 (N_35896,N_34960,N_34085);
nand U35897 (N_35897,N_34570,N_34872);
nand U35898 (N_35898,N_34926,N_34797);
or U35899 (N_35899,N_34418,N_34839);
xnor U35900 (N_35900,N_34885,N_34807);
or U35901 (N_35901,N_34165,N_34457);
nand U35902 (N_35902,N_34115,N_34001);
nand U35903 (N_35903,N_34640,N_34198);
and U35904 (N_35904,N_34820,N_34935);
or U35905 (N_35905,N_34291,N_34374);
xnor U35906 (N_35906,N_34519,N_34968);
or U35907 (N_35907,N_34602,N_34551);
and U35908 (N_35908,N_34803,N_34082);
and U35909 (N_35909,N_34975,N_34234);
or U35910 (N_35910,N_34079,N_34282);
or U35911 (N_35911,N_34600,N_34370);
xor U35912 (N_35912,N_34376,N_34127);
and U35913 (N_35913,N_34430,N_34147);
xor U35914 (N_35914,N_34907,N_34203);
or U35915 (N_35915,N_34268,N_34828);
or U35916 (N_35916,N_34413,N_34790);
nand U35917 (N_35917,N_34002,N_34409);
and U35918 (N_35918,N_34190,N_34143);
nand U35919 (N_35919,N_34376,N_34276);
or U35920 (N_35920,N_34325,N_34167);
and U35921 (N_35921,N_34342,N_34584);
nor U35922 (N_35922,N_34047,N_34155);
nor U35923 (N_35923,N_34249,N_34111);
xor U35924 (N_35924,N_34612,N_34994);
or U35925 (N_35925,N_34324,N_34930);
nand U35926 (N_35926,N_34386,N_34353);
nor U35927 (N_35927,N_34473,N_34651);
or U35928 (N_35928,N_34808,N_34838);
nor U35929 (N_35929,N_34866,N_34912);
nand U35930 (N_35930,N_34069,N_34469);
nor U35931 (N_35931,N_34641,N_34083);
and U35932 (N_35932,N_34023,N_34773);
and U35933 (N_35933,N_34700,N_34605);
xor U35934 (N_35934,N_34475,N_34046);
xor U35935 (N_35935,N_34606,N_34284);
or U35936 (N_35936,N_34570,N_34189);
nand U35937 (N_35937,N_34194,N_34630);
xnor U35938 (N_35938,N_34357,N_34371);
nand U35939 (N_35939,N_34160,N_34399);
or U35940 (N_35940,N_34136,N_34230);
and U35941 (N_35941,N_34268,N_34374);
nor U35942 (N_35942,N_34602,N_34877);
and U35943 (N_35943,N_34630,N_34279);
or U35944 (N_35944,N_34952,N_34150);
nand U35945 (N_35945,N_34563,N_34707);
or U35946 (N_35946,N_34221,N_34940);
nand U35947 (N_35947,N_34436,N_34047);
xor U35948 (N_35948,N_34444,N_34242);
or U35949 (N_35949,N_34273,N_34256);
xor U35950 (N_35950,N_34123,N_34728);
nor U35951 (N_35951,N_34910,N_34520);
or U35952 (N_35952,N_34775,N_34210);
nor U35953 (N_35953,N_34085,N_34002);
xor U35954 (N_35954,N_34317,N_34730);
xnor U35955 (N_35955,N_34282,N_34279);
nor U35956 (N_35956,N_34021,N_34458);
nand U35957 (N_35957,N_34094,N_34387);
xor U35958 (N_35958,N_34999,N_34564);
nor U35959 (N_35959,N_34342,N_34005);
nand U35960 (N_35960,N_34348,N_34116);
or U35961 (N_35961,N_34095,N_34692);
and U35962 (N_35962,N_34366,N_34135);
nand U35963 (N_35963,N_34596,N_34666);
xnor U35964 (N_35964,N_34524,N_34281);
or U35965 (N_35965,N_34368,N_34093);
and U35966 (N_35966,N_34309,N_34841);
nand U35967 (N_35967,N_34802,N_34128);
and U35968 (N_35968,N_34495,N_34368);
xor U35969 (N_35969,N_34533,N_34826);
nor U35970 (N_35970,N_34555,N_34739);
and U35971 (N_35971,N_34553,N_34297);
or U35972 (N_35972,N_34511,N_34705);
and U35973 (N_35973,N_34372,N_34158);
and U35974 (N_35974,N_34958,N_34374);
xor U35975 (N_35975,N_34751,N_34294);
and U35976 (N_35976,N_34659,N_34518);
and U35977 (N_35977,N_34888,N_34008);
nor U35978 (N_35978,N_34509,N_34274);
or U35979 (N_35979,N_34031,N_34249);
and U35980 (N_35980,N_34242,N_34835);
or U35981 (N_35981,N_34532,N_34716);
xnor U35982 (N_35982,N_34040,N_34814);
or U35983 (N_35983,N_34373,N_34119);
nand U35984 (N_35984,N_34424,N_34283);
and U35985 (N_35985,N_34464,N_34207);
xnor U35986 (N_35986,N_34508,N_34096);
or U35987 (N_35987,N_34958,N_34467);
nand U35988 (N_35988,N_34360,N_34103);
nand U35989 (N_35989,N_34458,N_34829);
and U35990 (N_35990,N_34143,N_34105);
and U35991 (N_35991,N_34724,N_34706);
and U35992 (N_35992,N_34526,N_34001);
nor U35993 (N_35993,N_34123,N_34251);
or U35994 (N_35994,N_34475,N_34664);
xor U35995 (N_35995,N_34177,N_34122);
nor U35996 (N_35996,N_34818,N_34273);
nor U35997 (N_35997,N_34133,N_34554);
or U35998 (N_35998,N_34281,N_34963);
nand U35999 (N_35999,N_34813,N_34997);
or U36000 (N_36000,N_35453,N_35790);
nor U36001 (N_36001,N_35205,N_35565);
nand U36002 (N_36002,N_35293,N_35979);
and U36003 (N_36003,N_35520,N_35639);
nor U36004 (N_36004,N_35577,N_35172);
and U36005 (N_36005,N_35466,N_35393);
nand U36006 (N_36006,N_35660,N_35890);
and U36007 (N_36007,N_35865,N_35170);
nand U36008 (N_36008,N_35544,N_35057);
nand U36009 (N_36009,N_35391,N_35826);
xnor U36010 (N_36010,N_35332,N_35338);
and U36011 (N_36011,N_35078,N_35808);
nand U36012 (N_36012,N_35440,N_35506);
nor U36013 (N_36013,N_35583,N_35745);
or U36014 (N_36014,N_35499,N_35355);
xor U36015 (N_36015,N_35299,N_35538);
xnor U36016 (N_36016,N_35292,N_35256);
or U36017 (N_36017,N_35262,N_35014);
nor U36018 (N_36018,N_35597,N_35714);
nor U36019 (N_36019,N_35581,N_35604);
nor U36020 (N_36020,N_35917,N_35168);
nor U36021 (N_36021,N_35752,N_35582);
xor U36022 (N_36022,N_35388,N_35495);
xor U36023 (N_36023,N_35615,N_35980);
or U36024 (N_36024,N_35514,N_35301);
or U36025 (N_36025,N_35215,N_35197);
nor U36026 (N_36026,N_35284,N_35525);
or U36027 (N_36027,N_35989,N_35611);
nand U36028 (N_36028,N_35427,N_35656);
nand U36029 (N_36029,N_35992,N_35113);
or U36030 (N_36030,N_35234,N_35037);
nand U36031 (N_36031,N_35713,N_35836);
nor U36032 (N_36032,N_35122,N_35066);
nand U36033 (N_36033,N_35661,N_35801);
nand U36034 (N_36034,N_35648,N_35456);
and U36035 (N_36035,N_35005,N_35006);
nand U36036 (N_36036,N_35557,N_35540);
nand U36037 (N_36037,N_35433,N_35494);
xnor U36038 (N_36038,N_35906,N_35861);
xor U36039 (N_36039,N_35441,N_35243);
nor U36040 (N_36040,N_35932,N_35396);
xor U36041 (N_36041,N_35950,N_35800);
nor U36042 (N_36042,N_35068,N_35276);
xor U36043 (N_36043,N_35000,N_35792);
and U36044 (N_36044,N_35579,N_35809);
nor U36045 (N_36045,N_35166,N_35106);
nand U36046 (N_36046,N_35802,N_35931);
xor U36047 (N_36047,N_35211,N_35373);
xnor U36048 (N_36048,N_35070,N_35318);
and U36049 (N_36049,N_35703,N_35846);
nand U36050 (N_36050,N_35786,N_35140);
xnor U36051 (N_36051,N_35271,N_35887);
or U36052 (N_36052,N_35058,N_35165);
or U36053 (N_36053,N_35636,N_35653);
nand U36054 (N_36054,N_35548,N_35144);
or U36055 (N_36055,N_35761,N_35784);
or U36056 (N_36056,N_35285,N_35358);
and U36057 (N_36057,N_35524,N_35295);
nor U36058 (N_36058,N_35126,N_35721);
and U36059 (N_36059,N_35125,N_35905);
nand U36060 (N_36060,N_35273,N_35720);
or U36061 (N_36061,N_35261,N_35501);
nor U36062 (N_36062,N_35092,N_35860);
and U36063 (N_36063,N_35425,N_35762);
nand U36064 (N_36064,N_35816,N_35606);
nand U36065 (N_36065,N_35807,N_35313);
nand U36066 (N_36066,N_35082,N_35851);
xnor U36067 (N_36067,N_35879,N_35194);
xnor U36068 (N_36068,N_35646,N_35754);
and U36069 (N_36069,N_35844,N_35287);
and U36070 (N_36070,N_35526,N_35707);
and U36071 (N_36071,N_35922,N_35715);
or U36072 (N_36072,N_35399,N_35300);
nor U36073 (N_36073,N_35502,N_35940);
xnor U36074 (N_36074,N_35823,N_35655);
or U36075 (N_36075,N_35320,N_35622);
nor U36076 (N_36076,N_35943,N_35020);
xnor U36077 (N_36077,N_35207,N_35146);
xnor U36078 (N_36078,N_35888,N_35830);
nor U36079 (N_36079,N_35048,N_35156);
nand U36080 (N_36080,N_35246,N_35145);
xnor U36081 (N_36081,N_35237,N_35695);
nand U36082 (N_36082,N_35055,N_35779);
or U36083 (N_36083,N_35665,N_35828);
or U36084 (N_36084,N_35105,N_35102);
nand U36085 (N_36085,N_35726,N_35326);
or U36086 (N_36086,N_35551,N_35177);
or U36087 (N_36087,N_35505,N_35983);
nor U36088 (N_36088,N_35833,N_35120);
nand U36089 (N_36089,N_35705,N_35231);
nor U36090 (N_36090,N_35824,N_35480);
nor U36091 (N_36091,N_35445,N_35982);
or U36092 (N_36092,N_35236,N_35668);
and U36093 (N_36093,N_35644,N_35666);
nand U36094 (N_36094,N_35563,N_35472);
nand U36095 (N_36095,N_35974,N_35119);
and U36096 (N_36096,N_35926,N_35924);
nor U36097 (N_36097,N_35739,N_35895);
and U36098 (N_36098,N_35111,N_35151);
nor U36099 (N_36099,N_35022,N_35507);
and U36100 (N_36100,N_35722,N_35148);
nor U36101 (N_36101,N_35336,N_35930);
nand U36102 (N_36102,N_35232,N_35406);
or U36103 (N_36103,N_35976,N_35039);
nand U36104 (N_36104,N_35378,N_35451);
or U36105 (N_36105,N_35530,N_35925);
nand U36106 (N_36106,N_35789,N_35171);
nor U36107 (N_36107,N_35324,N_35770);
and U36108 (N_36108,N_35134,N_35727);
xnor U36109 (N_36109,N_35936,N_35116);
nand U36110 (N_36110,N_35112,N_35229);
xor U36111 (N_36111,N_35783,N_35253);
and U36112 (N_36112,N_35028,N_35725);
nor U36113 (N_36113,N_35235,N_35374);
or U36114 (N_36114,N_35553,N_35904);
nor U36115 (N_36115,N_35700,N_35202);
xnor U36116 (N_36116,N_35303,N_35957);
or U36117 (N_36117,N_35054,N_35118);
xnor U36118 (N_36118,N_35288,N_35691);
and U36119 (N_36119,N_35755,N_35723);
xor U36120 (N_36120,N_35334,N_35994);
or U36121 (N_36121,N_35918,N_35690);
and U36122 (N_36122,N_35123,N_35845);
nor U36123 (N_36123,N_35651,N_35663);
nand U36124 (N_36124,N_35442,N_35843);
or U36125 (N_36125,N_35624,N_35874);
nor U36126 (N_36126,N_35489,N_35522);
or U36127 (N_36127,N_35882,N_35541);
and U36128 (N_36128,N_35605,N_35585);
or U36129 (N_36129,N_35309,N_35900);
or U36130 (N_36130,N_35626,N_35510);
nor U36131 (N_36131,N_35339,N_35361);
and U36132 (N_36132,N_35377,N_35363);
nand U36133 (N_36133,N_35104,N_35220);
and U36134 (N_36134,N_35897,N_35084);
nor U36135 (N_36135,N_35286,N_35731);
or U36136 (N_36136,N_35591,N_35912);
and U36137 (N_36137,N_35580,N_35121);
and U36138 (N_36138,N_35688,N_35777);
xnor U36139 (N_36139,N_35488,N_35264);
nand U36140 (N_36140,N_35697,N_35408);
nand U36141 (N_36141,N_35035,N_35294);
and U36142 (N_36142,N_35678,N_35956);
or U36143 (N_36143,N_35711,N_35012);
and U36144 (N_36144,N_35460,N_35062);
or U36145 (N_36145,N_35928,N_35840);
xnor U36146 (N_36146,N_35534,N_35481);
and U36147 (N_36147,N_35967,N_35199);
nand U36148 (N_36148,N_35881,N_35959);
xnor U36149 (N_36149,N_35196,N_35497);
or U36150 (N_36150,N_35073,N_35410);
nor U36151 (N_36151,N_35517,N_35610);
nor U36152 (N_36152,N_35944,N_35461);
nand U36153 (N_36153,N_35677,N_35975);
or U36154 (N_36154,N_35589,N_35476);
or U36155 (N_36155,N_35255,N_35079);
nor U36156 (N_36156,N_35002,N_35949);
xnor U36157 (N_36157,N_35307,N_35364);
and U36158 (N_36158,N_35474,N_35531);
or U36159 (N_36159,N_35439,N_35576);
or U36160 (N_36160,N_35618,N_35600);
or U36161 (N_36161,N_35328,N_35629);
nor U36162 (N_36162,N_35159,N_35018);
xor U36163 (N_36163,N_35225,N_35942);
nand U36164 (N_36164,N_35026,N_35335);
nor U36165 (N_36165,N_35056,N_35291);
xnor U36166 (N_36166,N_35536,N_35167);
and U36167 (N_36167,N_35650,N_35333);
nand U36168 (N_36168,N_35164,N_35350);
xor U36169 (N_36169,N_35212,N_35430);
or U36170 (N_36170,N_35732,N_35803);
nand U36171 (N_36171,N_35245,N_35637);
nand U36172 (N_36172,N_35386,N_35868);
and U36173 (N_36173,N_35927,N_35508);
nor U36174 (N_36174,N_35438,N_35896);
or U36175 (N_36175,N_35150,N_35669);
nor U36176 (N_36176,N_35866,N_35327);
and U36177 (N_36177,N_35870,N_35617);
nor U36178 (N_36178,N_35710,N_35405);
or U36179 (N_36179,N_35750,N_35033);
or U36180 (N_36180,N_35174,N_35913);
and U36181 (N_36181,N_35724,N_35632);
and U36182 (N_36182,N_35921,N_35322);
or U36183 (N_36183,N_35574,N_35011);
nand U36184 (N_36184,N_35201,N_35889);
and U36185 (N_36185,N_35869,N_35640);
nor U36186 (N_36186,N_35547,N_35687);
nor U36187 (N_36187,N_35465,N_35290);
nor U36188 (N_36188,N_35811,N_35457);
nand U36189 (N_36189,N_35834,N_35964);
nand U36190 (N_36190,N_35603,N_35218);
nor U36191 (N_36191,N_35024,N_35746);
and U36192 (N_36192,N_35588,N_35985);
and U36193 (N_36193,N_35572,N_35961);
xnor U36194 (N_36194,N_35417,N_35768);
xor U36195 (N_36195,N_35359,N_35643);
xnor U36196 (N_36196,N_35516,N_35209);
nand U36197 (N_36197,N_35392,N_35990);
nor U36198 (N_36198,N_35475,N_35652);
and U36199 (N_36199,N_35421,N_35878);
and U36200 (N_36200,N_35190,N_35741);
or U36201 (N_36201,N_35321,N_35088);
nand U36202 (N_36202,N_35914,N_35384);
xnor U36203 (N_36203,N_35749,N_35404);
nand U36204 (N_36204,N_35304,N_35160);
and U36205 (N_36205,N_35010,N_35001);
nand U36206 (N_36206,N_35772,N_35314);
or U36207 (N_36207,N_35089,N_35479);
xor U36208 (N_36208,N_35242,N_35991);
nand U36209 (N_36209,N_35892,N_35027);
or U36210 (N_36210,N_35416,N_35268);
and U36211 (N_36211,N_35858,N_35446);
or U36212 (N_36212,N_35157,N_35015);
and U36213 (N_36213,N_35751,N_35337);
nand U36214 (N_36214,N_35987,N_35331);
xnor U36215 (N_36215,N_35204,N_35319);
or U36216 (N_36216,N_35130,N_35186);
or U36217 (N_36217,N_35767,N_35701);
or U36218 (N_36218,N_35554,N_35228);
nand U36219 (N_36219,N_35176,N_35818);
xnor U36220 (N_36220,N_35933,N_35667);
nand U36221 (N_36221,N_35561,N_35623);
nand U36222 (N_36222,N_35244,N_35763);
nor U36223 (N_36223,N_35259,N_35042);
and U36224 (N_36224,N_35272,N_35744);
nand U36225 (N_36225,N_35712,N_35564);
nand U36226 (N_36226,N_35464,N_35077);
xnor U36227 (N_36227,N_35670,N_35616);
nand U36228 (N_36228,N_35794,N_35306);
or U36229 (N_36229,N_35674,N_35274);
and U36230 (N_36230,N_35627,N_35556);
xnor U36231 (N_36231,N_35437,N_35389);
nor U36232 (N_36232,N_35061,N_35743);
nand U36233 (N_36233,N_35275,N_35312);
and U36234 (N_36234,N_35490,N_35277);
or U36235 (N_36235,N_35997,N_35367);
or U36236 (N_36236,N_35612,N_35988);
or U36237 (N_36237,N_35305,N_35041);
nand U36238 (N_36238,N_35091,N_35482);
or U36239 (N_36239,N_35771,N_35411);
nor U36240 (N_36240,N_35469,N_35192);
nand U36241 (N_36241,N_35473,N_35704);
nor U36242 (N_36242,N_35594,N_35368);
xor U36243 (N_36243,N_35560,N_35103);
and U36244 (N_36244,N_35447,N_35060);
xor U36245 (N_36245,N_35853,N_35641);
or U36246 (N_36246,N_35127,N_35071);
nor U36247 (N_36247,N_35347,N_35296);
nand U36248 (N_36248,N_35550,N_35635);
nand U36249 (N_36249,N_35535,N_35013);
xnor U36250 (N_36250,N_35902,N_35289);
nand U36251 (N_36251,N_35671,N_35049);
xor U36252 (N_36252,N_35571,N_35596);
xnor U36253 (N_36253,N_35124,N_35598);
and U36254 (N_36254,N_35390,N_35269);
nand U36255 (N_36255,N_35920,N_35346);
xnor U36256 (N_36256,N_35864,N_35059);
nand U36257 (N_36257,N_35873,N_35310);
nor U36258 (N_36258,N_35647,N_35233);
xnor U36259 (N_36259,N_35040,N_35342);
xnor U36260 (N_36260,N_35593,N_35354);
and U36261 (N_36261,N_35095,N_35149);
nand U36262 (N_36262,N_35562,N_35978);
xor U36263 (N_36263,N_35543,N_35578);
nor U36264 (N_36264,N_35788,N_35135);
or U36265 (N_36265,N_35485,N_35297);
xnor U36266 (N_36266,N_35032,N_35267);
xor U36267 (N_36267,N_35847,N_35810);
nand U36268 (N_36268,N_35679,N_35302);
nor U36269 (N_36269,N_35702,N_35821);
nor U36270 (N_36270,N_35613,N_35766);
nor U36271 (N_36271,N_35774,N_35064);
nor U36272 (N_36272,N_35570,N_35325);
nand U36273 (N_36273,N_35848,N_35227);
nor U36274 (N_36274,N_35353,N_35587);
xnor U36275 (N_36275,N_35999,N_35708);
nand U36276 (N_36276,N_35098,N_35383);
nand U36277 (N_36277,N_35279,N_35155);
or U36278 (N_36278,N_35787,N_35136);
nand U36279 (N_36279,N_35179,N_35996);
xor U36280 (N_36280,N_35008,N_35935);
nand U36281 (N_36281,N_35831,N_35216);
xnor U36282 (N_36282,N_35625,N_35813);
xor U36283 (N_36283,N_35397,N_35759);
or U36284 (N_36284,N_35523,N_35402);
nor U36285 (N_36285,N_35282,N_35178);
and U36286 (N_36286,N_35518,N_35142);
and U36287 (N_36287,N_35521,N_35413);
xor U36288 (N_36288,N_35065,N_35947);
nand U36289 (N_36289,N_35778,N_35412);
nor U36290 (N_36290,N_35929,N_35050);
and U36291 (N_36291,N_35343,N_35131);
nor U36292 (N_36292,N_35854,N_35965);
nor U36293 (N_36293,N_35226,N_35814);
nor U36294 (N_36294,N_35907,N_35265);
nand U36295 (N_36295,N_35515,N_35398);
and U36296 (N_36296,N_35141,N_35395);
nand U36297 (N_36297,N_35529,N_35709);
or U36298 (N_36298,N_35654,N_35492);
nand U36299 (N_36299,N_35952,N_35909);
and U36300 (N_36300,N_35191,N_35590);
nor U36301 (N_36301,N_35658,N_35449);
nor U36302 (N_36302,N_35863,N_35699);
and U36303 (N_36303,N_35797,N_35184);
nand U36304 (N_36304,N_35498,N_35954);
xor U36305 (N_36305,N_35239,N_35962);
and U36306 (N_36306,N_35025,N_35340);
and U36307 (N_36307,N_35946,N_35747);
and U36308 (N_36308,N_35238,N_35638);
or U36309 (N_36309,N_35491,N_35675);
and U36310 (N_36310,N_35642,N_35349);
xnor U36311 (N_36311,N_35034,N_35298);
xor U36312 (N_36312,N_35742,N_35484);
or U36313 (N_36313,N_35376,N_35717);
nor U36314 (N_36314,N_35734,N_35162);
xor U36315 (N_36315,N_35716,N_35938);
and U36316 (N_36316,N_35819,N_35886);
nor U36317 (N_36317,N_35459,N_35528);
and U36318 (N_36318,N_35764,N_35981);
or U36319 (N_36319,N_35728,N_35407);
nand U36320 (N_36320,N_35036,N_35467);
nor U36321 (N_36321,N_35825,N_35428);
nor U36322 (N_36322,N_35317,N_35352);
and U36323 (N_36323,N_35208,N_35031);
nand U36324 (N_36324,N_35432,N_35757);
or U36325 (N_36325,N_35110,N_35085);
and U36326 (N_36326,N_35189,N_35953);
nand U36327 (N_36327,N_35213,N_35258);
nor U36328 (N_36328,N_35841,N_35486);
nand U36329 (N_36329,N_35487,N_35500);
and U36330 (N_36330,N_35607,N_35117);
xor U36331 (N_36331,N_35147,N_35069);
nand U36332 (N_36332,N_35210,N_35496);
nand U36333 (N_36333,N_35038,N_35153);
nand U36334 (N_36334,N_35586,N_35043);
nor U36335 (N_36335,N_35007,N_35086);
xor U36336 (N_36336,N_35545,N_35401);
nand U36337 (N_36337,N_35075,N_35884);
and U36338 (N_36338,N_35241,N_35369);
nand U36339 (N_36339,N_35738,N_35169);
nand U36340 (N_36340,N_35737,N_35682);
or U36341 (N_36341,N_35733,N_35867);
and U36342 (N_36342,N_35422,N_35356);
nor U36343 (N_36343,N_35649,N_35781);
nand U36344 (N_36344,N_35939,N_35076);
and U36345 (N_36345,N_35718,N_35128);
xor U36346 (N_36346,N_35375,N_35549);
nand U36347 (N_36347,N_35804,N_35817);
xnor U36348 (N_36348,N_35963,N_35195);
xor U36349 (N_36349,N_35765,N_35620);
and U36350 (N_36350,N_35758,N_35139);
and U36351 (N_36351,N_35672,N_35163);
nand U36352 (N_36352,N_35736,N_35849);
and U36353 (N_36353,N_35934,N_35250);
or U36354 (N_36354,N_35424,N_35512);
or U36355 (N_36355,N_35426,N_35219);
and U36356 (N_36356,N_35493,N_35628);
or U36357 (N_36357,N_35357,N_35815);
nand U36358 (N_36358,N_35532,N_35360);
and U36359 (N_36359,N_35948,N_35419);
and U36360 (N_36360,N_35542,N_35850);
nor U36361 (N_36361,N_35187,N_35684);
and U36362 (N_36362,N_35566,N_35394);
nand U36363 (N_36363,N_35081,N_35283);
and U36364 (N_36364,N_35161,N_35835);
xnor U36365 (N_36365,N_35030,N_35180);
and U36366 (N_36366,N_35837,N_35760);
or U36367 (N_36367,N_35748,N_35951);
nand U36368 (N_36368,N_35137,N_35021);
or U36369 (N_36369,N_35855,N_35871);
nand U36370 (N_36370,N_35051,N_35793);
and U36371 (N_36371,N_35645,N_35693);
nand U36372 (N_36372,N_35910,N_35698);
and U36373 (N_36373,N_35769,N_35254);
or U36374 (N_36374,N_35418,N_35753);
nand U36375 (N_36375,N_35370,N_35630);
xor U36376 (N_36376,N_35706,N_35595);
and U36377 (N_36377,N_35108,N_35152);
nor U36378 (N_36378,N_35972,N_35575);
or U36379 (N_36379,N_35842,N_35838);
xnor U36380 (N_36380,N_35045,N_35101);
nor U36381 (N_36381,N_35898,N_35047);
nand U36382 (N_36382,N_35053,N_35558);
xnor U36383 (N_36383,N_35478,N_35796);
or U36384 (N_36384,N_35614,N_35681);
or U36385 (N_36385,N_35455,N_35323);
or U36386 (N_36386,N_35567,N_35017);
nor U36387 (N_36387,N_35511,N_35569);
xnor U36388 (N_36388,N_35247,N_35692);
or U36389 (N_36389,N_35224,N_35903);
nand U36390 (N_36390,N_35533,N_35601);
xnor U36391 (N_36391,N_35381,N_35188);
or U36392 (N_36392,N_35885,N_35366);
and U36393 (N_36393,N_35181,N_35230);
nand U36394 (N_36394,N_35173,N_35602);
xor U36395 (N_36395,N_35740,N_35221);
or U36396 (N_36396,N_35513,N_35509);
or U36397 (N_36397,N_35504,N_35862);
xor U36398 (N_36398,N_35832,N_35877);
nand U36399 (N_36399,N_35270,N_35970);
nand U36400 (N_36400,N_35429,N_35090);
xnor U36401 (N_36401,N_35555,N_35436);
nor U36402 (N_36402,N_35217,N_35372);
and U36403 (N_36403,N_35072,N_35719);
and U36404 (N_36404,N_35799,N_35198);
or U36405 (N_36405,N_35968,N_35109);
xnor U36406 (N_36406,N_35138,N_35222);
xor U36407 (N_36407,N_35093,N_35689);
or U36408 (N_36408,N_35471,N_35894);
nor U36409 (N_36409,N_35046,N_35278);
or U36410 (N_36410,N_35351,N_35893);
and U36411 (N_36411,N_35004,N_35260);
and U36412 (N_36412,N_35984,N_35775);
and U36413 (N_36413,N_35608,N_35044);
nor U36414 (N_36414,N_35621,N_35132);
nor U36415 (N_36415,N_35158,N_35214);
nor U36416 (N_36416,N_35454,N_35609);
and U36417 (N_36417,N_35780,N_35052);
nand U36418 (N_36418,N_35385,N_35330);
and U36419 (N_36419,N_35263,N_35782);
xnor U36420 (N_36420,N_35067,N_35735);
nor U36421 (N_36421,N_35183,N_35546);
xor U36422 (N_36422,N_35776,N_35185);
nor U36423 (N_36423,N_35773,N_35443);
nand U36424 (N_36424,N_35908,N_35519);
or U36425 (N_36425,N_35584,N_35133);
nand U36426 (N_36426,N_35812,N_35114);
and U36427 (N_36427,N_35503,N_35659);
xnor U36428 (N_36428,N_35434,N_35899);
nor U36429 (N_36429,N_35345,N_35470);
or U36430 (N_36430,N_35955,N_35573);
nand U36431 (N_36431,N_35798,N_35099);
xnor U36432 (N_36432,N_35664,N_35685);
or U36433 (N_36433,N_35880,N_35941);
nand U36434 (N_36434,N_35450,N_35552);
or U36435 (N_36435,N_35248,N_35785);
nand U36436 (N_36436,N_35029,N_35795);
nor U36437 (N_36437,N_35009,N_35308);
or U36438 (N_36438,N_35696,N_35657);
or U36439 (N_36439,N_35129,N_35063);
xor U36440 (N_36440,N_35115,N_35414);
or U36441 (N_36441,N_35559,N_35859);
or U36442 (N_36442,N_35916,N_35633);
nor U36443 (N_36443,N_35182,N_35592);
and U36444 (N_36444,N_35986,N_35371);
and U36445 (N_36445,N_35019,N_35539);
xnor U36446 (N_36446,N_35568,N_35960);
nor U36447 (N_36447,N_35631,N_35382);
or U36448 (N_36448,N_35998,N_35100);
or U36449 (N_36449,N_35915,N_35839);
and U36450 (N_36450,N_35400,N_35958);
xor U36451 (N_36451,N_35362,N_35872);
or U36452 (N_36452,N_35329,N_35901);
or U36453 (N_36453,N_35756,N_35087);
nor U36454 (N_36454,N_35280,N_35805);
nand U36455 (N_36455,N_35316,N_35662);
and U36456 (N_36456,N_35966,N_35266);
nor U36457 (N_36457,N_35348,N_35937);
nand U36458 (N_36458,N_35730,N_35240);
nand U36459 (N_36459,N_35791,N_35420);
and U36460 (N_36460,N_35891,N_35252);
and U36461 (N_36461,N_35444,N_35993);
or U36462 (N_36462,N_35281,N_35680);
xnor U36463 (N_36463,N_35083,N_35074);
or U36464 (N_36464,N_35883,N_35452);
xor U36465 (N_36465,N_35694,N_35016);
or U36466 (N_36466,N_35686,N_35683);
xnor U36467 (N_36467,N_35249,N_35806);
xor U36468 (N_36468,N_35003,N_35200);
nor U36469 (N_36469,N_35458,N_35223);
nor U36470 (N_36470,N_35462,N_35468);
xor U36471 (N_36471,N_35969,N_35829);
nor U36472 (N_36472,N_35483,N_35094);
and U36473 (N_36473,N_35415,N_35857);
nor U36474 (N_36474,N_35203,N_35619);
xor U36475 (N_36475,N_35977,N_35676);
nand U36476 (N_36476,N_35107,N_35537);
nand U36477 (N_36477,N_35945,N_35409);
nand U36478 (N_36478,N_35097,N_35251);
nand U36479 (N_36479,N_35379,N_35527);
or U36480 (N_36480,N_35435,N_35154);
and U36481 (N_36481,N_35971,N_35634);
nand U36482 (N_36482,N_35023,N_35820);
nand U36483 (N_36483,N_35995,N_35852);
nor U36484 (N_36484,N_35080,N_35175);
or U36485 (N_36485,N_35463,N_35856);
or U36486 (N_36486,N_35827,N_35911);
nand U36487 (N_36487,N_35973,N_35403);
or U36488 (N_36488,N_35876,N_35193);
nor U36489 (N_36489,N_35729,N_35431);
or U36490 (N_36490,N_35477,N_35448);
xnor U36491 (N_36491,N_35923,N_35341);
nor U36492 (N_36492,N_35143,N_35315);
nand U36493 (N_36493,N_35257,N_35380);
nor U36494 (N_36494,N_35365,N_35673);
or U36495 (N_36495,N_35311,N_35822);
nand U36496 (N_36496,N_35599,N_35096);
nand U36497 (N_36497,N_35919,N_35387);
xnor U36498 (N_36498,N_35344,N_35206);
nand U36499 (N_36499,N_35423,N_35875);
and U36500 (N_36500,N_35205,N_35236);
xnor U36501 (N_36501,N_35594,N_35868);
nand U36502 (N_36502,N_35519,N_35383);
nor U36503 (N_36503,N_35735,N_35277);
and U36504 (N_36504,N_35900,N_35012);
nand U36505 (N_36505,N_35518,N_35513);
and U36506 (N_36506,N_35587,N_35601);
xnor U36507 (N_36507,N_35025,N_35757);
or U36508 (N_36508,N_35680,N_35557);
or U36509 (N_36509,N_35080,N_35816);
nand U36510 (N_36510,N_35510,N_35613);
xnor U36511 (N_36511,N_35635,N_35388);
nor U36512 (N_36512,N_35591,N_35211);
nor U36513 (N_36513,N_35191,N_35210);
nor U36514 (N_36514,N_35968,N_35382);
nor U36515 (N_36515,N_35993,N_35754);
and U36516 (N_36516,N_35281,N_35423);
xnor U36517 (N_36517,N_35517,N_35747);
or U36518 (N_36518,N_35849,N_35191);
and U36519 (N_36519,N_35812,N_35088);
and U36520 (N_36520,N_35624,N_35183);
or U36521 (N_36521,N_35393,N_35772);
nand U36522 (N_36522,N_35975,N_35052);
xnor U36523 (N_36523,N_35012,N_35499);
nor U36524 (N_36524,N_35639,N_35973);
and U36525 (N_36525,N_35679,N_35077);
nand U36526 (N_36526,N_35381,N_35143);
nand U36527 (N_36527,N_35957,N_35512);
and U36528 (N_36528,N_35320,N_35436);
and U36529 (N_36529,N_35904,N_35644);
nand U36530 (N_36530,N_35745,N_35079);
and U36531 (N_36531,N_35534,N_35239);
xor U36532 (N_36532,N_35040,N_35608);
xnor U36533 (N_36533,N_35028,N_35356);
nand U36534 (N_36534,N_35184,N_35166);
xnor U36535 (N_36535,N_35719,N_35100);
xor U36536 (N_36536,N_35762,N_35195);
xor U36537 (N_36537,N_35059,N_35930);
xor U36538 (N_36538,N_35848,N_35907);
or U36539 (N_36539,N_35443,N_35738);
nor U36540 (N_36540,N_35118,N_35155);
and U36541 (N_36541,N_35249,N_35945);
or U36542 (N_36542,N_35790,N_35108);
nor U36543 (N_36543,N_35880,N_35980);
nor U36544 (N_36544,N_35541,N_35180);
and U36545 (N_36545,N_35552,N_35183);
and U36546 (N_36546,N_35641,N_35050);
and U36547 (N_36547,N_35483,N_35339);
nand U36548 (N_36548,N_35464,N_35384);
xor U36549 (N_36549,N_35486,N_35455);
and U36550 (N_36550,N_35137,N_35858);
xor U36551 (N_36551,N_35770,N_35276);
or U36552 (N_36552,N_35086,N_35040);
xnor U36553 (N_36553,N_35193,N_35520);
xnor U36554 (N_36554,N_35540,N_35659);
nand U36555 (N_36555,N_35559,N_35590);
or U36556 (N_36556,N_35047,N_35819);
and U36557 (N_36557,N_35586,N_35809);
nand U36558 (N_36558,N_35166,N_35932);
and U36559 (N_36559,N_35859,N_35801);
nand U36560 (N_36560,N_35975,N_35277);
nor U36561 (N_36561,N_35965,N_35529);
xnor U36562 (N_36562,N_35591,N_35680);
nor U36563 (N_36563,N_35378,N_35220);
xnor U36564 (N_36564,N_35395,N_35109);
xor U36565 (N_36565,N_35319,N_35576);
and U36566 (N_36566,N_35941,N_35686);
and U36567 (N_36567,N_35277,N_35627);
and U36568 (N_36568,N_35018,N_35767);
nor U36569 (N_36569,N_35307,N_35224);
nor U36570 (N_36570,N_35173,N_35500);
xnor U36571 (N_36571,N_35117,N_35915);
and U36572 (N_36572,N_35662,N_35425);
or U36573 (N_36573,N_35740,N_35480);
nand U36574 (N_36574,N_35356,N_35994);
xor U36575 (N_36575,N_35196,N_35679);
xnor U36576 (N_36576,N_35832,N_35115);
nand U36577 (N_36577,N_35358,N_35459);
nand U36578 (N_36578,N_35146,N_35194);
nand U36579 (N_36579,N_35529,N_35304);
xnor U36580 (N_36580,N_35763,N_35581);
xor U36581 (N_36581,N_35439,N_35558);
and U36582 (N_36582,N_35960,N_35497);
and U36583 (N_36583,N_35118,N_35187);
nor U36584 (N_36584,N_35476,N_35313);
nand U36585 (N_36585,N_35642,N_35831);
nor U36586 (N_36586,N_35510,N_35539);
and U36587 (N_36587,N_35230,N_35220);
xor U36588 (N_36588,N_35404,N_35900);
nor U36589 (N_36589,N_35697,N_35169);
nor U36590 (N_36590,N_35929,N_35090);
nor U36591 (N_36591,N_35225,N_35197);
and U36592 (N_36592,N_35583,N_35595);
xor U36593 (N_36593,N_35952,N_35805);
nor U36594 (N_36594,N_35942,N_35341);
xor U36595 (N_36595,N_35527,N_35270);
nor U36596 (N_36596,N_35833,N_35719);
nand U36597 (N_36597,N_35854,N_35897);
and U36598 (N_36598,N_35350,N_35316);
or U36599 (N_36599,N_35801,N_35301);
or U36600 (N_36600,N_35013,N_35752);
xor U36601 (N_36601,N_35131,N_35464);
and U36602 (N_36602,N_35825,N_35222);
nand U36603 (N_36603,N_35141,N_35657);
nor U36604 (N_36604,N_35116,N_35422);
nand U36605 (N_36605,N_35720,N_35789);
nor U36606 (N_36606,N_35139,N_35330);
and U36607 (N_36607,N_35065,N_35025);
nor U36608 (N_36608,N_35470,N_35696);
and U36609 (N_36609,N_35071,N_35781);
nand U36610 (N_36610,N_35924,N_35672);
or U36611 (N_36611,N_35709,N_35998);
nand U36612 (N_36612,N_35385,N_35678);
xor U36613 (N_36613,N_35462,N_35118);
nand U36614 (N_36614,N_35980,N_35606);
or U36615 (N_36615,N_35763,N_35019);
and U36616 (N_36616,N_35633,N_35261);
and U36617 (N_36617,N_35312,N_35417);
nor U36618 (N_36618,N_35577,N_35141);
nand U36619 (N_36619,N_35030,N_35731);
nand U36620 (N_36620,N_35416,N_35312);
xor U36621 (N_36621,N_35106,N_35900);
nand U36622 (N_36622,N_35878,N_35596);
nand U36623 (N_36623,N_35270,N_35606);
or U36624 (N_36624,N_35997,N_35343);
nor U36625 (N_36625,N_35879,N_35286);
or U36626 (N_36626,N_35569,N_35092);
xor U36627 (N_36627,N_35498,N_35564);
or U36628 (N_36628,N_35375,N_35855);
or U36629 (N_36629,N_35434,N_35965);
or U36630 (N_36630,N_35615,N_35277);
nand U36631 (N_36631,N_35616,N_35076);
nand U36632 (N_36632,N_35720,N_35589);
xnor U36633 (N_36633,N_35771,N_35696);
and U36634 (N_36634,N_35653,N_35775);
or U36635 (N_36635,N_35805,N_35643);
xor U36636 (N_36636,N_35300,N_35386);
or U36637 (N_36637,N_35654,N_35432);
xor U36638 (N_36638,N_35083,N_35700);
or U36639 (N_36639,N_35046,N_35403);
nand U36640 (N_36640,N_35248,N_35529);
or U36641 (N_36641,N_35916,N_35045);
or U36642 (N_36642,N_35649,N_35384);
nor U36643 (N_36643,N_35745,N_35677);
nor U36644 (N_36644,N_35464,N_35351);
xnor U36645 (N_36645,N_35683,N_35752);
xor U36646 (N_36646,N_35240,N_35470);
nor U36647 (N_36647,N_35205,N_35645);
nand U36648 (N_36648,N_35480,N_35505);
and U36649 (N_36649,N_35758,N_35164);
or U36650 (N_36650,N_35128,N_35382);
nor U36651 (N_36651,N_35585,N_35547);
or U36652 (N_36652,N_35011,N_35490);
or U36653 (N_36653,N_35129,N_35080);
nand U36654 (N_36654,N_35823,N_35447);
nor U36655 (N_36655,N_35701,N_35033);
nor U36656 (N_36656,N_35522,N_35465);
nor U36657 (N_36657,N_35425,N_35897);
nand U36658 (N_36658,N_35481,N_35951);
nand U36659 (N_36659,N_35265,N_35982);
xnor U36660 (N_36660,N_35286,N_35543);
nor U36661 (N_36661,N_35343,N_35893);
xnor U36662 (N_36662,N_35945,N_35230);
nand U36663 (N_36663,N_35126,N_35899);
and U36664 (N_36664,N_35927,N_35901);
nand U36665 (N_36665,N_35793,N_35574);
and U36666 (N_36666,N_35160,N_35059);
or U36667 (N_36667,N_35632,N_35257);
nand U36668 (N_36668,N_35295,N_35594);
or U36669 (N_36669,N_35620,N_35911);
nand U36670 (N_36670,N_35376,N_35874);
or U36671 (N_36671,N_35319,N_35122);
or U36672 (N_36672,N_35187,N_35144);
nand U36673 (N_36673,N_35523,N_35098);
xor U36674 (N_36674,N_35085,N_35700);
xnor U36675 (N_36675,N_35257,N_35283);
nand U36676 (N_36676,N_35646,N_35922);
and U36677 (N_36677,N_35767,N_35053);
and U36678 (N_36678,N_35112,N_35377);
or U36679 (N_36679,N_35142,N_35575);
nand U36680 (N_36680,N_35000,N_35995);
nor U36681 (N_36681,N_35173,N_35307);
nand U36682 (N_36682,N_35859,N_35294);
nor U36683 (N_36683,N_35177,N_35232);
nor U36684 (N_36684,N_35296,N_35553);
xor U36685 (N_36685,N_35357,N_35558);
nand U36686 (N_36686,N_35450,N_35638);
nor U36687 (N_36687,N_35963,N_35549);
nor U36688 (N_36688,N_35044,N_35241);
or U36689 (N_36689,N_35458,N_35583);
nor U36690 (N_36690,N_35465,N_35568);
xor U36691 (N_36691,N_35734,N_35707);
nor U36692 (N_36692,N_35574,N_35497);
nor U36693 (N_36693,N_35944,N_35212);
nor U36694 (N_36694,N_35280,N_35322);
nand U36695 (N_36695,N_35514,N_35347);
xnor U36696 (N_36696,N_35809,N_35640);
nand U36697 (N_36697,N_35205,N_35513);
and U36698 (N_36698,N_35114,N_35473);
xor U36699 (N_36699,N_35468,N_35045);
or U36700 (N_36700,N_35513,N_35049);
xnor U36701 (N_36701,N_35265,N_35037);
nor U36702 (N_36702,N_35454,N_35903);
or U36703 (N_36703,N_35167,N_35216);
xnor U36704 (N_36704,N_35513,N_35743);
nand U36705 (N_36705,N_35413,N_35518);
xnor U36706 (N_36706,N_35199,N_35222);
nor U36707 (N_36707,N_35435,N_35151);
or U36708 (N_36708,N_35206,N_35602);
xnor U36709 (N_36709,N_35799,N_35515);
nor U36710 (N_36710,N_35019,N_35778);
nor U36711 (N_36711,N_35084,N_35661);
and U36712 (N_36712,N_35779,N_35435);
and U36713 (N_36713,N_35828,N_35300);
nor U36714 (N_36714,N_35259,N_35724);
xnor U36715 (N_36715,N_35682,N_35769);
or U36716 (N_36716,N_35377,N_35813);
and U36717 (N_36717,N_35260,N_35601);
nand U36718 (N_36718,N_35947,N_35311);
xor U36719 (N_36719,N_35446,N_35081);
and U36720 (N_36720,N_35084,N_35337);
xor U36721 (N_36721,N_35420,N_35207);
nand U36722 (N_36722,N_35830,N_35764);
xnor U36723 (N_36723,N_35414,N_35216);
nor U36724 (N_36724,N_35547,N_35120);
or U36725 (N_36725,N_35640,N_35669);
xnor U36726 (N_36726,N_35938,N_35953);
or U36727 (N_36727,N_35835,N_35504);
nand U36728 (N_36728,N_35323,N_35868);
nand U36729 (N_36729,N_35143,N_35276);
and U36730 (N_36730,N_35281,N_35011);
or U36731 (N_36731,N_35670,N_35964);
or U36732 (N_36732,N_35663,N_35466);
nand U36733 (N_36733,N_35088,N_35158);
and U36734 (N_36734,N_35627,N_35674);
xor U36735 (N_36735,N_35692,N_35257);
nand U36736 (N_36736,N_35721,N_35239);
xor U36737 (N_36737,N_35897,N_35791);
nand U36738 (N_36738,N_35784,N_35378);
or U36739 (N_36739,N_35275,N_35669);
xor U36740 (N_36740,N_35815,N_35323);
xnor U36741 (N_36741,N_35796,N_35872);
nand U36742 (N_36742,N_35095,N_35791);
and U36743 (N_36743,N_35562,N_35278);
xor U36744 (N_36744,N_35366,N_35708);
nor U36745 (N_36745,N_35889,N_35532);
xnor U36746 (N_36746,N_35277,N_35426);
nor U36747 (N_36747,N_35833,N_35094);
nand U36748 (N_36748,N_35200,N_35498);
nor U36749 (N_36749,N_35361,N_35491);
nand U36750 (N_36750,N_35494,N_35476);
nor U36751 (N_36751,N_35707,N_35092);
and U36752 (N_36752,N_35503,N_35946);
and U36753 (N_36753,N_35383,N_35254);
xnor U36754 (N_36754,N_35887,N_35834);
nor U36755 (N_36755,N_35438,N_35239);
nor U36756 (N_36756,N_35753,N_35358);
nor U36757 (N_36757,N_35548,N_35183);
nand U36758 (N_36758,N_35443,N_35341);
xor U36759 (N_36759,N_35041,N_35132);
nor U36760 (N_36760,N_35415,N_35506);
nand U36761 (N_36761,N_35788,N_35294);
and U36762 (N_36762,N_35513,N_35438);
xnor U36763 (N_36763,N_35878,N_35137);
or U36764 (N_36764,N_35404,N_35541);
or U36765 (N_36765,N_35937,N_35605);
nand U36766 (N_36766,N_35670,N_35309);
or U36767 (N_36767,N_35965,N_35476);
nand U36768 (N_36768,N_35806,N_35596);
and U36769 (N_36769,N_35047,N_35005);
and U36770 (N_36770,N_35308,N_35343);
nor U36771 (N_36771,N_35927,N_35299);
xor U36772 (N_36772,N_35536,N_35537);
or U36773 (N_36773,N_35863,N_35911);
or U36774 (N_36774,N_35813,N_35069);
or U36775 (N_36775,N_35843,N_35323);
nand U36776 (N_36776,N_35869,N_35266);
nand U36777 (N_36777,N_35479,N_35727);
and U36778 (N_36778,N_35862,N_35019);
and U36779 (N_36779,N_35470,N_35342);
or U36780 (N_36780,N_35046,N_35561);
and U36781 (N_36781,N_35144,N_35840);
xor U36782 (N_36782,N_35013,N_35595);
nand U36783 (N_36783,N_35392,N_35074);
xnor U36784 (N_36784,N_35121,N_35432);
nand U36785 (N_36785,N_35825,N_35335);
and U36786 (N_36786,N_35671,N_35840);
nand U36787 (N_36787,N_35778,N_35069);
and U36788 (N_36788,N_35636,N_35901);
and U36789 (N_36789,N_35436,N_35772);
or U36790 (N_36790,N_35543,N_35170);
nor U36791 (N_36791,N_35394,N_35046);
and U36792 (N_36792,N_35563,N_35327);
or U36793 (N_36793,N_35756,N_35305);
or U36794 (N_36794,N_35241,N_35132);
nor U36795 (N_36795,N_35401,N_35501);
nand U36796 (N_36796,N_35758,N_35503);
nand U36797 (N_36797,N_35369,N_35880);
or U36798 (N_36798,N_35605,N_35765);
and U36799 (N_36799,N_35591,N_35008);
and U36800 (N_36800,N_35632,N_35173);
nor U36801 (N_36801,N_35629,N_35786);
nand U36802 (N_36802,N_35204,N_35693);
xnor U36803 (N_36803,N_35189,N_35686);
and U36804 (N_36804,N_35524,N_35167);
or U36805 (N_36805,N_35569,N_35358);
and U36806 (N_36806,N_35614,N_35823);
xor U36807 (N_36807,N_35532,N_35847);
nand U36808 (N_36808,N_35126,N_35235);
or U36809 (N_36809,N_35174,N_35530);
nor U36810 (N_36810,N_35394,N_35963);
nand U36811 (N_36811,N_35548,N_35968);
and U36812 (N_36812,N_35807,N_35063);
and U36813 (N_36813,N_35644,N_35372);
xnor U36814 (N_36814,N_35010,N_35797);
nor U36815 (N_36815,N_35626,N_35031);
nor U36816 (N_36816,N_35204,N_35110);
xor U36817 (N_36817,N_35703,N_35004);
nand U36818 (N_36818,N_35282,N_35699);
nor U36819 (N_36819,N_35798,N_35406);
nor U36820 (N_36820,N_35877,N_35263);
nand U36821 (N_36821,N_35230,N_35437);
or U36822 (N_36822,N_35964,N_35293);
or U36823 (N_36823,N_35154,N_35743);
and U36824 (N_36824,N_35624,N_35259);
xnor U36825 (N_36825,N_35998,N_35593);
xnor U36826 (N_36826,N_35485,N_35868);
and U36827 (N_36827,N_35442,N_35022);
nor U36828 (N_36828,N_35085,N_35672);
nand U36829 (N_36829,N_35792,N_35064);
or U36830 (N_36830,N_35612,N_35861);
xnor U36831 (N_36831,N_35201,N_35757);
nor U36832 (N_36832,N_35547,N_35466);
nand U36833 (N_36833,N_35931,N_35554);
nor U36834 (N_36834,N_35132,N_35724);
and U36835 (N_36835,N_35765,N_35297);
and U36836 (N_36836,N_35816,N_35632);
nor U36837 (N_36837,N_35497,N_35202);
xor U36838 (N_36838,N_35323,N_35753);
xor U36839 (N_36839,N_35598,N_35255);
nor U36840 (N_36840,N_35155,N_35223);
nand U36841 (N_36841,N_35985,N_35560);
nand U36842 (N_36842,N_35405,N_35332);
nor U36843 (N_36843,N_35114,N_35882);
nor U36844 (N_36844,N_35730,N_35073);
and U36845 (N_36845,N_35153,N_35708);
nand U36846 (N_36846,N_35637,N_35387);
nor U36847 (N_36847,N_35962,N_35114);
nor U36848 (N_36848,N_35055,N_35780);
or U36849 (N_36849,N_35184,N_35040);
nor U36850 (N_36850,N_35091,N_35825);
nor U36851 (N_36851,N_35684,N_35590);
xor U36852 (N_36852,N_35210,N_35713);
and U36853 (N_36853,N_35777,N_35171);
nand U36854 (N_36854,N_35451,N_35542);
and U36855 (N_36855,N_35571,N_35434);
and U36856 (N_36856,N_35989,N_35041);
nand U36857 (N_36857,N_35851,N_35716);
and U36858 (N_36858,N_35818,N_35132);
xnor U36859 (N_36859,N_35291,N_35710);
xor U36860 (N_36860,N_35509,N_35763);
xor U36861 (N_36861,N_35938,N_35710);
nand U36862 (N_36862,N_35265,N_35051);
xor U36863 (N_36863,N_35988,N_35627);
nand U36864 (N_36864,N_35438,N_35706);
and U36865 (N_36865,N_35883,N_35727);
and U36866 (N_36866,N_35875,N_35397);
nand U36867 (N_36867,N_35519,N_35983);
or U36868 (N_36868,N_35934,N_35017);
xor U36869 (N_36869,N_35547,N_35768);
xor U36870 (N_36870,N_35120,N_35915);
xor U36871 (N_36871,N_35193,N_35072);
nand U36872 (N_36872,N_35904,N_35230);
xnor U36873 (N_36873,N_35857,N_35870);
xnor U36874 (N_36874,N_35133,N_35673);
xnor U36875 (N_36875,N_35373,N_35071);
xnor U36876 (N_36876,N_35462,N_35861);
and U36877 (N_36877,N_35993,N_35073);
or U36878 (N_36878,N_35619,N_35327);
nor U36879 (N_36879,N_35914,N_35666);
and U36880 (N_36880,N_35739,N_35488);
or U36881 (N_36881,N_35652,N_35011);
xnor U36882 (N_36882,N_35165,N_35582);
nand U36883 (N_36883,N_35458,N_35318);
xor U36884 (N_36884,N_35378,N_35044);
and U36885 (N_36885,N_35785,N_35132);
and U36886 (N_36886,N_35294,N_35926);
xnor U36887 (N_36887,N_35570,N_35587);
xor U36888 (N_36888,N_35529,N_35324);
and U36889 (N_36889,N_35741,N_35391);
or U36890 (N_36890,N_35190,N_35444);
and U36891 (N_36891,N_35023,N_35160);
or U36892 (N_36892,N_35908,N_35514);
nand U36893 (N_36893,N_35432,N_35085);
xnor U36894 (N_36894,N_35246,N_35961);
and U36895 (N_36895,N_35429,N_35542);
or U36896 (N_36896,N_35106,N_35450);
and U36897 (N_36897,N_35616,N_35285);
or U36898 (N_36898,N_35225,N_35839);
xnor U36899 (N_36899,N_35894,N_35736);
nor U36900 (N_36900,N_35510,N_35586);
or U36901 (N_36901,N_35384,N_35982);
and U36902 (N_36902,N_35369,N_35694);
nand U36903 (N_36903,N_35016,N_35491);
nand U36904 (N_36904,N_35989,N_35456);
nor U36905 (N_36905,N_35837,N_35059);
and U36906 (N_36906,N_35525,N_35747);
xnor U36907 (N_36907,N_35703,N_35022);
xor U36908 (N_36908,N_35624,N_35742);
nand U36909 (N_36909,N_35508,N_35952);
xor U36910 (N_36910,N_35240,N_35875);
or U36911 (N_36911,N_35371,N_35316);
and U36912 (N_36912,N_35481,N_35471);
and U36913 (N_36913,N_35609,N_35877);
nand U36914 (N_36914,N_35216,N_35332);
xor U36915 (N_36915,N_35268,N_35454);
nor U36916 (N_36916,N_35226,N_35010);
xor U36917 (N_36917,N_35456,N_35489);
and U36918 (N_36918,N_35113,N_35312);
or U36919 (N_36919,N_35326,N_35859);
nand U36920 (N_36920,N_35590,N_35822);
nor U36921 (N_36921,N_35854,N_35390);
and U36922 (N_36922,N_35918,N_35079);
and U36923 (N_36923,N_35239,N_35393);
xnor U36924 (N_36924,N_35014,N_35776);
nor U36925 (N_36925,N_35701,N_35411);
nand U36926 (N_36926,N_35372,N_35022);
xor U36927 (N_36927,N_35967,N_35182);
nand U36928 (N_36928,N_35613,N_35764);
xor U36929 (N_36929,N_35963,N_35526);
or U36930 (N_36930,N_35220,N_35120);
nand U36931 (N_36931,N_35019,N_35230);
xnor U36932 (N_36932,N_35377,N_35532);
or U36933 (N_36933,N_35035,N_35858);
xor U36934 (N_36934,N_35907,N_35168);
nand U36935 (N_36935,N_35458,N_35363);
and U36936 (N_36936,N_35764,N_35993);
and U36937 (N_36937,N_35227,N_35622);
or U36938 (N_36938,N_35500,N_35990);
nand U36939 (N_36939,N_35337,N_35299);
or U36940 (N_36940,N_35262,N_35342);
nor U36941 (N_36941,N_35997,N_35911);
and U36942 (N_36942,N_35882,N_35608);
nand U36943 (N_36943,N_35075,N_35946);
or U36944 (N_36944,N_35811,N_35260);
xnor U36945 (N_36945,N_35576,N_35818);
nor U36946 (N_36946,N_35585,N_35789);
nand U36947 (N_36947,N_35434,N_35426);
or U36948 (N_36948,N_35972,N_35704);
and U36949 (N_36949,N_35696,N_35897);
and U36950 (N_36950,N_35425,N_35269);
nor U36951 (N_36951,N_35090,N_35397);
xnor U36952 (N_36952,N_35431,N_35061);
and U36953 (N_36953,N_35557,N_35472);
or U36954 (N_36954,N_35761,N_35904);
nand U36955 (N_36955,N_35671,N_35669);
xor U36956 (N_36956,N_35040,N_35544);
xnor U36957 (N_36957,N_35005,N_35055);
or U36958 (N_36958,N_35443,N_35506);
nand U36959 (N_36959,N_35393,N_35438);
or U36960 (N_36960,N_35057,N_35403);
nor U36961 (N_36961,N_35588,N_35366);
or U36962 (N_36962,N_35011,N_35197);
and U36963 (N_36963,N_35417,N_35008);
or U36964 (N_36964,N_35907,N_35944);
nor U36965 (N_36965,N_35739,N_35665);
xnor U36966 (N_36966,N_35308,N_35455);
or U36967 (N_36967,N_35061,N_35573);
nand U36968 (N_36968,N_35583,N_35982);
xnor U36969 (N_36969,N_35644,N_35992);
nand U36970 (N_36970,N_35581,N_35071);
nand U36971 (N_36971,N_35977,N_35005);
or U36972 (N_36972,N_35322,N_35018);
or U36973 (N_36973,N_35047,N_35255);
nand U36974 (N_36974,N_35462,N_35188);
or U36975 (N_36975,N_35472,N_35834);
or U36976 (N_36976,N_35611,N_35782);
xor U36977 (N_36977,N_35345,N_35236);
and U36978 (N_36978,N_35380,N_35955);
and U36979 (N_36979,N_35204,N_35825);
xnor U36980 (N_36980,N_35215,N_35629);
xnor U36981 (N_36981,N_35266,N_35213);
or U36982 (N_36982,N_35470,N_35300);
or U36983 (N_36983,N_35169,N_35213);
nand U36984 (N_36984,N_35441,N_35819);
or U36985 (N_36985,N_35740,N_35697);
nor U36986 (N_36986,N_35249,N_35503);
nand U36987 (N_36987,N_35835,N_35206);
nand U36988 (N_36988,N_35510,N_35892);
nand U36989 (N_36989,N_35523,N_35123);
or U36990 (N_36990,N_35490,N_35311);
and U36991 (N_36991,N_35750,N_35157);
nor U36992 (N_36992,N_35318,N_35627);
nand U36993 (N_36993,N_35077,N_35291);
or U36994 (N_36994,N_35301,N_35257);
nand U36995 (N_36995,N_35504,N_35852);
nand U36996 (N_36996,N_35955,N_35097);
or U36997 (N_36997,N_35899,N_35456);
and U36998 (N_36998,N_35863,N_35027);
nand U36999 (N_36999,N_35382,N_35689);
nand U37000 (N_37000,N_36842,N_36069);
or U37001 (N_37001,N_36327,N_36345);
xor U37002 (N_37002,N_36170,N_36473);
nor U37003 (N_37003,N_36831,N_36340);
nand U37004 (N_37004,N_36962,N_36822);
or U37005 (N_37005,N_36821,N_36852);
nand U37006 (N_37006,N_36702,N_36902);
nor U37007 (N_37007,N_36577,N_36164);
and U37008 (N_37008,N_36974,N_36736);
and U37009 (N_37009,N_36518,N_36669);
nor U37010 (N_37010,N_36712,N_36717);
xor U37011 (N_37011,N_36427,N_36064);
and U37012 (N_37012,N_36253,N_36217);
or U37013 (N_37013,N_36344,N_36651);
or U37014 (N_37014,N_36222,N_36351);
or U37015 (N_37015,N_36237,N_36142);
xnor U37016 (N_37016,N_36050,N_36215);
xor U37017 (N_37017,N_36868,N_36529);
xor U37018 (N_37018,N_36662,N_36203);
or U37019 (N_37019,N_36022,N_36711);
and U37020 (N_37020,N_36040,N_36490);
xor U37021 (N_37021,N_36795,N_36915);
nor U37022 (N_37022,N_36090,N_36864);
and U37023 (N_37023,N_36007,N_36005);
and U37024 (N_37024,N_36656,N_36113);
or U37025 (N_37025,N_36003,N_36184);
or U37026 (N_37026,N_36636,N_36401);
or U37027 (N_37027,N_36104,N_36804);
nand U37028 (N_37028,N_36983,N_36212);
nor U37029 (N_37029,N_36209,N_36716);
nand U37030 (N_37030,N_36840,N_36861);
nor U37031 (N_37031,N_36749,N_36377);
xor U37032 (N_37032,N_36457,N_36423);
or U37033 (N_37033,N_36533,N_36476);
or U37034 (N_37034,N_36694,N_36833);
xor U37035 (N_37035,N_36337,N_36798);
nand U37036 (N_37036,N_36495,N_36396);
or U37037 (N_37037,N_36670,N_36838);
and U37038 (N_37038,N_36775,N_36191);
and U37039 (N_37039,N_36443,N_36665);
xnor U37040 (N_37040,N_36470,N_36044);
nor U37041 (N_37041,N_36683,N_36031);
nand U37042 (N_37042,N_36455,N_36135);
or U37043 (N_37043,N_36324,N_36865);
nor U37044 (N_37044,N_36467,N_36579);
nand U37045 (N_37045,N_36674,N_36765);
and U37046 (N_37046,N_36549,N_36823);
xnor U37047 (N_37047,N_36952,N_36048);
xnor U37048 (N_37048,N_36611,N_36060);
nand U37049 (N_37049,N_36723,N_36091);
xnor U37050 (N_37050,N_36872,N_36413);
nand U37051 (N_37051,N_36746,N_36496);
xor U37052 (N_37052,N_36273,N_36353);
and U37053 (N_37053,N_36517,N_36737);
and U37054 (N_37054,N_36834,N_36985);
nand U37055 (N_37055,N_36507,N_36828);
and U37056 (N_37056,N_36678,N_36130);
xnor U37057 (N_37057,N_36475,N_36978);
xor U37058 (N_37058,N_36829,N_36163);
nor U37059 (N_37059,N_36082,N_36332);
xnor U37060 (N_37060,N_36235,N_36479);
xor U37061 (N_37061,N_36891,N_36311);
and U37062 (N_37062,N_36863,N_36627);
and U37063 (N_37063,N_36274,N_36036);
nor U37064 (N_37064,N_36922,N_36446);
and U37065 (N_37065,N_36889,N_36799);
nand U37066 (N_37066,N_36792,N_36227);
and U37067 (N_37067,N_36596,N_36238);
and U37068 (N_37068,N_36807,N_36508);
or U37069 (N_37069,N_36866,N_36271);
xnor U37070 (N_37070,N_36001,N_36563);
and U37071 (N_37071,N_36472,N_36751);
nor U37072 (N_37072,N_36830,N_36367);
nor U37073 (N_37073,N_36127,N_36638);
xnor U37074 (N_37074,N_36888,N_36439);
or U37075 (N_37075,N_36643,N_36188);
nand U37076 (N_37076,N_36703,N_36767);
or U37077 (N_37077,N_36996,N_36339);
or U37078 (N_37078,N_36027,N_36748);
and U37079 (N_37079,N_36881,N_36484);
and U37080 (N_37080,N_36705,N_36286);
xnor U37081 (N_37081,N_36161,N_36464);
xnor U37082 (N_37082,N_36081,N_36644);
or U37083 (N_37083,N_36741,N_36254);
nor U37084 (N_37084,N_36975,N_36486);
and U37085 (N_37085,N_36305,N_36310);
nor U37086 (N_37086,N_36350,N_36174);
nand U37087 (N_37087,N_36160,N_36885);
nor U37088 (N_37088,N_36120,N_36420);
nand U37089 (N_37089,N_36898,N_36900);
nand U37090 (N_37090,N_36440,N_36946);
nor U37091 (N_37091,N_36673,N_36870);
or U37092 (N_37092,N_36941,N_36086);
nor U37093 (N_37093,N_36619,N_36356);
and U37094 (N_37094,N_36832,N_36213);
or U37095 (N_37095,N_36782,N_36522);
and U37096 (N_37096,N_36541,N_36732);
nand U37097 (N_37097,N_36270,N_36148);
and U37098 (N_37098,N_36956,N_36502);
nor U37099 (N_37099,N_36854,N_36528);
nand U37100 (N_37100,N_36580,N_36818);
xnor U37101 (N_37101,N_36550,N_36575);
nor U37102 (N_37102,N_36002,N_36250);
or U37103 (N_37103,N_36330,N_36848);
or U37104 (N_37104,N_36505,N_36412);
or U37105 (N_37105,N_36282,N_36061);
or U37106 (N_37106,N_36591,N_36616);
and U37107 (N_37107,N_36093,N_36945);
xor U37108 (N_37108,N_36520,N_36309);
nand U37109 (N_37109,N_36368,N_36721);
xnor U37110 (N_37110,N_36570,N_36333);
xor U37111 (N_37111,N_36547,N_36536);
or U37112 (N_37112,N_36882,N_36199);
or U37113 (N_37113,N_36021,N_36903);
nand U37114 (N_37114,N_36229,N_36109);
or U37115 (N_37115,N_36033,N_36145);
xor U37116 (N_37116,N_36291,N_36790);
nor U37117 (N_37117,N_36038,N_36498);
nand U37118 (N_37118,N_36598,N_36998);
nor U37119 (N_37119,N_36453,N_36430);
nor U37120 (N_37120,N_36346,N_36910);
and U37121 (N_37121,N_36450,N_36449);
nand U37122 (N_37122,N_36202,N_36483);
and U37123 (N_37123,N_36304,N_36460);
and U37124 (N_37124,N_36223,N_36672);
xnor U37125 (N_37125,N_36789,N_36970);
and U37126 (N_37126,N_36133,N_36421);
or U37127 (N_37127,N_36482,N_36690);
xnor U37128 (N_37128,N_36940,N_36796);
xnor U37129 (N_37129,N_36108,N_36512);
and U37130 (N_37130,N_36728,N_36500);
nand U37131 (N_37131,N_36935,N_36675);
nand U37132 (N_37132,N_36451,N_36255);
nor U37133 (N_37133,N_36784,N_36811);
nand U37134 (N_37134,N_36844,N_36463);
and U37135 (N_37135,N_36402,N_36609);
nand U37136 (N_37136,N_36648,N_36562);
and U37137 (N_37137,N_36560,N_36165);
or U37138 (N_37138,N_36637,N_36664);
nand U37139 (N_37139,N_36601,N_36835);
xor U37140 (N_37140,N_36141,N_36953);
xor U37141 (N_37141,N_36752,N_36603);
or U37142 (N_37142,N_36817,N_36147);
xnor U37143 (N_37143,N_36297,N_36851);
nand U37144 (N_37144,N_36681,N_36907);
xnor U37145 (N_37145,N_36599,N_36041);
and U37146 (N_37146,N_36265,N_36565);
nand U37147 (N_37147,N_36629,N_36369);
nand U37148 (N_37148,N_36454,N_36808);
nand U37149 (N_37149,N_36076,N_36408);
nor U37150 (N_37150,N_36667,N_36319);
nor U37151 (N_37151,N_36836,N_36251);
or U37152 (N_37152,N_36106,N_36269);
or U37153 (N_37153,N_36196,N_36745);
nand U37154 (N_37154,N_36029,N_36267);
or U37155 (N_37155,N_36383,N_36151);
xnor U37156 (N_37156,N_36358,N_36252);
xor U37157 (N_37157,N_36666,N_36663);
or U37158 (N_37158,N_36862,N_36359);
and U37159 (N_37159,N_36491,N_36175);
or U37160 (N_37160,N_36198,N_36458);
or U37161 (N_37161,N_36306,N_36967);
nor U37162 (N_37162,N_36645,N_36559);
or U37163 (N_37163,N_36492,N_36760);
xnor U37164 (N_37164,N_36375,N_36824);
xnor U37165 (N_37165,N_36249,N_36065);
or U37166 (N_37166,N_36682,N_36901);
or U37167 (N_37167,N_36162,N_36288);
and U37168 (N_37168,N_36438,N_36510);
or U37169 (N_37169,N_36926,N_36139);
or U37170 (N_37170,N_36999,N_36099);
and U37171 (N_37171,N_36660,N_36553);
nand U37172 (N_37172,N_36374,N_36893);
nor U37173 (N_37173,N_36986,N_36769);
or U37174 (N_37174,N_36006,N_36246);
nor U37175 (N_37175,N_36268,N_36341);
xor U37176 (N_37176,N_36382,N_36039);
or U37177 (N_37177,N_36921,N_36624);
xor U37178 (N_37178,N_36294,N_36261);
nor U37179 (N_37179,N_36258,N_36630);
nor U37180 (N_37180,N_36317,N_36011);
and U37181 (N_37181,N_36315,N_36372);
nor U37182 (N_37182,N_36461,N_36462);
nor U37183 (N_37183,N_36015,N_36720);
and U37184 (N_37184,N_36523,N_36552);
xor U37185 (N_37185,N_36302,N_36904);
nor U37186 (N_37186,N_36853,N_36688);
nor U37187 (N_37187,N_36614,N_36590);
xnor U37188 (N_37188,N_36931,N_36689);
nand U37189 (N_37189,N_36623,N_36275);
nand U37190 (N_37190,N_36328,N_36392);
nor U37191 (N_37191,N_36966,N_36806);
nand U37192 (N_37192,N_36617,N_36704);
nor U37193 (N_37193,N_36588,N_36247);
xnor U37194 (N_37194,N_36386,N_36049);
or U37195 (N_37195,N_36477,N_36587);
nor U37196 (N_37196,N_36696,N_36894);
xor U37197 (N_37197,N_36322,N_36905);
and U37198 (N_37198,N_36149,N_36024);
nor U37199 (N_37199,N_36739,N_36063);
xnor U37200 (N_37200,N_36859,N_36092);
and U37201 (N_37201,N_36805,N_36260);
and U37202 (N_37202,N_36032,N_36187);
and U37203 (N_37203,N_36243,N_36542);
nand U37204 (N_37204,N_36084,N_36146);
xnor U37205 (N_37205,N_36384,N_36583);
xnor U37206 (N_37206,N_36216,N_36228);
and U37207 (N_37207,N_36296,N_36390);
or U37208 (N_37208,N_36586,N_36958);
nor U37209 (N_37209,N_36173,N_36925);
xor U37210 (N_37210,N_36794,N_36558);
or U37211 (N_37211,N_36571,N_36157);
xor U37212 (N_37212,N_36432,N_36534);
nand U37213 (N_37213,N_36131,N_36548);
and U37214 (N_37214,N_36772,N_36348);
xnor U37215 (N_37215,N_36544,N_36232);
xor U37216 (N_37216,N_36025,N_36691);
or U37217 (N_37217,N_36070,N_36773);
and U37218 (N_37218,N_36963,N_36428);
nand U37219 (N_37219,N_36699,N_36088);
nor U37220 (N_37220,N_36679,N_36594);
nor U37221 (N_37221,N_36774,N_36761);
and U37222 (N_37222,N_36763,N_36887);
xor U37223 (N_37223,N_36431,N_36973);
nor U37224 (N_37224,N_36207,N_36400);
and U37225 (N_37225,N_36004,N_36787);
xnor U37226 (N_37226,N_36730,N_36743);
xor U37227 (N_37227,N_36422,N_36159);
and U37228 (N_37228,N_36468,N_36290);
nand U37229 (N_37229,N_36493,N_36494);
and U37230 (N_37230,N_36551,N_36981);
or U37231 (N_37231,N_36018,N_36204);
nand U37232 (N_37232,N_36334,N_36564);
or U37233 (N_37233,N_36930,N_36554);
nor U37234 (N_37234,N_36785,N_36233);
nand U37235 (N_37235,N_36715,N_36442);
nor U37236 (N_37236,N_36697,N_36182);
or U37237 (N_37237,N_36530,N_36110);
nand U37238 (N_37238,N_36079,N_36726);
xor U37239 (N_37239,N_36964,N_36574);
nand U37240 (N_37240,N_36465,N_36722);
or U37241 (N_37241,N_36404,N_36869);
nor U37242 (N_37242,N_36074,N_36205);
and U37243 (N_37243,N_36719,N_36000);
xor U37244 (N_37244,N_36521,N_36325);
xor U37245 (N_37245,N_36653,N_36155);
xor U37246 (N_37246,N_36718,N_36391);
and U37247 (N_37247,N_36220,N_36071);
or U37248 (N_37248,N_36698,N_36613);
or U37249 (N_37249,N_36389,N_36168);
and U37250 (N_37250,N_36123,N_36119);
nor U37251 (N_37251,N_36117,N_36841);
and U37252 (N_37252,N_36747,N_36181);
nand U37253 (N_37253,N_36009,N_36993);
xor U37254 (N_37254,N_36932,N_36912);
nand U37255 (N_37255,N_36067,N_36097);
nor U37256 (N_37256,N_36979,N_36410);
xnor U37257 (N_37257,N_36729,N_36416);
xnor U37258 (N_37258,N_36292,N_36708);
nand U37259 (N_37259,N_36783,N_36171);
xor U37260 (N_37260,N_36307,N_36019);
nor U37261 (N_37261,N_36028,N_36179);
or U37262 (N_37262,N_36756,N_36951);
nand U37263 (N_37263,N_36053,N_36045);
and U37264 (N_37264,N_36801,N_36687);
and U37265 (N_37265,N_36409,N_36183);
or U37266 (N_37266,N_36511,N_36733);
nor U37267 (N_37267,N_36231,N_36085);
nor U37268 (N_37268,N_36892,N_36437);
nand U37269 (N_37269,N_36879,N_36519);
nor U37270 (N_37270,N_36913,N_36128);
or U37271 (N_37271,N_36621,N_36362);
xnor U37272 (N_37272,N_36489,N_36239);
nand U37273 (N_37273,N_36814,N_36649);
nand U37274 (N_37274,N_36444,N_36397);
or U37275 (N_37275,N_36526,N_36293);
or U37276 (N_37276,N_36289,N_36059);
and U37277 (N_37277,N_36210,N_36827);
and U37278 (N_37278,N_36928,N_36035);
nor U37279 (N_37279,N_36277,N_36661);
and U37280 (N_37280,N_36156,N_36855);
or U37281 (N_37281,N_36096,N_36103);
nand U37282 (N_37282,N_36837,N_36977);
nor U37283 (N_37283,N_36057,N_36676);
or U37284 (N_37284,N_36378,N_36077);
xnor U37285 (N_37285,N_36635,N_36965);
nand U37286 (N_37286,N_36016,N_36435);
and U37287 (N_37287,N_36424,N_36014);
or U37288 (N_37288,N_36724,N_36323);
nor U37289 (N_37289,N_36899,N_36102);
and U37290 (N_37290,N_36895,N_36628);
xor U37291 (N_37291,N_36398,N_36411);
xor U37292 (N_37292,N_36008,N_36136);
xnor U37293 (N_37293,N_36370,N_36366);
nor U37294 (N_37294,N_36256,N_36602);
and U37295 (N_37295,N_36488,N_36919);
nor U37296 (N_37296,N_36121,N_36820);
or U37297 (N_37297,N_36927,N_36939);
or U37298 (N_37298,N_36154,N_36620);
and U37299 (N_37299,N_36797,N_36581);
or U37300 (N_37300,N_36062,N_36725);
xnor U37301 (N_37301,N_36447,N_36757);
nand U37302 (N_37302,N_36226,N_36567);
or U37303 (N_37303,N_36278,N_36608);
nand U37304 (N_37304,N_36871,N_36364);
or U37305 (N_37305,N_36285,N_36877);
and U37306 (N_37306,N_36755,N_36849);
or U37307 (N_37307,N_36349,N_36639);
nor U37308 (N_37308,N_36095,N_36321);
and U37309 (N_37309,N_36569,N_36407);
or U37310 (N_37310,N_36178,N_36284);
xnor U37311 (N_37311,N_36192,N_36101);
nor U37312 (N_37312,N_36230,N_36994);
nand U37313 (N_37313,N_36744,N_36122);
or U37314 (N_37314,N_36556,N_36094);
xor U37315 (N_37315,N_36497,N_36194);
nand U37316 (N_37316,N_36873,N_36361);
or U37317 (N_37317,N_36954,N_36320);
xor U37318 (N_37318,N_36190,N_36221);
or U37319 (N_37319,N_36373,N_36381);
and U37320 (N_37320,N_36023,N_36026);
nand U37321 (N_37321,N_36335,N_36343);
nand U37322 (N_37322,N_36896,N_36176);
or U37323 (N_37323,N_36112,N_36684);
or U37324 (N_37324,N_36758,N_36316);
xor U37325 (N_37325,N_36355,N_36659);
nor U37326 (N_37326,N_36118,N_36078);
nor U37327 (N_37327,N_36802,N_36186);
nand U37328 (N_37328,N_36537,N_36707);
and U37329 (N_37329,N_36020,N_36527);
xnor U37330 (N_37330,N_36933,N_36539);
nor U37331 (N_37331,N_36425,N_36605);
nand U37332 (N_37332,N_36989,N_36860);
and U37333 (N_37333,N_36515,N_36546);
or U37334 (N_37334,N_36770,N_36701);
nand U37335 (N_37335,N_36780,N_36525);
and U37336 (N_37336,N_36754,N_36607);
nor U37337 (N_37337,N_36318,N_36778);
xnor U37338 (N_37338,N_36481,N_36813);
nand U37339 (N_37339,N_36363,N_36480);
nand U37340 (N_37340,N_36949,N_36441);
nand U37341 (N_37341,N_36365,N_36279);
and U37342 (N_37342,N_36692,N_36326);
and U37343 (N_37343,N_36485,N_36272);
nor U37344 (N_37344,N_36582,N_36615);
xor U37345 (N_37345,N_36555,N_36781);
xnor U37346 (N_37346,N_36566,N_36972);
and U37347 (N_37347,N_36080,N_36906);
and U37348 (N_37348,N_36166,N_36917);
nor U37349 (N_37349,N_36961,N_36734);
xor U37350 (N_37350,N_36943,N_36169);
xor U37351 (N_37351,N_36300,N_36301);
nand U37352 (N_37352,N_36677,N_36845);
and U37353 (N_37353,N_36405,N_36944);
or U37354 (N_37354,N_36955,N_36777);
or U37355 (N_37355,N_36589,N_36631);
nand U37356 (N_37356,N_36089,N_36538);
and U37357 (N_37357,N_36995,N_36650);
and U37358 (N_37358,N_36395,N_36948);
and U37359 (N_37359,N_36980,N_36680);
nor U37360 (N_37360,N_36686,N_36695);
and U37361 (N_37361,N_36087,N_36634);
and U37362 (N_37362,N_36017,N_36585);
xor U37363 (N_37363,N_36991,N_36456);
and U37364 (N_37364,N_36762,N_36144);
nor U37365 (N_37365,N_36809,N_36387);
or U37366 (N_37366,N_36371,N_36241);
and U37367 (N_37367,N_36997,N_36668);
nand U37368 (N_37368,N_36779,N_36208);
xor U37369 (N_37369,N_36240,N_36800);
xnor U37370 (N_37370,N_36655,N_36911);
xnor U37371 (N_37371,N_36576,N_36657);
or U37372 (N_37372,N_36143,N_36641);
and U37373 (N_37373,N_36013,N_36478);
and U37374 (N_37374,N_36815,N_36503);
or U37375 (N_37375,N_36936,N_36742);
or U37376 (N_37376,N_36499,N_36846);
nand U37377 (N_37377,N_36047,N_36988);
or U37378 (N_37378,N_36360,N_36839);
and U37379 (N_37379,N_36600,N_36058);
xor U37380 (N_37380,N_36283,N_36399);
and U37381 (N_37381,N_36776,N_36257);
or U37382 (N_37382,N_36597,N_36987);
nor U37383 (N_37383,N_36934,N_36509);
or U37384 (N_37384,N_36380,N_36066);
and U37385 (N_37385,N_36394,N_36206);
or U37386 (N_37386,N_36137,N_36393);
nand U37387 (N_37387,N_36052,N_36714);
xnor U37388 (N_37388,N_36415,N_36593);
nor U37389 (N_37389,N_36874,N_36129);
or U37390 (N_37390,N_36298,N_36030);
and U37391 (N_37391,N_36347,N_36125);
and U37392 (N_37392,N_36916,N_36299);
xor U37393 (N_37393,N_36654,N_36376);
and U37394 (N_37394,N_36584,N_36242);
or U37395 (N_37395,N_36234,N_36622);
nor U37396 (N_37396,N_36731,N_36403);
and U37397 (N_37397,N_36068,N_36924);
nor U37398 (N_37398,N_36418,N_36201);
nor U37399 (N_37399,N_36342,N_36764);
xor U37400 (N_37400,N_36766,N_36858);
and U37401 (N_37401,N_36098,N_36646);
nand U37402 (N_37402,N_36693,N_36920);
xnor U37403 (N_37403,N_36513,N_36075);
nor U37404 (N_37404,N_36211,N_36969);
nor U37405 (N_37405,N_36264,N_36786);
xor U37406 (N_37406,N_36942,N_36524);
and U37407 (N_37407,N_36557,N_36990);
nand U37408 (N_37408,N_36385,N_36950);
and U37409 (N_37409,N_36132,N_36843);
nor U37410 (N_37410,N_36713,N_36436);
and U37411 (N_37411,N_36706,N_36469);
nor U37412 (N_37412,N_36647,N_36959);
nor U37413 (N_37413,N_36504,N_36561);
and U37414 (N_37414,N_36610,N_36727);
xor U37415 (N_37415,N_36632,N_36735);
nor U37416 (N_37416,N_36312,N_36768);
and U37417 (N_37417,N_36897,N_36012);
nor U37418 (N_37418,N_36073,N_36700);
xor U37419 (N_37419,N_36115,N_36434);
and U37420 (N_37420,N_36189,N_36452);
or U37421 (N_37421,N_36338,N_36788);
nor U37422 (N_37422,N_36506,N_36466);
nor U37423 (N_37423,N_36612,N_36540);
nor U37424 (N_37424,N_36158,N_36816);
nor U37425 (N_37425,N_36592,N_36248);
xor U37426 (N_37426,N_36197,N_36875);
nand U37427 (N_37427,N_36532,N_36709);
and U37428 (N_37428,N_36034,N_36037);
xnor U37429 (N_37429,N_36010,N_36051);
nand U37430 (N_37430,N_36193,N_36357);
or U37431 (N_37431,N_36336,N_36314);
nand U37432 (N_37432,N_36329,N_36124);
xnor U37433 (N_37433,N_36918,N_36826);
and U37434 (N_37434,N_36114,N_36793);
or U37435 (N_37435,N_36545,N_36295);
and U37436 (N_37436,N_36100,N_36971);
xnor U37437 (N_37437,N_36474,N_36263);
nand U37438 (N_37438,N_36625,N_36054);
or U37439 (N_37439,N_36957,N_36352);
xnor U37440 (N_37440,N_36150,N_36225);
nor U37441 (N_37441,N_36406,N_36262);
nand U37442 (N_37442,N_36459,N_36046);
and U37443 (N_37443,N_36429,N_36448);
or U37444 (N_37444,N_36890,N_36652);
nor U37445 (N_37445,N_36633,N_36111);
nor U37446 (N_37446,N_36172,N_36604);
nand U37447 (N_37447,N_36671,N_36259);
or U37448 (N_37448,N_36245,N_36759);
xor U37449 (N_37449,N_36984,N_36880);
nand U37450 (N_37450,N_36908,N_36883);
or U37451 (N_37451,N_36738,N_36976);
or U37452 (N_37452,N_36218,N_36938);
nand U37453 (N_37453,N_36923,N_36244);
nor U37454 (N_37454,N_36578,N_36471);
nand U37455 (N_37455,N_36857,N_36419);
or U37456 (N_37456,N_36572,N_36710);
or U37457 (N_37457,N_36153,N_36685);
nand U37458 (N_37458,N_36043,N_36200);
or U37459 (N_37459,N_36803,N_36992);
or U37460 (N_37460,N_36847,N_36947);
nor U37461 (N_37461,N_36167,N_36126);
xnor U37462 (N_37462,N_36266,N_36276);
xnor U37463 (N_37463,N_36968,N_36740);
or U37464 (N_37464,N_36152,N_36812);
or U37465 (N_37465,N_36568,N_36195);
nand U37466 (N_37466,N_36313,N_36884);
and U37467 (N_37467,N_36929,N_36287);
or U37468 (N_37468,N_36642,N_36626);
nand U37469 (N_37469,N_36595,N_36281);
xor U37470 (N_37470,N_36876,N_36771);
nand U37471 (N_37471,N_36856,N_36914);
or U37472 (N_37472,N_36867,N_36219);
and U37473 (N_37473,N_36055,N_36280);
nor U37474 (N_37474,N_36083,N_36878);
or U37475 (N_37475,N_36982,N_36487);
nor U37476 (N_37476,N_36354,N_36514);
nor U37477 (N_37477,N_36543,N_36331);
and U37478 (N_37478,N_36303,N_36531);
xnor U37479 (N_37479,N_36214,N_36606);
and U37480 (N_37480,N_36618,N_36414);
and U37481 (N_37481,N_36417,N_36433);
xor U37482 (N_37482,N_36224,N_36105);
and U37483 (N_37483,N_36180,N_36850);
nand U37484 (N_37484,N_36810,N_36825);
nand U37485 (N_37485,N_36134,N_36573);
and U37486 (N_37486,N_36308,N_36445);
nor U37487 (N_37487,N_36116,N_36909);
and U37488 (N_37488,N_36056,N_36236);
xnor U37489 (N_37489,N_36501,N_36426);
nand U37490 (N_37490,N_36750,N_36379);
or U37491 (N_37491,N_36140,N_36516);
nor U37492 (N_37492,N_36107,N_36042);
xnor U37493 (N_37493,N_36388,N_36791);
nor U37494 (N_37494,N_36177,N_36072);
nand U37495 (N_37495,N_36185,N_36960);
or U37496 (N_37496,N_36535,N_36138);
or U37497 (N_37497,N_36937,N_36886);
nand U37498 (N_37498,N_36640,N_36658);
xor U37499 (N_37499,N_36819,N_36753);
or U37500 (N_37500,N_36341,N_36594);
nand U37501 (N_37501,N_36042,N_36099);
nor U37502 (N_37502,N_36648,N_36559);
nor U37503 (N_37503,N_36372,N_36834);
and U37504 (N_37504,N_36642,N_36481);
xnor U37505 (N_37505,N_36972,N_36051);
and U37506 (N_37506,N_36485,N_36654);
and U37507 (N_37507,N_36916,N_36364);
nor U37508 (N_37508,N_36123,N_36695);
or U37509 (N_37509,N_36202,N_36236);
and U37510 (N_37510,N_36760,N_36906);
and U37511 (N_37511,N_36184,N_36141);
xor U37512 (N_37512,N_36795,N_36188);
and U37513 (N_37513,N_36309,N_36515);
nand U37514 (N_37514,N_36453,N_36954);
and U37515 (N_37515,N_36330,N_36416);
and U37516 (N_37516,N_36394,N_36296);
or U37517 (N_37517,N_36860,N_36785);
nor U37518 (N_37518,N_36890,N_36817);
xor U37519 (N_37519,N_36255,N_36699);
xor U37520 (N_37520,N_36955,N_36362);
or U37521 (N_37521,N_36671,N_36909);
or U37522 (N_37522,N_36370,N_36110);
nand U37523 (N_37523,N_36821,N_36061);
xnor U37524 (N_37524,N_36887,N_36631);
xor U37525 (N_37525,N_36826,N_36751);
nand U37526 (N_37526,N_36015,N_36517);
nor U37527 (N_37527,N_36747,N_36686);
or U37528 (N_37528,N_36578,N_36634);
nor U37529 (N_37529,N_36672,N_36399);
nor U37530 (N_37530,N_36142,N_36999);
or U37531 (N_37531,N_36630,N_36680);
and U37532 (N_37532,N_36073,N_36983);
nor U37533 (N_37533,N_36988,N_36050);
or U37534 (N_37534,N_36425,N_36061);
nor U37535 (N_37535,N_36039,N_36545);
nor U37536 (N_37536,N_36070,N_36108);
xor U37537 (N_37537,N_36833,N_36347);
and U37538 (N_37538,N_36537,N_36904);
or U37539 (N_37539,N_36606,N_36429);
xor U37540 (N_37540,N_36459,N_36947);
or U37541 (N_37541,N_36225,N_36411);
xnor U37542 (N_37542,N_36164,N_36229);
nor U37543 (N_37543,N_36455,N_36670);
xor U37544 (N_37544,N_36560,N_36963);
or U37545 (N_37545,N_36185,N_36914);
xor U37546 (N_37546,N_36238,N_36860);
nand U37547 (N_37547,N_36479,N_36386);
nand U37548 (N_37548,N_36087,N_36261);
and U37549 (N_37549,N_36310,N_36068);
nand U37550 (N_37550,N_36516,N_36098);
nor U37551 (N_37551,N_36215,N_36473);
nor U37552 (N_37552,N_36166,N_36765);
nor U37553 (N_37553,N_36595,N_36258);
xor U37554 (N_37554,N_36590,N_36626);
or U37555 (N_37555,N_36797,N_36147);
or U37556 (N_37556,N_36654,N_36620);
nor U37557 (N_37557,N_36429,N_36072);
and U37558 (N_37558,N_36883,N_36968);
xnor U37559 (N_37559,N_36562,N_36287);
xnor U37560 (N_37560,N_36412,N_36619);
nor U37561 (N_37561,N_36476,N_36779);
nor U37562 (N_37562,N_36034,N_36556);
and U37563 (N_37563,N_36458,N_36419);
nand U37564 (N_37564,N_36320,N_36975);
xor U37565 (N_37565,N_36625,N_36856);
nand U37566 (N_37566,N_36416,N_36275);
or U37567 (N_37567,N_36580,N_36023);
nand U37568 (N_37568,N_36078,N_36563);
nand U37569 (N_37569,N_36276,N_36698);
nand U37570 (N_37570,N_36626,N_36120);
and U37571 (N_37571,N_36663,N_36880);
and U37572 (N_37572,N_36439,N_36660);
nand U37573 (N_37573,N_36603,N_36560);
and U37574 (N_37574,N_36352,N_36319);
xor U37575 (N_37575,N_36654,N_36940);
and U37576 (N_37576,N_36580,N_36508);
and U37577 (N_37577,N_36298,N_36018);
nor U37578 (N_37578,N_36733,N_36404);
or U37579 (N_37579,N_36316,N_36806);
and U37580 (N_37580,N_36092,N_36231);
nor U37581 (N_37581,N_36504,N_36575);
or U37582 (N_37582,N_36907,N_36616);
and U37583 (N_37583,N_36125,N_36448);
or U37584 (N_37584,N_36619,N_36370);
or U37585 (N_37585,N_36695,N_36614);
xor U37586 (N_37586,N_36404,N_36373);
nand U37587 (N_37587,N_36390,N_36710);
or U37588 (N_37588,N_36048,N_36895);
or U37589 (N_37589,N_36943,N_36268);
xor U37590 (N_37590,N_36290,N_36659);
and U37591 (N_37591,N_36025,N_36804);
xor U37592 (N_37592,N_36327,N_36032);
xor U37593 (N_37593,N_36264,N_36643);
nor U37594 (N_37594,N_36741,N_36248);
and U37595 (N_37595,N_36109,N_36411);
and U37596 (N_37596,N_36364,N_36132);
nand U37597 (N_37597,N_36566,N_36871);
or U37598 (N_37598,N_36581,N_36276);
or U37599 (N_37599,N_36415,N_36679);
xnor U37600 (N_37600,N_36219,N_36518);
xor U37601 (N_37601,N_36188,N_36372);
nand U37602 (N_37602,N_36270,N_36687);
nand U37603 (N_37603,N_36201,N_36295);
xor U37604 (N_37604,N_36770,N_36577);
xnor U37605 (N_37605,N_36711,N_36671);
and U37606 (N_37606,N_36847,N_36007);
xnor U37607 (N_37607,N_36401,N_36487);
xor U37608 (N_37608,N_36891,N_36953);
nor U37609 (N_37609,N_36595,N_36421);
and U37610 (N_37610,N_36046,N_36418);
or U37611 (N_37611,N_36107,N_36893);
or U37612 (N_37612,N_36056,N_36658);
xor U37613 (N_37613,N_36023,N_36311);
xnor U37614 (N_37614,N_36296,N_36031);
nand U37615 (N_37615,N_36234,N_36322);
nor U37616 (N_37616,N_36826,N_36444);
or U37617 (N_37617,N_36282,N_36512);
or U37618 (N_37618,N_36136,N_36953);
xor U37619 (N_37619,N_36622,N_36023);
nand U37620 (N_37620,N_36188,N_36631);
nand U37621 (N_37621,N_36661,N_36525);
and U37622 (N_37622,N_36929,N_36930);
nor U37623 (N_37623,N_36980,N_36527);
nand U37624 (N_37624,N_36886,N_36985);
nor U37625 (N_37625,N_36893,N_36862);
nand U37626 (N_37626,N_36640,N_36651);
xor U37627 (N_37627,N_36195,N_36888);
xnor U37628 (N_37628,N_36415,N_36719);
nor U37629 (N_37629,N_36196,N_36728);
or U37630 (N_37630,N_36846,N_36311);
nand U37631 (N_37631,N_36994,N_36574);
or U37632 (N_37632,N_36470,N_36832);
and U37633 (N_37633,N_36891,N_36916);
xor U37634 (N_37634,N_36132,N_36366);
nor U37635 (N_37635,N_36405,N_36634);
xor U37636 (N_37636,N_36052,N_36899);
nand U37637 (N_37637,N_36999,N_36449);
nand U37638 (N_37638,N_36146,N_36225);
or U37639 (N_37639,N_36346,N_36848);
nand U37640 (N_37640,N_36502,N_36144);
nor U37641 (N_37641,N_36980,N_36993);
or U37642 (N_37642,N_36221,N_36970);
and U37643 (N_37643,N_36148,N_36980);
xnor U37644 (N_37644,N_36631,N_36149);
nor U37645 (N_37645,N_36725,N_36703);
xor U37646 (N_37646,N_36021,N_36101);
or U37647 (N_37647,N_36607,N_36271);
or U37648 (N_37648,N_36191,N_36631);
nor U37649 (N_37649,N_36979,N_36489);
nor U37650 (N_37650,N_36021,N_36946);
and U37651 (N_37651,N_36886,N_36507);
nor U37652 (N_37652,N_36506,N_36318);
or U37653 (N_37653,N_36071,N_36227);
xor U37654 (N_37654,N_36274,N_36908);
nand U37655 (N_37655,N_36077,N_36996);
xnor U37656 (N_37656,N_36371,N_36673);
xor U37657 (N_37657,N_36880,N_36782);
and U37658 (N_37658,N_36529,N_36598);
nand U37659 (N_37659,N_36110,N_36923);
nand U37660 (N_37660,N_36976,N_36151);
nand U37661 (N_37661,N_36020,N_36849);
xor U37662 (N_37662,N_36791,N_36796);
nand U37663 (N_37663,N_36918,N_36439);
xor U37664 (N_37664,N_36439,N_36881);
nand U37665 (N_37665,N_36553,N_36667);
nand U37666 (N_37666,N_36274,N_36023);
xnor U37667 (N_37667,N_36479,N_36616);
nand U37668 (N_37668,N_36921,N_36105);
xor U37669 (N_37669,N_36401,N_36904);
and U37670 (N_37670,N_36319,N_36014);
nor U37671 (N_37671,N_36435,N_36681);
nand U37672 (N_37672,N_36639,N_36124);
or U37673 (N_37673,N_36421,N_36682);
and U37674 (N_37674,N_36626,N_36188);
nor U37675 (N_37675,N_36100,N_36409);
and U37676 (N_37676,N_36206,N_36462);
or U37677 (N_37677,N_36540,N_36229);
nand U37678 (N_37678,N_36620,N_36818);
nor U37679 (N_37679,N_36973,N_36924);
nand U37680 (N_37680,N_36477,N_36656);
xnor U37681 (N_37681,N_36978,N_36571);
xor U37682 (N_37682,N_36680,N_36506);
nor U37683 (N_37683,N_36352,N_36269);
and U37684 (N_37684,N_36937,N_36391);
nor U37685 (N_37685,N_36412,N_36884);
or U37686 (N_37686,N_36561,N_36908);
and U37687 (N_37687,N_36534,N_36968);
or U37688 (N_37688,N_36916,N_36311);
nor U37689 (N_37689,N_36178,N_36535);
nor U37690 (N_37690,N_36388,N_36184);
or U37691 (N_37691,N_36935,N_36190);
xnor U37692 (N_37692,N_36749,N_36950);
nor U37693 (N_37693,N_36396,N_36082);
or U37694 (N_37694,N_36087,N_36811);
xnor U37695 (N_37695,N_36447,N_36248);
nand U37696 (N_37696,N_36732,N_36313);
or U37697 (N_37697,N_36562,N_36141);
or U37698 (N_37698,N_36336,N_36162);
and U37699 (N_37699,N_36014,N_36508);
or U37700 (N_37700,N_36284,N_36752);
nor U37701 (N_37701,N_36090,N_36681);
xor U37702 (N_37702,N_36566,N_36983);
xnor U37703 (N_37703,N_36255,N_36322);
and U37704 (N_37704,N_36277,N_36792);
nor U37705 (N_37705,N_36112,N_36601);
nor U37706 (N_37706,N_36178,N_36327);
nor U37707 (N_37707,N_36724,N_36532);
nor U37708 (N_37708,N_36906,N_36740);
and U37709 (N_37709,N_36529,N_36359);
nor U37710 (N_37710,N_36761,N_36545);
xor U37711 (N_37711,N_36864,N_36681);
and U37712 (N_37712,N_36866,N_36082);
xnor U37713 (N_37713,N_36331,N_36324);
nor U37714 (N_37714,N_36744,N_36241);
nand U37715 (N_37715,N_36006,N_36512);
or U37716 (N_37716,N_36780,N_36724);
nand U37717 (N_37717,N_36219,N_36057);
and U37718 (N_37718,N_36409,N_36104);
nor U37719 (N_37719,N_36949,N_36904);
xor U37720 (N_37720,N_36801,N_36718);
nand U37721 (N_37721,N_36008,N_36751);
nor U37722 (N_37722,N_36820,N_36125);
and U37723 (N_37723,N_36792,N_36647);
or U37724 (N_37724,N_36357,N_36075);
nor U37725 (N_37725,N_36949,N_36048);
and U37726 (N_37726,N_36626,N_36810);
or U37727 (N_37727,N_36667,N_36606);
and U37728 (N_37728,N_36168,N_36557);
and U37729 (N_37729,N_36536,N_36004);
xnor U37730 (N_37730,N_36095,N_36232);
and U37731 (N_37731,N_36746,N_36650);
xor U37732 (N_37732,N_36591,N_36282);
nor U37733 (N_37733,N_36562,N_36788);
and U37734 (N_37734,N_36732,N_36744);
nand U37735 (N_37735,N_36570,N_36838);
xor U37736 (N_37736,N_36909,N_36576);
xor U37737 (N_37737,N_36655,N_36671);
nor U37738 (N_37738,N_36210,N_36688);
nand U37739 (N_37739,N_36953,N_36558);
nor U37740 (N_37740,N_36017,N_36460);
nand U37741 (N_37741,N_36596,N_36429);
nand U37742 (N_37742,N_36015,N_36513);
and U37743 (N_37743,N_36214,N_36419);
nor U37744 (N_37744,N_36668,N_36853);
xnor U37745 (N_37745,N_36547,N_36991);
nand U37746 (N_37746,N_36622,N_36188);
or U37747 (N_37747,N_36234,N_36597);
xor U37748 (N_37748,N_36116,N_36616);
nand U37749 (N_37749,N_36270,N_36005);
and U37750 (N_37750,N_36118,N_36191);
nor U37751 (N_37751,N_36663,N_36501);
or U37752 (N_37752,N_36900,N_36254);
and U37753 (N_37753,N_36973,N_36140);
nor U37754 (N_37754,N_36070,N_36400);
nand U37755 (N_37755,N_36733,N_36197);
nand U37756 (N_37756,N_36049,N_36518);
nor U37757 (N_37757,N_36006,N_36563);
or U37758 (N_37758,N_36153,N_36196);
or U37759 (N_37759,N_36634,N_36276);
nor U37760 (N_37760,N_36692,N_36993);
xor U37761 (N_37761,N_36645,N_36137);
xnor U37762 (N_37762,N_36063,N_36255);
nor U37763 (N_37763,N_36520,N_36997);
xor U37764 (N_37764,N_36457,N_36096);
and U37765 (N_37765,N_36283,N_36453);
nand U37766 (N_37766,N_36836,N_36721);
or U37767 (N_37767,N_36342,N_36758);
nand U37768 (N_37768,N_36962,N_36434);
and U37769 (N_37769,N_36658,N_36609);
xnor U37770 (N_37770,N_36089,N_36119);
or U37771 (N_37771,N_36688,N_36329);
nor U37772 (N_37772,N_36303,N_36372);
or U37773 (N_37773,N_36632,N_36305);
nand U37774 (N_37774,N_36433,N_36526);
xor U37775 (N_37775,N_36417,N_36670);
xnor U37776 (N_37776,N_36338,N_36301);
nor U37777 (N_37777,N_36686,N_36470);
or U37778 (N_37778,N_36954,N_36035);
nor U37779 (N_37779,N_36721,N_36354);
nor U37780 (N_37780,N_36694,N_36334);
or U37781 (N_37781,N_36551,N_36890);
or U37782 (N_37782,N_36026,N_36360);
and U37783 (N_37783,N_36880,N_36548);
nand U37784 (N_37784,N_36898,N_36701);
nor U37785 (N_37785,N_36462,N_36329);
and U37786 (N_37786,N_36639,N_36110);
and U37787 (N_37787,N_36770,N_36138);
nor U37788 (N_37788,N_36658,N_36679);
and U37789 (N_37789,N_36928,N_36895);
xnor U37790 (N_37790,N_36221,N_36159);
and U37791 (N_37791,N_36514,N_36510);
xor U37792 (N_37792,N_36461,N_36974);
nand U37793 (N_37793,N_36472,N_36264);
xnor U37794 (N_37794,N_36977,N_36445);
or U37795 (N_37795,N_36026,N_36898);
xor U37796 (N_37796,N_36488,N_36171);
and U37797 (N_37797,N_36931,N_36323);
or U37798 (N_37798,N_36049,N_36985);
nand U37799 (N_37799,N_36595,N_36120);
xnor U37800 (N_37800,N_36111,N_36789);
xor U37801 (N_37801,N_36173,N_36383);
nand U37802 (N_37802,N_36477,N_36166);
or U37803 (N_37803,N_36409,N_36396);
and U37804 (N_37804,N_36660,N_36569);
or U37805 (N_37805,N_36362,N_36590);
nand U37806 (N_37806,N_36134,N_36733);
xnor U37807 (N_37807,N_36439,N_36852);
xor U37808 (N_37808,N_36026,N_36100);
and U37809 (N_37809,N_36812,N_36505);
xnor U37810 (N_37810,N_36851,N_36487);
or U37811 (N_37811,N_36478,N_36325);
nor U37812 (N_37812,N_36485,N_36200);
nor U37813 (N_37813,N_36302,N_36340);
and U37814 (N_37814,N_36989,N_36827);
nor U37815 (N_37815,N_36144,N_36041);
xor U37816 (N_37816,N_36774,N_36553);
and U37817 (N_37817,N_36577,N_36542);
and U37818 (N_37818,N_36860,N_36085);
nor U37819 (N_37819,N_36900,N_36716);
and U37820 (N_37820,N_36559,N_36726);
nor U37821 (N_37821,N_36508,N_36529);
and U37822 (N_37822,N_36679,N_36739);
nand U37823 (N_37823,N_36435,N_36614);
or U37824 (N_37824,N_36100,N_36231);
nand U37825 (N_37825,N_36907,N_36455);
or U37826 (N_37826,N_36041,N_36392);
and U37827 (N_37827,N_36885,N_36227);
or U37828 (N_37828,N_36614,N_36854);
or U37829 (N_37829,N_36927,N_36413);
nor U37830 (N_37830,N_36489,N_36530);
nand U37831 (N_37831,N_36916,N_36113);
xnor U37832 (N_37832,N_36219,N_36607);
xnor U37833 (N_37833,N_36027,N_36155);
xnor U37834 (N_37834,N_36018,N_36761);
nand U37835 (N_37835,N_36119,N_36366);
or U37836 (N_37836,N_36842,N_36480);
nand U37837 (N_37837,N_36561,N_36597);
and U37838 (N_37838,N_36109,N_36289);
nand U37839 (N_37839,N_36218,N_36072);
and U37840 (N_37840,N_36872,N_36981);
and U37841 (N_37841,N_36545,N_36043);
nor U37842 (N_37842,N_36796,N_36039);
xor U37843 (N_37843,N_36480,N_36295);
or U37844 (N_37844,N_36307,N_36679);
xor U37845 (N_37845,N_36304,N_36159);
or U37846 (N_37846,N_36524,N_36682);
and U37847 (N_37847,N_36214,N_36674);
nor U37848 (N_37848,N_36398,N_36969);
nor U37849 (N_37849,N_36973,N_36394);
or U37850 (N_37850,N_36468,N_36961);
xor U37851 (N_37851,N_36027,N_36313);
or U37852 (N_37852,N_36358,N_36498);
or U37853 (N_37853,N_36584,N_36510);
nand U37854 (N_37854,N_36034,N_36579);
nand U37855 (N_37855,N_36534,N_36832);
or U37856 (N_37856,N_36458,N_36730);
or U37857 (N_37857,N_36686,N_36423);
nand U37858 (N_37858,N_36753,N_36026);
nand U37859 (N_37859,N_36749,N_36472);
and U37860 (N_37860,N_36004,N_36318);
nor U37861 (N_37861,N_36605,N_36615);
and U37862 (N_37862,N_36562,N_36021);
or U37863 (N_37863,N_36946,N_36714);
nor U37864 (N_37864,N_36929,N_36544);
or U37865 (N_37865,N_36906,N_36956);
nand U37866 (N_37866,N_36686,N_36879);
or U37867 (N_37867,N_36562,N_36762);
nand U37868 (N_37868,N_36748,N_36079);
or U37869 (N_37869,N_36912,N_36645);
xor U37870 (N_37870,N_36667,N_36343);
nor U37871 (N_37871,N_36615,N_36465);
xor U37872 (N_37872,N_36148,N_36883);
nor U37873 (N_37873,N_36389,N_36834);
nor U37874 (N_37874,N_36840,N_36778);
xnor U37875 (N_37875,N_36709,N_36153);
xnor U37876 (N_37876,N_36490,N_36223);
and U37877 (N_37877,N_36587,N_36804);
nor U37878 (N_37878,N_36315,N_36758);
xor U37879 (N_37879,N_36090,N_36915);
nand U37880 (N_37880,N_36403,N_36179);
and U37881 (N_37881,N_36810,N_36266);
nand U37882 (N_37882,N_36515,N_36575);
nand U37883 (N_37883,N_36245,N_36154);
xor U37884 (N_37884,N_36447,N_36168);
nor U37885 (N_37885,N_36817,N_36472);
xor U37886 (N_37886,N_36638,N_36769);
xnor U37887 (N_37887,N_36746,N_36575);
and U37888 (N_37888,N_36667,N_36533);
or U37889 (N_37889,N_36330,N_36888);
and U37890 (N_37890,N_36682,N_36411);
nand U37891 (N_37891,N_36867,N_36583);
nor U37892 (N_37892,N_36804,N_36831);
nor U37893 (N_37893,N_36774,N_36003);
or U37894 (N_37894,N_36402,N_36336);
and U37895 (N_37895,N_36744,N_36065);
nor U37896 (N_37896,N_36233,N_36828);
xnor U37897 (N_37897,N_36442,N_36082);
and U37898 (N_37898,N_36196,N_36881);
or U37899 (N_37899,N_36922,N_36550);
xnor U37900 (N_37900,N_36633,N_36829);
xnor U37901 (N_37901,N_36103,N_36162);
xnor U37902 (N_37902,N_36256,N_36772);
xor U37903 (N_37903,N_36897,N_36058);
nor U37904 (N_37904,N_36396,N_36577);
xor U37905 (N_37905,N_36057,N_36173);
xnor U37906 (N_37906,N_36971,N_36695);
xor U37907 (N_37907,N_36403,N_36501);
and U37908 (N_37908,N_36771,N_36605);
or U37909 (N_37909,N_36165,N_36284);
xor U37910 (N_37910,N_36079,N_36120);
and U37911 (N_37911,N_36406,N_36471);
nand U37912 (N_37912,N_36573,N_36227);
nor U37913 (N_37913,N_36370,N_36621);
and U37914 (N_37914,N_36074,N_36070);
nand U37915 (N_37915,N_36480,N_36364);
nand U37916 (N_37916,N_36457,N_36227);
and U37917 (N_37917,N_36241,N_36890);
nor U37918 (N_37918,N_36172,N_36810);
nand U37919 (N_37919,N_36599,N_36348);
and U37920 (N_37920,N_36884,N_36021);
and U37921 (N_37921,N_36969,N_36244);
xor U37922 (N_37922,N_36277,N_36426);
xor U37923 (N_37923,N_36376,N_36473);
nor U37924 (N_37924,N_36575,N_36520);
or U37925 (N_37925,N_36684,N_36770);
and U37926 (N_37926,N_36236,N_36124);
nor U37927 (N_37927,N_36057,N_36902);
nand U37928 (N_37928,N_36119,N_36831);
or U37929 (N_37929,N_36022,N_36414);
or U37930 (N_37930,N_36587,N_36625);
nand U37931 (N_37931,N_36059,N_36061);
nand U37932 (N_37932,N_36719,N_36601);
xnor U37933 (N_37933,N_36400,N_36549);
nor U37934 (N_37934,N_36705,N_36045);
xnor U37935 (N_37935,N_36840,N_36372);
nand U37936 (N_37936,N_36167,N_36523);
and U37937 (N_37937,N_36391,N_36470);
or U37938 (N_37938,N_36084,N_36809);
and U37939 (N_37939,N_36550,N_36995);
and U37940 (N_37940,N_36231,N_36044);
and U37941 (N_37941,N_36316,N_36125);
nand U37942 (N_37942,N_36793,N_36962);
and U37943 (N_37943,N_36065,N_36381);
or U37944 (N_37944,N_36894,N_36138);
or U37945 (N_37945,N_36688,N_36982);
nand U37946 (N_37946,N_36563,N_36427);
and U37947 (N_37947,N_36815,N_36134);
and U37948 (N_37948,N_36028,N_36247);
xor U37949 (N_37949,N_36574,N_36747);
nor U37950 (N_37950,N_36638,N_36062);
and U37951 (N_37951,N_36049,N_36533);
xnor U37952 (N_37952,N_36114,N_36615);
or U37953 (N_37953,N_36841,N_36205);
nand U37954 (N_37954,N_36018,N_36474);
nand U37955 (N_37955,N_36494,N_36059);
nand U37956 (N_37956,N_36906,N_36021);
xnor U37957 (N_37957,N_36286,N_36408);
nor U37958 (N_37958,N_36793,N_36990);
nand U37959 (N_37959,N_36090,N_36922);
nor U37960 (N_37960,N_36038,N_36735);
or U37961 (N_37961,N_36041,N_36468);
and U37962 (N_37962,N_36524,N_36489);
or U37963 (N_37963,N_36758,N_36533);
xor U37964 (N_37964,N_36245,N_36034);
or U37965 (N_37965,N_36911,N_36748);
xor U37966 (N_37966,N_36618,N_36213);
and U37967 (N_37967,N_36734,N_36289);
xor U37968 (N_37968,N_36127,N_36352);
nand U37969 (N_37969,N_36484,N_36522);
nor U37970 (N_37970,N_36016,N_36765);
xnor U37971 (N_37971,N_36637,N_36104);
xor U37972 (N_37972,N_36807,N_36301);
and U37973 (N_37973,N_36099,N_36567);
xnor U37974 (N_37974,N_36571,N_36039);
nand U37975 (N_37975,N_36227,N_36686);
nand U37976 (N_37976,N_36520,N_36181);
xnor U37977 (N_37977,N_36975,N_36984);
nor U37978 (N_37978,N_36426,N_36778);
nor U37979 (N_37979,N_36264,N_36507);
or U37980 (N_37980,N_36421,N_36537);
nor U37981 (N_37981,N_36534,N_36896);
and U37982 (N_37982,N_36052,N_36477);
nand U37983 (N_37983,N_36177,N_36657);
xor U37984 (N_37984,N_36768,N_36788);
xor U37985 (N_37985,N_36963,N_36972);
xnor U37986 (N_37986,N_36163,N_36436);
nand U37987 (N_37987,N_36782,N_36196);
xnor U37988 (N_37988,N_36233,N_36991);
and U37989 (N_37989,N_36764,N_36432);
nor U37990 (N_37990,N_36699,N_36023);
nor U37991 (N_37991,N_36367,N_36193);
or U37992 (N_37992,N_36564,N_36711);
nor U37993 (N_37993,N_36058,N_36029);
xor U37994 (N_37994,N_36504,N_36802);
and U37995 (N_37995,N_36257,N_36223);
xnor U37996 (N_37996,N_36798,N_36076);
nand U37997 (N_37997,N_36743,N_36309);
and U37998 (N_37998,N_36034,N_36736);
nand U37999 (N_37999,N_36388,N_36236);
xnor U38000 (N_38000,N_37081,N_37517);
nor U38001 (N_38001,N_37891,N_37624);
xnor U38002 (N_38002,N_37697,N_37144);
or U38003 (N_38003,N_37414,N_37955);
or U38004 (N_38004,N_37751,N_37605);
and U38005 (N_38005,N_37808,N_37723);
nor U38006 (N_38006,N_37028,N_37371);
xor U38007 (N_38007,N_37173,N_37689);
or U38008 (N_38008,N_37405,N_37893);
nor U38009 (N_38009,N_37107,N_37187);
and U38010 (N_38010,N_37454,N_37256);
or U38011 (N_38011,N_37630,N_37312);
or U38012 (N_38012,N_37411,N_37557);
and U38013 (N_38013,N_37135,N_37428);
nor U38014 (N_38014,N_37858,N_37920);
nor U38015 (N_38015,N_37492,N_37047);
or U38016 (N_38016,N_37325,N_37544);
and U38017 (N_38017,N_37532,N_37345);
or U38018 (N_38018,N_37155,N_37842);
nor U38019 (N_38019,N_37732,N_37967);
nand U38020 (N_38020,N_37277,N_37621);
nor U38021 (N_38021,N_37828,N_37318);
or U38022 (N_38022,N_37314,N_37847);
nor U38023 (N_38023,N_37044,N_37190);
and U38024 (N_38024,N_37211,N_37394);
and U38025 (N_38025,N_37498,N_37522);
nand U38026 (N_38026,N_37323,N_37613);
or U38027 (N_38027,N_37442,N_37865);
nor U38028 (N_38028,N_37840,N_37953);
or U38029 (N_38029,N_37871,N_37565);
xor U38030 (N_38030,N_37749,N_37238);
and U38031 (N_38031,N_37964,N_37679);
nand U38032 (N_38032,N_37823,N_37341);
or U38033 (N_38033,N_37734,N_37014);
and U38034 (N_38034,N_37108,N_37322);
nor U38035 (N_38035,N_37872,N_37569);
nand U38036 (N_38036,N_37397,N_37129);
xor U38037 (N_38037,N_37777,N_37590);
or U38038 (N_38038,N_37052,N_37868);
nand U38039 (N_38039,N_37539,N_37938);
or U38040 (N_38040,N_37609,N_37564);
nand U38041 (N_38041,N_37034,N_37064);
and U38042 (N_38042,N_37744,N_37655);
nor U38043 (N_38043,N_37490,N_37857);
nor U38044 (N_38044,N_37151,N_37281);
nor U38045 (N_38045,N_37758,N_37015);
or U38046 (N_38046,N_37352,N_37705);
and U38047 (N_38047,N_37321,N_37547);
or U38048 (N_38048,N_37250,N_37461);
nand U38049 (N_38049,N_37805,N_37313);
nor U38050 (N_38050,N_37368,N_37178);
nand U38051 (N_38051,N_37780,N_37257);
and U38052 (N_38052,N_37692,N_37104);
nand U38053 (N_38053,N_37924,N_37320);
xnor U38054 (N_38054,N_37551,N_37217);
nand U38055 (N_38055,N_37680,N_37410);
or U38056 (N_38056,N_37853,N_37119);
xor U38057 (N_38057,N_37543,N_37328);
nor U38058 (N_38058,N_37068,N_37272);
nor U38059 (N_38059,N_37648,N_37709);
xor U38060 (N_38060,N_37804,N_37619);
nor U38061 (N_38061,N_37737,N_37818);
nor U38062 (N_38062,N_37084,N_37399);
or U38063 (N_38063,N_37691,N_37851);
xnor U38064 (N_38064,N_37819,N_37741);
and U38065 (N_38065,N_37251,N_37164);
or U38066 (N_38066,N_37293,N_37997);
nand U38067 (N_38067,N_37562,N_37688);
xnor U38068 (N_38068,N_37229,N_37100);
xor U38069 (N_38069,N_37659,N_37887);
or U38070 (N_38070,N_37472,N_37426);
or U38071 (N_38071,N_37483,N_37286);
nand U38072 (N_38072,N_37413,N_37957);
nor U38073 (N_38073,N_37676,N_37861);
and U38074 (N_38074,N_37127,N_37403);
or U38075 (N_38075,N_37380,N_37167);
and U38076 (N_38076,N_37448,N_37530);
nor U38077 (N_38077,N_37574,N_37290);
xnor U38078 (N_38078,N_37841,N_37273);
xor U38079 (N_38079,N_37439,N_37264);
xnor U38080 (N_38080,N_37158,N_37126);
and U38081 (N_38081,N_37446,N_37702);
nor U38082 (N_38082,N_37572,N_37480);
nand U38083 (N_38083,N_37141,N_37351);
nand U38084 (N_38084,N_37360,N_37332);
xor U38085 (N_38085,N_37247,N_37188);
or U38086 (N_38086,N_37087,N_37346);
and U38087 (N_38087,N_37591,N_37958);
xor U38088 (N_38088,N_37379,N_37388);
and U38089 (N_38089,N_37166,N_37019);
nor U38090 (N_38090,N_37474,N_37215);
and U38091 (N_38091,N_37752,N_37079);
or U38092 (N_38092,N_37202,N_37627);
nand U38093 (N_38093,N_37932,N_37497);
nor U38094 (N_38094,N_37879,N_37401);
and U38095 (N_38095,N_37469,N_37903);
xnor U38096 (N_38096,N_37799,N_37935);
nor U38097 (N_38097,N_37189,N_37227);
nor U38098 (N_38098,N_37349,N_37424);
and U38099 (N_38099,N_37468,N_37241);
nand U38100 (N_38100,N_37310,N_37886);
nand U38101 (N_38101,N_37478,N_37011);
and U38102 (N_38102,N_37287,N_37364);
nor U38103 (N_38103,N_37059,N_37512);
and U38104 (N_38104,N_37025,N_37161);
xnor U38105 (N_38105,N_37456,N_37113);
or U38106 (N_38106,N_37396,N_37973);
xor U38107 (N_38107,N_37800,N_37832);
nor U38108 (N_38108,N_37546,N_37276);
nand U38109 (N_38109,N_37894,N_37746);
nand U38110 (N_38110,N_37010,N_37003);
xor U38111 (N_38111,N_37600,N_37145);
and U38112 (N_38112,N_37668,N_37101);
and U38113 (N_38113,N_37038,N_37802);
or U38114 (N_38114,N_37431,N_37897);
nor U38115 (N_38115,N_37634,N_37369);
and U38116 (N_38116,N_37131,N_37146);
or U38117 (N_38117,N_37707,N_37859);
xor U38118 (N_38118,N_37441,N_37766);
and U38119 (N_38119,N_37745,N_37343);
xnor U38120 (N_38120,N_37993,N_37631);
and U38121 (N_38121,N_37420,N_37996);
or U38122 (N_38122,N_37685,N_37669);
and U38123 (N_38123,N_37806,N_37999);
xnor U38124 (N_38124,N_37282,N_37502);
nand U38125 (N_38125,N_37421,N_37391);
or U38126 (N_38126,N_37743,N_37826);
xor U38127 (N_38127,N_37644,N_37724);
nand U38128 (N_38128,N_37460,N_37181);
nor U38129 (N_38129,N_37514,N_37665);
nor U38130 (N_38130,N_37533,N_37370);
xnor U38131 (N_38131,N_37537,N_37389);
or U38132 (N_38132,N_37226,N_37831);
xor U38133 (N_38133,N_37026,N_37417);
nor U38134 (N_38134,N_37348,N_37309);
or U38135 (N_38135,N_37169,N_37798);
and U38136 (N_38136,N_37425,N_37560);
nor U38137 (N_38137,N_37984,N_37147);
xnor U38138 (N_38138,N_37719,N_37355);
xnor U38139 (N_38139,N_37880,N_37177);
or U38140 (N_38140,N_37713,N_37022);
or U38141 (N_38141,N_37906,N_37392);
nand U38142 (N_38142,N_37636,N_37577);
or U38143 (N_38143,N_37239,N_37070);
nand U38144 (N_38144,N_37357,N_37266);
or U38145 (N_38145,N_37753,N_37850);
and U38146 (N_38146,N_37032,N_37130);
nand U38147 (N_38147,N_37657,N_37715);
xnor U38148 (N_38148,N_37299,N_37316);
and U38149 (N_38149,N_37513,N_37526);
nand U38150 (N_38150,N_37944,N_37548);
xor U38151 (N_38151,N_37268,N_37013);
or U38152 (N_38152,N_37267,N_37855);
nand U38153 (N_38153,N_37890,N_37742);
nor U38154 (N_38154,N_37733,N_37934);
and U38155 (N_38155,N_37765,N_37757);
xnor U38156 (N_38156,N_37788,N_37252);
nand U38157 (N_38157,N_37910,N_37035);
and U38158 (N_38158,N_37465,N_37782);
nand U38159 (N_38159,N_37128,N_37001);
nor U38160 (N_38160,N_37589,N_37201);
nor U38161 (N_38161,N_37311,N_37793);
nor U38162 (N_38162,N_37053,N_37327);
nor U38163 (N_38163,N_37595,N_37464);
or U38164 (N_38164,N_37307,N_37043);
nor U38165 (N_38165,N_37000,N_37885);
xnor U38166 (N_38166,N_37024,N_37970);
or U38167 (N_38167,N_37610,N_37249);
nor U38168 (N_38168,N_37489,N_37284);
and U38169 (N_38169,N_37869,N_37342);
xnor U38170 (N_38170,N_37712,N_37139);
nor U38171 (N_38171,N_37274,N_37566);
nand U38172 (N_38172,N_37763,N_37518);
nor U38173 (N_38173,N_37196,N_37720);
nor U38174 (N_38174,N_37585,N_37020);
xnor U38175 (N_38175,N_37940,N_37491);
nor U38176 (N_38176,N_37695,N_37142);
nor U38177 (N_38177,N_37338,N_37481);
and U38178 (N_38178,N_37193,N_37330);
nand U38179 (N_38179,N_37567,N_37783);
nand U38180 (N_38180,N_37913,N_37942);
and U38181 (N_38181,N_37750,N_37344);
or U38182 (N_38182,N_37242,N_37466);
or U38183 (N_38183,N_37398,N_37545);
and U38184 (N_38184,N_37255,N_37384);
or U38185 (N_38185,N_37748,N_37303);
nor U38186 (N_38186,N_37083,N_37874);
and U38187 (N_38187,N_37138,N_37747);
xnor U38188 (N_38188,N_37604,N_37559);
xnor U38189 (N_38189,N_37103,N_37736);
and U38190 (N_38190,N_37023,N_37649);
xor U38191 (N_38191,N_37701,N_37515);
or U38192 (N_38192,N_37837,N_37687);
xor U38193 (N_38193,N_37404,N_37952);
nor U38194 (N_38194,N_37110,N_37538);
or U38195 (N_38195,N_37521,N_37407);
nand U38196 (N_38196,N_37243,N_37007);
or U38197 (N_38197,N_37041,N_37834);
xor U38198 (N_38198,N_37774,N_37835);
nand U38199 (N_38199,N_37764,N_37914);
and U38200 (N_38200,N_37294,N_37246);
nor U38201 (N_38201,N_37280,N_37881);
nand U38202 (N_38202,N_37009,N_37825);
nor U38203 (N_38203,N_37488,N_37817);
and U38204 (N_38204,N_37236,N_37896);
or U38205 (N_38205,N_37909,N_37160);
or U38206 (N_38206,N_37708,N_37959);
and U38207 (N_38207,N_37063,N_37224);
xnor U38208 (N_38208,N_37437,N_37663);
xor U38209 (N_38209,N_37755,N_37986);
nand U38210 (N_38210,N_37773,N_37152);
xnor U38211 (N_38211,N_37867,N_37058);
and U38212 (N_38212,N_37664,N_37253);
xor U38213 (N_38213,N_37184,N_37596);
xnor U38214 (N_38214,N_37159,N_37419);
nand U38215 (N_38215,N_37939,N_37651);
or U38216 (N_38216,N_37143,N_37698);
or U38217 (N_38217,N_37077,N_37406);
and U38218 (N_38218,N_37194,N_37045);
nand U38219 (N_38219,N_37091,N_37434);
nand U38220 (N_38220,N_37218,N_37754);
xor U38221 (N_38221,N_37315,N_37527);
and U38222 (N_38222,N_37361,N_37639);
nor U38223 (N_38223,N_37990,N_37699);
nand U38224 (N_38224,N_37499,N_37915);
and U38225 (N_38225,N_37040,N_37899);
xor U38226 (N_38226,N_37186,N_37204);
xor U38227 (N_38227,N_37452,N_37830);
xnor U38228 (N_38228,N_37536,N_37995);
or U38229 (N_38229,N_37171,N_37012);
or U38230 (N_38230,N_37607,N_37317);
nand U38231 (N_38231,N_37535,N_37801);
and U38232 (N_38232,N_37580,N_37500);
nand U38233 (N_38233,N_37073,N_37505);
or U38234 (N_38234,N_37501,N_37653);
nand U38235 (N_38235,N_37597,N_37008);
and U38236 (N_38236,N_37761,N_37212);
nand U38237 (N_38237,N_37978,N_37432);
nand U38238 (N_38238,N_37016,N_37833);
or U38239 (N_38239,N_37195,N_37714);
and U38240 (N_38240,N_37172,N_37976);
and U38241 (N_38241,N_37767,N_37443);
and U38242 (N_38242,N_37279,N_37592);
nand U38243 (N_38243,N_37198,N_37122);
or U38244 (N_38244,N_37980,N_37156);
or U38245 (N_38245,N_37390,N_37907);
or U38246 (N_38246,N_37839,N_37561);
and U38247 (N_38247,N_37082,N_37436);
nand U38248 (N_38248,N_37092,N_37951);
or U38249 (N_38249,N_37162,N_37163);
and U38250 (N_38250,N_37416,N_37118);
and U38251 (N_38251,N_37529,N_37381);
xor U38252 (N_38252,N_37922,N_37670);
and U38253 (N_38253,N_37947,N_37694);
nor U38254 (N_38254,N_37180,N_37508);
nand U38255 (N_38255,N_37453,N_37376);
xor U38256 (N_38256,N_37223,N_37852);
nand U38257 (N_38257,N_37509,N_37516);
nand U38258 (N_38258,N_37233,N_37095);
xnor U38259 (N_38259,N_37039,N_37816);
nand U38260 (N_38260,N_37027,N_37221);
and U38261 (N_38261,N_37475,N_37088);
and U38262 (N_38262,N_37696,N_37271);
nand U38263 (N_38263,N_37372,N_37111);
and U38264 (N_38264,N_37354,N_37966);
xnor U38265 (N_38265,N_37191,N_37813);
nand U38266 (N_38266,N_37296,N_37060);
and U38267 (N_38267,N_37150,N_37347);
or U38268 (N_38268,N_37678,N_37430);
and U38269 (N_38269,N_37412,N_37598);
nand U38270 (N_38270,N_37329,N_37568);
nor U38271 (N_38271,N_37882,N_37807);
or U38272 (N_38272,N_37033,N_37046);
nand U38273 (N_38273,N_37956,N_37080);
xor U38274 (N_38274,N_37220,N_37706);
xnor U38275 (N_38275,N_37735,N_37511);
nor U38276 (N_38276,N_37074,N_37962);
nand U38277 (N_38277,N_37950,N_37941);
xor U38278 (N_38278,N_37614,N_37050);
and U38279 (N_38279,N_37427,N_37667);
nor U38280 (N_38280,N_37408,N_37477);
and U38281 (N_38281,N_37339,N_37207);
nor U38282 (N_38282,N_37261,N_37458);
nand U38283 (N_38283,N_37030,N_37586);
or U38284 (N_38284,N_37730,N_37048);
and U38285 (N_38285,N_37288,N_37640);
nor U38286 (N_38286,N_37541,N_37495);
nor U38287 (N_38287,N_37635,N_37504);
xor U38288 (N_38288,N_37213,N_37057);
or U38289 (N_38289,N_37165,N_37042);
xnor U38290 (N_38290,N_37245,N_37445);
nand U38291 (N_38291,N_37927,N_37090);
and U38292 (N_38292,N_37554,N_37216);
nor U38293 (N_38293,N_37656,N_37176);
xor U38294 (N_38294,N_37270,N_37291);
and U38295 (N_38295,N_37843,N_37588);
nand U38296 (N_38296,N_37623,N_37056);
and U38297 (N_38297,N_37301,N_37275);
nand U38298 (N_38298,N_37779,N_37968);
and U38299 (N_38299,N_37331,N_37051);
or U38300 (N_38300,N_37983,N_37677);
nor U38301 (N_38301,N_37866,N_37812);
xnor U38302 (N_38302,N_37094,N_37615);
or U38303 (N_38303,N_37974,N_37049);
or U38304 (N_38304,N_37726,N_37998);
xnor U38305 (N_38305,N_37228,N_37827);
xor U38306 (N_38306,N_37525,N_37963);
or U38307 (N_38307,N_37375,N_37862);
nor U38308 (N_38308,N_37089,N_37931);
xnor U38309 (N_38309,N_37948,N_37289);
and U38310 (N_38310,N_37031,N_37977);
xor U38311 (N_38311,N_37612,N_37877);
nand U38312 (N_38312,N_37440,N_37618);
nand U38313 (N_38313,N_37383,N_37029);
or U38314 (N_38314,N_37520,N_37298);
nand U38315 (N_38315,N_37455,N_37916);
xor U38316 (N_38316,N_37462,N_37558);
nand U38317 (N_38317,N_37192,N_37377);
nand U38318 (N_38318,N_37768,N_37304);
and U38319 (N_38319,N_37674,N_37148);
nand U38320 (N_38320,N_37098,N_37811);
and U38321 (N_38321,N_37433,N_37785);
or U38322 (N_38322,N_37225,N_37901);
nor U38323 (N_38323,N_37484,N_37265);
xor U38324 (N_38324,N_37153,N_37949);
xor U38325 (N_38325,N_37373,N_37124);
nand U38326 (N_38326,N_37334,N_37260);
or U38327 (N_38327,N_37673,N_37638);
or U38328 (N_38328,N_37283,N_37926);
nor U38329 (N_38329,N_37863,N_37494);
or U38330 (N_38330,N_37895,N_37097);
nor U38331 (N_38331,N_37704,N_37654);
and U38332 (N_38332,N_37711,N_37203);
nor U38333 (N_38333,N_37982,N_37601);
nand U38334 (N_38334,N_37581,N_37102);
xor U38335 (N_38335,N_37864,N_37510);
or U38336 (N_38336,N_37632,N_37259);
nand U38337 (N_38337,N_37550,N_37486);
xnor U38338 (N_38338,N_37583,N_37718);
nand U38339 (N_38339,N_37933,N_37686);
nor U38340 (N_38340,N_37285,N_37844);
xor U38341 (N_38341,N_37382,N_37506);
nor U38342 (N_38342,N_37797,N_37200);
xor U38343 (N_38343,N_37810,N_37625);
nand U38344 (N_38344,N_37071,N_37771);
and U38345 (N_38345,N_37240,N_37675);
or U38346 (N_38346,N_37523,N_37463);
nand U38347 (N_38347,N_37820,N_37792);
nor U38348 (N_38348,N_37326,N_37232);
or U38349 (N_38349,N_37386,N_37912);
xnor U38350 (N_38350,N_37450,N_37769);
or U38351 (N_38351,N_37929,N_37727);
or U38352 (N_38352,N_37519,N_37555);
nor U38353 (N_38353,N_37231,N_37721);
or U38354 (N_38354,N_37305,N_37295);
or U38355 (N_38355,N_37762,N_37870);
or U38356 (N_38356,N_37672,N_37888);
nand U38357 (N_38357,N_37900,N_37658);
or U38358 (N_38358,N_37086,N_37584);
and U38359 (N_38359,N_37336,N_37004);
nand U38360 (N_38360,N_37333,N_37571);
xor U38361 (N_38361,N_37503,N_37660);
or U38362 (N_38362,N_37292,N_37447);
xor U38363 (N_38363,N_37061,N_37902);
or U38364 (N_38364,N_37919,N_37067);
xnor U38365 (N_38365,N_37085,N_37395);
or U38366 (N_38366,N_37739,N_37829);
and U38367 (N_38367,N_37133,N_37994);
and U38368 (N_38368,N_37356,N_37845);
xnor U38369 (N_38369,N_37722,N_37482);
xnor U38370 (N_38370,N_37123,N_37197);
nand U38371 (N_38371,N_37066,N_37848);
nand U38372 (N_38372,N_37796,N_37770);
or U38373 (N_38373,N_37824,N_37740);
and U38374 (N_38374,N_37054,N_37205);
and U38375 (N_38375,N_37781,N_37496);
nand U38376 (N_38376,N_37873,N_37471);
nor U38377 (N_38377,N_37593,N_37815);
or U38378 (N_38378,N_37069,N_37269);
xnor U38379 (N_38379,N_37553,N_37531);
nand U38380 (N_38380,N_37803,N_37563);
nor U38381 (N_38381,N_37981,N_37789);
nor U38382 (N_38382,N_37006,N_37470);
nand U38383 (N_38383,N_37787,N_37620);
nand U38384 (N_38384,N_37552,N_37476);
or U38385 (N_38385,N_37182,N_37629);
nor U38386 (N_38386,N_37363,N_37928);
xor U38387 (N_38387,N_37822,N_37716);
nor U38388 (N_38388,N_37703,N_37617);
nand U38389 (N_38389,N_37418,N_37608);
nand U38390 (N_38390,N_37365,N_37300);
nor U38391 (N_38391,N_37875,N_37116);
and U38392 (N_38392,N_37093,N_37836);
or U38393 (N_38393,N_37661,N_37979);
nand U38394 (N_38394,N_37449,N_37175);
nand U38395 (N_38395,N_37002,N_37725);
nand U38396 (N_38396,N_37209,N_37775);
and U38397 (N_38397,N_37641,N_37650);
and U38398 (N_38398,N_37262,N_37402);
xnor U38399 (N_38399,N_37507,N_37791);
xnor U38400 (N_38400,N_37120,N_37248);
nor U38401 (N_38401,N_37918,N_37170);
or U38402 (N_38402,N_37645,N_37109);
xor U38403 (N_38403,N_37115,N_37021);
nand U38404 (N_38404,N_37611,N_37908);
xnor U38405 (N_38405,N_37278,N_37731);
and U38406 (N_38406,N_37930,N_37234);
xor U38407 (N_38407,N_37297,N_37892);
nand U38408 (N_38408,N_37263,N_37018);
nand U38409 (N_38409,N_37991,N_37444);
xnor U38410 (N_38410,N_37105,N_37965);
and U38411 (N_38411,N_37905,N_37235);
nand U38412 (N_38412,N_37786,N_37208);
or U38413 (N_38413,N_37121,N_37622);
or U38414 (N_38414,N_37992,N_37524);
nor U38415 (N_38415,N_37072,N_37710);
and U38416 (N_38416,N_37666,N_37222);
nand U38417 (N_38417,N_37626,N_37075);
and U38418 (N_38418,N_37633,N_37549);
xnor U38419 (N_38419,N_37700,N_37989);
nand U38420 (N_38420,N_37760,N_37671);
and U38421 (N_38421,N_37374,N_37065);
nand U38422 (N_38422,N_37237,N_37756);
xnor U38423 (N_38423,N_37578,N_37975);
xnor U38424 (N_38424,N_37878,N_37451);
or U38425 (N_38425,N_37717,N_37340);
and U38426 (N_38426,N_37599,N_37814);
nand U38427 (N_38427,N_37302,N_37157);
nand U38428 (N_38428,N_37540,N_37438);
nor U38429 (N_38429,N_37911,N_37062);
and U38430 (N_38430,N_37971,N_37206);
nand U38431 (N_38431,N_37628,N_37324);
and U38432 (N_38432,N_37112,N_37140);
xor U38433 (N_38433,N_37643,N_37219);
or U38434 (N_38434,N_37210,N_37795);
nor U38435 (N_38435,N_37961,N_37076);
and U38436 (N_38436,N_37467,N_37602);
xor U38437 (N_38437,N_37969,N_37943);
nand U38438 (N_38438,N_37078,N_37778);
or U38439 (N_38439,N_37214,N_37923);
xor U38440 (N_38440,N_37573,N_37898);
and U38441 (N_38441,N_37662,N_37359);
or U38442 (N_38442,N_37579,N_37772);
xor U38443 (N_38443,N_37616,N_37179);
nor U38444 (N_38444,N_37335,N_37821);
nand U38445 (N_38445,N_37642,N_37244);
nor U38446 (N_38446,N_37435,N_37925);
nand U38447 (N_38447,N_37759,N_37693);
xnor U38448 (N_38448,N_37684,N_37917);
or U38449 (N_38449,N_37846,N_37136);
nand U38450 (N_38450,N_37485,N_37682);
nand U38451 (N_38451,N_37556,N_37308);
and U38452 (N_38452,N_37594,N_37729);
nor U38453 (N_38453,N_37528,N_37921);
xor U38454 (N_38454,N_37603,N_37776);
or U38455 (N_38455,N_37385,N_37037);
or U38456 (N_38456,N_37936,N_37473);
or U38457 (N_38457,N_37415,N_37005);
xor U38458 (N_38458,N_37809,N_37849);
nor U38459 (N_38459,N_37429,N_37096);
xnor U38460 (N_38460,N_37125,N_37137);
nor U38461 (N_38461,N_37017,N_37972);
xor U38462 (N_38462,N_37884,N_37378);
nor U38463 (N_38463,N_37132,N_37790);
and U38464 (N_38464,N_37646,N_37937);
and U38465 (N_38465,N_37681,N_37183);
xor U38466 (N_38466,N_37606,N_37985);
nor U38467 (N_38467,N_37230,N_37362);
nand U38468 (N_38468,N_37946,N_37838);
and U38469 (N_38469,N_37784,N_37117);
nand U38470 (N_38470,N_37570,N_37367);
nand U38471 (N_38471,N_37690,N_37987);
or U38472 (N_38472,N_37587,N_37457);
nand U38473 (N_38473,N_37889,N_37954);
or U38474 (N_38474,N_37319,N_37306);
and U38475 (N_38475,N_37409,N_37960);
and U38476 (N_38476,N_37387,N_37199);
nor U38477 (N_38477,N_37988,N_37154);
nand U38478 (N_38478,N_37106,N_37254);
xnor U38479 (N_38479,N_37683,N_37794);
and U38480 (N_38480,N_37423,N_37149);
and U38481 (N_38481,N_37904,N_37493);
nand U38482 (N_38482,N_37353,N_37168);
nand U38483 (N_38483,N_37876,N_37534);
xor U38484 (N_38484,N_37174,N_37366);
xnor U38485 (N_38485,N_37055,N_37860);
and U38486 (N_38486,N_37350,N_37652);
nand U38487 (N_38487,N_37647,N_37728);
and U38488 (N_38488,N_37487,N_37400);
nor U38489 (N_38489,N_37542,N_37358);
nand U38490 (N_38490,N_37114,N_37582);
or U38491 (N_38491,N_37459,N_37393);
and U38492 (N_38492,N_37637,N_37337);
or U38493 (N_38493,N_37099,N_37258);
nor U38494 (N_38494,N_37036,N_37738);
and U38495 (N_38495,N_37134,N_37575);
nand U38496 (N_38496,N_37479,N_37576);
xnor U38497 (N_38497,N_37856,N_37185);
or U38498 (N_38498,N_37854,N_37883);
nand U38499 (N_38499,N_37422,N_37945);
xnor U38500 (N_38500,N_37079,N_37376);
nand U38501 (N_38501,N_37589,N_37699);
or U38502 (N_38502,N_37080,N_37703);
and U38503 (N_38503,N_37190,N_37975);
xnor U38504 (N_38504,N_37168,N_37157);
nand U38505 (N_38505,N_37761,N_37069);
xnor U38506 (N_38506,N_37006,N_37438);
or U38507 (N_38507,N_37473,N_37118);
xnor U38508 (N_38508,N_37165,N_37579);
nand U38509 (N_38509,N_37523,N_37514);
nand U38510 (N_38510,N_37280,N_37170);
nand U38511 (N_38511,N_37881,N_37146);
or U38512 (N_38512,N_37054,N_37267);
or U38513 (N_38513,N_37251,N_37792);
xnor U38514 (N_38514,N_37983,N_37646);
and U38515 (N_38515,N_37623,N_37261);
xor U38516 (N_38516,N_37707,N_37566);
nor U38517 (N_38517,N_37676,N_37318);
and U38518 (N_38518,N_37924,N_37517);
nand U38519 (N_38519,N_37201,N_37218);
or U38520 (N_38520,N_37687,N_37438);
and U38521 (N_38521,N_37088,N_37423);
xnor U38522 (N_38522,N_37026,N_37242);
xnor U38523 (N_38523,N_37904,N_37783);
nand U38524 (N_38524,N_37924,N_37520);
xnor U38525 (N_38525,N_37809,N_37768);
nand U38526 (N_38526,N_37601,N_37996);
nor U38527 (N_38527,N_37692,N_37429);
nand U38528 (N_38528,N_37097,N_37318);
xor U38529 (N_38529,N_37566,N_37298);
nand U38530 (N_38530,N_37584,N_37482);
nand U38531 (N_38531,N_37881,N_37645);
xnor U38532 (N_38532,N_37568,N_37731);
or U38533 (N_38533,N_37566,N_37670);
xor U38534 (N_38534,N_37884,N_37266);
xnor U38535 (N_38535,N_37192,N_37328);
nand U38536 (N_38536,N_37740,N_37126);
or U38537 (N_38537,N_37780,N_37904);
or U38538 (N_38538,N_37465,N_37275);
and U38539 (N_38539,N_37146,N_37708);
nand U38540 (N_38540,N_37478,N_37551);
nand U38541 (N_38541,N_37502,N_37000);
nor U38542 (N_38542,N_37378,N_37265);
and U38543 (N_38543,N_37474,N_37848);
nand U38544 (N_38544,N_37557,N_37731);
or U38545 (N_38545,N_37533,N_37242);
nor U38546 (N_38546,N_37120,N_37253);
nand U38547 (N_38547,N_37082,N_37671);
and U38548 (N_38548,N_37499,N_37579);
or U38549 (N_38549,N_37545,N_37546);
and U38550 (N_38550,N_37381,N_37626);
and U38551 (N_38551,N_37061,N_37884);
nand U38552 (N_38552,N_37910,N_37418);
or U38553 (N_38553,N_37089,N_37395);
xor U38554 (N_38554,N_37212,N_37677);
or U38555 (N_38555,N_37877,N_37617);
xor U38556 (N_38556,N_37101,N_37633);
xnor U38557 (N_38557,N_37031,N_37958);
or U38558 (N_38558,N_37750,N_37265);
or U38559 (N_38559,N_37060,N_37665);
or U38560 (N_38560,N_37453,N_37110);
and U38561 (N_38561,N_37229,N_37060);
nor U38562 (N_38562,N_37451,N_37701);
xnor U38563 (N_38563,N_37659,N_37801);
nand U38564 (N_38564,N_37072,N_37655);
nor U38565 (N_38565,N_37865,N_37744);
nor U38566 (N_38566,N_37833,N_37668);
nand U38567 (N_38567,N_37979,N_37281);
or U38568 (N_38568,N_37757,N_37578);
nand U38569 (N_38569,N_37331,N_37231);
and U38570 (N_38570,N_37963,N_37564);
and U38571 (N_38571,N_37823,N_37961);
or U38572 (N_38572,N_37452,N_37859);
nand U38573 (N_38573,N_37857,N_37163);
or U38574 (N_38574,N_37373,N_37782);
xnor U38575 (N_38575,N_37054,N_37546);
or U38576 (N_38576,N_37226,N_37242);
and U38577 (N_38577,N_37373,N_37771);
and U38578 (N_38578,N_37150,N_37803);
nand U38579 (N_38579,N_37945,N_37783);
and U38580 (N_38580,N_37912,N_37183);
or U38581 (N_38581,N_37012,N_37825);
or U38582 (N_38582,N_37263,N_37331);
nand U38583 (N_38583,N_37423,N_37099);
or U38584 (N_38584,N_37512,N_37219);
nand U38585 (N_38585,N_37135,N_37142);
or U38586 (N_38586,N_37863,N_37789);
nor U38587 (N_38587,N_37092,N_37408);
nor U38588 (N_38588,N_37378,N_37071);
and U38589 (N_38589,N_37455,N_37620);
or U38590 (N_38590,N_37172,N_37180);
nor U38591 (N_38591,N_37401,N_37660);
and U38592 (N_38592,N_37654,N_37370);
nor U38593 (N_38593,N_37159,N_37830);
xor U38594 (N_38594,N_37916,N_37575);
or U38595 (N_38595,N_37046,N_37353);
and U38596 (N_38596,N_37659,N_37357);
xor U38597 (N_38597,N_37584,N_37275);
nand U38598 (N_38598,N_37266,N_37731);
nor U38599 (N_38599,N_37044,N_37074);
xor U38600 (N_38600,N_37147,N_37860);
xnor U38601 (N_38601,N_37996,N_37567);
xor U38602 (N_38602,N_37914,N_37225);
xor U38603 (N_38603,N_37144,N_37591);
nand U38604 (N_38604,N_37789,N_37322);
or U38605 (N_38605,N_37894,N_37498);
and U38606 (N_38606,N_37320,N_37463);
nand U38607 (N_38607,N_37825,N_37295);
and U38608 (N_38608,N_37505,N_37346);
nor U38609 (N_38609,N_37782,N_37728);
or U38610 (N_38610,N_37260,N_37333);
nor U38611 (N_38611,N_37404,N_37307);
or U38612 (N_38612,N_37098,N_37616);
xnor U38613 (N_38613,N_37535,N_37995);
xnor U38614 (N_38614,N_37916,N_37903);
and U38615 (N_38615,N_37167,N_37009);
and U38616 (N_38616,N_37949,N_37045);
nand U38617 (N_38617,N_37897,N_37317);
and U38618 (N_38618,N_37418,N_37795);
or U38619 (N_38619,N_37844,N_37286);
and U38620 (N_38620,N_37438,N_37696);
xnor U38621 (N_38621,N_37084,N_37450);
xor U38622 (N_38622,N_37190,N_37088);
and U38623 (N_38623,N_37562,N_37730);
xnor U38624 (N_38624,N_37418,N_37843);
xnor U38625 (N_38625,N_37197,N_37259);
or U38626 (N_38626,N_37120,N_37381);
or U38627 (N_38627,N_37601,N_37067);
xnor U38628 (N_38628,N_37541,N_37115);
nand U38629 (N_38629,N_37089,N_37391);
or U38630 (N_38630,N_37316,N_37612);
or U38631 (N_38631,N_37919,N_37663);
or U38632 (N_38632,N_37889,N_37099);
nand U38633 (N_38633,N_37790,N_37016);
or U38634 (N_38634,N_37410,N_37243);
nor U38635 (N_38635,N_37776,N_37019);
and U38636 (N_38636,N_37104,N_37112);
and U38637 (N_38637,N_37433,N_37463);
nor U38638 (N_38638,N_37069,N_37821);
xor U38639 (N_38639,N_37189,N_37449);
nand U38640 (N_38640,N_37795,N_37616);
nand U38641 (N_38641,N_37148,N_37293);
xnor U38642 (N_38642,N_37140,N_37626);
and U38643 (N_38643,N_37137,N_37977);
nor U38644 (N_38644,N_37946,N_37124);
nand U38645 (N_38645,N_37927,N_37114);
nand U38646 (N_38646,N_37914,N_37847);
nor U38647 (N_38647,N_37571,N_37162);
and U38648 (N_38648,N_37944,N_37935);
or U38649 (N_38649,N_37527,N_37885);
nand U38650 (N_38650,N_37403,N_37884);
nor U38651 (N_38651,N_37724,N_37351);
xnor U38652 (N_38652,N_37007,N_37043);
xor U38653 (N_38653,N_37671,N_37219);
or U38654 (N_38654,N_37786,N_37890);
and U38655 (N_38655,N_37229,N_37684);
nor U38656 (N_38656,N_37625,N_37338);
nand U38657 (N_38657,N_37394,N_37559);
xor U38658 (N_38658,N_37959,N_37317);
and U38659 (N_38659,N_37540,N_37989);
nor U38660 (N_38660,N_37075,N_37553);
or U38661 (N_38661,N_37551,N_37992);
nor U38662 (N_38662,N_37302,N_37889);
xnor U38663 (N_38663,N_37380,N_37341);
nor U38664 (N_38664,N_37562,N_37629);
xor U38665 (N_38665,N_37863,N_37143);
nor U38666 (N_38666,N_37845,N_37000);
or U38667 (N_38667,N_37051,N_37236);
and U38668 (N_38668,N_37329,N_37937);
nand U38669 (N_38669,N_37225,N_37579);
or U38670 (N_38670,N_37323,N_37416);
xnor U38671 (N_38671,N_37419,N_37474);
nand U38672 (N_38672,N_37678,N_37520);
or U38673 (N_38673,N_37242,N_37057);
nand U38674 (N_38674,N_37480,N_37623);
xor U38675 (N_38675,N_37361,N_37722);
nand U38676 (N_38676,N_37936,N_37320);
nor U38677 (N_38677,N_37881,N_37068);
nand U38678 (N_38678,N_37975,N_37086);
xnor U38679 (N_38679,N_37068,N_37013);
nand U38680 (N_38680,N_37489,N_37051);
nand U38681 (N_38681,N_37934,N_37031);
nor U38682 (N_38682,N_37537,N_37949);
and U38683 (N_38683,N_37591,N_37440);
nor U38684 (N_38684,N_37480,N_37471);
xor U38685 (N_38685,N_37918,N_37341);
xor U38686 (N_38686,N_37965,N_37668);
or U38687 (N_38687,N_37966,N_37277);
and U38688 (N_38688,N_37178,N_37586);
nand U38689 (N_38689,N_37606,N_37632);
nand U38690 (N_38690,N_37515,N_37430);
nor U38691 (N_38691,N_37569,N_37292);
nand U38692 (N_38692,N_37714,N_37478);
nor U38693 (N_38693,N_37863,N_37899);
and U38694 (N_38694,N_37903,N_37501);
nor U38695 (N_38695,N_37412,N_37894);
xor U38696 (N_38696,N_37933,N_37961);
nand U38697 (N_38697,N_37432,N_37139);
or U38698 (N_38698,N_37078,N_37411);
xor U38699 (N_38699,N_37314,N_37306);
nand U38700 (N_38700,N_37570,N_37050);
nor U38701 (N_38701,N_37852,N_37755);
or U38702 (N_38702,N_37995,N_37189);
xnor U38703 (N_38703,N_37343,N_37530);
xnor U38704 (N_38704,N_37565,N_37675);
and U38705 (N_38705,N_37332,N_37045);
xor U38706 (N_38706,N_37884,N_37024);
and U38707 (N_38707,N_37782,N_37820);
nor U38708 (N_38708,N_37499,N_37560);
and U38709 (N_38709,N_37337,N_37978);
nand U38710 (N_38710,N_37343,N_37936);
xnor U38711 (N_38711,N_37320,N_37592);
nor U38712 (N_38712,N_37336,N_37550);
nor U38713 (N_38713,N_37236,N_37119);
and U38714 (N_38714,N_37967,N_37627);
or U38715 (N_38715,N_37558,N_37623);
nor U38716 (N_38716,N_37962,N_37307);
and U38717 (N_38717,N_37557,N_37675);
nor U38718 (N_38718,N_37125,N_37675);
and U38719 (N_38719,N_37358,N_37879);
or U38720 (N_38720,N_37577,N_37864);
xor U38721 (N_38721,N_37894,N_37906);
nor U38722 (N_38722,N_37975,N_37405);
xnor U38723 (N_38723,N_37470,N_37087);
nor U38724 (N_38724,N_37573,N_37621);
and U38725 (N_38725,N_37206,N_37169);
nand U38726 (N_38726,N_37013,N_37580);
nor U38727 (N_38727,N_37314,N_37846);
or U38728 (N_38728,N_37396,N_37467);
and U38729 (N_38729,N_37761,N_37675);
and U38730 (N_38730,N_37497,N_37724);
or U38731 (N_38731,N_37898,N_37280);
and U38732 (N_38732,N_37226,N_37673);
or U38733 (N_38733,N_37545,N_37563);
and U38734 (N_38734,N_37053,N_37428);
nor U38735 (N_38735,N_37839,N_37849);
and U38736 (N_38736,N_37442,N_37849);
nand U38737 (N_38737,N_37637,N_37240);
or U38738 (N_38738,N_37060,N_37722);
and U38739 (N_38739,N_37404,N_37588);
nor U38740 (N_38740,N_37749,N_37956);
or U38741 (N_38741,N_37046,N_37637);
nor U38742 (N_38742,N_37517,N_37295);
nand U38743 (N_38743,N_37032,N_37161);
or U38744 (N_38744,N_37172,N_37130);
nand U38745 (N_38745,N_37750,N_37921);
or U38746 (N_38746,N_37680,N_37153);
xnor U38747 (N_38747,N_37635,N_37774);
nor U38748 (N_38748,N_37129,N_37218);
nor U38749 (N_38749,N_37962,N_37293);
or U38750 (N_38750,N_37224,N_37015);
nand U38751 (N_38751,N_37612,N_37462);
nor U38752 (N_38752,N_37581,N_37343);
xnor U38753 (N_38753,N_37726,N_37854);
and U38754 (N_38754,N_37168,N_37507);
and U38755 (N_38755,N_37437,N_37544);
or U38756 (N_38756,N_37927,N_37596);
and U38757 (N_38757,N_37765,N_37340);
nand U38758 (N_38758,N_37385,N_37808);
and U38759 (N_38759,N_37688,N_37407);
nor U38760 (N_38760,N_37172,N_37872);
xor U38761 (N_38761,N_37480,N_37498);
and U38762 (N_38762,N_37022,N_37826);
xnor U38763 (N_38763,N_37808,N_37961);
xor U38764 (N_38764,N_37196,N_37217);
xor U38765 (N_38765,N_37260,N_37954);
or U38766 (N_38766,N_37855,N_37561);
nor U38767 (N_38767,N_37547,N_37658);
or U38768 (N_38768,N_37957,N_37394);
nand U38769 (N_38769,N_37785,N_37408);
or U38770 (N_38770,N_37904,N_37227);
and U38771 (N_38771,N_37918,N_37883);
and U38772 (N_38772,N_37272,N_37210);
xor U38773 (N_38773,N_37884,N_37337);
and U38774 (N_38774,N_37289,N_37852);
and U38775 (N_38775,N_37527,N_37005);
xnor U38776 (N_38776,N_37930,N_37873);
nand U38777 (N_38777,N_37610,N_37473);
and U38778 (N_38778,N_37967,N_37472);
nor U38779 (N_38779,N_37688,N_37293);
nand U38780 (N_38780,N_37343,N_37087);
nand U38781 (N_38781,N_37513,N_37928);
and U38782 (N_38782,N_37178,N_37136);
nand U38783 (N_38783,N_37076,N_37868);
nor U38784 (N_38784,N_37591,N_37744);
or U38785 (N_38785,N_37614,N_37084);
nand U38786 (N_38786,N_37608,N_37213);
nor U38787 (N_38787,N_37617,N_37610);
nor U38788 (N_38788,N_37093,N_37294);
and U38789 (N_38789,N_37085,N_37131);
or U38790 (N_38790,N_37035,N_37437);
xor U38791 (N_38791,N_37240,N_37271);
nor U38792 (N_38792,N_37791,N_37194);
nand U38793 (N_38793,N_37791,N_37678);
xor U38794 (N_38794,N_37071,N_37113);
and U38795 (N_38795,N_37643,N_37121);
or U38796 (N_38796,N_37666,N_37360);
nand U38797 (N_38797,N_37211,N_37311);
nand U38798 (N_38798,N_37120,N_37201);
or U38799 (N_38799,N_37833,N_37736);
nand U38800 (N_38800,N_37792,N_37399);
and U38801 (N_38801,N_37368,N_37733);
or U38802 (N_38802,N_37773,N_37832);
nand U38803 (N_38803,N_37721,N_37719);
xnor U38804 (N_38804,N_37804,N_37348);
and U38805 (N_38805,N_37269,N_37021);
nand U38806 (N_38806,N_37797,N_37874);
nor U38807 (N_38807,N_37125,N_37185);
nor U38808 (N_38808,N_37725,N_37254);
or U38809 (N_38809,N_37918,N_37266);
nor U38810 (N_38810,N_37355,N_37362);
and U38811 (N_38811,N_37242,N_37434);
and U38812 (N_38812,N_37628,N_37901);
and U38813 (N_38813,N_37090,N_37044);
nor U38814 (N_38814,N_37647,N_37288);
nand U38815 (N_38815,N_37127,N_37641);
nor U38816 (N_38816,N_37230,N_37587);
nor U38817 (N_38817,N_37218,N_37594);
or U38818 (N_38818,N_37433,N_37671);
and U38819 (N_38819,N_37404,N_37473);
and U38820 (N_38820,N_37733,N_37212);
and U38821 (N_38821,N_37819,N_37134);
xnor U38822 (N_38822,N_37421,N_37414);
nor U38823 (N_38823,N_37502,N_37786);
xor U38824 (N_38824,N_37827,N_37193);
or U38825 (N_38825,N_37551,N_37547);
xnor U38826 (N_38826,N_37808,N_37106);
and U38827 (N_38827,N_37340,N_37192);
nand U38828 (N_38828,N_37560,N_37177);
or U38829 (N_38829,N_37311,N_37605);
nor U38830 (N_38830,N_37020,N_37841);
or U38831 (N_38831,N_37437,N_37552);
nand U38832 (N_38832,N_37919,N_37928);
and U38833 (N_38833,N_37804,N_37860);
or U38834 (N_38834,N_37040,N_37952);
and U38835 (N_38835,N_37152,N_37603);
nand U38836 (N_38836,N_37650,N_37024);
or U38837 (N_38837,N_37381,N_37678);
or U38838 (N_38838,N_37895,N_37966);
nand U38839 (N_38839,N_37976,N_37571);
or U38840 (N_38840,N_37982,N_37651);
or U38841 (N_38841,N_37291,N_37592);
xnor U38842 (N_38842,N_37941,N_37217);
nand U38843 (N_38843,N_37701,N_37417);
or U38844 (N_38844,N_37752,N_37834);
or U38845 (N_38845,N_37594,N_37035);
or U38846 (N_38846,N_37817,N_37088);
or U38847 (N_38847,N_37646,N_37056);
xnor U38848 (N_38848,N_37401,N_37070);
xnor U38849 (N_38849,N_37214,N_37623);
nand U38850 (N_38850,N_37090,N_37317);
and U38851 (N_38851,N_37291,N_37362);
nor U38852 (N_38852,N_37575,N_37649);
xor U38853 (N_38853,N_37394,N_37994);
xnor U38854 (N_38854,N_37373,N_37389);
xnor U38855 (N_38855,N_37974,N_37284);
nor U38856 (N_38856,N_37177,N_37849);
or U38857 (N_38857,N_37869,N_37113);
or U38858 (N_38858,N_37854,N_37673);
and U38859 (N_38859,N_37742,N_37058);
or U38860 (N_38860,N_37738,N_37011);
or U38861 (N_38861,N_37384,N_37245);
nand U38862 (N_38862,N_37556,N_37010);
and U38863 (N_38863,N_37052,N_37609);
or U38864 (N_38864,N_37834,N_37590);
xnor U38865 (N_38865,N_37322,N_37426);
xnor U38866 (N_38866,N_37455,N_37838);
nand U38867 (N_38867,N_37570,N_37481);
nand U38868 (N_38868,N_37847,N_37303);
nand U38869 (N_38869,N_37875,N_37383);
xor U38870 (N_38870,N_37324,N_37049);
nor U38871 (N_38871,N_37304,N_37601);
and U38872 (N_38872,N_37801,N_37020);
or U38873 (N_38873,N_37458,N_37507);
nor U38874 (N_38874,N_37175,N_37239);
nand U38875 (N_38875,N_37694,N_37049);
or U38876 (N_38876,N_37766,N_37592);
and U38877 (N_38877,N_37022,N_37091);
nor U38878 (N_38878,N_37214,N_37043);
or U38879 (N_38879,N_37455,N_37068);
nand U38880 (N_38880,N_37013,N_37139);
nor U38881 (N_38881,N_37561,N_37568);
or U38882 (N_38882,N_37713,N_37018);
or U38883 (N_38883,N_37299,N_37762);
nor U38884 (N_38884,N_37373,N_37388);
xor U38885 (N_38885,N_37214,N_37827);
xor U38886 (N_38886,N_37562,N_37081);
nor U38887 (N_38887,N_37033,N_37201);
nand U38888 (N_38888,N_37070,N_37680);
xnor U38889 (N_38889,N_37640,N_37407);
or U38890 (N_38890,N_37785,N_37075);
nand U38891 (N_38891,N_37868,N_37112);
nor U38892 (N_38892,N_37573,N_37273);
or U38893 (N_38893,N_37764,N_37486);
nand U38894 (N_38894,N_37625,N_37886);
xnor U38895 (N_38895,N_37755,N_37805);
or U38896 (N_38896,N_37271,N_37248);
xnor U38897 (N_38897,N_37513,N_37705);
nor U38898 (N_38898,N_37741,N_37820);
or U38899 (N_38899,N_37224,N_37723);
nor U38900 (N_38900,N_37312,N_37001);
xor U38901 (N_38901,N_37157,N_37415);
or U38902 (N_38902,N_37795,N_37522);
xnor U38903 (N_38903,N_37949,N_37878);
nand U38904 (N_38904,N_37327,N_37462);
nand U38905 (N_38905,N_37021,N_37506);
nand U38906 (N_38906,N_37134,N_37192);
nor U38907 (N_38907,N_37280,N_37748);
and U38908 (N_38908,N_37281,N_37988);
nand U38909 (N_38909,N_37187,N_37399);
xor U38910 (N_38910,N_37449,N_37847);
nand U38911 (N_38911,N_37479,N_37257);
xor U38912 (N_38912,N_37426,N_37405);
nor U38913 (N_38913,N_37336,N_37725);
xor U38914 (N_38914,N_37253,N_37476);
xnor U38915 (N_38915,N_37853,N_37576);
nand U38916 (N_38916,N_37894,N_37843);
or U38917 (N_38917,N_37478,N_37248);
nor U38918 (N_38918,N_37589,N_37747);
or U38919 (N_38919,N_37121,N_37915);
or U38920 (N_38920,N_37355,N_37075);
xnor U38921 (N_38921,N_37521,N_37055);
nor U38922 (N_38922,N_37760,N_37656);
and U38923 (N_38923,N_37420,N_37527);
and U38924 (N_38924,N_37000,N_37335);
nor U38925 (N_38925,N_37317,N_37146);
nor U38926 (N_38926,N_37304,N_37643);
and U38927 (N_38927,N_37643,N_37867);
or U38928 (N_38928,N_37867,N_37707);
and U38929 (N_38929,N_37993,N_37350);
nand U38930 (N_38930,N_37022,N_37049);
xnor U38931 (N_38931,N_37854,N_37629);
nor U38932 (N_38932,N_37321,N_37969);
and U38933 (N_38933,N_37739,N_37556);
xnor U38934 (N_38934,N_37430,N_37978);
nand U38935 (N_38935,N_37466,N_37769);
nand U38936 (N_38936,N_37708,N_37776);
and U38937 (N_38937,N_37078,N_37940);
xnor U38938 (N_38938,N_37580,N_37115);
nor U38939 (N_38939,N_37803,N_37539);
nor U38940 (N_38940,N_37302,N_37971);
nand U38941 (N_38941,N_37759,N_37841);
nand U38942 (N_38942,N_37140,N_37806);
nor U38943 (N_38943,N_37625,N_37567);
xnor U38944 (N_38944,N_37758,N_37511);
nor U38945 (N_38945,N_37066,N_37150);
and U38946 (N_38946,N_37718,N_37778);
xor U38947 (N_38947,N_37137,N_37107);
nor U38948 (N_38948,N_37824,N_37328);
nor U38949 (N_38949,N_37486,N_37216);
xnor U38950 (N_38950,N_37490,N_37326);
or U38951 (N_38951,N_37051,N_37408);
xnor U38952 (N_38952,N_37344,N_37842);
and U38953 (N_38953,N_37699,N_37086);
xnor U38954 (N_38954,N_37393,N_37208);
nand U38955 (N_38955,N_37030,N_37785);
nand U38956 (N_38956,N_37357,N_37356);
and U38957 (N_38957,N_37072,N_37695);
nand U38958 (N_38958,N_37696,N_37992);
or U38959 (N_38959,N_37087,N_37120);
or U38960 (N_38960,N_37434,N_37012);
xnor U38961 (N_38961,N_37416,N_37296);
nand U38962 (N_38962,N_37068,N_37417);
xor U38963 (N_38963,N_37955,N_37679);
and U38964 (N_38964,N_37574,N_37277);
nor U38965 (N_38965,N_37603,N_37825);
nor U38966 (N_38966,N_37527,N_37692);
xor U38967 (N_38967,N_37305,N_37851);
xnor U38968 (N_38968,N_37961,N_37324);
nand U38969 (N_38969,N_37751,N_37280);
xnor U38970 (N_38970,N_37217,N_37400);
or U38971 (N_38971,N_37447,N_37104);
nand U38972 (N_38972,N_37261,N_37536);
nand U38973 (N_38973,N_37455,N_37349);
nand U38974 (N_38974,N_37839,N_37163);
or U38975 (N_38975,N_37440,N_37537);
and U38976 (N_38976,N_37292,N_37638);
nor U38977 (N_38977,N_37327,N_37349);
nand U38978 (N_38978,N_37399,N_37628);
or U38979 (N_38979,N_37875,N_37630);
nand U38980 (N_38980,N_37641,N_37114);
nand U38981 (N_38981,N_37451,N_37816);
and U38982 (N_38982,N_37552,N_37488);
nor U38983 (N_38983,N_37409,N_37807);
xnor U38984 (N_38984,N_37605,N_37531);
nand U38985 (N_38985,N_37428,N_37010);
or U38986 (N_38986,N_37063,N_37305);
nor U38987 (N_38987,N_37183,N_37273);
and U38988 (N_38988,N_37009,N_37966);
and U38989 (N_38989,N_37192,N_37010);
nor U38990 (N_38990,N_37672,N_37441);
and U38991 (N_38991,N_37835,N_37942);
xnor U38992 (N_38992,N_37616,N_37975);
nor U38993 (N_38993,N_37837,N_37739);
nor U38994 (N_38994,N_37446,N_37010);
nand U38995 (N_38995,N_37232,N_37833);
xor U38996 (N_38996,N_37532,N_37260);
and U38997 (N_38997,N_37947,N_37043);
and U38998 (N_38998,N_37825,N_37717);
nor U38999 (N_38999,N_37320,N_37959);
nor U39000 (N_39000,N_38183,N_38247);
xnor U39001 (N_39001,N_38105,N_38187);
or U39002 (N_39002,N_38744,N_38946);
or U39003 (N_39003,N_38035,N_38264);
or U39004 (N_39004,N_38535,N_38165);
or U39005 (N_39005,N_38170,N_38297);
nor U39006 (N_39006,N_38641,N_38850);
and U39007 (N_39007,N_38468,N_38409);
or U39008 (N_39008,N_38254,N_38756);
xor U39009 (N_39009,N_38869,N_38415);
nand U39010 (N_39010,N_38366,N_38001);
nand U39011 (N_39011,N_38633,N_38494);
or U39012 (N_39012,N_38392,N_38249);
nand U39013 (N_39013,N_38844,N_38050);
nand U39014 (N_39014,N_38899,N_38194);
nand U39015 (N_39015,N_38288,N_38999);
or U39016 (N_39016,N_38482,N_38060);
xor U39017 (N_39017,N_38752,N_38476);
or U39018 (N_39018,N_38630,N_38093);
or U39019 (N_39019,N_38370,N_38843);
xnor U39020 (N_39020,N_38250,N_38522);
and U39021 (N_39021,N_38296,N_38385);
xor U39022 (N_39022,N_38009,N_38189);
nand U39023 (N_39023,N_38957,N_38578);
nand U39024 (N_39024,N_38367,N_38809);
or U39025 (N_39025,N_38123,N_38348);
or U39026 (N_39026,N_38089,N_38424);
nand U39027 (N_39027,N_38386,N_38803);
nand U39028 (N_39028,N_38175,N_38567);
and U39029 (N_39029,N_38582,N_38776);
or U39030 (N_39030,N_38061,N_38629);
xor U39031 (N_39031,N_38785,N_38885);
and U39032 (N_39032,N_38239,N_38595);
nor U39033 (N_39033,N_38954,N_38458);
nor U39034 (N_39034,N_38882,N_38671);
and U39035 (N_39035,N_38573,N_38719);
and U39036 (N_39036,N_38903,N_38102);
nor U39037 (N_39037,N_38434,N_38717);
nor U39038 (N_39038,N_38975,N_38904);
xnor U39039 (N_39039,N_38352,N_38234);
nand U39040 (N_39040,N_38730,N_38678);
nand U39041 (N_39041,N_38268,N_38549);
or U39042 (N_39042,N_38265,N_38586);
and U39043 (N_39043,N_38881,N_38935);
or U39044 (N_39044,N_38474,N_38200);
or U39045 (N_39045,N_38451,N_38256);
nand U39046 (N_39046,N_38081,N_38351);
nand U39047 (N_39047,N_38116,N_38537);
nand U39048 (N_39048,N_38072,N_38188);
xnor U39049 (N_39049,N_38226,N_38006);
and U39050 (N_39050,N_38968,N_38158);
nand U39051 (N_39051,N_38435,N_38279);
and U39052 (N_39052,N_38360,N_38670);
and U39053 (N_39053,N_38777,N_38143);
xnor U39054 (N_39054,N_38651,N_38736);
xnor U39055 (N_39055,N_38594,N_38680);
xor U39056 (N_39056,N_38393,N_38475);
xnor U39057 (N_39057,N_38026,N_38673);
xnor U39058 (N_39058,N_38856,N_38179);
or U39059 (N_39059,N_38526,N_38363);
nor U39060 (N_39060,N_38862,N_38519);
and U39061 (N_39061,N_38337,N_38760);
or U39062 (N_39062,N_38318,N_38868);
nand U39063 (N_39063,N_38202,N_38379);
and U39064 (N_39064,N_38378,N_38119);
or U39065 (N_39065,N_38615,N_38577);
nor U39066 (N_39066,N_38263,N_38910);
nor U39067 (N_39067,N_38109,N_38912);
nor U39068 (N_39068,N_38837,N_38602);
and U39069 (N_39069,N_38665,N_38332);
nor U39070 (N_39070,N_38977,N_38255);
nor U39071 (N_39071,N_38502,N_38399);
nor U39072 (N_39072,N_38959,N_38137);
nor U39073 (N_39073,N_38388,N_38099);
nand U39074 (N_39074,N_38635,N_38056);
and U39075 (N_39075,N_38324,N_38932);
xnor U39076 (N_39076,N_38723,N_38949);
and U39077 (N_39077,N_38252,N_38446);
nor U39078 (N_39078,N_38224,N_38390);
xor U39079 (N_39079,N_38739,N_38996);
or U39080 (N_39080,N_38025,N_38427);
or U39081 (N_39081,N_38755,N_38317);
nand U39082 (N_39082,N_38127,N_38192);
and U39083 (N_39083,N_38811,N_38998);
and U39084 (N_39084,N_38005,N_38488);
and U39085 (N_39085,N_38548,N_38135);
xor U39086 (N_39086,N_38147,N_38293);
or U39087 (N_39087,N_38813,N_38425);
xor U39088 (N_39088,N_38128,N_38244);
nor U39089 (N_39089,N_38682,N_38889);
nand U39090 (N_39090,N_38753,N_38152);
or U39091 (N_39091,N_38375,N_38429);
nand U39092 (N_39092,N_38566,N_38693);
and U39093 (N_39093,N_38273,N_38171);
nand U39094 (N_39094,N_38489,N_38627);
or U39095 (N_39095,N_38692,N_38312);
nor U39096 (N_39096,N_38138,N_38213);
and U39097 (N_39097,N_38459,N_38598);
nand U39098 (N_39098,N_38536,N_38107);
nor U39099 (N_39099,N_38965,N_38111);
xor U39100 (N_39100,N_38068,N_38544);
xor U39101 (N_39101,N_38849,N_38788);
xnor U39102 (N_39102,N_38113,N_38369);
and U39103 (N_39103,N_38420,N_38880);
nor U39104 (N_39104,N_38883,N_38738);
nor U39105 (N_39105,N_38782,N_38745);
and U39106 (N_39106,N_38937,N_38770);
nor U39107 (N_39107,N_38098,N_38330);
xor U39108 (N_39108,N_38303,N_38087);
xor U39109 (N_39109,N_38555,N_38829);
nand U39110 (N_39110,N_38642,N_38896);
and U39111 (N_39111,N_38043,N_38951);
xor U39112 (N_39112,N_38416,N_38620);
xnor U39113 (N_39113,N_38477,N_38302);
nor U39114 (N_39114,N_38685,N_38162);
xor U39115 (N_39115,N_38078,N_38022);
nand U39116 (N_39116,N_38568,N_38705);
nand U39117 (N_39117,N_38810,N_38735);
nor U39118 (N_39118,N_38579,N_38948);
and U39119 (N_39119,N_38059,N_38701);
nand U39120 (N_39120,N_38824,N_38203);
and U39121 (N_39121,N_38789,N_38928);
and U39122 (N_39122,N_38306,N_38500);
nand U39123 (N_39123,N_38840,N_38146);
nor U39124 (N_39124,N_38501,N_38845);
xor U39125 (N_39125,N_38004,N_38181);
nor U39126 (N_39126,N_38758,N_38024);
or U39127 (N_39127,N_38356,N_38800);
nand U39128 (N_39128,N_38686,N_38497);
and U39129 (N_39129,N_38820,N_38492);
or U39130 (N_39130,N_38359,N_38724);
nor U39131 (N_39131,N_38246,N_38030);
and U39132 (N_39132,N_38301,N_38394);
or U39133 (N_39133,N_38761,N_38097);
nand U39134 (N_39134,N_38016,N_38877);
xor U39135 (N_39135,N_38623,N_38212);
nor U39136 (N_39136,N_38812,N_38511);
nor U39137 (N_39137,N_38963,N_38484);
nor U39138 (N_39138,N_38539,N_38606);
nand U39139 (N_39139,N_38503,N_38382);
nor U39140 (N_39140,N_38229,N_38792);
nor U39141 (N_39141,N_38180,N_38909);
and U39142 (N_39142,N_38504,N_38655);
or U39143 (N_39143,N_38865,N_38133);
xor U39144 (N_39144,N_38887,N_38900);
or U39145 (N_39145,N_38973,N_38626);
xnor U39146 (N_39146,N_38561,N_38797);
nor U39147 (N_39147,N_38986,N_38649);
nand U39148 (N_39148,N_38283,N_38190);
xor U39149 (N_39149,N_38086,N_38990);
or U39150 (N_39150,N_38600,N_38074);
nand U39151 (N_39151,N_38406,N_38534);
or U39152 (N_39152,N_38646,N_38095);
nor U39153 (N_39153,N_38275,N_38173);
nand U39154 (N_39154,N_38140,N_38601);
nand U39155 (N_39155,N_38523,N_38737);
nand U39156 (N_39156,N_38457,N_38679);
or U39157 (N_39157,N_38159,N_38510);
xor U39158 (N_39158,N_38884,N_38764);
or U39159 (N_39159,N_38478,N_38211);
and U39160 (N_39160,N_38463,N_38284);
nor U39161 (N_39161,N_38855,N_38778);
nand U39162 (N_39162,N_38647,N_38533);
nor U39163 (N_39163,N_38514,N_38821);
and U39164 (N_39164,N_38483,N_38790);
or U39165 (N_39165,N_38280,N_38470);
or U39166 (N_39166,N_38219,N_38253);
xor U39167 (N_39167,N_38709,N_38704);
or U39168 (N_39168,N_38417,N_38729);
nand U39169 (N_39169,N_38836,N_38643);
nor U39170 (N_39170,N_38319,N_38515);
nand U39171 (N_39171,N_38418,N_38530);
xor U39172 (N_39172,N_38982,N_38681);
nor U39173 (N_39173,N_38216,N_38498);
and U39174 (N_39174,N_38570,N_38795);
and U39175 (N_39175,N_38160,N_38334);
or U39176 (N_39176,N_38931,N_38859);
nand U39177 (N_39177,N_38532,N_38983);
or U39178 (N_39178,N_38167,N_38767);
or U39179 (N_39179,N_38267,N_38727);
xor U39180 (N_39180,N_38053,N_38412);
nand U39181 (N_39181,N_38543,N_38985);
or U39182 (N_39182,N_38374,N_38291);
nor U39183 (N_39183,N_38220,N_38277);
or U39184 (N_39184,N_38080,N_38471);
nor U39185 (N_39185,N_38395,N_38323);
xor U39186 (N_39186,N_38270,N_38636);
and U39187 (N_39187,N_38926,N_38624);
and U39188 (N_39188,N_38428,N_38310);
or U39189 (N_39189,N_38294,N_38460);
nand U39190 (N_39190,N_38553,N_38694);
nor U39191 (N_39191,N_38690,N_38631);
nor U39192 (N_39192,N_38018,N_38377);
xnor U39193 (N_39193,N_38058,N_38902);
and U39194 (N_39194,N_38886,N_38712);
xnor U39195 (N_39195,N_38151,N_38144);
and U39196 (N_39196,N_38657,N_38920);
or U39197 (N_39197,N_38611,N_38528);
or U39198 (N_39198,N_38227,N_38066);
nor U39199 (N_39199,N_38698,N_38002);
nand U39200 (N_39200,N_38632,N_38117);
nand U39201 (N_39201,N_38397,N_38852);
xor U39202 (N_39202,N_38734,N_38944);
nor U39203 (N_39203,N_38947,N_38974);
nand U39204 (N_39204,N_38833,N_38069);
nand U39205 (N_39205,N_38593,N_38667);
nor U39206 (N_39206,N_38401,N_38962);
xor U39207 (N_39207,N_38346,N_38972);
or U39208 (N_39208,N_38554,N_38992);
nor U39209 (N_39209,N_38913,N_38750);
or U39210 (N_39210,N_38929,N_38715);
xor U39211 (N_39211,N_38970,N_38766);
nand U39212 (N_39212,N_38333,N_38565);
nor U39213 (N_39213,N_38933,N_38012);
nand U39214 (N_39214,N_38114,N_38136);
or U39215 (N_39215,N_38347,N_38037);
nand U39216 (N_39216,N_38447,N_38207);
xor U39217 (N_39217,N_38104,N_38841);
or U39218 (N_39218,N_38871,N_38571);
or U39219 (N_39219,N_38485,N_38421);
and U39220 (N_39220,N_38232,N_38587);
or U39221 (N_39221,N_38380,N_38927);
or U39222 (N_39222,N_38112,N_38592);
or U39223 (N_39223,N_38976,N_38199);
and U39224 (N_39224,N_38979,N_38726);
xnor U39225 (N_39225,N_38082,N_38033);
or U39226 (N_39226,N_38325,N_38858);
or U39227 (N_39227,N_38307,N_38007);
and U39228 (N_39228,N_38469,N_38350);
or U39229 (N_39229,N_38453,N_38989);
xnor U39230 (N_39230,N_38689,N_38243);
xor U39231 (N_39231,N_38768,N_38349);
or U39232 (N_39232,N_38942,N_38749);
nor U39233 (N_39233,N_38662,N_38449);
nor U39234 (N_39234,N_38702,N_38966);
and U39235 (N_39235,N_38251,N_38124);
or U39236 (N_39236,N_38000,N_38540);
nor U39237 (N_39237,N_38915,N_38911);
nor U39238 (N_39238,N_38816,N_38861);
nor U39239 (N_39239,N_38121,N_38322);
and U39240 (N_39240,N_38174,N_38917);
or U39241 (N_39241,N_38298,N_38364);
or U39242 (N_39242,N_38148,N_38711);
nand U39243 (N_39243,N_38923,N_38563);
nor U39244 (N_39244,N_38088,N_38414);
nor U39245 (N_39245,N_38391,N_38625);
nand U39246 (N_39246,N_38826,N_38791);
xor U39247 (N_39247,N_38512,N_38430);
xnor U39248 (N_39248,N_38008,N_38077);
and U39249 (N_39249,N_38580,N_38142);
nor U39250 (N_39250,N_38266,N_38003);
or U39251 (N_39251,N_38805,N_38118);
or U39252 (N_39252,N_38940,N_38560);
nor U39253 (N_39253,N_38638,N_38656);
and U39254 (N_39254,N_38047,N_38908);
nand U39255 (N_39255,N_38605,N_38521);
nand U39256 (N_39256,N_38661,N_38496);
xnor U39257 (N_39257,N_38619,N_38423);
or U39258 (N_39258,N_38071,N_38747);
nand U39259 (N_39259,N_38315,N_38804);
nor U39260 (N_39260,N_38029,N_38164);
and U39261 (N_39261,N_38953,N_38495);
and U39262 (N_39262,N_38860,N_38688);
xor U39263 (N_39263,N_38672,N_38237);
and U39264 (N_39264,N_38839,N_38827);
and U39265 (N_39265,N_38010,N_38440);
or U39266 (N_39266,N_38806,N_38410);
and U39267 (N_39267,N_38898,N_38214);
nand U39268 (N_39268,N_38262,N_38716);
nor U39269 (N_39269,N_38467,N_38783);
nor U39270 (N_39270,N_38299,N_38076);
xor U39271 (N_39271,N_38103,N_38065);
nor U39272 (N_39272,N_38557,N_38848);
or U39273 (N_39273,N_38198,N_38832);
and U39274 (N_39274,N_38454,N_38696);
nand U39275 (N_39275,N_38404,N_38509);
nor U39276 (N_39276,N_38110,N_38336);
xnor U39277 (N_39277,N_38398,N_38326);
and U39278 (N_39278,N_38344,N_38308);
nand U39279 (N_39279,N_38674,N_38648);
nand U39280 (N_39280,N_38765,N_38581);
nand U39281 (N_39281,N_38235,N_38479);
nand U39282 (N_39282,N_38654,N_38722);
nand U39283 (N_39283,N_38564,N_38584);
or U39284 (N_39284,N_38939,N_38612);
xor U39285 (N_39285,N_38461,N_38823);
xor U39286 (N_39286,N_38967,N_38481);
or U39287 (N_39287,N_38916,N_38863);
nor U39288 (N_39288,N_38762,N_38697);
or U39289 (N_39289,N_38607,N_38486);
nor U39290 (N_39290,N_38652,N_38191);
nor U39291 (N_39291,N_38773,N_38960);
and U39292 (N_39292,N_38419,N_38621);
xor U39293 (N_39293,N_38338,N_38708);
and U39294 (N_39294,N_38371,N_38426);
nand U39295 (N_39295,N_38876,N_38387);
and U39296 (N_39296,N_38292,N_38400);
nor U39297 (N_39297,N_38320,N_38520);
nand U39298 (N_39298,N_38847,N_38732);
nand U39299 (N_39299,N_38311,N_38628);
and U39300 (N_39300,N_38721,N_38166);
nor U39301 (N_39301,N_38304,N_38201);
or U39302 (N_39302,N_38517,N_38134);
xnor U39303 (N_39303,N_38452,N_38125);
xnor U39304 (N_39304,N_38184,N_38432);
nand U39305 (N_39305,N_38772,N_38339);
and U39306 (N_39306,N_38044,N_38591);
or U39307 (N_39307,N_38609,N_38155);
nor U39308 (N_39308,N_38922,N_38589);
xnor U39309 (N_39309,N_38064,N_38096);
nor U39310 (N_39310,N_38892,N_38217);
nand U39311 (N_39311,N_38365,N_38676);
nand U39312 (N_39312,N_38906,N_38864);
xor U39313 (N_39313,N_38073,N_38309);
nor U39314 (N_39314,N_38300,N_38046);
xor U39315 (N_39315,N_38063,N_38700);
nor U39316 (N_39316,N_38368,N_38663);
or U39317 (N_39317,N_38780,N_38186);
nand U39318 (N_39318,N_38172,N_38126);
nor U39319 (N_39319,N_38328,N_38055);
xnor U39320 (N_39320,N_38129,N_38613);
and U39321 (N_39321,N_38094,N_38819);
xor U39322 (N_39322,N_38808,N_38984);
or U39323 (N_39323,N_38596,N_38023);
nand U39324 (N_39324,N_38585,N_38956);
nor U39325 (N_39325,N_38988,N_38575);
nor U39326 (N_39326,N_38622,N_38644);
or U39327 (N_39327,N_38817,N_38407);
nand U39328 (N_39328,N_38289,N_38987);
nor U39329 (N_39329,N_38699,N_38248);
xor U39330 (N_39330,N_38209,N_38507);
and U39331 (N_39331,N_38703,N_38185);
xor U39332 (N_39332,N_38466,N_38036);
xnor U39333 (N_39333,N_38257,N_38659);
nor U39334 (N_39334,N_38383,N_38603);
and U39335 (N_39335,N_38639,N_38610);
and U39336 (N_39336,N_38786,N_38048);
and U39337 (N_39337,N_38675,N_38070);
xor U39338 (N_39338,N_38794,N_38930);
xor U39339 (N_39339,N_38879,N_38431);
nor U39340 (N_39340,N_38028,N_38079);
xnor U39341 (N_39341,N_38618,N_38218);
nor U39342 (N_39342,N_38617,N_38822);
nor U39343 (N_39343,N_38994,N_38204);
or U39344 (N_39344,N_38355,N_38775);
and U39345 (N_39345,N_38981,N_38895);
or U39346 (N_39346,N_38853,N_38473);
and U39347 (N_39347,N_38925,N_38531);
xnor U39348 (N_39348,N_38634,N_38455);
xnor U39349 (N_39349,N_38153,N_38952);
or U39350 (N_39350,N_38851,N_38223);
nor U39351 (N_39351,N_38995,N_38381);
nor U39352 (N_39352,N_38616,N_38874);
nor U39353 (N_39353,N_38921,N_38083);
nor U39354 (N_39354,N_38329,N_38552);
xnor U39355 (N_39355,N_38950,N_38331);
nor U39356 (N_39356,N_38793,N_38480);
and U39357 (N_39357,N_38801,N_38748);
or U39358 (N_39358,N_38769,N_38964);
xor U39359 (N_39359,N_38545,N_38668);
nor U39360 (N_39360,N_38197,N_38051);
nand U39361 (N_39361,N_38866,N_38208);
nor U39362 (N_39362,N_38193,N_38205);
nor U39363 (N_39363,N_38450,N_38278);
and U39364 (N_39364,N_38541,N_38084);
or U39365 (N_39365,N_38891,N_38878);
nor U39366 (N_39366,N_38733,N_38506);
nor U39367 (N_39367,N_38546,N_38271);
and U39368 (N_39368,N_38588,N_38978);
xor U39369 (N_39369,N_38838,N_38842);
and U39370 (N_39370,N_38901,N_38695);
nand U39371 (N_39371,N_38031,N_38295);
or U39372 (N_39372,N_38490,N_38141);
nor U39373 (N_39373,N_38802,N_38345);
and U39374 (N_39374,N_38754,N_38873);
xor U39375 (N_39375,N_38017,N_38706);
and U39376 (N_39376,N_38650,N_38222);
or U39377 (N_39377,N_38313,N_38014);
or U39378 (N_39378,N_38487,N_38728);
nand U39379 (N_39379,N_38396,N_38286);
xnor U39380 (N_39380,N_38835,N_38934);
nor U39381 (N_39381,N_38870,N_38054);
or U39382 (N_39382,N_38236,N_38796);
xor U39383 (N_39383,N_38508,N_38269);
xor U39384 (N_39384,N_38353,N_38590);
xnor U39385 (N_39385,N_38261,N_38518);
nor U39386 (N_39386,N_38120,N_38746);
xnor U39387 (N_39387,N_38465,N_38814);
nand U39388 (N_39388,N_38441,N_38893);
nand U39389 (N_39389,N_38576,N_38145);
nand U39390 (N_39390,N_38759,N_38305);
xnor U39391 (N_39391,N_38493,N_38282);
or U39392 (N_39392,N_38505,N_38807);
or U39393 (N_39393,N_38335,N_38527);
or U39394 (N_39394,N_38720,N_38062);
nand U39395 (N_39395,N_38438,N_38042);
and U39396 (N_39396,N_38640,N_38402);
nor U39397 (N_39397,N_38740,N_38743);
nand U39398 (N_39398,N_38683,N_38614);
nor U39399 (N_39399,N_38945,N_38993);
nand U39400 (N_39400,N_38090,N_38660);
and U39401 (N_39401,N_38834,N_38677);
xor U39402 (N_39402,N_38343,N_38376);
and U39403 (N_39403,N_38091,N_38150);
xnor U39404 (N_39404,N_38405,N_38763);
xor U39405 (N_39405,N_38139,N_38547);
nand U39406 (N_39406,N_38774,N_38403);
or U39407 (N_39407,N_38448,N_38314);
nand U39408 (N_39408,N_38260,N_38085);
nand U39409 (N_39409,N_38574,N_38206);
and U39410 (N_39410,N_38499,N_38316);
nand U39411 (N_39411,N_38857,N_38408);
nand U39412 (N_39412,N_38936,N_38422);
or U39413 (N_39413,N_38941,N_38980);
or U39414 (N_39414,N_38444,N_38905);
and U39415 (N_39415,N_38013,N_38019);
or U39416 (N_39416,N_38437,N_38067);
and U39417 (N_39417,N_38154,N_38462);
nand U39418 (N_39418,N_38361,N_38854);
nand U39419 (N_39419,N_38290,N_38798);
nor U39420 (N_39420,N_38281,N_38442);
xor U39421 (N_39421,N_38100,N_38287);
and U39422 (N_39422,N_38516,N_38597);
and U39423 (N_39423,N_38559,N_38182);
nand U39424 (N_39424,N_38011,N_38818);
or U39425 (N_39425,N_38550,N_38049);
nor U39426 (N_39426,N_38831,N_38491);
and U39427 (N_39427,N_38357,N_38741);
nor U39428 (N_39428,N_38872,N_38245);
nand U39429 (N_39429,N_38943,N_38991);
nand U39430 (N_39430,N_38157,N_38196);
or U39431 (N_39431,N_38599,N_38714);
or U39432 (N_39432,N_38439,N_38389);
nand U39433 (N_39433,N_38846,N_38569);
or U39434 (N_39434,N_38272,N_38828);
xnor U39435 (N_39435,N_38015,N_38238);
nand U39436 (N_39436,N_38524,N_38231);
nand U39437 (N_39437,N_38362,N_38710);
nand U39438 (N_39438,N_38890,N_38034);
xnor U39439 (N_39439,N_38919,N_38525);
nor U39440 (N_39440,N_38358,N_38032);
or U39441 (N_39441,N_38342,N_38955);
nand U39442 (N_39442,N_38653,N_38551);
nor U39443 (N_39443,N_38666,N_38215);
nand U39444 (N_39444,N_38731,N_38725);
nor U39445 (N_39445,N_38513,N_38997);
or U39446 (N_39446,N_38961,N_38274);
or U39447 (N_39447,N_38027,N_38645);
nand U39448 (N_39448,N_38169,N_38556);
and U39449 (N_39449,N_38240,N_38604);
nand U39450 (N_39450,N_38258,N_38787);
or U39451 (N_39451,N_38195,N_38691);
nand U39452 (N_39452,N_38924,N_38529);
xor U39453 (N_39453,N_38340,N_38687);
nor U39454 (N_39454,N_38039,N_38225);
and U39455 (N_39455,N_38131,N_38938);
or U39456 (N_39456,N_38168,N_38221);
or U39457 (N_39457,N_38562,N_38608);
nand U39458 (N_39458,N_38875,N_38558);
and U39459 (N_39459,N_38156,N_38757);
nor U39460 (N_39460,N_38472,N_38464);
xnor U39461 (N_39461,N_38542,N_38276);
nor U39462 (N_39462,N_38894,N_38456);
xor U39463 (N_39463,N_38664,N_38210);
or U39464 (N_39464,N_38178,N_38230);
nand U39465 (N_39465,N_38411,N_38108);
or U39466 (N_39466,N_38433,N_38799);
nor U39467 (N_39467,N_38897,N_38718);
nor U39468 (N_39468,N_38038,N_38115);
xor U39469 (N_39469,N_38413,N_38784);
xor U39470 (N_39470,N_38969,N_38583);
or U39471 (N_39471,N_38233,N_38771);
and U39472 (N_39472,N_38122,N_38637);
or U39473 (N_39473,N_38781,N_38161);
xor U39474 (N_39474,N_38572,N_38106);
nor U39475 (N_39475,N_38057,N_38742);
nand U39476 (N_39476,N_38177,N_38163);
or U39477 (N_39477,N_38436,N_38867);
and U39478 (N_39478,N_38149,N_38958);
nand U39479 (N_39479,N_38045,N_38321);
and U39480 (N_39480,N_38130,N_38041);
nand U39481 (N_39481,N_38443,N_38132);
or U39482 (N_39482,N_38341,N_38242);
nand U39483 (N_39483,N_38373,N_38020);
or U39484 (N_39484,N_38228,N_38285);
xnor U39485 (N_39485,N_38713,N_38259);
and U39486 (N_39486,N_38241,N_38658);
nand U39487 (N_39487,N_38327,N_38538);
or U39488 (N_39488,N_38384,N_38021);
nand U39489 (N_39489,N_38052,N_38101);
nand U39490 (N_39490,N_38354,N_38176);
nand U39491 (N_39491,N_38825,N_38815);
and U39492 (N_39492,N_38040,N_38372);
nor U39493 (N_39493,N_38445,N_38918);
or U39494 (N_39494,N_38669,N_38075);
xnor U39495 (N_39495,N_38888,N_38907);
or U39496 (N_39496,N_38830,N_38092);
nor U39497 (N_39497,N_38971,N_38914);
nor U39498 (N_39498,N_38779,N_38707);
nor U39499 (N_39499,N_38751,N_38684);
nor U39500 (N_39500,N_38046,N_38100);
nand U39501 (N_39501,N_38948,N_38844);
xnor U39502 (N_39502,N_38406,N_38816);
or U39503 (N_39503,N_38686,N_38589);
nor U39504 (N_39504,N_38356,N_38172);
xor U39505 (N_39505,N_38640,N_38380);
and U39506 (N_39506,N_38292,N_38804);
nor U39507 (N_39507,N_38599,N_38937);
nor U39508 (N_39508,N_38620,N_38859);
xor U39509 (N_39509,N_38456,N_38948);
xnor U39510 (N_39510,N_38821,N_38104);
nand U39511 (N_39511,N_38899,N_38924);
and U39512 (N_39512,N_38424,N_38324);
nor U39513 (N_39513,N_38318,N_38725);
xnor U39514 (N_39514,N_38779,N_38905);
xor U39515 (N_39515,N_38063,N_38078);
nand U39516 (N_39516,N_38530,N_38089);
nand U39517 (N_39517,N_38487,N_38265);
nand U39518 (N_39518,N_38310,N_38738);
nand U39519 (N_39519,N_38133,N_38874);
or U39520 (N_39520,N_38549,N_38819);
xor U39521 (N_39521,N_38170,N_38713);
xor U39522 (N_39522,N_38043,N_38298);
nand U39523 (N_39523,N_38256,N_38585);
nor U39524 (N_39524,N_38450,N_38553);
nor U39525 (N_39525,N_38564,N_38587);
nand U39526 (N_39526,N_38475,N_38940);
or U39527 (N_39527,N_38237,N_38763);
or U39528 (N_39528,N_38175,N_38055);
nor U39529 (N_39529,N_38596,N_38293);
and U39530 (N_39530,N_38030,N_38035);
nor U39531 (N_39531,N_38589,N_38369);
or U39532 (N_39532,N_38172,N_38499);
nand U39533 (N_39533,N_38027,N_38230);
and U39534 (N_39534,N_38622,N_38255);
nor U39535 (N_39535,N_38592,N_38052);
nand U39536 (N_39536,N_38828,N_38985);
and U39537 (N_39537,N_38642,N_38418);
xor U39538 (N_39538,N_38338,N_38680);
nor U39539 (N_39539,N_38526,N_38978);
nor U39540 (N_39540,N_38144,N_38843);
nor U39541 (N_39541,N_38406,N_38143);
nand U39542 (N_39542,N_38070,N_38522);
nor U39543 (N_39543,N_38899,N_38276);
xor U39544 (N_39544,N_38754,N_38367);
xor U39545 (N_39545,N_38931,N_38473);
nor U39546 (N_39546,N_38230,N_38605);
nor U39547 (N_39547,N_38776,N_38337);
xnor U39548 (N_39548,N_38719,N_38140);
nor U39549 (N_39549,N_38901,N_38583);
nor U39550 (N_39550,N_38702,N_38062);
nand U39551 (N_39551,N_38883,N_38665);
nor U39552 (N_39552,N_38137,N_38591);
and U39553 (N_39553,N_38290,N_38067);
or U39554 (N_39554,N_38092,N_38708);
nor U39555 (N_39555,N_38576,N_38265);
nor U39556 (N_39556,N_38422,N_38308);
nor U39557 (N_39557,N_38176,N_38770);
and U39558 (N_39558,N_38743,N_38197);
and U39559 (N_39559,N_38147,N_38733);
xor U39560 (N_39560,N_38390,N_38559);
xor U39561 (N_39561,N_38458,N_38432);
nor U39562 (N_39562,N_38933,N_38940);
nor U39563 (N_39563,N_38165,N_38925);
and U39564 (N_39564,N_38216,N_38806);
or U39565 (N_39565,N_38152,N_38241);
nand U39566 (N_39566,N_38395,N_38810);
or U39567 (N_39567,N_38162,N_38321);
and U39568 (N_39568,N_38264,N_38985);
and U39569 (N_39569,N_38676,N_38857);
or U39570 (N_39570,N_38634,N_38450);
nor U39571 (N_39571,N_38068,N_38700);
xnor U39572 (N_39572,N_38370,N_38773);
nor U39573 (N_39573,N_38304,N_38331);
nor U39574 (N_39574,N_38147,N_38714);
nand U39575 (N_39575,N_38597,N_38342);
nor U39576 (N_39576,N_38085,N_38804);
and U39577 (N_39577,N_38722,N_38451);
or U39578 (N_39578,N_38175,N_38393);
xnor U39579 (N_39579,N_38455,N_38718);
nor U39580 (N_39580,N_38073,N_38226);
or U39581 (N_39581,N_38408,N_38708);
nor U39582 (N_39582,N_38326,N_38922);
xor U39583 (N_39583,N_38818,N_38373);
nand U39584 (N_39584,N_38217,N_38325);
nand U39585 (N_39585,N_38327,N_38303);
nor U39586 (N_39586,N_38568,N_38364);
nor U39587 (N_39587,N_38649,N_38888);
xnor U39588 (N_39588,N_38829,N_38553);
xnor U39589 (N_39589,N_38399,N_38043);
nor U39590 (N_39590,N_38236,N_38204);
and U39591 (N_39591,N_38039,N_38690);
nor U39592 (N_39592,N_38745,N_38716);
xor U39593 (N_39593,N_38169,N_38160);
or U39594 (N_39594,N_38009,N_38255);
or U39595 (N_39595,N_38815,N_38675);
nor U39596 (N_39596,N_38173,N_38674);
nor U39597 (N_39597,N_38877,N_38620);
and U39598 (N_39598,N_38689,N_38428);
nor U39599 (N_39599,N_38796,N_38094);
nor U39600 (N_39600,N_38267,N_38252);
xnor U39601 (N_39601,N_38259,N_38150);
nand U39602 (N_39602,N_38939,N_38173);
nor U39603 (N_39603,N_38377,N_38019);
xor U39604 (N_39604,N_38883,N_38888);
or U39605 (N_39605,N_38910,N_38714);
nand U39606 (N_39606,N_38799,N_38684);
and U39607 (N_39607,N_38699,N_38185);
or U39608 (N_39608,N_38608,N_38855);
nor U39609 (N_39609,N_38544,N_38220);
xor U39610 (N_39610,N_38874,N_38271);
nand U39611 (N_39611,N_38810,N_38516);
nor U39612 (N_39612,N_38817,N_38814);
nand U39613 (N_39613,N_38114,N_38140);
and U39614 (N_39614,N_38952,N_38861);
nand U39615 (N_39615,N_38564,N_38458);
and U39616 (N_39616,N_38744,N_38183);
nor U39617 (N_39617,N_38232,N_38373);
nand U39618 (N_39618,N_38074,N_38446);
nor U39619 (N_39619,N_38277,N_38839);
or U39620 (N_39620,N_38046,N_38317);
xor U39621 (N_39621,N_38875,N_38959);
xnor U39622 (N_39622,N_38792,N_38602);
nor U39623 (N_39623,N_38921,N_38793);
or U39624 (N_39624,N_38023,N_38665);
or U39625 (N_39625,N_38409,N_38896);
nor U39626 (N_39626,N_38392,N_38033);
xor U39627 (N_39627,N_38817,N_38564);
xnor U39628 (N_39628,N_38335,N_38571);
nor U39629 (N_39629,N_38317,N_38933);
nor U39630 (N_39630,N_38790,N_38813);
and U39631 (N_39631,N_38874,N_38031);
and U39632 (N_39632,N_38422,N_38652);
and U39633 (N_39633,N_38463,N_38083);
nor U39634 (N_39634,N_38184,N_38259);
and U39635 (N_39635,N_38167,N_38605);
nand U39636 (N_39636,N_38333,N_38751);
and U39637 (N_39637,N_38578,N_38979);
and U39638 (N_39638,N_38194,N_38392);
and U39639 (N_39639,N_38052,N_38716);
or U39640 (N_39640,N_38393,N_38542);
nand U39641 (N_39641,N_38326,N_38672);
and U39642 (N_39642,N_38915,N_38024);
or U39643 (N_39643,N_38023,N_38781);
and U39644 (N_39644,N_38312,N_38131);
and U39645 (N_39645,N_38864,N_38712);
xnor U39646 (N_39646,N_38437,N_38896);
xor U39647 (N_39647,N_38510,N_38866);
xnor U39648 (N_39648,N_38987,N_38460);
or U39649 (N_39649,N_38369,N_38235);
nand U39650 (N_39650,N_38593,N_38241);
xor U39651 (N_39651,N_38042,N_38851);
and U39652 (N_39652,N_38871,N_38138);
xnor U39653 (N_39653,N_38446,N_38763);
or U39654 (N_39654,N_38748,N_38983);
nor U39655 (N_39655,N_38646,N_38308);
or U39656 (N_39656,N_38513,N_38563);
or U39657 (N_39657,N_38035,N_38855);
nand U39658 (N_39658,N_38518,N_38060);
or U39659 (N_39659,N_38191,N_38545);
nor U39660 (N_39660,N_38741,N_38851);
and U39661 (N_39661,N_38466,N_38828);
or U39662 (N_39662,N_38288,N_38890);
xnor U39663 (N_39663,N_38903,N_38291);
xnor U39664 (N_39664,N_38753,N_38011);
nand U39665 (N_39665,N_38998,N_38977);
nor U39666 (N_39666,N_38650,N_38371);
nand U39667 (N_39667,N_38391,N_38716);
and U39668 (N_39668,N_38787,N_38210);
and U39669 (N_39669,N_38061,N_38539);
and U39670 (N_39670,N_38042,N_38421);
xnor U39671 (N_39671,N_38862,N_38141);
xor U39672 (N_39672,N_38753,N_38264);
nand U39673 (N_39673,N_38451,N_38265);
nor U39674 (N_39674,N_38495,N_38113);
xnor U39675 (N_39675,N_38557,N_38679);
nor U39676 (N_39676,N_38614,N_38585);
nor U39677 (N_39677,N_38846,N_38295);
or U39678 (N_39678,N_38816,N_38518);
nor U39679 (N_39679,N_38927,N_38867);
nand U39680 (N_39680,N_38642,N_38868);
or U39681 (N_39681,N_38116,N_38939);
nand U39682 (N_39682,N_38624,N_38496);
xnor U39683 (N_39683,N_38708,N_38838);
or U39684 (N_39684,N_38469,N_38810);
nand U39685 (N_39685,N_38130,N_38148);
nor U39686 (N_39686,N_38822,N_38517);
nand U39687 (N_39687,N_38940,N_38804);
nor U39688 (N_39688,N_38062,N_38672);
and U39689 (N_39689,N_38334,N_38998);
nand U39690 (N_39690,N_38693,N_38831);
and U39691 (N_39691,N_38377,N_38077);
xor U39692 (N_39692,N_38195,N_38849);
nor U39693 (N_39693,N_38767,N_38702);
nor U39694 (N_39694,N_38983,N_38692);
and U39695 (N_39695,N_38415,N_38147);
xor U39696 (N_39696,N_38549,N_38535);
nand U39697 (N_39697,N_38794,N_38945);
xor U39698 (N_39698,N_38808,N_38591);
and U39699 (N_39699,N_38059,N_38051);
and U39700 (N_39700,N_38927,N_38134);
nand U39701 (N_39701,N_38374,N_38224);
nand U39702 (N_39702,N_38918,N_38409);
xor U39703 (N_39703,N_38974,N_38748);
nor U39704 (N_39704,N_38752,N_38530);
nand U39705 (N_39705,N_38063,N_38367);
nor U39706 (N_39706,N_38281,N_38782);
and U39707 (N_39707,N_38735,N_38209);
nor U39708 (N_39708,N_38547,N_38404);
and U39709 (N_39709,N_38511,N_38746);
nor U39710 (N_39710,N_38117,N_38818);
nand U39711 (N_39711,N_38860,N_38260);
nand U39712 (N_39712,N_38041,N_38970);
and U39713 (N_39713,N_38975,N_38513);
nand U39714 (N_39714,N_38072,N_38467);
or U39715 (N_39715,N_38247,N_38121);
nor U39716 (N_39716,N_38625,N_38640);
xor U39717 (N_39717,N_38590,N_38204);
and U39718 (N_39718,N_38268,N_38384);
nand U39719 (N_39719,N_38567,N_38515);
or U39720 (N_39720,N_38968,N_38028);
or U39721 (N_39721,N_38465,N_38260);
or U39722 (N_39722,N_38246,N_38544);
nor U39723 (N_39723,N_38375,N_38494);
or U39724 (N_39724,N_38970,N_38220);
and U39725 (N_39725,N_38765,N_38345);
and U39726 (N_39726,N_38731,N_38026);
or U39727 (N_39727,N_38523,N_38726);
nor U39728 (N_39728,N_38530,N_38781);
nand U39729 (N_39729,N_38411,N_38868);
xor U39730 (N_39730,N_38727,N_38463);
and U39731 (N_39731,N_38579,N_38403);
nor U39732 (N_39732,N_38696,N_38016);
or U39733 (N_39733,N_38485,N_38014);
and U39734 (N_39734,N_38655,N_38638);
xnor U39735 (N_39735,N_38565,N_38875);
nor U39736 (N_39736,N_38291,N_38100);
or U39737 (N_39737,N_38811,N_38450);
nand U39738 (N_39738,N_38667,N_38591);
nand U39739 (N_39739,N_38640,N_38864);
nor U39740 (N_39740,N_38455,N_38275);
xnor U39741 (N_39741,N_38088,N_38527);
and U39742 (N_39742,N_38776,N_38336);
xnor U39743 (N_39743,N_38216,N_38926);
or U39744 (N_39744,N_38168,N_38556);
xor U39745 (N_39745,N_38361,N_38482);
and U39746 (N_39746,N_38454,N_38374);
or U39747 (N_39747,N_38765,N_38012);
xnor U39748 (N_39748,N_38093,N_38471);
and U39749 (N_39749,N_38116,N_38720);
nor U39750 (N_39750,N_38142,N_38567);
nand U39751 (N_39751,N_38932,N_38705);
and U39752 (N_39752,N_38617,N_38008);
nor U39753 (N_39753,N_38206,N_38113);
or U39754 (N_39754,N_38237,N_38245);
nor U39755 (N_39755,N_38080,N_38707);
nand U39756 (N_39756,N_38088,N_38958);
xnor U39757 (N_39757,N_38979,N_38824);
nand U39758 (N_39758,N_38533,N_38511);
xor U39759 (N_39759,N_38023,N_38544);
xnor U39760 (N_39760,N_38830,N_38792);
xor U39761 (N_39761,N_38292,N_38484);
nand U39762 (N_39762,N_38924,N_38420);
xor U39763 (N_39763,N_38448,N_38163);
nor U39764 (N_39764,N_38094,N_38597);
or U39765 (N_39765,N_38134,N_38200);
or U39766 (N_39766,N_38863,N_38384);
and U39767 (N_39767,N_38499,N_38804);
nand U39768 (N_39768,N_38675,N_38501);
nor U39769 (N_39769,N_38798,N_38192);
xnor U39770 (N_39770,N_38628,N_38091);
nor U39771 (N_39771,N_38676,N_38077);
nand U39772 (N_39772,N_38453,N_38283);
or U39773 (N_39773,N_38607,N_38166);
xor U39774 (N_39774,N_38925,N_38409);
nand U39775 (N_39775,N_38929,N_38713);
nor U39776 (N_39776,N_38469,N_38629);
or U39777 (N_39777,N_38265,N_38642);
or U39778 (N_39778,N_38252,N_38012);
nand U39779 (N_39779,N_38465,N_38873);
nor U39780 (N_39780,N_38692,N_38652);
or U39781 (N_39781,N_38062,N_38423);
nor U39782 (N_39782,N_38282,N_38425);
and U39783 (N_39783,N_38032,N_38555);
or U39784 (N_39784,N_38377,N_38614);
nand U39785 (N_39785,N_38263,N_38198);
nand U39786 (N_39786,N_38182,N_38602);
or U39787 (N_39787,N_38461,N_38749);
or U39788 (N_39788,N_38060,N_38415);
xnor U39789 (N_39789,N_38499,N_38123);
or U39790 (N_39790,N_38716,N_38498);
and U39791 (N_39791,N_38983,N_38121);
or U39792 (N_39792,N_38478,N_38692);
nor U39793 (N_39793,N_38543,N_38590);
or U39794 (N_39794,N_38810,N_38050);
nand U39795 (N_39795,N_38736,N_38824);
or U39796 (N_39796,N_38125,N_38150);
nand U39797 (N_39797,N_38832,N_38910);
nor U39798 (N_39798,N_38848,N_38659);
nand U39799 (N_39799,N_38052,N_38440);
and U39800 (N_39800,N_38732,N_38475);
nor U39801 (N_39801,N_38719,N_38102);
nand U39802 (N_39802,N_38515,N_38778);
nor U39803 (N_39803,N_38907,N_38339);
nand U39804 (N_39804,N_38241,N_38249);
or U39805 (N_39805,N_38337,N_38511);
or U39806 (N_39806,N_38131,N_38223);
nand U39807 (N_39807,N_38148,N_38493);
and U39808 (N_39808,N_38999,N_38364);
or U39809 (N_39809,N_38240,N_38875);
nor U39810 (N_39810,N_38927,N_38761);
and U39811 (N_39811,N_38315,N_38885);
xor U39812 (N_39812,N_38929,N_38107);
nor U39813 (N_39813,N_38710,N_38396);
nor U39814 (N_39814,N_38383,N_38691);
xnor U39815 (N_39815,N_38203,N_38490);
nor U39816 (N_39816,N_38352,N_38282);
xor U39817 (N_39817,N_38594,N_38065);
or U39818 (N_39818,N_38595,N_38768);
or U39819 (N_39819,N_38316,N_38256);
nor U39820 (N_39820,N_38260,N_38354);
and U39821 (N_39821,N_38134,N_38155);
and U39822 (N_39822,N_38633,N_38042);
xnor U39823 (N_39823,N_38015,N_38089);
or U39824 (N_39824,N_38364,N_38326);
nor U39825 (N_39825,N_38230,N_38231);
xnor U39826 (N_39826,N_38003,N_38894);
nand U39827 (N_39827,N_38766,N_38015);
or U39828 (N_39828,N_38661,N_38854);
nor U39829 (N_39829,N_38809,N_38978);
nand U39830 (N_39830,N_38373,N_38708);
nand U39831 (N_39831,N_38408,N_38942);
nor U39832 (N_39832,N_38031,N_38319);
or U39833 (N_39833,N_38201,N_38736);
nor U39834 (N_39834,N_38224,N_38346);
nand U39835 (N_39835,N_38058,N_38299);
nor U39836 (N_39836,N_38444,N_38549);
nand U39837 (N_39837,N_38531,N_38929);
xor U39838 (N_39838,N_38343,N_38654);
and U39839 (N_39839,N_38398,N_38632);
and U39840 (N_39840,N_38267,N_38869);
nand U39841 (N_39841,N_38505,N_38200);
xnor U39842 (N_39842,N_38815,N_38220);
nand U39843 (N_39843,N_38739,N_38785);
nor U39844 (N_39844,N_38026,N_38829);
nand U39845 (N_39845,N_38184,N_38360);
and U39846 (N_39846,N_38272,N_38222);
and U39847 (N_39847,N_38073,N_38554);
nand U39848 (N_39848,N_38364,N_38877);
and U39849 (N_39849,N_38287,N_38447);
or U39850 (N_39850,N_38677,N_38305);
and U39851 (N_39851,N_38018,N_38678);
xnor U39852 (N_39852,N_38941,N_38091);
and U39853 (N_39853,N_38947,N_38797);
nand U39854 (N_39854,N_38242,N_38302);
xnor U39855 (N_39855,N_38977,N_38687);
xnor U39856 (N_39856,N_38554,N_38389);
nor U39857 (N_39857,N_38048,N_38078);
xnor U39858 (N_39858,N_38200,N_38282);
and U39859 (N_39859,N_38438,N_38512);
or U39860 (N_39860,N_38687,N_38643);
and U39861 (N_39861,N_38368,N_38275);
nor U39862 (N_39862,N_38040,N_38248);
and U39863 (N_39863,N_38221,N_38361);
and U39864 (N_39864,N_38534,N_38028);
or U39865 (N_39865,N_38966,N_38605);
and U39866 (N_39866,N_38498,N_38674);
nand U39867 (N_39867,N_38527,N_38821);
and U39868 (N_39868,N_38149,N_38254);
or U39869 (N_39869,N_38678,N_38338);
xnor U39870 (N_39870,N_38379,N_38200);
nor U39871 (N_39871,N_38460,N_38267);
or U39872 (N_39872,N_38497,N_38032);
and U39873 (N_39873,N_38613,N_38644);
and U39874 (N_39874,N_38775,N_38154);
nand U39875 (N_39875,N_38969,N_38832);
xor U39876 (N_39876,N_38192,N_38029);
nor U39877 (N_39877,N_38468,N_38554);
xnor U39878 (N_39878,N_38944,N_38438);
or U39879 (N_39879,N_38803,N_38271);
and U39880 (N_39880,N_38131,N_38464);
nand U39881 (N_39881,N_38571,N_38123);
nand U39882 (N_39882,N_38364,N_38249);
or U39883 (N_39883,N_38862,N_38305);
and U39884 (N_39884,N_38544,N_38860);
xor U39885 (N_39885,N_38531,N_38240);
or U39886 (N_39886,N_38498,N_38126);
or U39887 (N_39887,N_38294,N_38614);
nor U39888 (N_39888,N_38358,N_38204);
nor U39889 (N_39889,N_38911,N_38579);
or U39890 (N_39890,N_38588,N_38019);
xnor U39891 (N_39891,N_38573,N_38020);
nor U39892 (N_39892,N_38000,N_38408);
nand U39893 (N_39893,N_38261,N_38152);
nand U39894 (N_39894,N_38250,N_38498);
nor U39895 (N_39895,N_38298,N_38799);
or U39896 (N_39896,N_38683,N_38298);
or U39897 (N_39897,N_38507,N_38357);
or U39898 (N_39898,N_38515,N_38680);
nand U39899 (N_39899,N_38728,N_38312);
or U39900 (N_39900,N_38670,N_38243);
and U39901 (N_39901,N_38728,N_38746);
nand U39902 (N_39902,N_38314,N_38775);
and U39903 (N_39903,N_38622,N_38349);
nor U39904 (N_39904,N_38743,N_38570);
nand U39905 (N_39905,N_38413,N_38811);
or U39906 (N_39906,N_38168,N_38605);
xnor U39907 (N_39907,N_38812,N_38765);
nor U39908 (N_39908,N_38209,N_38929);
nor U39909 (N_39909,N_38010,N_38215);
nand U39910 (N_39910,N_38145,N_38326);
nor U39911 (N_39911,N_38859,N_38819);
nand U39912 (N_39912,N_38922,N_38232);
and U39913 (N_39913,N_38738,N_38831);
nand U39914 (N_39914,N_38547,N_38271);
and U39915 (N_39915,N_38938,N_38712);
nand U39916 (N_39916,N_38415,N_38162);
nand U39917 (N_39917,N_38582,N_38070);
or U39918 (N_39918,N_38287,N_38261);
xnor U39919 (N_39919,N_38988,N_38349);
nand U39920 (N_39920,N_38895,N_38815);
nor U39921 (N_39921,N_38979,N_38862);
nor U39922 (N_39922,N_38172,N_38381);
xnor U39923 (N_39923,N_38592,N_38084);
and U39924 (N_39924,N_38043,N_38663);
or U39925 (N_39925,N_38907,N_38858);
or U39926 (N_39926,N_38742,N_38678);
nor U39927 (N_39927,N_38486,N_38241);
xor U39928 (N_39928,N_38363,N_38301);
or U39929 (N_39929,N_38610,N_38375);
xor U39930 (N_39930,N_38516,N_38917);
nor U39931 (N_39931,N_38988,N_38744);
xnor U39932 (N_39932,N_38551,N_38597);
and U39933 (N_39933,N_38780,N_38038);
or U39934 (N_39934,N_38589,N_38940);
nor U39935 (N_39935,N_38969,N_38239);
and U39936 (N_39936,N_38803,N_38502);
or U39937 (N_39937,N_38371,N_38741);
nor U39938 (N_39938,N_38699,N_38387);
and U39939 (N_39939,N_38799,N_38758);
nor U39940 (N_39940,N_38334,N_38134);
and U39941 (N_39941,N_38553,N_38539);
or U39942 (N_39942,N_38345,N_38058);
nand U39943 (N_39943,N_38996,N_38459);
nand U39944 (N_39944,N_38285,N_38005);
xor U39945 (N_39945,N_38885,N_38894);
nand U39946 (N_39946,N_38351,N_38204);
xor U39947 (N_39947,N_38863,N_38057);
nand U39948 (N_39948,N_38585,N_38264);
nand U39949 (N_39949,N_38470,N_38891);
nor U39950 (N_39950,N_38521,N_38657);
nand U39951 (N_39951,N_38588,N_38516);
nor U39952 (N_39952,N_38774,N_38084);
or U39953 (N_39953,N_38363,N_38115);
nor U39954 (N_39954,N_38417,N_38511);
and U39955 (N_39955,N_38101,N_38473);
nor U39956 (N_39956,N_38730,N_38106);
xor U39957 (N_39957,N_38823,N_38803);
or U39958 (N_39958,N_38647,N_38294);
xnor U39959 (N_39959,N_38610,N_38128);
or U39960 (N_39960,N_38619,N_38898);
or U39961 (N_39961,N_38766,N_38569);
nor U39962 (N_39962,N_38936,N_38146);
or U39963 (N_39963,N_38153,N_38605);
and U39964 (N_39964,N_38929,N_38603);
nand U39965 (N_39965,N_38495,N_38419);
or U39966 (N_39966,N_38937,N_38910);
and U39967 (N_39967,N_38005,N_38851);
and U39968 (N_39968,N_38146,N_38725);
nor U39969 (N_39969,N_38843,N_38024);
nor U39970 (N_39970,N_38894,N_38732);
nand U39971 (N_39971,N_38525,N_38641);
nor U39972 (N_39972,N_38859,N_38115);
or U39973 (N_39973,N_38914,N_38583);
xnor U39974 (N_39974,N_38270,N_38090);
xor U39975 (N_39975,N_38987,N_38015);
nor U39976 (N_39976,N_38071,N_38384);
nor U39977 (N_39977,N_38468,N_38264);
nor U39978 (N_39978,N_38033,N_38047);
or U39979 (N_39979,N_38761,N_38311);
or U39980 (N_39980,N_38330,N_38831);
or U39981 (N_39981,N_38802,N_38573);
nor U39982 (N_39982,N_38029,N_38391);
nand U39983 (N_39983,N_38145,N_38920);
nand U39984 (N_39984,N_38160,N_38060);
nor U39985 (N_39985,N_38397,N_38777);
or U39986 (N_39986,N_38850,N_38653);
or U39987 (N_39987,N_38633,N_38793);
nand U39988 (N_39988,N_38845,N_38763);
nand U39989 (N_39989,N_38058,N_38220);
and U39990 (N_39990,N_38800,N_38381);
and U39991 (N_39991,N_38292,N_38467);
nor U39992 (N_39992,N_38086,N_38361);
xnor U39993 (N_39993,N_38375,N_38565);
nor U39994 (N_39994,N_38975,N_38875);
or U39995 (N_39995,N_38457,N_38715);
or U39996 (N_39996,N_38118,N_38293);
and U39997 (N_39997,N_38573,N_38867);
nor U39998 (N_39998,N_38189,N_38634);
nor U39999 (N_39999,N_38022,N_38729);
nor U40000 (N_40000,N_39208,N_39706);
and U40001 (N_40001,N_39891,N_39227);
nor U40002 (N_40002,N_39164,N_39549);
nand U40003 (N_40003,N_39187,N_39550);
nor U40004 (N_40004,N_39845,N_39289);
nor U40005 (N_40005,N_39688,N_39517);
nand U40006 (N_40006,N_39580,N_39356);
nand U40007 (N_40007,N_39631,N_39016);
nor U40008 (N_40008,N_39717,N_39430);
nor U40009 (N_40009,N_39235,N_39104);
or U40010 (N_40010,N_39018,N_39751);
or U40011 (N_40011,N_39553,N_39163);
nor U40012 (N_40012,N_39593,N_39440);
and U40013 (N_40013,N_39438,N_39852);
nor U40014 (N_40014,N_39303,N_39800);
xor U40015 (N_40015,N_39762,N_39282);
nand U40016 (N_40016,N_39527,N_39510);
or U40017 (N_40017,N_39536,N_39474);
xnor U40018 (N_40018,N_39779,N_39721);
xor U40019 (N_40019,N_39903,N_39774);
or U40020 (N_40020,N_39743,N_39153);
or U40021 (N_40021,N_39613,N_39497);
and U40022 (N_40022,N_39341,N_39127);
and U40023 (N_40023,N_39649,N_39677);
and U40024 (N_40024,N_39606,N_39283);
xnor U40025 (N_40025,N_39477,N_39511);
xnor U40026 (N_40026,N_39548,N_39736);
and U40027 (N_40027,N_39874,N_39417);
or U40028 (N_40028,N_39067,N_39128);
xnor U40029 (N_40029,N_39376,N_39133);
nor U40030 (N_40030,N_39911,N_39772);
xor U40031 (N_40031,N_39698,N_39884);
nand U40032 (N_40032,N_39966,N_39795);
nor U40033 (N_40033,N_39419,N_39509);
xnor U40034 (N_40034,N_39111,N_39421);
and U40035 (N_40035,N_39730,N_39693);
and U40036 (N_40036,N_39820,N_39702);
nand U40037 (N_40037,N_39882,N_39997);
and U40038 (N_40038,N_39784,N_39264);
nand U40039 (N_40039,N_39337,N_39821);
xor U40040 (N_40040,N_39375,N_39562);
and U40041 (N_40041,N_39292,N_39589);
nand U40042 (N_40042,N_39240,N_39000);
and U40043 (N_40043,N_39718,N_39723);
or U40044 (N_40044,N_39359,N_39213);
and U40045 (N_40045,N_39501,N_39389);
nand U40046 (N_40046,N_39662,N_39678);
nand U40047 (N_40047,N_39447,N_39045);
nand U40048 (N_40048,N_39500,N_39099);
or U40049 (N_40049,N_39687,N_39014);
and U40050 (N_40050,N_39528,N_39707);
or U40051 (N_40051,N_39719,N_39373);
xnor U40052 (N_40052,N_39735,N_39568);
xnor U40053 (N_40053,N_39670,N_39770);
nand U40054 (N_40054,N_39973,N_39219);
nand U40055 (N_40055,N_39886,N_39675);
xnor U40056 (N_40056,N_39142,N_39609);
nor U40057 (N_40057,N_39679,N_39652);
nor U40058 (N_40058,N_39034,N_39027);
or U40059 (N_40059,N_39722,N_39291);
or U40060 (N_40060,N_39617,N_39334);
and U40061 (N_40061,N_39584,N_39007);
nor U40062 (N_40062,N_39600,N_39725);
xnor U40063 (N_40063,N_39185,N_39752);
or U40064 (N_40064,N_39004,N_39559);
or U40065 (N_40065,N_39308,N_39244);
and U40066 (N_40066,N_39854,N_39771);
and U40067 (N_40067,N_39392,N_39293);
xnor U40068 (N_40068,N_39801,N_39551);
nor U40069 (N_40069,N_39827,N_39573);
nor U40070 (N_40070,N_39407,N_39340);
nor U40071 (N_40071,N_39529,N_39778);
xor U40072 (N_40072,N_39790,N_39435);
and U40073 (N_40073,N_39567,N_39656);
or U40074 (N_40074,N_39913,N_39413);
or U40075 (N_40075,N_39462,N_39676);
xor U40076 (N_40076,N_39304,N_39794);
or U40077 (N_40077,N_39547,N_39898);
xnor U40078 (N_40078,N_39479,N_39313);
or U40079 (N_40079,N_39959,N_39864);
xnor U40080 (N_40080,N_39348,N_39483);
nor U40081 (N_40081,N_39563,N_39616);
xor U40082 (N_40082,N_39942,N_39165);
nand U40083 (N_40083,N_39076,N_39701);
and U40084 (N_40084,N_39871,N_39653);
or U40085 (N_40085,N_39082,N_39860);
or U40086 (N_40086,N_39121,N_39427);
xor U40087 (N_40087,N_39460,N_39829);
and U40088 (N_40088,N_39011,N_39089);
nor U40089 (N_40089,N_39019,N_39039);
or U40090 (N_40090,N_39126,N_39060);
or U40091 (N_40091,N_39144,N_39729);
xor U40092 (N_40092,N_39062,N_39250);
nor U40093 (N_40093,N_39176,N_39120);
nor U40094 (N_40094,N_39320,N_39644);
and U40095 (N_40095,N_39754,N_39070);
nand U40096 (N_40096,N_39482,N_39040);
xnor U40097 (N_40097,N_39423,N_39229);
and U40098 (N_40098,N_39443,N_39488);
or U40099 (N_40099,N_39628,N_39198);
or U40100 (N_40100,N_39967,N_39484);
xnor U40101 (N_40101,N_39444,N_39792);
or U40102 (N_40102,N_39934,N_39422);
nor U40103 (N_40103,N_39110,N_39808);
or U40104 (N_40104,N_39352,N_39668);
or U40105 (N_40105,N_39416,N_39734);
nor U40106 (N_40106,N_39543,N_39713);
and U40107 (N_40107,N_39639,N_39646);
xor U40108 (N_40108,N_39806,N_39057);
nor U40109 (N_40109,N_39494,N_39921);
nand U40110 (N_40110,N_39078,N_39931);
or U40111 (N_40111,N_39941,N_39759);
and U40112 (N_40112,N_39755,N_39115);
and U40113 (N_40113,N_39247,N_39393);
nor U40114 (N_40114,N_39385,N_39519);
and U40115 (N_40115,N_39432,N_39377);
nor U40116 (N_40116,N_39683,N_39892);
nor U40117 (N_40117,N_39516,N_39332);
xor U40118 (N_40118,N_39270,N_39611);
nor U40119 (N_40119,N_39175,N_39763);
xnor U40120 (N_40120,N_39271,N_39180);
xor U40121 (N_40121,N_39715,N_39703);
nand U40122 (N_40122,N_39306,N_39807);
or U40123 (N_40123,N_39437,N_39284);
or U40124 (N_40124,N_39002,N_39347);
nand U40125 (N_40125,N_39411,N_39712);
and U40126 (N_40126,N_39161,N_39281);
nand U40127 (N_40127,N_39415,N_39531);
or U40128 (N_40128,N_39990,N_39301);
xor U40129 (N_40129,N_39615,N_39674);
and U40130 (N_40130,N_39895,N_39956);
xnor U40131 (N_40131,N_39542,N_39075);
and U40132 (N_40132,N_39887,N_39358);
and U40133 (N_40133,N_39094,N_39026);
nand U40134 (N_40134,N_39445,N_39748);
nor U40135 (N_40135,N_39624,N_39579);
and U40136 (N_40136,N_39449,N_39414);
and U40137 (N_40137,N_39731,N_39962);
nor U40138 (N_40138,N_39824,N_39107);
nor U40139 (N_40139,N_39626,N_39345);
nand U40140 (N_40140,N_39455,N_39321);
nor U40141 (N_40141,N_39979,N_39614);
or U40142 (N_40142,N_39077,N_39470);
and U40143 (N_40143,N_39370,N_39836);
and U40144 (N_40144,N_39588,N_39192);
nand U40145 (N_40145,N_39109,N_39069);
xor U40146 (N_40146,N_39681,N_39645);
nand U40147 (N_40147,N_39196,N_39881);
nor U40148 (N_40148,N_39409,N_39556);
nor U40149 (N_40149,N_39124,N_39028);
nor U40150 (N_40150,N_39410,N_39080);
nor U40151 (N_40151,N_39158,N_39506);
and U40152 (N_40152,N_39051,N_39135);
nand U40153 (N_40153,N_39200,N_39159);
xnor U40154 (N_40154,N_39780,N_39276);
or U40155 (N_40155,N_39571,N_39318);
nor U40156 (N_40156,N_39487,N_39918);
and U40157 (N_40157,N_39908,N_39711);
nand U40158 (N_40158,N_39975,N_39946);
and U40159 (N_40159,N_39418,N_39193);
or U40160 (N_40160,N_39178,N_39812);
or U40161 (N_40161,N_39914,N_39042);
and U40162 (N_40162,N_39514,N_39714);
nand U40163 (N_40163,N_39184,N_39983);
xnor U40164 (N_40164,N_39765,N_39296);
nor U40165 (N_40165,N_39572,N_39541);
and U40166 (N_40166,N_39114,N_39189);
nand U40167 (N_40167,N_39183,N_39637);
nand U40168 (N_40168,N_39813,N_39117);
and U40169 (N_40169,N_39540,N_39793);
or U40170 (N_40170,N_39096,N_39238);
or U40171 (N_40171,N_39333,N_39464);
or U40172 (N_40172,N_39442,N_39869);
xor U40173 (N_40173,N_39401,N_39535);
or U40174 (N_40174,N_39204,N_39904);
and U40175 (N_40175,N_39275,N_39379);
xor U40176 (N_40176,N_39512,N_39651);
nand U40177 (N_40177,N_39576,N_39929);
xor U40178 (N_40178,N_39317,N_39634);
xnor U40179 (N_40179,N_39930,N_39181);
nand U40180 (N_40180,N_39149,N_39230);
or U40181 (N_40181,N_39953,N_39945);
nor U40182 (N_40182,N_39169,N_39658);
nor U40183 (N_40183,N_39322,N_39922);
and U40184 (N_40184,N_39650,N_39188);
or U40185 (N_40185,N_39545,N_39750);
and U40186 (N_40186,N_39134,N_39330);
nand U40187 (N_40187,N_39598,N_39367);
nand U40188 (N_40188,N_39587,N_39724);
or U40189 (N_40189,N_39037,N_39902);
nand U40190 (N_40190,N_39056,N_39091);
or U40191 (N_40191,N_39819,N_39520);
or U40192 (N_40192,N_39992,N_39157);
xnor U40193 (N_40193,N_39672,N_39234);
xnor U40194 (N_40194,N_39809,N_39307);
xor U40195 (N_40195,N_39205,N_39690);
nor U40196 (N_40196,N_39804,N_39980);
xnor U40197 (N_40197,N_39335,N_39280);
and U40198 (N_40198,N_39534,N_39129);
or U40199 (N_40199,N_39300,N_39465);
nor U40200 (N_40200,N_39459,N_39074);
nand U40201 (N_40201,N_39206,N_39025);
and U40202 (N_40202,N_39108,N_39673);
nor U40203 (N_40203,N_39311,N_39704);
nand U40204 (N_40204,N_39262,N_39597);
nor U40205 (N_40205,N_39171,N_39825);
nor U40206 (N_40206,N_39896,N_39977);
nor U40207 (N_40207,N_39994,N_39428);
or U40208 (N_40208,N_39602,N_39081);
xnor U40209 (N_40209,N_39601,N_39210);
xnor U40210 (N_40210,N_39446,N_39403);
nand U40211 (N_40211,N_39917,N_39831);
and U40212 (N_40212,N_39822,N_39139);
and U40213 (N_40213,N_39105,N_39486);
xor U40214 (N_40214,N_39302,N_39998);
nor U40215 (N_40215,N_39228,N_39346);
xor U40216 (N_40216,N_39102,N_39397);
and U40217 (N_40217,N_39739,N_39065);
and U40218 (N_40218,N_39740,N_39252);
and U40219 (N_40219,N_39399,N_39682);
and U40220 (N_40220,N_39978,N_39453);
xor U40221 (N_40221,N_39851,N_39505);
or U40222 (N_40222,N_39441,N_39315);
nor U40223 (N_40223,N_39325,N_39369);
nor U40224 (N_40224,N_39787,N_39231);
nor U40225 (N_40225,N_39761,N_39591);
nand U40226 (N_40226,N_39521,N_39297);
or U40227 (N_40227,N_39919,N_39518);
xnor U40228 (N_40228,N_39880,N_39136);
xnor U40229 (N_40229,N_39044,N_39802);
nand U40230 (N_40230,N_39555,N_39585);
and U40231 (N_40231,N_39380,N_39068);
xor U40232 (N_40232,N_39888,N_39118);
nor U40233 (N_40233,N_39872,N_39522);
and U40234 (N_40234,N_39850,N_39849);
nor U40235 (N_40235,N_39909,N_39156);
and U40236 (N_40236,N_39491,N_39485);
nand U40237 (N_40237,N_39982,N_39424);
nand U40238 (N_40238,N_39097,N_39863);
nand U40239 (N_40239,N_39939,N_39101);
nand U40240 (N_40240,N_39691,N_39298);
and U40241 (N_40241,N_39843,N_39781);
or U40242 (N_40242,N_39728,N_39661);
nor U40243 (N_40243,N_39249,N_39530);
xor U40244 (N_40244,N_39476,N_39457);
nor U40245 (N_40245,N_39876,N_39191);
or U40246 (N_40246,N_39396,N_39561);
nor U40247 (N_40247,N_39710,N_39893);
xor U40248 (N_40248,N_39757,N_39995);
nand U40249 (N_40249,N_39524,N_39390);
or U40250 (N_40250,N_39371,N_39776);
nand U40251 (N_40251,N_39894,N_39857);
and U40252 (N_40252,N_39190,N_39439);
xor U40253 (N_40253,N_39867,N_39243);
nor U40254 (N_40254,N_39148,N_39630);
or U40255 (N_40255,N_39935,N_39404);
or U40256 (N_40256,N_39203,N_39268);
nor U40257 (N_40257,N_39883,N_39013);
and U40258 (N_40258,N_39586,N_39504);
nor U40259 (N_40259,N_39478,N_39316);
nand U40260 (N_40260,N_39844,N_39059);
xor U40261 (N_40261,N_39685,N_39936);
or U40262 (N_40262,N_39452,N_39950);
nand U40263 (N_40263,N_39215,N_39777);
nor U40264 (N_40264,N_39029,N_39596);
or U40265 (N_40265,N_39595,N_39912);
nand U40266 (N_40266,N_39395,N_39948);
nor U40267 (N_40267,N_39263,N_39727);
xor U40268 (N_40268,N_39928,N_39607);
or U40269 (N_40269,N_39873,N_39603);
or U40270 (N_40270,N_39468,N_39218);
xnor U40271 (N_40271,N_39799,N_39684);
or U40272 (N_40272,N_39916,N_39100);
nand U40273 (N_40273,N_39055,N_39508);
or U40274 (N_40274,N_39368,N_39868);
or U40275 (N_40275,N_39467,N_39391);
nand U40276 (N_40276,N_39605,N_39574);
and U40277 (N_40277,N_39741,N_39747);
and U40278 (N_40278,N_39875,N_39008);
xor U40279 (N_40279,N_39236,N_39450);
nor U40280 (N_40280,N_39828,N_39570);
xor U40281 (N_40281,N_39733,N_39803);
or U40282 (N_40282,N_39116,N_39131);
or U40283 (N_40283,N_39323,N_39451);
xor U40284 (N_40284,N_39889,N_39558);
or U40285 (N_40285,N_39791,N_39473);
nor U40286 (N_40286,N_39964,N_39357);
nand U40287 (N_40287,N_39095,N_39363);
and U40288 (N_40288,N_39022,N_39463);
nand U40289 (N_40289,N_39899,N_39768);
and U40290 (N_40290,N_39223,N_39469);
or U40291 (N_40291,N_39830,N_39216);
nor U40292 (N_40292,N_39907,N_39012);
and U40293 (N_40293,N_39502,N_39620);
or U40294 (N_40294,N_39492,N_39906);
and U40295 (N_40295,N_39811,N_39195);
and U40296 (N_40296,N_39783,N_39940);
nor U40297 (N_40297,N_39141,N_39253);
and U40298 (N_40298,N_39855,N_39985);
xor U40299 (N_40299,N_39092,N_39805);
or U40300 (N_40300,N_39657,N_39539);
and U40301 (N_40301,N_39923,N_39336);
xnor U40302 (N_40302,N_39840,N_39745);
and U40303 (N_40303,N_39436,N_39020);
or U40304 (N_40304,N_39877,N_39279);
nor U40305 (N_40305,N_39031,N_39642);
or U40306 (N_40306,N_39061,N_39147);
xor U40307 (N_40307,N_39797,N_39388);
nand U40308 (N_40308,N_39211,N_39667);
or U40309 (N_40309,N_39608,N_39697);
and U40310 (N_40310,N_39789,N_39700);
and U40311 (N_40311,N_39901,N_39621);
or U40312 (N_40312,N_39277,N_39578);
and U40313 (N_40313,N_39041,N_39331);
or U40314 (N_40314,N_39048,N_39383);
xnor U40315 (N_40315,N_39366,N_39664);
or U40316 (N_40316,N_39145,N_39957);
nor U40317 (N_40317,N_39006,N_39949);
or U40318 (N_40318,N_39054,N_39622);
or U40319 (N_40319,N_39339,N_39566);
nor U40320 (N_40320,N_39659,N_39194);
nand U40321 (N_40321,N_39737,N_39405);
and U40322 (N_40322,N_39846,N_39927);
nand U40323 (N_40323,N_39999,N_39032);
and U40324 (N_40324,N_39648,N_39248);
xor U40325 (N_40325,N_39816,N_39538);
nand U40326 (N_40326,N_39564,N_39764);
xor U40327 (N_40327,N_39987,N_39636);
nand U40328 (N_40328,N_39692,N_39834);
xor U40329 (N_40329,N_39726,N_39746);
or U40330 (N_40330,N_39265,N_39285);
and U40331 (N_40331,N_39050,N_39015);
or U40332 (N_40332,N_39905,N_39256);
or U40333 (N_40333,N_39259,N_39386);
or U40334 (N_40334,N_39151,N_39853);
nand U40335 (N_40335,N_39552,N_39796);
and U40336 (N_40336,N_39058,N_39695);
or U40337 (N_40337,N_39245,N_39495);
nand U40338 (N_40338,N_39665,N_39503);
xor U40339 (N_40339,N_39989,N_39398);
or U40340 (N_40340,N_39753,N_39847);
xnor U40341 (N_40341,N_39560,N_39448);
nand U40342 (N_40342,N_39879,N_39749);
xnor U40343 (N_40343,N_39387,N_39954);
and U40344 (N_40344,N_39461,N_39046);
xnor U40345 (N_40345,N_39355,N_39496);
nand U40346 (N_40346,N_39705,N_39241);
nand U40347 (N_40347,N_39329,N_39841);
xor U40348 (N_40348,N_39402,N_39490);
nor U40349 (N_40349,N_39155,N_39047);
and U40350 (N_40350,N_39472,N_39372);
xnor U40351 (N_40351,N_39146,N_39212);
xor U40352 (N_40352,N_39420,N_39856);
nand U40353 (N_40353,N_39242,N_39666);
xnor U40354 (N_40354,N_39179,N_39350);
xor U40355 (N_40355,N_39098,N_39988);
and U40356 (N_40356,N_39033,N_39818);
xnor U40357 (N_40357,N_39635,N_39361);
nand U40358 (N_40358,N_39758,N_39848);
or U40359 (N_40359,N_39878,N_39258);
xnor U40360 (N_40360,N_39870,N_39214);
nand U40361 (N_40361,N_39456,N_39222);
or U40362 (N_40362,N_39143,N_39507);
xnor U40363 (N_40363,N_39865,N_39273);
and U40364 (N_40364,N_39592,N_39063);
xor U40365 (N_40365,N_39434,N_39996);
nand U40366 (N_40366,N_39970,N_39817);
and U40367 (N_40367,N_39663,N_39838);
nor U40368 (N_40368,N_39123,N_39009);
nand U40369 (N_40369,N_39569,N_39079);
and U40370 (N_40370,N_39699,N_39257);
and U40371 (N_40371,N_39991,N_39738);
and U40372 (N_40372,N_39475,N_39254);
nor U40373 (N_40373,N_39374,N_39986);
xnor U40374 (N_40374,N_39207,N_39182);
nor U40375 (N_40375,N_39960,N_39716);
nand U40376 (N_40376,N_39431,N_39351);
or U40377 (N_40377,N_39720,N_39064);
nor U40378 (N_40378,N_39024,N_39952);
and U40379 (N_40379,N_39278,N_39454);
and U40380 (N_40380,N_39364,N_39680);
nor U40381 (N_40381,N_39471,N_39833);
nand U40382 (N_40382,N_39272,N_39839);
or U40383 (N_40383,N_39172,N_39209);
xnor U40384 (N_40384,N_39837,N_39976);
and U40385 (N_40385,N_39005,N_39859);
xor U40386 (N_40386,N_39788,N_39537);
nand U40387 (N_40387,N_39327,N_39202);
nor U40388 (N_40388,N_39314,N_39610);
and U40389 (N_40389,N_39003,N_39618);
nor U40390 (N_40390,N_39217,N_39232);
and U40391 (N_40391,N_39150,N_39429);
and U40392 (N_40392,N_39910,N_39354);
nor U40393 (N_40393,N_39947,N_39251);
or U40394 (N_40394,N_39305,N_39342);
nor U40395 (N_40395,N_39085,N_39119);
or U40396 (N_40396,N_39433,N_39523);
nor U40397 (N_40397,N_39654,N_39640);
and U40398 (N_40398,N_39010,N_39290);
xnor U40399 (N_40399,N_39655,N_39708);
xor U40400 (N_40400,N_39038,N_39170);
nor U40401 (N_40401,N_39224,N_39766);
nand U40402 (N_40402,N_39832,N_39233);
or U40403 (N_40403,N_39632,N_39093);
or U40404 (N_40404,N_39220,N_39309);
nor U40405 (N_40405,N_39900,N_39971);
and U40406 (N_40406,N_39968,N_39944);
or U40407 (N_40407,N_39246,N_39400);
or U40408 (N_40408,N_39581,N_39362);
xor U40409 (N_40409,N_39288,N_39925);
xnor U40410 (N_40410,N_39152,N_39933);
nor U40411 (N_40411,N_39353,N_39338);
xnor U40412 (N_40412,N_39173,N_39577);
or U40413 (N_40413,N_39043,N_39174);
and U40414 (N_40414,N_39493,N_39360);
nor U40415 (N_40415,N_39575,N_39125);
xor U40416 (N_40416,N_39660,N_39590);
or U40417 (N_40417,N_39835,N_39073);
nand U40418 (N_40418,N_39286,N_39629);
xnor U40419 (N_40419,N_39623,N_39168);
nand U40420 (N_40420,N_39599,N_39546);
nor U40421 (N_40421,N_39083,N_39943);
or U40422 (N_40422,N_39862,N_39326);
nor U40423 (N_40423,N_39162,N_39972);
or U40424 (N_40424,N_39130,N_39647);
nand U40425 (N_40425,N_39324,N_39267);
xnor U40426 (N_40426,N_39294,N_39199);
nand U40427 (N_40427,N_39565,N_39090);
or U40428 (N_40428,N_39088,N_39641);
or U40429 (N_40429,N_39961,N_39915);
and U40430 (N_40430,N_39239,N_39381);
and U40431 (N_40431,N_39785,N_39544);
nor U40432 (N_40432,N_39103,N_39689);
xor U40433 (N_40433,N_39053,N_39255);
or U40434 (N_40434,N_39513,N_39937);
xnor U40435 (N_40435,N_39140,N_39525);
or U40436 (N_40436,N_39394,N_39633);
nor U40437 (N_40437,N_39237,N_39885);
nand U40438 (N_40438,N_39072,N_39963);
and U40439 (N_40439,N_39489,N_39343);
or U40440 (N_40440,N_39408,N_39627);
nand U40441 (N_40441,N_39295,N_39533);
or U40442 (N_40442,N_39106,N_39287);
xor U40443 (N_40443,N_39760,N_39426);
xnor U40444 (N_40444,N_39382,N_39365);
xnor U40445 (N_40445,N_39001,N_39035);
nand U40446 (N_40446,N_39932,N_39955);
nor U40447 (N_40447,N_39814,N_39269);
and U40448 (N_40448,N_39412,N_39160);
or U40449 (N_40449,N_39965,N_39557);
xor U40450 (N_40450,N_39481,N_39742);
or U40451 (N_40451,N_39052,N_39023);
or U40452 (N_40452,N_39686,N_39328);
nand U40453 (N_40453,N_39017,N_39349);
nand U40454 (N_40454,N_39669,N_39612);
nand U40455 (N_40455,N_39066,N_39225);
nand U40456 (N_40456,N_39071,N_39984);
nor U40457 (N_40457,N_39625,N_39260);
nand U40458 (N_40458,N_39638,N_39049);
or U40459 (N_40459,N_39981,N_39582);
or U40460 (N_40460,N_39866,N_39197);
nor U40461 (N_40461,N_39138,N_39696);
and U40462 (N_40462,N_39221,N_39384);
or U40463 (N_40463,N_39030,N_39226);
nor U40464 (N_40464,N_39951,N_39920);
xnor U40465 (N_40465,N_39773,N_39583);
xnor U40466 (N_40466,N_39154,N_39021);
and U40467 (N_40467,N_39466,N_39958);
or U40468 (N_40468,N_39594,N_39890);
xor U40469 (N_40469,N_39924,N_39186);
or U40470 (N_40470,N_39993,N_39084);
nand U40471 (N_40471,N_39406,N_39425);
and U40472 (N_40472,N_39974,N_39480);
or U40473 (N_40473,N_39767,N_39299);
nand U40474 (N_40474,N_39526,N_39732);
or U40475 (N_40475,N_39312,N_39515);
nor U40476 (N_40476,N_39086,N_39266);
xnor U40477 (N_40477,N_39897,N_39137);
and U40478 (N_40478,N_39113,N_39926);
xnor U40479 (N_40479,N_39166,N_39786);
or U40480 (N_40480,N_39938,N_39775);
nand U40481 (N_40481,N_39769,N_39604);
nand U40482 (N_40482,N_39554,N_39310);
nor U40483 (N_40483,N_39122,N_39815);
nor U40484 (N_40484,N_39823,N_39810);
nor U40485 (N_40485,N_39619,N_39087);
xor U40486 (N_40486,N_39344,N_39261);
nor U40487 (N_40487,N_39671,N_39274);
xnor U40488 (N_40488,N_39167,N_39756);
nand U40489 (N_40489,N_39798,N_39532);
or U40490 (N_40490,N_39458,N_39861);
nand U40491 (N_40491,N_39319,N_39498);
nor U40492 (N_40492,N_39709,N_39969);
nor U40493 (N_40493,N_39826,N_39842);
and U40494 (N_40494,N_39744,N_39177);
or U40495 (N_40495,N_39782,N_39694);
and U40496 (N_40496,N_39201,N_39643);
nand U40497 (N_40497,N_39112,N_39132);
and U40498 (N_40498,N_39036,N_39378);
nand U40499 (N_40499,N_39858,N_39499);
or U40500 (N_40500,N_39715,N_39430);
nand U40501 (N_40501,N_39743,N_39484);
and U40502 (N_40502,N_39028,N_39976);
xnor U40503 (N_40503,N_39667,N_39032);
xor U40504 (N_40504,N_39031,N_39247);
xor U40505 (N_40505,N_39731,N_39941);
xnor U40506 (N_40506,N_39242,N_39350);
and U40507 (N_40507,N_39604,N_39161);
nand U40508 (N_40508,N_39280,N_39424);
xor U40509 (N_40509,N_39717,N_39970);
xor U40510 (N_40510,N_39267,N_39901);
nor U40511 (N_40511,N_39957,N_39219);
xor U40512 (N_40512,N_39527,N_39642);
and U40513 (N_40513,N_39010,N_39805);
and U40514 (N_40514,N_39636,N_39302);
xnor U40515 (N_40515,N_39353,N_39797);
xor U40516 (N_40516,N_39082,N_39846);
and U40517 (N_40517,N_39972,N_39040);
and U40518 (N_40518,N_39271,N_39938);
xnor U40519 (N_40519,N_39604,N_39784);
xor U40520 (N_40520,N_39310,N_39968);
and U40521 (N_40521,N_39462,N_39132);
xor U40522 (N_40522,N_39969,N_39707);
xnor U40523 (N_40523,N_39390,N_39120);
xnor U40524 (N_40524,N_39254,N_39791);
nand U40525 (N_40525,N_39379,N_39654);
xnor U40526 (N_40526,N_39471,N_39951);
and U40527 (N_40527,N_39923,N_39458);
xnor U40528 (N_40528,N_39723,N_39918);
nand U40529 (N_40529,N_39876,N_39351);
or U40530 (N_40530,N_39569,N_39501);
nor U40531 (N_40531,N_39885,N_39830);
and U40532 (N_40532,N_39621,N_39408);
nor U40533 (N_40533,N_39487,N_39230);
or U40534 (N_40534,N_39948,N_39099);
xnor U40535 (N_40535,N_39519,N_39077);
and U40536 (N_40536,N_39782,N_39641);
and U40537 (N_40537,N_39595,N_39256);
and U40538 (N_40538,N_39412,N_39464);
or U40539 (N_40539,N_39047,N_39857);
nor U40540 (N_40540,N_39404,N_39890);
nand U40541 (N_40541,N_39288,N_39907);
nand U40542 (N_40542,N_39508,N_39775);
and U40543 (N_40543,N_39776,N_39100);
and U40544 (N_40544,N_39942,N_39796);
or U40545 (N_40545,N_39407,N_39591);
and U40546 (N_40546,N_39069,N_39727);
xor U40547 (N_40547,N_39376,N_39837);
nand U40548 (N_40548,N_39002,N_39732);
and U40549 (N_40549,N_39833,N_39446);
xnor U40550 (N_40550,N_39540,N_39646);
xor U40551 (N_40551,N_39690,N_39656);
and U40552 (N_40552,N_39226,N_39571);
and U40553 (N_40553,N_39287,N_39598);
xnor U40554 (N_40554,N_39971,N_39593);
nor U40555 (N_40555,N_39801,N_39437);
xor U40556 (N_40556,N_39094,N_39435);
or U40557 (N_40557,N_39890,N_39035);
nor U40558 (N_40558,N_39142,N_39451);
nand U40559 (N_40559,N_39918,N_39395);
xor U40560 (N_40560,N_39546,N_39623);
xnor U40561 (N_40561,N_39465,N_39486);
or U40562 (N_40562,N_39530,N_39807);
and U40563 (N_40563,N_39296,N_39050);
nor U40564 (N_40564,N_39019,N_39085);
or U40565 (N_40565,N_39463,N_39138);
nand U40566 (N_40566,N_39289,N_39022);
and U40567 (N_40567,N_39953,N_39821);
nor U40568 (N_40568,N_39651,N_39195);
and U40569 (N_40569,N_39396,N_39825);
or U40570 (N_40570,N_39543,N_39580);
nand U40571 (N_40571,N_39098,N_39542);
nor U40572 (N_40572,N_39990,N_39570);
xnor U40573 (N_40573,N_39919,N_39414);
nand U40574 (N_40574,N_39153,N_39372);
xnor U40575 (N_40575,N_39835,N_39772);
xor U40576 (N_40576,N_39488,N_39307);
nor U40577 (N_40577,N_39002,N_39261);
nor U40578 (N_40578,N_39884,N_39710);
xor U40579 (N_40579,N_39745,N_39592);
and U40580 (N_40580,N_39723,N_39777);
or U40581 (N_40581,N_39856,N_39998);
and U40582 (N_40582,N_39984,N_39104);
and U40583 (N_40583,N_39334,N_39161);
nor U40584 (N_40584,N_39272,N_39053);
nor U40585 (N_40585,N_39116,N_39743);
and U40586 (N_40586,N_39735,N_39738);
and U40587 (N_40587,N_39722,N_39298);
xor U40588 (N_40588,N_39640,N_39506);
nand U40589 (N_40589,N_39323,N_39512);
and U40590 (N_40590,N_39560,N_39951);
and U40591 (N_40591,N_39329,N_39973);
nand U40592 (N_40592,N_39617,N_39725);
and U40593 (N_40593,N_39948,N_39037);
nor U40594 (N_40594,N_39564,N_39237);
nand U40595 (N_40595,N_39644,N_39005);
xnor U40596 (N_40596,N_39378,N_39691);
or U40597 (N_40597,N_39045,N_39157);
nor U40598 (N_40598,N_39926,N_39477);
nand U40599 (N_40599,N_39029,N_39698);
nand U40600 (N_40600,N_39045,N_39412);
or U40601 (N_40601,N_39415,N_39707);
nand U40602 (N_40602,N_39648,N_39675);
or U40603 (N_40603,N_39078,N_39069);
or U40604 (N_40604,N_39207,N_39002);
or U40605 (N_40605,N_39169,N_39429);
and U40606 (N_40606,N_39856,N_39949);
and U40607 (N_40607,N_39888,N_39764);
and U40608 (N_40608,N_39090,N_39934);
and U40609 (N_40609,N_39985,N_39812);
nor U40610 (N_40610,N_39323,N_39290);
nand U40611 (N_40611,N_39015,N_39326);
or U40612 (N_40612,N_39479,N_39859);
xor U40613 (N_40613,N_39124,N_39081);
nor U40614 (N_40614,N_39679,N_39196);
or U40615 (N_40615,N_39728,N_39897);
or U40616 (N_40616,N_39937,N_39697);
and U40617 (N_40617,N_39972,N_39821);
nand U40618 (N_40618,N_39675,N_39383);
xnor U40619 (N_40619,N_39837,N_39285);
xnor U40620 (N_40620,N_39600,N_39576);
xor U40621 (N_40621,N_39061,N_39655);
nand U40622 (N_40622,N_39844,N_39656);
or U40623 (N_40623,N_39952,N_39709);
nand U40624 (N_40624,N_39672,N_39806);
xnor U40625 (N_40625,N_39826,N_39077);
and U40626 (N_40626,N_39418,N_39992);
nand U40627 (N_40627,N_39456,N_39744);
xnor U40628 (N_40628,N_39992,N_39657);
nand U40629 (N_40629,N_39590,N_39654);
and U40630 (N_40630,N_39315,N_39070);
xnor U40631 (N_40631,N_39994,N_39761);
xor U40632 (N_40632,N_39695,N_39239);
and U40633 (N_40633,N_39110,N_39768);
and U40634 (N_40634,N_39342,N_39285);
nand U40635 (N_40635,N_39216,N_39236);
nor U40636 (N_40636,N_39660,N_39200);
or U40637 (N_40637,N_39854,N_39512);
and U40638 (N_40638,N_39926,N_39980);
nor U40639 (N_40639,N_39746,N_39126);
nor U40640 (N_40640,N_39152,N_39707);
nand U40641 (N_40641,N_39712,N_39705);
xor U40642 (N_40642,N_39313,N_39433);
or U40643 (N_40643,N_39277,N_39718);
and U40644 (N_40644,N_39176,N_39861);
nor U40645 (N_40645,N_39156,N_39533);
nand U40646 (N_40646,N_39552,N_39761);
nor U40647 (N_40647,N_39914,N_39769);
or U40648 (N_40648,N_39098,N_39172);
xnor U40649 (N_40649,N_39851,N_39398);
xor U40650 (N_40650,N_39104,N_39876);
or U40651 (N_40651,N_39540,N_39205);
and U40652 (N_40652,N_39521,N_39803);
and U40653 (N_40653,N_39050,N_39212);
nand U40654 (N_40654,N_39498,N_39165);
nand U40655 (N_40655,N_39392,N_39109);
nand U40656 (N_40656,N_39623,N_39044);
and U40657 (N_40657,N_39725,N_39263);
xnor U40658 (N_40658,N_39642,N_39217);
nor U40659 (N_40659,N_39759,N_39040);
xnor U40660 (N_40660,N_39128,N_39866);
or U40661 (N_40661,N_39663,N_39384);
xor U40662 (N_40662,N_39238,N_39949);
xor U40663 (N_40663,N_39944,N_39877);
and U40664 (N_40664,N_39334,N_39018);
xnor U40665 (N_40665,N_39722,N_39994);
or U40666 (N_40666,N_39485,N_39012);
nand U40667 (N_40667,N_39820,N_39124);
and U40668 (N_40668,N_39283,N_39788);
nor U40669 (N_40669,N_39264,N_39527);
xnor U40670 (N_40670,N_39870,N_39560);
nor U40671 (N_40671,N_39879,N_39225);
or U40672 (N_40672,N_39912,N_39408);
nand U40673 (N_40673,N_39734,N_39069);
or U40674 (N_40674,N_39660,N_39340);
and U40675 (N_40675,N_39169,N_39800);
nand U40676 (N_40676,N_39614,N_39960);
and U40677 (N_40677,N_39916,N_39469);
and U40678 (N_40678,N_39190,N_39076);
or U40679 (N_40679,N_39341,N_39852);
nor U40680 (N_40680,N_39810,N_39513);
nand U40681 (N_40681,N_39677,N_39659);
xor U40682 (N_40682,N_39362,N_39645);
or U40683 (N_40683,N_39752,N_39222);
and U40684 (N_40684,N_39620,N_39295);
or U40685 (N_40685,N_39953,N_39395);
or U40686 (N_40686,N_39060,N_39273);
or U40687 (N_40687,N_39736,N_39012);
nor U40688 (N_40688,N_39900,N_39422);
xor U40689 (N_40689,N_39043,N_39904);
nand U40690 (N_40690,N_39841,N_39800);
nor U40691 (N_40691,N_39074,N_39710);
nor U40692 (N_40692,N_39414,N_39130);
xnor U40693 (N_40693,N_39131,N_39704);
and U40694 (N_40694,N_39398,N_39156);
and U40695 (N_40695,N_39145,N_39658);
or U40696 (N_40696,N_39065,N_39199);
or U40697 (N_40697,N_39907,N_39203);
nand U40698 (N_40698,N_39530,N_39919);
and U40699 (N_40699,N_39473,N_39483);
and U40700 (N_40700,N_39009,N_39998);
and U40701 (N_40701,N_39085,N_39598);
and U40702 (N_40702,N_39786,N_39848);
or U40703 (N_40703,N_39321,N_39505);
and U40704 (N_40704,N_39723,N_39640);
nor U40705 (N_40705,N_39114,N_39314);
xor U40706 (N_40706,N_39225,N_39119);
and U40707 (N_40707,N_39129,N_39435);
nand U40708 (N_40708,N_39140,N_39970);
or U40709 (N_40709,N_39788,N_39486);
and U40710 (N_40710,N_39815,N_39374);
and U40711 (N_40711,N_39775,N_39812);
nand U40712 (N_40712,N_39860,N_39444);
or U40713 (N_40713,N_39025,N_39075);
nor U40714 (N_40714,N_39580,N_39588);
xor U40715 (N_40715,N_39933,N_39223);
nor U40716 (N_40716,N_39142,N_39576);
and U40717 (N_40717,N_39063,N_39568);
or U40718 (N_40718,N_39735,N_39070);
nor U40719 (N_40719,N_39026,N_39191);
xor U40720 (N_40720,N_39178,N_39225);
xnor U40721 (N_40721,N_39835,N_39325);
or U40722 (N_40722,N_39770,N_39473);
or U40723 (N_40723,N_39167,N_39220);
xor U40724 (N_40724,N_39116,N_39988);
or U40725 (N_40725,N_39112,N_39499);
and U40726 (N_40726,N_39015,N_39963);
and U40727 (N_40727,N_39219,N_39023);
nor U40728 (N_40728,N_39435,N_39681);
nand U40729 (N_40729,N_39542,N_39697);
or U40730 (N_40730,N_39655,N_39358);
nor U40731 (N_40731,N_39570,N_39262);
xor U40732 (N_40732,N_39699,N_39851);
nor U40733 (N_40733,N_39414,N_39649);
xnor U40734 (N_40734,N_39236,N_39825);
or U40735 (N_40735,N_39673,N_39215);
nand U40736 (N_40736,N_39354,N_39741);
and U40737 (N_40737,N_39209,N_39796);
nor U40738 (N_40738,N_39956,N_39334);
and U40739 (N_40739,N_39126,N_39117);
or U40740 (N_40740,N_39249,N_39801);
or U40741 (N_40741,N_39875,N_39805);
or U40742 (N_40742,N_39856,N_39033);
or U40743 (N_40743,N_39525,N_39960);
nand U40744 (N_40744,N_39579,N_39553);
xor U40745 (N_40745,N_39179,N_39815);
or U40746 (N_40746,N_39793,N_39977);
or U40747 (N_40747,N_39643,N_39702);
nand U40748 (N_40748,N_39496,N_39015);
xor U40749 (N_40749,N_39764,N_39939);
nor U40750 (N_40750,N_39461,N_39118);
xor U40751 (N_40751,N_39749,N_39251);
or U40752 (N_40752,N_39641,N_39729);
or U40753 (N_40753,N_39453,N_39117);
nand U40754 (N_40754,N_39051,N_39721);
xor U40755 (N_40755,N_39742,N_39950);
nand U40756 (N_40756,N_39636,N_39404);
or U40757 (N_40757,N_39198,N_39085);
nand U40758 (N_40758,N_39157,N_39371);
xor U40759 (N_40759,N_39006,N_39550);
nand U40760 (N_40760,N_39060,N_39724);
xor U40761 (N_40761,N_39335,N_39137);
nand U40762 (N_40762,N_39919,N_39052);
nand U40763 (N_40763,N_39556,N_39878);
nand U40764 (N_40764,N_39042,N_39573);
nor U40765 (N_40765,N_39890,N_39532);
nor U40766 (N_40766,N_39046,N_39162);
nand U40767 (N_40767,N_39595,N_39609);
and U40768 (N_40768,N_39001,N_39996);
xor U40769 (N_40769,N_39078,N_39812);
xnor U40770 (N_40770,N_39632,N_39999);
xnor U40771 (N_40771,N_39882,N_39774);
or U40772 (N_40772,N_39475,N_39224);
and U40773 (N_40773,N_39051,N_39585);
nor U40774 (N_40774,N_39992,N_39919);
nor U40775 (N_40775,N_39227,N_39438);
nand U40776 (N_40776,N_39372,N_39897);
and U40777 (N_40777,N_39051,N_39495);
xnor U40778 (N_40778,N_39064,N_39370);
or U40779 (N_40779,N_39738,N_39240);
nor U40780 (N_40780,N_39342,N_39054);
or U40781 (N_40781,N_39180,N_39718);
nand U40782 (N_40782,N_39457,N_39342);
or U40783 (N_40783,N_39508,N_39118);
xor U40784 (N_40784,N_39476,N_39220);
or U40785 (N_40785,N_39395,N_39519);
xnor U40786 (N_40786,N_39014,N_39050);
nor U40787 (N_40787,N_39300,N_39635);
nor U40788 (N_40788,N_39821,N_39994);
or U40789 (N_40789,N_39581,N_39770);
or U40790 (N_40790,N_39824,N_39346);
or U40791 (N_40791,N_39955,N_39411);
nor U40792 (N_40792,N_39672,N_39693);
and U40793 (N_40793,N_39071,N_39405);
xor U40794 (N_40794,N_39237,N_39259);
xor U40795 (N_40795,N_39875,N_39571);
and U40796 (N_40796,N_39077,N_39290);
nor U40797 (N_40797,N_39366,N_39774);
xor U40798 (N_40798,N_39358,N_39918);
xnor U40799 (N_40799,N_39344,N_39479);
xnor U40800 (N_40800,N_39854,N_39965);
or U40801 (N_40801,N_39164,N_39305);
nor U40802 (N_40802,N_39205,N_39926);
nor U40803 (N_40803,N_39760,N_39396);
and U40804 (N_40804,N_39494,N_39020);
xnor U40805 (N_40805,N_39823,N_39101);
nor U40806 (N_40806,N_39048,N_39683);
xor U40807 (N_40807,N_39173,N_39285);
nand U40808 (N_40808,N_39042,N_39397);
xor U40809 (N_40809,N_39122,N_39331);
xor U40810 (N_40810,N_39456,N_39408);
nand U40811 (N_40811,N_39425,N_39285);
xnor U40812 (N_40812,N_39957,N_39479);
and U40813 (N_40813,N_39496,N_39133);
and U40814 (N_40814,N_39511,N_39488);
nand U40815 (N_40815,N_39496,N_39643);
and U40816 (N_40816,N_39312,N_39104);
or U40817 (N_40817,N_39172,N_39830);
xor U40818 (N_40818,N_39819,N_39020);
nand U40819 (N_40819,N_39437,N_39194);
nor U40820 (N_40820,N_39601,N_39639);
nor U40821 (N_40821,N_39483,N_39055);
nor U40822 (N_40822,N_39440,N_39653);
or U40823 (N_40823,N_39973,N_39365);
and U40824 (N_40824,N_39955,N_39901);
and U40825 (N_40825,N_39163,N_39140);
and U40826 (N_40826,N_39928,N_39315);
xnor U40827 (N_40827,N_39700,N_39425);
or U40828 (N_40828,N_39208,N_39384);
nor U40829 (N_40829,N_39269,N_39242);
xnor U40830 (N_40830,N_39165,N_39056);
or U40831 (N_40831,N_39263,N_39631);
xnor U40832 (N_40832,N_39802,N_39204);
nand U40833 (N_40833,N_39647,N_39155);
xor U40834 (N_40834,N_39477,N_39845);
nor U40835 (N_40835,N_39062,N_39029);
and U40836 (N_40836,N_39569,N_39944);
and U40837 (N_40837,N_39649,N_39322);
nor U40838 (N_40838,N_39830,N_39698);
or U40839 (N_40839,N_39241,N_39540);
nor U40840 (N_40840,N_39471,N_39010);
nand U40841 (N_40841,N_39991,N_39690);
nor U40842 (N_40842,N_39085,N_39915);
and U40843 (N_40843,N_39366,N_39981);
or U40844 (N_40844,N_39291,N_39536);
xor U40845 (N_40845,N_39792,N_39067);
and U40846 (N_40846,N_39308,N_39848);
nor U40847 (N_40847,N_39028,N_39667);
nor U40848 (N_40848,N_39754,N_39874);
and U40849 (N_40849,N_39279,N_39366);
or U40850 (N_40850,N_39582,N_39356);
nand U40851 (N_40851,N_39151,N_39765);
nand U40852 (N_40852,N_39148,N_39686);
xor U40853 (N_40853,N_39592,N_39515);
nor U40854 (N_40854,N_39459,N_39977);
nor U40855 (N_40855,N_39709,N_39643);
nor U40856 (N_40856,N_39482,N_39432);
or U40857 (N_40857,N_39985,N_39695);
xor U40858 (N_40858,N_39747,N_39225);
xor U40859 (N_40859,N_39271,N_39954);
nor U40860 (N_40860,N_39120,N_39221);
nand U40861 (N_40861,N_39487,N_39130);
xor U40862 (N_40862,N_39332,N_39277);
xor U40863 (N_40863,N_39839,N_39284);
nand U40864 (N_40864,N_39427,N_39024);
nor U40865 (N_40865,N_39165,N_39905);
and U40866 (N_40866,N_39100,N_39903);
or U40867 (N_40867,N_39586,N_39364);
nand U40868 (N_40868,N_39930,N_39041);
nand U40869 (N_40869,N_39738,N_39655);
xnor U40870 (N_40870,N_39307,N_39760);
xnor U40871 (N_40871,N_39548,N_39202);
or U40872 (N_40872,N_39489,N_39719);
xor U40873 (N_40873,N_39463,N_39438);
or U40874 (N_40874,N_39493,N_39414);
or U40875 (N_40875,N_39620,N_39031);
and U40876 (N_40876,N_39630,N_39918);
or U40877 (N_40877,N_39212,N_39578);
xor U40878 (N_40878,N_39964,N_39384);
nand U40879 (N_40879,N_39064,N_39185);
or U40880 (N_40880,N_39670,N_39440);
xnor U40881 (N_40881,N_39647,N_39306);
nor U40882 (N_40882,N_39291,N_39849);
xor U40883 (N_40883,N_39401,N_39039);
nor U40884 (N_40884,N_39501,N_39458);
xor U40885 (N_40885,N_39206,N_39334);
nand U40886 (N_40886,N_39952,N_39312);
nor U40887 (N_40887,N_39348,N_39938);
nor U40888 (N_40888,N_39735,N_39792);
nand U40889 (N_40889,N_39463,N_39120);
or U40890 (N_40890,N_39078,N_39077);
or U40891 (N_40891,N_39376,N_39583);
nor U40892 (N_40892,N_39873,N_39127);
nand U40893 (N_40893,N_39486,N_39773);
and U40894 (N_40894,N_39653,N_39514);
nor U40895 (N_40895,N_39187,N_39674);
and U40896 (N_40896,N_39287,N_39525);
nand U40897 (N_40897,N_39553,N_39188);
nand U40898 (N_40898,N_39444,N_39736);
or U40899 (N_40899,N_39613,N_39523);
xor U40900 (N_40900,N_39626,N_39417);
or U40901 (N_40901,N_39383,N_39545);
nor U40902 (N_40902,N_39658,N_39173);
or U40903 (N_40903,N_39235,N_39352);
nor U40904 (N_40904,N_39955,N_39607);
nor U40905 (N_40905,N_39207,N_39714);
nand U40906 (N_40906,N_39109,N_39288);
or U40907 (N_40907,N_39609,N_39418);
or U40908 (N_40908,N_39894,N_39029);
and U40909 (N_40909,N_39772,N_39905);
xor U40910 (N_40910,N_39742,N_39735);
and U40911 (N_40911,N_39631,N_39605);
and U40912 (N_40912,N_39630,N_39292);
nand U40913 (N_40913,N_39937,N_39289);
xor U40914 (N_40914,N_39796,N_39765);
or U40915 (N_40915,N_39471,N_39805);
xor U40916 (N_40916,N_39765,N_39605);
or U40917 (N_40917,N_39717,N_39146);
xnor U40918 (N_40918,N_39411,N_39275);
and U40919 (N_40919,N_39520,N_39886);
nor U40920 (N_40920,N_39850,N_39590);
nand U40921 (N_40921,N_39710,N_39066);
and U40922 (N_40922,N_39928,N_39587);
nand U40923 (N_40923,N_39005,N_39492);
and U40924 (N_40924,N_39516,N_39278);
and U40925 (N_40925,N_39291,N_39198);
xor U40926 (N_40926,N_39105,N_39727);
nand U40927 (N_40927,N_39986,N_39336);
xor U40928 (N_40928,N_39591,N_39966);
xor U40929 (N_40929,N_39033,N_39335);
nand U40930 (N_40930,N_39786,N_39047);
and U40931 (N_40931,N_39351,N_39451);
xnor U40932 (N_40932,N_39545,N_39857);
nand U40933 (N_40933,N_39734,N_39273);
nand U40934 (N_40934,N_39682,N_39073);
and U40935 (N_40935,N_39078,N_39217);
nand U40936 (N_40936,N_39883,N_39865);
and U40937 (N_40937,N_39102,N_39800);
xnor U40938 (N_40938,N_39877,N_39517);
xor U40939 (N_40939,N_39460,N_39067);
and U40940 (N_40940,N_39388,N_39582);
xor U40941 (N_40941,N_39765,N_39807);
xor U40942 (N_40942,N_39825,N_39120);
nand U40943 (N_40943,N_39763,N_39682);
xor U40944 (N_40944,N_39202,N_39352);
xor U40945 (N_40945,N_39344,N_39621);
nor U40946 (N_40946,N_39400,N_39856);
or U40947 (N_40947,N_39714,N_39505);
nor U40948 (N_40948,N_39904,N_39577);
or U40949 (N_40949,N_39513,N_39796);
nor U40950 (N_40950,N_39128,N_39786);
nor U40951 (N_40951,N_39115,N_39459);
and U40952 (N_40952,N_39211,N_39696);
xor U40953 (N_40953,N_39849,N_39336);
nand U40954 (N_40954,N_39665,N_39272);
nor U40955 (N_40955,N_39375,N_39975);
nor U40956 (N_40956,N_39752,N_39702);
or U40957 (N_40957,N_39416,N_39064);
nand U40958 (N_40958,N_39873,N_39235);
nand U40959 (N_40959,N_39964,N_39922);
or U40960 (N_40960,N_39750,N_39576);
or U40961 (N_40961,N_39937,N_39921);
nand U40962 (N_40962,N_39749,N_39121);
and U40963 (N_40963,N_39078,N_39459);
and U40964 (N_40964,N_39159,N_39229);
nand U40965 (N_40965,N_39270,N_39288);
and U40966 (N_40966,N_39064,N_39763);
nor U40967 (N_40967,N_39046,N_39856);
or U40968 (N_40968,N_39045,N_39383);
and U40969 (N_40969,N_39357,N_39329);
and U40970 (N_40970,N_39013,N_39620);
or U40971 (N_40971,N_39595,N_39186);
nand U40972 (N_40972,N_39120,N_39490);
nand U40973 (N_40973,N_39025,N_39382);
or U40974 (N_40974,N_39158,N_39087);
nor U40975 (N_40975,N_39054,N_39041);
nand U40976 (N_40976,N_39134,N_39572);
nor U40977 (N_40977,N_39507,N_39987);
xor U40978 (N_40978,N_39337,N_39718);
nand U40979 (N_40979,N_39115,N_39581);
xor U40980 (N_40980,N_39141,N_39953);
nor U40981 (N_40981,N_39804,N_39575);
and U40982 (N_40982,N_39266,N_39803);
and U40983 (N_40983,N_39551,N_39467);
nor U40984 (N_40984,N_39974,N_39302);
nor U40985 (N_40985,N_39592,N_39539);
or U40986 (N_40986,N_39730,N_39336);
nand U40987 (N_40987,N_39509,N_39726);
xor U40988 (N_40988,N_39807,N_39440);
and U40989 (N_40989,N_39423,N_39161);
nor U40990 (N_40990,N_39913,N_39157);
nor U40991 (N_40991,N_39849,N_39204);
nand U40992 (N_40992,N_39466,N_39506);
xnor U40993 (N_40993,N_39740,N_39085);
or U40994 (N_40994,N_39002,N_39597);
xor U40995 (N_40995,N_39022,N_39308);
xnor U40996 (N_40996,N_39496,N_39822);
xnor U40997 (N_40997,N_39572,N_39324);
or U40998 (N_40998,N_39841,N_39084);
and U40999 (N_40999,N_39775,N_39255);
and U41000 (N_41000,N_40497,N_40707);
xor U41001 (N_41001,N_40347,N_40157);
xor U41002 (N_41002,N_40668,N_40736);
and U41003 (N_41003,N_40795,N_40147);
nor U41004 (N_41004,N_40863,N_40273);
and U41005 (N_41005,N_40509,N_40426);
or U41006 (N_41006,N_40896,N_40304);
nand U41007 (N_41007,N_40044,N_40349);
xor U41008 (N_41008,N_40786,N_40012);
xor U41009 (N_41009,N_40139,N_40960);
or U41010 (N_41010,N_40965,N_40600);
or U41011 (N_41011,N_40845,N_40501);
or U41012 (N_41012,N_40335,N_40620);
nor U41013 (N_41013,N_40361,N_40872);
nand U41014 (N_41014,N_40033,N_40318);
or U41015 (N_41015,N_40913,N_40558);
or U41016 (N_41016,N_40907,N_40553);
or U41017 (N_41017,N_40594,N_40631);
nor U41018 (N_41018,N_40693,N_40161);
or U41019 (N_41019,N_40194,N_40251);
and U41020 (N_41020,N_40270,N_40485);
or U41021 (N_41021,N_40371,N_40592);
or U41022 (N_41022,N_40298,N_40534);
nand U41023 (N_41023,N_40019,N_40531);
xor U41024 (N_41024,N_40705,N_40290);
nor U41025 (N_41025,N_40819,N_40406);
or U41026 (N_41026,N_40908,N_40151);
xnor U41027 (N_41027,N_40843,N_40254);
and U41028 (N_41028,N_40543,N_40102);
xnor U41029 (N_41029,N_40510,N_40310);
xor U41030 (N_41030,N_40116,N_40419);
nor U41031 (N_41031,N_40765,N_40953);
nor U41032 (N_41032,N_40637,N_40894);
nand U41033 (N_41033,N_40153,N_40138);
nand U41034 (N_41034,N_40905,N_40587);
nand U41035 (N_41035,N_40833,N_40479);
and U41036 (N_41036,N_40740,N_40917);
and U41037 (N_41037,N_40458,N_40236);
xor U41038 (N_41038,N_40486,N_40517);
nand U41039 (N_41039,N_40932,N_40986);
xor U41040 (N_41040,N_40367,N_40372);
or U41041 (N_41041,N_40253,N_40459);
or U41042 (N_41042,N_40927,N_40959);
nand U41043 (N_41043,N_40149,N_40720);
or U41044 (N_41044,N_40520,N_40866);
nor U41045 (N_41045,N_40283,N_40137);
or U41046 (N_41046,N_40799,N_40989);
or U41047 (N_41047,N_40282,N_40280);
xor U41048 (N_41048,N_40985,N_40064);
nand U41049 (N_41049,N_40615,N_40067);
xnor U41050 (N_41050,N_40783,N_40537);
nand U41051 (N_41051,N_40784,N_40643);
nor U41052 (N_41052,N_40000,N_40040);
xor U41053 (N_41053,N_40011,N_40577);
nand U41054 (N_41054,N_40877,N_40548);
nor U41055 (N_41055,N_40164,N_40131);
nor U41056 (N_41056,N_40513,N_40195);
nand U41057 (N_41057,N_40460,N_40384);
xnor U41058 (N_41058,N_40902,N_40188);
nor U41059 (N_41059,N_40056,N_40591);
nand U41060 (N_41060,N_40689,N_40549);
or U41061 (N_41061,N_40821,N_40313);
nand U41062 (N_41062,N_40365,N_40136);
nand U41063 (N_41063,N_40632,N_40100);
and U41064 (N_41064,N_40084,N_40410);
xor U41065 (N_41065,N_40292,N_40690);
nand U41066 (N_41066,N_40070,N_40617);
nor U41067 (N_41067,N_40804,N_40774);
xnor U41068 (N_41068,N_40155,N_40465);
nand U41069 (N_41069,N_40876,N_40704);
nor U41070 (N_41070,N_40134,N_40619);
or U41071 (N_41071,N_40910,N_40996);
nand U41072 (N_41072,N_40726,N_40664);
nand U41073 (N_41073,N_40092,N_40235);
or U41074 (N_41074,N_40484,N_40069);
xnor U41075 (N_41075,N_40141,N_40453);
xnor U41076 (N_41076,N_40441,N_40108);
nor U41077 (N_41077,N_40246,N_40550);
and U41078 (N_41078,N_40432,N_40374);
and U41079 (N_41079,N_40091,N_40628);
and U41080 (N_41080,N_40807,N_40162);
nand U41081 (N_41081,N_40079,N_40608);
and U41082 (N_41082,N_40450,N_40709);
and U41083 (N_41083,N_40421,N_40754);
nor U41084 (N_41084,N_40182,N_40605);
and U41085 (N_41085,N_40115,N_40272);
xor U41086 (N_41086,N_40868,N_40013);
nor U41087 (N_41087,N_40507,N_40198);
nor U41088 (N_41088,N_40657,N_40424);
or U41089 (N_41089,N_40729,N_40023);
nor U41090 (N_41090,N_40455,N_40576);
nand U41091 (N_41091,N_40764,N_40593);
and U41092 (N_41092,N_40427,N_40468);
nor U41093 (N_41093,N_40284,N_40376);
or U41094 (N_41094,N_40275,N_40093);
xor U41095 (N_41095,N_40710,N_40206);
or U41096 (N_41096,N_40110,N_40768);
or U41097 (N_41097,N_40263,N_40487);
or U41098 (N_41098,N_40028,N_40844);
nand U41099 (N_41099,N_40052,N_40359);
and U41100 (N_41100,N_40285,N_40735);
nor U41101 (N_41101,N_40606,N_40538);
nor U41102 (N_41102,N_40966,N_40658);
xnor U41103 (N_41103,N_40350,N_40278);
or U41104 (N_41104,N_40626,N_40733);
and U41105 (N_41105,N_40076,N_40170);
and U41106 (N_41106,N_40224,N_40977);
nand U41107 (N_41107,N_40639,N_40914);
nand U41108 (N_41108,N_40680,N_40247);
nor U41109 (N_41109,N_40767,N_40055);
nand U41110 (N_41110,N_40345,N_40408);
nor U41111 (N_41111,N_40496,N_40926);
or U41112 (N_41112,N_40219,N_40482);
and U41113 (N_41113,N_40281,N_40015);
nand U41114 (N_41114,N_40744,N_40382);
or U41115 (N_41115,N_40622,N_40492);
nand U41116 (N_41116,N_40393,N_40677);
nor U41117 (N_41117,N_40941,N_40976);
and U41118 (N_41118,N_40422,N_40958);
nand U41119 (N_41119,N_40239,N_40429);
xor U41120 (N_41120,N_40603,N_40597);
nand U41121 (N_41121,N_40685,N_40679);
xor U41122 (N_41122,N_40732,N_40791);
xnor U41123 (N_41123,N_40536,N_40377);
and U41124 (N_41124,N_40113,N_40250);
or U41125 (N_41125,N_40823,N_40464);
or U41126 (N_41126,N_40030,N_40998);
xnor U41127 (N_41127,N_40261,N_40041);
and U41128 (N_41128,N_40363,N_40245);
nand U41129 (N_41129,N_40630,N_40865);
nand U41130 (N_41130,N_40255,N_40542);
nor U41131 (N_41131,N_40884,N_40666);
or U41132 (N_41132,N_40524,N_40994);
and U41133 (N_41133,N_40648,N_40301);
nand U41134 (N_41134,N_40293,N_40992);
xnor U41135 (N_41135,N_40925,N_40703);
or U41136 (N_41136,N_40739,N_40073);
and U41137 (N_41137,N_40330,N_40444);
and U41138 (N_41138,N_40808,N_40633);
or U41139 (N_41139,N_40718,N_40388);
nor U41140 (N_41140,N_40647,N_40706);
or U41141 (N_41141,N_40260,N_40470);
or U41142 (N_41142,N_40126,N_40233);
nor U41143 (N_41143,N_40081,N_40473);
and U41144 (N_41144,N_40665,N_40885);
nor U41145 (N_41145,N_40816,N_40319);
nand U41146 (N_41146,N_40955,N_40920);
nor U41147 (N_41147,N_40890,N_40584);
and U41148 (N_41148,N_40747,N_40200);
nand U41149 (N_41149,N_40752,N_40934);
and U41150 (N_41150,N_40915,N_40337);
nand U41151 (N_41151,N_40058,N_40922);
or U41152 (N_41152,N_40567,N_40080);
nor U41153 (N_41153,N_40849,N_40196);
nand U41154 (N_41154,N_40037,N_40189);
and U41155 (N_41155,N_40095,N_40174);
or U41156 (N_41156,N_40456,N_40984);
nand U41157 (N_41157,N_40667,N_40477);
or U41158 (N_41158,N_40684,N_40981);
xnor U41159 (N_41159,N_40858,N_40602);
nand U41160 (N_41160,N_40644,N_40949);
or U41161 (N_41161,N_40532,N_40651);
xnor U41162 (N_41162,N_40903,N_40105);
and U41163 (N_41163,N_40656,N_40692);
xnor U41164 (N_41164,N_40936,N_40771);
or U41165 (N_41165,N_40918,N_40888);
xor U41166 (N_41166,N_40880,N_40302);
and U41167 (N_41167,N_40225,N_40853);
nand U41168 (N_41168,N_40017,N_40323);
and U41169 (N_41169,N_40051,N_40488);
or U41170 (N_41170,N_40423,N_40066);
and U41171 (N_41171,N_40314,N_40268);
xnor U41172 (N_41172,N_40226,N_40154);
or U41173 (N_41173,N_40940,N_40860);
xor U41174 (N_41174,N_40653,N_40944);
nor U41175 (N_41175,N_40546,N_40118);
or U41176 (N_41176,N_40824,N_40589);
xor U41177 (N_41177,N_40386,N_40217);
and U41178 (N_41178,N_40851,N_40185);
nor U41179 (N_41179,N_40207,N_40036);
xnor U41180 (N_41180,N_40414,N_40878);
nor U41181 (N_41181,N_40463,N_40090);
or U41182 (N_41182,N_40541,N_40489);
nand U41183 (N_41183,N_40405,N_40794);
or U41184 (N_41184,N_40742,N_40063);
or U41185 (N_41185,N_40289,N_40930);
nand U41186 (N_41186,N_40906,N_40390);
or U41187 (N_41187,N_40010,N_40939);
or U41188 (N_41188,N_40336,N_40948);
and U41189 (N_41189,N_40223,N_40106);
and U41190 (N_41190,N_40760,N_40560);
and U41191 (N_41191,N_40448,N_40950);
nand U41192 (N_41192,N_40904,N_40383);
nand U41193 (N_41193,N_40249,N_40428);
xnor U41194 (N_41194,N_40723,N_40675);
or U41195 (N_41195,N_40053,N_40616);
nand U41196 (N_41196,N_40971,N_40176);
nand U41197 (N_41197,N_40837,N_40190);
nor U41198 (N_41198,N_40355,N_40697);
nand U41199 (N_41199,N_40215,N_40552);
and U41200 (N_41200,N_40535,N_40873);
nor U41201 (N_41201,N_40050,N_40924);
nor U41202 (N_41202,N_40623,N_40700);
nand U41203 (N_41203,N_40875,N_40121);
nor U41204 (N_41204,N_40687,N_40320);
xor U41205 (N_41205,N_40963,N_40334);
nand U41206 (N_41206,N_40835,N_40262);
and U41207 (N_41207,N_40610,N_40530);
nor U41208 (N_41208,N_40898,N_40775);
nor U41209 (N_41209,N_40714,N_40027);
xor U41210 (N_41210,N_40083,N_40803);
nor U41211 (N_41211,N_40437,N_40129);
nand U41212 (N_41212,N_40266,N_40022);
or U41213 (N_41213,N_40491,N_40598);
nor U41214 (N_41214,N_40395,N_40476);
nor U41215 (N_41215,N_40294,N_40269);
or U41216 (N_41216,N_40387,N_40018);
or U41217 (N_41217,N_40745,N_40978);
or U41218 (N_41218,N_40232,N_40451);
nor U41219 (N_41219,N_40974,N_40566);
and U41220 (N_41220,N_40523,N_40502);
and U41221 (N_41221,N_40208,N_40467);
nor U41222 (N_41222,N_40544,N_40681);
or U41223 (N_41223,N_40086,N_40369);
xor U41224 (N_41224,N_40825,N_40267);
or U41225 (N_41225,N_40344,N_40075);
xnor U41226 (N_41226,N_40452,N_40793);
nor U41227 (N_41227,N_40887,N_40564);
nand U41228 (N_41228,N_40306,N_40032);
and U41229 (N_41229,N_40391,N_40074);
nand U41230 (N_41230,N_40937,N_40466);
nor U41231 (N_41231,N_40234,N_40169);
nor U41232 (N_41232,N_40125,N_40662);
or U41233 (N_41233,N_40404,N_40059);
and U41234 (N_41234,N_40046,N_40265);
nor U41235 (N_41235,N_40181,N_40874);
nand U41236 (N_41236,N_40357,N_40407);
and U41237 (N_41237,N_40300,N_40440);
or U41238 (N_41238,N_40676,N_40750);
or U41239 (N_41239,N_40942,N_40144);
or U41240 (N_41240,N_40400,N_40039);
xor U41241 (N_41241,N_40859,N_40527);
xor U41242 (N_41242,N_40128,N_40228);
or U41243 (N_41243,N_40338,N_40385);
nand U41244 (N_41244,N_40691,N_40609);
nand U41245 (N_41245,N_40088,N_40834);
and U41246 (N_41246,N_40204,N_40167);
nor U41247 (N_41247,N_40140,N_40991);
xor U41248 (N_41248,N_40048,N_40831);
nand U41249 (N_41249,N_40921,N_40607);
nor U41250 (N_41250,N_40756,N_40431);
nand U41251 (N_41251,N_40462,N_40299);
and U41252 (N_41252,N_40127,N_40857);
nor U41253 (N_41253,N_40802,N_40743);
and U41254 (N_41254,N_40848,N_40413);
and U41255 (N_41255,N_40652,N_40326);
nand U41256 (N_41256,N_40499,N_40135);
or U41257 (N_41257,N_40746,N_40870);
and U41258 (N_41258,N_40686,N_40983);
or U41259 (N_41259,N_40852,N_40199);
and U41260 (N_41260,N_40782,N_40142);
and U41261 (N_41261,N_40979,N_40434);
and U41262 (N_41262,N_40370,N_40480);
nand U41263 (N_41263,N_40867,N_40026);
or U41264 (N_41264,N_40892,N_40505);
and U41265 (N_41265,N_40003,N_40340);
or U41266 (N_41266,N_40187,N_40449);
nand U41267 (N_41267,N_40655,N_40640);
nor U41268 (N_41268,N_40883,N_40230);
xor U41269 (N_41269,N_40715,N_40737);
xor U41270 (N_41270,N_40773,N_40798);
xor U41271 (N_41271,N_40586,N_40191);
and U41272 (N_41272,N_40415,N_40493);
or U41273 (N_41273,N_40165,N_40311);
nor U41274 (N_41274,N_40351,N_40087);
nor U41275 (N_41275,N_40258,N_40506);
xor U41276 (N_41276,N_40946,N_40826);
nor U41277 (N_41277,N_40214,N_40420);
xnor U41278 (N_41278,N_40529,N_40588);
xnor U41279 (N_41279,N_40178,N_40399);
nor U41280 (N_41280,N_40016,N_40346);
nor U41281 (N_41281,N_40721,N_40561);
or U41282 (N_41282,N_40177,N_40569);
or U41283 (N_41283,N_40820,N_40964);
nand U41284 (N_41284,N_40288,N_40730);
nor U41285 (N_41285,N_40297,N_40525);
nor U41286 (N_41286,N_40916,N_40518);
nor U41287 (N_41287,N_40770,N_40425);
xnor U41288 (N_41288,N_40559,N_40439);
or U41289 (N_41289,N_40728,N_40698);
nor U41290 (N_41290,N_40882,N_40057);
xor U41291 (N_41291,N_40585,N_40124);
or U41292 (N_41292,N_40815,N_40956);
nor U41293 (N_41293,N_40122,N_40741);
nand U41294 (N_41294,N_40114,N_40999);
or U41295 (N_41295,N_40007,N_40305);
and U41296 (N_41296,N_40160,N_40443);
and U41297 (N_41297,N_40861,N_40216);
xor U41298 (N_41298,N_40222,N_40919);
xor U41299 (N_41299,N_40243,N_40259);
or U41300 (N_41300,N_40333,N_40975);
nand U41301 (N_41301,N_40575,N_40389);
xnor U41302 (N_41302,N_40104,N_40909);
and U41303 (N_41303,N_40646,N_40929);
or U41304 (N_41304,N_40098,N_40009);
nor U41305 (N_41305,N_40143,N_40035);
and U41306 (N_41306,N_40001,N_40923);
xnor U41307 (N_41307,N_40341,N_40358);
and U41308 (N_41308,N_40495,N_40901);
xor U41309 (N_41309,N_40522,N_40082);
or U41310 (N_41310,N_40526,N_40547);
or U41311 (N_41311,N_40579,N_40990);
xnor U41312 (N_41312,N_40881,N_40213);
and U41313 (N_41313,N_40099,N_40928);
nor U41314 (N_41314,N_40781,N_40572);
nand U41315 (N_41315,N_40711,N_40797);
nand U41316 (N_41316,N_40461,N_40481);
nand U41317 (N_41317,N_40396,N_40331);
xor U41318 (N_41318,N_40109,N_40071);
or U41319 (N_41319,N_40248,N_40891);
nor U41320 (N_41320,N_40494,N_40378);
or U41321 (N_41321,N_40995,N_40308);
nand U41322 (N_41322,N_40047,N_40511);
xor U41323 (N_41323,N_40945,N_40734);
and U41324 (N_41324,N_40702,N_40997);
and U41325 (N_41325,N_40045,N_40533);
xor U41326 (N_41326,N_40869,N_40871);
nand U41327 (N_41327,N_40411,N_40968);
and U41328 (N_41328,N_40738,N_40899);
nor U41329 (N_41329,N_40972,N_40554);
xor U41330 (N_41330,N_40601,N_40096);
or U41331 (N_41331,N_40327,N_40307);
or U41332 (N_41332,N_40183,N_40551);
nand U41333 (N_41333,N_40660,N_40800);
nor U41334 (N_41334,N_40889,N_40111);
or U41335 (N_41335,N_40952,N_40197);
or U41336 (N_41336,N_40418,N_40672);
nand U41337 (N_41337,N_40596,N_40031);
xor U41338 (N_41338,N_40077,N_40211);
nor U41339 (N_41339,N_40573,N_40339);
nand U41340 (N_41340,N_40673,N_40570);
and U41341 (N_41341,N_40578,N_40792);
or U41342 (N_41342,N_40814,N_40171);
or U41343 (N_41343,N_40879,N_40366);
nand U41344 (N_41344,N_40829,N_40683);
nand U41345 (N_41345,N_40168,N_40352);
nand U41346 (N_41346,N_40315,N_40445);
xnor U41347 (N_41347,N_40678,N_40785);
nor U41348 (N_41348,N_40042,N_40840);
nand U41349 (N_41349,N_40483,N_40221);
and U41350 (N_41350,N_40173,N_40582);
and U41351 (N_41351,N_40145,N_40618);
and U41352 (N_41352,N_40716,N_40402);
nor U41353 (N_41353,N_40911,N_40724);
nor U41354 (N_41354,N_40779,N_40392);
and U41355 (N_41355,N_40296,N_40670);
nor U41356 (N_41356,N_40836,N_40172);
nor U41357 (N_41357,N_40242,N_40827);
and U41358 (N_41358,N_40627,N_40353);
xor U41359 (N_41359,N_40103,N_40694);
xnor U41360 (N_41360,N_40712,N_40212);
or U41361 (N_41361,N_40514,N_40830);
xor U41362 (N_41362,N_40629,N_40625);
or U41363 (N_41363,N_40777,N_40969);
and U41364 (N_41364,N_40749,N_40813);
nand U41365 (N_41365,N_40580,N_40847);
and U41366 (N_41366,N_40403,N_40380);
nor U41367 (N_41367,N_40810,N_40961);
and U41368 (N_41368,N_40809,N_40271);
nor U41369 (N_41369,N_40412,N_40818);
nor U41370 (N_41370,N_40364,N_40368);
nor U41371 (N_41371,N_40150,N_40220);
nor U41372 (N_41372,N_40611,N_40938);
or U41373 (N_41373,N_40446,N_40231);
xor U41374 (N_41374,N_40801,N_40264);
and U41375 (N_41375,N_40839,N_40838);
nor U41376 (N_41376,N_40695,N_40638);
nand U41377 (N_41377,N_40822,N_40708);
or U41378 (N_41378,N_40613,N_40563);
or U41379 (N_41379,N_40850,N_40701);
xnor U41380 (N_41380,N_40900,N_40642);
or U41381 (N_41381,N_40789,N_40897);
or U41382 (N_41382,N_40430,N_40021);
nand U41383 (N_41383,N_40763,N_40787);
nor U41384 (N_41384,N_40943,N_40540);
xnor U41385 (N_41385,N_40846,N_40133);
or U41386 (N_41386,N_40409,N_40256);
nand U41387 (N_41387,N_40811,N_40024);
or U41388 (N_41388,N_40158,N_40442);
nand U41389 (N_41389,N_40841,N_40332);
and U41390 (N_41390,N_40295,N_40806);
and U41391 (N_41391,N_40152,N_40038);
or U41392 (N_41392,N_40817,N_40842);
nor U41393 (N_41393,N_40731,N_40186);
or U41394 (N_41394,N_40062,N_40776);
xor U41395 (N_41395,N_40982,N_40855);
or U41396 (N_41396,N_40790,N_40490);
xnor U41397 (N_41397,N_40394,N_40061);
nor U41398 (N_41398,N_40277,N_40356);
or U41399 (N_41399,N_40004,N_40895);
or U41400 (N_41400,N_40089,N_40659);
xor U41401 (N_41401,N_40474,N_40179);
nor U41402 (N_41402,N_40498,N_40674);
nand U41403 (N_41403,N_40504,N_40025);
xor U41404 (N_41404,N_40328,N_40931);
nor U41405 (N_41405,N_40148,N_40166);
nor U41406 (N_41406,N_40130,N_40362);
and U41407 (N_41407,N_40469,N_40893);
and U41408 (N_41408,N_40006,N_40634);
nor U41409 (N_41409,N_40621,N_40962);
nor U41410 (N_41410,N_40805,N_40645);
nand U41411 (N_41411,N_40360,N_40175);
xnor U41412 (N_41412,N_40973,N_40590);
and U41413 (N_41413,N_40316,N_40661);
nor U41414 (N_41414,N_40119,N_40508);
nor U41415 (N_41415,N_40097,N_40227);
nor U41416 (N_41416,N_40276,N_40322);
xnor U41417 (N_41417,N_40755,N_40274);
nor U41418 (N_41418,N_40780,N_40252);
nand U41419 (N_41419,N_40286,N_40688);
and U41420 (N_41420,N_40257,N_40205);
nor U41421 (N_41421,N_40132,N_40663);
xnor U41422 (N_41422,N_40475,N_40641);
nor U41423 (N_41423,N_40184,N_40988);
nor U41424 (N_41424,N_40049,N_40581);
and U41425 (N_41425,N_40951,N_40719);
nand U41426 (N_41426,N_40107,N_40472);
and U41427 (N_41427,N_40669,N_40515);
nand U41428 (N_41428,N_40457,N_40717);
nor U41429 (N_41429,N_40085,N_40555);
nor U41430 (N_41430,N_40202,N_40008);
nor U41431 (N_41431,N_40503,N_40065);
xnor U41432 (N_41432,N_40112,N_40654);
or U41433 (N_41433,N_40317,N_40970);
nor U41434 (N_41434,N_40325,N_40287);
and U41435 (N_41435,N_40571,N_40757);
nand U41436 (N_41436,N_40636,N_40020);
nand U41437 (N_41437,N_40722,N_40545);
nand U41438 (N_41438,N_40373,N_40072);
xnor U41439 (N_41439,N_40671,N_40398);
and U41440 (N_41440,N_40002,N_40324);
and U41441 (N_41441,N_40624,N_40240);
and U41442 (N_41442,N_40604,N_40614);
and U41443 (N_41443,N_40416,N_40696);
nor U41444 (N_41444,N_40238,N_40060);
nand U41445 (N_41445,N_40862,N_40778);
and U41446 (N_41446,N_40761,N_40699);
or U41447 (N_41447,N_40753,N_40123);
xnor U41448 (N_41448,N_40599,N_40980);
and U41449 (N_41449,N_40713,N_40832);
xnor U41450 (N_41450,N_40528,N_40967);
nand U41451 (N_41451,N_40438,N_40583);
and U41452 (N_41452,N_40192,N_40772);
nand U41453 (N_41453,N_40854,N_40557);
nand U41454 (N_41454,N_40516,N_40034);
nor U41455 (N_41455,N_40649,N_40159);
or U41456 (N_41456,N_40279,N_40433);
or U41457 (N_41457,N_40912,N_40471);
or U41458 (N_41458,N_40078,N_40987);
nor U41459 (N_41459,N_40241,N_40957);
xor U41460 (N_41460,N_40068,N_40054);
xor U41461 (N_41461,N_40193,N_40436);
and U41462 (N_41462,N_40203,N_40180);
or U41463 (N_41463,N_40635,N_40727);
and U41464 (N_41464,N_40120,N_40556);
nand U41465 (N_41465,N_40303,N_40343);
and U41466 (N_41466,N_40954,N_40725);
nor U41467 (N_41467,N_40864,N_40828);
xor U41468 (N_41468,N_40612,N_40146);
nor U41469 (N_41469,N_40650,N_40682);
xor U41470 (N_41470,N_40201,N_40321);
or U41471 (N_41471,N_40993,N_40568);
and U41472 (N_41472,N_40117,N_40156);
xnor U41473 (N_41473,N_40500,N_40521);
or U41474 (N_41474,N_40435,N_40947);
xor U41475 (N_41475,N_40574,N_40244);
and U41476 (N_41476,N_40762,N_40478);
xnor U41477 (N_41477,N_40595,N_40401);
and U41478 (N_41478,N_40229,N_40397);
nor U41479 (N_41479,N_40043,N_40447);
nand U41480 (N_41480,N_40291,N_40812);
or U41481 (N_41481,N_40375,N_40933);
nor U41482 (N_41482,N_40539,N_40562);
or U41483 (N_41483,N_40748,N_40512);
or U41484 (N_41484,N_40014,N_40519);
nand U41485 (N_41485,N_40935,N_40101);
and U41486 (N_41486,N_40005,N_40796);
nand U41487 (N_41487,N_40856,N_40094);
xor U41488 (N_41488,N_40218,N_40210);
and U41489 (N_41489,N_40237,N_40759);
and U41490 (N_41490,N_40381,N_40342);
or U41491 (N_41491,N_40788,N_40329);
nand U41492 (N_41492,N_40886,N_40312);
xor U41493 (N_41493,N_40029,N_40309);
xnor U41494 (N_41494,N_40354,N_40209);
nor U41495 (N_41495,N_40348,N_40454);
xnor U41496 (N_41496,N_40565,N_40769);
nand U41497 (N_41497,N_40163,N_40379);
xor U41498 (N_41498,N_40758,N_40766);
and U41499 (N_41499,N_40417,N_40751);
xnor U41500 (N_41500,N_40546,N_40915);
nor U41501 (N_41501,N_40570,N_40386);
nand U41502 (N_41502,N_40168,N_40885);
nor U41503 (N_41503,N_40916,N_40133);
nor U41504 (N_41504,N_40176,N_40756);
and U41505 (N_41505,N_40723,N_40419);
nor U41506 (N_41506,N_40379,N_40287);
xor U41507 (N_41507,N_40499,N_40119);
nand U41508 (N_41508,N_40323,N_40081);
nor U41509 (N_41509,N_40239,N_40541);
or U41510 (N_41510,N_40113,N_40852);
xnor U41511 (N_41511,N_40617,N_40511);
xnor U41512 (N_41512,N_40449,N_40212);
nand U41513 (N_41513,N_40530,N_40700);
or U41514 (N_41514,N_40714,N_40399);
and U41515 (N_41515,N_40570,N_40646);
and U41516 (N_41516,N_40583,N_40348);
nand U41517 (N_41517,N_40300,N_40579);
nand U41518 (N_41518,N_40713,N_40537);
or U41519 (N_41519,N_40911,N_40956);
nand U41520 (N_41520,N_40211,N_40237);
or U41521 (N_41521,N_40965,N_40762);
nor U41522 (N_41522,N_40724,N_40701);
nor U41523 (N_41523,N_40114,N_40970);
nand U41524 (N_41524,N_40149,N_40845);
nor U41525 (N_41525,N_40072,N_40588);
xnor U41526 (N_41526,N_40839,N_40515);
xor U41527 (N_41527,N_40798,N_40727);
or U41528 (N_41528,N_40853,N_40612);
nor U41529 (N_41529,N_40788,N_40461);
and U41530 (N_41530,N_40611,N_40845);
nor U41531 (N_41531,N_40751,N_40515);
nor U41532 (N_41532,N_40320,N_40796);
nand U41533 (N_41533,N_40891,N_40992);
or U41534 (N_41534,N_40522,N_40047);
xor U41535 (N_41535,N_40273,N_40883);
nor U41536 (N_41536,N_40649,N_40353);
or U41537 (N_41537,N_40894,N_40979);
xnor U41538 (N_41538,N_40841,N_40880);
nand U41539 (N_41539,N_40054,N_40195);
nand U41540 (N_41540,N_40772,N_40536);
xor U41541 (N_41541,N_40114,N_40158);
and U41542 (N_41542,N_40614,N_40458);
nand U41543 (N_41543,N_40177,N_40630);
nand U41544 (N_41544,N_40943,N_40968);
nor U41545 (N_41545,N_40665,N_40286);
nor U41546 (N_41546,N_40669,N_40291);
nor U41547 (N_41547,N_40542,N_40122);
nor U41548 (N_41548,N_40440,N_40954);
nand U41549 (N_41549,N_40091,N_40263);
and U41550 (N_41550,N_40057,N_40394);
nand U41551 (N_41551,N_40822,N_40539);
nor U41552 (N_41552,N_40724,N_40912);
nor U41553 (N_41553,N_40668,N_40260);
nand U41554 (N_41554,N_40707,N_40559);
xor U41555 (N_41555,N_40357,N_40459);
and U41556 (N_41556,N_40498,N_40817);
nand U41557 (N_41557,N_40397,N_40773);
nor U41558 (N_41558,N_40144,N_40136);
nor U41559 (N_41559,N_40852,N_40884);
xor U41560 (N_41560,N_40145,N_40851);
and U41561 (N_41561,N_40342,N_40077);
or U41562 (N_41562,N_40630,N_40831);
or U41563 (N_41563,N_40269,N_40160);
nand U41564 (N_41564,N_40196,N_40839);
nand U41565 (N_41565,N_40024,N_40481);
and U41566 (N_41566,N_40334,N_40515);
or U41567 (N_41567,N_40432,N_40451);
nor U41568 (N_41568,N_40372,N_40196);
nand U41569 (N_41569,N_40754,N_40702);
and U41570 (N_41570,N_40565,N_40429);
nand U41571 (N_41571,N_40790,N_40198);
or U41572 (N_41572,N_40254,N_40392);
nor U41573 (N_41573,N_40910,N_40292);
xnor U41574 (N_41574,N_40186,N_40149);
nor U41575 (N_41575,N_40912,N_40441);
and U41576 (N_41576,N_40675,N_40820);
or U41577 (N_41577,N_40368,N_40937);
xor U41578 (N_41578,N_40549,N_40179);
and U41579 (N_41579,N_40205,N_40382);
nand U41580 (N_41580,N_40175,N_40946);
or U41581 (N_41581,N_40459,N_40967);
nor U41582 (N_41582,N_40687,N_40166);
and U41583 (N_41583,N_40312,N_40403);
xor U41584 (N_41584,N_40640,N_40474);
or U41585 (N_41585,N_40805,N_40243);
xor U41586 (N_41586,N_40274,N_40645);
and U41587 (N_41587,N_40321,N_40916);
nor U41588 (N_41588,N_40246,N_40901);
xnor U41589 (N_41589,N_40846,N_40865);
and U41590 (N_41590,N_40670,N_40010);
and U41591 (N_41591,N_40733,N_40653);
nor U41592 (N_41592,N_40699,N_40563);
nor U41593 (N_41593,N_40401,N_40195);
nand U41594 (N_41594,N_40707,N_40542);
xnor U41595 (N_41595,N_40787,N_40824);
nand U41596 (N_41596,N_40926,N_40801);
nor U41597 (N_41597,N_40763,N_40826);
nor U41598 (N_41598,N_40802,N_40056);
nor U41599 (N_41599,N_40000,N_40225);
xor U41600 (N_41600,N_40335,N_40714);
nor U41601 (N_41601,N_40217,N_40780);
or U41602 (N_41602,N_40886,N_40557);
or U41603 (N_41603,N_40961,N_40354);
xor U41604 (N_41604,N_40603,N_40008);
nand U41605 (N_41605,N_40062,N_40220);
nand U41606 (N_41606,N_40749,N_40216);
or U41607 (N_41607,N_40913,N_40625);
nor U41608 (N_41608,N_40986,N_40322);
nand U41609 (N_41609,N_40454,N_40227);
or U41610 (N_41610,N_40317,N_40896);
xor U41611 (N_41611,N_40885,N_40720);
nand U41612 (N_41612,N_40520,N_40675);
nor U41613 (N_41613,N_40871,N_40996);
xnor U41614 (N_41614,N_40791,N_40716);
nand U41615 (N_41615,N_40917,N_40083);
or U41616 (N_41616,N_40093,N_40003);
or U41617 (N_41617,N_40688,N_40460);
nand U41618 (N_41618,N_40266,N_40905);
or U41619 (N_41619,N_40817,N_40588);
xor U41620 (N_41620,N_40665,N_40172);
and U41621 (N_41621,N_40490,N_40090);
xnor U41622 (N_41622,N_40071,N_40942);
nor U41623 (N_41623,N_40036,N_40721);
and U41624 (N_41624,N_40034,N_40074);
nand U41625 (N_41625,N_40362,N_40430);
nand U41626 (N_41626,N_40341,N_40274);
nand U41627 (N_41627,N_40147,N_40330);
nor U41628 (N_41628,N_40525,N_40982);
or U41629 (N_41629,N_40643,N_40704);
xnor U41630 (N_41630,N_40805,N_40372);
or U41631 (N_41631,N_40131,N_40266);
nor U41632 (N_41632,N_40578,N_40647);
or U41633 (N_41633,N_40341,N_40782);
or U41634 (N_41634,N_40981,N_40735);
and U41635 (N_41635,N_40903,N_40059);
or U41636 (N_41636,N_40863,N_40529);
xor U41637 (N_41637,N_40032,N_40366);
nand U41638 (N_41638,N_40231,N_40269);
nand U41639 (N_41639,N_40514,N_40627);
or U41640 (N_41640,N_40436,N_40169);
nor U41641 (N_41641,N_40320,N_40390);
or U41642 (N_41642,N_40906,N_40720);
or U41643 (N_41643,N_40942,N_40516);
nand U41644 (N_41644,N_40513,N_40328);
nor U41645 (N_41645,N_40111,N_40323);
xor U41646 (N_41646,N_40251,N_40359);
nand U41647 (N_41647,N_40895,N_40545);
xor U41648 (N_41648,N_40038,N_40795);
xnor U41649 (N_41649,N_40729,N_40582);
and U41650 (N_41650,N_40407,N_40599);
xnor U41651 (N_41651,N_40023,N_40442);
and U41652 (N_41652,N_40467,N_40695);
and U41653 (N_41653,N_40680,N_40332);
xnor U41654 (N_41654,N_40347,N_40084);
or U41655 (N_41655,N_40165,N_40227);
nor U41656 (N_41656,N_40966,N_40766);
and U41657 (N_41657,N_40814,N_40846);
and U41658 (N_41658,N_40641,N_40771);
xor U41659 (N_41659,N_40699,N_40343);
nor U41660 (N_41660,N_40095,N_40722);
or U41661 (N_41661,N_40796,N_40938);
xnor U41662 (N_41662,N_40116,N_40278);
or U41663 (N_41663,N_40739,N_40284);
nand U41664 (N_41664,N_40991,N_40428);
nor U41665 (N_41665,N_40724,N_40672);
or U41666 (N_41666,N_40750,N_40253);
xnor U41667 (N_41667,N_40717,N_40084);
nor U41668 (N_41668,N_40328,N_40052);
nor U41669 (N_41669,N_40730,N_40895);
xnor U41670 (N_41670,N_40380,N_40783);
or U41671 (N_41671,N_40478,N_40216);
nor U41672 (N_41672,N_40681,N_40412);
nor U41673 (N_41673,N_40865,N_40266);
nand U41674 (N_41674,N_40293,N_40533);
or U41675 (N_41675,N_40800,N_40730);
xnor U41676 (N_41676,N_40885,N_40052);
or U41677 (N_41677,N_40234,N_40014);
xor U41678 (N_41678,N_40253,N_40332);
or U41679 (N_41679,N_40715,N_40177);
and U41680 (N_41680,N_40878,N_40527);
nand U41681 (N_41681,N_40403,N_40959);
nand U41682 (N_41682,N_40435,N_40960);
nand U41683 (N_41683,N_40897,N_40636);
xnor U41684 (N_41684,N_40980,N_40800);
xor U41685 (N_41685,N_40189,N_40136);
and U41686 (N_41686,N_40494,N_40812);
or U41687 (N_41687,N_40090,N_40841);
and U41688 (N_41688,N_40644,N_40732);
xnor U41689 (N_41689,N_40346,N_40361);
or U41690 (N_41690,N_40927,N_40676);
xnor U41691 (N_41691,N_40317,N_40140);
nor U41692 (N_41692,N_40583,N_40483);
xor U41693 (N_41693,N_40807,N_40120);
xnor U41694 (N_41694,N_40773,N_40913);
nand U41695 (N_41695,N_40883,N_40552);
or U41696 (N_41696,N_40963,N_40674);
and U41697 (N_41697,N_40138,N_40130);
and U41698 (N_41698,N_40830,N_40448);
and U41699 (N_41699,N_40499,N_40684);
xnor U41700 (N_41700,N_40076,N_40522);
nand U41701 (N_41701,N_40954,N_40951);
nor U41702 (N_41702,N_40406,N_40109);
nand U41703 (N_41703,N_40542,N_40050);
or U41704 (N_41704,N_40759,N_40069);
or U41705 (N_41705,N_40216,N_40888);
nand U41706 (N_41706,N_40361,N_40549);
xnor U41707 (N_41707,N_40447,N_40498);
xnor U41708 (N_41708,N_40796,N_40570);
nor U41709 (N_41709,N_40563,N_40046);
nor U41710 (N_41710,N_40775,N_40452);
xor U41711 (N_41711,N_40122,N_40613);
nand U41712 (N_41712,N_40383,N_40068);
and U41713 (N_41713,N_40182,N_40445);
or U41714 (N_41714,N_40773,N_40818);
nand U41715 (N_41715,N_40615,N_40033);
or U41716 (N_41716,N_40840,N_40642);
and U41717 (N_41717,N_40592,N_40873);
nor U41718 (N_41718,N_40050,N_40263);
xnor U41719 (N_41719,N_40747,N_40321);
or U41720 (N_41720,N_40960,N_40758);
or U41721 (N_41721,N_40555,N_40820);
nand U41722 (N_41722,N_40973,N_40555);
nor U41723 (N_41723,N_40100,N_40975);
nand U41724 (N_41724,N_40842,N_40690);
xor U41725 (N_41725,N_40754,N_40579);
xor U41726 (N_41726,N_40243,N_40928);
or U41727 (N_41727,N_40909,N_40492);
nand U41728 (N_41728,N_40976,N_40140);
nand U41729 (N_41729,N_40799,N_40368);
nor U41730 (N_41730,N_40850,N_40693);
nor U41731 (N_41731,N_40573,N_40539);
nand U41732 (N_41732,N_40310,N_40352);
or U41733 (N_41733,N_40896,N_40804);
xnor U41734 (N_41734,N_40370,N_40464);
or U41735 (N_41735,N_40021,N_40799);
or U41736 (N_41736,N_40523,N_40542);
xor U41737 (N_41737,N_40485,N_40872);
xor U41738 (N_41738,N_40933,N_40287);
nor U41739 (N_41739,N_40631,N_40657);
xnor U41740 (N_41740,N_40615,N_40958);
and U41741 (N_41741,N_40197,N_40541);
nor U41742 (N_41742,N_40359,N_40960);
and U41743 (N_41743,N_40409,N_40664);
or U41744 (N_41744,N_40336,N_40370);
nor U41745 (N_41745,N_40486,N_40578);
and U41746 (N_41746,N_40931,N_40565);
nor U41747 (N_41747,N_40808,N_40793);
nor U41748 (N_41748,N_40634,N_40250);
nand U41749 (N_41749,N_40535,N_40405);
and U41750 (N_41750,N_40261,N_40495);
nand U41751 (N_41751,N_40243,N_40672);
xnor U41752 (N_41752,N_40721,N_40850);
nor U41753 (N_41753,N_40878,N_40485);
xor U41754 (N_41754,N_40204,N_40379);
xor U41755 (N_41755,N_40310,N_40263);
xor U41756 (N_41756,N_40888,N_40954);
or U41757 (N_41757,N_40316,N_40871);
or U41758 (N_41758,N_40769,N_40634);
or U41759 (N_41759,N_40289,N_40456);
nor U41760 (N_41760,N_40592,N_40385);
xnor U41761 (N_41761,N_40270,N_40723);
or U41762 (N_41762,N_40579,N_40893);
nor U41763 (N_41763,N_40959,N_40745);
nand U41764 (N_41764,N_40161,N_40137);
and U41765 (N_41765,N_40194,N_40496);
or U41766 (N_41766,N_40712,N_40647);
and U41767 (N_41767,N_40930,N_40400);
xnor U41768 (N_41768,N_40441,N_40222);
nor U41769 (N_41769,N_40679,N_40925);
or U41770 (N_41770,N_40468,N_40923);
nand U41771 (N_41771,N_40741,N_40021);
nor U41772 (N_41772,N_40315,N_40761);
nor U41773 (N_41773,N_40898,N_40283);
nand U41774 (N_41774,N_40299,N_40377);
nand U41775 (N_41775,N_40924,N_40191);
nor U41776 (N_41776,N_40093,N_40401);
nor U41777 (N_41777,N_40143,N_40902);
and U41778 (N_41778,N_40515,N_40100);
nor U41779 (N_41779,N_40901,N_40869);
xnor U41780 (N_41780,N_40010,N_40351);
nand U41781 (N_41781,N_40062,N_40591);
nor U41782 (N_41782,N_40868,N_40974);
xor U41783 (N_41783,N_40596,N_40585);
nand U41784 (N_41784,N_40749,N_40390);
or U41785 (N_41785,N_40961,N_40302);
and U41786 (N_41786,N_40029,N_40640);
and U41787 (N_41787,N_40812,N_40483);
xor U41788 (N_41788,N_40401,N_40784);
nand U41789 (N_41789,N_40268,N_40058);
nand U41790 (N_41790,N_40387,N_40653);
nand U41791 (N_41791,N_40535,N_40413);
nor U41792 (N_41792,N_40800,N_40874);
xor U41793 (N_41793,N_40119,N_40837);
nand U41794 (N_41794,N_40978,N_40915);
or U41795 (N_41795,N_40737,N_40224);
and U41796 (N_41796,N_40963,N_40910);
xnor U41797 (N_41797,N_40013,N_40663);
xnor U41798 (N_41798,N_40160,N_40180);
and U41799 (N_41799,N_40012,N_40279);
nor U41800 (N_41800,N_40083,N_40004);
or U41801 (N_41801,N_40556,N_40500);
or U41802 (N_41802,N_40492,N_40757);
nand U41803 (N_41803,N_40666,N_40489);
nor U41804 (N_41804,N_40679,N_40724);
nand U41805 (N_41805,N_40084,N_40177);
nand U41806 (N_41806,N_40298,N_40541);
nand U41807 (N_41807,N_40470,N_40786);
and U41808 (N_41808,N_40904,N_40846);
or U41809 (N_41809,N_40510,N_40790);
nor U41810 (N_41810,N_40849,N_40842);
xor U41811 (N_41811,N_40499,N_40260);
nand U41812 (N_41812,N_40172,N_40887);
nand U41813 (N_41813,N_40415,N_40853);
or U41814 (N_41814,N_40319,N_40535);
nor U41815 (N_41815,N_40768,N_40637);
and U41816 (N_41816,N_40455,N_40991);
nand U41817 (N_41817,N_40065,N_40486);
and U41818 (N_41818,N_40439,N_40040);
or U41819 (N_41819,N_40837,N_40789);
nand U41820 (N_41820,N_40087,N_40841);
nand U41821 (N_41821,N_40522,N_40616);
xor U41822 (N_41822,N_40378,N_40207);
nand U41823 (N_41823,N_40805,N_40236);
nand U41824 (N_41824,N_40724,N_40016);
nor U41825 (N_41825,N_40283,N_40490);
nor U41826 (N_41826,N_40065,N_40366);
and U41827 (N_41827,N_40689,N_40019);
or U41828 (N_41828,N_40943,N_40521);
nand U41829 (N_41829,N_40911,N_40535);
nor U41830 (N_41830,N_40345,N_40637);
nor U41831 (N_41831,N_40866,N_40288);
nand U41832 (N_41832,N_40031,N_40540);
nor U41833 (N_41833,N_40138,N_40572);
or U41834 (N_41834,N_40357,N_40786);
nand U41835 (N_41835,N_40838,N_40636);
nand U41836 (N_41836,N_40785,N_40024);
xnor U41837 (N_41837,N_40885,N_40022);
xor U41838 (N_41838,N_40206,N_40398);
or U41839 (N_41839,N_40286,N_40753);
xor U41840 (N_41840,N_40925,N_40774);
nor U41841 (N_41841,N_40499,N_40354);
and U41842 (N_41842,N_40592,N_40001);
xnor U41843 (N_41843,N_40291,N_40428);
xnor U41844 (N_41844,N_40431,N_40534);
or U41845 (N_41845,N_40762,N_40366);
xnor U41846 (N_41846,N_40874,N_40193);
and U41847 (N_41847,N_40988,N_40343);
or U41848 (N_41848,N_40265,N_40023);
xnor U41849 (N_41849,N_40559,N_40807);
or U41850 (N_41850,N_40606,N_40609);
and U41851 (N_41851,N_40001,N_40073);
or U41852 (N_41852,N_40900,N_40342);
nor U41853 (N_41853,N_40834,N_40609);
nor U41854 (N_41854,N_40836,N_40042);
or U41855 (N_41855,N_40267,N_40376);
nand U41856 (N_41856,N_40237,N_40004);
nor U41857 (N_41857,N_40593,N_40392);
nand U41858 (N_41858,N_40697,N_40690);
nand U41859 (N_41859,N_40032,N_40962);
nand U41860 (N_41860,N_40217,N_40530);
or U41861 (N_41861,N_40633,N_40929);
and U41862 (N_41862,N_40237,N_40190);
or U41863 (N_41863,N_40997,N_40449);
and U41864 (N_41864,N_40893,N_40280);
nor U41865 (N_41865,N_40412,N_40193);
or U41866 (N_41866,N_40723,N_40205);
or U41867 (N_41867,N_40103,N_40773);
nand U41868 (N_41868,N_40190,N_40252);
and U41869 (N_41869,N_40057,N_40575);
nor U41870 (N_41870,N_40675,N_40999);
nand U41871 (N_41871,N_40058,N_40077);
xor U41872 (N_41872,N_40823,N_40277);
nand U41873 (N_41873,N_40434,N_40168);
nor U41874 (N_41874,N_40960,N_40854);
xnor U41875 (N_41875,N_40560,N_40495);
nor U41876 (N_41876,N_40519,N_40101);
nor U41877 (N_41877,N_40644,N_40294);
nor U41878 (N_41878,N_40926,N_40687);
or U41879 (N_41879,N_40174,N_40484);
xor U41880 (N_41880,N_40389,N_40704);
or U41881 (N_41881,N_40842,N_40141);
xor U41882 (N_41882,N_40692,N_40923);
xnor U41883 (N_41883,N_40670,N_40331);
nor U41884 (N_41884,N_40536,N_40945);
nor U41885 (N_41885,N_40607,N_40102);
or U41886 (N_41886,N_40309,N_40053);
nand U41887 (N_41887,N_40664,N_40820);
and U41888 (N_41888,N_40731,N_40100);
xor U41889 (N_41889,N_40173,N_40537);
and U41890 (N_41890,N_40617,N_40527);
nor U41891 (N_41891,N_40694,N_40416);
xor U41892 (N_41892,N_40568,N_40387);
nand U41893 (N_41893,N_40249,N_40533);
nand U41894 (N_41894,N_40377,N_40683);
and U41895 (N_41895,N_40150,N_40148);
xor U41896 (N_41896,N_40610,N_40896);
and U41897 (N_41897,N_40402,N_40233);
nand U41898 (N_41898,N_40347,N_40011);
nor U41899 (N_41899,N_40386,N_40238);
xnor U41900 (N_41900,N_40300,N_40805);
xnor U41901 (N_41901,N_40779,N_40699);
nor U41902 (N_41902,N_40683,N_40954);
nand U41903 (N_41903,N_40139,N_40668);
or U41904 (N_41904,N_40697,N_40406);
and U41905 (N_41905,N_40427,N_40594);
nor U41906 (N_41906,N_40761,N_40894);
or U41907 (N_41907,N_40921,N_40221);
nand U41908 (N_41908,N_40379,N_40416);
nand U41909 (N_41909,N_40814,N_40258);
nor U41910 (N_41910,N_40177,N_40044);
or U41911 (N_41911,N_40024,N_40283);
nand U41912 (N_41912,N_40045,N_40733);
nand U41913 (N_41913,N_40785,N_40185);
nand U41914 (N_41914,N_40137,N_40868);
and U41915 (N_41915,N_40278,N_40638);
nand U41916 (N_41916,N_40085,N_40995);
and U41917 (N_41917,N_40834,N_40007);
or U41918 (N_41918,N_40165,N_40714);
nor U41919 (N_41919,N_40909,N_40187);
nor U41920 (N_41920,N_40473,N_40927);
xor U41921 (N_41921,N_40331,N_40726);
and U41922 (N_41922,N_40507,N_40315);
xnor U41923 (N_41923,N_40407,N_40277);
nor U41924 (N_41924,N_40717,N_40508);
nand U41925 (N_41925,N_40712,N_40922);
nor U41926 (N_41926,N_40896,N_40195);
and U41927 (N_41927,N_40215,N_40299);
nand U41928 (N_41928,N_40277,N_40408);
and U41929 (N_41929,N_40093,N_40315);
nand U41930 (N_41930,N_40403,N_40046);
and U41931 (N_41931,N_40380,N_40754);
xor U41932 (N_41932,N_40835,N_40983);
xor U41933 (N_41933,N_40065,N_40601);
xnor U41934 (N_41934,N_40007,N_40891);
or U41935 (N_41935,N_40506,N_40238);
and U41936 (N_41936,N_40871,N_40241);
xnor U41937 (N_41937,N_40703,N_40244);
nand U41938 (N_41938,N_40354,N_40125);
and U41939 (N_41939,N_40625,N_40941);
and U41940 (N_41940,N_40550,N_40548);
and U41941 (N_41941,N_40211,N_40800);
nor U41942 (N_41942,N_40642,N_40941);
xnor U41943 (N_41943,N_40364,N_40522);
nor U41944 (N_41944,N_40591,N_40498);
xnor U41945 (N_41945,N_40238,N_40129);
and U41946 (N_41946,N_40966,N_40517);
and U41947 (N_41947,N_40043,N_40674);
nor U41948 (N_41948,N_40181,N_40252);
or U41949 (N_41949,N_40741,N_40498);
nor U41950 (N_41950,N_40717,N_40184);
and U41951 (N_41951,N_40473,N_40239);
xor U41952 (N_41952,N_40574,N_40439);
nand U41953 (N_41953,N_40721,N_40994);
and U41954 (N_41954,N_40077,N_40266);
or U41955 (N_41955,N_40278,N_40001);
nand U41956 (N_41956,N_40818,N_40051);
nor U41957 (N_41957,N_40900,N_40690);
and U41958 (N_41958,N_40457,N_40349);
or U41959 (N_41959,N_40487,N_40776);
nand U41960 (N_41960,N_40138,N_40073);
nand U41961 (N_41961,N_40317,N_40234);
nor U41962 (N_41962,N_40961,N_40514);
nor U41963 (N_41963,N_40272,N_40325);
nor U41964 (N_41964,N_40738,N_40458);
xor U41965 (N_41965,N_40504,N_40065);
nand U41966 (N_41966,N_40836,N_40765);
and U41967 (N_41967,N_40264,N_40184);
nand U41968 (N_41968,N_40825,N_40601);
xor U41969 (N_41969,N_40718,N_40795);
or U41970 (N_41970,N_40453,N_40156);
xnor U41971 (N_41971,N_40237,N_40872);
or U41972 (N_41972,N_40032,N_40973);
and U41973 (N_41973,N_40830,N_40822);
nand U41974 (N_41974,N_40934,N_40009);
or U41975 (N_41975,N_40303,N_40723);
or U41976 (N_41976,N_40341,N_40149);
or U41977 (N_41977,N_40879,N_40499);
and U41978 (N_41978,N_40527,N_40054);
and U41979 (N_41979,N_40499,N_40553);
and U41980 (N_41980,N_40350,N_40536);
nor U41981 (N_41981,N_40058,N_40484);
nand U41982 (N_41982,N_40688,N_40764);
nor U41983 (N_41983,N_40884,N_40592);
xor U41984 (N_41984,N_40224,N_40633);
nor U41985 (N_41985,N_40083,N_40825);
xnor U41986 (N_41986,N_40313,N_40605);
or U41987 (N_41987,N_40689,N_40882);
and U41988 (N_41988,N_40030,N_40843);
and U41989 (N_41989,N_40236,N_40700);
nand U41990 (N_41990,N_40976,N_40789);
nor U41991 (N_41991,N_40680,N_40112);
nor U41992 (N_41992,N_40563,N_40305);
xnor U41993 (N_41993,N_40620,N_40521);
nor U41994 (N_41994,N_40857,N_40598);
nor U41995 (N_41995,N_40296,N_40200);
or U41996 (N_41996,N_40108,N_40552);
and U41997 (N_41997,N_40061,N_40810);
nor U41998 (N_41998,N_40764,N_40044);
nor U41999 (N_41999,N_40280,N_40815);
nand U42000 (N_42000,N_41239,N_41416);
and U42001 (N_42001,N_41789,N_41230);
nand U42002 (N_42002,N_41391,N_41659);
and U42003 (N_42003,N_41144,N_41559);
nand U42004 (N_42004,N_41870,N_41014);
and U42005 (N_42005,N_41622,N_41235);
xor U42006 (N_42006,N_41042,N_41977);
or U42007 (N_42007,N_41054,N_41823);
or U42008 (N_42008,N_41343,N_41061);
nor U42009 (N_42009,N_41139,N_41904);
nor U42010 (N_42010,N_41248,N_41808);
nor U42011 (N_42011,N_41147,N_41861);
nand U42012 (N_42012,N_41240,N_41133);
and U42013 (N_42013,N_41306,N_41847);
nor U42014 (N_42014,N_41153,N_41205);
xnor U42015 (N_42015,N_41202,N_41975);
nor U42016 (N_42016,N_41357,N_41413);
and U42017 (N_42017,N_41925,N_41916);
nor U42018 (N_42018,N_41191,N_41149);
and U42019 (N_42019,N_41873,N_41041);
and U42020 (N_42020,N_41378,N_41024);
nand U42021 (N_42021,N_41456,N_41472);
nand U42022 (N_42022,N_41022,N_41715);
nor U42023 (N_42023,N_41933,N_41803);
nand U42024 (N_42024,N_41955,N_41327);
and U42025 (N_42025,N_41880,N_41409);
and U42026 (N_42026,N_41914,N_41613);
and U42027 (N_42027,N_41320,N_41027);
nor U42028 (N_42028,N_41814,N_41636);
or U42029 (N_42029,N_41523,N_41148);
or U42030 (N_42030,N_41099,N_41401);
xnor U42031 (N_42031,N_41295,N_41232);
nand U42032 (N_42032,N_41690,N_41893);
nor U42033 (N_42033,N_41768,N_41918);
nor U42034 (N_42034,N_41967,N_41249);
or U42035 (N_42035,N_41921,N_41553);
nor U42036 (N_42036,N_41582,N_41540);
nor U42037 (N_42037,N_41811,N_41079);
xor U42038 (N_42038,N_41113,N_41822);
nand U42039 (N_42039,N_41476,N_41457);
xor U42040 (N_42040,N_41062,N_41741);
nand U42041 (N_42041,N_41432,N_41009);
nand U42042 (N_42042,N_41256,N_41560);
xnor U42043 (N_42043,N_41723,N_41517);
and U42044 (N_42044,N_41542,N_41280);
or U42045 (N_42045,N_41450,N_41213);
nand U42046 (N_42046,N_41546,N_41005);
nand U42047 (N_42047,N_41352,N_41096);
and U42048 (N_42048,N_41274,N_41544);
and U42049 (N_42049,N_41111,N_41217);
nor U42050 (N_42050,N_41677,N_41052);
xor U42051 (N_42051,N_41045,N_41912);
nor U42052 (N_42052,N_41123,N_41455);
or U42053 (N_42053,N_41349,N_41596);
xor U42054 (N_42054,N_41736,N_41614);
or U42055 (N_42055,N_41120,N_41093);
nand U42056 (N_42056,N_41944,N_41576);
nor U42057 (N_42057,N_41851,N_41465);
nand U42058 (N_42058,N_41109,N_41531);
nand U42059 (N_42059,N_41229,N_41072);
or U42060 (N_42060,N_41490,N_41081);
nor U42061 (N_42061,N_41877,N_41335);
and U42062 (N_42062,N_41610,N_41818);
nor U42063 (N_42063,N_41070,N_41000);
and U42064 (N_42064,N_41685,N_41473);
nor U42065 (N_42065,N_41999,N_41819);
xor U42066 (N_42066,N_41684,N_41404);
xnor U42067 (N_42067,N_41458,N_41693);
or U42068 (N_42068,N_41063,N_41292);
nand U42069 (N_42069,N_41786,N_41155);
and U42070 (N_42070,N_41645,N_41508);
or U42071 (N_42071,N_41825,N_41928);
nand U42072 (N_42072,N_41121,N_41480);
nor U42073 (N_42073,N_41640,N_41087);
or U42074 (N_42074,N_41958,N_41122);
and U42075 (N_42075,N_41011,N_41824);
xnor U42076 (N_42076,N_41915,N_41954);
xor U42077 (N_42077,N_41503,N_41772);
nor U42078 (N_42078,N_41784,N_41058);
nand U42079 (N_42079,N_41782,N_41896);
nor U42080 (N_42080,N_41676,N_41983);
nor U42081 (N_42081,N_41400,N_41262);
or U42082 (N_42082,N_41351,N_41555);
xor U42083 (N_42083,N_41408,N_41737);
or U42084 (N_42084,N_41244,N_41632);
and U42085 (N_42085,N_41639,N_41648);
and U42086 (N_42086,N_41342,N_41220);
and U42087 (N_42087,N_41442,N_41922);
nand U42088 (N_42088,N_41747,N_41510);
xnor U42089 (N_42089,N_41835,N_41010);
nand U42090 (N_42090,N_41477,N_41203);
and U42091 (N_42091,N_41478,N_41209);
xor U42092 (N_42092,N_41359,N_41946);
nand U42093 (N_42093,N_41623,N_41279);
nand U42094 (N_42094,N_41941,N_41278);
or U42095 (N_42095,N_41056,N_41399);
nand U42096 (N_42096,N_41688,N_41532);
or U42097 (N_42097,N_41892,N_41770);
xnor U42098 (N_42098,N_41794,N_41980);
xnor U42099 (N_42099,N_41127,N_41829);
and U42100 (N_42100,N_41382,N_41501);
nor U42101 (N_42101,N_41194,N_41593);
or U42102 (N_42102,N_41034,N_41906);
nor U42103 (N_42103,N_41333,N_41956);
and U42104 (N_42104,N_41475,N_41316);
or U42105 (N_42105,N_41481,N_41700);
nor U42106 (N_42106,N_41431,N_41972);
and U42107 (N_42107,N_41923,N_41579);
or U42108 (N_42108,N_41900,N_41200);
or U42109 (N_42109,N_41107,N_41309);
nand U42110 (N_42110,N_41634,N_41361);
or U42111 (N_42111,N_41360,N_41289);
nor U42112 (N_42112,N_41631,N_41658);
xnor U42113 (N_42113,N_41702,N_41520);
xnor U42114 (N_42114,N_41871,N_41447);
nor U42115 (N_42115,N_41682,N_41545);
nor U42116 (N_42116,N_41143,N_41036);
nor U42117 (N_42117,N_41687,N_41182);
or U42118 (N_42118,N_41304,N_41539);
xnor U42119 (N_42119,N_41943,N_41488);
and U42120 (N_42120,N_41383,N_41964);
nor U42121 (N_42121,N_41367,N_41541);
or U42122 (N_42122,N_41657,N_41603);
and U42123 (N_42123,N_41529,N_41562);
and U42124 (N_42124,N_41298,N_41161);
xnor U42125 (N_42125,N_41722,N_41710);
or U42126 (N_42126,N_41467,N_41032);
nand U42127 (N_42127,N_41831,N_41725);
nand U42128 (N_42128,N_41714,N_41995);
and U42129 (N_42129,N_41841,N_41328);
or U42130 (N_42130,N_41238,N_41565);
xor U42131 (N_42131,N_41556,N_41389);
nand U42132 (N_42132,N_41942,N_41713);
and U42133 (N_42133,N_41988,N_41996);
xnor U42134 (N_42134,N_41007,N_41004);
or U42135 (N_42135,N_41680,N_41176);
xnor U42136 (N_42136,N_41574,N_41745);
or U42137 (N_42137,N_41040,N_41668);
and U42138 (N_42138,N_41805,N_41973);
nor U42139 (N_42139,N_41976,N_41809);
or U42140 (N_42140,N_41064,N_41651);
or U42141 (N_42141,N_41524,N_41245);
nor U42142 (N_42142,N_41842,N_41994);
or U42143 (N_42143,N_41231,N_41429);
xnor U42144 (N_42144,N_41258,N_41718);
and U42145 (N_42145,N_41931,N_41398);
nor U42146 (N_42146,N_41815,N_41852);
nor U42147 (N_42147,N_41655,N_41598);
nand U42148 (N_42148,N_41820,N_41797);
nand U42149 (N_42149,N_41430,N_41885);
nor U42150 (N_42150,N_41577,N_41353);
xor U42151 (N_42151,N_41427,N_41184);
or U42152 (N_42152,N_41635,N_41118);
or U42153 (N_42153,N_41119,N_41165);
nor U42154 (N_42154,N_41204,N_41299);
nor U42155 (N_42155,N_41172,N_41595);
nor U42156 (N_42156,N_41387,N_41750);
and U42157 (N_42157,N_41902,N_41169);
xnor U42158 (N_42158,N_41448,N_41649);
xnor U42159 (N_42159,N_41197,N_41372);
xor U42160 (N_42160,N_41265,N_41028);
nor U42161 (N_42161,N_41834,N_41438);
or U42162 (N_42162,N_41857,N_41901);
nand U42163 (N_42163,N_41526,N_41192);
xnor U42164 (N_42164,N_41848,N_41538);
or U42165 (N_42165,N_41415,N_41908);
or U42166 (N_42166,N_41607,N_41341);
nor U42167 (N_42167,N_41319,N_41307);
nand U42168 (N_42168,N_41895,N_41633);
and U42169 (N_42169,N_41385,N_41969);
xor U42170 (N_42170,N_41729,N_41406);
nand U42171 (N_42171,N_41935,N_41242);
nand U42172 (N_42172,N_41462,N_41832);
or U42173 (N_42173,N_41586,N_41201);
nor U42174 (N_42174,N_41599,N_41074);
xor U42175 (N_42175,N_41086,N_41957);
nand U42176 (N_42176,N_41084,N_41251);
nand U42177 (N_42177,N_41301,N_41218);
or U42178 (N_42178,N_41624,N_41846);
or U42179 (N_42179,N_41920,N_41263);
nor U42180 (N_42180,N_41686,N_41615);
nor U42181 (N_42181,N_41364,N_41717);
xor U42182 (N_42182,N_41154,N_41025);
and U42183 (N_42183,N_41654,N_41215);
nor U42184 (N_42184,N_41573,N_41758);
or U42185 (N_42185,N_41151,N_41816);
nand U42186 (N_42186,N_41570,N_41185);
xor U42187 (N_42187,N_41827,N_41909);
nor U42188 (N_42188,N_41053,N_41675);
nand U42189 (N_42189,N_41105,N_41344);
nand U42190 (N_42190,N_41883,N_41646);
nand U42191 (N_42191,N_41384,N_41392);
and U42192 (N_42192,N_41507,N_41673);
or U42193 (N_42193,N_41858,N_41115);
nor U42194 (N_42194,N_41495,N_41683);
nor U42195 (N_42195,N_41937,N_41754);
nand U42196 (N_42196,N_41002,N_41740);
nand U42197 (N_42197,N_41511,N_41951);
or U42198 (N_42198,N_41311,N_41324);
nor U42199 (N_42199,N_41641,N_41746);
nor U42200 (N_42200,N_41092,N_41696);
and U42201 (N_42201,N_41001,N_41377);
and U42202 (N_42202,N_41221,N_41268);
xor U42203 (N_42203,N_41500,N_41605);
nor U42204 (N_42204,N_41379,N_41939);
nor U42205 (N_42205,N_41496,N_41211);
nand U42206 (N_42206,N_41261,N_41514);
nor U42207 (N_42207,N_41733,N_41046);
nand U42208 (N_42208,N_41287,N_41934);
nor U42209 (N_42209,N_41332,N_41029);
nor U42210 (N_42210,N_41302,N_41876);
nor U42211 (N_42211,N_41469,N_41974);
nor U42212 (N_42212,N_41875,N_41591);
or U42213 (N_42213,N_41358,N_41878);
nor U42214 (N_42214,N_41077,N_41468);
nor U42215 (N_42215,N_41173,N_41106);
xnor U42216 (N_42216,N_41188,N_41076);
or U42217 (N_42217,N_41761,N_41619);
nor U42218 (N_42218,N_41525,N_41608);
and U42219 (N_42219,N_41020,N_41773);
and U42220 (N_42220,N_41826,N_41606);
and U42221 (N_42221,N_41345,N_41348);
nand U42222 (N_42222,N_41919,N_41336);
nand U42223 (N_42223,N_41666,N_41800);
nand U42224 (N_42224,N_41887,N_41466);
xnor U42225 (N_42225,N_41771,N_41869);
and U42226 (N_42226,N_41537,N_41065);
nand U42227 (N_42227,N_41003,N_41445);
nor U42228 (N_42228,N_41752,N_41290);
nand U42229 (N_42229,N_41482,N_41795);
nand U42230 (N_42230,N_41402,N_41435);
nor U42231 (N_42231,N_41990,N_41059);
nand U42232 (N_42232,N_41617,N_41069);
nand U42233 (N_42233,N_41163,N_41927);
xor U42234 (N_42234,N_41938,N_41692);
nor U42235 (N_42235,N_41528,N_41699);
or U42236 (N_42236,N_41769,N_41026);
nor U42237 (N_42237,N_41936,N_41601);
and U42238 (N_42238,N_41303,N_41868);
nor U42239 (N_42239,N_41038,N_41671);
xor U42240 (N_42240,N_41845,N_41561);
or U42241 (N_42241,N_41549,N_41285);
xnor U42242 (N_42242,N_41674,N_41078);
nand U42243 (N_42243,N_41267,N_41724);
and U42244 (N_42244,N_41804,N_41355);
nor U42245 (N_42245,N_41727,N_41798);
xor U42246 (N_42246,N_41899,N_41665);
and U42247 (N_42247,N_41897,N_41571);
nand U42248 (N_42248,N_41732,N_41618);
or U42249 (N_42249,N_41452,N_41864);
and U42250 (N_42250,N_41459,N_41777);
and U42251 (N_42251,N_41247,N_41890);
nor U42252 (N_42252,N_41474,N_41548);
and U42253 (N_42253,N_41305,N_41611);
or U42254 (N_42254,N_41329,N_41283);
or U42255 (N_42255,N_41381,N_41451);
nor U42256 (N_42256,N_41253,N_41720);
xor U42257 (N_42257,N_41584,N_41886);
nor U42258 (N_42258,N_41670,N_41371);
and U42259 (N_42259,N_41494,N_41626);
or U42260 (N_42260,N_41600,N_41806);
xor U42261 (N_42261,N_41222,N_41297);
and U42262 (N_42262,N_41839,N_41663);
or U42263 (N_42263,N_41160,N_41604);
xnor U42264 (N_42264,N_41530,N_41156);
nor U42265 (N_42265,N_41971,N_41136);
or U42266 (N_42266,N_41879,N_41356);
and U42267 (N_42267,N_41021,N_41294);
xnor U42268 (N_42268,N_41694,N_41037);
and U42269 (N_42269,N_41853,N_41346);
nand U42270 (N_42270,N_41872,N_41366);
and U42271 (N_42271,N_41100,N_41585);
or U42272 (N_42272,N_41380,N_41150);
xor U42273 (N_42273,N_41778,N_41592);
xnor U42274 (N_42274,N_41339,N_41254);
xor U42275 (N_42275,N_41266,N_41678);
or U42276 (N_42276,N_41743,N_41330);
nand U42277 (N_42277,N_41763,N_41505);
xnor U42278 (N_42278,N_41110,N_41463);
and U42279 (N_42279,N_41397,N_41924);
xor U42280 (N_42280,N_41479,N_41932);
nand U42281 (N_42281,N_41499,N_41728);
and U42282 (N_42282,N_41891,N_41629);
nand U42283 (N_42283,N_41354,N_41708);
nand U42284 (N_42284,N_41224,N_41566);
nor U42285 (N_42285,N_41533,N_41536);
nand U42286 (N_42286,N_41180,N_41446);
xnor U42287 (N_42287,N_41862,N_41882);
nor U42288 (N_42288,N_41968,N_41170);
nor U42289 (N_42289,N_41206,N_41369);
xnor U42290 (N_42290,N_41102,N_41103);
nand U42291 (N_42291,N_41066,N_41790);
and U42292 (N_42292,N_41198,N_41486);
or U42293 (N_42293,N_41863,N_41216);
nand U42294 (N_42294,N_41581,N_41660);
nand U42295 (N_42295,N_41181,N_41396);
nor U42296 (N_42296,N_41340,N_41228);
nor U42297 (N_42297,N_41960,N_41966);
xor U42298 (N_42298,N_41802,N_41131);
and U42299 (N_42299,N_41594,N_41567);
and U42300 (N_42300,N_41376,N_41347);
and U42301 (N_42301,N_41709,N_41843);
nand U42302 (N_42302,N_41703,N_41855);
or U42303 (N_42303,N_41748,N_41866);
and U42304 (N_42304,N_41874,N_41226);
nor U42305 (N_42305,N_41273,N_41716);
nand U42306 (N_42306,N_41088,N_41705);
and U42307 (N_42307,N_41554,N_41612);
nand U42308 (N_42308,N_41735,N_41774);
xnor U42309 (N_42309,N_41300,N_41669);
or U42310 (N_42310,N_41195,N_41214);
nor U42311 (N_42311,N_41929,N_41625);
nand U42312 (N_42312,N_41141,N_41518);
and U42313 (N_42313,N_41187,N_41425);
xor U42314 (N_42314,N_41410,N_41779);
or U42315 (N_42315,N_41854,N_41982);
or U42316 (N_42316,N_41812,N_41984);
and U42317 (N_42317,N_41656,N_41337);
or U42318 (N_42318,N_41756,N_41453);
and U42319 (N_42319,N_41414,N_41913);
and U42320 (N_42320,N_41753,N_41903);
xor U42321 (N_42321,N_41836,N_41979);
nor U42322 (N_42322,N_41765,N_41085);
and U42323 (N_42323,N_41564,N_41437);
or U42324 (N_42324,N_41580,N_41757);
nor U42325 (N_42325,N_41721,N_41749);
nand U42326 (N_42326,N_41487,N_41365);
nand U42327 (N_42327,N_41998,N_41791);
and U42328 (N_42328,N_41125,N_41023);
xor U42329 (N_42329,N_41859,N_41035);
nor U42330 (N_42330,N_41090,N_41726);
xor U42331 (N_42331,N_41813,N_41807);
or U42332 (N_42332,N_41522,N_41706);
nand U42333 (N_42333,N_41193,N_41830);
or U42334 (N_42334,N_41464,N_41953);
and U42335 (N_42335,N_41884,N_41167);
nand U42336 (N_42336,N_41177,N_41679);
and U42337 (N_42337,N_41428,N_41212);
and U42338 (N_42338,N_41313,N_41697);
nor U42339 (N_42339,N_41060,N_41535);
xor U42340 (N_42340,N_41288,N_41637);
and U42341 (N_42341,N_41403,N_41989);
nand U42342 (N_42342,N_41751,N_41801);
and U42343 (N_42343,N_41949,N_41572);
xnor U42344 (N_42344,N_41616,N_41097);
nand U42345 (N_42345,N_41281,N_41412);
nor U42346 (N_42346,N_41759,N_41276);
nor U42347 (N_42347,N_41208,N_41374);
and U42348 (N_42348,N_41698,N_41436);
and U42349 (N_42349,N_41323,N_41094);
or U42350 (N_42350,N_41134,N_41250);
or U42351 (N_42351,N_41704,N_41417);
nand U42352 (N_42352,N_41158,N_41043);
nor U42353 (N_42353,N_41781,N_41130);
and U42354 (N_42354,N_41867,N_41460);
and U42355 (N_42355,N_41439,N_41444);
xnor U42356 (N_42356,N_41817,N_41098);
and U42357 (N_42357,N_41502,N_41449);
and U42358 (N_42358,N_41661,N_41483);
nand U42359 (N_42359,N_41712,N_41075);
nor U42360 (N_42360,N_41515,N_41521);
nand U42361 (N_42361,N_41563,N_41981);
or U42362 (N_42362,N_41850,N_41926);
or U42363 (N_42363,N_41434,N_41386);
nor U42364 (N_42364,N_41643,N_41057);
xnor U42365 (N_42365,N_41948,N_41575);
nor U42366 (N_42366,N_41609,N_41189);
nand U42367 (N_42367,N_41405,N_41534);
xor U42368 (N_42368,N_41810,N_41856);
nand U42369 (N_42369,N_41650,N_41050);
nor U42370 (N_42370,N_41796,N_41767);
xor U42371 (N_42371,N_41129,N_41785);
nand U42372 (N_42372,N_41159,N_41055);
or U42373 (N_42373,N_41766,N_41498);
nand U42374 (N_42374,N_41260,N_41286);
xor U42375 (N_42375,N_41073,N_41291);
and U42376 (N_42376,N_41638,N_41128);
or U42377 (N_42377,N_41833,N_41373);
xor U42378 (N_42378,N_41089,N_41091);
nor U42379 (N_42379,N_41762,N_41190);
nor U42380 (N_42380,N_41210,N_41621);
or U42381 (N_42381,N_41587,N_41881);
and U42382 (N_42382,N_41667,N_41375);
nor U42383 (N_42383,N_41145,N_41162);
and U42384 (N_42384,N_41219,N_41257);
nand U42385 (N_42385,N_41308,N_41962);
or U42386 (N_42386,N_41742,N_41945);
nor U42387 (N_42387,N_41993,N_41334);
xor U42388 (N_42388,N_41433,N_41992);
xor U42389 (N_42389,N_41997,N_41174);
or U42390 (N_42390,N_41506,N_41930);
nand U42391 (N_42391,N_41178,N_41048);
or U42392 (N_42392,N_41331,N_41558);
nor U42393 (N_42393,N_41828,N_41411);
or U42394 (N_42394,N_41443,N_41047);
nand U42395 (N_42395,N_41440,N_41662);
nor U42396 (N_42396,N_41760,N_41888);
nor U42397 (N_42397,N_41543,N_41689);
or U42398 (N_42398,N_41509,N_41788);
or U42399 (N_42399,N_41252,N_41764);
or U42400 (N_42400,N_41317,N_41039);
xor U42401 (N_42401,N_41272,N_41597);
nor U42402 (N_42402,N_41142,N_41114);
and U42403 (N_42403,N_41860,N_41326);
nor U42404 (N_42404,N_41513,N_41905);
nand U42405 (N_42405,N_41196,N_41424);
and U42406 (N_42406,N_41227,N_41620);
nand U42407 (N_42407,N_41393,N_41321);
nor U42408 (N_42408,N_41739,N_41602);
xor U42409 (N_42409,N_41101,N_41312);
xnor U42410 (N_42410,N_41550,N_41083);
nor U42411 (N_42411,N_41461,N_41527);
or U42412 (N_42412,N_41071,N_41421);
xor U42413 (N_42413,N_41551,N_41259);
or U42414 (N_42414,N_41695,N_41961);
nand U42415 (N_42415,N_41112,N_41454);
xnor U42416 (N_42416,N_41067,N_41277);
and U42417 (N_42417,N_41731,N_41910);
nor U42418 (N_42418,N_41223,N_41783);
nand U42419 (N_42419,N_41730,N_41051);
or U42420 (N_42420,N_41325,N_41590);
nand U42421 (N_42421,N_41171,N_41241);
nor U42422 (N_42422,N_41044,N_41137);
and U42423 (N_42423,N_41865,N_41255);
or U42424 (N_42424,N_41138,N_41246);
or U42425 (N_42425,N_41207,N_41907);
nor U42426 (N_42426,N_41844,N_41168);
nor U42427 (N_42427,N_41030,N_41959);
or U42428 (N_42428,N_41799,N_41965);
xnor U42429 (N_42429,N_41793,N_41963);
nand U42430 (N_42430,N_41701,N_41236);
xnor U42431 (N_42431,N_41950,N_41940);
nor U42432 (N_42432,N_41420,N_41264);
nand U42433 (N_42433,N_41164,N_41707);
and U42434 (N_42434,N_41271,N_41146);
nand U42435 (N_42435,N_41552,N_41653);
nand U42436 (N_42436,N_41642,N_41419);
nand U42437 (N_42437,N_41894,N_41978);
or U42438 (N_42438,N_41837,N_41284);
nand U42439 (N_42439,N_41318,N_41491);
nand U42440 (N_42440,N_41422,N_41987);
nand U42441 (N_42441,N_41719,N_41275);
xnor U42442 (N_42442,N_41080,N_41293);
xor U42443 (N_42443,N_41395,N_41568);
nand U42444 (N_42444,N_41441,N_41296);
xor U42445 (N_42445,N_41183,N_41519);
xnor U42446 (N_42446,N_41407,N_41821);
and U42447 (N_42447,N_41033,N_41787);
xnor U42448 (N_42448,N_41017,N_41755);
or U42449 (N_42449,N_41991,N_41426);
or U42450 (N_42450,N_41484,N_41578);
or U42451 (N_42451,N_41008,N_41124);
or U42452 (N_42452,N_41225,N_41362);
nand U42453 (N_42453,N_41370,N_41985);
and U42454 (N_42454,N_41179,N_41711);
nand U42455 (N_42455,N_41016,N_41497);
or U42456 (N_42456,N_41492,N_41166);
xnor U42457 (N_42457,N_41647,N_41388);
and U42458 (N_42458,N_41776,N_41199);
and U42459 (N_42459,N_41911,N_41282);
nand U42460 (N_42460,N_41547,N_41175);
and U42461 (N_42461,N_41691,N_41006);
and U42462 (N_42462,N_41780,N_41237);
and U42463 (N_42463,N_41234,N_41838);
xor U42464 (N_42464,N_41233,N_41390);
and U42465 (N_42465,N_41588,N_41157);
xnor U42466 (N_42466,N_41350,N_41589);
and U42467 (N_42467,N_41504,N_41117);
xor U42468 (N_42468,N_41310,N_41569);
or U42469 (N_42469,N_41322,N_41630);
nor U42470 (N_42470,N_41644,N_41314);
nor U42471 (N_42471,N_41368,N_41018);
and U42472 (N_42472,N_41917,N_41135);
nor U42473 (N_42473,N_41775,N_41338);
nand U42474 (N_42474,N_41470,N_41840);
or U42475 (N_42475,N_41489,N_41243);
or U42476 (N_42476,N_41418,N_41015);
nand U42477 (N_42477,N_41013,N_41672);
nand U42478 (N_42478,N_41889,N_41898);
xor U42479 (N_42479,N_41628,N_41116);
and U42480 (N_42480,N_41986,N_41792);
or U42481 (N_42481,N_41394,N_41152);
xor U42482 (N_42482,N_41095,N_41140);
and U42483 (N_42483,N_41471,N_41652);
nor U42484 (N_42484,N_41947,N_41315);
nor U42485 (N_42485,N_41132,N_41512);
nand U42486 (N_42486,N_41734,N_41664);
or U42487 (N_42487,N_41849,N_41068);
nand U42488 (N_42488,N_41485,N_41681);
xnor U42489 (N_42489,N_41557,N_41186);
nor U42490 (N_42490,N_41952,N_41049);
nand U42491 (N_42491,N_41031,N_41744);
and U42492 (N_42492,N_41104,N_41423);
and U42493 (N_42493,N_41270,N_41516);
xor U42494 (N_42494,N_41269,N_41493);
xnor U42495 (N_42495,N_41012,N_41970);
and U42496 (N_42496,N_41363,N_41583);
nor U42497 (N_42497,N_41082,N_41738);
nor U42498 (N_42498,N_41126,N_41108);
and U42499 (N_42499,N_41019,N_41627);
or U42500 (N_42500,N_41963,N_41080);
xor U42501 (N_42501,N_41487,N_41311);
and U42502 (N_42502,N_41281,N_41749);
and U42503 (N_42503,N_41888,N_41728);
or U42504 (N_42504,N_41938,N_41720);
and U42505 (N_42505,N_41965,N_41730);
or U42506 (N_42506,N_41800,N_41472);
nor U42507 (N_42507,N_41339,N_41720);
nand U42508 (N_42508,N_41040,N_41932);
and U42509 (N_42509,N_41487,N_41071);
nand U42510 (N_42510,N_41029,N_41919);
nand U42511 (N_42511,N_41306,N_41389);
xnor U42512 (N_42512,N_41101,N_41726);
nand U42513 (N_42513,N_41085,N_41080);
or U42514 (N_42514,N_41073,N_41530);
and U42515 (N_42515,N_41384,N_41144);
and U42516 (N_42516,N_41573,N_41457);
nor U42517 (N_42517,N_41305,N_41733);
or U42518 (N_42518,N_41096,N_41853);
nor U42519 (N_42519,N_41203,N_41381);
nor U42520 (N_42520,N_41395,N_41309);
or U42521 (N_42521,N_41942,N_41568);
xor U42522 (N_42522,N_41473,N_41016);
nand U42523 (N_42523,N_41730,N_41251);
nand U42524 (N_42524,N_41309,N_41577);
xnor U42525 (N_42525,N_41248,N_41094);
and U42526 (N_42526,N_41598,N_41161);
xnor U42527 (N_42527,N_41126,N_41380);
nor U42528 (N_42528,N_41040,N_41058);
xor U42529 (N_42529,N_41199,N_41434);
xor U42530 (N_42530,N_41045,N_41107);
nor U42531 (N_42531,N_41274,N_41950);
nand U42532 (N_42532,N_41983,N_41906);
nor U42533 (N_42533,N_41327,N_41047);
and U42534 (N_42534,N_41824,N_41488);
and U42535 (N_42535,N_41284,N_41370);
and U42536 (N_42536,N_41768,N_41270);
and U42537 (N_42537,N_41281,N_41843);
or U42538 (N_42538,N_41770,N_41584);
xnor U42539 (N_42539,N_41693,N_41334);
nand U42540 (N_42540,N_41414,N_41764);
and U42541 (N_42541,N_41660,N_41821);
xor U42542 (N_42542,N_41814,N_41392);
xnor U42543 (N_42543,N_41143,N_41789);
xor U42544 (N_42544,N_41221,N_41478);
and U42545 (N_42545,N_41162,N_41229);
nor U42546 (N_42546,N_41523,N_41675);
nor U42547 (N_42547,N_41429,N_41965);
or U42548 (N_42548,N_41147,N_41551);
nand U42549 (N_42549,N_41134,N_41903);
and U42550 (N_42550,N_41913,N_41728);
nor U42551 (N_42551,N_41096,N_41874);
xor U42552 (N_42552,N_41367,N_41057);
nor U42553 (N_42553,N_41656,N_41168);
xnor U42554 (N_42554,N_41878,N_41406);
nor U42555 (N_42555,N_41990,N_41141);
nor U42556 (N_42556,N_41339,N_41479);
xnor U42557 (N_42557,N_41771,N_41261);
nand U42558 (N_42558,N_41445,N_41224);
and U42559 (N_42559,N_41981,N_41180);
nor U42560 (N_42560,N_41280,N_41055);
and U42561 (N_42561,N_41641,N_41674);
and U42562 (N_42562,N_41520,N_41168);
nand U42563 (N_42563,N_41710,N_41787);
xor U42564 (N_42564,N_41907,N_41637);
and U42565 (N_42565,N_41549,N_41962);
nor U42566 (N_42566,N_41497,N_41121);
xor U42567 (N_42567,N_41828,N_41180);
or U42568 (N_42568,N_41426,N_41405);
nor U42569 (N_42569,N_41866,N_41045);
or U42570 (N_42570,N_41160,N_41552);
xor U42571 (N_42571,N_41380,N_41188);
nand U42572 (N_42572,N_41697,N_41011);
nand U42573 (N_42573,N_41435,N_41880);
or U42574 (N_42574,N_41916,N_41187);
and U42575 (N_42575,N_41254,N_41559);
nand U42576 (N_42576,N_41320,N_41244);
or U42577 (N_42577,N_41429,N_41230);
xor U42578 (N_42578,N_41465,N_41820);
or U42579 (N_42579,N_41360,N_41886);
or U42580 (N_42580,N_41840,N_41374);
and U42581 (N_42581,N_41444,N_41010);
nor U42582 (N_42582,N_41528,N_41406);
xnor U42583 (N_42583,N_41640,N_41657);
nor U42584 (N_42584,N_41273,N_41943);
or U42585 (N_42585,N_41726,N_41907);
and U42586 (N_42586,N_41707,N_41723);
and U42587 (N_42587,N_41481,N_41519);
xor U42588 (N_42588,N_41806,N_41582);
xor U42589 (N_42589,N_41763,N_41199);
nand U42590 (N_42590,N_41813,N_41871);
nor U42591 (N_42591,N_41448,N_41118);
nand U42592 (N_42592,N_41501,N_41303);
xor U42593 (N_42593,N_41765,N_41492);
xor U42594 (N_42594,N_41722,N_41966);
nand U42595 (N_42595,N_41744,N_41017);
nor U42596 (N_42596,N_41031,N_41289);
xnor U42597 (N_42597,N_41120,N_41234);
nand U42598 (N_42598,N_41242,N_41071);
or U42599 (N_42599,N_41306,N_41797);
nand U42600 (N_42600,N_41162,N_41343);
and U42601 (N_42601,N_41608,N_41153);
xor U42602 (N_42602,N_41433,N_41915);
nor U42603 (N_42603,N_41121,N_41223);
or U42604 (N_42604,N_41158,N_41264);
xor U42605 (N_42605,N_41550,N_41595);
nor U42606 (N_42606,N_41991,N_41807);
nor U42607 (N_42607,N_41826,N_41815);
nor U42608 (N_42608,N_41447,N_41529);
nand U42609 (N_42609,N_41104,N_41535);
nand U42610 (N_42610,N_41480,N_41040);
or U42611 (N_42611,N_41932,N_41460);
xnor U42612 (N_42612,N_41882,N_41928);
and U42613 (N_42613,N_41036,N_41083);
or U42614 (N_42614,N_41319,N_41765);
nor U42615 (N_42615,N_41255,N_41867);
nor U42616 (N_42616,N_41876,N_41021);
and U42617 (N_42617,N_41786,N_41757);
xor U42618 (N_42618,N_41031,N_41329);
or U42619 (N_42619,N_41956,N_41784);
and U42620 (N_42620,N_41218,N_41769);
and U42621 (N_42621,N_41154,N_41042);
or U42622 (N_42622,N_41044,N_41857);
and U42623 (N_42623,N_41856,N_41045);
xnor U42624 (N_42624,N_41161,N_41963);
nor U42625 (N_42625,N_41198,N_41936);
nor U42626 (N_42626,N_41442,N_41189);
nand U42627 (N_42627,N_41984,N_41114);
nor U42628 (N_42628,N_41712,N_41503);
xor U42629 (N_42629,N_41545,N_41090);
xnor U42630 (N_42630,N_41096,N_41105);
nor U42631 (N_42631,N_41677,N_41346);
nand U42632 (N_42632,N_41422,N_41333);
or U42633 (N_42633,N_41874,N_41654);
xnor U42634 (N_42634,N_41671,N_41102);
and U42635 (N_42635,N_41236,N_41458);
nand U42636 (N_42636,N_41383,N_41027);
or U42637 (N_42637,N_41066,N_41429);
and U42638 (N_42638,N_41473,N_41218);
nand U42639 (N_42639,N_41014,N_41184);
xnor U42640 (N_42640,N_41385,N_41479);
xor U42641 (N_42641,N_41260,N_41368);
or U42642 (N_42642,N_41862,N_41093);
or U42643 (N_42643,N_41693,N_41630);
nor U42644 (N_42644,N_41012,N_41517);
nor U42645 (N_42645,N_41759,N_41301);
and U42646 (N_42646,N_41486,N_41842);
nand U42647 (N_42647,N_41050,N_41617);
or U42648 (N_42648,N_41836,N_41873);
xor U42649 (N_42649,N_41441,N_41472);
nor U42650 (N_42650,N_41782,N_41900);
xnor U42651 (N_42651,N_41366,N_41717);
nor U42652 (N_42652,N_41337,N_41679);
nand U42653 (N_42653,N_41039,N_41593);
or U42654 (N_42654,N_41022,N_41654);
nor U42655 (N_42655,N_41329,N_41490);
nand U42656 (N_42656,N_41121,N_41353);
nor U42657 (N_42657,N_41653,N_41676);
or U42658 (N_42658,N_41370,N_41934);
nand U42659 (N_42659,N_41729,N_41901);
xnor U42660 (N_42660,N_41935,N_41460);
nor U42661 (N_42661,N_41445,N_41155);
nor U42662 (N_42662,N_41027,N_41095);
and U42663 (N_42663,N_41047,N_41590);
nor U42664 (N_42664,N_41482,N_41242);
nor U42665 (N_42665,N_41784,N_41405);
nand U42666 (N_42666,N_41290,N_41178);
xnor U42667 (N_42667,N_41569,N_41585);
xor U42668 (N_42668,N_41861,N_41067);
nand U42669 (N_42669,N_41402,N_41064);
or U42670 (N_42670,N_41666,N_41896);
xnor U42671 (N_42671,N_41833,N_41907);
and U42672 (N_42672,N_41457,N_41776);
and U42673 (N_42673,N_41039,N_41360);
xnor U42674 (N_42674,N_41528,N_41659);
nand U42675 (N_42675,N_41736,N_41161);
or U42676 (N_42676,N_41548,N_41374);
nand U42677 (N_42677,N_41400,N_41266);
nor U42678 (N_42678,N_41190,N_41998);
nor U42679 (N_42679,N_41697,N_41030);
nor U42680 (N_42680,N_41131,N_41740);
and U42681 (N_42681,N_41107,N_41586);
or U42682 (N_42682,N_41700,N_41031);
and U42683 (N_42683,N_41898,N_41872);
nor U42684 (N_42684,N_41566,N_41812);
nor U42685 (N_42685,N_41478,N_41823);
and U42686 (N_42686,N_41023,N_41686);
xor U42687 (N_42687,N_41568,N_41699);
and U42688 (N_42688,N_41546,N_41971);
and U42689 (N_42689,N_41666,N_41500);
or U42690 (N_42690,N_41843,N_41195);
xor U42691 (N_42691,N_41167,N_41688);
and U42692 (N_42692,N_41625,N_41276);
and U42693 (N_42693,N_41325,N_41825);
or U42694 (N_42694,N_41740,N_41233);
and U42695 (N_42695,N_41838,N_41081);
nor U42696 (N_42696,N_41470,N_41254);
nand U42697 (N_42697,N_41681,N_41226);
nand U42698 (N_42698,N_41157,N_41168);
nor U42699 (N_42699,N_41880,N_41163);
nand U42700 (N_42700,N_41362,N_41116);
and U42701 (N_42701,N_41736,N_41441);
nor U42702 (N_42702,N_41191,N_41224);
nand U42703 (N_42703,N_41372,N_41468);
nand U42704 (N_42704,N_41729,N_41465);
xnor U42705 (N_42705,N_41094,N_41744);
nor U42706 (N_42706,N_41289,N_41780);
nand U42707 (N_42707,N_41013,N_41032);
and U42708 (N_42708,N_41942,N_41272);
or U42709 (N_42709,N_41057,N_41548);
nand U42710 (N_42710,N_41958,N_41959);
or U42711 (N_42711,N_41670,N_41026);
xnor U42712 (N_42712,N_41189,N_41648);
or U42713 (N_42713,N_41045,N_41138);
and U42714 (N_42714,N_41658,N_41115);
nand U42715 (N_42715,N_41598,N_41719);
or U42716 (N_42716,N_41218,N_41319);
xnor U42717 (N_42717,N_41946,N_41971);
nor U42718 (N_42718,N_41511,N_41907);
nor U42719 (N_42719,N_41713,N_41073);
or U42720 (N_42720,N_41597,N_41218);
xnor U42721 (N_42721,N_41329,N_41301);
xnor U42722 (N_42722,N_41799,N_41564);
nand U42723 (N_42723,N_41104,N_41698);
and U42724 (N_42724,N_41166,N_41692);
nor U42725 (N_42725,N_41299,N_41826);
or U42726 (N_42726,N_41446,N_41344);
or U42727 (N_42727,N_41617,N_41056);
xnor U42728 (N_42728,N_41525,N_41004);
xnor U42729 (N_42729,N_41387,N_41219);
nand U42730 (N_42730,N_41953,N_41927);
nand U42731 (N_42731,N_41216,N_41117);
nand U42732 (N_42732,N_41822,N_41255);
xnor U42733 (N_42733,N_41519,N_41862);
or U42734 (N_42734,N_41368,N_41646);
nor U42735 (N_42735,N_41616,N_41200);
nor U42736 (N_42736,N_41538,N_41362);
xor U42737 (N_42737,N_41428,N_41209);
and U42738 (N_42738,N_41857,N_41397);
and U42739 (N_42739,N_41726,N_41711);
or U42740 (N_42740,N_41001,N_41596);
xnor U42741 (N_42741,N_41043,N_41085);
nor U42742 (N_42742,N_41904,N_41370);
and U42743 (N_42743,N_41099,N_41965);
and U42744 (N_42744,N_41913,N_41619);
xnor U42745 (N_42745,N_41440,N_41116);
nor U42746 (N_42746,N_41176,N_41119);
or U42747 (N_42747,N_41873,N_41909);
or U42748 (N_42748,N_41448,N_41513);
nor U42749 (N_42749,N_41581,N_41049);
and U42750 (N_42750,N_41965,N_41164);
and U42751 (N_42751,N_41496,N_41316);
nor U42752 (N_42752,N_41086,N_41589);
or U42753 (N_42753,N_41194,N_41815);
nor U42754 (N_42754,N_41841,N_41682);
nor U42755 (N_42755,N_41154,N_41545);
nor U42756 (N_42756,N_41270,N_41992);
nor U42757 (N_42757,N_41670,N_41329);
nor U42758 (N_42758,N_41782,N_41850);
and U42759 (N_42759,N_41914,N_41173);
xnor U42760 (N_42760,N_41858,N_41828);
xnor U42761 (N_42761,N_41999,N_41398);
nor U42762 (N_42762,N_41963,N_41302);
and U42763 (N_42763,N_41094,N_41163);
nand U42764 (N_42764,N_41939,N_41789);
nand U42765 (N_42765,N_41967,N_41929);
nor U42766 (N_42766,N_41563,N_41081);
nand U42767 (N_42767,N_41733,N_41536);
or U42768 (N_42768,N_41197,N_41359);
and U42769 (N_42769,N_41320,N_41290);
nand U42770 (N_42770,N_41593,N_41160);
nor U42771 (N_42771,N_41387,N_41776);
nand U42772 (N_42772,N_41267,N_41582);
nand U42773 (N_42773,N_41534,N_41984);
xor U42774 (N_42774,N_41880,N_41230);
xor U42775 (N_42775,N_41724,N_41016);
nor U42776 (N_42776,N_41925,N_41630);
or U42777 (N_42777,N_41556,N_41540);
and U42778 (N_42778,N_41976,N_41786);
nand U42779 (N_42779,N_41022,N_41496);
xor U42780 (N_42780,N_41764,N_41654);
nor U42781 (N_42781,N_41832,N_41826);
and U42782 (N_42782,N_41004,N_41342);
or U42783 (N_42783,N_41427,N_41784);
and U42784 (N_42784,N_41971,N_41627);
xor U42785 (N_42785,N_41114,N_41700);
or U42786 (N_42786,N_41720,N_41949);
xor U42787 (N_42787,N_41446,N_41800);
or U42788 (N_42788,N_41551,N_41308);
nor U42789 (N_42789,N_41275,N_41564);
nor U42790 (N_42790,N_41965,N_41976);
or U42791 (N_42791,N_41098,N_41039);
and U42792 (N_42792,N_41251,N_41780);
or U42793 (N_42793,N_41304,N_41834);
nor U42794 (N_42794,N_41876,N_41913);
or U42795 (N_42795,N_41384,N_41746);
or U42796 (N_42796,N_41586,N_41837);
nand U42797 (N_42797,N_41290,N_41430);
xor U42798 (N_42798,N_41638,N_41494);
xor U42799 (N_42799,N_41711,N_41543);
xnor U42800 (N_42800,N_41841,N_41853);
nand U42801 (N_42801,N_41739,N_41402);
nor U42802 (N_42802,N_41610,N_41820);
xor U42803 (N_42803,N_41702,N_41618);
or U42804 (N_42804,N_41328,N_41413);
nor U42805 (N_42805,N_41353,N_41039);
nand U42806 (N_42806,N_41032,N_41456);
or U42807 (N_42807,N_41577,N_41275);
or U42808 (N_42808,N_41145,N_41692);
nor U42809 (N_42809,N_41175,N_41091);
nand U42810 (N_42810,N_41076,N_41268);
nand U42811 (N_42811,N_41089,N_41120);
and U42812 (N_42812,N_41611,N_41307);
nor U42813 (N_42813,N_41109,N_41587);
xnor U42814 (N_42814,N_41414,N_41775);
or U42815 (N_42815,N_41274,N_41535);
nor U42816 (N_42816,N_41297,N_41351);
nand U42817 (N_42817,N_41133,N_41951);
and U42818 (N_42818,N_41518,N_41990);
or U42819 (N_42819,N_41859,N_41553);
and U42820 (N_42820,N_41757,N_41865);
or U42821 (N_42821,N_41436,N_41272);
xnor U42822 (N_42822,N_41014,N_41370);
or U42823 (N_42823,N_41865,N_41327);
or U42824 (N_42824,N_41760,N_41092);
xor U42825 (N_42825,N_41788,N_41499);
or U42826 (N_42826,N_41181,N_41106);
or U42827 (N_42827,N_41740,N_41972);
or U42828 (N_42828,N_41360,N_41983);
and U42829 (N_42829,N_41879,N_41461);
and U42830 (N_42830,N_41061,N_41014);
nor U42831 (N_42831,N_41044,N_41621);
and U42832 (N_42832,N_41063,N_41436);
nand U42833 (N_42833,N_41924,N_41508);
nor U42834 (N_42834,N_41492,N_41480);
and U42835 (N_42835,N_41771,N_41947);
xor U42836 (N_42836,N_41600,N_41389);
nand U42837 (N_42837,N_41637,N_41291);
xor U42838 (N_42838,N_41270,N_41752);
and U42839 (N_42839,N_41561,N_41481);
nor U42840 (N_42840,N_41474,N_41970);
xnor U42841 (N_42841,N_41103,N_41884);
and U42842 (N_42842,N_41240,N_41354);
nand U42843 (N_42843,N_41530,N_41174);
or U42844 (N_42844,N_41152,N_41710);
and U42845 (N_42845,N_41039,N_41279);
nor U42846 (N_42846,N_41167,N_41324);
and U42847 (N_42847,N_41585,N_41453);
and U42848 (N_42848,N_41835,N_41645);
xnor U42849 (N_42849,N_41212,N_41648);
xnor U42850 (N_42850,N_41323,N_41288);
xor U42851 (N_42851,N_41428,N_41442);
nor U42852 (N_42852,N_41454,N_41581);
or U42853 (N_42853,N_41426,N_41876);
nand U42854 (N_42854,N_41452,N_41635);
nand U42855 (N_42855,N_41685,N_41144);
xnor U42856 (N_42856,N_41566,N_41474);
nor U42857 (N_42857,N_41831,N_41193);
nor U42858 (N_42858,N_41221,N_41611);
nor U42859 (N_42859,N_41162,N_41026);
nand U42860 (N_42860,N_41253,N_41191);
and U42861 (N_42861,N_41420,N_41192);
nor U42862 (N_42862,N_41711,N_41097);
and U42863 (N_42863,N_41374,N_41527);
and U42864 (N_42864,N_41672,N_41637);
and U42865 (N_42865,N_41120,N_41005);
nand U42866 (N_42866,N_41902,N_41237);
nand U42867 (N_42867,N_41912,N_41079);
or U42868 (N_42868,N_41447,N_41532);
nor U42869 (N_42869,N_41719,N_41961);
and U42870 (N_42870,N_41721,N_41362);
nor U42871 (N_42871,N_41374,N_41512);
nor U42872 (N_42872,N_41719,N_41625);
nor U42873 (N_42873,N_41922,N_41256);
or U42874 (N_42874,N_41864,N_41483);
and U42875 (N_42875,N_41292,N_41248);
and U42876 (N_42876,N_41403,N_41798);
and U42877 (N_42877,N_41817,N_41023);
nor U42878 (N_42878,N_41505,N_41825);
and U42879 (N_42879,N_41805,N_41103);
xnor U42880 (N_42880,N_41119,N_41261);
nor U42881 (N_42881,N_41003,N_41897);
or U42882 (N_42882,N_41556,N_41727);
nor U42883 (N_42883,N_41173,N_41062);
nand U42884 (N_42884,N_41342,N_41515);
nand U42885 (N_42885,N_41762,N_41035);
and U42886 (N_42886,N_41917,N_41000);
and U42887 (N_42887,N_41571,N_41794);
nand U42888 (N_42888,N_41489,N_41512);
xor U42889 (N_42889,N_41347,N_41416);
and U42890 (N_42890,N_41008,N_41299);
or U42891 (N_42891,N_41942,N_41428);
nor U42892 (N_42892,N_41540,N_41532);
nor U42893 (N_42893,N_41421,N_41860);
and U42894 (N_42894,N_41522,N_41908);
and U42895 (N_42895,N_41767,N_41305);
and U42896 (N_42896,N_41044,N_41252);
or U42897 (N_42897,N_41505,N_41060);
xnor U42898 (N_42898,N_41379,N_41239);
nor U42899 (N_42899,N_41075,N_41271);
nor U42900 (N_42900,N_41063,N_41585);
or U42901 (N_42901,N_41289,N_41340);
or U42902 (N_42902,N_41849,N_41307);
nand U42903 (N_42903,N_41873,N_41956);
nand U42904 (N_42904,N_41549,N_41214);
xnor U42905 (N_42905,N_41325,N_41980);
xnor U42906 (N_42906,N_41190,N_41545);
and U42907 (N_42907,N_41622,N_41915);
nor U42908 (N_42908,N_41360,N_41098);
xor U42909 (N_42909,N_41354,N_41010);
nor U42910 (N_42910,N_41270,N_41525);
nand U42911 (N_42911,N_41161,N_41908);
and U42912 (N_42912,N_41517,N_41125);
nand U42913 (N_42913,N_41651,N_41154);
nor U42914 (N_42914,N_41034,N_41314);
and U42915 (N_42915,N_41632,N_41207);
or U42916 (N_42916,N_41740,N_41763);
and U42917 (N_42917,N_41059,N_41185);
nor U42918 (N_42918,N_41152,N_41781);
nand U42919 (N_42919,N_41201,N_41113);
nor U42920 (N_42920,N_41709,N_41628);
nand U42921 (N_42921,N_41096,N_41688);
and U42922 (N_42922,N_41162,N_41228);
and U42923 (N_42923,N_41220,N_41145);
xnor U42924 (N_42924,N_41574,N_41067);
nor U42925 (N_42925,N_41235,N_41399);
nand U42926 (N_42926,N_41643,N_41922);
and U42927 (N_42927,N_41108,N_41750);
xor U42928 (N_42928,N_41717,N_41433);
xor U42929 (N_42929,N_41547,N_41917);
or U42930 (N_42930,N_41373,N_41392);
or U42931 (N_42931,N_41771,N_41782);
and U42932 (N_42932,N_41655,N_41081);
nand U42933 (N_42933,N_41869,N_41750);
and U42934 (N_42934,N_41779,N_41968);
nor U42935 (N_42935,N_41459,N_41244);
and U42936 (N_42936,N_41538,N_41049);
nor U42937 (N_42937,N_41058,N_41595);
or U42938 (N_42938,N_41747,N_41143);
and U42939 (N_42939,N_41105,N_41713);
xnor U42940 (N_42940,N_41414,N_41440);
nor U42941 (N_42941,N_41458,N_41423);
and U42942 (N_42942,N_41962,N_41918);
nand U42943 (N_42943,N_41720,N_41107);
nor U42944 (N_42944,N_41528,N_41972);
nand U42945 (N_42945,N_41643,N_41177);
nor U42946 (N_42946,N_41625,N_41128);
nor U42947 (N_42947,N_41138,N_41732);
xnor U42948 (N_42948,N_41907,N_41555);
xnor U42949 (N_42949,N_41428,N_41910);
or U42950 (N_42950,N_41730,N_41717);
nand U42951 (N_42951,N_41047,N_41589);
and U42952 (N_42952,N_41696,N_41677);
nor U42953 (N_42953,N_41003,N_41940);
and U42954 (N_42954,N_41841,N_41034);
and U42955 (N_42955,N_41687,N_41166);
xor U42956 (N_42956,N_41667,N_41941);
nand U42957 (N_42957,N_41869,N_41019);
nor U42958 (N_42958,N_41658,N_41791);
nor U42959 (N_42959,N_41274,N_41668);
nor U42960 (N_42960,N_41170,N_41007);
xnor U42961 (N_42961,N_41933,N_41461);
nor U42962 (N_42962,N_41717,N_41424);
xor U42963 (N_42963,N_41376,N_41888);
xor U42964 (N_42964,N_41371,N_41212);
or U42965 (N_42965,N_41846,N_41867);
or U42966 (N_42966,N_41560,N_41699);
nand U42967 (N_42967,N_41153,N_41393);
xor U42968 (N_42968,N_41712,N_41086);
or U42969 (N_42969,N_41701,N_41655);
or U42970 (N_42970,N_41705,N_41774);
or U42971 (N_42971,N_41993,N_41972);
nand U42972 (N_42972,N_41853,N_41192);
nor U42973 (N_42973,N_41490,N_41461);
nor U42974 (N_42974,N_41603,N_41154);
nor U42975 (N_42975,N_41753,N_41650);
or U42976 (N_42976,N_41072,N_41313);
nor U42977 (N_42977,N_41613,N_41697);
and U42978 (N_42978,N_41882,N_41883);
and U42979 (N_42979,N_41291,N_41536);
nand U42980 (N_42980,N_41055,N_41386);
xnor U42981 (N_42981,N_41427,N_41465);
or U42982 (N_42982,N_41573,N_41747);
nor U42983 (N_42983,N_41310,N_41773);
and U42984 (N_42984,N_41022,N_41648);
or U42985 (N_42985,N_41198,N_41638);
nor U42986 (N_42986,N_41548,N_41117);
and U42987 (N_42987,N_41207,N_41610);
nand U42988 (N_42988,N_41096,N_41716);
nand U42989 (N_42989,N_41047,N_41724);
nor U42990 (N_42990,N_41552,N_41847);
or U42991 (N_42991,N_41338,N_41459);
or U42992 (N_42992,N_41212,N_41845);
or U42993 (N_42993,N_41674,N_41381);
nor U42994 (N_42994,N_41758,N_41587);
nand U42995 (N_42995,N_41819,N_41247);
and U42996 (N_42996,N_41495,N_41223);
nand U42997 (N_42997,N_41905,N_41976);
nor U42998 (N_42998,N_41207,N_41758);
or U42999 (N_42999,N_41447,N_41632);
or U43000 (N_43000,N_42552,N_42455);
nand U43001 (N_43001,N_42219,N_42404);
nand U43002 (N_43002,N_42502,N_42220);
and U43003 (N_43003,N_42900,N_42886);
nor U43004 (N_43004,N_42114,N_42718);
or U43005 (N_43005,N_42462,N_42363);
nand U43006 (N_43006,N_42332,N_42223);
nor U43007 (N_43007,N_42018,N_42344);
or U43008 (N_43008,N_42720,N_42947);
nand U43009 (N_43009,N_42382,N_42784);
xor U43010 (N_43010,N_42724,N_42187);
xor U43011 (N_43011,N_42513,N_42293);
and U43012 (N_43012,N_42297,N_42110);
nand U43013 (N_43013,N_42674,N_42567);
xor U43014 (N_43014,N_42695,N_42470);
xor U43015 (N_43015,N_42681,N_42159);
and U43016 (N_43016,N_42291,N_42744);
and U43017 (N_43017,N_42890,N_42052);
and U43018 (N_43018,N_42583,N_42551);
xor U43019 (N_43019,N_42571,N_42079);
nor U43020 (N_43020,N_42026,N_42765);
or U43021 (N_43021,N_42895,N_42614);
nand U43022 (N_43022,N_42236,N_42168);
nor U43023 (N_43023,N_42885,N_42206);
and U43024 (N_43024,N_42454,N_42190);
nor U43025 (N_43025,N_42202,N_42871);
or U43026 (N_43026,N_42425,N_42437);
nor U43027 (N_43027,N_42867,N_42330);
nand U43028 (N_43028,N_42690,N_42860);
nor U43029 (N_43029,N_42290,N_42530);
xor U43030 (N_43030,N_42682,N_42624);
xnor U43031 (N_43031,N_42420,N_42915);
xnor U43032 (N_43032,N_42034,N_42509);
or U43033 (N_43033,N_42239,N_42679);
nor U43034 (N_43034,N_42800,N_42403);
nor U43035 (N_43035,N_42974,N_42651);
and U43036 (N_43036,N_42556,N_42664);
or U43037 (N_43037,N_42602,N_42625);
and U43038 (N_43038,N_42818,N_42074);
or U43039 (N_43039,N_42268,N_42497);
or U43040 (N_43040,N_42395,N_42662);
xor U43041 (N_43041,N_42192,N_42708);
nor U43042 (N_43042,N_42002,N_42843);
or U43043 (N_43043,N_42914,N_42276);
or U43044 (N_43044,N_42357,N_42542);
or U43045 (N_43045,N_42935,N_42968);
nor U43046 (N_43046,N_42029,N_42274);
or U43047 (N_43047,N_42294,N_42610);
nor U43048 (N_43048,N_42089,N_42253);
nor U43049 (N_43049,N_42468,N_42902);
nand U43050 (N_43050,N_42631,N_42491);
nand U43051 (N_43051,N_42004,N_42917);
and U43052 (N_43052,N_42770,N_42421);
nand U43053 (N_43053,N_42554,N_42036);
nor U43054 (N_43054,N_42921,N_42246);
xor U43055 (N_43055,N_42241,N_42577);
or U43056 (N_43056,N_42597,N_42957);
and U43057 (N_43057,N_42845,N_42217);
or U43058 (N_43058,N_42489,N_42085);
xnor U43059 (N_43059,N_42318,N_42535);
nor U43060 (N_43060,N_42128,N_42066);
nand U43061 (N_43061,N_42482,N_42013);
nand U43062 (N_43062,N_42616,N_42920);
and U43063 (N_43063,N_42989,N_42719);
or U43064 (N_43064,N_42386,N_42568);
nand U43065 (N_43065,N_42317,N_42858);
xor U43066 (N_43066,N_42031,N_42557);
and U43067 (N_43067,N_42229,N_42265);
nand U43068 (N_43068,N_42954,N_42771);
nor U43069 (N_43069,N_42508,N_42767);
nor U43070 (N_43070,N_42832,N_42780);
nor U43071 (N_43071,N_42798,N_42792);
xnor U43072 (N_43072,N_42005,N_42195);
and U43073 (N_43073,N_42545,N_42051);
nand U43074 (N_43074,N_42777,N_42933);
nand U43075 (N_43075,N_42001,N_42901);
xnor U43076 (N_43076,N_42083,N_42151);
or U43077 (N_43077,N_42356,N_42723);
and U43078 (N_43078,N_42650,N_42450);
nand U43079 (N_43079,N_42147,N_42855);
nor U43080 (N_43080,N_42523,N_42279);
nor U43081 (N_43081,N_42918,N_42984);
nand U43082 (N_43082,N_42227,N_42758);
nand U43083 (N_43083,N_42387,N_42113);
nand U43084 (N_43084,N_42562,N_42243);
and U43085 (N_43085,N_42361,N_42928);
and U43086 (N_43086,N_42782,N_42865);
nor U43087 (N_43087,N_42626,N_42053);
xnor U43088 (N_43088,N_42418,N_42775);
and U43089 (N_43089,N_42366,N_42605);
nand U43090 (N_43090,N_42337,N_42995);
or U43091 (N_43091,N_42752,N_42977);
nor U43092 (N_43092,N_42911,N_42226);
or U43093 (N_43093,N_42250,N_42856);
and U43094 (N_43094,N_42133,N_42897);
or U43095 (N_43095,N_42970,N_42656);
xor U43096 (N_43096,N_42586,N_42727);
and U43097 (N_43097,N_42952,N_42949);
xor U43098 (N_43098,N_42547,N_42963);
and U43099 (N_43099,N_42352,N_42678);
nor U43100 (N_43100,N_42641,N_42819);
xor U43101 (N_43101,N_42275,N_42796);
and U43102 (N_43102,N_42177,N_42833);
nor U43103 (N_43103,N_42082,N_42864);
nand U43104 (N_43104,N_42804,N_42311);
nor U43105 (N_43105,N_42196,N_42827);
and U43106 (N_43106,N_42848,N_42390);
xnor U43107 (N_43107,N_42838,N_42010);
or U43108 (N_43108,N_42740,N_42866);
xor U43109 (N_43109,N_42980,N_42126);
nand U43110 (N_43110,N_42966,N_42328);
nor U43111 (N_43111,N_42907,N_42015);
and U43112 (N_43112,N_42197,N_42785);
and U43113 (N_43113,N_42872,N_42267);
or U43114 (N_43114,N_42973,N_42376);
nand U43115 (N_43115,N_42847,N_42378);
xor U43116 (N_43116,N_42255,N_42991);
nor U43117 (N_43117,N_42550,N_42876);
or U43118 (N_43118,N_42590,N_42527);
and U43119 (N_43119,N_42904,N_42913);
xor U43120 (N_43120,N_42233,N_42449);
nor U43121 (N_43121,N_42483,N_42365);
or U43122 (N_43122,N_42433,N_42415);
or U43123 (N_43123,N_42284,N_42086);
nor U43124 (N_43124,N_42639,N_42687);
and U43125 (N_43125,N_42546,N_42116);
or U43126 (N_43126,N_42863,N_42305);
or U43127 (N_43127,N_42242,N_42043);
and U43128 (N_43128,N_42286,N_42228);
and U43129 (N_43129,N_42916,N_42312);
nand U43130 (N_43130,N_42697,N_42071);
nand U43131 (N_43131,N_42014,N_42105);
or U43132 (N_43132,N_42321,N_42417);
and U43133 (N_43133,N_42742,N_42167);
xnor U43134 (N_43134,N_42335,N_42058);
and U43135 (N_43135,N_42778,N_42998);
xnor U43136 (N_43136,N_42214,N_42408);
nand U43137 (N_43137,N_42955,N_42170);
or U43138 (N_43138,N_42982,N_42721);
or U43139 (N_43139,N_42429,N_42373);
nor U43140 (N_43140,N_42346,N_42729);
nor U43141 (N_43141,N_42204,N_42065);
or U43142 (N_43142,N_42815,N_42561);
xor U43143 (N_43143,N_42810,N_42282);
nor U43144 (N_43144,N_42903,N_42097);
xnor U43145 (N_43145,N_42237,N_42288);
nand U43146 (N_43146,N_42306,N_42473);
nor U43147 (N_43147,N_42092,N_42654);
xor U43148 (N_43148,N_42673,N_42983);
nand U43149 (N_43149,N_42038,N_42319);
nor U43150 (N_43150,N_42117,N_42230);
or U43151 (N_43151,N_42613,N_42452);
and U43152 (N_43152,N_42012,N_42157);
or U43153 (N_43153,N_42313,N_42962);
nor U43154 (N_43154,N_42600,N_42943);
or U43155 (N_43155,N_42137,N_42910);
nand U43156 (N_43156,N_42923,N_42559);
nand U43157 (N_43157,N_42340,N_42776);
nand U43158 (N_43158,N_42316,N_42277);
nand U43159 (N_43159,N_42389,N_42440);
and U43160 (N_43160,N_42174,N_42388);
nor U43161 (N_43161,N_42779,N_42503);
or U43162 (N_43162,N_42564,N_42009);
nor U43163 (N_43163,N_42205,N_42802);
nor U43164 (N_43164,N_42033,N_42746);
or U43165 (N_43165,N_42700,N_42121);
nand U43166 (N_43166,N_42385,N_42090);
and U43167 (N_43167,N_42553,N_42353);
or U43168 (N_43168,N_42589,N_42591);
xnor U43169 (N_43169,N_42743,N_42099);
or U43170 (N_43170,N_42495,N_42768);
xor U43171 (N_43171,N_42985,N_42643);
nand U43172 (N_43172,N_42048,N_42181);
nand U43173 (N_43173,N_42381,N_42409);
xor U43174 (N_43174,N_42601,N_42812);
xnor U43175 (N_43175,N_42299,N_42371);
nand U43176 (N_43176,N_42615,N_42272);
xnor U43177 (N_43177,N_42080,N_42307);
nand U43178 (N_43178,N_42140,N_42111);
xor U43179 (N_43179,N_42481,N_42500);
xor U43180 (N_43180,N_42134,N_42176);
xor U43181 (N_43181,N_42262,N_42574);
nand U43182 (N_43182,N_42278,N_42908);
nand U43183 (N_43183,N_42056,N_42607);
and U43184 (N_43184,N_42400,N_42772);
nor U43185 (N_43185,N_42789,N_42880);
nand U43186 (N_43186,N_42541,N_42537);
xnor U43187 (N_43187,N_42100,N_42712);
nand U43188 (N_43188,N_42139,N_42479);
nand U43189 (N_43189,N_42726,N_42380);
or U43190 (N_43190,N_42831,N_42446);
nand U43191 (N_43191,N_42285,N_42922);
nor U43192 (N_43192,N_42103,N_42273);
nor U43193 (N_43193,N_42645,N_42189);
nor U43194 (N_43194,N_42606,N_42135);
or U43195 (N_43195,N_42068,N_42257);
nor U43196 (N_43196,N_42466,N_42788);
and U43197 (N_43197,N_42835,N_42617);
nor U43198 (N_43198,N_42894,N_42016);
or U43199 (N_43199,N_42416,N_42098);
nor U43200 (N_43200,N_42238,N_42830);
and U43201 (N_43201,N_42163,N_42670);
xnor U43202 (N_43202,N_42201,N_42691);
or U43203 (N_43203,N_42837,N_42715);
nand U43204 (N_43204,N_42925,N_42245);
nand U43205 (N_43205,N_42109,N_42164);
and U43206 (N_43206,N_42484,N_42732);
xor U43207 (N_43207,N_42993,N_42347);
and U43208 (N_43208,N_42680,N_42360);
nand U43209 (N_43209,N_42823,N_42608);
nand U43210 (N_43210,N_42839,N_42951);
nand U43211 (N_43211,N_42570,N_42022);
or U43212 (N_43212,N_42756,N_42797);
and U43213 (N_43213,N_42428,N_42999);
nor U43214 (N_43214,N_42851,N_42207);
xnor U43215 (N_43215,N_42899,N_42326);
or U43216 (N_43216,N_42950,N_42534);
and U43217 (N_43217,N_42745,N_42447);
nor U43218 (N_43218,N_42940,N_42668);
and U43219 (N_43219,N_42524,N_42604);
xor U43220 (N_43220,N_42392,N_42735);
and U43221 (N_43221,N_42573,N_42760);
and U43222 (N_43222,N_42493,N_42936);
nand U43223 (N_43223,N_42857,N_42350);
or U43224 (N_43224,N_42424,N_42939);
and U43225 (N_43225,N_42836,N_42741);
xnor U43226 (N_43226,N_42094,N_42076);
nor U43227 (N_43227,N_42292,N_42398);
nor U43228 (N_43228,N_42069,N_42351);
nand U43229 (N_43229,N_42992,N_42423);
xnor U43230 (N_43230,N_42512,N_42793);
or U43231 (N_43231,N_42405,N_42000);
nand U43232 (N_43232,N_42584,N_42208);
nand U43233 (N_43233,N_42023,N_42125);
or U43234 (N_43234,N_42104,N_42677);
xnor U43235 (N_43235,N_42997,N_42507);
and U43236 (N_43236,N_42345,N_42081);
nor U43237 (N_43237,N_42072,N_42006);
nand U43238 (N_43238,N_42302,N_42160);
xnor U43239 (N_43239,N_42769,N_42795);
nand U43240 (N_43240,N_42260,N_42349);
xnor U43241 (N_43241,N_42224,N_42528);
nand U43242 (N_43242,N_42480,N_42419);
nor U43243 (N_43243,N_42870,N_42453);
nor U43244 (N_43244,N_42924,N_42757);
nor U43245 (N_43245,N_42762,N_42790);
and U43246 (N_43246,N_42323,N_42874);
and U43247 (N_43247,N_42598,N_42883);
xor U43248 (N_43248,N_42948,N_42127);
nand U43249 (N_43249,N_42661,N_42298);
nand U43250 (N_43250,N_42696,N_42445);
nand U43251 (N_43251,N_42536,N_42384);
or U43252 (N_43252,N_42088,N_42787);
or U43253 (N_43253,N_42359,N_42548);
or U43254 (N_43254,N_42402,N_42129);
nor U43255 (N_43255,N_42945,N_42410);
or U43256 (N_43256,N_42234,N_42505);
nand U43257 (N_43257,N_42477,N_42039);
nor U43258 (N_43258,N_42158,N_42582);
nand U43259 (N_43259,N_42248,N_42490);
nor U43260 (N_43260,N_42372,N_42969);
nand U43261 (N_43261,N_42426,N_42180);
nor U43262 (N_43262,N_42811,N_42565);
nor U43263 (N_43263,N_42488,N_42879);
nand U43264 (N_43264,N_42136,N_42703);
or U43265 (N_43265,N_42078,N_42967);
or U43266 (N_43266,N_42544,N_42251);
and U43267 (N_43267,N_42165,N_42494);
xnor U43268 (N_43268,N_42225,N_42702);
nor U43269 (N_43269,N_42816,N_42075);
nand U43270 (N_43270,N_42222,N_42689);
or U43271 (N_43271,N_42632,N_42576);
xor U43272 (N_43272,N_42188,N_42522);
xnor U43273 (N_43273,N_42063,N_42514);
nor U43274 (N_43274,N_42432,N_42055);
xor U43275 (N_43275,N_42834,N_42166);
xor U43276 (N_43276,N_42683,N_42152);
or U43277 (N_43277,N_42693,N_42020);
xor U43278 (N_43278,N_42701,N_42976);
and U43279 (N_43279,N_42733,N_42007);
and U43280 (N_43280,N_42391,N_42821);
nand U43281 (N_43281,N_42367,N_42799);
or U43282 (N_43282,N_42132,N_42642);
nor U43283 (N_43283,N_42504,N_42946);
xnor U43284 (N_43284,N_42707,N_42754);
xnor U43285 (N_43285,N_42826,N_42722);
nor U43286 (N_43286,N_42634,N_42774);
and U43287 (N_43287,N_42280,N_42603);
nor U43288 (N_43288,N_42841,N_42411);
and U43289 (N_43289,N_42981,N_42501);
nand U43290 (N_43290,N_42849,N_42336);
nand U43291 (N_43291,N_42394,N_42362);
and U43292 (N_43292,N_42655,N_42252);
nand U43293 (N_43293,N_42711,N_42975);
and U43294 (N_43294,N_42325,N_42518);
nand U43295 (N_43295,N_42049,N_42853);
nor U43296 (N_43296,N_42003,N_42254);
and U43297 (N_43297,N_42783,N_42271);
nor U43298 (N_43298,N_42759,N_42442);
nor U43299 (N_43299,N_42463,N_42266);
or U43300 (N_43300,N_42801,N_42859);
nand U43301 (N_43301,N_42996,N_42964);
and U43302 (N_43302,N_42024,N_42891);
and U43303 (N_43303,N_42730,N_42264);
xnor U43304 (N_43304,N_42327,N_42640);
xnor U43305 (N_43305,N_42706,N_42663);
xnor U43306 (N_43306,N_42169,N_42817);
nor U43307 (N_43307,N_42882,N_42540);
and U43308 (N_43308,N_42084,N_42443);
and U43309 (N_43309,N_42059,N_42764);
or U43310 (N_43310,N_42191,N_42560);
nor U43311 (N_43311,N_42611,N_42295);
and U43312 (N_43312,N_42520,N_42124);
and U43313 (N_43313,N_42358,N_42032);
xor U43314 (N_43314,N_42379,N_42301);
or U43315 (N_43315,N_42814,N_42073);
xnor U43316 (N_43316,N_42529,N_42062);
nor U43317 (N_43317,N_42748,N_42808);
or U43318 (N_43318,N_42183,N_42296);
nor U43319 (N_43319,N_42324,N_42162);
and U43320 (N_43320,N_42587,N_42203);
xnor U43321 (N_43321,N_42101,N_42261);
or U43322 (N_43322,N_42596,N_42216);
or U43323 (N_43323,N_42990,N_42927);
or U43324 (N_43324,N_42822,N_42154);
and U43325 (N_43325,N_42511,N_42460);
nand U43326 (N_43326,N_42657,N_42960);
nand U43327 (N_43327,N_42467,N_42487);
and U43328 (N_43328,N_42303,N_42283);
or U43329 (N_43329,N_42994,N_42829);
or U43330 (N_43330,N_42888,N_42609);
xor U43331 (N_43331,N_42644,N_42308);
nand U43332 (N_43332,N_42093,N_42912);
nor U43333 (N_43333,N_42263,N_42806);
xor U43334 (N_43334,N_42738,N_42348);
nand U43335 (N_43335,N_42413,N_42926);
and U43336 (N_43336,N_42828,N_42739);
and U43337 (N_43337,N_42182,N_42469);
or U43338 (N_43338,N_42566,N_42107);
or U43339 (N_43339,N_42434,N_42892);
or U43340 (N_43340,N_42041,N_42944);
nor U43341 (N_43341,N_42728,N_42737);
nor U43342 (N_43342,N_42593,N_42736);
nand U43343 (N_43343,N_42893,N_42046);
and U43344 (N_43344,N_42304,N_42231);
nor U43345 (N_43345,N_42142,N_42877);
nor U43346 (N_43346,N_42119,N_42212);
nor U43347 (N_43347,N_42377,N_42713);
nor U43348 (N_43348,N_42717,N_42334);
nand U43349 (N_43349,N_42412,N_42199);
nor U43350 (N_43350,N_42025,N_42725);
and U43351 (N_43351,N_42173,N_42149);
or U43352 (N_43352,N_42931,N_42338);
xor U43353 (N_43353,N_42675,N_42840);
or U43354 (N_43354,N_42517,N_42179);
nor U43355 (N_43355,N_42131,N_42569);
nor U43356 (N_43356,N_42249,N_42130);
nor U43357 (N_43357,N_42685,N_42842);
nor U43358 (N_43358,N_42218,N_42145);
or U43359 (N_43359,N_42627,N_42064);
nand U43360 (N_43360,N_42106,N_42956);
or U43361 (N_43361,N_42850,N_42658);
nor U43362 (N_43362,N_42047,N_42716);
nand U43363 (N_43363,N_42499,N_42881);
and U43364 (N_43364,N_42476,N_42938);
and U43365 (N_43365,N_42112,N_42846);
and U43366 (N_43366,N_42986,N_42652);
nand U43367 (N_43367,N_42150,N_42749);
nor U43368 (N_43368,N_42622,N_42676);
nand U43369 (N_43369,N_42269,N_42731);
xnor U43370 (N_43370,N_42057,N_42171);
and U43371 (N_43371,N_42198,N_42809);
or U43372 (N_43372,N_42070,N_42521);
xor U43373 (N_43373,N_42435,N_42232);
or U43374 (N_43374,N_42971,N_42289);
nor U43375 (N_43375,N_42258,N_42118);
nand U43376 (N_43376,N_42035,N_42934);
xor U43377 (N_43377,N_42008,N_42959);
nand U43378 (N_43378,N_42406,N_42077);
and U43379 (N_43379,N_42456,N_42341);
nor U43380 (N_43380,N_42102,N_42786);
and U43381 (N_43381,N_42669,N_42472);
or U43382 (N_43382,N_42138,N_42200);
or U43383 (N_43383,N_42095,N_42813);
xnor U43384 (N_43384,N_42953,N_42464);
or U43385 (N_43385,N_42209,N_42862);
xnor U43386 (N_43386,N_42506,N_42475);
nand U43387 (N_43387,N_42750,N_42580);
nor U43388 (N_43388,N_42988,N_42905);
xor U43389 (N_43389,N_42558,N_42595);
nand U43390 (N_43390,N_42027,N_42710);
nand U43391 (N_43391,N_42623,N_42320);
and U43392 (N_43392,N_42331,N_42630);
xnor U43393 (N_43393,N_42087,N_42649);
and U43394 (N_43394,N_42578,N_42531);
nand U43395 (N_43395,N_42459,N_42184);
nor U43396 (N_43396,N_42734,N_42909);
or U43397 (N_43397,N_42824,N_42898);
nand U43398 (N_43398,N_42144,N_42067);
and U43399 (N_43399,N_42714,N_42213);
xor U43400 (N_43400,N_42875,N_42592);
and U43401 (N_43401,N_42868,N_42575);
nor U43402 (N_43402,N_42538,N_42044);
nor U43403 (N_43403,N_42300,N_42820);
nand U43404 (N_43404,N_42618,N_42021);
xnor U43405 (N_43405,N_42979,N_42873);
or U43406 (N_43406,N_42919,N_42329);
nand U43407 (N_43407,N_42937,N_42515);
and U43408 (N_43408,N_42309,N_42060);
and U43409 (N_43409,N_42599,N_42461);
or U43410 (N_43410,N_42314,N_42671);
nor U43411 (N_43411,N_42355,N_42887);
nor U43412 (N_43412,N_42751,N_42030);
or U43413 (N_43413,N_42343,N_42396);
nor U43414 (N_43414,N_42878,N_42146);
or U43415 (N_43415,N_42186,N_42987);
xor U43416 (N_43416,N_42930,N_42629);
nor U43417 (N_43417,N_42698,N_42122);
or U43418 (N_43418,N_42441,N_42896);
xor U43419 (N_43419,N_42492,N_42439);
nand U43420 (N_43420,N_42761,N_42037);
nand U43421 (N_43421,N_42665,N_42028);
nand U43422 (N_43422,N_42572,N_42854);
nand U43423 (N_43423,N_42638,N_42594);
or U43424 (N_43424,N_42375,N_42451);
or U43425 (N_43425,N_42322,N_42486);
or U43426 (N_43426,N_42436,N_42256);
or U43427 (N_43427,N_42369,N_42247);
xnor U43428 (N_43428,N_42555,N_42393);
or U43429 (N_43429,N_42619,N_42906);
and U43430 (N_43430,N_42210,N_42215);
and U43431 (N_43431,N_42686,N_42794);
xor U43432 (N_43432,N_42667,N_42869);
xnor U43433 (N_43433,N_42444,N_42148);
xnor U43434 (N_43434,N_42143,N_42585);
xor U43435 (N_43435,N_42635,N_42852);
nand U43436 (N_43436,N_42791,N_42496);
nand U43437 (N_43437,N_42120,N_42478);
xor U43438 (N_43438,N_42175,N_42519);
xnor U43439 (N_43439,N_42510,N_42807);
nor U43440 (N_43440,N_42040,N_42108);
and U43441 (N_43441,N_42368,N_42660);
and U43442 (N_43442,N_42684,N_42096);
nand U43443 (N_43443,N_42766,N_42342);
nand U43444 (N_43444,N_42637,N_42978);
nand U43445 (N_43445,N_42932,N_42705);
nor U43446 (N_43446,N_42525,N_42647);
and U43447 (N_43447,N_42045,N_42563);
xor U43448 (N_43448,N_42017,N_42123);
nor U43449 (N_43449,N_42672,N_42763);
nand U43450 (N_43450,N_42235,N_42310);
nand U43451 (N_43451,N_42448,N_42958);
or U43452 (N_43452,N_42339,N_42803);
xnor U43453 (N_43453,N_42471,N_42755);
nand U43454 (N_43454,N_42699,N_42753);
and U43455 (N_43455,N_42153,N_42709);
and U43456 (N_43456,N_42688,N_42704);
xor U43457 (N_43457,N_42884,N_42941);
nand U43458 (N_43458,N_42485,N_42539);
xor U43459 (N_43459,N_42579,N_42648);
nand U43460 (N_43460,N_42370,N_42091);
nand U43461 (N_43461,N_42354,N_42636);
nand U43462 (N_43462,N_42588,N_42465);
nor U43463 (N_43463,N_42178,N_42194);
xnor U43464 (N_43464,N_42430,N_42965);
and U43465 (N_43465,N_42549,N_42621);
nor U43466 (N_43466,N_42259,N_42281);
nand U43467 (N_43467,N_42694,N_42431);
xnor U43468 (N_43468,N_42161,N_42773);
and U43469 (N_43469,N_42414,N_42141);
or U43470 (N_43470,N_42427,N_42516);
nand U43471 (N_43471,N_42155,N_42397);
nand U43472 (N_43472,N_42747,N_42333);
nand U43473 (N_43473,N_42422,N_42438);
nor U43474 (N_43474,N_42399,N_42972);
nor U43475 (N_43475,N_42172,N_42620);
xor U43476 (N_43476,N_42666,N_42861);
and U43477 (N_43477,N_42115,N_42646);
and U43478 (N_43478,N_42458,N_42244);
nand U43479 (N_43479,N_42287,N_42929);
and U43480 (N_43480,N_42193,N_42533);
or U43481 (N_43481,N_42315,N_42211);
xor U43482 (N_43482,N_42532,N_42019);
or U43483 (N_43483,N_42889,N_42054);
xnor U43484 (N_43484,N_42474,N_42612);
and U43485 (N_43485,N_42659,N_42653);
or U43486 (N_43486,N_42270,N_42581);
nand U43487 (N_43487,N_42011,N_42401);
or U43488 (N_43488,N_42383,N_42526);
nor U43489 (N_43489,N_42781,N_42692);
xnor U43490 (N_43490,N_42942,N_42844);
or U43491 (N_43491,N_42628,N_42961);
nand U43492 (N_43492,N_42805,N_42050);
xnor U43493 (N_43493,N_42457,N_42633);
xnor U43494 (N_43494,N_42825,N_42364);
or U43495 (N_43495,N_42042,N_42061);
or U43496 (N_43496,N_42498,N_42221);
and U43497 (N_43497,N_42374,N_42543);
xnor U43498 (N_43498,N_42185,N_42240);
nor U43499 (N_43499,N_42156,N_42407);
nand U43500 (N_43500,N_42427,N_42420);
and U43501 (N_43501,N_42069,N_42236);
or U43502 (N_43502,N_42616,N_42910);
or U43503 (N_43503,N_42633,N_42758);
or U43504 (N_43504,N_42928,N_42340);
and U43505 (N_43505,N_42263,N_42342);
nor U43506 (N_43506,N_42183,N_42241);
xnor U43507 (N_43507,N_42359,N_42081);
or U43508 (N_43508,N_42432,N_42158);
or U43509 (N_43509,N_42159,N_42208);
or U43510 (N_43510,N_42265,N_42594);
or U43511 (N_43511,N_42823,N_42701);
nand U43512 (N_43512,N_42280,N_42279);
or U43513 (N_43513,N_42643,N_42261);
and U43514 (N_43514,N_42988,N_42093);
or U43515 (N_43515,N_42496,N_42079);
xnor U43516 (N_43516,N_42310,N_42978);
xnor U43517 (N_43517,N_42110,N_42177);
nor U43518 (N_43518,N_42085,N_42654);
or U43519 (N_43519,N_42859,N_42957);
or U43520 (N_43520,N_42127,N_42774);
xor U43521 (N_43521,N_42394,N_42679);
nand U43522 (N_43522,N_42322,N_42406);
xor U43523 (N_43523,N_42462,N_42910);
or U43524 (N_43524,N_42303,N_42466);
xor U43525 (N_43525,N_42805,N_42548);
xnor U43526 (N_43526,N_42276,N_42160);
nand U43527 (N_43527,N_42008,N_42273);
xnor U43528 (N_43528,N_42979,N_42658);
and U43529 (N_43529,N_42870,N_42324);
nor U43530 (N_43530,N_42681,N_42431);
or U43531 (N_43531,N_42587,N_42926);
nand U43532 (N_43532,N_42976,N_42317);
nand U43533 (N_43533,N_42976,N_42906);
and U43534 (N_43534,N_42237,N_42572);
or U43535 (N_43535,N_42430,N_42405);
nor U43536 (N_43536,N_42890,N_42256);
or U43537 (N_43537,N_42638,N_42852);
nor U43538 (N_43538,N_42370,N_42328);
xnor U43539 (N_43539,N_42763,N_42003);
nor U43540 (N_43540,N_42215,N_42879);
xnor U43541 (N_43541,N_42477,N_42768);
and U43542 (N_43542,N_42078,N_42854);
nand U43543 (N_43543,N_42838,N_42528);
nor U43544 (N_43544,N_42131,N_42673);
nand U43545 (N_43545,N_42790,N_42861);
nor U43546 (N_43546,N_42747,N_42349);
xor U43547 (N_43547,N_42034,N_42124);
xnor U43548 (N_43548,N_42514,N_42824);
nor U43549 (N_43549,N_42903,N_42048);
xnor U43550 (N_43550,N_42003,N_42289);
xor U43551 (N_43551,N_42128,N_42373);
xor U43552 (N_43552,N_42476,N_42481);
nand U43553 (N_43553,N_42991,N_42851);
xnor U43554 (N_43554,N_42521,N_42710);
nor U43555 (N_43555,N_42582,N_42237);
nor U43556 (N_43556,N_42191,N_42002);
and U43557 (N_43557,N_42025,N_42347);
or U43558 (N_43558,N_42724,N_42253);
xnor U43559 (N_43559,N_42458,N_42864);
nand U43560 (N_43560,N_42195,N_42052);
or U43561 (N_43561,N_42936,N_42114);
and U43562 (N_43562,N_42940,N_42110);
xnor U43563 (N_43563,N_42953,N_42993);
nand U43564 (N_43564,N_42672,N_42865);
nand U43565 (N_43565,N_42019,N_42500);
or U43566 (N_43566,N_42584,N_42813);
nor U43567 (N_43567,N_42161,N_42156);
and U43568 (N_43568,N_42591,N_42850);
nor U43569 (N_43569,N_42328,N_42899);
xor U43570 (N_43570,N_42446,N_42062);
xor U43571 (N_43571,N_42017,N_42893);
and U43572 (N_43572,N_42232,N_42918);
xnor U43573 (N_43573,N_42789,N_42312);
nand U43574 (N_43574,N_42119,N_42199);
nand U43575 (N_43575,N_42503,N_42559);
and U43576 (N_43576,N_42501,N_42067);
nand U43577 (N_43577,N_42684,N_42780);
and U43578 (N_43578,N_42852,N_42675);
nor U43579 (N_43579,N_42874,N_42864);
nand U43580 (N_43580,N_42838,N_42517);
and U43581 (N_43581,N_42861,N_42285);
nor U43582 (N_43582,N_42677,N_42415);
nor U43583 (N_43583,N_42653,N_42270);
nand U43584 (N_43584,N_42822,N_42782);
nand U43585 (N_43585,N_42437,N_42084);
xnor U43586 (N_43586,N_42648,N_42600);
nor U43587 (N_43587,N_42915,N_42482);
xor U43588 (N_43588,N_42444,N_42780);
and U43589 (N_43589,N_42543,N_42103);
nand U43590 (N_43590,N_42107,N_42130);
xor U43591 (N_43591,N_42073,N_42779);
nand U43592 (N_43592,N_42955,N_42163);
nor U43593 (N_43593,N_42165,N_42452);
nor U43594 (N_43594,N_42913,N_42321);
or U43595 (N_43595,N_42981,N_42770);
xnor U43596 (N_43596,N_42960,N_42189);
and U43597 (N_43597,N_42532,N_42642);
xnor U43598 (N_43598,N_42224,N_42435);
nand U43599 (N_43599,N_42179,N_42986);
or U43600 (N_43600,N_42514,N_42918);
and U43601 (N_43601,N_42387,N_42401);
and U43602 (N_43602,N_42517,N_42629);
nor U43603 (N_43603,N_42822,N_42956);
xor U43604 (N_43604,N_42487,N_42274);
nand U43605 (N_43605,N_42457,N_42427);
and U43606 (N_43606,N_42900,N_42481);
or U43607 (N_43607,N_42168,N_42139);
and U43608 (N_43608,N_42583,N_42553);
nor U43609 (N_43609,N_42676,N_42885);
nand U43610 (N_43610,N_42869,N_42935);
xor U43611 (N_43611,N_42060,N_42398);
nand U43612 (N_43612,N_42015,N_42994);
nand U43613 (N_43613,N_42872,N_42095);
nor U43614 (N_43614,N_42001,N_42805);
nand U43615 (N_43615,N_42959,N_42697);
nor U43616 (N_43616,N_42956,N_42035);
xor U43617 (N_43617,N_42771,N_42213);
xnor U43618 (N_43618,N_42128,N_42453);
and U43619 (N_43619,N_42223,N_42356);
xor U43620 (N_43620,N_42892,N_42244);
or U43621 (N_43621,N_42231,N_42458);
or U43622 (N_43622,N_42879,N_42162);
xor U43623 (N_43623,N_42565,N_42601);
nor U43624 (N_43624,N_42198,N_42080);
nand U43625 (N_43625,N_42675,N_42359);
and U43626 (N_43626,N_42490,N_42247);
nor U43627 (N_43627,N_42149,N_42320);
nand U43628 (N_43628,N_42359,N_42302);
or U43629 (N_43629,N_42444,N_42142);
or U43630 (N_43630,N_42272,N_42789);
nand U43631 (N_43631,N_42454,N_42935);
and U43632 (N_43632,N_42143,N_42570);
or U43633 (N_43633,N_42191,N_42253);
nor U43634 (N_43634,N_42648,N_42322);
xnor U43635 (N_43635,N_42249,N_42325);
nor U43636 (N_43636,N_42838,N_42670);
nor U43637 (N_43637,N_42075,N_42941);
or U43638 (N_43638,N_42561,N_42769);
or U43639 (N_43639,N_42198,N_42948);
nor U43640 (N_43640,N_42849,N_42461);
or U43641 (N_43641,N_42021,N_42456);
and U43642 (N_43642,N_42765,N_42067);
nand U43643 (N_43643,N_42676,N_42223);
or U43644 (N_43644,N_42190,N_42145);
and U43645 (N_43645,N_42602,N_42657);
and U43646 (N_43646,N_42292,N_42579);
nor U43647 (N_43647,N_42992,N_42016);
nor U43648 (N_43648,N_42196,N_42007);
or U43649 (N_43649,N_42871,N_42996);
and U43650 (N_43650,N_42436,N_42866);
nor U43651 (N_43651,N_42232,N_42903);
and U43652 (N_43652,N_42078,N_42808);
nand U43653 (N_43653,N_42641,N_42856);
nor U43654 (N_43654,N_42202,N_42550);
or U43655 (N_43655,N_42179,N_42204);
and U43656 (N_43656,N_42499,N_42699);
or U43657 (N_43657,N_42502,N_42787);
and U43658 (N_43658,N_42431,N_42408);
or U43659 (N_43659,N_42215,N_42358);
nor U43660 (N_43660,N_42575,N_42783);
xor U43661 (N_43661,N_42997,N_42821);
and U43662 (N_43662,N_42912,N_42515);
xnor U43663 (N_43663,N_42833,N_42482);
nor U43664 (N_43664,N_42425,N_42565);
and U43665 (N_43665,N_42600,N_42893);
nor U43666 (N_43666,N_42929,N_42184);
nor U43667 (N_43667,N_42226,N_42711);
xnor U43668 (N_43668,N_42659,N_42555);
nor U43669 (N_43669,N_42095,N_42396);
xnor U43670 (N_43670,N_42858,N_42095);
nor U43671 (N_43671,N_42759,N_42626);
nor U43672 (N_43672,N_42055,N_42128);
or U43673 (N_43673,N_42350,N_42517);
xor U43674 (N_43674,N_42651,N_42479);
nand U43675 (N_43675,N_42322,N_42659);
nor U43676 (N_43676,N_42617,N_42606);
nor U43677 (N_43677,N_42013,N_42769);
nor U43678 (N_43678,N_42505,N_42694);
nand U43679 (N_43679,N_42300,N_42877);
or U43680 (N_43680,N_42160,N_42140);
xor U43681 (N_43681,N_42906,N_42337);
xnor U43682 (N_43682,N_42671,N_42655);
nor U43683 (N_43683,N_42601,N_42376);
xnor U43684 (N_43684,N_42954,N_42956);
xnor U43685 (N_43685,N_42489,N_42763);
or U43686 (N_43686,N_42803,N_42946);
nor U43687 (N_43687,N_42891,N_42763);
and U43688 (N_43688,N_42080,N_42012);
nand U43689 (N_43689,N_42884,N_42943);
xnor U43690 (N_43690,N_42783,N_42243);
xor U43691 (N_43691,N_42105,N_42715);
or U43692 (N_43692,N_42061,N_42152);
and U43693 (N_43693,N_42508,N_42844);
nor U43694 (N_43694,N_42112,N_42994);
and U43695 (N_43695,N_42275,N_42045);
nand U43696 (N_43696,N_42928,N_42378);
or U43697 (N_43697,N_42497,N_42237);
xor U43698 (N_43698,N_42960,N_42698);
nand U43699 (N_43699,N_42871,N_42761);
nor U43700 (N_43700,N_42637,N_42233);
nor U43701 (N_43701,N_42693,N_42248);
and U43702 (N_43702,N_42119,N_42944);
xnor U43703 (N_43703,N_42764,N_42454);
and U43704 (N_43704,N_42114,N_42672);
or U43705 (N_43705,N_42931,N_42190);
or U43706 (N_43706,N_42352,N_42561);
nor U43707 (N_43707,N_42783,N_42374);
and U43708 (N_43708,N_42071,N_42954);
nor U43709 (N_43709,N_42123,N_42586);
xnor U43710 (N_43710,N_42612,N_42988);
nor U43711 (N_43711,N_42856,N_42236);
xor U43712 (N_43712,N_42166,N_42381);
or U43713 (N_43713,N_42379,N_42716);
nand U43714 (N_43714,N_42479,N_42400);
nand U43715 (N_43715,N_42956,N_42413);
nor U43716 (N_43716,N_42454,N_42276);
xor U43717 (N_43717,N_42857,N_42074);
and U43718 (N_43718,N_42227,N_42424);
nor U43719 (N_43719,N_42181,N_42030);
or U43720 (N_43720,N_42595,N_42930);
or U43721 (N_43721,N_42208,N_42739);
nand U43722 (N_43722,N_42302,N_42982);
nor U43723 (N_43723,N_42282,N_42352);
xor U43724 (N_43724,N_42262,N_42697);
nand U43725 (N_43725,N_42312,N_42992);
nand U43726 (N_43726,N_42782,N_42649);
or U43727 (N_43727,N_42384,N_42948);
xnor U43728 (N_43728,N_42312,N_42174);
or U43729 (N_43729,N_42477,N_42542);
nor U43730 (N_43730,N_42337,N_42361);
nor U43731 (N_43731,N_42764,N_42637);
nor U43732 (N_43732,N_42841,N_42516);
nor U43733 (N_43733,N_42610,N_42118);
or U43734 (N_43734,N_42463,N_42051);
nor U43735 (N_43735,N_42104,N_42729);
nand U43736 (N_43736,N_42088,N_42933);
or U43737 (N_43737,N_42474,N_42165);
nand U43738 (N_43738,N_42030,N_42300);
nand U43739 (N_43739,N_42036,N_42297);
nor U43740 (N_43740,N_42979,N_42047);
nand U43741 (N_43741,N_42462,N_42901);
xor U43742 (N_43742,N_42650,N_42691);
nand U43743 (N_43743,N_42477,N_42174);
nor U43744 (N_43744,N_42677,N_42887);
xnor U43745 (N_43745,N_42081,N_42286);
or U43746 (N_43746,N_42496,N_42377);
or U43747 (N_43747,N_42462,N_42102);
nor U43748 (N_43748,N_42033,N_42368);
xnor U43749 (N_43749,N_42105,N_42783);
nor U43750 (N_43750,N_42870,N_42294);
nor U43751 (N_43751,N_42868,N_42283);
nand U43752 (N_43752,N_42464,N_42758);
or U43753 (N_43753,N_42457,N_42994);
nor U43754 (N_43754,N_42025,N_42072);
and U43755 (N_43755,N_42893,N_42938);
and U43756 (N_43756,N_42047,N_42421);
xor U43757 (N_43757,N_42734,N_42963);
nor U43758 (N_43758,N_42344,N_42551);
nor U43759 (N_43759,N_42075,N_42238);
xor U43760 (N_43760,N_42850,N_42823);
nand U43761 (N_43761,N_42894,N_42390);
or U43762 (N_43762,N_42077,N_42084);
xor U43763 (N_43763,N_42174,N_42517);
or U43764 (N_43764,N_42086,N_42478);
nand U43765 (N_43765,N_42848,N_42095);
xnor U43766 (N_43766,N_42966,N_42343);
or U43767 (N_43767,N_42575,N_42773);
or U43768 (N_43768,N_42199,N_42098);
and U43769 (N_43769,N_42051,N_42082);
and U43770 (N_43770,N_42896,N_42254);
nor U43771 (N_43771,N_42605,N_42109);
nand U43772 (N_43772,N_42780,N_42792);
nor U43773 (N_43773,N_42739,N_42753);
xnor U43774 (N_43774,N_42659,N_42854);
nand U43775 (N_43775,N_42860,N_42793);
nand U43776 (N_43776,N_42735,N_42225);
nand U43777 (N_43777,N_42143,N_42223);
nor U43778 (N_43778,N_42996,N_42805);
nand U43779 (N_43779,N_42667,N_42304);
nand U43780 (N_43780,N_42478,N_42827);
nand U43781 (N_43781,N_42574,N_42428);
xor U43782 (N_43782,N_42187,N_42345);
nor U43783 (N_43783,N_42892,N_42354);
nand U43784 (N_43784,N_42682,N_42189);
or U43785 (N_43785,N_42867,N_42626);
or U43786 (N_43786,N_42061,N_42564);
nand U43787 (N_43787,N_42807,N_42161);
nor U43788 (N_43788,N_42877,N_42581);
xnor U43789 (N_43789,N_42341,N_42576);
xnor U43790 (N_43790,N_42912,N_42023);
nand U43791 (N_43791,N_42682,N_42683);
nand U43792 (N_43792,N_42230,N_42026);
and U43793 (N_43793,N_42693,N_42958);
or U43794 (N_43794,N_42539,N_42230);
nor U43795 (N_43795,N_42147,N_42828);
and U43796 (N_43796,N_42255,N_42908);
nand U43797 (N_43797,N_42945,N_42974);
xor U43798 (N_43798,N_42497,N_42590);
or U43799 (N_43799,N_42654,N_42048);
and U43800 (N_43800,N_42676,N_42391);
nand U43801 (N_43801,N_42410,N_42759);
or U43802 (N_43802,N_42940,N_42123);
and U43803 (N_43803,N_42013,N_42418);
xor U43804 (N_43804,N_42540,N_42530);
and U43805 (N_43805,N_42438,N_42227);
xnor U43806 (N_43806,N_42638,N_42891);
xor U43807 (N_43807,N_42325,N_42062);
xor U43808 (N_43808,N_42878,N_42952);
xnor U43809 (N_43809,N_42729,N_42872);
or U43810 (N_43810,N_42333,N_42752);
or U43811 (N_43811,N_42345,N_42158);
nand U43812 (N_43812,N_42653,N_42873);
xnor U43813 (N_43813,N_42887,N_42559);
nand U43814 (N_43814,N_42387,N_42092);
nor U43815 (N_43815,N_42942,N_42175);
nand U43816 (N_43816,N_42794,N_42621);
nand U43817 (N_43817,N_42605,N_42242);
nand U43818 (N_43818,N_42529,N_42210);
xnor U43819 (N_43819,N_42195,N_42635);
nor U43820 (N_43820,N_42010,N_42007);
and U43821 (N_43821,N_42399,N_42689);
or U43822 (N_43822,N_42475,N_42892);
or U43823 (N_43823,N_42974,N_42319);
and U43824 (N_43824,N_42650,N_42381);
and U43825 (N_43825,N_42793,N_42952);
or U43826 (N_43826,N_42207,N_42428);
and U43827 (N_43827,N_42226,N_42776);
or U43828 (N_43828,N_42309,N_42036);
nor U43829 (N_43829,N_42753,N_42471);
xor U43830 (N_43830,N_42794,N_42259);
nand U43831 (N_43831,N_42283,N_42040);
nor U43832 (N_43832,N_42279,N_42737);
and U43833 (N_43833,N_42170,N_42752);
xor U43834 (N_43834,N_42018,N_42644);
nand U43835 (N_43835,N_42270,N_42958);
and U43836 (N_43836,N_42833,N_42400);
and U43837 (N_43837,N_42716,N_42771);
nand U43838 (N_43838,N_42633,N_42638);
or U43839 (N_43839,N_42770,N_42917);
nor U43840 (N_43840,N_42557,N_42045);
nor U43841 (N_43841,N_42553,N_42442);
and U43842 (N_43842,N_42262,N_42924);
and U43843 (N_43843,N_42283,N_42062);
and U43844 (N_43844,N_42232,N_42397);
nor U43845 (N_43845,N_42263,N_42065);
and U43846 (N_43846,N_42796,N_42885);
nand U43847 (N_43847,N_42357,N_42781);
xor U43848 (N_43848,N_42505,N_42109);
nor U43849 (N_43849,N_42632,N_42370);
nand U43850 (N_43850,N_42915,N_42831);
nor U43851 (N_43851,N_42431,N_42432);
nand U43852 (N_43852,N_42939,N_42363);
or U43853 (N_43853,N_42662,N_42251);
nand U43854 (N_43854,N_42989,N_42185);
xnor U43855 (N_43855,N_42345,N_42890);
xnor U43856 (N_43856,N_42013,N_42965);
nand U43857 (N_43857,N_42412,N_42517);
nand U43858 (N_43858,N_42123,N_42104);
xnor U43859 (N_43859,N_42078,N_42868);
xor U43860 (N_43860,N_42235,N_42221);
or U43861 (N_43861,N_42830,N_42367);
and U43862 (N_43862,N_42938,N_42990);
nand U43863 (N_43863,N_42760,N_42046);
xnor U43864 (N_43864,N_42154,N_42555);
xor U43865 (N_43865,N_42470,N_42001);
nor U43866 (N_43866,N_42456,N_42243);
and U43867 (N_43867,N_42499,N_42393);
nor U43868 (N_43868,N_42905,N_42062);
and U43869 (N_43869,N_42619,N_42801);
nor U43870 (N_43870,N_42815,N_42095);
nand U43871 (N_43871,N_42043,N_42706);
nor U43872 (N_43872,N_42303,N_42319);
xnor U43873 (N_43873,N_42844,N_42873);
xnor U43874 (N_43874,N_42426,N_42991);
nand U43875 (N_43875,N_42620,N_42870);
xnor U43876 (N_43876,N_42775,N_42782);
or U43877 (N_43877,N_42820,N_42368);
or U43878 (N_43878,N_42525,N_42236);
xor U43879 (N_43879,N_42500,N_42981);
xnor U43880 (N_43880,N_42185,N_42492);
or U43881 (N_43881,N_42292,N_42996);
nand U43882 (N_43882,N_42201,N_42014);
xnor U43883 (N_43883,N_42899,N_42817);
nor U43884 (N_43884,N_42685,N_42031);
nor U43885 (N_43885,N_42129,N_42904);
xnor U43886 (N_43886,N_42154,N_42160);
xnor U43887 (N_43887,N_42509,N_42711);
xnor U43888 (N_43888,N_42211,N_42937);
and U43889 (N_43889,N_42097,N_42848);
xnor U43890 (N_43890,N_42981,N_42557);
nand U43891 (N_43891,N_42004,N_42141);
nand U43892 (N_43892,N_42913,N_42849);
nor U43893 (N_43893,N_42792,N_42542);
and U43894 (N_43894,N_42812,N_42207);
and U43895 (N_43895,N_42314,N_42140);
and U43896 (N_43896,N_42539,N_42238);
nor U43897 (N_43897,N_42183,N_42777);
nor U43898 (N_43898,N_42366,N_42775);
nand U43899 (N_43899,N_42576,N_42754);
nor U43900 (N_43900,N_42342,N_42266);
nor U43901 (N_43901,N_42858,N_42186);
or U43902 (N_43902,N_42786,N_42469);
xor U43903 (N_43903,N_42548,N_42553);
nor U43904 (N_43904,N_42194,N_42649);
nor U43905 (N_43905,N_42127,N_42662);
nor U43906 (N_43906,N_42985,N_42837);
nor U43907 (N_43907,N_42407,N_42072);
nand U43908 (N_43908,N_42667,N_42099);
or U43909 (N_43909,N_42397,N_42036);
and U43910 (N_43910,N_42263,N_42637);
nor U43911 (N_43911,N_42389,N_42252);
or U43912 (N_43912,N_42709,N_42804);
and U43913 (N_43913,N_42262,N_42585);
and U43914 (N_43914,N_42567,N_42511);
xnor U43915 (N_43915,N_42310,N_42136);
and U43916 (N_43916,N_42239,N_42624);
or U43917 (N_43917,N_42213,N_42078);
or U43918 (N_43918,N_42177,N_42813);
nand U43919 (N_43919,N_42947,N_42866);
xor U43920 (N_43920,N_42491,N_42628);
and U43921 (N_43921,N_42923,N_42825);
nand U43922 (N_43922,N_42628,N_42547);
nor U43923 (N_43923,N_42260,N_42576);
or U43924 (N_43924,N_42861,N_42234);
xor U43925 (N_43925,N_42239,N_42916);
nor U43926 (N_43926,N_42344,N_42944);
or U43927 (N_43927,N_42668,N_42432);
nor U43928 (N_43928,N_42784,N_42584);
nand U43929 (N_43929,N_42954,N_42923);
and U43930 (N_43930,N_42605,N_42994);
nand U43931 (N_43931,N_42646,N_42559);
xor U43932 (N_43932,N_42907,N_42280);
nand U43933 (N_43933,N_42163,N_42225);
xnor U43934 (N_43934,N_42374,N_42430);
and U43935 (N_43935,N_42122,N_42303);
and U43936 (N_43936,N_42877,N_42498);
xnor U43937 (N_43937,N_42769,N_42969);
and U43938 (N_43938,N_42134,N_42408);
and U43939 (N_43939,N_42456,N_42045);
nand U43940 (N_43940,N_42141,N_42979);
and U43941 (N_43941,N_42064,N_42201);
or U43942 (N_43942,N_42342,N_42654);
xor U43943 (N_43943,N_42859,N_42239);
xnor U43944 (N_43944,N_42513,N_42433);
nand U43945 (N_43945,N_42538,N_42541);
nand U43946 (N_43946,N_42886,N_42149);
or U43947 (N_43947,N_42067,N_42738);
xnor U43948 (N_43948,N_42086,N_42681);
or U43949 (N_43949,N_42182,N_42468);
and U43950 (N_43950,N_42096,N_42833);
nor U43951 (N_43951,N_42145,N_42992);
xnor U43952 (N_43952,N_42454,N_42577);
xnor U43953 (N_43953,N_42367,N_42113);
nand U43954 (N_43954,N_42977,N_42997);
or U43955 (N_43955,N_42149,N_42254);
nor U43956 (N_43956,N_42031,N_42228);
or U43957 (N_43957,N_42045,N_42631);
xor U43958 (N_43958,N_42714,N_42793);
xor U43959 (N_43959,N_42103,N_42472);
and U43960 (N_43960,N_42847,N_42905);
nor U43961 (N_43961,N_42100,N_42963);
xor U43962 (N_43962,N_42512,N_42273);
nor U43963 (N_43963,N_42521,N_42634);
xor U43964 (N_43964,N_42821,N_42729);
nand U43965 (N_43965,N_42996,N_42478);
nand U43966 (N_43966,N_42049,N_42513);
and U43967 (N_43967,N_42733,N_42439);
and U43968 (N_43968,N_42377,N_42900);
or U43969 (N_43969,N_42239,N_42592);
nand U43970 (N_43970,N_42632,N_42768);
nor U43971 (N_43971,N_42880,N_42442);
or U43972 (N_43972,N_42348,N_42186);
or U43973 (N_43973,N_42142,N_42019);
nor U43974 (N_43974,N_42037,N_42958);
xor U43975 (N_43975,N_42668,N_42470);
or U43976 (N_43976,N_42214,N_42131);
nor U43977 (N_43977,N_42578,N_42707);
and U43978 (N_43978,N_42666,N_42681);
nand U43979 (N_43979,N_42043,N_42132);
and U43980 (N_43980,N_42803,N_42756);
nand U43981 (N_43981,N_42823,N_42507);
and U43982 (N_43982,N_42609,N_42082);
nand U43983 (N_43983,N_42807,N_42046);
nand U43984 (N_43984,N_42084,N_42777);
xor U43985 (N_43985,N_42956,N_42312);
nor U43986 (N_43986,N_42781,N_42156);
and U43987 (N_43987,N_42592,N_42490);
or U43988 (N_43988,N_42738,N_42570);
nand U43989 (N_43989,N_42297,N_42134);
and U43990 (N_43990,N_42509,N_42739);
and U43991 (N_43991,N_42875,N_42504);
and U43992 (N_43992,N_42417,N_42538);
and U43993 (N_43993,N_42000,N_42151);
and U43994 (N_43994,N_42210,N_42000);
or U43995 (N_43995,N_42815,N_42195);
or U43996 (N_43996,N_42454,N_42397);
and U43997 (N_43997,N_42116,N_42502);
and U43998 (N_43998,N_42465,N_42600);
or U43999 (N_43999,N_42092,N_42356);
or U44000 (N_44000,N_43817,N_43628);
nand U44001 (N_44001,N_43756,N_43582);
or U44002 (N_44002,N_43503,N_43463);
nor U44003 (N_44003,N_43173,N_43118);
and U44004 (N_44004,N_43231,N_43102);
nor U44005 (N_44005,N_43474,N_43732);
nand U44006 (N_44006,N_43432,N_43986);
nand U44007 (N_44007,N_43194,N_43998);
and U44008 (N_44008,N_43225,N_43674);
nand U44009 (N_44009,N_43764,N_43807);
nor U44010 (N_44010,N_43854,N_43548);
xor U44011 (N_44011,N_43252,N_43535);
and U44012 (N_44012,N_43838,N_43268);
nand U44013 (N_44013,N_43845,N_43660);
xnor U44014 (N_44014,N_43920,N_43909);
xnor U44015 (N_44015,N_43755,N_43819);
xnor U44016 (N_44016,N_43300,N_43523);
and U44017 (N_44017,N_43192,N_43399);
or U44018 (N_44018,N_43462,N_43919);
xor U44019 (N_44019,N_43643,N_43861);
nor U44020 (N_44020,N_43293,N_43078);
and U44021 (N_44021,N_43196,N_43486);
or U44022 (N_44022,N_43084,N_43559);
nand U44023 (N_44023,N_43789,N_43925);
and U44024 (N_44024,N_43355,N_43809);
and U44025 (N_44025,N_43771,N_43276);
and U44026 (N_44026,N_43536,N_43524);
xor U44027 (N_44027,N_43450,N_43792);
nor U44028 (N_44028,N_43151,N_43226);
xor U44029 (N_44029,N_43250,N_43240);
nand U44030 (N_44030,N_43859,N_43769);
xor U44031 (N_44031,N_43784,N_43798);
xor U44032 (N_44032,N_43496,N_43826);
nor U44033 (N_44033,N_43454,N_43765);
nor U44034 (N_44034,N_43867,N_43741);
nor U44035 (N_44035,N_43583,N_43483);
nand U44036 (N_44036,N_43824,N_43951);
and U44037 (N_44037,N_43692,N_43640);
or U44038 (N_44038,N_43887,N_43725);
xor U44039 (N_44039,N_43487,N_43239);
xor U44040 (N_44040,N_43747,N_43544);
xnor U44041 (N_44041,N_43199,N_43728);
and U44042 (N_44042,N_43855,N_43629);
xnor U44043 (N_44043,N_43195,N_43733);
and U44044 (N_44044,N_43338,N_43851);
nand U44045 (N_44045,N_43967,N_43106);
xor U44046 (N_44046,N_43073,N_43219);
and U44047 (N_44047,N_43651,N_43934);
or U44048 (N_44048,N_43618,N_43184);
and U44049 (N_44049,N_43892,N_43721);
nor U44050 (N_44050,N_43472,N_43395);
or U44051 (N_44051,N_43011,N_43475);
nor U44052 (N_44052,N_43269,N_43017);
xnor U44053 (N_44053,N_43349,N_43460);
and U44054 (N_44054,N_43437,N_43259);
nand U44055 (N_44055,N_43963,N_43596);
and U44056 (N_44056,N_43014,N_43329);
nor U44057 (N_44057,N_43976,N_43871);
nand U44058 (N_44058,N_43661,N_43669);
nand U44059 (N_44059,N_43632,N_43930);
and U44060 (N_44060,N_43666,N_43558);
xnor U44061 (N_44061,N_43221,N_43551);
or U44062 (N_44062,N_43823,N_43623);
or U44063 (N_44063,N_43987,N_43303);
and U44064 (N_44064,N_43012,N_43519);
or U44065 (N_44065,N_43145,N_43082);
or U44066 (N_44066,N_43389,N_43274);
nor U44067 (N_44067,N_43726,N_43822);
and U44068 (N_44068,N_43198,N_43080);
nor U44069 (N_44069,N_43490,N_43754);
nand U44070 (N_44070,N_43790,N_43163);
nand U44071 (N_44071,N_43370,N_43321);
and U44072 (N_44072,N_43970,N_43580);
nor U44073 (N_44073,N_43023,N_43204);
or U44074 (N_44074,N_43206,N_43129);
or U44075 (N_44075,N_43641,N_43698);
xnor U44076 (N_44076,N_43626,N_43077);
and U44077 (N_44077,N_43600,N_43279);
and U44078 (N_44078,N_43015,N_43943);
xor U44079 (N_44079,N_43254,N_43757);
or U44080 (N_44080,N_43786,N_43974);
or U44081 (N_44081,N_43683,N_43103);
xor U44082 (N_44082,N_43470,N_43616);
and U44083 (N_44083,N_43801,N_43458);
and U44084 (N_44084,N_43227,N_43128);
xor U44085 (N_44085,N_43713,N_43575);
xnor U44086 (N_44086,N_43703,N_43690);
nand U44087 (N_44087,N_43135,N_43176);
nor U44088 (N_44088,N_43915,N_43372);
nand U44089 (N_44089,N_43762,N_43979);
nor U44090 (N_44090,N_43004,N_43562);
or U44091 (N_44091,N_43079,N_43260);
nor U44092 (N_44092,N_43440,N_43895);
nor U44093 (N_44093,N_43820,N_43639);
nand U44094 (N_44094,N_43933,N_43401);
and U44095 (N_44095,N_43479,N_43506);
and U44096 (N_44096,N_43697,N_43526);
xnor U44097 (N_44097,N_43185,N_43694);
xor U44098 (N_44098,N_43180,N_43876);
or U44099 (N_44099,N_43299,N_43730);
nor U44100 (N_44100,N_43803,N_43492);
nor U44101 (N_44101,N_43289,N_43325);
and U44102 (N_44102,N_43530,N_43656);
nand U44103 (N_44103,N_43423,N_43534);
or U44104 (N_44104,N_43120,N_43283);
nand U44105 (N_44105,N_43386,N_43687);
nor U44106 (N_44106,N_43108,N_43055);
and U44107 (N_44107,N_43316,N_43527);
or U44108 (N_44108,N_43944,N_43946);
xor U44109 (N_44109,N_43997,N_43680);
or U44110 (N_44110,N_43150,N_43636);
nand U44111 (N_44111,N_43610,N_43126);
or U44112 (N_44112,N_43183,N_43200);
nor U44113 (N_44113,N_43652,N_43353);
or U44114 (N_44114,N_43650,N_43388);
or U44115 (N_44115,N_43996,N_43298);
and U44116 (N_44116,N_43043,N_43744);
nand U44117 (N_44117,N_43465,N_43121);
nor U44118 (N_44118,N_43203,N_43913);
xor U44119 (N_44119,N_43222,N_43659);
and U44120 (N_44120,N_43917,N_43517);
xor U44121 (N_44121,N_43761,N_43988);
and U44122 (N_44122,N_43242,N_43480);
nor U44123 (N_44123,N_43696,N_43210);
nor U44124 (N_44124,N_43856,N_43760);
xor U44125 (N_44125,N_43770,N_43785);
xnor U44126 (N_44126,N_43029,N_43606);
xnor U44127 (N_44127,N_43123,N_43658);
and U44128 (N_44128,N_43094,N_43104);
and U44129 (N_44129,N_43396,N_43352);
nor U44130 (N_44130,N_43264,N_43599);
nor U44131 (N_44131,N_43904,N_43686);
nand U44132 (N_44132,N_43648,N_43540);
nor U44133 (N_44133,N_43751,N_43516);
nand U44134 (N_44134,N_43350,N_43339);
or U44135 (N_44135,N_43369,N_43074);
nor U44136 (N_44136,N_43868,N_43209);
nand U44137 (N_44137,N_43403,N_43211);
xnor U44138 (N_44138,N_43049,N_43985);
and U44139 (N_44139,N_43024,N_43097);
nor U44140 (N_44140,N_43810,N_43064);
nor U44141 (N_44141,N_43238,N_43175);
nand U44142 (N_44142,N_43363,N_43502);
xor U44143 (N_44143,N_43685,N_43670);
nor U44144 (N_44144,N_43020,N_43453);
nand U44145 (N_44145,N_43679,N_43869);
and U44146 (N_44146,N_43076,N_43570);
or U44147 (N_44147,N_43164,N_43107);
nor U44148 (N_44148,N_43335,N_43627);
nand U44149 (N_44149,N_43815,N_43287);
nor U44150 (N_44150,N_43019,N_43662);
nand U44151 (N_44151,N_43565,N_43039);
or U44152 (N_44152,N_43032,N_43262);
nor U44153 (N_44153,N_43099,N_43310);
nor U44154 (N_44154,N_43553,N_43301);
and U44155 (N_44155,N_43707,N_43667);
nand U44156 (N_44156,N_43360,N_43655);
or U44157 (N_44157,N_43441,N_43290);
and U44158 (N_44158,N_43953,N_43980);
or U44159 (N_44159,N_43307,N_43962);
nand U44160 (N_44160,N_43091,N_43808);
and U44161 (N_44161,N_43843,N_43605);
nand U44162 (N_44162,N_43588,N_43607);
or U44163 (N_44163,N_43532,N_43417);
nor U44164 (N_44164,N_43139,N_43497);
nor U44165 (N_44165,N_43695,N_43291);
xor U44166 (N_44166,N_43846,N_43675);
nor U44167 (N_44167,N_43407,N_43724);
or U44168 (N_44168,N_43812,N_43383);
or U44169 (N_44169,N_43796,N_43347);
xnor U44170 (N_44170,N_43921,N_43545);
xor U44171 (N_44171,N_43603,N_43883);
xor U44172 (N_44172,N_43438,N_43853);
and U44173 (N_44173,N_43923,N_43657);
nor U44174 (N_44174,N_43275,N_43215);
or U44175 (N_44175,N_43218,N_43070);
xor U44176 (N_44176,N_43277,N_43935);
nor U44177 (N_44177,N_43469,N_43366);
and U44178 (N_44178,N_43172,N_43763);
nand U44179 (N_44179,N_43237,N_43499);
or U44180 (N_44180,N_43059,N_43518);
xnor U44181 (N_44181,N_43612,N_43729);
and U44182 (N_44182,N_43167,N_43112);
or U44183 (N_44183,N_43689,N_43897);
or U44184 (N_44184,N_43447,N_43054);
or U44185 (N_44185,N_43704,N_43343);
xnor U44186 (N_44186,N_43966,N_43473);
or U44187 (N_44187,N_43870,N_43842);
xnor U44188 (N_44188,N_43874,N_43813);
nand U44189 (N_44189,N_43711,N_43031);
nand U44190 (N_44190,N_43642,N_43543);
and U44191 (N_44191,N_43320,N_43088);
xor U44192 (N_44192,N_43302,N_43331);
or U44193 (N_44193,N_43863,N_43739);
nor U44194 (N_44194,N_43385,N_43306);
or U44195 (N_44195,N_43886,N_43394);
nor U44196 (N_44196,N_43356,N_43836);
and U44197 (N_44197,N_43515,N_43026);
and U44198 (N_44198,N_43865,N_43914);
xnor U44199 (N_44199,N_43504,N_43900);
xnor U44200 (N_44200,N_43554,N_43811);
nor U44201 (N_44201,N_43945,N_43214);
and U44202 (N_44202,N_43577,N_43926);
xnor U44203 (N_44203,N_43034,N_43560);
xnor U44204 (N_44204,N_43124,N_43875);
and U44205 (N_44205,N_43574,N_43405);
or U44206 (N_44206,N_43902,N_43891);
nand U44207 (N_44207,N_43702,N_43783);
nor U44208 (N_44208,N_43528,N_43062);
nand U44209 (N_44209,N_43825,N_43731);
or U44210 (N_44210,N_43994,N_43390);
and U44211 (N_44211,N_43529,N_43485);
nand U44212 (N_44212,N_43681,N_43244);
and U44213 (N_44213,N_43533,N_43512);
nand U44214 (N_44214,N_43371,N_43814);
or U44215 (N_44215,N_43734,N_43456);
nor U44216 (N_44216,N_43481,N_43578);
nor U44217 (N_44217,N_43255,N_43758);
xnor U44218 (N_44218,N_43896,N_43952);
nand U44219 (N_44219,N_43188,N_43443);
nand U44220 (N_44220,N_43426,N_43162);
xnor U44221 (N_44221,N_43625,N_43873);
nand U44222 (N_44222,N_43999,N_43592);
xor U44223 (N_44223,N_43452,N_43593);
nand U44224 (N_44224,N_43514,N_43380);
xor U44225 (N_44225,N_43931,N_43066);
xnor U44226 (N_44226,N_43271,N_43100);
nand U44227 (N_44227,N_43878,N_43067);
and U44228 (N_44228,N_43359,N_43482);
and U44229 (N_44229,N_43672,N_43978);
xor U44230 (N_44230,N_43157,N_43522);
and U44231 (N_44231,N_43959,N_43631);
nand U44232 (N_44232,N_43468,N_43950);
and U44233 (N_44233,N_43833,N_43849);
nand U44234 (N_44234,N_43791,N_43367);
nor U44235 (N_44235,N_43484,N_43940);
or U44236 (N_44236,N_43585,N_43701);
xor U44237 (N_44237,N_43954,N_43649);
and U44238 (N_44238,N_43323,N_43511);
and U44239 (N_44239,N_43056,N_43042);
nand U44240 (N_44240,N_43982,N_43147);
nand U44241 (N_44241,N_43364,N_43332);
xor U44242 (N_44242,N_43142,N_43948);
nor U44243 (N_44243,N_43712,N_43907);
or U44244 (N_44244,N_43361,N_43408);
or U44245 (N_44245,N_43146,N_43615);
and U44246 (N_44246,N_43916,N_43956);
nand U44247 (N_44247,N_43132,N_43095);
nor U44248 (N_44248,N_43774,N_43805);
or U44249 (N_44249,N_43041,N_43451);
nand U44250 (N_44250,N_43313,N_43673);
and U44251 (N_44251,N_43889,N_43190);
and U44252 (N_44252,N_43633,N_43096);
nand U44253 (N_44253,N_43884,N_43280);
or U44254 (N_44254,N_43937,N_43348);
nand U44255 (N_44255,N_43936,N_43620);
or U44256 (N_44256,N_43068,N_43572);
or U44257 (N_44257,N_43576,N_43416);
and U44258 (N_44258,N_43341,N_43051);
nor U44259 (N_44259,N_43797,N_43158);
and U44260 (N_44260,N_43182,N_43243);
nand U44261 (N_44261,N_43375,N_43717);
nand U44262 (N_44262,N_43333,N_43893);
and U44263 (N_44263,N_43412,N_43414);
and U44264 (N_44264,N_43839,N_43425);
nor U44265 (N_44265,N_43973,N_43075);
nand U44266 (N_44266,N_43688,N_43109);
xnor U44267 (N_44267,N_43767,N_43903);
nand U44268 (N_44268,N_43415,N_43033);
xnor U44269 (N_44269,N_43140,N_43156);
nor U44270 (N_44270,N_43705,N_43847);
or U44271 (N_44271,N_43579,N_43406);
nor U44272 (N_44272,N_43130,N_43776);
xnor U44273 (N_44273,N_43028,N_43787);
and U44274 (N_44274,N_43477,N_43816);
nand U44275 (N_44275,N_43714,N_43086);
nand U44276 (N_44276,N_43205,N_43581);
xnor U44277 (N_44277,N_43598,N_43802);
nor U44278 (N_44278,N_43500,N_43773);
nor U44279 (N_44279,N_43566,N_43089);
xnor U44280 (N_44280,N_43236,N_43977);
or U44281 (N_44281,N_43362,N_43471);
nor U44282 (N_44282,N_43358,N_43898);
and U44283 (N_44283,N_43430,N_43961);
xor U44284 (N_44284,N_43317,N_43327);
nand U44285 (N_44285,N_43782,N_43573);
nor U44286 (N_44286,N_43495,N_43928);
or U44287 (N_44287,N_43737,N_43233);
nand U44288 (N_44288,N_43968,N_43932);
nor U44289 (N_44289,N_43949,N_43110);
nand U44290 (N_44290,N_43664,N_43964);
nand U44291 (N_44291,N_43382,N_43398);
xnor U44292 (N_44292,N_43265,N_43491);
nand U44293 (N_44293,N_43131,N_43409);
xnor U44294 (N_44294,N_43324,N_43419);
nor U44295 (N_44295,N_43908,N_43745);
or U44296 (N_44296,N_43924,N_43044);
and U44297 (N_44297,N_43992,N_43821);
nand U44298 (N_44298,N_43965,N_43174);
nor U44299 (N_44299,N_43159,N_43594);
nor U44300 (N_44300,N_43906,N_43245);
nor U44301 (N_44301,N_43336,N_43637);
xor U44302 (N_44302,N_43834,N_43251);
xnor U44303 (N_44303,N_43141,N_43911);
and U44304 (N_44304,N_43852,N_43759);
or U44305 (N_44305,N_43002,N_43220);
or U44306 (N_44306,N_43677,N_43624);
nor U44307 (N_44307,N_43645,N_43030);
nand U44308 (N_44308,N_43166,N_43983);
or U44309 (N_44309,N_43840,N_43866);
and U44310 (N_44310,N_43045,N_43181);
xnor U44311 (N_44311,N_43050,N_43421);
or U44312 (N_44312,N_43716,N_43161);
xor U44313 (N_44313,N_43153,N_43314);
xor U44314 (N_44314,N_43571,N_43635);
nand U44315 (N_44315,N_43105,N_43736);
and U44316 (N_44316,N_43488,N_43601);
nor U44317 (N_44317,N_43160,N_43521);
nand U44318 (N_44318,N_43989,N_43595);
or U44319 (N_44319,N_43531,N_43609);
xor U44320 (N_44320,N_43549,N_43114);
nor U44321 (N_44321,N_43614,N_43171);
xor U44322 (N_44322,N_43248,N_43547);
xnor U44323 (N_44323,N_43111,N_43378);
nand U44324 (N_44324,N_43273,N_43296);
nor U44325 (N_44325,N_43006,N_43848);
xor U44326 (N_44326,N_43288,N_43189);
nand U44327 (N_44327,N_43253,N_43351);
nand U44328 (N_44328,N_43742,N_43178);
xor U44329 (N_44329,N_43376,N_43308);
or U44330 (N_44330,N_43021,N_43975);
nor U44331 (N_44331,N_43493,N_43455);
nand U44332 (N_44332,N_43442,N_43431);
or U44333 (N_44333,N_43284,N_43727);
nand U44334 (N_44334,N_43127,N_43563);
nand U44335 (N_44335,N_43459,N_43234);
nor U44336 (N_44336,N_43835,N_43918);
xor U44337 (N_44337,N_43768,N_43263);
and U44338 (N_44338,N_43971,N_43735);
nand U44339 (N_44339,N_43427,N_43040);
nor U44340 (N_44340,N_43410,N_43402);
nand U44341 (N_44341,N_43613,N_43235);
and U44342 (N_44342,N_43827,N_43001);
nand U44343 (N_44343,N_43539,N_43960);
and U44344 (N_44344,N_43311,N_43546);
nor U44345 (N_44345,N_43144,N_43116);
and U44346 (N_44346,N_43397,N_43795);
nor U44347 (N_44347,N_43027,N_43719);
nand U44348 (N_44348,N_43723,N_43653);
nand U44349 (N_44349,N_43586,N_43009);
and U44350 (N_44350,N_43990,N_43213);
nor U44351 (N_44351,N_43993,N_43429);
xor U44352 (N_44352,N_43346,N_43047);
nand U44353 (N_44353,N_43207,N_43750);
or U44354 (N_44354,N_43899,N_43556);
nor U44355 (N_44355,N_43972,N_43799);
nand U44356 (N_44356,N_43864,N_43446);
nand U44357 (N_44357,N_43788,N_43910);
and U44358 (N_44358,N_43374,N_43115);
and U44359 (N_44359,N_43046,N_43831);
xor U44360 (N_44360,N_43510,N_43537);
and U44361 (N_44361,N_43258,N_43439);
and U44362 (N_44362,N_43354,N_43525);
and U44363 (N_44363,N_43319,N_43434);
nor U44364 (N_44364,N_43958,N_43381);
or U44365 (N_44365,N_43148,N_43400);
nor U44366 (N_44366,N_43743,N_43008);
and U44367 (N_44367,N_43092,N_43927);
xor U44368 (N_44368,N_43619,N_43186);
nor U44369 (N_44369,N_43589,N_43038);
nand U44370 (N_44370,N_43671,N_43602);
nand U44371 (N_44371,N_43684,N_43800);
and U44372 (N_44372,N_43804,N_43230);
and U44373 (N_44373,N_43093,N_43016);
or U44374 (N_44374,N_43830,N_43445);
nor U44375 (N_44375,N_43393,N_43201);
xor U44376 (N_44376,N_43229,N_43035);
xnor U44377 (N_44377,N_43505,N_43337);
and U44378 (N_44378,N_43885,N_43538);
xor U44379 (N_44379,N_43053,N_43941);
nor U44380 (N_44380,N_43257,N_43777);
nor U44381 (N_44381,N_43706,N_43413);
nand U44382 (N_44382,N_43860,N_43748);
nand U44383 (N_44383,N_43654,N_43793);
or U44384 (N_44384,N_43622,N_43753);
nand U44385 (N_44385,N_43202,N_43567);
nand U44386 (N_44386,N_43330,N_43678);
xor U44387 (N_44387,N_43718,N_43326);
nor U44388 (N_44388,N_43342,N_43090);
or U44389 (N_44389,N_43844,N_43555);
or U44390 (N_44390,N_43905,N_43422);
and U44391 (N_44391,N_43850,N_43297);
nor U44392 (N_44392,N_43191,N_43249);
or U44393 (N_44393,N_43942,N_43520);
nand U44394 (N_44394,N_43464,N_43604);
and U44395 (N_44395,N_43278,N_43022);
nand U44396 (N_44396,N_43818,N_43740);
xor U44397 (N_44397,N_43995,N_43435);
nor U44398 (N_44398,N_43057,N_43591);
xnor U44399 (N_44399,N_43781,N_43929);
nor U44400 (N_44400,N_43246,N_43010);
nand U44401 (N_44401,N_43507,N_43541);
or U44402 (N_44402,N_43466,N_43224);
and U44403 (N_44403,N_43444,N_43749);
nand U44404 (N_44404,N_43113,N_43890);
nor U44405 (N_44405,N_43862,N_43122);
nand U44406 (N_44406,N_43478,N_43557);
xor U44407 (N_44407,N_43428,N_43018);
nor U44408 (N_44408,N_43305,N_43119);
or U44409 (N_44409,N_43715,N_43508);
and U44410 (N_44410,N_43779,N_43552);
and U44411 (N_44411,N_43286,N_43368);
nand U44412 (N_44412,N_43901,N_43304);
nand U44413 (N_44413,N_43256,N_43069);
and U44414 (N_44414,N_43154,N_43025);
or U44415 (N_44415,N_43832,N_43433);
and U44416 (N_44416,N_43969,N_43003);
or U44417 (N_44417,N_43879,N_43668);
and U44418 (N_44418,N_43647,N_43138);
nor U44419 (N_44419,N_43778,N_43134);
nand U44420 (N_44420,N_43170,N_43387);
or U44421 (N_44421,N_43420,N_43117);
or U44422 (N_44422,N_43912,N_43880);
and U44423 (N_44423,N_43569,N_43261);
and U44424 (N_44424,N_43266,N_43328);
and U44425 (N_44425,N_43072,N_43665);
and U44426 (N_44426,N_43197,N_43568);
nor U44427 (N_44427,N_43208,N_43133);
or U44428 (N_44428,N_43125,N_43584);
nor U44429 (N_44429,N_43065,N_43165);
xnor U44430 (N_44430,N_43212,N_43424);
or U44431 (N_44431,N_43663,N_43738);
or U44432 (N_44432,N_43476,N_43775);
xor U44433 (N_44433,N_43007,N_43691);
or U44434 (N_44434,N_43693,N_43318);
xor U44435 (N_44435,N_43611,N_43149);
nor U44436 (N_44436,N_43947,N_43981);
and U44437 (N_44437,N_43646,N_43177);
or U44438 (N_44438,N_43391,N_43489);
or U44439 (N_44439,N_43058,N_43780);
and U44440 (N_44440,N_43766,N_43841);
nor U44441 (N_44441,N_43060,N_43882);
nand U44442 (N_44442,N_43621,N_43193);
nor U44443 (N_44443,N_43136,N_43340);
nor U44444 (N_44444,N_43270,N_43071);
and U44445 (N_44445,N_43063,N_43168);
nor U44446 (N_44446,N_43561,N_43098);
nand U44447 (N_44447,N_43377,N_43772);
xor U44448 (N_44448,N_43984,N_43564);
nor U44449 (N_44449,N_43322,N_43411);
nand U44450 (N_44450,N_43232,N_43137);
and U44451 (N_44451,N_43888,N_43597);
xor U44452 (N_44452,N_43081,N_43282);
nor U44453 (N_44453,N_43991,N_43083);
xor U44454 (N_44454,N_43700,N_43436);
nor U44455 (N_44455,N_43644,N_43682);
xnor U44456 (N_44456,N_43267,N_43179);
xnor U44457 (N_44457,N_43052,N_43000);
nand U44458 (N_44458,N_43143,N_43404);
or U44459 (N_44459,N_43344,N_43013);
nor U44460 (N_44460,N_43676,N_43085);
or U44461 (N_44461,N_43216,N_43228);
and U44462 (N_44462,N_43638,N_43457);
xnor U44463 (N_44463,N_43630,N_43285);
nand U44464 (N_44464,N_43881,N_43872);
nor U44465 (N_44465,N_43315,N_43939);
xor U44466 (N_44466,N_43461,N_43379);
or U44467 (N_44467,N_43384,N_43509);
or U44468 (N_44468,N_43708,N_43152);
nor U44469 (N_44469,N_43247,N_43837);
xor U44470 (N_44470,N_43722,N_43036);
xor U44471 (N_44471,N_43217,N_43806);
and U44472 (N_44472,N_43501,N_43922);
and U44473 (N_44473,N_43357,N_43345);
nor U44474 (N_44474,N_43542,N_43187);
and U44475 (N_44475,N_43857,N_43746);
nor U44476 (N_44476,N_43294,N_43365);
nand U44477 (N_44477,N_43037,N_43449);
nor U44478 (N_44478,N_43169,N_43550);
nand U44479 (N_44479,N_43048,N_43295);
xnor U44480 (N_44480,N_43957,N_43223);
or U44481 (N_44481,N_43877,N_43710);
and U44482 (N_44482,N_43467,N_43955);
and U44483 (N_44483,N_43709,N_43061);
nor U44484 (N_44484,N_43281,N_43894);
nor U44485 (N_44485,N_43513,N_43587);
nand U44486 (N_44486,N_43608,N_43829);
xor U44487 (N_44487,N_43155,N_43272);
or U44488 (N_44488,N_43392,N_43418);
nand U44489 (N_44489,N_43938,N_43241);
nor U44490 (N_44490,N_43494,N_43309);
and U44491 (N_44491,N_43720,N_43794);
or U44492 (N_44492,N_43373,N_43312);
or U44493 (N_44493,N_43334,N_43448);
and U44494 (N_44494,N_43699,N_43858);
or U44495 (N_44495,N_43828,N_43292);
xnor U44496 (N_44496,N_43498,N_43087);
and U44497 (N_44497,N_43634,N_43617);
and U44498 (N_44498,N_43590,N_43101);
and U44499 (N_44499,N_43005,N_43752);
nand U44500 (N_44500,N_43219,N_43935);
or U44501 (N_44501,N_43494,N_43658);
or U44502 (N_44502,N_43276,N_43127);
and U44503 (N_44503,N_43758,N_43325);
or U44504 (N_44504,N_43021,N_43962);
xor U44505 (N_44505,N_43901,N_43616);
and U44506 (N_44506,N_43380,N_43502);
or U44507 (N_44507,N_43368,N_43028);
nor U44508 (N_44508,N_43367,N_43729);
and U44509 (N_44509,N_43863,N_43653);
xnor U44510 (N_44510,N_43068,N_43490);
nor U44511 (N_44511,N_43409,N_43977);
nor U44512 (N_44512,N_43155,N_43650);
or U44513 (N_44513,N_43660,N_43217);
and U44514 (N_44514,N_43823,N_43618);
xnor U44515 (N_44515,N_43216,N_43760);
xnor U44516 (N_44516,N_43130,N_43089);
xor U44517 (N_44517,N_43014,N_43952);
or U44518 (N_44518,N_43200,N_43839);
nand U44519 (N_44519,N_43460,N_43612);
nor U44520 (N_44520,N_43140,N_43958);
and U44521 (N_44521,N_43191,N_43748);
xor U44522 (N_44522,N_43780,N_43556);
and U44523 (N_44523,N_43423,N_43283);
nand U44524 (N_44524,N_43031,N_43585);
nand U44525 (N_44525,N_43941,N_43023);
xnor U44526 (N_44526,N_43617,N_43915);
nand U44527 (N_44527,N_43358,N_43873);
or U44528 (N_44528,N_43136,N_43987);
nand U44529 (N_44529,N_43279,N_43112);
nand U44530 (N_44530,N_43657,N_43424);
xor U44531 (N_44531,N_43679,N_43443);
or U44532 (N_44532,N_43949,N_43948);
nand U44533 (N_44533,N_43457,N_43509);
nand U44534 (N_44534,N_43599,N_43987);
or U44535 (N_44535,N_43525,N_43246);
nand U44536 (N_44536,N_43758,N_43063);
or U44537 (N_44537,N_43528,N_43845);
or U44538 (N_44538,N_43101,N_43695);
and U44539 (N_44539,N_43369,N_43308);
nand U44540 (N_44540,N_43614,N_43587);
nor U44541 (N_44541,N_43014,N_43008);
and U44542 (N_44542,N_43302,N_43231);
nand U44543 (N_44543,N_43126,N_43837);
or U44544 (N_44544,N_43862,N_43900);
xor U44545 (N_44545,N_43273,N_43942);
and U44546 (N_44546,N_43042,N_43364);
or U44547 (N_44547,N_43145,N_43347);
nor U44548 (N_44548,N_43264,N_43267);
and U44549 (N_44549,N_43398,N_43469);
nand U44550 (N_44550,N_43522,N_43774);
nor U44551 (N_44551,N_43516,N_43062);
nor U44552 (N_44552,N_43484,N_43878);
nor U44553 (N_44553,N_43038,N_43487);
or U44554 (N_44554,N_43197,N_43790);
and U44555 (N_44555,N_43627,N_43412);
xnor U44556 (N_44556,N_43773,N_43150);
xor U44557 (N_44557,N_43363,N_43412);
or U44558 (N_44558,N_43031,N_43668);
nor U44559 (N_44559,N_43565,N_43462);
or U44560 (N_44560,N_43798,N_43664);
or U44561 (N_44561,N_43091,N_43322);
xnor U44562 (N_44562,N_43108,N_43653);
and U44563 (N_44563,N_43857,N_43328);
and U44564 (N_44564,N_43487,N_43449);
and U44565 (N_44565,N_43939,N_43621);
xnor U44566 (N_44566,N_43877,N_43329);
or U44567 (N_44567,N_43574,N_43637);
and U44568 (N_44568,N_43939,N_43463);
and U44569 (N_44569,N_43055,N_43670);
xnor U44570 (N_44570,N_43079,N_43304);
and U44571 (N_44571,N_43667,N_43858);
nor U44572 (N_44572,N_43898,N_43608);
or U44573 (N_44573,N_43881,N_43825);
nor U44574 (N_44574,N_43006,N_43741);
and U44575 (N_44575,N_43622,N_43538);
nor U44576 (N_44576,N_43032,N_43810);
nand U44577 (N_44577,N_43974,N_43971);
nor U44578 (N_44578,N_43264,N_43309);
xor U44579 (N_44579,N_43335,N_43480);
nor U44580 (N_44580,N_43523,N_43110);
nand U44581 (N_44581,N_43290,N_43821);
or U44582 (N_44582,N_43917,N_43174);
or U44583 (N_44583,N_43629,N_43464);
or U44584 (N_44584,N_43457,N_43325);
nand U44585 (N_44585,N_43829,N_43069);
and U44586 (N_44586,N_43196,N_43646);
or U44587 (N_44587,N_43878,N_43256);
nor U44588 (N_44588,N_43868,N_43433);
xor U44589 (N_44589,N_43463,N_43663);
and U44590 (N_44590,N_43179,N_43693);
nor U44591 (N_44591,N_43866,N_43821);
nand U44592 (N_44592,N_43523,N_43989);
nor U44593 (N_44593,N_43726,N_43324);
xor U44594 (N_44594,N_43721,N_43411);
nor U44595 (N_44595,N_43576,N_43488);
or U44596 (N_44596,N_43649,N_43849);
nor U44597 (N_44597,N_43393,N_43028);
nand U44598 (N_44598,N_43681,N_43670);
and U44599 (N_44599,N_43660,N_43901);
nand U44600 (N_44600,N_43509,N_43685);
and U44601 (N_44601,N_43068,N_43047);
or U44602 (N_44602,N_43075,N_43024);
and U44603 (N_44603,N_43045,N_43768);
nand U44604 (N_44604,N_43589,N_43782);
xor U44605 (N_44605,N_43244,N_43597);
or U44606 (N_44606,N_43345,N_43966);
nand U44607 (N_44607,N_43230,N_43512);
nor U44608 (N_44608,N_43727,N_43118);
and U44609 (N_44609,N_43152,N_43157);
nor U44610 (N_44610,N_43597,N_43031);
or U44611 (N_44611,N_43841,N_43973);
or U44612 (N_44612,N_43947,N_43613);
xor U44613 (N_44613,N_43297,N_43545);
nor U44614 (N_44614,N_43933,N_43315);
and U44615 (N_44615,N_43822,N_43596);
or U44616 (N_44616,N_43144,N_43573);
or U44617 (N_44617,N_43658,N_43795);
or U44618 (N_44618,N_43896,N_43058);
and U44619 (N_44619,N_43182,N_43111);
and U44620 (N_44620,N_43747,N_43214);
nand U44621 (N_44621,N_43122,N_43050);
and U44622 (N_44622,N_43345,N_43923);
and U44623 (N_44623,N_43763,N_43179);
nor U44624 (N_44624,N_43286,N_43980);
nand U44625 (N_44625,N_43926,N_43675);
nor U44626 (N_44626,N_43623,N_43669);
or U44627 (N_44627,N_43546,N_43938);
nor U44628 (N_44628,N_43513,N_43498);
nand U44629 (N_44629,N_43538,N_43548);
nor U44630 (N_44630,N_43002,N_43285);
xnor U44631 (N_44631,N_43897,N_43253);
nor U44632 (N_44632,N_43539,N_43961);
nor U44633 (N_44633,N_43553,N_43935);
or U44634 (N_44634,N_43364,N_43367);
and U44635 (N_44635,N_43357,N_43153);
nor U44636 (N_44636,N_43441,N_43421);
nor U44637 (N_44637,N_43343,N_43490);
nor U44638 (N_44638,N_43066,N_43668);
or U44639 (N_44639,N_43826,N_43579);
xor U44640 (N_44640,N_43459,N_43398);
xor U44641 (N_44641,N_43874,N_43831);
nor U44642 (N_44642,N_43317,N_43098);
xnor U44643 (N_44643,N_43808,N_43888);
nor U44644 (N_44644,N_43923,N_43693);
or U44645 (N_44645,N_43714,N_43273);
and U44646 (N_44646,N_43901,N_43011);
xor U44647 (N_44647,N_43347,N_43242);
and U44648 (N_44648,N_43176,N_43056);
nor U44649 (N_44649,N_43763,N_43370);
and U44650 (N_44650,N_43887,N_43015);
nor U44651 (N_44651,N_43552,N_43969);
nor U44652 (N_44652,N_43263,N_43910);
xnor U44653 (N_44653,N_43915,N_43756);
or U44654 (N_44654,N_43931,N_43721);
xor U44655 (N_44655,N_43968,N_43116);
or U44656 (N_44656,N_43966,N_43230);
and U44657 (N_44657,N_43997,N_43377);
nand U44658 (N_44658,N_43552,N_43458);
nand U44659 (N_44659,N_43063,N_43402);
xor U44660 (N_44660,N_43906,N_43312);
nand U44661 (N_44661,N_43940,N_43080);
nand U44662 (N_44662,N_43131,N_43872);
xnor U44663 (N_44663,N_43563,N_43410);
nor U44664 (N_44664,N_43278,N_43624);
or U44665 (N_44665,N_43959,N_43968);
or U44666 (N_44666,N_43727,N_43014);
nor U44667 (N_44667,N_43428,N_43994);
or U44668 (N_44668,N_43469,N_43013);
xor U44669 (N_44669,N_43479,N_43470);
and U44670 (N_44670,N_43756,N_43696);
nor U44671 (N_44671,N_43583,N_43658);
xor U44672 (N_44672,N_43701,N_43034);
nor U44673 (N_44673,N_43445,N_43545);
nor U44674 (N_44674,N_43997,N_43165);
nand U44675 (N_44675,N_43295,N_43779);
nor U44676 (N_44676,N_43967,N_43893);
xnor U44677 (N_44677,N_43025,N_43939);
and U44678 (N_44678,N_43025,N_43089);
and U44679 (N_44679,N_43757,N_43833);
nand U44680 (N_44680,N_43422,N_43828);
nand U44681 (N_44681,N_43021,N_43610);
nand U44682 (N_44682,N_43857,N_43166);
xnor U44683 (N_44683,N_43303,N_43275);
nand U44684 (N_44684,N_43973,N_43693);
xor U44685 (N_44685,N_43160,N_43921);
xnor U44686 (N_44686,N_43214,N_43347);
nor U44687 (N_44687,N_43837,N_43622);
and U44688 (N_44688,N_43869,N_43983);
nor U44689 (N_44689,N_43072,N_43088);
nor U44690 (N_44690,N_43314,N_43028);
and U44691 (N_44691,N_43775,N_43561);
nor U44692 (N_44692,N_43471,N_43449);
nand U44693 (N_44693,N_43946,N_43182);
and U44694 (N_44694,N_43331,N_43567);
nand U44695 (N_44695,N_43737,N_43647);
and U44696 (N_44696,N_43907,N_43634);
and U44697 (N_44697,N_43881,N_43611);
xnor U44698 (N_44698,N_43452,N_43567);
nor U44699 (N_44699,N_43428,N_43640);
xor U44700 (N_44700,N_43204,N_43288);
or U44701 (N_44701,N_43461,N_43444);
and U44702 (N_44702,N_43310,N_43698);
nand U44703 (N_44703,N_43779,N_43643);
nor U44704 (N_44704,N_43074,N_43211);
nor U44705 (N_44705,N_43950,N_43512);
and U44706 (N_44706,N_43287,N_43198);
xor U44707 (N_44707,N_43444,N_43776);
nor U44708 (N_44708,N_43275,N_43891);
xor U44709 (N_44709,N_43455,N_43891);
xnor U44710 (N_44710,N_43079,N_43531);
and U44711 (N_44711,N_43222,N_43168);
nor U44712 (N_44712,N_43774,N_43371);
or U44713 (N_44713,N_43823,N_43630);
or U44714 (N_44714,N_43714,N_43765);
xnor U44715 (N_44715,N_43371,N_43305);
and U44716 (N_44716,N_43649,N_43301);
or U44717 (N_44717,N_43273,N_43640);
and U44718 (N_44718,N_43449,N_43439);
xnor U44719 (N_44719,N_43886,N_43148);
nand U44720 (N_44720,N_43567,N_43899);
nand U44721 (N_44721,N_43921,N_43961);
or U44722 (N_44722,N_43762,N_43336);
and U44723 (N_44723,N_43525,N_43212);
xor U44724 (N_44724,N_43553,N_43479);
or U44725 (N_44725,N_43421,N_43711);
or U44726 (N_44726,N_43590,N_43279);
xnor U44727 (N_44727,N_43255,N_43642);
nor U44728 (N_44728,N_43079,N_43792);
nor U44729 (N_44729,N_43230,N_43776);
and U44730 (N_44730,N_43450,N_43398);
nor U44731 (N_44731,N_43055,N_43489);
and U44732 (N_44732,N_43767,N_43501);
nand U44733 (N_44733,N_43844,N_43541);
nand U44734 (N_44734,N_43402,N_43126);
or U44735 (N_44735,N_43974,N_43142);
and U44736 (N_44736,N_43372,N_43433);
nor U44737 (N_44737,N_43015,N_43343);
nor U44738 (N_44738,N_43821,N_43525);
nand U44739 (N_44739,N_43436,N_43225);
xnor U44740 (N_44740,N_43141,N_43151);
and U44741 (N_44741,N_43445,N_43538);
nand U44742 (N_44742,N_43368,N_43920);
and U44743 (N_44743,N_43716,N_43489);
xnor U44744 (N_44744,N_43036,N_43091);
nand U44745 (N_44745,N_43326,N_43957);
nor U44746 (N_44746,N_43886,N_43345);
nand U44747 (N_44747,N_43679,N_43090);
and U44748 (N_44748,N_43411,N_43403);
nand U44749 (N_44749,N_43102,N_43190);
nand U44750 (N_44750,N_43001,N_43794);
or U44751 (N_44751,N_43937,N_43389);
or U44752 (N_44752,N_43610,N_43102);
nand U44753 (N_44753,N_43209,N_43610);
xnor U44754 (N_44754,N_43665,N_43463);
xnor U44755 (N_44755,N_43928,N_43153);
xnor U44756 (N_44756,N_43970,N_43246);
xor U44757 (N_44757,N_43843,N_43924);
and U44758 (N_44758,N_43947,N_43009);
or U44759 (N_44759,N_43186,N_43311);
nor U44760 (N_44760,N_43932,N_43391);
xnor U44761 (N_44761,N_43028,N_43783);
nor U44762 (N_44762,N_43374,N_43075);
xor U44763 (N_44763,N_43315,N_43439);
nand U44764 (N_44764,N_43956,N_43505);
nand U44765 (N_44765,N_43517,N_43833);
and U44766 (N_44766,N_43877,N_43713);
nor U44767 (N_44767,N_43072,N_43851);
nor U44768 (N_44768,N_43008,N_43272);
or U44769 (N_44769,N_43441,N_43965);
nor U44770 (N_44770,N_43734,N_43860);
xor U44771 (N_44771,N_43401,N_43617);
xor U44772 (N_44772,N_43923,N_43145);
nand U44773 (N_44773,N_43431,N_43099);
nor U44774 (N_44774,N_43912,N_43824);
nor U44775 (N_44775,N_43430,N_43781);
and U44776 (N_44776,N_43646,N_43358);
xor U44777 (N_44777,N_43651,N_43221);
or U44778 (N_44778,N_43578,N_43547);
nand U44779 (N_44779,N_43178,N_43296);
or U44780 (N_44780,N_43588,N_43979);
and U44781 (N_44781,N_43107,N_43048);
nor U44782 (N_44782,N_43587,N_43597);
nor U44783 (N_44783,N_43750,N_43486);
and U44784 (N_44784,N_43598,N_43325);
and U44785 (N_44785,N_43640,N_43802);
xnor U44786 (N_44786,N_43140,N_43506);
and U44787 (N_44787,N_43628,N_43252);
nand U44788 (N_44788,N_43456,N_43756);
and U44789 (N_44789,N_43498,N_43268);
nor U44790 (N_44790,N_43574,N_43577);
nor U44791 (N_44791,N_43447,N_43071);
or U44792 (N_44792,N_43604,N_43491);
nor U44793 (N_44793,N_43853,N_43009);
and U44794 (N_44794,N_43805,N_43031);
and U44795 (N_44795,N_43968,N_43559);
nand U44796 (N_44796,N_43434,N_43284);
or U44797 (N_44797,N_43973,N_43221);
nor U44798 (N_44798,N_43073,N_43855);
xnor U44799 (N_44799,N_43983,N_43218);
nor U44800 (N_44800,N_43474,N_43608);
xor U44801 (N_44801,N_43282,N_43146);
xnor U44802 (N_44802,N_43039,N_43986);
xnor U44803 (N_44803,N_43030,N_43660);
and U44804 (N_44804,N_43626,N_43782);
and U44805 (N_44805,N_43959,N_43853);
nand U44806 (N_44806,N_43677,N_43048);
and U44807 (N_44807,N_43005,N_43699);
xnor U44808 (N_44808,N_43166,N_43572);
nand U44809 (N_44809,N_43340,N_43575);
and U44810 (N_44810,N_43738,N_43514);
and U44811 (N_44811,N_43167,N_43080);
nand U44812 (N_44812,N_43465,N_43215);
or U44813 (N_44813,N_43331,N_43938);
nand U44814 (N_44814,N_43236,N_43136);
or U44815 (N_44815,N_43941,N_43987);
or U44816 (N_44816,N_43811,N_43010);
nor U44817 (N_44817,N_43613,N_43497);
xnor U44818 (N_44818,N_43235,N_43989);
nand U44819 (N_44819,N_43850,N_43061);
or U44820 (N_44820,N_43383,N_43267);
or U44821 (N_44821,N_43771,N_43824);
xor U44822 (N_44822,N_43499,N_43006);
or U44823 (N_44823,N_43613,N_43385);
xnor U44824 (N_44824,N_43976,N_43263);
nand U44825 (N_44825,N_43624,N_43740);
or U44826 (N_44826,N_43852,N_43159);
nor U44827 (N_44827,N_43121,N_43073);
nor U44828 (N_44828,N_43641,N_43265);
and U44829 (N_44829,N_43624,N_43848);
nor U44830 (N_44830,N_43418,N_43161);
xor U44831 (N_44831,N_43765,N_43464);
xnor U44832 (N_44832,N_43934,N_43806);
nand U44833 (N_44833,N_43822,N_43104);
or U44834 (N_44834,N_43249,N_43724);
and U44835 (N_44835,N_43536,N_43151);
xor U44836 (N_44836,N_43942,N_43076);
nand U44837 (N_44837,N_43311,N_43152);
xnor U44838 (N_44838,N_43472,N_43024);
nor U44839 (N_44839,N_43555,N_43530);
xnor U44840 (N_44840,N_43766,N_43239);
nand U44841 (N_44841,N_43621,N_43241);
xor U44842 (N_44842,N_43613,N_43699);
xor U44843 (N_44843,N_43854,N_43572);
xor U44844 (N_44844,N_43515,N_43968);
or U44845 (N_44845,N_43600,N_43719);
or U44846 (N_44846,N_43187,N_43035);
nor U44847 (N_44847,N_43124,N_43361);
and U44848 (N_44848,N_43073,N_43742);
or U44849 (N_44849,N_43281,N_43098);
nand U44850 (N_44850,N_43523,N_43887);
xnor U44851 (N_44851,N_43856,N_43535);
and U44852 (N_44852,N_43499,N_43624);
and U44853 (N_44853,N_43267,N_43369);
xor U44854 (N_44854,N_43558,N_43181);
and U44855 (N_44855,N_43749,N_43644);
or U44856 (N_44856,N_43509,N_43622);
or U44857 (N_44857,N_43737,N_43311);
xor U44858 (N_44858,N_43652,N_43794);
nand U44859 (N_44859,N_43101,N_43086);
or U44860 (N_44860,N_43509,N_43613);
nand U44861 (N_44861,N_43696,N_43979);
or U44862 (N_44862,N_43459,N_43571);
or U44863 (N_44863,N_43100,N_43001);
xnor U44864 (N_44864,N_43682,N_43994);
nor U44865 (N_44865,N_43219,N_43306);
and U44866 (N_44866,N_43364,N_43785);
xnor U44867 (N_44867,N_43667,N_43268);
nor U44868 (N_44868,N_43008,N_43950);
nor U44869 (N_44869,N_43776,N_43089);
xor U44870 (N_44870,N_43802,N_43055);
or U44871 (N_44871,N_43091,N_43022);
nand U44872 (N_44872,N_43954,N_43666);
or U44873 (N_44873,N_43041,N_43786);
and U44874 (N_44874,N_43553,N_43193);
nand U44875 (N_44875,N_43129,N_43699);
and U44876 (N_44876,N_43835,N_43047);
nor U44877 (N_44877,N_43583,N_43898);
nand U44878 (N_44878,N_43693,N_43605);
or U44879 (N_44879,N_43986,N_43020);
xor U44880 (N_44880,N_43500,N_43255);
nand U44881 (N_44881,N_43397,N_43406);
nor U44882 (N_44882,N_43987,N_43638);
nor U44883 (N_44883,N_43504,N_43430);
nand U44884 (N_44884,N_43855,N_43447);
nand U44885 (N_44885,N_43294,N_43916);
or U44886 (N_44886,N_43058,N_43112);
xnor U44887 (N_44887,N_43924,N_43220);
nor U44888 (N_44888,N_43106,N_43157);
nor U44889 (N_44889,N_43523,N_43540);
nand U44890 (N_44890,N_43915,N_43252);
and U44891 (N_44891,N_43175,N_43960);
or U44892 (N_44892,N_43546,N_43715);
nand U44893 (N_44893,N_43311,N_43904);
and U44894 (N_44894,N_43630,N_43366);
nor U44895 (N_44895,N_43639,N_43985);
xnor U44896 (N_44896,N_43294,N_43192);
xor U44897 (N_44897,N_43310,N_43081);
or U44898 (N_44898,N_43011,N_43567);
nand U44899 (N_44899,N_43836,N_43871);
nand U44900 (N_44900,N_43959,N_43237);
nor U44901 (N_44901,N_43946,N_43918);
nor U44902 (N_44902,N_43113,N_43404);
xor U44903 (N_44903,N_43159,N_43445);
nand U44904 (N_44904,N_43475,N_43467);
xor U44905 (N_44905,N_43061,N_43001);
and U44906 (N_44906,N_43752,N_43320);
nor U44907 (N_44907,N_43903,N_43017);
nor U44908 (N_44908,N_43227,N_43377);
xor U44909 (N_44909,N_43413,N_43021);
or U44910 (N_44910,N_43729,N_43113);
or U44911 (N_44911,N_43777,N_43425);
nand U44912 (N_44912,N_43729,N_43691);
and U44913 (N_44913,N_43614,N_43807);
nor U44914 (N_44914,N_43117,N_43396);
or U44915 (N_44915,N_43774,N_43890);
nor U44916 (N_44916,N_43961,N_43491);
nand U44917 (N_44917,N_43119,N_43729);
or U44918 (N_44918,N_43447,N_43653);
nor U44919 (N_44919,N_43957,N_43483);
xnor U44920 (N_44920,N_43696,N_43482);
nor U44921 (N_44921,N_43469,N_43519);
or U44922 (N_44922,N_43966,N_43351);
or U44923 (N_44923,N_43365,N_43656);
nor U44924 (N_44924,N_43353,N_43477);
or U44925 (N_44925,N_43598,N_43697);
xnor U44926 (N_44926,N_43243,N_43204);
or U44927 (N_44927,N_43289,N_43271);
or U44928 (N_44928,N_43359,N_43101);
xor U44929 (N_44929,N_43468,N_43609);
nor U44930 (N_44930,N_43281,N_43647);
nand U44931 (N_44931,N_43019,N_43637);
nand U44932 (N_44932,N_43594,N_43548);
and U44933 (N_44933,N_43725,N_43826);
or U44934 (N_44934,N_43763,N_43341);
or U44935 (N_44935,N_43455,N_43189);
nor U44936 (N_44936,N_43668,N_43199);
and U44937 (N_44937,N_43839,N_43841);
or U44938 (N_44938,N_43677,N_43707);
and U44939 (N_44939,N_43334,N_43773);
nand U44940 (N_44940,N_43357,N_43814);
nor U44941 (N_44941,N_43748,N_43079);
or U44942 (N_44942,N_43583,N_43791);
nor U44943 (N_44943,N_43185,N_43156);
or U44944 (N_44944,N_43294,N_43571);
nor U44945 (N_44945,N_43836,N_43817);
xnor U44946 (N_44946,N_43599,N_43661);
xnor U44947 (N_44947,N_43711,N_43661);
xor U44948 (N_44948,N_43276,N_43482);
nor U44949 (N_44949,N_43278,N_43845);
and U44950 (N_44950,N_43906,N_43447);
or U44951 (N_44951,N_43421,N_43226);
nand U44952 (N_44952,N_43519,N_43181);
or U44953 (N_44953,N_43889,N_43267);
and U44954 (N_44954,N_43008,N_43285);
or U44955 (N_44955,N_43263,N_43561);
nand U44956 (N_44956,N_43943,N_43143);
and U44957 (N_44957,N_43104,N_43600);
nand U44958 (N_44958,N_43895,N_43620);
or U44959 (N_44959,N_43249,N_43053);
and U44960 (N_44960,N_43878,N_43569);
nor U44961 (N_44961,N_43487,N_43724);
xor U44962 (N_44962,N_43568,N_43631);
or U44963 (N_44963,N_43609,N_43030);
xnor U44964 (N_44964,N_43553,N_43368);
nand U44965 (N_44965,N_43708,N_43435);
nor U44966 (N_44966,N_43043,N_43364);
xor U44967 (N_44967,N_43852,N_43181);
xnor U44968 (N_44968,N_43720,N_43174);
nand U44969 (N_44969,N_43875,N_43272);
xnor U44970 (N_44970,N_43981,N_43966);
xnor U44971 (N_44971,N_43923,N_43805);
and U44972 (N_44972,N_43764,N_43032);
and U44973 (N_44973,N_43810,N_43065);
xor U44974 (N_44974,N_43475,N_43186);
or U44975 (N_44975,N_43732,N_43936);
nor U44976 (N_44976,N_43996,N_43503);
and U44977 (N_44977,N_43980,N_43088);
and U44978 (N_44978,N_43745,N_43930);
xnor U44979 (N_44979,N_43937,N_43387);
nand U44980 (N_44980,N_43984,N_43007);
xor U44981 (N_44981,N_43835,N_43541);
and U44982 (N_44982,N_43346,N_43036);
and U44983 (N_44983,N_43968,N_43134);
nor U44984 (N_44984,N_43387,N_43298);
and U44985 (N_44985,N_43543,N_43365);
or U44986 (N_44986,N_43683,N_43737);
and U44987 (N_44987,N_43046,N_43905);
and U44988 (N_44988,N_43931,N_43325);
nor U44989 (N_44989,N_43179,N_43071);
xnor U44990 (N_44990,N_43228,N_43215);
nand U44991 (N_44991,N_43660,N_43090);
and U44992 (N_44992,N_43166,N_43139);
nand U44993 (N_44993,N_43365,N_43385);
and U44994 (N_44994,N_43191,N_43964);
and U44995 (N_44995,N_43980,N_43992);
nor U44996 (N_44996,N_43622,N_43889);
xor U44997 (N_44997,N_43179,N_43741);
nor U44998 (N_44998,N_43355,N_43518);
xnor U44999 (N_44999,N_43895,N_43880);
nand U45000 (N_45000,N_44227,N_44226);
xor U45001 (N_45001,N_44687,N_44719);
xnor U45002 (N_45002,N_44834,N_44580);
and U45003 (N_45003,N_44981,N_44488);
and U45004 (N_45004,N_44955,N_44318);
xor U45005 (N_45005,N_44983,N_44200);
nand U45006 (N_45006,N_44904,N_44038);
nand U45007 (N_45007,N_44600,N_44937);
nor U45008 (N_45008,N_44124,N_44250);
and U45009 (N_45009,N_44511,N_44872);
xor U45010 (N_45010,N_44712,N_44796);
nand U45011 (N_45011,N_44662,N_44728);
nand U45012 (N_45012,N_44032,N_44592);
or U45013 (N_45013,N_44008,N_44210);
nor U45014 (N_45014,N_44532,N_44251);
and U45015 (N_45015,N_44099,N_44493);
xnor U45016 (N_45016,N_44054,N_44860);
xor U45017 (N_45017,N_44500,N_44522);
nand U45018 (N_45018,N_44174,N_44512);
xor U45019 (N_45019,N_44805,N_44982);
or U45020 (N_45020,N_44946,N_44173);
or U45021 (N_45021,N_44517,N_44507);
nand U45022 (N_45022,N_44827,N_44768);
and U45023 (N_45023,N_44783,N_44132);
xnor U45024 (N_45024,N_44801,N_44667);
nor U45025 (N_45025,N_44207,N_44420);
nor U45026 (N_45026,N_44128,N_44323);
nor U45027 (N_45027,N_44826,N_44903);
and U45028 (N_45028,N_44656,N_44570);
nand U45029 (N_45029,N_44997,N_44182);
nor U45030 (N_45030,N_44304,N_44724);
and U45031 (N_45031,N_44705,N_44336);
and U45032 (N_45032,N_44079,N_44635);
or U45033 (N_45033,N_44461,N_44327);
and U45034 (N_45034,N_44943,N_44622);
or U45035 (N_45035,N_44811,N_44542);
and U45036 (N_45036,N_44373,N_44450);
xor U45037 (N_45037,N_44579,N_44219);
and U45038 (N_45038,N_44411,N_44704);
xnor U45039 (N_45039,N_44252,N_44673);
and U45040 (N_45040,N_44764,N_44268);
xnor U45041 (N_45041,N_44028,N_44171);
and U45042 (N_45042,N_44134,N_44191);
nand U45043 (N_45043,N_44912,N_44299);
xor U45044 (N_45044,N_44740,N_44973);
or U45045 (N_45045,N_44264,N_44385);
nor U45046 (N_45046,N_44927,N_44059);
and U45047 (N_45047,N_44998,N_44524);
and U45048 (N_45048,N_44555,N_44310);
xor U45049 (N_45049,N_44588,N_44708);
and U45050 (N_45050,N_44302,N_44272);
nand U45051 (N_45051,N_44415,N_44193);
nor U45052 (N_45052,N_44989,N_44986);
and U45053 (N_45053,N_44551,N_44840);
nor U45054 (N_45054,N_44727,N_44694);
nand U45055 (N_45055,N_44976,N_44259);
xnor U45056 (N_45056,N_44154,N_44934);
nand U45057 (N_45057,N_44971,N_44351);
nor U45058 (N_45058,N_44926,N_44464);
and U45059 (N_45059,N_44473,N_44322);
xnor U45060 (N_45060,N_44942,N_44412);
xnor U45061 (N_45061,N_44651,N_44188);
nand U45062 (N_45062,N_44345,N_44342);
nor U45063 (N_45063,N_44218,N_44771);
or U45064 (N_45064,N_44388,N_44798);
and U45065 (N_45065,N_44626,N_44498);
or U45066 (N_45066,N_44557,N_44138);
and U45067 (N_45067,N_44936,N_44806);
and U45068 (N_45068,N_44329,N_44891);
nor U45069 (N_45069,N_44590,N_44599);
nand U45070 (N_45070,N_44325,N_44895);
nor U45071 (N_45071,N_44486,N_44122);
xor U45072 (N_45072,N_44562,N_44392);
nor U45073 (N_45073,N_44240,N_44568);
or U45074 (N_45074,N_44495,N_44567);
and U45075 (N_45075,N_44569,N_44540);
and U45076 (N_45076,N_44812,N_44841);
xor U45077 (N_45077,N_44100,N_44925);
nor U45078 (N_45078,N_44549,N_44383);
nand U45079 (N_45079,N_44509,N_44556);
and U45080 (N_45080,N_44108,N_44107);
nor U45081 (N_45081,N_44550,N_44781);
xor U45082 (N_45082,N_44497,N_44423);
and U45083 (N_45083,N_44065,N_44699);
nor U45084 (N_45084,N_44526,N_44095);
or U45085 (N_45085,N_44504,N_44893);
nor U45086 (N_45086,N_44166,N_44939);
or U45087 (N_45087,N_44127,N_44287);
xor U45088 (N_45088,N_44313,N_44445);
nand U45089 (N_45089,N_44585,N_44346);
xor U45090 (N_45090,N_44832,N_44915);
or U45091 (N_45091,N_44275,N_44571);
nor U45092 (N_45092,N_44399,N_44309);
xor U45093 (N_45093,N_44460,N_44073);
nor U45094 (N_45094,N_44503,N_44822);
xnor U45095 (N_45095,N_44737,N_44746);
nand U45096 (N_45096,N_44089,N_44485);
and U45097 (N_45097,N_44417,N_44959);
nand U45098 (N_45098,N_44804,N_44396);
nand U45099 (N_45099,N_44916,N_44470);
xor U45100 (N_45100,N_44075,N_44772);
or U45101 (N_45101,N_44372,N_44199);
nand U45102 (N_45102,N_44594,N_44255);
nand U45103 (N_45103,N_44917,N_44401);
and U45104 (N_45104,N_44713,N_44839);
or U45105 (N_45105,N_44686,N_44766);
nor U45106 (N_45106,N_44559,N_44755);
and U45107 (N_45107,N_44231,N_44456);
nand U45108 (N_45108,N_44378,N_44204);
xor U45109 (N_45109,N_44198,N_44665);
nand U45110 (N_45110,N_44121,N_44865);
nand U45111 (N_45111,N_44036,N_44640);
nand U45112 (N_45112,N_44066,N_44744);
xor U45113 (N_45113,N_44723,N_44950);
nor U45114 (N_45114,N_44326,N_44466);
nand U45115 (N_45115,N_44085,N_44448);
xor U45116 (N_45116,N_44162,N_44043);
xor U45117 (N_45117,N_44969,N_44717);
and U45118 (N_45118,N_44220,N_44985);
xnor U45119 (N_45119,N_44364,N_44753);
nor U45120 (N_45120,N_44087,N_44561);
or U45121 (N_45121,N_44483,N_44523);
or U45122 (N_45122,N_44676,N_44301);
nand U45123 (N_45123,N_44340,N_44024);
and U45124 (N_45124,N_44633,N_44775);
nor U45125 (N_45125,N_44106,N_44685);
xor U45126 (N_45126,N_44047,N_44894);
nor U45127 (N_45127,N_44869,N_44823);
or U45128 (N_45128,N_44791,N_44945);
nor U45129 (N_45129,N_44238,N_44745);
nor U45130 (N_45130,N_44501,N_44896);
and U45131 (N_45131,N_44076,N_44765);
nor U45132 (N_45132,N_44332,N_44666);
or U45133 (N_45133,N_44920,N_44877);
and U45134 (N_45134,N_44867,N_44232);
or U45135 (N_45135,N_44019,N_44115);
xor U45136 (N_45136,N_44289,N_44111);
nand U45137 (N_45137,N_44056,N_44664);
xnor U45138 (N_45138,N_44844,N_44416);
xnor U45139 (N_45139,N_44990,N_44968);
or U45140 (N_45140,N_44938,N_44695);
nand U45141 (N_45141,N_44725,N_44082);
and U45142 (N_45142,N_44675,N_44113);
nor U45143 (N_45143,N_44975,N_44808);
and U45144 (N_45144,N_44021,N_44952);
xnor U45145 (N_45145,N_44991,N_44129);
or U45146 (N_45146,N_44184,N_44492);
xor U45147 (N_45147,N_44478,N_44649);
and U45148 (N_45148,N_44465,N_44978);
nor U45149 (N_45149,N_44148,N_44018);
or U45150 (N_45150,N_44350,N_44883);
nand U45151 (N_45151,N_44928,N_44145);
xnor U45152 (N_45152,N_44449,N_44209);
or U45153 (N_45153,N_44335,N_44546);
xnor U45154 (N_45154,N_44026,N_44947);
xor U45155 (N_45155,N_44352,N_44842);
nand U45156 (N_45156,N_44609,N_44314);
or U45157 (N_45157,N_44317,N_44064);
nor U45158 (N_45158,N_44042,N_44119);
nor U45159 (N_45159,N_44888,N_44677);
and U45160 (N_45160,N_44636,N_44838);
or U45161 (N_45161,N_44126,N_44970);
nor U45162 (N_45162,N_44147,N_44203);
nor U45163 (N_45163,N_44312,N_44527);
nand U45164 (N_45164,N_44341,N_44587);
and U45165 (N_45165,N_44573,N_44566);
or U45166 (N_45166,N_44446,N_44881);
nor U45167 (N_45167,N_44797,N_44157);
nor U45168 (N_45168,N_44631,N_44670);
and U45169 (N_45169,N_44830,N_44294);
nand U45170 (N_45170,N_44786,N_44691);
or U45171 (N_45171,N_44280,N_44821);
xor U45172 (N_45172,N_44052,N_44980);
and U45173 (N_45173,N_44290,N_44552);
or U45174 (N_45174,N_44790,N_44363);
or U45175 (N_45175,N_44593,N_44529);
or U45176 (N_45176,N_44836,N_44105);
nor U45177 (N_45177,N_44776,N_44964);
nor U45178 (N_45178,N_44703,N_44907);
and U45179 (N_45179,N_44576,N_44288);
nand U45180 (N_45180,N_44505,N_44647);
nor U45181 (N_45181,N_44544,N_44164);
or U45182 (N_45182,N_44262,N_44393);
xnor U45183 (N_45183,N_44086,N_44884);
and U45184 (N_45184,N_44453,N_44381);
nor U45185 (N_45185,N_44878,N_44586);
nand U45186 (N_45186,N_44109,N_44992);
and U45187 (N_45187,N_44469,N_44192);
and U45188 (N_45188,N_44330,N_44815);
or U45189 (N_45189,N_44595,N_44131);
nor U45190 (N_45190,N_44333,N_44875);
or U45191 (N_45191,N_44077,N_44924);
nand U45192 (N_45192,N_44400,N_44856);
xnor U45193 (N_45193,N_44053,N_44023);
or U45194 (N_45194,N_44063,N_44539);
nand U45195 (N_45195,N_44168,N_44607);
nor U45196 (N_45196,N_44291,N_44040);
or U45197 (N_45197,N_44833,N_44092);
or U45198 (N_45198,N_44117,N_44030);
and U45199 (N_45199,N_44462,N_44621);
xor U45200 (N_45200,N_44463,N_44484);
nor U45201 (N_45201,N_44361,N_44663);
xor U45202 (N_45202,N_44810,N_44426);
xnor U45203 (N_45203,N_44496,N_44792);
nand U45204 (N_45204,N_44906,N_44919);
nand U45205 (N_45205,N_44818,N_44292);
or U45206 (N_45206,N_44515,N_44305);
xor U45207 (N_45207,N_44929,N_44404);
or U45208 (N_45208,N_44679,N_44747);
or U45209 (N_45209,N_44851,N_44222);
xor U45210 (N_45210,N_44311,N_44398);
or U45211 (N_45211,N_44560,N_44799);
xnor U45212 (N_45212,N_44530,N_44254);
nand U45213 (N_45213,N_44265,N_44338);
or U45214 (N_45214,N_44803,N_44889);
and U45215 (N_45215,N_44375,N_44366);
xor U45216 (N_45216,N_44433,N_44974);
or U45217 (N_45217,N_44002,N_44468);
or U45218 (N_45218,N_44178,N_44369);
nand U45219 (N_45219,N_44435,N_44578);
and U45220 (N_45220,N_44324,N_44853);
nand U45221 (N_45221,N_44951,N_44247);
and U45222 (N_45222,N_44732,N_44103);
nor U45223 (N_45223,N_44655,N_44613);
and U45224 (N_45224,N_44236,N_44538);
or U45225 (N_45225,N_44116,N_44283);
nand U45226 (N_45226,N_44244,N_44359);
xor U45227 (N_45227,N_44591,N_44558);
nand U45228 (N_45228,N_44758,N_44293);
and U45229 (N_45229,N_44189,N_44885);
or U45230 (N_45230,N_44239,N_44221);
xnor U45231 (N_45231,N_44431,N_44554);
nand U45232 (N_45232,N_44223,N_44582);
and U45233 (N_45233,N_44152,N_44405);
and U45234 (N_45234,N_44669,N_44807);
nor U45235 (N_45235,N_44697,N_44390);
and U45236 (N_45236,N_44279,N_44020);
nor U45237 (N_45237,N_44824,N_44348);
nand U45238 (N_45238,N_44093,N_44958);
or U45239 (N_45239,N_44306,N_44360);
or U45240 (N_45240,N_44682,N_44577);
or U45241 (N_45241,N_44729,N_44535);
xnor U45242 (N_45242,N_44545,N_44726);
xor U45243 (N_45243,N_44909,N_44614);
xnor U45244 (N_45244,N_44611,N_44606);
xor U45245 (N_45245,N_44049,N_44035);
xor U45246 (N_45246,N_44062,N_44274);
or U45247 (N_45247,N_44357,N_44961);
nor U45248 (N_45248,N_44996,N_44094);
xor U45249 (N_45249,N_44374,N_44637);
or U45250 (N_45250,N_44718,N_44706);
nand U45251 (N_45251,N_44006,N_44295);
nand U45252 (N_45252,N_44347,N_44045);
nor U45253 (N_45253,N_44604,N_44197);
or U45254 (N_45254,N_44900,N_44443);
xor U45255 (N_45255,N_44419,N_44646);
xor U45256 (N_45256,N_44722,N_44521);
or U45257 (N_45257,N_44457,N_44367);
nor U45258 (N_45258,N_44653,N_44855);
nand U45259 (N_45259,N_44658,N_44858);
xnor U45260 (N_45260,N_44584,N_44785);
and U45261 (N_45261,N_44954,N_44337);
xnor U45262 (N_45262,N_44245,N_44410);
and U45263 (N_45263,N_44910,N_44782);
nor U45264 (N_45264,N_44080,N_44820);
or U45265 (N_45265,N_44300,N_44413);
or U45266 (N_45266,N_44321,N_44652);
and U45267 (N_45267,N_44487,N_44137);
xor U45268 (N_45268,N_44356,N_44763);
or U45269 (N_45269,N_44146,N_44931);
or U45270 (N_45270,N_44257,N_44169);
or U45271 (N_45271,N_44050,N_44683);
xnor U45272 (N_45272,N_44183,N_44537);
and U45273 (N_45273,N_44948,N_44155);
nand U45274 (N_45274,N_44001,N_44143);
xor U45275 (N_45275,N_44354,N_44848);
and U45276 (N_45276,N_44102,N_44194);
nor U45277 (N_45277,N_44418,N_44380);
nand U45278 (N_45278,N_44657,N_44778);
nand U45279 (N_45279,N_44344,N_44572);
xor U45280 (N_45280,N_44794,N_44767);
or U45281 (N_45281,N_44861,N_44510);
and U45282 (N_45282,N_44260,N_44328);
xnor U45283 (N_45283,N_44068,N_44632);
xnor U45284 (N_45284,N_44849,N_44010);
nor U45285 (N_45285,N_44692,N_44882);
nor U45286 (N_45286,N_44932,N_44273);
or U45287 (N_45287,N_44266,N_44714);
nand U45288 (N_45288,N_44541,N_44874);
nand U45289 (N_45289,N_44972,N_44034);
or U45290 (N_45290,N_44616,N_44857);
and U45291 (N_45291,N_44846,N_44014);
nor U45292 (N_45292,N_44368,N_44905);
nor U45293 (N_45293,N_44436,N_44644);
xnor U45294 (N_45294,N_44430,N_44788);
xor U45295 (N_45295,N_44196,N_44620);
or U45296 (N_45296,N_44270,N_44721);
or U45297 (N_45297,N_44009,N_44455);
or U45298 (N_45298,N_44596,N_44170);
nand U45299 (N_45299,N_44256,N_44422);
xor U45300 (N_45300,N_44165,N_44012);
xor U45301 (N_45301,N_44271,N_44731);
nor U45302 (N_45302,N_44136,N_44612);
xor U45303 (N_45303,N_44852,N_44733);
and U45304 (N_45304,N_44060,N_44118);
and U45305 (N_45305,N_44097,N_44144);
nand U45306 (N_45306,N_44475,N_44589);
nand U45307 (N_45307,N_44355,N_44862);
nor U45308 (N_45308,N_44711,N_44130);
or U45309 (N_45309,N_44802,N_44847);
xor U45310 (N_45310,N_44984,N_44813);
nand U45311 (N_45311,N_44605,N_44941);
nand U45312 (N_45312,N_44837,N_44243);
xor U45313 (N_45313,N_44298,N_44843);
xnor U45314 (N_45314,N_44513,N_44402);
nand U45315 (N_45315,N_44003,N_44071);
xor U45316 (N_45316,N_44048,N_44819);
and U45317 (N_45317,N_44701,N_44278);
or U45318 (N_45318,N_44681,N_44756);
nand U45319 (N_45319,N_44707,N_44615);
nor U45320 (N_45320,N_44979,N_44583);
nand U45321 (N_45321,N_44242,N_44353);
xor U45322 (N_45322,N_44751,N_44386);
nand U45323 (N_45323,N_44993,N_44994);
xnor U45324 (N_45324,N_44966,N_44142);
xor U45325 (N_45325,N_44999,N_44514);
nor U45326 (N_45326,N_44565,N_44234);
nand U45327 (N_45327,N_44736,N_44689);
and U45328 (N_45328,N_44151,N_44389);
or U45329 (N_45329,N_44634,N_44957);
xnor U45330 (N_45330,N_44519,N_44286);
and U45331 (N_45331,N_44141,N_44114);
nand U45332 (N_45332,N_44516,N_44334);
xor U45333 (N_45333,N_44602,N_44025);
nor U45334 (N_45334,N_44308,N_44447);
nor U45335 (N_45335,N_44007,N_44960);
and U45336 (N_45336,N_44525,N_44437);
or U45337 (N_45337,N_44414,N_44956);
nand U45338 (N_45338,N_44693,N_44000);
and U45339 (N_45339,N_44090,N_44454);
xnor U45340 (N_45340,N_44949,N_44135);
nor U45341 (N_45341,N_44285,N_44284);
and U45342 (N_45342,N_44228,N_44391);
or U45343 (N_45343,N_44809,N_44702);
or U45344 (N_45344,N_44491,N_44015);
xor U45345 (N_45345,N_44828,N_44490);
and U45346 (N_45346,N_44603,N_44214);
nor U45347 (N_45347,N_44112,N_44215);
or U45348 (N_45348,N_44133,N_44459);
nor U45349 (N_45349,N_44269,N_44033);
xnor U45350 (N_45350,N_44617,N_44027);
or U45351 (N_45351,N_44850,N_44547);
or U45352 (N_45352,N_44678,N_44738);
xor U45353 (N_45353,N_44988,N_44930);
xor U45354 (N_45354,N_44779,N_44749);
nor U45355 (N_45355,N_44403,N_44267);
or U45356 (N_45356,N_44349,N_44476);
and U45357 (N_45357,N_44083,N_44235);
or U45358 (N_45358,N_44752,N_44660);
and U45359 (N_45359,N_44377,N_44709);
nand U45360 (N_45360,N_44831,N_44069);
nor U45361 (N_45361,N_44520,N_44246);
nand U45362 (N_45362,N_44777,N_44908);
xor U45363 (N_45363,N_44070,N_44923);
nand U45364 (N_45364,N_44854,N_44225);
or U45365 (N_45365,N_44716,N_44471);
and U45366 (N_45366,N_44690,N_44379);
nor U45367 (N_45367,N_44784,N_44172);
xnor U45368 (N_45368,N_44201,N_44870);
and U45369 (N_45369,N_44987,N_44084);
and U45370 (N_45370,N_44759,N_44921);
nand U45371 (N_45371,N_44125,N_44481);
xnor U45372 (N_45372,N_44918,N_44425);
nand U45373 (N_45373,N_44659,N_44452);
nor U45374 (N_45374,N_44922,N_44276);
and U45375 (N_45375,N_44187,N_44123);
nand U45376 (N_45376,N_44742,N_44902);
and U45377 (N_45377,N_44494,N_44444);
nor U45378 (N_45378,N_44536,N_44029);
and U45379 (N_45379,N_44741,N_44041);
xor U45380 (N_45380,N_44757,N_44163);
nor U45381 (N_45381,N_44773,N_44899);
nand U45382 (N_45382,N_44409,N_44533);
xnor U45383 (N_45383,N_44627,N_44362);
nor U45384 (N_45384,N_44382,N_44153);
xnor U45385 (N_45385,N_44654,N_44962);
nor U45386 (N_45386,N_44179,N_44057);
nor U45387 (N_45387,N_44046,N_44205);
or U45388 (N_45388,N_44864,N_44940);
nor U45389 (N_45389,N_44307,N_44074);
nand U45390 (N_45390,N_44261,N_44508);
xor U45391 (N_45391,N_44574,N_44316);
nor U45392 (N_45392,N_44282,N_44743);
or U45393 (N_45393,N_44458,N_44671);
nand U45394 (N_45394,N_44072,N_44158);
and U45395 (N_45395,N_44249,N_44868);
xnor U45396 (N_45396,N_44110,N_44022);
nand U45397 (N_45397,N_44467,N_44428);
and U45398 (N_45398,N_44720,N_44630);
xnor U45399 (N_45399,N_44429,N_44296);
or U45400 (N_45400,N_44281,N_44167);
nand U45401 (N_45401,N_44237,N_44224);
xnor U45402 (N_45402,N_44977,N_44104);
and U45403 (N_45403,N_44387,N_44963);
nand U45404 (N_45404,N_44780,N_44177);
and U45405 (N_45405,N_44610,N_44700);
and U45406 (N_45406,N_44863,N_44186);
or U45407 (N_45407,N_44175,N_44553);
and U45408 (N_45408,N_44639,N_44217);
and U45409 (N_45409,N_44037,N_44031);
and U45410 (N_45410,N_44421,N_44795);
or U45411 (N_45411,N_44735,N_44672);
and U45412 (N_45412,N_44575,N_44879);
nand U45413 (N_45413,N_44674,N_44935);
nor U45414 (N_45414,N_44543,N_44208);
or U45415 (N_45415,N_44160,N_44734);
and U45416 (N_45416,N_44394,N_44371);
xnor U45417 (N_45417,N_44581,N_44098);
and U45418 (N_45418,N_44176,N_44845);
and U45419 (N_45419,N_44432,N_44642);
nor U45420 (N_45420,N_44370,N_44880);
nor U45421 (N_45421,N_44156,N_44897);
or U45422 (N_45422,N_44814,N_44442);
nor U45423 (N_45423,N_44750,N_44229);
nand U45424 (N_45424,N_44898,N_44715);
xnor U45425 (N_45425,N_44339,N_44206);
nor U45426 (N_45426,N_44303,N_44619);
and U45427 (N_45427,N_44608,N_44518);
or U45428 (N_45428,N_44039,N_44629);
nor U45429 (N_45429,N_44887,N_44424);
nor U45430 (N_45430,N_44597,N_44789);
and U45431 (N_45431,N_44078,N_44835);
nand U45432 (N_45432,N_44953,N_44185);
or U45433 (N_45433,N_44531,N_44866);
xnor U45434 (N_45434,N_44161,N_44051);
nand U45435 (N_45435,N_44004,N_44451);
xnor U45436 (N_45436,N_44564,N_44598);
nor U45437 (N_45437,N_44438,N_44623);
nand U45438 (N_45438,N_44376,N_44101);
xnor U45439 (N_45439,N_44216,N_44648);
nor U45440 (N_45440,N_44770,N_44624);
and U45441 (N_45441,N_44253,N_44825);
xnor U45442 (N_45442,N_44965,N_44358);
xnor U45443 (N_45443,N_44913,N_44774);
nand U45444 (N_45444,N_44650,N_44159);
nand U45445 (N_45445,N_44195,N_44061);
nand U45446 (N_45446,N_44914,N_44748);
or U45447 (N_45447,N_44933,N_44876);
and U45448 (N_45448,N_44044,N_44408);
and U45449 (N_45449,N_44761,N_44730);
and U45450 (N_45450,N_44213,N_44793);
nor U45451 (N_45451,N_44739,N_44427);
xor U45452 (N_45452,N_44331,N_44440);
or U45453 (N_45453,N_44625,N_44890);
nand U45454 (N_45454,N_44754,N_44474);
xor U45455 (N_45455,N_44397,N_44055);
xnor U45456 (N_45456,N_44067,N_44871);
or U45457 (N_45457,N_44482,N_44563);
or U45458 (N_45458,N_44762,N_44150);
and U45459 (N_45459,N_44181,N_44091);
xor U45460 (N_45460,N_44011,N_44944);
xor U45461 (N_45461,N_44816,N_44016);
nand U45462 (N_45462,N_44698,N_44502);
xnor U45463 (N_45463,N_44829,N_44233);
or U45464 (N_45464,N_44548,N_44787);
nor U45465 (N_45465,N_44241,N_44995);
and U45466 (N_45466,N_44297,N_44439);
nor U45467 (N_45467,N_44489,N_44661);
xor U45468 (N_45468,N_44441,N_44534);
or U45469 (N_45469,N_44202,N_44760);
and U45470 (N_45470,N_44499,N_44017);
nor U45471 (N_45471,N_44277,N_44601);
xor U45472 (N_45472,N_44472,N_44013);
or U45473 (N_45473,N_44696,N_44149);
or U45474 (N_45474,N_44190,N_44479);
xor U45475 (N_45475,N_44406,N_44506);
and U45476 (N_45476,N_44628,N_44480);
nor U45477 (N_45477,N_44096,N_44817);
nand U45478 (N_45478,N_44873,N_44365);
or U45479 (N_45479,N_44407,N_44320);
nand U45480 (N_45480,N_44230,N_44319);
xor U45481 (N_45481,N_44081,N_44248);
nand U45482 (N_45482,N_44892,N_44211);
nand U45483 (N_45483,N_44005,N_44139);
or U45484 (N_45484,N_44859,N_44800);
or U45485 (N_45485,N_44688,N_44180);
and U45486 (N_45486,N_44684,N_44088);
nor U45487 (N_45487,N_44901,N_44434);
nand U45488 (N_45488,N_44710,N_44668);
nand U45489 (N_45489,N_44911,N_44618);
or U45490 (N_45490,N_44769,N_44120);
or U45491 (N_45491,N_44258,N_44395);
or U45492 (N_45492,N_44886,N_44343);
and U45493 (N_45493,N_44645,N_44384);
xor U45494 (N_45494,N_44638,N_44212);
and U45495 (N_45495,N_44140,N_44528);
or U45496 (N_45496,N_44477,N_44967);
or U45497 (N_45497,N_44680,N_44643);
nand U45498 (N_45498,N_44315,N_44058);
nand U45499 (N_45499,N_44641,N_44263);
nor U45500 (N_45500,N_44646,N_44157);
and U45501 (N_45501,N_44601,N_44979);
nand U45502 (N_45502,N_44478,N_44180);
nor U45503 (N_45503,N_44134,N_44669);
or U45504 (N_45504,N_44753,N_44641);
nor U45505 (N_45505,N_44026,N_44591);
nand U45506 (N_45506,N_44711,N_44807);
nor U45507 (N_45507,N_44029,N_44499);
xor U45508 (N_45508,N_44695,N_44352);
nand U45509 (N_45509,N_44149,N_44243);
and U45510 (N_45510,N_44855,N_44514);
xnor U45511 (N_45511,N_44753,N_44234);
nor U45512 (N_45512,N_44964,N_44364);
xor U45513 (N_45513,N_44016,N_44142);
and U45514 (N_45514,N_44437,N_44527);
nor U45515 (N_45515,N_44974,N_44641);
nor U45516 (N_45516,N_44708,N_44444);
or U45517 (N_45517,N_44644,N_44324);
nor U45518 (N_45518,N_44287,N_44422);
or U45519 (N_45519,N_44302,N_44288);
and U45520 (N_45520,N_44853,N_44241);
nor U45521 (N_45521,N_44507,N_44109);
xor U45522 (N_45522,N_44760,N_44612);
nor U45523 (N_45523,N_44207,N_44858);
xor U45524 (N_45524,N_44467,N_44582);
nor U45525 (N_45525,N_44464,N_44493);
and U45526 (N_45526,N_44492,N_44671);
nor U45527 (N_45527,N_44948,N_44259);
or U45528 (N_45528,N_44573,N_44639);
and U45529 (N_45529,N_44355,N_44962);
nand U45530 (N_45530,N_44624,N_44368);
nor U45531 (N_45531,N_44644,N_44137);
nor U45532 (N_45532,N_44767,N_44662);
nand U45533 (N_45533,N_44819,N_44552);
xnor U45534 (N_45534,N_44666,N_44368);
nand U45535 (N_45535,N_44020,N_44458);
nor U45536 (N_45536,N_44474,N_44531);
nand U45537 (N_45537,N_44836,N_44610);
nand U45538 (N_45538,N_44074,N_44883);
or U45539 (N_45539,N_44613,N_44706);
and U45540 (N_45540,N_44722,N_44204);
nand U45541 (N_45541,N_44403,N_44390);
and U45542 (N_45542,N_44668,N_44977);
nor U45543 (N_45543,N_44124,N_44370);
or U45544 (N_45544,N_44358,N_44488);
and U45545 (N_45545,N_44272,N_44181);
nor U45546 (N_45546,N_44459,N_44775);
nand U45547 (N_45547,N_44007,N_44103);
nor U45548 (N_45548,N_44341,N_44655);
nor U45549 (N_45549,N_44506,N_44129);
nand U45550 (N_45550,N_44783,N_44963);
xor U45551 (N_45551,N_44040,N_44490);
nand U45552 (N_45552,N_44279,N_44869);
or U45553 (N_45553,N_44268,N_44631);
nor U45554 (N_45554,N_44219,N_44677);
and U45555 (N_45555,N_44448,N_44566);
and U45556 (N_45556,N_44042,N_44669);
nor U45557 (N_45557,N_44753,N_44987);
nand U45558 (N_45558,N_44139,N_44290);
or U45559 (N_45559,N_44373,N_44853);
xnor U45560 (N_45560,N_44510,N_44562);
or U45561 (N_45561,N_44365,N_44031);
and U45562 (N_45562,N_44942,N_44425);
nand U45563 (N_45563,N_44746,N_44533);
or U45564 (N_45564,N_44380,N_44979);
and U45565 (N_45565,N_44850,N_44829);
and U45566 (N_45566,N_44432,N_44482);
and U45567 (N_45567,N_44771,N_44126);
xor U45568 (N_45568,N_44109,N_44307);
nand U45569 (N_45569,N_44996,N_44857);
nor U45570 (N_45570,N_44904,N_44528);
nor U45571 (N_45571,N_44395,N_44354);
nor U45572 (N_45572,N_44722,N_44439);
or U45573 (N_45573,N_44229,N_44168);
nand U45574 (N_45574,N_44770,N_44060);
or U45575 (N_45575,N_44598,N_44592);
nor U45576 (N_45576,N_44019,N_44248);
nor U45577 (N_45577,N_44301,N_44870);
nor U45578 (N_45578,N_44141,N_44738);
nand U45579 (N_45579,N_44581,N_44577);
nand U45580 (N_45580,N_44515,N_44616);
xor U45581 (N_45581,N_44644,N_44009);
and U45582 (N_45582,N_44573,N_44904);
nor U45583 (N_45583,N_44824,N_44828);
xnor U45584 (N_45584,N_44521,N_44131);
and U45585 (N_45585,N_44220,N_44979);
and U45586 (N_45586,N_44525,N_44267);
xor U45587 (N_45587,N_44842,N_44878);
and U45588 (N_45588,N_44556,N_44734);
and U45589 (N_45589,N_44841,N_44895);
or U45590 (N_45590,N_44070,N_44456);
and U45591 (N_45591,N_44437,N_44379);
or U45592 (N_45592,N_44576,N_44313);
or U45593 (N_45593,N_44665,N_44421);
nor U45594 (N_45594,N_44155,N_44653);
and U45595 (N_45595,N_44317,N_44676);
or U45596 (N_45596,N_44574,N_44002);
nor U45597 (N_45597,N_44481,N_44861);
or U45598 (N_45598,N_44471,N_44014);
nor U45599 (N_45599,N_44898,N_44636);
xnor U45600 (N_45600,N_44704,N_44660);
nor U45601 (N_45601,N_44449,N_44921);
and U45602 (N_45602,N_44129,N_44013);
xor U45603 (N_45603,N_44062,N_44043);
or U45604 (N_45604,N_44030,N_44157);
xor U45605 (N_45605,N_44252,N_44475);
or U45606 (N_45606,N_44212,N_44260);
nor U45607 (N_45607,N_44438,N_44232);
xor U45608 (N_45608,N_44026,N_44703);
nor U45609 (N_45609,N_44423,N_44566);
and U45610 (N_45610,N_44421,N_44817);
nand U45611 (N_45611,N_44078,N_44196);
nand U45612 (N_45612,N_44588,N_44753);
and U45613 (N_45613,N_44871,N_44004);
and U45614 (N_45614,N_44458,N_44284);
or U45615 (N_45615,N_44890,N_44301);
or U45616 (N_45616,N_44806,N_44840);
xor U45617 (N_45617,N_44350,N_44050);
or U45618 (N_45618,N_44009,N_44836);
xor U45619 (N_45619,N_44895,N_44216);
nand U45620 (N_45620,N_44094,N_44117);
nand U45621 (N_45621,N_44852,N_44602);
and U45622 (N_45622,N_44398,N_44131);
nor U45623 (N_45623,N_44070,N_44397);
and U45624 (N_45624,N_44926,N_44558);
and U45625 (N_45625,N_44035,N_44525);
nand U45626 (N_45626,N_44948,N_44554);
xnor U45627 (N_45627,N_44746,N_44532);
and U45628 (N_45628,N_44958,N_44187);
or U45629 (N_45629,N_44533,N_44131);
nor U45630 (N_45630,N_44734,N_44250);
nand U45631 (N_45631,N_44341,N_44726);
nor U45632 (N_45632,N_44216,N_44837);
and U45633 (N_45633,N_44975,N_44465);
and U45634 (N_45634,N_44285,N_44644);
nor U45635 (N_45635,N_44904,N_44674);
or U45636 (N_45636,N_44484,N_44233);
nor U45637 (N_45637,N_44528,N_44550);
and U45638 (N_45638,N_44018,N_44496);
nand U45639 (N_45639,N_44411,N_44100);
xnor U45640 (N_45640,N_44883,N_44849);
xnor U45641 (N_45641,N_44468,N_44985);
xor U45642 (N_45642,N_44301,N_44493);
or U45643 (N_45643,N_44868,N_44779);
nor U45644 (N_45644,N_44913,N_44069);
or U45645 (N_45645,N_44029,N_44045);
nand U45646 (N_45646,N_44750,N_44718);
and U45647 (N_45647,N_44366,N_44093);
or U45648 (N_45648,N_44062,N_44499);
and U45649 (N_45649,N_44651,N_44408);
nand U45650 (N_45650,N_44105,N_44679);
and U45651 (N_45651,N_44264,N_44378);
or U45652 (N_45652,N_44976,N_44225);
and U45653 (N_45653,N_44429,N_44835);
nand U45654 (N_45654,N_44122,N_44629);
or U45655 (N_45655,N_44434,N_44630);
xnor U45656 (N_45656,N_44857,N_44646);
xor U45657 (N_45657,N_44341,N_44725);
and U45658 (N_45658,N_44936,N_44706);
nor U45659 (N_45659,N_44362,N_44285);
xnor U45660 (N_45660,N_44180,N_44630);
nor U45661 (N_45661,N_44326,N_44922);
nand U45662 (N_45662,N_44212,N_44956);
nand U45663 (N_45663,N_44070,N_44844);
or U45664 (N_45664,N_44396,N_44229);
and U45665 (N_45665,N_44965,N_44773);
and U45666 (N_45666,N_44921,N_44770);
and U45667 (N_45667,N_44300,N_44381);
nand U45668 (N_45668,N_44280,N_44873);
and U45669 (N_45669,N_44473,N_44389);
nand U45670 (N_45670,N_44294,N_44846);
nor U45671 (N_45671,N_44984,N_44933);
xnor U45672 (N_45672,N_44916,N_44548);
nand U45673 (N_45673,N_44398,N_44119);
nor U45674 (N_45674,N_44123,N_44839);
xor U45675 (N_45675,N_44693,N_44301);
or U45676 (N_45676,N_44410,N_44545);
and U45677 (N_45677,N_44886,N_44469);
nand U45678 (N_45678,N_44309,N_44403);
nor U45679 (N_45679,N_44031,N_44731);
xor U45680 (N_45680,N_44845,N_44831);
and U45681 (N_45681,N_44064,N_44354);
nor U45682 (N_45682,N_44840,N_44738);
nand U45683 (N_45683,N_44662,N_44920);
xnor U45684 (N_45684,N_44756,N_44797);
or U45685 (N_45685,N_44068,N_44754);
xnor U45686 (N_45686,N_44242,N_44757);
xor U45687 (N_45687,N_44877,N_44761);
and U45688 (N_45688,N_44762,N_44248);
nand U45689 (N_45689,N_44249,N_44944);
nor U45690 (N_45690,N_44088,N_44924);
and U45691 (N_45691,N_44556,N_44888);
or U45692 (N_45692,N_44170,N_44911);
nor U45693 (N_45693,N_44912,N_44573);
xnor U45694 (N_45694,N_44657,N_44223);
or U45695 (N_45695,N_44089,N_44958);
nor U45696 (N_45696,N_44711,N_44783);
nand U45697 (N_45697,N_44562,N_44542);
and U45698 (N_45698,N_44193,N_44642);
xnor U45699 (N_45699,N_44900,N_44698);
xor U45700 (N_45700,N_44479,N_44364);
or U45701 (N_45701,N_44881,N_44274);
nand U45702 (N_45702,N_44786,N_44040);
xnor U45703 (N_45703,N_44551,N_44490);
nand U45704 (N_45704,N_44847,N_44512);
nor U45705 (N_45705,N_44936,N_44275);
or U45706 (N_45706,N_44347,N_44942);
nand U45707 (N_45707,N_44550,N_44262);
xnor U45708 (N_45708,N_44930,N_44345);
or U45709 (N_45709,N_44100,N_44588);
nor U45710 (N_45710,N_44518,N_44082);
xnor U45711 (N_45711,N_44338,N_44200);
xnor U45712 (N_45712,N_44139,N_44598);
or U45713 (N_45713,N_44225,N_44830);
xnor U45714 (N_45714,N_44251,N_44531);
xnor U45715 (N_45715,N_44908,N_44155);
and U45716 (N_45716,N_44040,N_44478);
nor U45717 (N_45717,N_44289,N_44784);
nand U45718 (N_45718,N_44779,N_44063);
nand U45719 (N_45719,N_44449,N_44320);
or U45720 (N_45720,N_44592,N_44881);
or U45721 (N_45721,N_44563,N_44457);
nor U45722 (N_45722,N_44482,N_44097);
or U45723 (N_45723,N_44200,N_44423);
nand U45724 (N_45724,N_44541,N_44751);
nor U45725 (N_45725,N_44004,N_44941);
or U45726 (N_45726,N_44929,N_44979);
nand U45727 (N_45727,N_44403,N_44584);
or U45728 (N_45728,N_44679,N_44794);
and U45729 (N_45729,N_44856,N_44466);
nand U45730 (N_45730,N_44094,N_44731);
nor U45731 (N_45731,N_44549,N_44236);
xnor U45732 (N_45732,N_44594,N_44565);
nor U45733 (N_45733,N_44992,N_44281);
nand U45734 (N_45734,N_44231,N_44950);
nor U45735 (N_45735,N_44083,N_44847);
xor U45736 (N_45736,N_44093,N_44448);
nand U45737 (N_45737,N_44568,N_44533);
xnor U45738 (N_45738,N_44933,N_44071);
and U45739 (N_45739,N_44343,N_44399);
and U45740 (N_45740,N_44383,N_44697);
xnor U45741 (N_45741,N_44490,N_44337);
and U45742 (N_45742,N_44591,N_44399);
xnor U45743 (N_45743,N_44351,N_44519);
nand U45744 (N_45744,N_44019,N_44131);
and U45745 (N_45745,N_44398,N_44958);
nor U45746 (N_45746,N_44048,N_44552);
and U45747 (N_45747,N_44904,N_44129);
and U45748 (N_45748,N_44314,N_44996);
and U45749 (N_45749,N_44229,N_44882);
nor U45750 (N_45750,N_44608,N_44373);
nor U45751 (N_45751,N_44140,N_44643);
xnor U45752 (N_45752,N_44333,N_44808);
nor U45753 (N_45753,N_44404,N_44504);
or U45754 (N_45754,N_44382,N_44925);
or U45755 (N_45755,N_44985,N_44289);
nor U45756 (N_45756,N_44366,N_44696);
or U45757 (N_45757,N_44418,N_44665);
nor U45758 (N_45758,N_44408,N_44634);
or U45759 (N_45759,N_44265,N_44331);
or U45760 (N_45760,N_44878,N_44727);
and U45761 (N_45761,N_44960,N_44058);
or U45762 (N_45762,N_44711,N_44366);
nor U45763 (N_45763,N_44049,N_44645);
xnor U45764 (N_45764,N_44585,N_44355);
or U45765 (N_45765,N_44095,N_44004);
nand U45766 (N_45766,N_44984,N_44760);
and U45767 (N_45767,N_44968,N_44448);
nand U45768 (N_45768,N_44709,N_44530);
and U45769 (N_45769,N_44090,N_44651);
nand U45770 (N_45770,N_44361,N_44305);
nand U45771 (N_45771,N_44484,N_44433);
nor U45772 (N_45772,N_44633,N_44612);
and U45773 (N_45773,N_44974,N_44367);
nand U45774 (N_45774,N_44227,N_44016);
or U45775 (N_45775,N_44166,N_44518);
or U45776 (N_45776,N_44042,N_44947);
xor U45777 (N_45777,N_44023,N_44443);
nor U45778 (N_45778,N_44654,N_44435);
or U45779 (N_45779,N_44775,N_44835);
or U45780 (N_45780,N_44108,N_44051);
nand U45781 (N_45781,N_44930,N_44682);
and U45782 (N_45782,N_44998,N_44262);
nand U45783 (N_45783,N_44269,N_44222);
or U45784 (N_45784,N_44005,N_44291);
or U45785 (N_45785,N_44257,N_44716);
or U45786 (N_45786,N_44290,N_44647);
xor U45787 (N_45787,N_44136,N_44261);
nand U45788 (N_45788,N_44785,N_44431);
nand U45789 (N_45789,N_44735,N_44909);
nand U45790 (N_45790,N_44505,N_44510);
or U45791 (N_45791,N_44708,N_44971);
nor U45792 (N_45792,N_44982,N_44470);
or U45793 (N_45793,N_44387,N_44462);
and U45794 (N_45794,N_44199,N_44338);
nor U45795 (N_45795,N_44667,N_44143);
and U45796 (N_45796,N_44127,N_44329);
nor U45797 (N_45797,N_44200,N_44383);
or U45798 (N_45798,N_44841,N_44324);
nor U45799 (N_45799,N_44204,N_44808);
xor U45800 (N_45800,N_44463,N_44545);
or U45801 (N_45801,N_44959,N_44501);
or U45802 (N_45802,N_44864,N_44814);
or U45803 (N_45803,N_44613,N_44230);
xnor U45804 (N_45804,N_44725,N_44456);
and U45805 (N_45805,N_44994,N_44981);
xnor U45806 (N_45806,N_44072,N_44903);
nor U45807 (N_45807,N_44787,N_44956);
nor U45808 (N_45808,N_44759,N_44111);
or U45809 (N_45809,N_44666,N_44775);
nand U45810 (N_45810,N_44181,N_44378);
and U45811 (N_45811,N_44381,N_44163);
and U45812 (N_45812,N_44858,N_44991);
or U45813 (N_45813,N_44389,N_44744);
xnor U45814 (N_45814,N_44133,N_44350);
or U45815 (N_45815,N_44420,N_44483);
and U45816 (N_45816,N_44079,N_44828);
xor U45817 (N_45817,N_44974,N_44072);
xor U45818 (N_45818,N_44773,N_44591);
nor U45819 (N_45819,N_44533,N_44942);
nor U45820 (N_45820,N_44851,N_44036);
or U45821 (N_45821,N_44397,N_44695);
nand U45822 (N_45822,N_44511,N_44008);
xnor U45823 (N_45823,N_44565,N_44906);
nor U45824 (N_45824,N_44295,N_44009);
or U45825 (N_45825,N_44549,N_44618);
xnor U45826 (N_45826,N_44576,N_44567);
nand U45827 (N_45827,N_44590,N_44013);
and U45828 (N_45828,N_44562,N_44010);
nor U45829 (N_45829,N_44368,N_44318);
nor U45830 (N_45830,N_44889,N_44644);
or U45831 (N_45831,N_44137,N_44374);
or U45832 (N_45832,N_44529,N_44555);
or U45833 (N_45833,N_44545,N_44854);
or U45834 (N_45834,N_44061,N_44339);
or U45835 (N_45835,N_44099,N_44141);
and U45836 (N_45836,N_44674,N_44622);
nor U45837 (N_45837,N_44683,N_44259);
and U45838 (N_45838,N_44127,N_44641);
or U45839 (N_45839,N_44402,N_44057);
xor U45840 (N_45840,N_44054,N_44871);
nor U45841 (N_45841,N_44224,N_44815);
nor U45842 (N_45842,N_44841,N_44881);
or U45843 (N_45843,N_44573,N_44622);
or U45844 (N_45844,N_44183,N_44628);
and U45845 (N_45845,N_44538,N_44861);
and U45846 (N_45846,N_44295,N_44235);
and U45847 (N_45847,N_44559,N_44082);
or U45848 (N_45848,N_44701,N_44030);
and U45849 (N_45849,N_44936,N_44630);
nor U45850 (N_45850,N_44795,N_44065);
and U45851 (N_45851,N_44431,N_44396);
xnor U45852 (N_45852,N_44224,N_44251);
xor U45853 (N_45853,N_44627,N_44289);
xor U45854 (N_45854,N_44001,N_44542);
or U45855 (N_45855,N_44501,N_44595);
nor U45856 (N_45856,N_44090,N_44650);
or U45857 (N_45857,N_44994,N_44775);
nand U45858 (N_45858,N_44340,N_44313);
nor U45859 (N_45859,N_44759,N_44279);
nor U45860 (N_45860,N_44382,N_44200);
and U45861 (N_45861,N_44051,N_44872);
nor U45862 (N_45862,N_44561,N_44788);
and U45863 (N_45863,N_44534,N_44283);
nand U45864 (N_45864,N_44206,N_44395);
and U45865 (N_45865,N_44553,N_44210);
nor U45866 (N_45866,N_44050,N_44834);
xnor U45867 (N_45867,N_44239,N_44820);
and U45868 (N_45868,N_44855,N_44332);
and U45869 (N_45869,N_44491,N_44503);
and U45870 (N_45870,N_44220,N_44118);
xnor U45871 (N_45871,N_44055,N_44277);
xor U45872 (N_45872,N_44657,N_44364);
xnor U45873 (N_45873,N_44701,N_44926);
xor U45874 (N_45874,N_44979,N_44337);
xnor U45875 (N_45875,N_44624,N_44740);
nor U45876 (N_45876,N_44797,N_44573);
or U45877 (N_45877,N_44084,N_44626);
nand U45878 (N_45878,N_44222,N_44162);
nor U45879 (N_45879,N_44026,N_44790);
or U45880 (N_45880,N_44214,N_44586);
and U45881 (N_45881,N_44019,N_44092);
and U45882 (N_45882,N_44602,N_44648);
or U45883 (N_45883,N_44537,N_44777);
or U45884 (N_45884,N_44244,N_44747);
and U45885 (N_45885,N_44731,N_44693);
xnor U45886 (N_45886,N_44886,N_44638);
nand U45887 (N_45887,N_44366,N_44024);
xnor U45888 (N_45888,N_44702,N_44825);
and U45889 (N_45889,N_44337,N_44825);
and U45890 (N_45890,N_44945,N_44511);
and U45891 (N_45891,N_44917,N_44313);
nor U45892 (N_45892,N_44676,N_44198);
nor U45893 (N_45893,N_44798,N_44211);
and U45894 (N_45894,N_44301,N_44525);
nor U45895 (N_45895,N_44949,N_44763);
nand U45896 (N_45896,N_44606,N_44954);
nor U45897 (N_45897,N_44000,N_44857);
and U45898 (N_45898,N_44447,N_44981);
or U45899 (N_45899,N_44455,N_44718);
xor U45900 (N_45900,N_44814,N_44532);
or U45901 (N_45901,N_44559,N_44572);
xor U45902 (N_45902,N_44199,N_44536);
and U45903 (N_45903,N_44166,N_44602);
and U45904 (N_45904,N_44553,N_44902);
xnor U45905 (N_45905,N_44302,N_44462);
or U45906 (N_45906,N_44222,N_44052);
xnor U45907 (N_45907,N_44040,N_44797);
xnor U45908 (N_45908,N_44806,N_44227);
xnor U45909 (N_45909,N_44614,N_44509);
and U45910 (N_45910,N_44283,N_44772);
nand U45911 (N_45911,N_44855,N_44383);
and U45912 (N_45912,N_44208,N_44820);
nand U45913 (N_45913,N_44603,N_44227);
or U45914 (N_45914,N_44145,N_44820);
and U45915 (N_45915,N_44598,N_44407);
nand U45916 (N_45916,N_44474,N_44973);
or U45917 (N_45917,N_44540,N_44228);
or U45918 (N_45918,N_44823,N_44019);
xnor U45919 (N_45919,N_44780,N_44545);
nor U45920 (N_45920,N_44526,N_44508);
nor U45921 (N_45921,N_44765,N_44306);
nor U45922 (N_45922,N_44007,N_44345);
nor U45923 (N_45923,N_44447,N_44139);
and U45924 (N_45924,N_44002,N_44805);
or U45925 (N_45925,N_44890,N_44797);
and U45926 (N_45926,N_44362,N_44369);
nand U45927 (N_45927,N_44299,N_44476);
nor U45928 (N_45928,N_44232,N_44231);
nor U45929 (N_45929,N_44728,N_44353);
and U45930 (N_45930,N_44086,N_44825);
xor U45931 (N_45931,N_44226,N_44587);
or U45932 (N_45932,N_44391,N_44928);
nor U45933 (N_45933,N_44717,N_44817);
or U45934 (N_45934,N_44029,N_44371);
or U45935 (N_45935,N_44873,N_44323);
nor U45936 (N_45936,N_44140,N_44031);
nand U45937 (N_45937,N_44270,N_44415);
or U45938 (N_45938,N_44516,N_44392);
nor U45939 (N_45939,N_44607,N_44846);
nor U45940 (N_45940,N_44541,N_44260);
or U45941 (N_45941,N_44316,N_44913);
nor U45942 (N_45942,N_44182,N_44236);
or U45943 (N_45943,N_44024,N_44331);
xor U45944 (N_45944,N_44552,N_44071);
nand U45945 (N_45945,N_44602,N_44638);
nor U45946 (N_45946,N_44829,N_44515);
and U45947 (N_45947,N_44223,N_44889);
nand U45948 (N_45948,N_44769,N_44773);
xor U45949 (N_45949,N_44133,N_44889);
xor U45950 (N_45950,N_44670,N_44381);
nand U45951 (N_45951,N_44334,N_44278);
and U45952 (N_45952,N_44984,N_44907);
nand U45953 (N_45953,N_44533,N_44758);
nor U45954 (N_45954,N_44786,N_44974);
nand U45955 (N_45955,N_44172,N_44634);
or U45956 (N_45956,N_44041,N_44942);
xor U45957 (N_45957,N_44347,N_44112);
xnor U45958 (N_45958,N_44875,N_44935);
or U45959 (N_45959,N_44085,N_44775);
nand U45960 (N_45960,N_44176,N_44628);
nor U45961 (N_45961,N_44285,N_44693);
xnor U45962 (N_45962,N_44421,N_44029);
and U45963 (N_45963,N_44530,N_44418);
and U45964 (N_45964,N_44432,N_44174);
or U45965 (N_45965,N_44365,N_44360);
xnor U45966 (N_45966,N_44162,N_44735);
or U45967 (N_45967,N_44210,N_44965);
xor U45968 (N_45968,N_44846,N_44593);
nand U45969 (N_45969,N_44833,N_44610);
nand U45970 (N_45970,N_44238,N_44093);
or U45971 (N_45971,N_44232,N_44251);
nand U45972 (N_45972,N_44086,N_44965);
xnor U45973 (N_45973,N_44937,N_44940);
and U45974 (N_45974,N_44904,N_44245);
or U45975 (N_45975,N_44541,N_44025);
nand U45976 (N_45976,N_44328,N_44252);
or U45977 (N_45977,N_44558,N_44605);
nand U45978 (N_45978,N_44633,N_44730);
nor U45979 (N_45979,N_44195,N_44108);
xnor U45980 (N_45980,N_44066,N_44094);
xor U45981 (N_45981,N_44872,N_44357);
and U45982 (N_45982,N_44683,N_44626);
and U45983 (N_45983,N_44637,N_44919);
and U45984 (N_45984,N_44236,N_44478);
nand U45985 (N_45985,N_44509,N_44148);
xnor U45986 (N_45986,N_44415,N_44110);
or U45987 (N_45987,N_44496,N_44332);
and U45988 (N_45988,N_44097,N_44391);
nor U45989 (N_45989,N_44175,N_44670);
and U45990 (N_45990,N_44249,N_44201);
or U45991 (N_45991,N_44842,N_44684);
nor U45992 (N_45992,N_44934,N_44581);
nor U45993 (N_45993,N_44650,N_44404);
nand U45994 (N_45994,N_44217,N_44337);
or U45995 (N_45995,N_44957,N_44248);
or U45996 (N_45996,N_44766,N_44017);
or U45997 (N_45997,N_44266,N_44476);
or U45998 (N_45998,N_44605,N_44659);
nor U45999 (N_45999,N_44087,N_44678);
xnor U46000 (N_46000,N_45969,N_45989);
nor U46001 (N_46001,N_45215,N_45450);
xor U46002 (N_46002,N_45996,N_45231);
nand U46003 (N_46003,N_45785,N_45058);
and U46004 (N_46004,N_45282,N_45073);
or U46005 (N_46005,N_45919,N_45766);
nor U46006 (N_46006,N_45893,N_45788);
and U46007 (N_46007,N_45367,N_45583);
or U46008 (N_46008,N_45471,N_45546);
nor U46009 (N_46009,N_45025,N_45502);
xor U46010 (N_46010,N_45200,N_45030);
or U46011 (N_46011,N_45466,N_45125);
nand U46012 (N_46012,N_45258,N_45596);
xor U46013 (N_46013,N_45250,N_45652);
nand U46014 (N_46014,N_45216,N_45878);
or U46015 (N_46015,N_45089,N_45486);
xnor U46016 (N_46016,N_45889,N_45709);
nor U46017 (N_46017,N_45463,N_45864);
nand U46018 (N_46018,N_45036,N_45808);
and U46019 (N_46019,N_45449,N_45980);
nor U46020 (N_46020,N_45854,N_45422);
and U46021 (N_46021,N_45802,N_45316);
xor U46022 (N_46022,N_45225,N_45409);
nand U46023 (N_46023,N_45222,N_45848);
xor U46024 (N_46024,N_45865,N_45883);
nand U46025 (N_46025,N_45798,N_45845);
and U46026 (N_46026,N_45885,N_45273);
nor U46027 (N_46027,N_45140,N_45941);
xnor U46028 (N_46028,N_45704,N_45375);
or U46029 (N_46029,N_45625,N_45789);
and U46030 (N_46030,N_45850,N_45942);
nand U46031 (N_46031,N_45890,N_45803);
xor U46032 (N_46032,N_45610,N_45142);
nor U46033 (N_46033,N_45742,N_45710);
or U46034 (N_46034,N_45618,N_45204);
nor U46035 (N_46035,N_45696,N_45473);
or U46036 (N_46036,N_45267,N_45272);
nand U46037 (N_46037,N_45485,N_45555);
and U46038 (N_46038,N_45500,N_45038);
and U46039 (N_46039,N_45522,N_45894);
nor U46040 (N_46040,N_45554,N_45100);
and U46041 (N_46041,N_45966,N_45037);
and U46042 (N_46042,N_45619,N_45926);
nor U46043 (N_46043,N_45227,N_45171);
nor U46044 (N_46044,N_45531,N_45237);
nor U46045 (N_46045,N_45192,N_45564);
nand U46046 (N_46046,N_45491,N_45768);
nand U46047 (N_46047,N_45069,N_45925);
nor U46048 (N_46048,N_45039,N_45141);
nand U46049 (N_46049,N_45355,N_45532);
xor U46050 (N_46050,N_45795,N_45573);
nand U46051 (N_46051,N_45791,N_45041);
nor U46052 (N_46052,N_45859,N_45226);
and U46053 (N_46053,N_45081,N_45310);
xor U46054 (N_46054,N_45595,N_45621);
nor U46055 (N_46055,N_45718,N_45332);
xnor U46056 (N_46056,N_45957,N_45689);
and U46057 (N_46057,N_45043,N_45498);
and U46058 (N_46058,N_45642,N_45339);
nor U46059 (N_46059,N_45430,N_45018);
xnor U46060 (N_46060,N_45862,N_45399);
and U46061 (N_46061,N_45390,N_45458);
xnor U46062 (N_46062,N_45602,N_45211);
or U46063 (N_46063,N_45098,N_45732);
nor U46064 (N_46064,N_45270,N_45229);
nor U46065 (N_46065,N_45816,N_45724);
or U46066 (N_46066,N_45976,N_45769);
nand U46067 (N_46067,N_45285,N_45361);
nor U46068 (N_46068,N_45584,N_45138);
nand U46069 (N_46069,N_45074,N_45149);
or U46070 (N_46070,N_45717,N_45353);
or U46071 (N_46071,N_45824,N_45002);
and U46072 (N_46072,N_45708,N_45245);
and U46073 (N_46073,N_45699,N_45161);
and U46074 (N_46074,N_45933,N_45320);
nand U46075 (N_46075,N_45715,N_45374);
nor U46076 (N_46076,N_45494,N_45042);
or U46077 (N_46077,N_45014,N_45992);
nand U46078 (N_46078,N_45951,N_45068);
and U46079 (N_46079,N_45464,N_45291);
xor U46080 (N_46080,N_45369,N_45207);
nand U46081 (N_46081,N_45830,N_45467);
nor U46082 (N_46082,N_45358,N_45947);
nor U46083 (N_46083,N_45840,N_45406);
and U46084 (N_46084,N_45444,N_45421);
and U46085 (N_46085,N_45110,N_45755);
nor U46086 (N_46086,N_45553,N_45213);
xnor U46087 (N_46087,N_45900,N_45566);
nand U46088 (N_46088,N_45576,N_45603);
xnor U46089 (N_46089,N_45266,N_45301);
nand U46090 (N_46090,N_45695,N_45896);
or U46091 (N_46091,N_45462,N_45934);
nor U46092 (N_46092,N_45021,N_45313);
and U46093 (N_46093,N_45080,N_45870);
xnor U46094 (N_46094,N_45626,N_45882);
and U46095 (N_46095,N_45876,N_45295);
xnor U46096 (N_46096,N_45857,N_45283);
nor U46097 (N_46097,N_45106,N_45530);
xnor U46098 (N_46098,N_45087,N_45286);
xor U46099 (N_46099,N_45040,N_45852);
xnor U46100 (N_46100,N_45760,N_45303);
nand U46101 (N_46101,N_45304,N_45033);
nor U46102 (N_46102,N_45815,N_45078);
and U46103 (N_46103,N_45103,N_45912);
nor U46104 (N_46104,N_45688,N_45317);
nand U46105 (N_46105,N_45481,N_45725);
nor U46106 (N_46106,N_45565,N_45509);
or U46107 (N_46107,N_45356,N_45836);
nor U46108 (N_46108,N_45115,N_45235);
or U46109 (N_46109,N_45578,N_45180);
or U46110 (N_46110,N_45257,N_45929);
nand U46111 (N_46111,N_45147,N_45507);
and U46112 (N_46112,N_45646,N_45423);
or U46113 (N_46113,N_45800,N_45370);
and U46114 (N_46114,N_45753,N_45220);
and U46115 (N_46115,N_45210,N_45927);
nor U46116 (N_46116,N_45945,N_45413);
or U46117 (N_46117,N_45524,N_45964);
or U46118 (N_46118,N_45241,N_45178);
xnor U46119 (N_46119,N_45160,N_45681);
xor U46120 (N_46120,N_45453,N_45244);
nor U46121 (N_46121,N_45682,N_45612);
xor U46122 (N_46122,N_45228,N_45672);
nand U46123 (N_46123,N_45337,N_45948);
or U46124 (N_46124,N_45392,N_45117);
nor U46125 (N_46125,N_45813,N_45028);
nand U46126 (N_46126,N_45774,N_45383);
or U46127 (N_46127,N_45787,N_45762);
xnor U46128 (N_46128,N_45045,N_45635);
and U46129 (N_46129,N_45261,N_45977);
xor U46130 (N_46130,N_45661,N_45015);
xor U46131 (N_46131,N_45720,N_45506);
or U46132 (N_46132,N_45129,N_45079);
nor U46133 (N_46133,N_45232,N_45405);
and U46134 (N_46134,N_45656,N_45759);
nor U46135 (N_46135,N_45032,N_45460);
nor U46136 (N_46136,N_45122,N_45575);
nor U46137 (N_46137,N_45671,N_45297);
nand U46138 (N_46138,N_45913,N_45641);
nand U46139 (N_46139,N_45362,N_45159);
nand U46140 (N_46140,N_45535,N_45735);
nor U46141 (N_46141,N_45675,N_45606);
nor U46142 (N_46142,N_45104,N_45658);
and U46143 (N_46143,N_45891,N_45861);
and U46144 (N_46144,N_45806,N_45744);
and U46145 (N_46145,N_45263,N_45842);
nor U46146 (N_46146,N_45404,N_45846);
and U46147 (N_46147,N_45936,N_45090);
xnor U46148 (N_46148,N_45182,N_45468);
and U46149 (N_46149,N_45408,N_45278);
or U46150 (N_46150,N_45561,N_45548);
or U46151 (N_46151,N_45434,N_45959);
or U46152 (N_46152,N_45909,N_45910);
and U46153 (N_46153,N_45252,N_45587);
xor U46154 (N_46154,N_45442,N_45072);
xor U46155 (N_46155,N_45731,N_45132);
or U46156 (N_46156,N_45007,N_45887);
nand U46157 (N_46157,N_45684,N_45938);
or U46158 (N_46158,N_45047,N_45677);
xnor U46159 (N_46159,N_45549,N_45526);
xor U46160 (N_46160,N_45218,N_45930);
xor U46161 (N_46161,N_45607,N_45348);
or U46162 (N_46162,N_45264,N_45116);
and U46163 (N_46163,N_45020,N_45551);
nor U46164 (N_46164,N_45664,N_45590);
nand U46165 (N_46165,N_45853,N_45962);
or U46166 (N_46166,N_45611,N_45822);
and U46167 (N_46167,N_45702,N_45924);
nor U46168 (N_46168,N_45654,N_45991);
and U46169 (N_46169,N_45364,N_45493);
and U46170 (N_46170,N_45224,N_45446);
nand U46171 (N_46171,N_45567,N_45443);
and U46172 (N_46172,N_45761,N_45376);
and U46173 (N_46173,N_45338,N_45749);
xor U46174 (N_46174,N_45819,N_45954);
xor U46175 (N_46175,N_45144,N_45238);
nor U46176 (N_46176,N_45582,N_45403);
xor U46177 (N_46177,N_45624,N_45354);
nor U46178 (N_46178,N_45424,N_45923);
nor U46179 (N_46179,N_45714,N_45503);
and U46180 (N_46180,N_45153,N_45118);
or U46181 (N_46181,N_45428,N_45175);
nor U46182 (N_46182,N_45837,N_45351);
nor U46183 (N_46183,N_45734,N_45740);
or U46184 (N_46184,N_45372,N_45330);
nand U46185 (N_46185,N_45165,N_45647);
or U46186 (N_46186,N_45569,N_45793);
or U46187 (N_46187,N_45064,N_45949);
or U46188 (N_46188,N_45600,N_45345);
xor U46189 (N_46189,N_45637,N_45203);
nand U46190 (N_46190,N_45414,N_45181);
and U46191 (N_46191,N_45308,N_45001);
xor U46192 (N_46192,N_45679,N_45342);
nor U46193 (N_46193,N_45176,N_45209);
nor U46194 (N_46194,N_45169,N_45461);
nand U46195 (N_46195,N_45139,N_45693);
nand U46196 (N_46196,N_45779,N_45031);
or U46197 (N_46197,N_45757,N_45897);
or U46198 (N_46198,N_45311,N_45119);
nand U46199 (N_46199,N_45000,N_45823);
or U46200 (N_46200,N_45197,N_45541);
nand U46201 (N_46201,N_45188,N_45128);
nand U46202 (N_46202,N_45673,N_45643);
nor U46203 (N_46203,N_45478,N_45868);
or U46204 (N_46204,N_45516,N_45721);
xnor U46205 (N_46205,N_45183,N_45052);
and U46206 (N_46206,N_45419,N_45756);
nand U46207 (N_46207,N_45552,N_45628);
xor U46208 (N_46208,N_45236,N_45810);
and U46209 (N_46209,N_45205,N_45177);
xnor U46210 (N_46210,N_45382,N_45917);
or U46211 (N_46211,N_45636,N_45655);
xnor U46212 (N_46212,N_45248,N_45741);
xnor U46213 (N_46213,N_45151,N_45016);
xnor U46214 (N_46214,N_45651,N_45490);
nand U46215 (N_46215,N_45112,N_45847);
xnor U46216 (N_46216,N_45003,N_45605);
or U46217 (N_46217,N_45880,N_45520);
and U46218 (N_46218,N_45821,N_45420);
nor U46219 (N_46219,N_45558,N_45812);
xor U46220 (N_46220,N_45591,N_45136);
nand U46221 (N_46221,N_45008,N_45085);
xnor U46222 (N_46222,N_45747,N_45440);
and U46223 (N_46223,N_45946,N_45508);
or U46224 (N_46224,N_45918,N_45111);
nand U46225 (N_46225,N_45448,N_45315);
nor U46226 (N_46226,N_45006,N_45095);
xor U46227 (N_46227,N_45776,N_45084);
nand U46228 (N_46228,N_45495,N_45748);
xor U46229 (N_46229,N_45196,N_45700);
nor U46230 (N_46230,N_45187,N_45269);
xor U46231 (N_46231,N_45649,N_45726);
or U46232 (N_46232,N_45872,N_45687);
and U46233 (N_46233,N_45055,N_45034);
or U46234 (N_46234,N_45379,N_45035);
nor U46235 (N_46235,N_45307,N_45288);
or U46236 (N_46236,N_45445,N_45432);
nor U46237 (N_46237,N_45814,N_45289);
xnor U46238 (N_46238,N_45046,N_45719);
or U46239 (N_46239,N_45556,N_45557);
nor U46240 (N_46240,N_45324,N_45662);
xnor U46241 (N_46241,N_45519,N_45378);
or U46242 (N_46242,N_45685,N_45214);
and U46243 (N_46243,N_45799,N_45539);
xnor U46244 (N_46244,N_45581,N_45402);
and U46245 (N_46245,N_45166,N_45381);
or U46246 (N_46246,N_45251,N_45154);
or U46247 (N_46247,N_45163,N_45066);
or U46248 (N_46248,N_45497,N_45133);
xor U46249 (N_46249,N_45186,N_45838);
and U46250 (N_46250,N_45427,N_45805);
xnor U46251 (N_46251,N_45426,N_45327);
or U46252 (N_46252,N_45256,N_45212);
or U46253 (N_46253,N_45436,N_45242);
nor U46254 (N_46254,N_45054,N_45185);
nand U46255 (N_46255,N_45780,N_45986);
xnor U46256 (N_46256,N_45952,N_45727);
nor U46257 (N_46257,N_45645,N_45172);
and U46258 (N_46258,N_45091,N_45616);
and U46259 (N_46259,N_45410,N_45869);
xor U46260 (N_46260,N_45255,N_45387);
xor U46261 (N_46261,N_45648,N_45851);
nand U46262 (N_46262,N_45060,N_45781);
xnor U46263 (N_46263,N_45230,N_45908);
or U46264 (N_46264,N_45538,N_45873);
nor U46265 (N_46265,N_45521,N_45730);
and U46266 (N_46266,N_45048,N_45750);
nand U46267 (N_46267,N_45157,N_45431);
nand U46268 (N_46268,N_45331,N_45660);
nor U46269 (N_46269,N_45164,N_45827);
nor U46270 (N_46270,N_45150,N_45886);
or U46271 (N_46271,N_45412,N_45124);
or U46272 (N_46272,N_45825,N_45457);
and U46273 (N_46273,N_45638,N_45683);
and U46274 (N_46274,N_45544,N_45429);
xnor U46275 (N_46275,N_45640,N_45737);
and U46276 (N_46276,N_45973,N_45279);
nand U46277 (N_46277,N_45540,N_45983);
xor U46278 (N_46278,N_45219,N_45371);
nand U46279 (N_46279,N_45614,N_45657);
nand U46280 (N_46280,N_45318,N_45944);
and U46281 (N_46281,N_45574,N_45801);
and U46282 (N_46282,N_45786,N_45899);
nand U46283 (N_46283,N_45504,N_45223);
and U46284 (N_46284,N_45026,N_45298);
xnor U46285 (N_46285,N_45697,N_45170);
or U46286 (N_46286,N_45920,N_45905);
and U46287 (N_46287,N_45928,N_45650);
xor U46288 (N_46288,N_45492,N_45010);
nor U46289 (N_46289,N_45137,N_45009);
nand U46290 (N_46290,N_45243,N_45686);
and U46291 (N_46291,N_45895,N_45995);
xor U46292 (N_46292,N_45189,N_45547);
and U46293 (N_46293,N_45293,N_45208);
or U46294 (N_46294,N_45764,N_45961);
nand U46295 (N_46295,N_45083,N_45765);
and U46296 (N_46296,N_45617,N_45127);
or U46297 (N_46297,N_45592,N_45588);
xor U46298 (N_46298,N_45694,N_45206);
or U46299 (N_46299,N_45004,N_45488);
nor U46300 (N_46300,N_45470,N_45571);
nand U46301 (N_46301,N_45875,N_45901);
nand U46302 (N_46302,N_45593,N_45738);
and U46303 (N_46303,N_45290,N_45322);
xnor U46304 (N_46304,N_45703,N_45334);
or U46305 (N_46305,N_45902,N_45505);
and U46306 (N_46306,N_45300,N_45743);
nor U46307 (N_46307,N_45094,N_45415);
nand U46308 (N_46308,N_45368,N_45314);
xor U46309 (N_46309,N_45701,N_45433);
and U46310 (N_46310,N_45221,N_45400);
nand U46311 (N_46311,N_45134,N_45782);
and U46312 (N_46312,N_45537,N_45644);
nand U46313 (N_46313,N_45347,N_45828);
nand U46314 (N_46314,N_45063,N_45993);
nand U46315 (N_46315,N_45579,N_45965);
or U46316 (N_46316,N_45416,N_45967);
nand U46317 (N_46317,N_45517,N_45296);
nor U46318 (N_46318,N_45712,N_45771);
nand U46319 (N_46319,N_45623,N_45629);
or U46320 (N_46320,N_45148,N_45982);
nand U46321 (N_46321,N_45156,N_45953);
or U46322 (N_46322,N_45086,N_45676);
nor U46323 (N_46323,N_45523,N_45667);
xor U46324 (N_46324,N_45772,N_45723);
or U46325 (N_46325,N_45634,N_45126);
nand U46326 (N_46326,N_45292,N_45550);
and U46327 (N_46327,N_45609,N_45326);
nor U46328 (N_46328,N_45247,N_45811);
or U46329 (N_46329,N_45922,N_45758);
and U46330 (N_46330,N_45968,N_45385);
nand U46331 (N_46331,N_45931,N_45542);
xnor U46332 (N_46332,N_45784,N_45733);
and U46333 (N_46333,N_45305,N_45971);
or U46334 (N_46334,N_45484,N_45455);
nor U46335 (N_46335,N_45287,N_45013);
nand U46336 (N_46336,N_45678,N_45056);
xor U46337 (N_46337,N_45259,N_45511);
xor U46338 (N_46338,N_45023,N_45572);
nor U46339 (N_46339,N_45174,N_45262);
xnor U46340 (N_46340,N_45198,N_45114);
nor U46341 (N_46341,N_45994,N_45601);
or U46342 (N_46342,N_45254,N_45829);
nor U46343 (N_46343,N_45341,N_45082);
nor U46344 (N_46344,N_45459,N_45067);
or U46345 (N_46345,N_45594,N_45359);
xor U46346 (N_46346,N_45745,N_45386);
xor U46347 (N_46347,N_45158,N_45670);
xnor U46348 (N_46348,N_45577,N_45630);
or U46349 (N_46349,N_45570,N_45184);
or U46350 (N_46350,N_45411,N_45998);
or U46351 (N_46351,N_45906,N_45975);
and U46352 (N_46352,N_45866,N_45510);
and U46353 (N_46353,N_45194,N_45487);
and U46354 (N_46354,N_45005,N_45604);
nand U46355 (N_46355,N_45131,N_45560);
and U46356 (N_46356,N_45022,N_45050);
nand U46357 (N_46357,N_45044,N_45956);
xnor U46358 (N_46358,N_45077,N_45352);
xnor U46359 (N_46359,N_45987,N_45146);
xor U46360 (N_46360,N_45775,N_45997);
xnor U46361 (N_46361,N_45281,N_45527);
and U46362 (N_46362,N_45767,N_45482);
nand U46363 (N_46363,N_45792,N_45479);
or U46364 (N_46364,N_45346,N_45395);
and U46365 (N_46365,N_45391,N_45384);
nor U46366 (N_46366,N_45988,N_45397);
nor U46367 (N_46367,N_45388,N_45807);
xnor U46368 (N_46368,N_45284,N_45666);
and U46369 (N_46369,N_45984,N_45613);
nor U46370 (N_46370,N_45191,N_45012);
xor U46371 (N_46371,N_45937,N_45729);
nand U46372 (N_46372,N_45120,N_45716);
nand U46373 (N_46373,N_45820,N_45168);
and U46374 (N_46374,N_45107,N_45620);
and U46375 (N_46375,N_45974,N_45017);
xnor U46376 (N_46376,N_45525,N_45465);
xor U46377 (N_46377,N_45328,N_45143);
or U46378 (N_46378,N_45585,N_45474);
nand U46379 (N_46379,N_45075,N_45407);
nand U46380 (N_46380,N_45960,N_45349);
xnor U46381 (N_46381,N_45329,N_45751);
and U46382 (N_46382,N_45597,N_45877);
or U46383 (N_46383,N_45691,N_45451);
nor U46384 (N_46384,N_45309,N_45323);
nand U46385 (N_46385,N_45253,N_45518);
or U46386 (N_46386,N_45179,N_45778);
and U46387 (N_46387,N_45668,N_45489);
nand U46388 (N_46388,N_45543,N_45804);
or U46389 (N_46389,N_45477,N_45841);
nand U46390 (N_46390,N_45860,N_45135);
or U46391 (N_46391,N_45515,N_45871);
nand U46392 (N_46392,N_45070,N_45631);
or U46393 (N_46393,N_45271,N_45325);
xnor U46394 (N_46394,N_45108,N_45162);
and U46395 (N_46395,N_45915,N_45916);
xnor U46396 (N_46396,N_45855,N_45340);
xor U46397 (N_46397,N_45622,N_45884);
nor U46398 (N_46398,N_45109,N_45053);
nand U46399 (N_46399,N_45790,N_45783);
or U46400 (N_46400,N_45881,N_45336);
and U46401 (N_46401,N_45447,N_45739);
nand U46402 (N_46402,N_45155,N_45061);
or U46403 (N_46403,N_45469,N_45389);
and U46404 (N_46404,N_45746,N_45377);
and U46405 (N_46405,N_45728,N_45277);
or U46406 (N_46406,N_45999,N_45190);
nor U46407 (N_46407,N_45011,N_45568);
and U46408 (N_46408,N_45113,N_45483);
nand U46409 (N_46409,N_45480,N_45863);
nand U46410 (N_46410,N_45580,N_45380);
or U46411 (N_46411,N_45195,N_45396);
xnor U46412 (N_46412,N_45514,N_45797);
xor U46413 (N_46413,N_45059,N_45586);
and U46414 (N_46414,N_45663,N_45598);
xor U46415 (N_46415,N_45076,N_45393);
nand U46416 (N_46416,N_45456,N_45268);
xor U46417 (N_46417,N_45401,N_45921);
and U46418 (N_46418,N_45972,N_45680);
nand U46419 (N_46419,N_45722,N_45335);
nor U46420 (N_46420,N_45249,N_45888);
or U46421 (N_46421,N_45096,N_45319);
nor U46422 (N_46422,N_45898,N_45990);
or U46423 (N_46423,N_45705,N_45599);
nand U46424 (N_46424,N_45935,N_45849);
and U46425 (N_46425,N_45659,N_45476);
or U46426 (N_46426,N_45152,N_45763);
nand U46427 (N_46427,N_45911,N_45425);
nand U46428 (N_46428,N_45102,N_45513);
xor U46429 (N_46429,N_45167,N_45713);
nor U46430 (N_46430,N_45499,N_45496);
or U46431 (N_46431,N_45692,N_45123);
nor U46432 (N_46432,N_45394,N_45698);
nor U46433 (N_46433,N_45832,N_45418);
nor U46434 (N_46434,N_45233,N_45333);
nand U46435 (N_46435,N_45101,N_45843);
xor U46436 (N_46436,N_45097,N_45438);
xnor U46437 (N_46437,N_45559,N_45690);
xor U46438 (N_46438,N_45280,N_45536);
xnor U46439 (N_46439,N_45653,N_45130);
nand U46440 (N_46440,N_45265,N_45970);
nand U46441 (N_46441,N_45019,N_45939);
nor U46442 (N_46442,N_45958,N_45512);
or U46443 (N_46443,N_45796,N_45439);
nand U46444 (N_46444,N_45940,N_45202);
nand U46445 (N_46445,N_45357,N_45441);
nor U46446 (N_46446,N_45193,N_45302);
xnor U46447 (N_46447,N_45665,N_45057);
nand U46448 (N_46448,N_45024,N_45027);
nor U46449 (N_46449,N_45563,N_45321);
and U46450 (N_46450,N_45344,N_45274);
or U46451 (N_46451,N_45306,N_45246);
nor U46452 (N_46452,N_45834,N_45817);
nor U46453 (N_46453,N_45343,N_45363);
or U46454 (N_46454,N_45844,N_45299);
or U46455 (N_46455,N_45145,N_45093);
nand U46456 (N_46456,N_45528,N_45029);
and U46457 (N_46457,N_45475,N_45562);
xor U46458 (N_46458,N_45833,N_45099);
nor U46459 (N_46459,N_45932,N_45534);
nand U46460 (N_46460,N_45809,N_45435);
xnor U46461 (N_46461,N_45217,N_45201);
or U46462 (N_46462,N_45173,N_45831);
xnor U46463 (N_46463,N_45879,N_45979);
and U46464 (N_46464,N_45674,N_45417);
and U46465 (N_46465,N_45955,N_45234);
or U46466 (N_46466,N_45049,N_45065);
or U46467 (N_46467,N_45062,N_45312);
xor U46468 (N_46468,N_45950,N_45366);
nand U46469 (N_46469,N_45350,N_45589);
or U46470 (N_46470,N_45501,N_45963);
nor U46471 (N_46471,N_45892,N_45639);
nor U46472 (N_46472,N_45874,N_45706);
and U46473 (N_46473,N_45633,N_45903);
nor U46474 (N_46474,N_45051,N_45545);
nand U46475 (N_46475,N_45533,N_45105);
xnor U46476 (N_46476,N_45529,N_45121);
and U46477 (N_46477,N_45373,N_45632);
xnor U46478 (N_46478,N_45707,N_45839);
nor U46479 (N_46479,N_45669,N_45736);
and U46480 (N_46480,N_45627,N_45835);
nor U46481 (N_46481,N_45452,N_45907);
nor U46482 (N_46482,N_45826,N_45276);
or U46483 (N_46483,N_45240,N_45856);
xnor U46484 (N_46484,N_45275,N_45472);
nand U46485 (N_46485,N_45360,N_45773);
nor U46486 (N_46486,N_45092,N_45260);
or U46487 (N_46487,N_45454,N_45858);
nand U46488 (N_46488,N_45754,N_45777);
and U46489 (N_46489,N_45365,N_45294);
and U46490 (N_46490,N_45398,N_45711);
xor U46491 (N_46491,N_45752,N_45437);
nand U46492 (N_46492,N_45978,N_45199);
nand U46493 (N_46493,N_45943,N_45615);
or U46494 (N_46494,N_45818,N_45794);
xnor U46495 (N_46495,N_45914,N_45981);
nand U46496 (N_46496,N_45904,N_45867);
and U46497 (N_46497,N_45770,N_45985);
nor U46498 (N_46498,N_45608,N_45071);
nor U46499 (N_46499,N_45239,N_45088);
or U46500 (N_46500,N_45412,N_45634);
nand U46501 (N_46501,N_45896,N_45519);
and U46502 (N_46502,N_45379,N_45061);
nor U46503 (N_46503,N_45501,N_45225);
xnor U46504 (N_46504,N_45221,N_45285);
and U46505 (N_46505,N_45245,N_45228);
nor U46506 (N_46506,N_45280,N_45930);
or U46507 (N_46507,N_45361,N_45546);
xnor U46508 (N_46508,N_45852,N_45210);
or U46509 (N_46509,N_45082,N_45632);
nor U46510 (N_46510,N_45910,N_45103);
xor U46511 (N_46511,N_45160,N_45246);
nor U46512 (N_46512,N_45119,N_45989);
or U46513 (N_46513,N_45404,N_45462);
nor U46514 (N_46514,N_45615,N_45175);
nand U46515 (N_46515,N_45692,N_45275);
and U46516 (N_46516,N_45413,N_45006);
and U46517 (N_46517,N_45233,N_45946);
or U46518 (N_46518,N_45206,N_45279);
and U46519 (N_46519,N_45032,N_45339);
xor U46520 (N_46520,N_45820,N_45545);
or U46521 (N_46521,N_45070,N_45422);
nand U46522 (N_46522,N_45725,N_45620);
xor U46523 (N_46523,N_45944,N_45077);
nor U46524 (N_46524,N_45402,N_45842);
or U46525 (N_46525,N_45264,N_45872);
and U46526 (N_46526,N_45027,N_45815);
and U46527 (N_46527,N_45332,N_45466);
or U46528 (N_46528,N_45092,N_45111);
and U46529 (N_46529,N_45625,N_45682);
or U46530 (N_46530,N_45802,N_45002);
or U46531 (N_46531,N_45155,N_45304);
xnor U46532 (N_46532,N_45179,N_45758);
nand U46533 (N_46533,N_45244,N_45193);
nor U46534 (N_46534,N_45193,N_45761);
nor U46535 (N_46535,N_45785,N_45492);
or U46536 (N_46536,N_45046,N_45595);
nand U46537 (N_46537,N_45110,N_45626);
nand U46538 (N_46538,N_45658,N_45574);
nor U46539 (N_46539,N_45376,N_45457);
nand U46540 (N_46540,N_45797,N_45112);
or U46541 (N_46541,N_45047,N_45676);
or U46542 (N_46542,N_45030,N_45369);
and U46543 (N_46543,N_45866,N_45558);
or U46544 (N_46544,N_45832,N_45254);
xor U46545 (N_46545,N_45069,N_45027);
xor U46546 (N_46546,N_45980,N_45907);
nor U46547 (N_46547,N_45924,N_45662);
and U46548 (N_46548,N_45504,N_45164);
nand U46549 (N_46549,N_45302,N_45624);
and U46550 (N_46550,N_45487,N_45557);
xor U46551 (N_46551,N_45253,N_45997);
and U46552 (N_46552,N_45936,N_45347);
or U46553 (N_46553,N_45835,N_45759);
or U46554 (N_46554,N_45691,N_45227);
nor U46555 (N_46555,N_45144,N_45765);
nand U46556 (N_46556,N_45715,N_45961);
nor U46557 (N_46557,N_45505,N_45108);
xnor U46558 (N_46558,N_45649,N_45611);
xnor U46559 (N_46559,N_45856,N_45510);
or U46560 (N_46560,N_45152,N_45510);
or U46561 (N_46561,N_45679,N_45035);
and U46562 (N_46562,N_45008,N_45694);
nand U46563 (N_46563,N_45464,N_45204);
or U46564 (N_46564,N_45197,N_45262);
nand U46565 (N_46565,N_45391,N_45033);
nand U46566 (N_46566,N_45906,N_45220);
nand U46567 (N_46567,N_45841,N_45206);
nor U46568 (N_46568,N_45847,N_45433);
nand U46569 (N_46569,N_45153,N_45324);
nand U46570 (N_46570,N_45276,N_45043);
nor U46571 (N_46571,N_45503,N_45057);
xor U46572 (N_46572,N_45944,N_45759);
nor U46573 (N_46573,N_45401,N_45707);
nor U46574 (N_46574,N_45981,N_45246);
nor U46575 (N_46575,N_45471,N_45515);
and U46576 (N_46576,N_45967,N_45214);
nor U46577 (N_46577,N_45980,N_45048);
or U46578 (N_46578,N_45745,N_45678);
xor U46579 (N_46579,N_45821,N_45750);
nand U46580 (N_46580,N_45561,N_45856);
nand U46581 (N_46581,N_45279,N_45800);
nand U46582 (N_46582,N_45627,N_45513);
or U46583 (N_46583,N_45719,N_45377);
xnor U46584 (N_46584,N_45414,N_45077);
or U46585 (N_46585,N_45584,N_45250);
and U46586 (N_46586,N_45775,N_45126);
nor U46587 (N_46587,N_45192,N_45561);
and U46588 (N_46588,N_45165,N_45576);
or U46589 (N_46589,N_45247,N_45375);
nor U46590 (N_46590,N_45705,N_45501);
xor U46591 (N_46591,N_45117,N_45087);
xnor U46592 (N_46592,N_45051,N_45400);
xnor U46593 (N_46593,N_45457,N_45337);
nand U46594 (N_46594,N_45217,N_45906);
nor U46595 (N_46595,N_45968,N_45267);
xor U46596 (N_46596,N_45272,N_45979);
or U46597 (N_46597,N_45052,N_45454);
or U46598 (N_46598,N_45028,N_45239);
xor U46599 (N_46599,N_45121,N_45253);
xnor U46600 (N_46600,N_45818,N_45018);
xor U46601 (N_46601,N_45508,N_45828);
nor U46602 (N_46602,N_45578,N_45163);
xor U46603 (N_46603,N_45206,N_45731);
or U46604 (N_46604,N_45399,N_45583);
xor U46605 (N_46605,N_45935,N_45193);
and U46606 (N_46606,N_45341,N_45651);
nor U46607 (N_46607,N_45482,N_45504);
or U46608 (N_46608,N_45389,N_45582);
nor U46609 (N_46609,N_45111,N_45657);
and U46610 (N_46610,N_45405,N_45098);
and U46611 (N_46611,N_45822,N_45620);
or U46612 (N_46612,N_45807,N_45819);
and U46613 (N_46613,N_45762,N_45810);
or U46614 (N_46614,N_45083,N_45610);
or U46615 (N_46615,N_45369,N_45611);
or U46616 (N_46616,N_45411,N_45437);
or U46617 (N_46617,N_45391,N_45439);
and U46618 (N_46618,N_45521,N_45135);
nand U46619 (N_46619,N_45847,N_45482);
nand U46620 (N_46620,N_45838,N_45137);
nand U46621 (N_46621,N_45947,N_45696);
xor U46622 (N_46622,N_45756,N_45042);
nand U46623 (N_46623,N_45140,N_45726);
and U46624 (N_46624,N_45830,N_45455);
nand U46625 (N_46625,N_45990,N_45421);
or U46626 (N_46626,N_45724,N_45829);
nand U46627 (N_46627,N_45943,N_45749);
nand U46628 (N_46628,N_45351,N_45518);
xnor U46629 (N_46629,N_45371,N_45363);
and U46630 (N_46630,N_45099,N_45251);
or U46631 (N_46631,N_45718,N_45874);
or U46632 (N_46632,N_45822,N_45158);
nand U46633 (N_46633,N_45023,N_45108);
xnor U46634 (N_46634,N_45978,N_45029);
nand U46635 (N_46635,N_45500,N_45030);
and U46636 (N_46636,N_45755,N_45298);
or U46637 (N_46637,N_45778,N_45163);
nand U46638 (N_46638,N_45056,N_45865);
nand U46639 (N_46639,N_45004,N_45218);
or U46640 (N_46640,N_45899,N_45089);
nor U46641 (N_46641,N_45788,N_45845);
or U46642 (N_46642,N_45198,N_45972);
and U46643 (N_46643,N_45691,N_45580);
and U46644 (N_46644,N_45274,N_45891);
nand U46645 (N_46645,N_45042,N_45014);
nor U46646 (N_46646,N_45462,N_45581);
xor U46647 (N_46647,N_45370,N_45881);
nand U46648 (N_46648,N_45341,N_45068);
xnor U46649 (N_46649,N_45784,N_45457);
nor U46650 (N_46650,N_45918,N_45839);
nand U46651 (N_46651,N_45838,N_45821);
xor U46652 (N_46652,N_45233,N_45711);
nor U46653 (N_46653,N_45221,N_45484);
or U46654 (N_46654,N_45825,N_45689);
nand U46655 (N_46655,N_45271,N_45390);
nor U46656 (N_46656,N_45765,N_45136);
xnor U46657 (N_46657,N_45552,N_45009);
xnor U46658 (N_46658,N_45465,N_45404);
or U46659 (N_46659,N_45339,N_45073);
nand U46660 (N_46660,N_45835,N_45245);
xnor U46661 (N_46661,N_45522,N_45841);
xnor U46662 (N_46662,N_45944,N_45549);
and U46663 (N_46663,N_45689,N_45322);
xnor U46664 (N_46664,N_45955,N_45880);
and U46665 (N_46665,N_45791,N_45623);
and U46666 (N_46666,N_45477,N_45832);
xnor U46667 (N_46667,N_45458,N_45082);
or U46668 (N_46668,N_45476,N_45579);
or U46669 (N_46669,N_45193,N_45933);
nor U46670 (N_46670,N_45177,N_45173);
nand U46671 (N_46671,N_45503,N_45974);
nand U46672 (N_46672,N_45264,N_45196);
or U46673 (N_46673,N_45566,N_45752);
xor U46674 (N_46674,N_45765,N_45041);
nand U46675 (N_46675,N_45380,N_45996);
nor U46676 (N_46676,N_45838,N_45153);
nor U46677 (N_46677,N_45347,N_45228);
xor U46678 (N_46678,N_45216,N_45053);
nor U46679 (N_46679,N_45442,N_45755);
nand U46680 (N_46680,N_45001,N_45200);
nand U46681 (N_46681,N_45296,N_45388);
nor U46682 (N_46682,N_45050,N_45997);
nor U46683 (N_46683,N_45155,N_45669);
and U46684 (N_46684,N_45036,N_45381);
and U46685 (N_46685,N_45841,N_45405);
or U46686 (N_46686,N_45429,N_45186);
xor U46687 (N_46687,N_45905,N_45706);
xnor U46688 (N_46688,N_45428,N_45659);
and U46689 (N_46689,N_45281,N_45224);
or U46690 (N_46690,N_45493,N_45494);
xnor U46691 (N_46691,N_45638,N_45455);
xnor U46692 (N_46692,N_45330,N_45498);
or U46693 (N_46693,N_45390,N_45793);
or U46694 (N_46694,N_45774,N_45084);
nor U46695 (N_46695,N_45426,N_45191);
nor U46696 (N_46696,N_45715,N_45769);
xor U46697 (N_46697,N_45737,N_45278);
or U46698 (N_46698,N_45398,N_45164);
nand U46699 (N_46699,N_45700,N_45432);
xnor U46700 (N_46700,N_45670,N_45804);
and U46701 (N_46701,N_45306,N_45582);
or U46702 (N_46702,N_45901,N_45574);
and U46703 (N_46703,N_45253,N_45251);
and U46704 (N_46704,N_45749,N_45174);
xor U46705 (N_46705,N_45471,N_45054);
or U46706 (N_46706,N_45817,N_45135);
xnor U46707 (N_46707,N_45088,N_45280);
and U46708 (N_46708,N_45921,N_45770);
nand U46709 (N_46709,N_45785,N_45003);
and U46710 (N_46710,N_45598,N_45254);
and U46711 (N_46711,N_45421,N_45300);
nand U46712 (N_46712,N_45383,N_45854);
nor U46713 (N_46713,N_45226,N_45694);
nand U46714 (N_46714,N_45208,N_45131);
nor U46715 (N_46715,N_45464,N_45349);
or U46716 (N_46716,N_45368,N_45462);
and U46717 (N_46717,N_45823,N_45659);
nor U46718 (N_46718,N_45271,N_45590);
nor U46719 (N_46719,N_45574,N_45609);
xnor U46720 (N_46720,N_45098,N_45723);
nor U46721 (N_46721,N_45260,N_45209);
and U46722 (N_46722,N_45282,N_45936);
and U46723 (N_46723,N_45372,N_45804);
nand U46724 (N_46724,N_45430,N_45977);
nand U46725 (N_46725,N_45174,N_45464);
and U46726 (N_46726,N_45034,N_45080);
or U46727 (N_46727,N_45045,N_45599);
nand U46728 (N_46728,N_45305,N_45747);
nor U46729 (N_46729,N_45057,N_45595);
nand U46730 (N_46730,N_45906,N_45115);
nand U46731 (N_46731,N_45612,N_45158);
nor U46732 (N_46732,N_45318,N_45040);
nor U46733 (N_46733,N_45643,N_45731);
xnor U46734 (N_46734,N_45183,N_45955);
nor U46735 (N_46735,N_45353,N_45867);
or U46736 (N_46736,N_45046,N_45090);
and U46737 (N_46737,N_45538,N_45595);
and U46738 (N_46738,N_45032,N_45480);
and U46739 (N_46739,N_45551,N_45768);
nor U46740 (N_46740,N_45503,N_45125);
nand U46741 (N_46741,N_45425,N_45233);
and U46742 (N_46742,N_45877,N_45372);
xor U46743 (N_46743,N_45167,N_45697);
nor U46744 (N_46744,N_45761,N_45826);
nor U46745 (N_46745,N_45313,N_45876);
nand U46746 (N_46746,N_45879,N_45880);
and U46747 (N_46747,N_45941,N_45322);
and U46748 (N_46748,N_45013,N_45747);
xor U46749 (N_46749,N_45091,N_45341);
nor U46750 (N_46750,N_45148,N_45939);
nor U46751 (N_46751,N_45827,N_45319);
and U46752 (N_46752,N_45106,N_45582);
nor U46753 (N_46753,N_45799,N_45056);
nand U46754 (N_46754,N_45538,N_45266);
nor U46755 (N_46755,N_45022,N_45660);
and U46756 (N_46756,N_45349,N_45766);
nor U46757 (N_46757,N_45001,N_45735);
nand U46758 (N_46758,N_45399,N_45892);
nand U46759 (N_46759,N_45499,N_45284);
or U46760 (N_46760,N_45811,N_45901);
nor U46761 (N_46761,N_45473,N_45337);
or U46762 (N_46762,N_45656,N_45498);
or U46763 (N_46763,N_45301,N_45750);
and U46764 (N_46764,N_45641,N_45759);
nand U46765 (N_46765,N_45792,N_45075);
or U46766 (N_46766,N_45108,N_45038);
or U46767 (N_46767,N_45820,N_45031);
xor U46768 (N_46768,N_45130,N_45198);
xnor U46769 (N_46769,N_45360,N_45735);
or U46770 (N_46770,N_45423,N_45323);
nand U46771 (N_46771,N_45052,N_45702);
or U46772 (N_46772,N_45997,N_45452);
and U46773 (N_46773,N_45388,N_45757);
xnor U46774 (N_46774,N_45912,N_45300);
xor U46775 (N_46775,N_45143,N_45924);
and U46776 (N_46776,N_45783,N_45139);
nand U46777 (N_46777,N_45503,N_45323);
and U46778 (N_46778,N_45357,N_45253);
nand U46779 (N_46779,N_45674,N_45686);
or U46780 (N_46780,N_45752,N_45303);
xnor U46781 (N_46781,N_45397,N_45722);
xor U46782 (N_46782,N_45602,N_45449);
xnor U46783 (N_46783,N_45127,N_45745);
xor U46784 (N_46784,N_45237,N_45446);
and U46785 (N_46785,N_45270,N_45141);
nor U46786 (N_46786,N_45007,N_45148);
nand U46787 (N_46787,N_45737,N_45503);
and U46788 (N_46788,N_45114,N_45558);
and U46789 (N_46789,N_45648,N_45528);
nor U46790 (N_46790,N_45463,N_45196);
nor U46791 (N_46791,N_45065,N_45414);
or U46792 (N_46792,N_45089,N_45418);
or U46793 (N_46793,N_45723,N_45113);
nand U46794 (N_46794,N_45263,N_45150);
nor U46795 (N_46795,N_45777,N_45544);
or U46796 (N_46796,N_45936,N_45875);
and U46797 (N_46797,N_45433,N_45616);
nand U46798 (N_46798,N_45656,N_45348);
nor U46799 (N_46799,N_45312,N_45837);
nor U46800 (N_46800,N_45126,N_45469);
or U46801 (N_46801,N_45682,N_45867);
and U46802 (N_46802,N_45047,N_45790);
nand U46803 (N_46803,N_45474,N_45840);
nor U46804 (N_46804,N_45228,N_45580);
nor U46805 (N_46805,N_45817,N_45160);
xnor U46806 (N_46806,N_45621,N_45267);
nor U46807 (N_46807,N_45671,N_45448);
and U46808 (N_46808,N_45415,N_45029);
or U46809 (N_46809,N_45286,N_45472);
and U46810 (N_46810,N_45547,N_45676);
nand U46811 (N_46811,N_45076,N_45022);
nor U46812 (N_46812,N_45200,N_45248);
and U46813 (N_46813,N_45936,N_45011);
xnor U46814 (N_46814,N_45931,N_45509);
nand U46815 (N_46815,N_45712,N_45696);
nor U46816 (N_46816,N_45203,N_45328);
xnor U46817 (N_46817,N_45779,N_45476);
nand U46818 (N_46818,N_45100,N_45885);
nor U46819 (N_46819,N_45766,N_45690);
nor U46820 (N_46820,N_45304,N_45416);
nor U46821 (N_46821,N_45040,N_45966);
xor U46822 (N_46822,N_45877,N_45270);
nand U46823 (N_46823,N_45928,N_45707);
and U46824 (N_46824,N_45695,N_45152);
xor U46825 (N_46825,N_45318,N_45977);
nor U46826 (N_46826,N_45323,N_45813);
nand U46827 (N_46827,N_45947,N_45034);
nor U46828 (N_46828,N_45442,N_45450);
nor U46829 (N_46829,N_45765,N_45112);
xnor U46830 (N_46830,N_45678,N_45467);
or U46831 (N_46831,N_45332,N_45183);
xor U46832 (N_46832,N_45294,N_45100);
xor U46833 (N_46833,N_45476,N_45230);
and U46834 (N_46834,N_45153,N_45411);
or U46835 (N_46835,N_45527,N_45471);
nand U46836 (N_46836,N_45079,N_45820);
and U46837 (N_46837,N_45720,N_45341);
nor U46838 (N_46838,N_45173,N_45987);
xor U46839 (N_46839,N_45806,N_45704);
or U46840 (N_46840,N_45353,N_45015);
or U46841 (N_46841,N_45390,N_45123);
nor U46842 (N_46842,N_45043,N_45900);
or U46843 (N_46843,N_45429,N_45869);
nor U46844 (N_46844,N_45461,N_45358);
nor U46845 (N_46845,N_45658,N_45291);
or U46846 (N_46846,N_45095,N_45951);
nor U46847 (N_46847,N_45990,N_45999);
nor U46848 (N_46848,N_45269,N_45765);
nor U46849 (N_46849,N_45032,N_45313);
xor U46850 (N_46850,N_45984,N_45722);
nand U46851 (N_46851,N_45669,N_45881);
xor U46852 (N_46852,N_45534,N_45118);
nor U46853 (N_46853,N_45616,N_45620);
or U46854 (N_46854,N_45416,N_45984);
nand U46855 (N_46855,N_45136,N_45421);
or U46856 (N_46856,N_45196,N_45928);
and U46857 (N_46857,N_45652,N_45858);
and U46858 (N_46858,N_45276,N_45204);
nand U46859 (N_46859,N_45187,N_45553);
or U46860 (N_46860,N_45204,N_45069);
and U46861 (N_46861,N_45947,N_45280);
xor U46862 (N_46862,N_45850,N_45252);
nor U46863 (N_46863,N_45174,N_45774);
and U46864 (N_46864,N_45939,N_45132);
or U46865 (N_46865,N_45452,N_45095);
or U46866 (N_46866,N_45128,N_45336);
xnor U46867 (N_46867,N_45857,N_45032);
xor U46868 (N_46868,N_45125,N_45948);
and U46869 (N_46869,N_45181,N_45887);
nor U46870 (N_46870,N_45750,N_45508);
nand U46871 (N_46871,N_45344,N_45396);
xor U46872 (N_46872,N_45143,N_45691);
xor U46873 (N_46873,N_45731,N_45279);
nor U46874 (N_46874,N_45330,N_45507);
xnor U46875 (N_46875,N_45414,N_45236);
and U46876 (N_46876,N_45812,N_45259);
and U46877 (N_46877,N_45500,N_45166);
nand U46878 (N_46878,N_45892,N_45073);
xor U46879 (N_46879,N_45403,N_45964);
nand U46880 (N_46880,N_45121,N_45655);
and U46881 (N_46881,N_45127,N_45536);
or U46882 (N_46882,N_45038,N_45909);
and U46883 (N_46883,N_45456,N_45567);
nor U46884 (N_46884,N_45428,N_45004);
nand U46885 (N_46885,N_45838,N_45478);
nor U46886 (N_46886,N_45543,N_45441);
xor U46887 (N_46887,N_45608,N_45787);
and U46888 (N_46888,N_45405,N_45819);
and U46889 (N_46889,N_45520,N_45888);
nand U46890 (N_46890,N_45676,N_45046);
or U46891 (N_46891,N_45552,N_45689);
xnor U46892 (N_46892,N_45489,N_45861);
nor U46893 (N_46893,N_45968,N_45511);
xor U46894 (N_46894,N_45066,N_45660);
nand U46895 (N_46895,N_45121,N_45786);
xnor U46896 (N_46896,N_45923,N_45838);
and U46897 (N_46897,N_45143,N_45042);
and U46898 (N_46898,N_45215,N_45894);
or U46899 (N_46899,N_45358,N_45056);
nor U46900 (N_46900,N_45929,N_45268);
xnor U46901 (N_46901,N_45566,N_45535);
xor U46902 (N_46902,N_45666,N_45313);
xnor U46903 (N_46903,N_45869,N_45639);
or U46904 (N_46904,N_45668,N_45393);
nor U46905 (N_46905,N_45743,N_45706);
nor U46906 (N_46906,N_45866,N_45808);
xor U46907 (N_46907,N_45036,N_45880);
nor U46908 (N_46908,N_45803,N_45952);
xnor U46909 (N_46909,N_45701,N_45847);
and U46910 (N_46910,N_45381,N_45316);
nor U46911 (N_46911,N_45471,N_45311);
nor U46912 (N_46912,N_45496,N_45215);
or U46913 (N_46913,N_45920,N_45890);
nand U46914 (N_46914,N_45173,N_45794);
nand U46915 (N_46915,N_45900,N_45314);
xnor U46916 (N_46916,N_45429,N_45709);
and U46917 (N_46917,N_45535,N_45687);
nand U46918 (N_46918,N_45908,N_45195);
and U46919 (N_46919,N_45105,N_45692);
nor U46920 (N_46920,N_45299,N_45183);
nor U46921 (N_46921,N_45664,N_45489);
nor U46922 (N_46922,N_45138,N_45990);
nand U46923 (N_46923,N_45260,N_45047);
nor U46924 (N_46924,N_45643,N_45678);
xnor U46925 (N_46925,N_45355,N_45705);
nand U46926 (N_46926,N_45957,N_45686);
nor U46927 (N_46927,N_45744,N_45306);
nor U46928 (N_46928,N_45442,N_45407);
nand U46929 (N_46929,N_45247,N_45109);
nand U46930 (N_46930,N_45086,N_45654);
xor U46931 (N_46931,N_45370,N_45640);
nor U46932 (N_46932,N_45732,N_45798);
nor U46933 (N_46933,N_45488,N_45029);
or U46934 (N_46934,N_45606,N_45105);
xor U46935 (N_46935,N_45187,N_45570);
nor U46936 (N_46936,N_45198,N_45086);
or U46937 (N_46937,N_45231,N_45565);
nor U46938 (N_46938,N_45634,N_45733);
nor U46939 (N_46939,N_45511,N_45232);
nand U46940 (N_46940,N_45206,N_45761);
or U46941 (N_46941,N_45329,N_45996);
nor U46942 (N_46942,N_45418,N_45445);
nor U46943 (N_46943,N_45431,N_45464);
nor U46944 (N_46944,N_45577,N_45201);
nor U46945 (N_46945,N_45553,N_45026);
nand U46946 (N_46946,N_45021,N_45030);
nor U46947 (N_46947,N_45506,N_45560);
nor U46948 (N_46948,N_45524,N_45808);
and U46949 (N_46949,N_45229,N_45629);
xor U46950 (N_46950,N_45583,N_45416);
and U46951 (N_46951,N_45142,N_45982);
xnor U46952 (N_46952,N_45389,N_45329);
nor U46953 (N_46953,N_45515,N_45299);
nand U46954 (N_46954,N_45260,N_45448);
nor U46955 (N_46955,N_45985,N_45992);
nor U46956 (N_46956,N_45086,N_45494);
xnor U46957 (N_46957,N_45982,N_45862);
xnor U46958 (N_46958,N_45088,N_45172);
nand U46959 (N_46959,N_45916,N_45727);
nand U46960 (N_46960,N_45927,N_45733);
or U46961 (N_46961,N_45005,N_45709);
nor U46962 (N_46962,N_45884,N_45303);
nor U46963 (N_46963,N_45864,N_45793);
or U46964 (N_46964,N_45668,N_45148);
nor U46965 (N_46965,N_45891,N_45933);
xor U46966 (N_46966,N_45269,N_45872);
or U46967 (N_46967,N_45117,N_45566);
nand U46968 (N_46968,N_45789,N_45311);
and U46969 (N_46969,N_45375,N_45507);
nor U46970 (N_46970,N_45232,N_45585);
xor U46971 (N_46971,N_45846,N_45798);
and U46972 (N_46972,N_45613,N_45151);
xnor U46973 (N_46973,N_45252,N_45383);
or U46974 (N_46974,N_45206,N_45869);
nor U46975 (N_46975,N_45483,N_45047);
xor U46976 (N_46976,N_45340,N_45720);
nor U46977 (N_46977,N_45740,N_45056);
xnor U46978 (N_46978,N_45871,N_45891);
or U46979 (N_46979,N_45934,N_45560);
or U46980 (N_46980,N_45423,N_45488);
nor U46981 (N_46981,N_45192,N_45084);
and U46982 (N_46982,N_45921,N_45614);
nand U46983 (N_46983,N_45210,N_45943);
and U46984 (N_46984,N_45664,N_45766);
or U46985 (N_46985,N_45383,N_45650);
and U46986 (N_46986,N_45850,N_45228);
and U46987 (N_46987,N_45661,N_45534);
or U46988 (N_46988,N_45633,N_45242);
xnor U46989 (N_46989,N_45918,N_45486);
nand U46990 (N_46990,N_45090,N_45109);
or U46991 (N_46991,N_45190,N_45700);
and U46992 (N_46992,N_45443,N_45884);
xor U46993 (N_46993,N_45764,N_45073);
nor U46994 (N_46994,N_45106,N_45307);
nor U46995 (N_46995,N_45872,N_45913);
or U46996 (N_46996,N_45918,N_45772);
xnor U46997 (N_46997,N_45098,N_45860);
nand U46998 (N_46998,N_45760,N_45034);
or U46999 (N_46999,N_45134,N_45174);
nor U47000 (N_47000,N_46626,N_46515);
xor U47001 (N_47001,N_46675,N_46663);
xnor U47002 (N_47002,N_46208,N_46696);
nor U47003 (N_47003,N_46300,N_46597);
xnor U47004 (N_47004,N_46790,N_46376);
and U47005 (N_47005,N_46531,N_46665);
or U47006 (N_47006,N_46335,N_46113);
nand U47007 (N_47007,N_46709,N_46939);
xor U47008 (N_47008,N_46510,N_46087);
or U47009 (N_47009,N_46913,N_46119);
and U47010 (N_47010,N_46930,N_46845);
nand U47011 (N_47011,N_46179,N_46792);
or U47012 (N_47012,N_46071,N_46981);
xnor U47013 (N_47013,N_46023,N_46272);
nor U47014 (N_47014,N_46992,N_46002);
or U47015 (N_47015,N_46761,N_46834);
or U47016 (N_47016,N_46132,N_46828);
or U47017 (N_47017,N_46338,N_46240);
or U47018 (N_47018,N_46484,N_46890);
xor U47019 (N_47019,N_46362,N_46829);
nor U47020 (N_47020,N_46588,N_46610);
xor U47021 (N_47021,N_46267,N_46157);
nand U47022 (N_47022,N_46012,N_46786);
nand U47023 (N_47023,N_46088,N_46823);
and U47024 (N_47024,N_46681,N_46202);
or U47025 (N_47025,N_46396,N_46566);
nor U47026 (N_47026,N_46833,N_46098);
or U47027 (N_47027,N_46228,N_46747);
nand U47028 (N_47028,N_46928,N_46985);
nor U47029 (N_47029,N_46135,N_46476);
nor U47030 (N_47030,N_46882,N_46975);
or U47031 (N_47031,N_46474,N_46957);
or U47032 (N_47032,N_46863,N_46400);
nor U47033 (N_47033,N_46371,N_46598);
nand U47034 (N_47034,N_46674,N_46806);
nor U47035 (N_47035,N_46117,N_46528);
nor U47036 (N_47036,N_46082,N_46770);
xnor U47037 (N_47037,N_46751,N_46648);
nor U47038 (N_47038,N_46193,N_46838);
nand U47039 (N_47039,N_46501,N_46775);
and U47040 (N_47040,N_46144,N_46561);
and U47041 (N_47041,N_46105,N_46938);
xnor U47042 (N_47042,N_46329,N_46931);
xor U47043 (N_47043,N_46655,N_46980);
xnor U47044 (N_47044,N_46427,N_46698);
nor U47045 (N_47045,N_46497,N_46437);
and U47046 (N_47046,N_46430,N_46115);
or U47047 (N_47047,N_46918,N_46298);
or U47048 (N_47048,N_46529,N_46488);
nand U47049 (N_47049,N_46956,N_46988);
and U47050 (N_47050,N_46435,N_46051);
nor U47051 (N_47051,N_46707,N_46814);
xor U47052 (N_47052,N_46892,N_46408);
or U47053 (N_47053,N_46316,N_46619);
nor U47054 (N_47054,N_46263,N_46916);
or U47055 (N_47055,N_46120,N_46409);
nand U47056 (N_47056,N_46744,N_46702);
xnor U47057 (N_47057,N_46024,N_46965);
or U47058 (N_47058,N_46549,N_46962);
nor U47059 (N_47059,N_46780,N_46246);
and U47060 (N_47060,N_46230,N_46537);
nor U47061 (N_47061,N_46213,N_46449);
nor U47062 (N_47062,N_46539,N_46204);
nor U47063 (N_47063,N_46960,N_46124);
and U47064 (N_47064,N_46948,N_46363);
xnor U47065 (N_47065,N_46609,N_46274);
nor U47066 (N_47066,N_46705,N_46116);
or U47067 (N_47067,N_46130,N_46061);
nor U47068 (N_47068,N_46617,N_46827);
nor U47069 (N_47069,N_46391,N_46065);
nand U47070 (N_47070,N_46028,N_46731);
xor U47071 (N_47071,N_46352,N_46565);
or U47072 (N_47072,N_46434,N_46909);
or U47073 (N_47073,N_46982,N_46604);
nor U47074 (N_47074,N_46669,N_46540);
and U47075 (N_47075,N_46252,N_46643);
or U47076 (N_47076,N_46802,N_46671);
or U47077 (N_47077,N_46191,N_46111);
nand U47078 (N_47078,N_46134,N_46893);
nor U47079 (N_47079,N_46929,N_46189);
and U47080 (N_47080,N_46219,N_46884);
xor U47081 (N_47081,N_46425,N_46746);
nand U47082 (N_47082,N_46046,N_46820);
nor U47083 (N_47083,N_46270,N_46322);
nand U47084 (N_47084,N_46968,N_46294);
and U47085 (N_47085,N_46078,N_46354);
or U47086 (N_47086,N_46718,N_46291);
nand U47087 (N_47087,N_46852,N_46587);
or U47088 (N_47088,N_46795,N_46390);
nor U47089 (N_47089,N_46879,N_46868);
and U47090 (N_47090,N_46021,N_46771);
nor U47091 (N_47091,N_46285,N_46000);
nand U47092 (N_47092,N_46320,N_46813);
nand U47093 (N_47093,N_46011,N_46997);
xnor U47094 (N_47094,N_46872,N_46612);
nor U47095 (N_47095,N_46282,N_46108);
or U47096 (N_47096,N_46367,N_46420);
and U47097 (N_47097,N_46917,N_46682);
and U47098 (N_47098,N_46613,N_46504);
nor U47099 (N_47099,N_46060,N_46458);
nand U47100 (N_47100,N_46001,N_46791);
nand U47101 (N_47101,N_46239,N_46182);
xnor U47102 (N_47102,N_46265,N_46532);
xor U47103 (N_47103,N_46723,N_46278);
and U47104 (N_47104,N_46689,N_46570);
nand U47105 (N_47105,N_46932,N_46704);
and U47106 (N_47106,N_46417,N_46512);
and U47107 (N_47107,N_46952,N_46197);
nand U47108 (N_47108,N_46480,N_46624);
or U47109 (N_47109,N_46336,N_46749);
nor U47110 (N_47110,N_46978,N_46853);
and U47111 (N_47111,N_46547,N_46620);
xor U47112 (N_47112,N_46946,N_46578);
nor U47113 (N_47113,N_46866,N_46407);
nor U47114 (N_47114,N_46092,N_46927);
nand U47115 (N_47115,N_46936,N_46653);
and U47116 (N_47116,N_46573,N_46846);
and U47117 (N_47117,N_46594,N_46154);
nor U47118 (N_47118,N_46045,N_46777);
xor U47119 (N_47119,N_46646,N_46990);
and U47120 (N_47120,N_46217,N_46768);
nand U47121 (N_47121,N_46100,N_46888);
or U47122 (N_47122,N_46050,N_46779);
and U47123 (N_47123,N_46279,N_46178);
nand U47124 (N_47124,N_46171,N_46589);
or U47125 (N_47125,N_46077,N_46805);
xor U47126 (N_47126,N_46824,N_46926);
xnor U47127 (N_47127,N_46373,N_46538);
or U47128 (N_47128,N_46740,N_46089);
xor U47129 (N_47129,N_46614,N_46688);
and U47130 (N_47130,N_46439,N_46207);
and U47131 (N_47131,N_46348,N_46526);
xor U47132 (N_47132,N_46977,N_46013);
and U47133 (N_47133,N_46621,N_46037);
or U47134 (N_47134,N_46163,N_46462);
xor U47135 (N_47135,N_46642,N_46634);
or U47136 (N_47136,N_46714,N_46104);
nand U47137 (N_47137,N_46495,N_46787);
xor U47138 (N_47138,N_46843,N_46874);
or U47139 (N_47139,N_46752,N_46081);
and U47140 (N_47140,N_46861,N_46577);
nor U47141 (N_47141,N_46954,N_46034);
and U47142 (N_47142,N_46247,N_46914);
nor U47143 (N_47143,N_46582,N_46891);
and U47144 (N_47144,N_46235,N_46195);
and U47145 (N_47145,N_46651,N_46138);
or U47146 (N_47146,N_46428,N_46881);
nor U47147 (N_47147,N_46708,N_46542);
and U47148 (N_47148,N_46374,N_46772);
xor U47149 (N_47149,N_46382,N_46266);
nand U47150 (N_47150,N_46377,N_46900);
nor U47151 (N_47151,N_46623,N_46911);
and U47152 (N_47152,N_46052,N_46993);
nor U47153 (N_47153,N_46122,N_46940);
or U47154 (N_47154,N_46935,N_46636);
or U47155 (N_47155,N_46148,N_46769);
nand U47156 (N_47156,N_46137,N_46221);
xor U47157 (N_47157,N_46330,N_46155);
or U47158 (N_47158,N_46210,N_46840);
or U47159 (N_47159,N_46543,N_46386);
and U47160 (N_47160,N_46344,N_46712);
and U47161 (N_47161,N_46477,N_46019);
and U47162 (N_47162,N_46234,N_46987);
nand U47163 (N_47163,N_46678,N_46258);
and U47164 (N_47164,N_46466,N_46033);
xor U47165 (N_47165,N_46017,N_46699);
nand U47166 (N_47166,N_46307,N_46158);
or U47167 (N_47167,N_46557,N_46735);
xnor U47168 (N_47168,N_46128,N_46575);
nand U47169 (N_47169,N_46465,N_46535);
xnor U47170 (N_47170,N_46516,N_46209);
nor U47171 (N_47171,N_46405,N_46722);
and U47172 (N_47172,N_46734,N_46030);
xnor U47173 (N_47173,N_46273,N_46485);
xnor U47174 (N_47174,N_46924,N_46706);
nand U47175 (N_47175,N_46225,N_46763);
and U47176 (N_47176,N_46831,N_46934);
or U47177 (N_47177,N_46743,N_46072);
or U47178 (N_47178,N_46850,N_46103);
nor U47179 (N_47179,N_46498,N_46507);
nor U47180 (N_47180,N_46378,N_46166);
and U47181 (N_47181,N_46093,N_46313);
nand U47182 (N_47182,N_46441,N_46862);
nor U47183 (N_47183,N_46821,N_46905);
nand U47184 (N_47184,N_46963,N_46585);
xnor U47185 (N_47185,N_46438,N_46793);
nor U47186 (N_47186,N_46762,N_46967);
nor U47187 (N_47187,N_46925,N_46715);
nand U47188 (N_47188,N_46174,N_46640);
nor U47189 (N_47189,N_46416,N_46605);
nand U47190 (N_47190,N_46342,N_46830);
xnor U47191 (N_47191,N_46309,N_46851);
nand U47192 (N_47192,N_46680,N_46842);
nand U47193 (N_47193,N_46295,N_46555);
xnor U47194 (N_47194,N_46513,N_46522);
nor U47195 (N_47195,N_46215,N_46090);
or U47196 (N_47196,N_46574,N_46679);
and U47197 (N_47197,N_46016,N_46327);
nand U47198 (N_47198,N_46350,N_46053);
nor U47199 (N_47199,N_46760,N_46541);
and U47200 (N_47200,N_46844,N_46554);
nor U47201 (N_47201,N_46020,N_46937);
or U47202 (N_47202,N_46256,N_46657);
and U47203 (N_47203,N_46281,N_46717);
nand U47204 (N_47204,N_46901,N_46347);
nand U47205 (N_47205,N_46553,N_46062);
and U47206 (N_47206,N_46955,N_46592);
and U47207 (N_47207,N_46687,N_46175);
and U47208 (N_47208,N_46206,N_46452);
xnor U47209 (N_47209,N_46530,N_46737);
nor U47210 (N_47210,N_46661,N_46798);
nand U47211 (N_47211,N_46470,N_46750);
xor U47212 (N_47212,N_46136,N_46857);
and U47213 (N_47213,N_46563,N_46880);
nand U47214 (N_47214,N_46271,N_46066);
nor U47215 (N_47215,N_46152,N_46738);
nand U47216 (N_47216,N_46920,N_46625);
xnor U47217 (N_47217,N_46943,N_46630);
nor U47218 (N_47218,N_46287,N_46616);
xor U47219 (N_47219,N_46710,N_46442);
nor U47220 (N_47220,N_46736,N_46748);
nand U47221 (N_47221,N_46603,N_46472);
nand U47222 (N_47222,N_46248,N_46701);
nand U47223 (N_47223,N_46164,N_46172);
xnor U47224 (N_47224,N_46035,N_46499);
xor U47225 (N_47225,N_46895,N_46832);
or U47226 (N_47226,N_46633,N_46724);
xor U47227 (N_47227,N_46010,N_46533);
nand U47228 (N_47228,N_46318,N_46835);
xor U47229 (N_47229,N_46292,N_46290);
nand U47230 (N_47230,N_46397,N_46475);
and U47231 (N_47231,N_46875,N_46162);
and U47232 (N_47232,N_46922,N_46123);
nand U47233 (N_47233,N_46886,N_46903);
nor U47234 (N_47234,N_46058,N_46500);
xor U47235 (N_47235,N_46536,N_46101);
nand U47236 (N_47236,N_46983,N_46455);
and U47237 (N_47237,N_46085,N_46907);
or U47238 (N_47238,N_46898,N_46096);
or U47239 (N_47239,N_46331,N_46126);
and U47240 (N_47240,N_46807,N_46356);
or U47241 (N_47241,N_46146,N_46402);
nand U47242 (N_47242,N_46725,N_46676);
and U47243 (N_47243,N_46794,N_46068);
and U47244 (N_47244,N_46871,N_46176);
and U47245 (N_47245,N_46112,N_46431);
nand U47246 (N_47246,N_46200,N_46190);
or U47247 (N_47247,N_46027,N_46127);
xor U47248 (N_47248,N_46659,N_46423);
xor U47249 (N_47249,N_46328,N_46481);
nor U47250 (N_47250,N_46494,N_46305);
and U47251 (N_47251,N_46662,N_46569);
and U47252 (N_47252,N_46550,N_46581);
xnor U47253 (N_47253,N_46783,N_46995);
and U47254 (N_47254,N_46479,N_46042);
and U47255 (N_47255,N_46600,N_46877);
nand U47256 (N_47256,N_46118,N_46556);
or U47257 (N_47257,N_46627,N_46493);
nor U47258 (N_47258,N_46008,N_46804);
xor U47259 (N_47259,N_46822,N_46873);
and U47260 (N_47260,N_46047,N_46385);
xnor U47261 (N_47261,N_46583,N_46076);
nor U47262 (N_47262,N_46357,N_46375);
nor U47263 (N_47263,N_46406,N_46694);
xor U47264 (N_47264,N_46684,N_46099);
nand U47265 (N_47265,N_46319,N_46433);
and U47266 (N_47266,N_46383,N_46448);
nand U47267 (N_47267,N_46816,N_46534);
nor U47268 (N_47268,N_46564,N_46854);
xnor U47269 (N_47269,N_46260,N_46482);
and U47270 (N_47270,N_46490,N_46505);
xnor U47271 (N_47271,N_46576,N_46847);
nand U47272 (N_47272,N_46489,N_46227);
or U47273 (N_47273,N_46629,N_46183);
and U47274 (N_47274,N_46341,N_46483);
and U47275 (N_47275,N_46048,N_46959);
nand U47276 (N_47276,N_46593,N_46766);
or U47277 (N_47277,N_46635,N_46022);
or U47278 (N_47278,N_46140,N_46083);
and U47279 (N_47279,N_46170,N_46496);
xor U47280 (N_47280,N_46692,N_46237);
nand U47281 (N_47281,N_46360,N_46222);
xnor U47282 (N_47282,N_46075,N_46067);
and U47283 (N_47283,N_46401,N_46301);
nand U47284 (N_47284,N_46459,N_46333);
or U47285 (N_47285,N_46325,N_46141);
nand U47286 (N_47286,N_46580,N_46364);
nand U47287 (N_47287,N_46859,N_46226);
nor U47288 (N_47288,N_46520,N_46941);
xnor U47289 (N_47289,N_46224,N_46837);
nand U47290 (N_47290,N_46177,N_46860);
nor U47291 (N_47291,N_46976,N_46796);
nand U47292 (N_47292,N_46615,N_46055);
and U47293 (N_47293,N_46186,N_46006);
and U47294 (N_47294,N_46685,N_46317);
and U47295 (N_47295,N_46789,N_46973);
and U47296 (N_47296,N_46720,N_46242);
xnor U47297 (N_47297,N_46690,N_46080);
xor U47298 (N_47298,N_46032,N_46180);
and U47299 (N_47299,N_46131,N_46218);
nor U47300 (N_47300,N_46697,N_46848);
xnor U47301 (N_47301,N_46801,N_46054);
or U47302 (N_47302,N_46194,N_46953);
and U47303 (N_47303,N_46889,N_46369);
or U47304 (N_47304,N_46173,N_46057);
nand U47305 (N_47305,N_46043,N_46713);
nor U47306 (N_47306,N_46602,N_46314);
nor U47307 (N_47307,N_46579,N_46921);
nor U47308 (N_47308,N_46168,N_46346);
and U47309 (N_47309,N_46064,N_46961);
nand U47310 (N_47310,N_46560,N_46964);
and U47311 (N_47311,N_46185,N_46184);
or U47312 (N_47312,N_46109,N_46996);
or U47313 (N_47313,N_46899,N_46800);
nand U47314 (N_47314,N_46711,N_46897);
nand U47315 (N_47315,N_46029,N_46393);
nor U47316 (N_47316,N_46232,N_46611);
nor U47317 (N_47317,N_46492,N_46461);
or U47318 (N_47318,N_46915,N_46716);
and U47319 (N_47319,N_46729,N_46261);
xnor U47320 (N_47320,N_46359,N_46608);
nor U47321 (N_47321,N_46403,N_46858);
xnor U47322 (N_47322,N_46151,N_46381);
and U47323 (N_47323,N_46432,N_46644);
or U47324 (N_47324,N_46686,N_46264);
xnor U47325 (N_47325,N_46788,N_46632);
nand U47326 (N_47326,N_46421,N_46870);
or U47327 (N_47327,N_46815,N_46436);
xor U47328 (N_47328,N_46638,N_46041);
xor U47329 (N_47329,N_46277,N_46003);
or U47330 (N_47330,N_46262,N_46398);
or U47331 (N_47331,N_46049,N_46097);
and U47332 (N_47332,N_46323,N_46074);
xnor U47333 (N_47333,N_46836,N_46351);
nor U47334 (N_47334,N_46031,N_46269);
xnor U47335 (N_47335,N_46739,N_46683);
xor U47336 (N_47336,N_46399,N_46220);
nor U47337 (N_47337,N_46456,N_46203);
or U47338 (N_47338,N_46673,N_46551);
xnor U47339 (N_47339,N_46241,N_46293);
nand U47340 (N_47340,N_46389,N_46809);
or U47341 (N_47341,N_46776,N_46312);
or U47342 (N_47342,N_46084,N_46424);
or U47343 (N_47343,N_46753,N_46114);
nand U47344 (N_47344,N_46559,N_46243);
and U47345 (N_47345,N_46149,N_46044);
xnor U47346 (N_47346,N_46728,N_46147);
nand U47347 (N_47347,N_46949,N_46288);
nand U47348 (N_47348,N_46667,N_46308);
or U47349 (N_47349,N_46971,N_46810);
nand U47350 (N_47350,N_46797,N_46365);
or U47351 (N_47351,N_46649,N_46896);
nor U47352 (N_47352,N_46411,N_46999);
nor U47353 (N_47353,N_46631,N_46572);
or U47354 (N_47354,N_46009,N_46394);
xnor U47355 (N_47355,N_46742,N_46414);
nand U47356 (N_47356,N_46658,N_46601);
nor U47357 (N_47357,N_46785,N_46599);
or U47358 (N_47358,N_46595,N_46250);
nor U47359 (N_47359,N_46395,N_46527);
and U47360 (N_47360,N_46906,N_46759);
nand U47361 (N_47361,N_46422,N_46639);
and U47362 (N_47362,N_46018,N_46102);
xor U47363 (N_47363,N_46201,N_46388);
xnor U47364 (N_47364,N_46869,N_46817);
or U47365 (N_47365,N_46606,N_46110);
or U47366 (N_47366,N_46571,N_46511);
xnor U47367 (N_47367,N_46418,N_46473);
or U47368 (N_47368,N_46641,N_46666);
and U47369 (N_47369,N_46703,N_46645);
and U47370 (N_47370,N_46894,N_46544);
xor U47371 (N_47371,N_46463,N_46453);
xnor U47372 (N_47372,N_46091,N_46904);
and U47373 (N_47373,N_46984,N_46345);
and U47374 (N_47374,N_46404,N_46289);
and U47375 (N_47375,N_46826,N_46998);
and U47376 (N_47376,N_46259,N_46958);
nand U47377 (N_47377,N_46966,N_46214);
or U47378 (N_47378,N_46303,N_46812);
nor U47379 (N_47379,N_46370,N_46015);
or U47380 (N_47380,N_46864,N_46159);
nor U47381 (N_47381,N_46412,N_46656);
and U47382 (N_47382,N_46519,N_46025);
or U47383 (N_47383,N_46244,N_46637);
and U47384 (N_47384,N_46811,N_46517);
and U47385 (N_47385,N_46150,N_46036);
xnor U47386 (N_47386,N_46677,N_46161);
and U47387 (N_47387,N_46302,N_46469);
or U47388 (N_47388,N_46143,N_46231);
and U47389 (N_47389,N_46361,N_46415);
nor U47390 (N_47390,N_46670,N_46951);
nand U47391 (N_47391,N_46607,N_46254);
xnor U47392 (N_47392,N_46086,N_46908);
xor U47393 (N_47393,N_46945,N_46764);
nor U47394 (N_47394,N_46596,N_46063);
and U47395 (N_47395,N_46196,N_46387);
nor U47396 (N_47396,N_46919,N_46169);
or U47397 (N_47397,N_46070,N_46622);
nand U47398 (N_47398,N_46545,N_46216);
xor U47399 (N_47399,N_46107,N_46974);
nor U47400 (N_47400,N_46306,N_46767);
xnor U47401 (N_47401,N_46876,N_46487);
and U47402 (N_47402,N_46745,N_46211);
and U47403 (N_47403,N_46558,N_46521);
xor U47404 (N_47404,N_46758,N_46145);
or U47405 (N_47405,N_46887,N_46839);
nor U47406 (N_47406,N_46310,N_46756);
nor U47407 (N_47407,N_46584,N_46368);
or U47408 (N_47408,N_46525,N_46503);
xnor U47409 (N_47409,N_46774,N_46353);
xnor U47410 (N_47410,N_46446,N_46719);
xnor U47411 (N_47411,N_46865,N_46546);
nor U47412 (N_47412,N_46133,N_46491);
nand U47413 (N_47413,N_46276,N_46129);
and U47414 (N_47414,N_46095,N_46855);
and U47415 (N_47415,N_46552,N_46808);
xnor U47416 (N_47416,N_46524,N_46972);
nand U47417 (N_47417,N_46384,N_46647);
or U47418 (N_47418,N_46486,N_46343);
xor U47419 (N_47419,N_46073,N_46590);
nor U47420 (N_47420,N_46450,N_46268);
and U47421 (N_47421,N_46094,N_46334);
xor U47422 (N_47422,N_46502,N_46355);
and U47423 (N_47423,N_46280,N_46568);
xor U47424 (N_47424,N_46125,N_46142);
xor U47425 (N_47425,N_46754,N_46618);
or U47426 (N_47426,N_46199,N_46192);
xnor U47427 (N_47427,N_46315,N_46650);
nor U47428 (N_47428,N_46726,N_46304);
nor U47429 (N_47429,N_46160,N_46257);
nand U47430 (N_47430,N_46167,N_46284);
and U47431 (N_47431,N_46757,N_46950);
nor U47432 (N_47432,N_46885,N_46471);
or U47433 (N_47433,N_46039,N_46467);
and U47434 (N_47434,N_46188,N_46730);
nand U47435 (N_47435,N_46181,N_46591);
nor U47436 (N_47436,N_46040,N_46198);
and U47437 (N_47437,N_46562,N_46668);
xnor U47438 (N_47438,N_46238,N_46819);
xor U47439 (N_47439,N_46825,N_46139);
nand U47440 (N_47440,N_46392,N_46508);
nand U47441 (N_47441,N_46379,N_46229);
nor U47442 (N_47442,N_46784,N_46969);
or U47443 (N_47443,N_46443,N_46339);
nand U47444 (N_47444,N_46841,N_46007);
nor U47445 (N_47445,N_46933,N_46165);
xnor U47446 (N_47446,N_46912,N_46445);
or U47447 (N_47447,N_46514,N_46233);
or U47448 (N_47448,N_46283,N_46223);
nor U47449 (N_47449,N_46297,N_46741);
or U47450 (N_47450,N_46755,N_46253);
xor U47451 (N_47451,N_46358,N_46380);
and U47452 (N_47452,N_46251,N_46413);
nand U47453 (N_47453,N_46332,N_46447);
xnor U47454 (N_47454,N_46444,N_46468);
nand U47455 (N_47455,N_46700,N_46153);
or U47456 (N_47456,N_46156,N_46994);
and U47457 (N_47457,N_46245,N_46349);
nand U47458 (N_47458,N_46340,N_46773);
nor U47459 (N_47459,N_46454,N_46778);
nand U47460 (N_47460,N_46026,N_46628);
and U47461 (N_47461,N_46464,N_46321);
nor U47462 (N_47462,N_46275,N_46249);
nor U47463 (N_47463,N_46986,N_46014);
and U47464 (N_47464,N_46296,N_46038);
or U47465 (N_47465,N_46652,N_46799);
or U47466 (N_47466,N_46672,N_46664);
nand U47467 (N_47467,N_46732,N_46947);
xnor U47468 (N_47468,N_46457,N_46944);
nor U47469 (N_47469,N_46326,N_46069);
xor U47470 (N_47470,N_46460,N_46372);
nand U47471 (N_47471,N_46849,N_46883);
nor U47472 (N_47472,N_46366,N_46781);
xor U47473 (N_47473,N_46299,N_46255);
xor U47474 (N_47474,N_46187,N_46989);
nand U47475 (N_47475,N_46324,N_46782);
or U47476 (N_47476,N_46212,N_46506);
or U47477 (N_47477,N_46440,N_46970);
nand U47478 (N_47478,N_46004,N_46518);
and U47479 (N_47479,N_46733,N_46079);
or U47480 (N_47480,N_46056,N_46691);
nand U47481 (N_47481,N_46567,N_46586);
xnor U47482 (N_47482,N_46523,N_46721);
xnor U47483 (N_47483,N_46878,N_46451);
and U47484 (N_47484,N_46236,N_46942);
nor U47485 (N_47485,N_46205,N_46121);
xor U47486 (N_47486,N_46910,N_46695);
nor U47487 (N_47487,N_46654,N_46991);
nand U47488 (N_47488,N_46059,N_46311);
xnor U47489 (N_47489,N_46979,N_46856);
or U47490 (N_47490,N_46548,N_46803);
or U47491 (N_47491,N_46509,N_46429);
or U47492 (N_47492,N_46419,N_46923);
xor U47493 (N_47493,N_46727,N_46005);
nand U47494 (N_47494,N_46660,N_46867);
nor U47495 (N_47495,N_46765,N_46478);
nor U47496 (N_47496,N_46337,N_46693);
and U47497 (N_47497,N_46410,N_46818);
nor U47498 (N_47498,N_46286,N_46902);
or U47499 (N_47499,N_46106,N_46426);
and U47500 (N_47500,N_46469,N_46859);
nor U47501 (N_47501,N_46771,N_46143);
xnor U47502 (N_47502,N_46292,N_46931);
nand U47503 (N_47503,N_46899,N_46153);
nand U47504 (N_47504,N_46098,N_46405);
and U47505 (N_47505,N_46227,N_46130);
xnor U47506 (N_47506,N_46165,N_46442);
nor U47507 (N_47507,N_46690,N_46862);
or U47508 (N_47508,N_46718,N_46578);
nand U47509 (N_47509,N_46525,N_46509);
xnor U47510 (N_47510,N_46075,N_46650);
nor U47511 (N_47511,N_46309,N_46140);
or U47512 (N_47512,N_46707,N_46722);
or U47513 (N_47513,N_46844,N_46458);
nand U47514 (N_47514,N_46246,N_46700);
or U47515 (N_47515,N_46498,N_46238);
and U47516 (N_47516,N_46882,N_46395);
nand U47517 (N_47517,N_46475,N_46414);
nand U47518 (N_47518,N_46138,N_46562);
or U47519 (N_47519,N_46062,N_46241);
or U47520 (N_47520,N_46489,N_46492);
xnor U47521 (N_47521,N_46022,N_46352);
xor U47522 (N_47522,N_46349,N_46958);
or U47523 (N_47523,N_46608,N_46274);
nand U47524 (N_47524,N_46623,N_46327);
nor U47525 (N_47525,N_46855,N_46414);
nand U47526 (N_47526,N_46152,N_46530);
nor U47527 (N_47527,N_46310,N_46380);
xor U47528 (N_47528,N_46418,N_46724);
nor U47529 (N_47529,N_46944,N_46008);
or U47530 (N_47530,N_46220,N_46226);
xnor U47531 (N_47531,N_46351,N_46821);
xor U47532 (N_47532,N_46875,N_46894);
nor U47533 (N_47533,N_46425,N_46467);
nor U47534 (N_47534,N_46278,N_46362);
xnor U47535 (N_47535,N_46502,N_46640);
nand U47536 (N_47536,N_46995,N_46748);
and U47537 (N_47537,N_46823,N_46668);
and U47538 (N_47538,N_46337,N_46729);
and U47539 (N_47539,N_46883,N_46404);
or U47540 (N_47540,N_46393,N_46987);
nand U47541 (N_47541,N_46765,N_46751);
nor U47542 (N_47542,N_46735,N_46473);
and U47543 (N_47543,N_46995,N_46521);
or U47544 (N_47544,N_46732,N_46189);
and U47545 (N_47545,N_46289,N_46260);
xnor U47546 (N_47546,N_46726,N_46953);
nand U47547 (N_47547,N_46702,N_46971);
and U47548 (N_47548,N_46943,N_46972);
or U47549 (N_47549,N_46060,N_46108);
xnor U47550 (N_47550,N_46644,N_46223);
or U47551 (N_47551,N_46765,N_46312);
xor U47552 (N_47552,N_46705,N_46158);
and U47553 (N_47553,N_46313,N_46477);
nand U47554 (N_47554,N_46498,N_46947);
xnor U47555 (N_47555,N_46175,N_46139);
and U47556 (N_47556,N_46091,N_46267);
nand U47557 (N_47557,N_46713,N_46781);
xor U47558 (N_47558,N_46767,N_46502);
nand U47559 (N_47559,N_46206,N_46140);
nor U47560 (N_47560,N_46583,N_46424);
nor U47561 (N_47561,N_46661,N_46626);
and U47562 (N_47562,N_46579,N_46571);
nor U47563 (N_47563,N_46679,N_46278);
or U47564 (N_47564,N_46815,N_46124);
xor U47565 (N_47565,N_46120,N_46181);
nor U47566 (N_47566,N_46438,N_46579);
nor U47567 (N_47567,N_46242,N_46443);
nand U47568 (N_47568,N_46092,N_46516);
xor U47569 (N_47569,N_46012,N_46520);
nand U47570 (N_47570,N_46866,N_46991);
and U47571 (N_47571,N_46561,N_46211);
nand U47572 (N_47572,N_46722,N_46442);
nor U47573 (N_47573,N_46924,N_46340);
and U47574 (N_47574,N_46605,N_46809);
and U47575 (N_47575,N_46299,N_46908);
nand U47576 (N_47576,N_46084,N_46800);
or U47577 (N_47577,N_46161,N_46786);
or U47578 (N_47578,N_46411,N_46496);
nand U47579 (N_47579,N_46459,N_46187);
and U47580 (N_47580,N_46611,N_46643);
nor U47581 (N_47581,N_46841,N_46563);
xnor U47582 (N_47582,N_46839,N_46938);
xnor U47583 (N_47583,N_46387,N_46648);
and U47584 (N_47584,N_46112,N_46441);
or U47585 (N_47585,N_46827,N_46568);
and U47586 (N_47586,N_46855,N_46483);
nor U47587 (N_47587,N_46111,N_46941);
xnor U47588 (N_47588,N_46157,N_46473);
or U47589 (N_47589,N_46922,N_46169);
and U47590 (N_47590,N_46005,N_46892);
nand U47591 (N_47591,N_46368,N_46064);
and U47592 (N_47592,N_46207,N_46734);
or U47593 (N_47593,N_46478,N_46612);
or U47594 (N_47594,N_46928,N_46894);
or U47595 (N_47595,N_46232,N_46412);
xnor U47596 (N_47596,N_46475,N_46898);
or U47597 (N_47597,N_46891,N_46084);
and U47598 (N_47598,N_46745,N_46432);
nor U47599 (N_47599,N_46123,N_46370);
and U47600 (N_47600,N_46895,N_46176);
and U47601 (N_47601,N_46588,N_46445);
or U47602 (N_47602,N_46435,N_46903);
nand U47603 (N_47603,N_46997,N_46082);
and U47604 (N_47604,N_46560,N_46935);
or U47605 (N_47605,N_46814,N_46904);
xnor U47606 (N_47606,N_46375,N_46421);
and U47607 (N_47607,N_46260,N_46235);
nor U47608 (N_47608,N_46111,N_46370);
nor U47609 (N_47609,N_46171,N_46731);
xor U47610 (N_47610,N_46988,N_46305);
xor U47611 (N_47611,N_46869,N_46794);
or U47612 (N_47612,N_46649,N_46845);
and U47613 (N_47613,N_46344,N_46068);
or U47614 (N_47614,N_46708,N_46782);
xnor U47615 (N_47615,N_46057,N_46974);
nor U47616 (N_47616,N_46138,N_46056);
nor U47617 (N_47617,N_46841,N_46181);
nor U47618 (N_47618,N_46779,N_46276);
nor U47619 (N_47619,N_46252,N_46462);
and U47620 (N_47620,N_46382,N_46339);
or U47621 (N_47621,N_46637,N_46574);
xor U47622 (N_47622,N_46483,N_46578);
and U47623 (N_47623,N_46535,N_46829);
xnor U47624 (N_47624,N_46630,N_46458);
nor U47625 (N_47625,N_46997,N_46796);
nor U47626 (N_47626,N_46033,N_46640);
or U47627 (N_47627,N_46655,N_46659);
xor U47628 (N_47628,N_46532,N_46307);
and U47629 (N_47629,N_46103,N_46574);
xor U47630 (N_47630,N_46168,N_46920);
or U47631 (N_47631,N_46122,N_46229);
nor U47632 (N_47632,N_46437,N_46862);
and U47633 (N_47633,N_46885,N_46650);
xor U47634 (N_47634,N_46551,N_46710);
and U47635 (N_47635,N_46888,N_46831);
or U47636 (N_47636,N_46338,N_46885);
nand U47637 (N_47637,N_46698,N_46764);
nand U47638 (N_47638,N_46530,N_46778);
or U47639 (N_47639,N_46378,N_46285);
nand U47640 (N_47640,N_46791,N_46924);
nor U47641 (N_47641,N_46094,N_46463);
nand U47642 (N_47642,N_46778,N_46242);
xnor U47643 (N_47643,N_46075,N_46184);
nor U47644 (N_47644,N_46509,N_46293);
nand U47645 (N_47645,N_46843,N_46441);
xnor U47646 (N_47646,N_46228,N_46766);
or U47647 (N_47647,N_46561,N_46779);
xor U47648 (N_47648,N_46970,N_46297);
or U47649 (N_47649,N_46095,N_46624);
nor U47650 (N_47650,N_46518,N_46194);
xor U47651 (N_47651,N_46754,N_46818);
or U47652 (N_47652,N_46294,N_46499);
nand U47653 (N_47653,N_46992,N_46923);
nand U47654 (N_47654,N_46603,N_46033);
nor U47655 (N_47655,N_46218,N_46329);
or U47656 (N_47656,N_46001,N_46678);
or U47657 (N_47657,N_46453,N_46010);
nand U47658 (N_47658,N_46548,N_46512);
nand U47659 (N_47659,N_46310,N_46336);
or U47660 (N_47660,N_46486,N_46942);
or U47661 (N_47661,N_46546,N_46077);
nand U47662 (N_47662,N_46325,N_46715);
nand U47663 (N_47663,N_46311,N_46611);
and U47664 (N_47664,N_46688,N_46792);
nand U47665 (N_47665,N_46047,N_46168);
xnor U47666 (N_47666,N_46397,N_46041);
nor U47667 (N_47667,N_46004,N_46780);
and U47668 (N_47668,N_46292,N_46311);
xnor U47669 (N_47669,N_46053,N_46123);
nor U47670 (N_47670,N_46403,N_46128);
or U47671 (N_47671,N_46194,N_46205);
nand U47672 (N_47672,N_46632,N_46679);
xnor U47673 (N_47673,N_46297,N_46986);
or U47674 (N_47674,N_46821,N_46283);
xnor U47675 (N_47675,N_46139,N_46389);
xnor U47676 (N_47676,N_46497,N_46491);
or U47677 (N_47677,N_46566,N_46868);
nor U47678 (N_47678,N_46805,N_46680);
or U47679 (N_47679,N_46296,N_46668);
and U47680 (N_47680,N_46925,N_46940);
xor U47681 (N_47681,N_46978,N_46262);
xnor U47682 (N_47682,N_46892,N_46772);
nand U47683 (N_47683,N_46500,N_46837);
or U47684 (N_47684,N_46750,N_46806);
nor U47685 (N_47685,N_46506,N_46331);
xor U47686 (N_47686,N_46373,N_46356);
nand U47687 (N_47687,N_46017,N_46520);
and U47688 (N_47688,N_46662,N_46147);
nand U47689 (N_47689,N_46986,N_46316);
or U47690 (N_47690,N_46429,N_46112);
nand U47691 (N_47691,N_46953,N_46805);
or U47692 (N_47692,N_46345,N_46289);
nand U47693 (N_47693,N_46657,N_46168);
nand U47694 (N_47694,N_46062,N_46672);
nand U47695 (N_47695,N_46699,N_46544);
nand U47696 (N_47696,N_46056,N_46864);
or U47697 (N_47697,N_46008,N_46622);
and U47698 (N_47698,N_46476,N_46167);
or U47699 (N_47699,N_46190,N_46693);
and U47700 (N_47700,N_46297,N_46823);
or U47701 (N_47701,N_46793,N_46403);
and U47702 (N_47702,N_46701,N_46120);
xnor U47703 (N_47703,N_46356,N_46663);
nand U47704 (N_47704,N_46353,N_46030);
and U47705 (N_47705,N_46419,N_46090);
nor U47706 (N_47706,N_46460,N_46662);
nand U47707 (N_47707,N_46281,N_46310);
and U47708 (N_47708,N_46374,N_46862);
nand U47709 (N_47709,N_46374,N_46538);
nand U47710 (N_47710,N_46713,N_46376);
or U47711 (N_47711,N_46361,N_46482);
and U47712 (N_47712,N_46604,N_46714);
xnor U47713 (N_47713,N_46641,N_46593);
xor U47714 (N_47714,N_46800,N_46131);
nor U47715 (N_47715,N_46709,N_46003);
nand U47716 (N_47716,N_46144,N_46903);
nand U47717 (N_47717,N_46841,N_46343);
and U47718 (N_47718,N_46669,N_46086);
and U47719 (N_47719,N_46517,N_46585);
xnor U47720 (N_47720,N_46481,N_46094);
or U47721 (N_47721,N_46047,N_46381);
xor U47722 (N_47722,N_46919,N_46207);
nand U47723 (N_47723,N_46137,N_46800);
xnor U47724 (N_47724,N_46181,N_46008);
or U47725 (N_47725,N_46528,N_46573);
nor U47726 (N_47726,N_46714,N_46846);
or U47727 (N_47727,N_46092,N_46826);
and U47728 (N_47728,N_46513,N_46447);
nor U47729 (N_47729,N_46859,N_46752);
and U47730 (N_47730,N_46329,N_46582);
or U47731 (N_47731,N_46752,N_46187);
nand U47732 (N_47732,N_46848,N_46918);
xnor U47733 (N_47733,N_46693,N_46010);
nand U47734 (N_47734,N_46983,N_46075);
or U47735 (N_47735,N_46322,N_46931);
nor U47736 (N_47736,N_46353,N_46633);
nand U47737 (N_47737,N_46501,N_46189);
or U47738 (N_47738,N_46356,N_46048);
or U47739 (N_47739,N_46421,N_46774);
or U47740 (N_47740,N_46971,N_46032);
or U47741 (N_47741,N_46520,N_46022);
xnor U47742 (N_47742,N_46724,N_46205);
and U47743 (N_47743,N_46791,N_46620);
or U47744 (N_47744,N_46105,N_46610);
nand U47745 (N_47745,N_46456,N_46139);
nand U47746 (N_47746,N_46963,N_46708);
or U47747 (N_47747,N_46528,N_46932);
nand U47748 (N_47748,N_46717,N_46610);
xnor U47749 (N_47749,N_46425,N_46304);
or U47750 (N_47750,N_46401,N_46493);
nor U47751 (N_47751,N_46250,N_46847);
and U47752 (N_47752,N_46559,N_46595);
nand U47753 (N_47753,N_46960,N_46396);
nand U47754 (N_47754,N_46190,N_46911);
and U47755 (N_47755,N_46847,N_46530);
xnor U47756 (N_47756,N_46922,N_46407);
and U47757 (N_47757,N_46390,N_46478);
nand U47758 (N_47758,N_46368,N_46195);
or U47759 (N_47759,N_46492,N_46584);
xor U47760 (N_47760,N_46206,N_46280);
xor U47761 (N_47761,N_46209,N_46383);
or U47762 (N_47762,N_46395,N_46644);
xnor U47763 (N_47763,N_46123,N_46769);
nor U47764 (N_47764,N_46587,N_46808);
nor U47765 (N_47765,N_46764,N_46467);
nor U47766 (N_47766,N_46441,N_46160);
xnor U47767 (N_47767,N_46179,N_46394);
xnor U47768 (N_47768,N_46171,N_46353);
or U47769 (N_47769,N_46205,N_46198);
xnor U47770 (N_47770,N_46480,N_46052);
nand U47771 (N_47771,N_46823,N_46138);
nand U47772 (N_47772,N_46886,N_46432);
xor U47773 (N_47773,N_46249,N_46497);
or U47774 (N_47774,N_46696,N_46030);
xor U47775 (N_47775,N_46081,N_46437);
nand U47776 (N_47776,N_46199,N_46355);
nor U47777 (N_47777,N_46137,N_46365);
and U47778 (N_47778,N_46602,N_46069);
and U47779 (N_47779,N_46289,N_46658);
nor U47780 (N_47780,N_46508,N_46138);
or U47781 (N_47781,N_46922,N_46001);
nor U47782 (N_47782,N_46832,N_46601);
xnor U47783 (N_47783,N_46479,N_46663);
or U47784 (N_47784,N_46495,N_46312);
and U47785 (N_47785,N_46010,N_46229);
and U47786 (N_47786,N_46623,N_46290);
and U47787 (N_47787,N_46492,N_46425);
xnor U47788 (N_47788,N_46237,N_46411);
nor U47789 (N_47789,N_46538,N_46984);
or U47790 (N_47790,N_46605,N_46651);
nand U47791 (N_47791,N_46787,N_46942);
and U47792 (N_47792,N_46294,N_46155);
nor U47793 (N_47793,N_46456,N_46178);
nand U47794 (N_47794,N_46736,N_46168);
or U47795 (N_47795,N_46703,N_46634);
or U47796 (N_47796,N_46341,N_46168);
nor U47797 (N_47797,N_46348,N_46187);
xnor U47798 (N_47798,N_46201,N_46674);
xor U47799 (N_47799,N_46742,N_46620);
or U47800 (N_47800,N_46957,N_46758);
nand U47801 (N_47801,N_46409,N_46399);
xnor U47802 (N_47802,N_46555,N_46565);
or U47803 (N_47803,N_46171,N_46174);
and U47804 (N_47804,N_46465,N_46303);
nor U47805 (N_47805,N_46466,N_46192);
nand U47806 (N_47806,N_46819,N_46660);
nor U47807 (N_47807,N_46571,N_46541);
and U47808 (N_47808,N_46494,N_46695);
xor U47809 (N_47809,N_46956,N_46538);
and U47810 (N_47810,N_46884,N_46860);
and U47811 (N_47811,N_46923,N_46540);
or U47812 (N_47812,N_46780,N_46740);
xor U47813 (N_47813,N_46005,N_46331);
nand U47814 (N_47814,N_46248,N_46472);
or U47815 (N_47815,N_46554,N_46160);
nand U47816 (N_47816,N_46847,N_46777);
and U47817 (N_47817,N_46799,N_46783);
nor U47818 (N_47818,N_46051,N_46189);
nor U47819 (N_47819,N_46761,N_46916);
nand U47820 (N_47820,N_46384,N_46328);
and U47821 (N_47821,N_46869,N_46548);
xnor U47822 (N_47822,N_46933,N_46237);
nand U47823 (N_47823,N_46268,N_46847);
nand U47824 (N_47824,N_46466,N_46870);
and U47825 (N_47825,N_46075,N_46120);
and U47826 (N_47826,N_46899,N_46491);
and U47827 (N_47827,N_46569,N_46978);
nor U47828 (N_47828,N_46803,N_46848);
xor U47829 (N_47829,N_46789,N_46476);
or U47830 (N_47830,N_46258,N_46147);
nand U47831 (N_47831,N_46177,N_46973);
xor U47832 (N_47832,N_46679,N_46289);
nand U47833 (N_47833,N_46323,N_46587);
nor U47834 (N_47834,N_46481,N_46084);
nand U47835 (N_47835,N_46102,N_46247);
nor U47836 (N_47836,N_46395,N_46155);
nor U47837 (N_47837,N_46329,N_46057);
nand U47838 (N_47838,N_46826,N_46807);
nor U47839 (N_47839,N_46768,N_46066);
and U47840 (N_47840,N_46654,N_46248);
nor U47841 (N_47841,N_46296,N_46106);
nand U47842 (N_47842,N_46132,N_46930);
and U47843 (N_47843,N_46716,N_46897);
nor U47844 (N_47844,N_46985,N_46150);
nand U47845 (N_47845,N_46274,N_46268);
nand U47846 (N_47846,N_46562,N_46106);
xnor U47847 (N_47847,N_46302,N_46251);
xor U47848 (N_47848,N_46314,N_46756);
or U47849 (N_47849,N_46519,N_46866);
xnor U47850 (N_47850,N_46949,N_46005);
xnor U47851 (N_47851,N_46942,N_46424);
xor U47852 (N_47852,N_46170,N_46474);
or U47853 (N_47853,N_46327,N_46809);
or U47854 (N_47854,N_46882,N_46226);
xnor U47855 (N_47855,N_46813,N_46221);
nand U47856 (N_47856,N_46298,N_46218);
xor U47857 (N_47857,N_46685,N_46305);
and U47858 (N_47858,N_46783,N_46853);
and U47859 (N_47859,N_46681,N_46071);
xnor U47860 (N_47860,N_46832,N_46522);
nor U47861 (N_47861,N_46152,N_46923);
and U47862 (N_47862,N_46242,N_46812);
xor U47863 (N_47863,N_46047,N_46096);
xor U47864 (N_47864,N_46661,N_46451);
nand U47865 (N_47865,N_46548,N_46143);
and U47866 (N_47866,N_46457,N_46771);
xor U47867 (N_47867,N_46588,N_46392);
xnor U47868 (N_47868,N_46874,N_46685);
and U47869 (N_47869,N_46526,N_46582);
nand U47870 (N_47870,N_46711,N_46859);
xor U47871 (N_47871,N_46612,N_46274);
or U47872 (N_47872,N_46089,N_46633);
and U47873 (N_47873,N_46106,N_46587);
nand U47874 (N_47874,N_46946,N_46944);
xnor U47875 (N_47875,N_46254,N_46031);
or U47876 (N_47876,N_46135,N_46098);
nand U47877 (N_47877,N_46449,N_46442);
nand U47878 (N_47878,N_46152,N_46156);
nor U47879 (N_47879,N_46236,N_46811);
nor U47880 (N_47880,N_46259,N_46058);
nor U47881 (N_47881,N_46990,N_46843);
xor U47882 (N_47882,N_46145,N_46698);
and U47883 (N_47883,N_46941,N_46002);
or U47884 (N_47884,N_46267,N_46567);
xor U47885 (N_47885,N_46900,N_46141);
and U47886 (N_47886,N_46829,N_46983);
and U47887 (N_47887,N_46043,N_46541);
xnor U47888 (N_47888,N_46730,N_46586);
xnor U47889 (N_47889,N_46107,N_46412);
and U47890 (N_47890,N_46518,N_46092);
or U47891 (N_47891,N_46508,N_46280);
nor U47892 (N_47892,N_46218,N_46478);
and U47893 (N_47893,N_46027,N_46236);
xor U47894 (N_47894,N_46590,N_46990);
or U47895 (N_47895,N_46372,N_46910);
nor U47896 (N_47896,N_46646,N_46631);
or U47897 (N_47897,N_46238,N_46957);
and U47898 (N_47898,N_46281,N_46411);
or U47899 (N_47899,N_46622,N_46980);
and U47900 (N_47900,N_46590,N_46009);
xnor U47901 (N_47901,N_46942,N_46152);
nor U47902 (N_47902,N_46013,N_46911);
and U47903 (N_47903,N_46637,N_46635);
and U47904 (N_47904,N_46555,N_46077);
or U47905 (N_47905,N_46893,N_46542);
xor U47906 (N_47906,N_46194,N_46667);
xor U47907 (N_47907,N_46918,N_46000);
nor U47908 (N_47908,N_46223,N_46633);
nand U47909 (N_47909,N_46354,N_46115);
nand U47910 (N_47910,N_46937,N_46341);
or U47911 (N_47911,N_46633,N_46943);
nor U47912 (N_47912,N_46619,N_46409);
or U47913 (N_47913,N_46708,N_46863);
and U47914 (N_47914,N_46731,N_46114);
nand U47915 (N_47915,N_46013,N_46332);
xor U47916 (N_47916,N_46664,N_46813);
xor U47917 (N_47917,N_46003,N_46714);
xnor U47918 (N_47918,N_46703,N_46256);
nand U47919 (N_47919,N_46470,N_46834);
xor U47920 (N_47920,N_46555,N_46032);
and U47921 (N_47921,N_46502,N_46289);
xnor U47922 (N_47922,N_46323,N_46255);
and U47923 (N_47923,N_46358,N_46053);
and U47924 (N_47924,N_46357,N_46484);
xnor U47925 (N_47925,N_46885,N_46811);
nand U47926 (N_47926,N_46221,N_46241);
xor U47927 (N_47927,N_46984,N_46894);
nand U47928 (N_47928,N_46050,N_46220);
and U47929 (N_47929,N_46536,N_46035);
xnor U47930 (N_47930,N_46746,N_46802);
or U47931 (N_47931,N_46832,N_46632);
and U47932 (N_47932,N_46272,N_46401);
nand U47933 (N_47933,N_46939,N_46366);
and U47934 (N_47934,N_46933,N_46694);
nand U47935 (N_47935,N_46062,N_46995);
and U47936 (N_47936,N_46205,N_46033);
xor U47937 (N_47937,N_46452,N_46927);
or U47938 (N_47938,N_46468,N_46843);
or U47939 (N_47939,N_46189,N_46622);
nand U47940 (N_47940,N_46535,N_46644);
or U47941 (N_47941,N_46937,N_46293);
nand U47942 (N_47942,N_46545,N_46600);
or U47943 (N_47943,N_46613,N_46513);
nand U47944 (N_47944,N_46531,N_46890);
and U47945 (N_47945,N_46771,N_46647);
nand U47946 (N_47946,N_46206,N_46258);
xnor U47947 (N_47947,N_46554,N_46411);
nor U47948 (N_47948,N_46599,N_46198);
nand U47949 (N_47949,N_46074,N_46689);
nor U47950 (N_47950,N_46384,N_46269);
or U47951 (N_47951,N_46580,N_46312);
or U47952 (N_47952,N_46943,N_46846);
nand U47953 (N_47953,N_46061,N_46748);
and U47954 (N_47954,N_46447,N_46322);
and U47955 (N_47955,N_46244,N_46149);
nor U47956 (N_47956,N_46976,N_46360);
nor U47957 (N_47957,N_46984,N_46930);
nand U47958 (N_47958,N_46711,N_46672);
nand U47959 (N_47959,N_46250,N_46385);
nor U47960 (N_47960,N_46525,N_46014);
and U47961 (N_47961,N_46012,N_46529);
nor U47962 (N_47962,N_46502,N_46893);
or U47963 (N_47963,N_46919,N_46605);
nor U47964 (N_47964,N_46249,N_46548);
nor U47965 (N_47965,N_46688,N_46031);
or U47966 (N_47966,N_46431,N_46647);
nor U47967 (N_47967,N_46437,N_46987);
nor U47968 (N_47968,N_46197,N_46310);
xnor U47969 (N_47969,N_46726,N_46212);
or U47970 (N_47970,N_46559,N_46371);
xor U47971 (N_47971,N_46741,N_46213);
xor U47972 (N_47972,N_46802,N_46073);
nor U47973 (N_47973,N_46750,N_46005);
nor U47974 (N_47974,N_46745,N_46339);
nor U47975 (N_47975,N_46498,N_46864);
xor U47976 (N_47976,N_46694,N_46155);
nand U47977 (N_47977,N_46881,N_46644);
nand U47978 (N_47978,N_46099,N_46134);
and U47979 (N_47979,N_46443,N_46766);
xor U47980 (N_47980,N_46745,N_46282);
and U47981 (N_47981,N_46966,N_46066);
and U47982 (N_47982,N_46940,N_46014);
nand U47983 (N_47983,N_46320,N_46922);
nor U47984 (N_47984,N_46448,N_46150);
and U47985 (N_47985,N_46614,N_46746);
nor U47986 (N_47986,N_46219,N_46108);
and U47987 (N_47987,N_46014,N_46154);
nand U47988 (N_47988,N_46886,N_46781);
and U47989 (N_47989,N_46383,N_46009);
nand U47990 (N_47990,N_46217,N_46156);
or U47991 (N_47991,N_46929,N_46129);
or U47992 (N_47992,N_46524,N_46730);
and U47993 (N_47993,N_46922,N_46592);
xor U47994 (N_47994,N_46267,N_46875);
nand U47995 (N_47995,N_46167,N_46593);
and U47996 (N_47996,N_46118,N_46736);
or U47997 (N_47997,N_46262,N_46090);
nand U47998 (N_47998,N_46897,N_46794);
or U47999 (N_47999,N_46278,N_46095);
nand U48000 (N_48000,N_47203,N_47551);
xor U48001 (N_48001,N_47262,N_47119);
and U48002 (N_48002,N_47162,N_47984);
xnor U48003 (N_48003,N_47165,N_47781);
xor U48004 (N_48004,N_47032,N_47259);
xnor U48005 (N_48005,N_47773,N_47652);
or U48006 (N_48006,N_47454,N_47601);
or U48007 (N_48007,N_47382,N_47877);
nor U48008 (N_48008,N_47332,N_47820);
and U48009 (N_48009,N_47330,N_47139);
nor U48010 (N_48010,N_47358,N_47033);
or U48011 (N_48011,N_47501,N_47573);
nor U48012 (N_48012,N_47605,N_47222);
nand U48013 (N_48013,N_47530,N_47420);
and U48014 (N_48014,N_47643,N_47866);
nand U48015 (N_48015,N_47166,N_47449);
nor U48016 (N_48016,N_47253,N_47765);
xor U48017 (N_48017,N_47168,N_47925);
or U48018 (N_48018,N_47649,N_47541);
xor U48019 (N_48019,N_47475,N_47702);
xnor U48020 (N_48020,N_47658,N_47027);
and U48021 (N_48021,N_47405,N_47800);
xor U48022 (N_48022,N_47572,N_47432);
nor U48023 (N_48023,N_47574,N_47582);
xnor U48024 (N_48024,N_47410,N_47282);
and U48025 (N_48025,N_47609,N_47660);
or U48026 (N_48026,N_47948,N_47395);
nand U48027 (N_48027,N_47183,N_47163);
xnor U48028 (N_48028,N_47958,N_47860);
or U48029 (N_48029,N_47337,N_47007);
nor U48030 (N_48030,N_47568,N_47899);
nand U48031 (N_48031,N_47206,N_47876);
nor U48032 (N_48032,N_47034,N_47585);
nand U48033 (N_48033,N_47536,N_47741);
and U48034 (N_48034,N_47959,N_47224);
nor U48035 (N_48035,N_47350,N_47736);
nor U48036 (N_48036,N_47028,N_47078);
nor U48037 (N_48037,N_47468,N_47969);
or U48038 (N_48038,N_47399,N_47836);
and U48039 (N_48039,N_47193,N_47415);
nor U48040 (N_48040,N_47728,N_47005);
xor U48041 (N_48041,N_47359,N_47323);
nand U48042 (N_48042,N_47552,N_47662);
or U48043 (N_48043,N_47956,N_47608);
or U48044 (N_48044,N_47830,N_47386);
and U48045 (N_48045,N_47022,N_47264);
nand U48046 (N_48046,N_47255,N_47616);
nor U48047 (N_48047,N_47931,N_47493);
nand U48048 (N_48048,N_47819,N_47850);
nor U48049 (N_48049,N_47790,N_47451);
and U48050 (N_48050,N_47117,N_47376);
nor U48051 (N_48051,N_47476,N_47136);
and U48052 (N_48052,N_47550,N_47149);
or U48053 (N_48053,N_47708,N_47983);
or U48054 (N_48054,N_47887,N_47062);
nor U48055 (N_48055,N_47351,N_47391);
nor U48056 (N_48056,N_47654,N_47625);
xor U48057 (N_48057,N_47277,N_47327);
or U48058 (N_48058,N_47215,N_47780);
nor U48059 (N_48059,N_47578,N_47243);
and U48060 (N_48060,N_47767,N_47118);
nor U48061 (N_48061,N_47151,N_47895);
nand U48062 (N_48062,N_47651,N_47134);
nor U48063 (N_48063,N_47535,N_47706);
nor U48064 (N_48064,N_47871,N_47380);
xnor U48065 (N_48065,N_47024,N_47645);
nor U48066 (N_48066,N_47637,N_47722);
and U48067 (N_48067,N_47621,N_47875);
nor U48068 (N_48068,N_47318,N_47406);
or U48069 (N_48069,N_47065,N_47127);
nor U48070 (N_48070,N_47241,N_47029);
and U48071 (N_48071,N_47826,N_47299);
or U48072 (N_48072,N_47963,N_47999);
nor U48073 (N_48073,N_47385,N_47158);
xor U48074 (N_48074,N_47414,N_47626);
nand U48075 (N_48075,N_47281,N_47191);
and U48076 (N_48076,N_47960,N_47870);
nor U48077 (N_48077,N_47344,N_47808);
nand U48078 (N_48078,N_47863,N_47363);
nor U48079 (N_48079,N_47333,N_47310);
or U48080 (N_48080,N_47091,N_47209);
nor U48081 (N_48081,N_47976,N_47482);
or U48082 (N_48082,N_47093,N_47430);
and U48083 (N_48083,N_47140,N_47546);
nand U48084 (N_48084,N_47013,N_47031);
nor U48085 (N_48085,N_47288,N_47205);
xnor U48086 (N_48086,N_47774,N_47159);
nand U48087 (N_48087,N_47724,N_47648);
nor U48088 (N_48088,N_47698,N_47693);
and U48089 (N_48089,N_47392,N_47804);
xor U48090 (N_48090,N_47856,N_47884);
or U48091 (N_48091,N_47074,N_47740);
and U48092 (N_48092,N_47369,N_47903);
xor U48093 (N_48093,N_47153,N_47307);
and U48094 (N_48094,N_47816,N_47602);
or U48095 (N_48095,N_47575,N_47997);
and U48096 (N_48096,N_47907,N_47661);
or U48097 (N_48097,N_47686,N_47674);
and U48098 (N_48098,N_47297,N_47061);
nor U48099 (N_48099,N_47044,N_47302);
or U48100 (N_48100,N_47152,N_47272);
nor U48101 (N_48101,N_47707,N_47566);
xor U48102 (N_48102,N_47828,N_47939);
nor U48103 (N_48103,N_47064,N_47050);
nand U48104 (N_48104,N_47271,N_47635);
nor U48105 (N_48105,N_47340,N_47111);
xor U48106 (N_48106,N_47755,N_47104);
nor U48107 (N_48107,N_47279,N_47655);
or U48108 (N_48108,N_47972,N_47040);
or U48109 (N_48109,N_47135,N_47026);
and U48110 (N_48110,N_47321,N_47219);
or U48111 (N_48111,N_47371,N_47711);
and U48112 (N_48112,N_47496,N_47284);
or U48113 (N_48113,N_47543,N_47269);
or U48114 (N_48114,N_47980,N_47456);
xnor U48115 (N_48115,N_47125,N_47529);
xnor U48116 (N_48116,N_47100,N_47483);
nand U48117 (N_48117,N_47315,N_47910);
or U48118 (N_48118,N_47020,N_47717);
and U48119 (N_48119,N_47954,N_47971);
nand U48120 (N_48120,N_47250,N_47146);
or U48121 (N_48121,N_47786,N_47436);
nor U48122 (N_48122,N_47642,N_47835);
xor U48123 (N_48123,N_47996,N_47896);
or U48124 (N_48124,N_47945,N_47933);
xnor U48125 (N_48125,N_47114,N_47052);
xor U48126 (N_48126,N_47942,N_47670);
and U48127 (N_48127,N_47760,N_47977);
xor U48128 (N_48128,N_47304,N_47964);
nor U48129 (N_48129,N_47400,N_47822);
nand U48130 (N_48130,N_47782,N_47756);
nand U48131 (N_48131,N_47690,N_47677);
xor U48132 (N_48132,N_47479,N_47214);
and U48133 (N_48133,N_47116,N_47455);
or U48134 (N_48134,N_47544,N_47260);
nand U48135 (N_48135,N_47811,N_47533);
nor U48136 (N_48136,N_47054,N_47944);
xnor U48137 (N_48137,N_47081,N_47576);
nand U48138 (N_48138,N_47628,N_47060);
xor U48139 (N_48139,N_47240,N_47772);
nand U48140 (N_48140,N_47935,N_47603);
and U48141 (N_48141,N_47266,N_47700);
or U48142 (N_48142,N_47901,N_47413);
nand U48143 (N_48143,N_47107,N_47727);
or U48144 (N_48144,N_47633,N_47018);
xor U48145 (N_48145,N_47236,N_47577);
nand U48146 (N_48146,N_47370,N_47920);
or U48147 (N_48147,N_47930,N_47710);
nand U48148 (N_48148,N_47787,N_47784);
nor U48149 (N_48149,N_47893,N_47672);
and U48150 (N_48150,N_47381,N_47067);
nor U48151 (N_48151,N_47101,N_47926);
nor U48152 (N_48152,N_47505,N_47619);
nor U48153 (N_48153,N_47199,N_47594);
xor U48154 (N_48154,N_47810,N_47882);
nand U48155 (N_48155,N_47495,N_47775);
xnor U48156 (N_48156,N_47831,N_47268);
nand U48157 (N_48157,N_47053,N_47748);
xor U48158 (N_48158,N_47604,N_47957);
nor U48159 (N_48159,N_47319,N_47187);
nor U48160 (N_48160,N_47172,N_47657);
nor U48161 (N_48161,N_47390,N_47889);
nand U48162 (N_48162,N_47004,N_47730);
nor U48163 (N_48163,N_47975,N_47834);
nand U48164 (N_48164,N_47331,N_47967);
nand U48165 (N_48165,N_47562,N_47929);
xnor U48166 (N_48166,N_47868,N_47750);
or U48167 (N_48167,N_47557,N_47325);
and U48168 (N_48168,N_47886,N_47154);
and U48169 (N_48169,N_47865,N_47416);
nor U48170 (N_48170,N_47195,N_47854);
xor U48171 (N_48171,N_47855,N_47225);
xnor U48172 (N_48172,N_47946,N_47444);
xor U48173 (N_48173,N_47442,N_47192);
nand U48174 (N_48174,N_47144,N_47766);
or U48175 (N_48175,N_47681,N_47785);
xor U48176 (N_48176,N_47885,N_47547);
and U48177 (N_48177,N_47070,N_47611);
nand U48178 (N_48178,N_47063,N_47564);
nor U48179 (N_48179,N_47082,N_47035);
and U48180 (N_48180,N_47129,N_47313);
xnor U48181 (N_48181,N_47825,N_47844);
nor U48182 (N_48182,N_47751,N_47675);
nor U48183 (N_48183,N_47764,N_47968);
xnor U48184 (N_48184,N_47987,N_47937);
nor U48185 (N_48185,N_47261,N_47368);
nand U48186 (N_48186,N_47754,N_47487);
nand U48187 (N_48187,N_47394,N_47752);
xnor U48188 (N_48188,N_47174,N_47056);
xnor U48189 (N_48189,N_47098,N_47057);
and U48190 (N_48190,N_47915,N_47913);
and U48191 (N_48191,N_47460,N_47008);
nand U48192 (N_48192,N_47596,N_47273);
or U48193 (N_48193,N_47248,N_47580);
xnor U48194 (N_48194,N_47528,N_47458);
and U48195 (N_48195,N_47612,N_47988);
and U48196 (N_48196,N_47106,N_47579);
xor U48197 (N_48197,N_47881,N_47978);
nor U48198 (N_48198,N_47510,N_47296);
xor U48199 (N_48199,N_47000,N_47137);
or U48200 (N_48200,N_47590,N_47631);
nor U48201 (N_48201,N_47953,N_47570);
nor U48202 (N_48202,N_47068,N_47803);
xor U48203 (N_48203,N_47320,N_47840);
xor U48204 (N_48204,N_47077,N_47791);
xnor U48205 (N_48205,N_47108,N_47716);
nand U48206 (N_48206,N_47650,N_47328);
xor U48207 (N_48207,N_47169,N_47559);
or U48208 (N_48208,N_47897,N_47936);
or U48209 (N_48209,N_47778,N_47848);
or U48210 (N_48210,N_47898,N_47373);
nor U48211 (N_48211,N_47472,N_47179);
xnor U48212 (N_48212,N_47869,N_47814);
xnor U48213 (N_48213,N_47818,N_47586);
and U48214 (N_48214,N_47779,N_47753);
xor U48215 (N_48215,N_47744,N_47506);
nor U48216 (N_48216,N_47150,N_47883);
xor U48217 (N_48217,N_47457,N_47287);
or U48218 (N_48218,N_47290,N_47439);
nor U48219 (N_48219,N_47833,N_47538);
and U48220 (N_48220,N_47197,N_47141);
or U48221 (N_48221,N_47435,N_47667);
xnor U48222 (N_48222,N_47364,N_47220);
xor U48223 (N_48223,N_47425,N_47204);
nand U48224 (N_48224,N_47839,N_47384);
or U48225 (N_48225,N_47402,N_47914);
nor U48226 (N_48226,N_47237,N_47862);
nor U48227 (N_48227,N_47792,N_47326);
or U48228 (N_48228,N_47389,N_47673);
and U48229 (N_48229,N_47481,N_47979);
nand U48230 (N_48230,N_47143,N_47469);
nor U48231 (N_48231,N_47951,N_47096);
nand U48232 (N_48232,N_47419,N_47503);
or U48233 (N_48233,N_47847,N_47746);
xor U48234 (N_48234,N_47275,N_47689);
xnor U48235 (N_48235,N_47905,N_47294);
nor U48236 (N_48236,N_47429,N_47488);
or U48237 (N_48237,N_47556,N_47545);
or U48238 (N_48238,N_47265,N_47995);
nand U48239 (N_48239,N_47059,N_47335);
nand U48240 (N_48240,N_47043,N_47042);
nor U48241 (N_48241,N_47170,N_47998);
nor U48242 (N_48242,N_47726,N_47156);
xnor U48243 (N_48243,N_47485,N_47176);
or U48244 (N_48244,N_47086,N_47598);
and U48245 (N_48245,N_47798,N_47807);
xnor U48246 (N_48246,N_47103,N_47037);
xor U48247 (N_48247,N_47902,N_47286);
and U48248 (N_48248,N_47521,N_47525);
and U48249 (N_48249,N_47298,N_47409);
and U48250 (N_48250,N_47084,N_47880);
nand U48251 (N_48251,N_47947,N_47105);
xor U48252 (N_48252,N_47424,N_47437);
and U48253 (N_48253,N_47555,N_47721);
xnor U48254 (N_48254,N_47934,N_47355);
xnor U48255 (N_48255,N_47445,N_47571);
and U48256 (N_48256,N_47614,N_47189);
xor U48257 (N_48257,N_47663,N_47591);
nor U48258 (N_48258,N_47349,N_47665);
nor U48259 (N_48259,N_47745,N_47908);
nor U48260 (N_48260,N_47314,N_47874);
xor U48261 (N_48261,N_47450,N_47190);
and U48262 (N_48262,N_47821,N_47789);
or U48263 (N_48263,N_47478,N_47095);
nand U48264 (N_48264,N_47348,N_47185);
xnor U48265 (N_48265,N_47486,N_47687);
or U48266 (N_48266,N_47588,N_47597);
nand U48267 (N_48267,N_47859,N_47256);
and U48268 (N_48268,N_47431,N_47595);
nor U48269 (N_48269,N_47270,N_47563);
and U48270 (N_48270,N_47632,N_47113);
nor U48271 (N_48271,N_47465,N_47990);
or U48272 (N_48272,N_47066,N_47051);
nand U48273 (N_48273,N_47511,N_47733);
nor U48274 (N_48274,N_47961,N_47223);
nand U48275 (N_48275,N_47678,N_47993);
and U48276 (N_48276,N_47202,N_47474);
and U48277 (N_48277,N_47593,N_47467);
nand U48278 (N_48278,N_47459,N_47233);
nor U48279 (N_48279,N_47180,N_47723);
nand U48280 (N_48280,N_47211,N_47213);
or U48281 (N_48281,N_47366,N_47341);
nor U48282 (N_48282,N_47788,N_47438);
nor U48283 (N_48283,N_47989,N_47247);
nand U48284 (N_48284,N_47512,N_47155);
nand U48285 (N_48285,N_47749,N_47620);
nand U48286 (N_48286,N_47339,N_47696);
nand U48287 (N_48287,N_47461,N_47131);
nand U48288 (N_48288,N_47561,N_47523);
nor U48289 (N_48289,N_47704,N_47542);
nor U48290 (N_48290,N_47049,N_47966);
nand U48291 (N_48291,N_47311,N_47184);
or U48292 (N_48292,N_47398,N_47703);
xnor U48293 (N_48293,N_47861,N_47200);
nor U48294 (N_48294,N_47217,N_47046);
nor U48295 (N_48295,N_47705,N_47809);
or U48296 (N_48296,N_47242,N_47216);
or U48297 (N_48297,N_47890,N_47293);
or U48298 (N_48298,N_47181,N_47829);
xnor U48299 (N_48299,N_47904,N_47699);
nor U48300 (N_48300,N_47653,N_47110);
nand U48301 (N_48301,N_47336,N_47329);
xnor U48302 (N_48302,N_47888,N_47161);
or U48303 (N_48303,N_47629,N_47403);
and U48304 (N_48304,N_47072,N_47433);
nand U48305 (N_48305,N_47201,N_47210);
or U48306 (N_48306,N_47167,N_47701);
nand U48307 (N_48307,N_47531,N_47841);
nor U48308 (N_48308,N_47776,N_47226);
nand U48309 (N_48309,N_47407,N_47949);
nor U48310 (N_48310,N_47514,N_47923);
and U48311 (N_48311,N_47322,N_47085);
or U48312 (N_48312,N_47375,N_47346);
nor U48313 (N_48313,N_47507,N_47138);
nor U48314 (N_48314,N_47554,N_47684);
xnor U48315 (N_48315,N_47306,N_47490);
and U48316 (N_48316,N_47017,N_47891);
nand U48317 (N_48317,N_47709,N_47267);
or U48318 (N_48318,N_47099,N_47725);
and U48319 (N_48319,N_47196,N_47613);
and U48320 (N_48320,N_47919,N_47470);
or U48321 (N_48321,N_47817,N_47522);
and U48322 (N_48322,N_47894,N_47229);
or U48323 (N_48323,N_47048,N_47565);
or U48324 (N_48324,N_47447,N_47088);
xnor U48325 (N_48325,N_47016,N_47802);
and U48326 (N_48326,N_47112,N_47504);
nor U48327 (N_48327,N_47837,N_47055);
or U48328 (N_48328,N_47770,N_47659);
or U48329 (N_48329,N_47301,N_47769);
and U48330 (N_48330,N_47857,N_47795);
or U48331 (N_48331,N_47911,N_47365);
xor U48332 (N_48332,N_47524,N_47805);
xnor U48333 (N_48333,N_47589,N_47126);
nor U48334 (N_48334,N_47122,N_47940);
or U48335 (N_48335,N_47917,N_47361);
and U48336 (N_48336,N_47207,N_47938);
or U48337 (N_48337,N_47238,N_47671);
nand U48338 (N_48338,N_47345,N_47950);
and U48339 (N_48339,N_47694,N_47735);
nand U48340 (N_48340,N_47087,N_47257);
and U48341 (N_48341,N_47777,N_47234);
nand U48342 (N_48342,N_47038,N_47994);
nor U48343 (N_48343,N_47194,N_47669);
nor U48344 (N_48344,N_47965,N_47627);
nor U48345 (N_48345,N_47362,N_47010);
or U48346 (N_48346,N_47845,N_47441);
or U48347 (N_48347,N_47985,N_47668);
xor U48348 (N_48348,N_47509,N_47757);
nor U48349 (N_48349,N_47970,N_47303);
nand U48350 (N_48350,N_47079,N_47367);
xnor U48351 (N_48351,N_47244,N_47160);
or U48352 (N_48352,N_47801,N_47421);
xnor U48353 (N_48353,N_47513,N_47872);
and U48354 (N_48354,N_47041,N_47396);
or U48355 (N_48355,N_47644,N_47397);
nand U48356 (N_48356,N_47393,N_47592);
xor U48357 (N_48357,N_47630,N_47489);
and U48358 (N_48358,N_47679,N_47832);
nand U48359 (N_48359,N_47477,N_47734);
nor U48360 (N_48360,N_47685,N_47291);
xnor U48361 (N_48361,N_47473,N_47500);
and U48362 (N_48362,N_47606,N_47218);
and U48363 (N_48363,N_47617,N_47006);
or U48364 (N_48364,N_47426,N_47285);
nor U48365 (N_48365,N_47607,N_47404);
and U48366 (N_48366,N_47615,N_47517);
xnor U48367 (N_48367,N_47480,N_47249);
nand U48368 (N_48368,N_47123,N_47824);
and U48369 (N_48369,N_47747,N_47742);
nand U48370 (N_48370,N_47712,N_47853);
and U48371 (N_48371,N_47173,N_47494);
nor U48372 (N_48372,N_47758,N_47235);
nand U48373 (N_48373,N_47428,N_47714);
and U48374 (N_48374,N_47879,N_47133);
or U48375 (N_48375,N_47502,N_47794);
or U48376 (N_48376,N_47377,N_47813);
or U48377 (N_48377,N_47353,N_47878);
or U48378 (N_48378,N_47638,N_47440);
or U48379 (N_48379,N_47001,N_47812);
nor U48380 (N_48380,N_47618,N_47423);
or U48381 (N_48381,N_47090,N_47581);
xnor U48382 (N_48382,N_47928,N_47021);
nor U48383 (N_48383,N_47761,N_47646);
xor U48384 (N_48384,N_47873,N_47012);
and U48385 (N_48385,N_47768,N_47316);
or U48386 (N_48386,N_47497,N_47357);
or U48387 (N_48387,N_47540,N_47360);
or U48388 (N_48388,N_47036,N_47278);
xnor U48389 (N_48389,N_47843,N_47906);
nand U48390 (N_48390,N_47498,N_47434);
xnor U48391 (N_48391,N_47737,N_47073);
or U48392 (N_48392,N_47231,N_47796);
and U48393 (N_48393,N_47148,N_47676);
xor U48394 (N_48394,N_47583,N_47815);
nand U48395 (N_48395,N_47102,N_47089);
or U48396 (N_48396,N_47227,N_47312);
and U48397 (N_48397,N_47527,N_47352);
nor U48398 (N_48398,N_47900,N_47534);
nand U48399 (N_48399,N_47157,N_47520);
nand U48400 (N_48400,N_47239,N_47992);
nor U48401 (N_48401,N_47009,N_47932);
or U48402 (N_48402,N_47516,N_47378);
and U48403 (N_48403,N_47030,N_47974);
xor U48404 (N_48404,N_47732,N_47718);
and U48405 (N_48405,N_47952,N_47759);
nand U48406 (N_48406,N_47418,N_47688);
or U48407 (N_48407,N_47295,N_47208);
and U48408 (N_48408,N_47383,N_47526);
nand U48409 (N_48409,N_47622,N_47537);
xnor U48410 (N_48410,N_47263,N_47014);
nand U48411 (N_48411,N_47508,N_47921);
nor U48412 (N_48412,N_47466,N_47411);
nor U48413 (N_48413,N_47539,N_47015);
xor U48414 (N_48414,N_47462,N_47692);
and U48415 (N_48415,N_47254,N_47912);
nand U48416 (N_48416,N_47317,N_47587);
nand U48417 (N_48417,N_47739,N_47729);
nor U48418 (N_48418,N_47300,N_47075);
and U48419 (N_48419,N_47356,N_47918);
nand U48420 (N_48420,N_47308,N_47412);
xor U48421 (N_48421,N_47519,N_47324);
nor U48422 (N_48422,N_47715,N_47838);
nand U48423 (N_48423,N_47491,N_47719);
xnor U48424 (N_48424,N_47453,N_47076);
nand U48425 (N_48425,N_47198,N_47634);
xnor U48426 (N_48426,N_47664,N_47600);
nor U48427 (N_48427,N_47656,N_47083);
nand U48428 (N_48428,N_47846,N_47955);
and U48429 (N_48429,N_47443,N_47372);
xor U48430 (N_48430,N_47851,N_47289);
nand U48431 (N_48431,N_47124,N_47258);
nand U48432 (N_48432,N_47981,N_47274);
or U48433 (N_48433,N_47973,N_47343);
or U48434 (N_48434,N_47023,N_47379);
xnor U48435 (N_48435,N_47471,N_47178);
or U48436 (N_48436,N_47080,N_47823);
nand U48437 (N_48437,N_47058,N_47639);
and U48438 (N_48438,N_47842,N_47232);
nor U48439 (N_48439,N_47045,N_47695);
nand U48440 (N_48440,N_47647,N_47186);
nand U48441 (N_48441,N_47071,N_47251);
and U48442 (N_48442,N_47680,N_47109);
nand U48443 (N_48443,N_47130,N_47783);
xor U48444 (N_48444,N_47182,N_47852);
nor U48445 (N_48445,N_47560,N_47922);
and U48446 (N_48446,N_47599,N_47941);
or U48447 (N_48447,N_47147,N_47697);
or U48448 (N_48448,N_47094,N_47763);
nor U48449 (N_48449,N_47986,N_47228);
and U48450 (N_48450,N_47991,N_47188);
nor U48451 (N_48451,N_47338,N_47682);
and U48452 (N_48452,N_47422,N_47569);
and U48453 (N_48453,N_47246,N_47401);
nor U48454 (N_48454,N_47142,N_47132);
xor U48455 (N_48455,N_47623,N_47115);
nand U48456 (N_48456,N_47128,N_47515);
or U48457 (N_48457,N_47492,N_47683);
or U48458 (N_48458,N_47025,N_47743);
or U48459 (N_48459,N_47771,N_47858);
or U48460 (N_48460,N_47221,N_47092);
and U48461 (N_48461,N_47175,N_47982);
nor U48462 (N_48462,N_47069,N_47212);
xor U48463 (N_48463,N_47171,N_47097);
nand U48464 (N_48464,N_47484,N_47720);
xnor U48465 (N_48465,N_47558,N_47305);
nand U48466 (N_48466,N_47549,N_47666);
nand U48467 (N_48467,N_47464,N_47276);
or U48468 (N_48468,N_47003,N_47047);
xnor U48469 (N_48469,N_47691,N_47892);
or U48470 (N_48470,N_47292,N_47408);
nand U48471 (N_48471,N_47387,N_47374);
or U48472 (N_48472,N_47624,N_47762);
nor U48473 (N_48473,N_47334,N_47280);
nand U48474 (N_48474,N_47499,N_47799);
and U48475 (N_48475,N_47446,N_47943);
or U48476 (N_48476,N_47463,N_47567);
nand U48477 (N_48477,N_47584,N_47548);
nand U48478 (N_48478,N_47806,N_47164);
or U48479 (N_48479,N_47354,N_47011);
nand U48480 (N_48480,N_47177,N_47738);
nand U48481 (N_48481,N_47827,N_47002);
and U48482 (N_48482,N_47309,N_47283);
xor U48483 (N_48483,N_47909,N_47518);
or U48484 (N_48484,N_47864,N_47252);
and U48485 (N_48485,N_47640,N_47916);
xnor U48486 (N_48486,N_47039,N_47448);
and U48487 (N_48487,N_47452,N_47532);
nor U48488 (N_48488,N_47417,N_47797);
and U48489 (N_48489,N_47019,N_47230);
xor U48490 (N_48490,N_47610,N_47927);
and U48491 (N_48491,N_47121,N_47427);
or U48492 (N_48492,N_47713,N_47553);
nor U48493 (N_48493,N_47793,N_47120);
or U48494 (N_48494,N_47636,N_47962);
and U48495 (N_48495,N_47145,N_47245);
nand U48496 (N_48496,N_47731,N_47867);
and U48497 (N_48497,N_47388,N_47641);
or U48498 (N_48498,N_47347,N_47342);
or U48499 (N_48499,N_47849,N_47924);
xor U48500 (N_48500,N_47876,N_47584);
nor U48501 (N_48501,N_47146,N_47957);
xor U48502 (N_48502,N_47051,N_47722);
nand U48503 (N_48503,N_47213,N_47931);
nor U48504 (N_48504,N_47037,N_47853);
nand U48505 (N_48505,N_47272,N_47632);
and U48506 (N_48506,N_47268,N_47755);
nand U48507 (N_48507,N_47660,N_47722);
or U48508 (N_48508,N_47059,N_47947);
xnor U48509 (N_48509,N_47938,N_47162);
or U48510 (N_48510,N_47353,N_47490);
or U48511 (N_48511,N_47321,N_47382);
xnor U48512 (N_48512,N_47654,N_47780);
and U48513 (N_48513,N_47509,N_47665);
or U48514 (N_48514,N_47681,N_47840);
nor U48515 (N_48515,N_47348,N_47186);
nor U48516 (N_48516,N_47160,N_47983);
nand U48517 (N_48517,N_47375,N_47612);
and U48518 (N_48518,N_47379,N_47670);
nand U48519 (N_48519,N_47546,N_47235);
or U48520 (N_48520,N_47048,N_47385);
xnor U48521 (N_48521,N_47437,N_47350);
xor U48522 (N_48522,N_47723,N_47051);
nand U48523 (N_48523,N_47067,N_47839);
nand U48524 (N_48524,N_47053,N_47850);
nand U48525 (N_48525,N_47177,N_47215);
xnor U48526 (N_48526,N_47640,N_47645);
xor U48527 (N_48527,N_47141,N_47322);
nor U48528 (N_48528,N_47927,N_47954);
nor U48529 (N_48529,N_47527,N_47019);
and U48530 (N_48530,N_47354,N_47605);
or U48531 (N_48531,N_47957,N_47785);
or U48532 (N_48532,N_47912,N_47163);
nor U48533 (N_48533,N_47888,N_47518);
nand U48534 (N_48534,N_47399,N_47973);
nand U48535 (N_48535,N_47470,N_47454);
and U48536 (N_48536,N_47631,N_47273);
nor U48537 (N_48537,N_47440,N_47022);
xnor U48538 (N_48538,N_47549,N_47853);
and U48539 (N_48539,N_47715,N_47474);
or U48540 (N_48540,N_47679,N_47248);
nor U48541 (N_48541,N_47660,N_47552);
nor U48542 (N_48542,N_47607,N_47667);
or U48543 (N_48543,N_47563,N_47392);
nand U48544 (N_48544,N_47231,N_47554);
and U48545 (N_48545,N_47348,N_47875);
nor U48546 (N_48546,N_47036,N_47439);
and U48547 (N_48547,N_47130,N_47407);
nand U48548 (N_48548,N_47529,N_47704);
nor U48549 (N_48549,N_47193,N_47340);
nor U48550 (N_48550,N_47333,N_47236);
or U48551 (N_48551,N_47087,N_47640);
and U48552 (N_48552,N_47630,N_47063);
xnor U48553 (N_48553,N_47238,N_47945);
nand U48554 (N_48554,N_47060,N_47886);
xor U48555 (N_48555,N_47730,N_47572);
and U48556 (N_48556,N_47916,N_47410);
or U48557 (N_48557,N_47778,N_47814);
nand U48558 (N_48558,N_47937,N_47439);
and U48559 (N_48559,N_47253,N_47180);
or U48560 (N_48560,N_47192,N_47620);
nand U48561 (N_48561,N_47313,N_47879);
nand U48562 (N_48562,N_47938,N_47044);
or U48563 (N_48563,N_47300,N_47859);
and U48564 (N_48564,N_47765,N_47917);
nand U48565 (N_48565,N_47790,N_47709);
and U48566 (N_48566,N_47025,N_47788);
nor U48567 (N_48567,N_47423,N_47519);
or U48568 (N_48568,N_47211,N_47919);
and U48569 (N_48569,N_47568,N_47837);
xnor U48570 (N_48570,N_47251,N_47977);
xnor U48571 (N_48571,N_47745,N_47089);
nor U48572 (N_48572,N_47988,N_47595);
xor U48573 (N_48573,N_47059,N_47602);
xor U48574 (N_48574,N_47037,N_47424);
or U48575 (N_48575,N_47883,N_47727);
xor U48576 (N_48576,N_47260,N_47442);
or U48577 (N_48577,N_47822,N_47764);
xnor U48578 (N_48578,N_47447,N_47952);
xor U48579 (N_48579,N_47171,N_47008);
and U48580 (N_48580,N_47326,N_47015);
nand U48581 (N_48581,N_47746,N_47591);
or U48582 (N_48582,N_47810,N_47788);
nand U48583 (N_48583,N_47145,N_47491);
or U48584 (N_48584,N_47453,N_47409);
and U48585 (N_48585,N_47985,N_47052);
or U48586 (N_48586,N_47789,N_47260);
or U48587 (N_48587,N_47556,N_47499);
or U48588 (N_48588,N_47809,N_47432);
xnor U48589 (N_48589,N_47042,N_47940);
or U48590 (N_48590,N_47482,N_47346);
nor U48591 (N_48591,N_47042,N_47192);
nand U48592 (N_48592,N_47541,N_47044);
or U48593 (N_48593,N_47740,N_47161);
or U48594 (N_48594,N_47961,N_47789);
nand U48595 (N_48595,N_47498,N_47970);
or U48596 (N_48596,N_47534,N_47783);
nand U48597 (N_48597,N_47925,N_47769);
and U48598 (N_48598,N_47588,N_47101);
and U48599 (N_48599,N_47851,N_47797);
xnor U48600 (N_48600,N_47078,N_47474);
nor U48601 (N_48601,N_47254,N_47444);
and U48602 (N_48602,N_47500,N_47660);
nor U48603 (N_48603,N_47913,N_47562);
and U48604 (N_48604,N_47721,N_47413);
xor U48605 (N_48605,N_47433,N_47181);
nand U48606 (N_48606,N_47594,N_47887);
or U48607 (N_48607,N_47742,N_47637);
nor U48608 (N_48608,N_47623,N_47638);
xnor U48609 (N_48609,N_47272,N_47890);
xnor U48610 (N_48610,N_47768,N_47279);
nand U48611 (N_48611,N_47746,N_47216);
xor U48612 (N_48612,N_47433,N_47359);
and U48613 (N_48613,N_47716,N_47277);
or U48614 (N_48614,N_47796,N_47950);
or U48615 (N_48615,N_47538,N_47758);
nand U48616 (N_48616,N_47164,N_47246);
nand U48617 (N_48617,N_47816,N_47129);
nor U48618 (N_48618,N_47844,N_47222);
or U48619 (N_48619,N_47326,N_47994);
xnor U48620 (N_48620,N_47898,N_47770);
xor U48621 (N_48621,N_47491,N_47840);
nor U48622 (N_48622,N_47334,N_47516);
or U48623 (N_48623,N_47629,N_47195);
xnor U48624 (N_48624,N_47004,N_47006);
xor U48625 (N_48625,N_47014,N_47503);
and U48626 (N_48626,N_47580,N_47454);
nand U48627 (N_48627,N_47746,N_47683);
nand U48628 (N_48628,N_47893,N_47925);
nor U48629 (N_48629,N_47558,N_47750);
nor U48630 (N_48630,N_47632,N_47867);
nor U48631 (N_48631,N_47061,N_47477);
nor U48632 (N_48632,N_47068,N_47121);
xor U48633 (N_48633,N_47577,N_47045);
nand U48634 (N_48634,N_47088,N_47744);
xor U48635 (N_48635,N_47282,N_47219);
nand U48636 (N_48636,N_47352,N_47248);
and U48637 (N_48637,N_47280,N_47808);
and U48638 (N_48638,N_47369,N_47323);
and U48639 (N_48639,N_47958,N_47148);
or U48640 (N_48640,N_47814,N_47015);
xnor U48641 (N_48641,N_47953,N_47762);
nand U48642 (N_48642,N_47625,N_47808);
and U48643 (N_48643,N_47712,N_47161);
nor U48644 (N_48644,N_47918,N_47360);
xnor U48645 (N_48645,N_47134,N_47054);
or U48646 (N_48646,N_47306,N_47090);
and U48647 (N_48647,N_47340,N_47960);
nand U48648 (N_48648,N_47700,N_47762);
or U48649 (N_48649,N_47089,N_47237);
or U48650 (N_48650,N_47228,N_47725);
nor U48651 (N_48651,N_47271,N_47055);
nand U48652 (N_48652,N_47619,N_47360);
xor U48653 (N_48653,N_47087,N_47465);
xor U48654 (N_48654,N_47639,N_47811);
nand U48655 (N_48655,N_47947,N_47562);
or U48656 (N_48656,N_47008,N_47240);
xnor U48657 (N_48657,N_47231,N_47790);
and U48658 (N_48658,N_47714,N_47885);
xor U48659 (N_48659,N_47968,N_47371);
nand U48660 (N_48660,N_47748,N_47200);
or U48661 (N_48661,N_47578,N_47394);
xnor U48662 (N_48662,N_47947,N_47099);
nand U48663 (N_48663,N_47927,N_47525);
nor U48664 (N_48664,N_47662,N_47984);
nor U48665 (N_48665,N_47729,N_47304);
and U48666 (N_48666,N_47191,N_47823);
xnor U48667 (N_48667,N_47092,N_47526);
or U48668 (N_48668,N_47734,N_47697);
and U48669 (N_48669,N_47482,N_47144);
or U48670 (N_48670,N_47802,N_47499);
or U48671 (N_48671,N_47392,N_47564);
xnor U48672 (N_48672,N_47718,N_47658);
or U48673 (N_48673,N_47307,N_47531);
nand U48674 (N_48674,N_47899,N_47711);
and U48675 (N_48675,N_47799,N_47276);
and U48676 (N_48676,N_47071,N_47833);
xor U48677 (N_48677,N_47504,N_47256);
or U48678 (N_48678,N_47559,N_47202);
nor U48679 (N_48679,N_47267,N_47823);
xor U48680 (N_48680,N_47823,N_47007);
nor U48681 (N_48681,N_47081,N_47019);
nand U48682 (N_48682,N_47998,N_47613);
or U48683 (N_48683,N_47232,N_47807);
and U48684 (N_48684,N_47962,N_47061);
or U48685 (N_48685,N_47366,N_47888);
or U48686 (N_48686,N_47075,N_47650);
xnor U48687 (N_48687,N_47655,N_47287);
and U48688 (N_48688,N_47972,N_47822);
nand U48689 (N_48689,N_47506,N_47612);
nor U48690 (N_48690,N_47885,N_47673);
nand U48691 (N_48691,N_47350,N_47214);
and U48692 (N_48692,N_47547,N_47687);
and U48693 (N_48693,N_47134,N_47664);
xnor U48694 (N_48694,N_47830,N_47614);
xnor U48695 (N_48695,N_47907,N_47594);
or U48696 (N_48696,N_47133,N_47642);
nand U48697 (N_48697,N_47925,N_47785);
and U48698 (N_48698,N_47892,N_47373);
nor U48699 (N_48699,N_47308,N_47365);
nand U48700 (N_48700,N_47805,N_47569);
xnor U48701 (N_48701,N_47364,N_47340);
or U48702 (N_48702,N_47469,N_47336);
xor U48703 (N_48703,N_47721,N_47248);
nor U48704 (N_48704,N_47116,N_47498);
xor U48705 (N_48705,N_47898,N_47552);
and U48706 (N_48706,N_47637,N_47644);
or U48707 (N_48707,N_47899,N_47560);
and U48708 (N_48708,N_47335,N_47080);
and U48709 (N_48709,N_47703,N_47540);
and U48710 (N_48710,N_47269,N_47485);
or U48711 (N_48711,N_47820,N_47346);
or U48712 (N_48712,N_47286,N_47917);
or U48713 (N_48713,N_47515,N_47402);
nand U48714 (N_48714,N_47651,N_47663);
nor U48715 (N_48715,N_47356,N_47282);
nor U48716 (N_48716,N_47446,N_47684);
xnor U48717 (N_48717,N_47941,N_47479);
xor U48718 (N_48718,N_47088,N_47406);
nand U48719 (N_48719,N_47715,N_47926);
or U48720 (N_48720,N_47450,N_47779);
or U48721 (N_48721,N_47798,N_47552);
xor U48722 (N_48722,N_47660,N_47134);
and U48723 (N_48723,N_47942,N_47951);
nand U48724 (N_48724,N_47935,N_47694);
and U48725 (N_48725,N_47760,N_47740);
and U48726 (N_48726,N_47328,N_47556);
nor U48727 (N_48727,N_47837,N_47954);
nor U48728 (N_48728,N_47795,N_47701);
or U48729 (N_48729,N_47386,N_47297);
or U48730 (N_48730,N_47138,N_47961);
xnor U48731 (N_48731,N_47238,N_47021);
nand U48732 (N_48732,N_47848,N_47414);
nand U48733 (N_48733,N_47757,N_47324);
nand U48734 (N_48734,N_47960,N_47949);
xnor U48735 (N_48735,N_47198,N_47192);
nand U48736 (N_48736,N_47006,N_47048);
nor U48737 (N_48737,N_47074,N_47323);
or U48738 (N_48738,N_47030,N_47363);
nand U48739 (N_48739,N_47380,N_47611);
and U48740 (N_48740,N_47821,N_47849);
or U48741 (N_48741,N_47554,N_47278);
and U48742 (N_48742,N_47320,N_47934);
nand U48743 (N_48743,N_47659,N_47894);
and U48744 (N_48744,N_47802,N_47692);
or U48745 (N_48745,N_47489,N_47521);
or U48746 (N_48746,N_47478,N_47027);
nor U48747 (N_48747,N_47615,N_47232);
nor U48748 (N_48748,N_47312,N_47037);
nor U48749 (N_48749,N_47161,N_47237);
or U48750 (N_48750,N_47137,N_47674);
and U48751 (N_48751,N_47722,N_47023);
and U48752 (N_48752,N_47691,N_47640);
xnor U48753 (N_48753,N_47471,N_47139);
and U48754 (N_48754,N_47078,N_47414);
xor U48755 (N_48755,N_47673,N_47419);
nand U48756 (N_48756,N_47029,N_47777);
xor U48757 (N_48757,N_47770,N_47540);
nor U48758 (N_48758,N_47919,N_47019);
nand U48759 (N_48759,N_47552,N_47458);
xnor U48760 (N_48760,N_47763,N_47102);
nand U48761 (N_48761,N_47829,N_47186);
nand U48762 (N_48762,N_47483,N_47043);
and U48763 (N_48763,N_47267,N_47013);
nor U48764 (N_48764,N_47550,N_47440);
and U48765 (N_48765,N_47941,N_47143);
and U48766 (N_48766,N_47780,N_47465);
or U48767 (N_48767,N_47190,N_47849);
and U48768 (N_48768,N_47798,N_47238);
or U48769 (N_48769,N_47019,N_47696);
nand U48770 (N_48770,N_47510,N_47334);
and U48771 (N_48771,N_47841,N_47327);
and U48772 (N_48772,N_47543,N_47746);
or U48773 (N_48773,N_47701,N_47324);
nor U48774 (N_48774,N_47764,N_47123);
nor U48775 (N_48775,N_47788,N_47437);
xnor U48776 (N_48776,N_47305,N_47147);
xnor U48777 (N_48777,N_47201,N_47684);
or U48778 (N_48778,N_47336,N_47729);
and U48779 (N_48779,N_47751,N_47817);
nor U48780 (N_48780,N_47828,N_47588);
or U48781 (N_48781,N_47280,N_47555);
xor U48782 (N_48782,N_47397,N_47409);
and U48783 (N_48783,N_47328,N_47609);
nand U48784 (N_48784,N_47892,N_47698);
nand U48785 (N_48785,N_47443,N_47304);
and U48786 (N_48786,N_47422,N_47405);
xnor U48787 (N_48787,N_47328,N_47917);
or U48788 (N_48788,N_47148,N_47014);
nand U48789 (N_48789,N_47704,N_47624);
nor U48790 (N_48790,N_47608,N_47810);
and U48791 (N_48791,N_47576,N_47842);
or U48792 (N_48792,N_47267,N_47591);
xor U48793 (N_48793,N_47202,N_47640);
and U48794 (N_48794,N_47742,N_47649);
nand U48795 (N_48795,N_47297,N_47923);
and U48796 (N_48796,N_47044,N_47260);
xor U48797 (N_48797,N_47340,N_47445);
xnor U48798 (N_48798,N_47091,N_47146);
xor U48799 (N_48799,N_47983,N_47237);
xor U48800 (N_48800,N_47239,N_47588);
and U48801 (N_48801,N_47439,N_47887);
nand U48802 (N_48802,N_47203,N_47082);
and U48803 (N_48803,N_47485,N_47728);
nand U48804 (N_48804,N_47617,N_47162);
and U48805 (N_48805,N_47417,N_47843);
and U48806 (N_48806,N_47506,N_47564);
xnor U48807 (N_48807,N_47742,N_47893);
and U48808 (N_48808,N_47874,N_47891);
and U48809 (N_48809,N_47653,N_47507);
nand U48810 (N_48810,N_47776,N_47173);
xnor U48811 (N_48811,N_47977,N_47327);
or U48812 (N_48812,N_47305,N_47859);
nand U48813 (N_48813,N_47935,N_47879);
and U48814 (N_48814,N_47284,N_47733);
xor U48815 (N_48815,N_47248,N_47908);
nor U48816 (N_48816,N_47353,N_47441);
nand U48817 (N_48817,N_47141,N_47154);
xor U48818 (N_48818,N_47189,N_47092);
or U48819 (N_48819,N_47234,N_47850);
and U48820 (N_48820,N_47011,N_47704);
xor U48821 (N_48821,N_47434,N_47443);
xor U48822 (N_48822,N_47646,N_47801);
xnor U48823 (N_48823,N_47992,N_47728);
nor U48824 (N_48824,N_47685,N_47694);
nand U48825 (N_48825,N_47634,N_47511);
nor U48826 (N_48826,N_47620,N_47627);
nor U48827 (N_48827,N_47690,N_47279);
and U48828 (N_48828,N_47460,N_47480);
or U48829 (N_48829,N_47317,N_47951);
nor U48830 (N_48830,N_47423,N_47736);
nor U48831 (N_48831,N_47629,N_47140);
nand U48832 (N_48832,N_47384,N_47968);
or U48833 (N_48833,N_47940,N_47864);
and U48834 (N_48834,N_47305,N_47942);
xor U48835 (N_48835,N_47190,N_47029);
xor U48836 (N_48836,N_47937,N_47409);
nand U48837 (N_48837,N_47317,N_47984);
or U48838 (N_48838,N_47729,N_47560);
or U48839 (N_48839,N_47680,N_47116);
and U48840 (N_48840,N_47093,N_47983);
or U48841 (N_48841,N_47619,N_47082);
xor U48842 (N_48842,N_47418,N_47643);
nand U48843 (N_48843,N_47598,N_47449);
nand U48844 (N_48844,N_47490,N_47497);
xnor U48845 (N_48845,N_47485,N_47661);
or U48846 (N_48846,N_47761,N_47470);
or U48847 (N_48847,N_47732,N_47576);
nor U48848 (N_48848,N_47353,N_47447);
nand U48849 (N_48849,N_47432,N_47837);
nand U48850 (N_48850,N_47115,N_47468);
nand U48851 (N_48851,N_47988,N_47513);
xnor U48852 (N_48852,N_47274,N_47878);
or U48853 (N_48853,N_47699,N_47935);
and U48854 (N_48854,N_47010,N_47024);
and U48855 (N_48855,N_47993,N_47423);
nand U48856 (N_48856,N_47827,N_47985);
and U48857 (N_48857,N_47419,N_47726);
or U48858 (N_48858,N_47593,N_47649);
nand U48859 (N_48859,N_47125,N_47547);
or U48860 (N_48860,N_47337,N_47996);
nor U48861 (N_48861,N_47423,N_47335);
and U48862 (N_48862,N_47888,N_47769);
xnor U48863 (N_48863,N_47771,N_47015);
and U48864 (N_48864,N_47245,N_47891);
and U48865 (N_48865,N_47900,N_47671);
xnor U48866 (N_48866,N_47519,N_47934);
nand U48867 (N_48867,N_47895,N_47653);
nand U48868 (N_48868,N_47574,N_47810);
nand U48869 (N_48869,N_47056,N_47595);
nand U48870 (N_48870,N_47285,N_47590);
or U48871 (N_48871,N_47761,N_47251);
nand U48872 (N_48872,N_47838,N_47320);
xnor U48873 (N_48873,N_47073,N_47691);
and U48874 (N_48874,N_47360,N_47268);
and U48875 (N_48875,N_47596,N_47183);
xnor U48876 (N_48876,N_47577,N_47807);
nand U48877 (N_48877,N_47612,N_47752);
nand U48878 (N_48878,N_47566,N_47244);
nand U48879 (N_48879,N_47310,N_47584);
and U48880 (N_48880,N_47363,N_47744);
or U48881 (N_48881,N_47445,N_47353);
and U48882 (N_48882,N_47046,N_47989);
or U48883 (N_48883,N_47603,N_47507);
nand U48884 (N_48884,N_47545,N_47719);
or U48885 (N_48885,N_47336,N_47697);
nand U48886 (N_48886,N_47143,N_47580);
xor U48887 (N_48887,N_47226,N_47174);
or U48888 (N_48888,N_47684,N_47644);
nand U48889 (N_48889,N_47026,N_47507);
and U48890 (N_48890,N_47200,N_47236);
xnor U48891 (N_48891,N_47325,N_47099);
nand U48892 (N_48892,N_47583,N_47790);
nand U48893 (N_48893,N_47456,N_47166);
xnor U48894 (N_48894,N_47668,N_47784);
nor U48895 (N_48895,N_47067,N_47315);
nand U48896 (N_48896,N_47211,N_47000);
nor U48897 (N_48897,N_47941,N_47997);
xnor U48898 (N_48898,N_47158,N_47690);
xor U48899 (N_48899,N_47188,N_47829);
or U48900 (N_48900,N_47884,N_47515);
or U48901 (N_48901,N_47251,N_47168);
or U48902 (N_48902,N_47298,N_47173);
nand U48903 (N_48903,N_47390,N_47583);
nor U48904 (N_48904,N_47788,N_47762);
or U48905 (N_48905,N_47417,N_47616);
nor U48906 (N_48906,N_47751,N_47395);
xnor U48907 (N_48907,N_47097,N_47745);
and U48908 (N_48908,N_47572,N_47814);
xnor U48909 (N_48909,N_47180,N_47467);
nor U48910 (N_48910,N_47665,N_47942);
nand U48911 (N_48911,N_47616,N_47207);
or U48912 (N_48912,N_47508,N_47768);
or U48913 (N_48913,N_47890,N_47332);
xnor U48914 (N_48914,N_47400,N_47053);
xor U48915 (N_48915,N_47746,N_47086);
nand U48916 (N_48916,N_47541,N_47010);
xnor U48917 (N_48917,N_47402,N_47907);
nor U48918 (N_48918,N_47684,N_47418);
and U48919 (N_48919,N_47029,N_47982);
xor U48920 (N_48920,N_47021,N_47948);
or U48921 (N_48921,N_47317,N_47545);
nor U48922 (N_48922,N_47829,N_47396);
nor U48923 (N_48923,N_47443,N_47973);
xnor U48924 (N_48924,N_47458,N_47759);
and U48925 (N_48925,N_47169,N_47657);
and U48926 (N_48926,N_47957,N_47499);
and U48927 (N_48927,N_47931,N_47109);
nand U48928 (N_48928,N_47304,N_47528);
nand U48929 (N_48929,N_47683,N_47778);
or U48930 (N_48930,N_47190,N_47875);
xnor U48931 (N_48931,N_47173,N_47998);
or U48932 (N_48932,N_47603,N_47803);
nand U48933 (N_48933,N_47991,N_47247);
xor U48934 (N_48934,N_47975,N_47918);
nor U48935 (N_48935,N_47727,N_47533);
or U48936 (N_48936,N_47139,N_47579);
nor U48937 (N_48937,N_47159,N_47228);
or U48938 (N_48938,N_47207,N_47987);
xor U48939 (N_48939,N_47736,N_47437);
xnor U48940 (N_48940,N_47517,N_47378);
nand U48941 (N_48941,N_47814,N_47618);
and U48942 (N_48942,N_47147,N_47856);
xor U48943 (N_48943,N_47396,N_47986);
nand U48944 (N_48944,N_47593,N_47474);
or U48945 (N_48945,N_47059,N_47052);
xnor U48946 (N_48946,N_47931,N_47424);
nand U48947 (N_48947,N_47511,N_47899);
and U48948 (N_48948,N_47325,N_47798);
nand U48949 (N_48949,N_47281,N_47792);
xnor U48950 (N_48950,N_47760,N_47094);
and U48951 (N_48951,N_47986,N_47757);
xor U48952 (N_48952,N_47549,N_47845);
and U48953 (N_48953,N_47140,N_47374);
nand U48954 (N_48954,N_47941,N_47008);
and U48955 (N_48955,N_47284,N_47690);
and U48956 (N_48956,N_47457,N_47629);
nand U48957 (N_48957,N_47867,N_47760);
xor U48958 (N_48958,N_47391,N_47323);
nor U48959 (N_48959,N_47347,N_47848);
nor U48960 (N_48960,N_47085,N_47880);
and U48961 (N_48961,N_47480,N_47428);
or U48962 (N_48962,N_47757,N_47447);
nor U48963 (N_48963,N_47512,N_47766);
nand U48964 (N_48964,N_47276,N_47632);
nand U48965 (N_48965,N_47631,N_47313);
nor U48966 (N_48966,N_47890,N_47719);
and U48967 (N_48967,N_47270,N_47455);
or U48968 (N_48968,N_47220,N_47303);
and U48969 (N_48969,N_47002,N_47205);
or U48970 (N_48970,N_47162,N_47653);
nand U48971 (N_48971,N_47726,N_47005);
nand U48972 (N_48972,N_47774,N_47889);
nand U48973 (N_48973,N_47251,N_47549);
or U48974 (N_48974,N_47366,N_47740);
nor U48975 (N_48975,N_47687,N_47491);
nand U48976 (N_48976,N_47220,N_47380);
nand U48977 (N_48977,N_47737,N_47411);
nand U48978 (N_48978,N_47283,N_47692);
nand U48979 (N_48979,N_47202,N_47778);
nand U48980 (N_48980,N_47868,N_47265);
or U48981 (N_48981,N_47916,N_47386);
xnor U48982 (N_48982,N_47848,N_47787);
nor U48983 (N_48983,N_47840,N_47021);
and U48984 (N_48984,N_47016,N_47442);
or U48985 (N_48985,N_47666,N_47330);
and U48986 (N_48986,N_47075,N_47383);
xor U48987 (N_48987,N_47257,N_47250);
xnor U48988 (N_48988,N_47985,N_47422);
and U48989 (N_48989,N_47092,N_47764);
or U48990 (N_48990,N_47120,N_47934);
or U48991 (N_48991,N_47013,N_47287);
xnor U48992 (N_48992,N_47518,N_47917);
nand U48993 (N_48993,N_47215,N_47340);
nor U48994 (N_48994,N_47689,N_47985);
nand U48995 (N_48995,N_47046,N_47711);
xor U48996 (N_48996,N_47470,N_47981);
or U48997 (N_48997,N_47799,N_47440);
and U48998 (N_48998,N_47755,N_47901);
and U48999 (N_48999,N_47562,N_47346);
and U49000 (N_49000,N_48673,N_48074);
or U49001 (N_49001,N_48776,N_48773);
xnor U49002 (N_49002,N_48784,N_48031);
or U49003 (N_49003,N_48957,N_48455);
or U49004 (N_49004,N_48215,N_48188);
xnor U49005 (N_49005,N_48449,N_48518);
xor U49006 (N_49006,N_48841,N_48242);
and U49007 (N_49007,N_48736,N_48321);
nor U49008 (N_49008,N_48436,N_48853);
nand U49009 (N_49009,N_48716,N_48207);
xnor U49010 (N_49010,N_48767,N_48503);
nor U49011 (N_49011,N_48501,N_48569);
nor U49012 (N_49012,N_48761,N_48221);
xnor U49013 (N_49013,N_48465,N_48828);
and U49014 (N_49014,N_48839,N_48912);
or U49015 (N_49015,N_48566,N_48932);
or U49016 (N_49016,N_48750,N_48661);
and U49017 (N_49017,N_48553,N_48804);
and U49018 (N_49018,N_48950,N_48026);
and U49019 (N_49019,N_48586,N_48641);
xor U49020 (N_49020,N_48140,N_48818);
xnor U49021 (N_49021,N_48005,N_48398);
or U49022 (N_49022,N_48241,N_48129);
nor U49023 (N_49023,N_48010,N_48835);
or U49024 (N_49024,N_48534,N_48210);
xnor U49025 (N_49025,N_48965,N_48459);
and U49026 (N_49026,N_48665,N_48970);
xnor U49027 (N_49027,N_48994,N_48992);
nand U49028 (N_49028,N_48190,N_48675);
or U49029 (N_49029,N_48380,N_48557);
nor U49030 (N_49030,N_48953,N_48947);
nand U49031 (N_49031,N_48682,N_48642);
or U49032 (N_49032,N_48173,N_48087);
nor U49033 (N_49033,N_48126,N_48464);
nand U49034 (N_49034,N_48332,N_48703);
and U49035 (N_49035,N_48421,N_48601);
xnor U49036 (N_49036,N_48561,N_48669);
nand U49037 (N_49037,N_48591,N_48892);
nand U49038 (N_49038,N_48516,N_48680);
and U49039 (N_49039,N_48089,N_48496);
nand U49040 (N_49040,N_48630,N_48610);
and U49041 (N_49041,N_48977,N_48709);
or U49042 (N_49042,N_48481,N_48741);
xor U49043 (N_49043,N_48753,N_48510);
or U49044 (N_49044,N_48695,N_48563);
nand U49045 (N_49045,N_48521,N_48280);
and U49046 (N_49046,N_48136,N_48824);
and U49047 (N_49047,N_48391,N_48420);
nand U49048 (N_49048,N_48158,N_48621);
nand U49049 (N_49049,N_48971,N_48823);
xor U49050 (N_49050,N_48806,N_48915);
or U49051 (N_49051,N_48989,N_48531);
and U49052 (N_49052,N_48628,N_48184);
nor U49053 (N_49053,N_48279,N_48663);
and U49054 (N_49054,N_48759,N_48727);
nand U49055 (N_49055,N_48133,N_48018);
or U49056 (N_49056,N_48228,N_48049);
and U49057 (N_49057,N_48497,N_48080);
xnor U49058 (N_49058,N_48577,N_48822);
or U49059 (N_49059,N_48118,N_48875);
nor U49060 (N_49060,N_48775,N_48615);
nor U49061 (N_49061,N_48012,N_48803);
xor U49062 (N_49062,N_48769,N_48523);
or U49063 (N_49063,N_48081,N_48282);
nor U49064 (N_49064,N_48402,N_48248);
nor U49065 (N_49065,N_48772,N_48019);
xor U49066 (N_49066,N_48124,N_48872);
or U49067 (N_49067,N_48612,N_48145);
nand U49068 (N_49068,N_48331,N_48346);
nor U49069 (N_49069,N_48528,N_48274);
nand U49070 (N_49070,N_48698,N_48293);
or U49071 (N_49071,N_48942,N_48052);
nor U49072 (N_49072,N_48762,N_48370);
and U49073 (N_49073,N_48424,N_48473);
nor U49074 (N_49074,N_48537,N_48379);
nand U49075 (N_49075,N_48798,N_48494);
and U49076 (N_49076,N_48737,N_48840);
and U49077 (N_49077,N_48177,N_48431);
and U49078 (N_49078,N_48690,N_48789);
nor U49079 (N_49079,N_48498,N_48482);
and U49080 (N_49080,N_48995,N_48653);
nand U49081 (N_49081,N_48434,N_48117);
nor U49082 (N_49082,N_48639,N_48832);
nor U49083 (N_49083,N_48194,N_48372);
xnor U49084 (N_49084,N_48713,N_48471);
and U49085 (N_49085,N_48991,N_48768);
and U49086 (N_49086,N_48352,N_48251);
or U49087 (N_49087,N_48134,N_48856);
nand U49088 (N_49088,N_48002,N_48000);
and U49089 (N_49089,N_48072,N_48966);
nor U49090 (N_49090,N_48351,N_48006);
or U49091 (N_49091,N_48978,N_48324);
and U49092 (N_49092,N_48618,N_48707);
or U49093 (N_49093,N_48038,N_48422);
nand U49094 (N_49094,N_48652,N_48842);
nor U49095 (N_49095,N_48908,N_48302);
xor U49096 (N_49096,N_48339,N_48606);
xor U49097 (N_49097,N_48760,N_48587);
nand U49098 (N_49098,N_48046,N_48148);
xor U49099 (N_49099,N_48743,N_48677);
nor U49100 (N_49100,N_48114,N_48972);
nand U49101 (N_49101,N_48342,N_48616);
and U49102 (N_49102,N_48224,N_48524);
and U49103 (N_49103,N_48595,N_48020);
nor U49104 (N_49104,N_48440,N_48530);
or U49105 (N_49105,N_48156,N_48259);
xor U49106 (N_49106,N_48968,N_48325);
nand U49107 (N_49107,N_48462,N_48163);
xnor U49108 (N_49108,N_48594,N_48644);
nand U49109 (N_49109,N_48917,N_48260);
nand U49110 (N_49110,N_48113,N_48122);
xnor U49111 (N_49111,N_48726,N_48626);
or U49112 (N_49112,N_48137,N_48104);
nor U49113 (N_49113,N_48419,N_48394);
xnor U49114 (N_49114,N_48547,N_48106);
nand U49115 (N_49115,N_48799,N_48416);
xor U49116 (N_49116,N_48714,N_48738);
and U49117 (N_49117,N_48880,N_48252);
nand U49118 (N_49118,N_48959,N_48763);
or U49119 (N_49119,N_48167,N_48627);
nand U49120 (N_49120,N_48231,N_48893);
or U49121 (N_49121,N_48801,N_48890);
xor U49122 (N_49122,N_48958,N_48410);
or U49123 (N_49123,N_48024,N_48648);
nand U49124 (N_49124,N_48405,N_48624);
nand U49125 (N_49125,N_48904,N_48474);
or U49126 (N_49126,N_48825,N_48884);
nor U49127 (N_49127,N_48838,N_48082);
nand U49128 (N_49128,N_48802,N_48583);
xnor U49129 (N_49129,N_48862,N_48445);
nor U49130 (N_49130,N_48375,N_48740);
nand U49131 (N_49131,N_48461,N_48334);
and U49132 (N_49132,N_48197,N_48388);
or U49133 (N_49133,N_48152,N_48895);
xnor U49134 (N_49134,N_48281,N_48907);
or U49135 (N_49135,N_48559,N_48437);
and U49136 (N_49136,N_48429,N_48797);
xnor U49137 (N_49137,N_48830,N_48902);
nor U49138 (N_49138,N_48415,N_48899);
xor U49139 (N_49139,N_48980,N_48732);
nand U49140 (N_49140,N_48666,N_48460);
and U49141 (N_49141,N_48373,N_48597);
xor U49142 (N_49142,N_48257,N_48165);
nand U49143 (N_49143,N_48285,N_48751);
nor U49144 (N_49144,N_48452,N_48887);
and U49145 (N_49145,N_48358,N_48288);
or U49146 (N_49146,N_48312,N_48993);
or U49147 (N_49147,N_48724,N_48418);
or U49148 (N_49148,N_48131,N_48094);
and U49149 (N_49149,N_48655,N_48670);
nand U49150 (N_49150,N_48335,N_48463);
and U49151 (N_49151,N_48812,N_48034);
or U49152 (N_49152,N_48403,N_48593);
nand U49153 (N_49153,N_48084,N_48647);
nand U49154 (N_49154,N_48159,N_48196);
or U49155 (N_49155,N_48349,N_48969);
nor U49156 (N_49156,N_48790,N_48039);
nor U49157 (N_49157,N_48320,N_48023);
nand U49158 (N_49158,N_48105,N_48264);
and U49159 (N_49159,N_48044,N_48064);
nor U49160 (N_49160,N_48683,N_48693);
xnor U49161 (N_49161,N_48393,N_48008);
nor U49162 (N_49162,N_48668,N_48217);
nor U49163 (N_49163,N_48088,N_48042);
xor U49164 (N_49164,N_48142,N_48292);
nor U49165 (N_49165,N_48674,N_48045);
or U49166 (N_49166,N_48934,N_48585);
nand U49167 (N_49167,N_48700,N_48870);
and U49168 (N_49168,N_48232,N_48141);
xor U49169 (N_49169,N_48174,N_48780);
xor U49170 (N_49170,N_48720,N_48658);
or U49171 (N_49171,N_48651,N_48356);
and U49172 (N_49172,N_48679,N_48913);
and U49173 (N_49173,N_48108,N_48843);
nor U49174 (N_49174,N_48861,N_48121);
xnor U49175 (N_49175,N_48392,N_48879);
nand U49176 (N_49176,N_48604,N_48643);
or U49177 (N_49177,N_48598,N_48846);
nor U49178 (N_49178,N_48466,N_48502);
or U49179 (N_49179,N_48886,N_48395);
xor U49180 (N_49180,N_48238,N_48589);
or U49181 (N_49181,N_48574,N_48314);
nand U49182 (N_49182,N_48013,N_48535);
or U49183 (N_49183,N_48611,N_48213);
nor U49184 (N_49184,N_48036,N_48287);
xnor U49185 (N_49185,N_48381,N_48514);
nand U49186 (N_49186,N_48564,N_48764);
xnor U49187 (N_49187,N_48386,N_48809);
nand U49188 (N_49188,N_48273,N_48997);
nand U49189 (N_49189,N_48929,N_48849);
and U49190 (N_49190,N_48945,N_48428);
xnor U49191 (N_49191,N_48729,N_48245);
and U49192 (N_49192,N_48077,N_48278);
nor U49193 (N_49193,N_48816,N_48291);
or U49194 (N_49194,N_48580,N_48027);
and U49195 (N_49195,N_48609,N_48526);
or U49196 (N_49196,N_48244,N_48891);
and U49197 (N_49197,N_48781,N_48341);
and U49198 (N_49198,N_48927,N_48329);
or U49199 (N_49199,N_48065,N_48962);
or U49200 (N_49200,N_48536,N_48191);
or U49201 (N_49201,N_48284,N_48485);
nor U49202 (N_49202,N_48901,N_48817);
nand U49203 (N_49203,N_48542,N_48691);
xor U49204 (N_49204,N_48607,N_48914);
nand U49205 (N_49205,N_48617,N_48227);
and U49206 (N_49206,N_48130,N_48963);
and U49207 (N_49207,N_48718,N_48638);
xnor U49208 (N_49208,N_48376,N_48169);
nor U49209 (N_49209,N_48059,N_48304);
xnor U49210 (N_49210,N_48230,N_48692);
xor U49211 (N_49211,N_48337,N_48425);
xor U49212 (N_49212,N_48488,N_48990);
nand U49213 (N_49213,N_48295,N_48988);
nand U49214 (N_49214,N_48097,N_48246);
xnor U49215 (N_49215,N_48722,N_48359);
nand U49216 (N_49216,N_48694,N_48579);
and U49217 (N_49217,N_48378,N_48888);
or U49218 (N_49218,N_48400,N_48176);
nor U49219 (N_49219,N_48066,N_48101);
xor U49220 (N_49220,N_48125,N_48505);
nor U49221 (N_49221,N_48486,N_48664);
or U49222 (N_49222,N_48258,N_48814);
nor U49223 (N_49223,N_48366,N_48330);
and U49224 (N_49224,N_48793,N_48941);
nand U49225 (N_49225,N_48863,N_48795);
nand U49226 (N_49226,N_48930,N_48900);
and U49227 (N_49227,N_48057,N_48786);
nand U49228 (N_49228,N_48571,N_48556);
and U49229 (N_49229,N_48353,N_48877);
and U49230 (N_49230,N_48476,N_48864);
or U49231 (N_49231,N_48413,N_48656);
nand U49232 (N_49232,N_48596,N_48640);
or U49233 (N_49233,N_48964,N_48175);
nand U49234 (N_49234,N_48361,N_48149);
nand U49235 (N_49235,N_48202,N_48570);
nand U49236 (N_49236,N_48983,N_48735);
nor U49237 (N_49237,N_48987,N_48662);
or U49238 (N_49238,N_48225,N_48960);
nand U49239 (N_49239,N_48622,N_48578);
xnor U49240 (N_49240,N_48456,N_48549);
and U49241 (N_49241,N_48671,N_48322);
nand U49242 (N_49242,N_48371,N_48483);
nand U49243 (N_49243,N_48834,N_48198);
and U49244 (N_49244,N_48103,N_48233);
and U49245 (N_49245,N_48676,N_48432);
or U49246 (N_49246,N_48286,N_48948);
or U49247 (N_49247,N_48602,N_48389);
or U49248 (N_49248,N_48178,N_48756);
nor U49249 (N_49249,N_48717,N_48056);
or U49250 (N_49250,N_48266,N_48766);
xnor U49251 (N_49251,N_48973,N_48078);
nand U49252 (N_49252,N_48397,N_48406);
and U49253 (N_49253,N_48147,N_48015);
nand U49254 (N_49254,N_48447,N_48811);
nor U49255 (N_49255,N_48300,N_48146);
xor U49256 (N_49256,N_48928,N_48851);
and U49257 (N_49257,N_48116,N_48755);
and U49258 (N_49258,N_48697,N_48193);
nand U49259 (N_49259,N_48200,N_48299);
or U49260 (N_49260,N_48385,N_48268);
nor U49261 (N_49261,N_48778,N_48099);
nor U49262 (N_49262,N_48032,N_48276);
nand U49263 (N_49263,N_48792,N_48565);
or U49264 (N_49264,N_48199,N_48060);
and U49265 (N_49265,N_48527,N_48477);
and U49266 (N_49266,N_48180,N_48409);
nand U49267 (N_49267,N_48603,N_48954);
or U49268 (N_49268,N_48310,N_48272);
and U49269 (N_49269,N_48367,N_48047);
and U49270 (N_49270,N_48508,N_48368);
or U49271 (N_49271,N_48939,N_48007);
or U49272 (N_49272,N_48765,N_48926);
xnor U49273 (N_49273,N_48438,N_48430);
and U49274 (N_49274,N_48777,N_48667);
nand U49275 (N_49275,N_48984,N_48747);
nor U49276 (N_49276,N_48857,N_48127);
or U49277 (N_49277,N_48532,N_48634);
nand U49278 (N_49278,N_48450,N_48160);
or U49279 (N_49279,N_48029,N_48555);
xor U49280 (N_49280,N_48519,N_48728);
and U49281 (N_49281,N_48572,N_48195);
nor U49282 (N_49282,N_48319,N_48710);
or U49283 (N_49283,N_48889,N_48135);
and U49284 (N_49284,N_48701,N_48263);
or U49285 (N_49285,N_48216,N_48115);
nand U49286 (N_49286,N_48446,N_48599);
xnor U49287 (N_49287,N_48058,N_48487);
or U49288 (N_49288,N_48920,N_48981);
nor U49289 (N_49289,N_48646,N_48067);
xor U49290 (N_49290,N_48247,N_48181);
nor U49291 (N_49291,N_48894,N_48309);
nand U49292 (N_49292,N_48758,N_48909);
nand U49293 (N_49293,N_48858,N_48704);
and U49294 (N_49294,N_48068,N_48629);
xnor U49295 (N_49295,N_48850,N_48470);
or U49296 (N_49296,N_48063,N_48313);
and U49297 (N_49297,N_48326,N_48054);
nor U49298 (N_49298,N_48678,N_48507);
nor U49299 (N_49299,N_48092,N_48820);
nor U49300 (N_49300,N_48998,N_48623);
and U49301 (N_49301,N_48350,N_48390);
nand U49302 (N_49302,N_48363,N_48550);
and U49303 (N_49303,N_48733,N_48243);
nor U49304 (N_49304,N_48573,N_48696);
xor U49305 (N_49305,N_48985,N_48513);
or U49306 (N_49306,N_48808,N_48151);
nand U49307 (N_49307,N_48576,N_48845);
or U49308 (N_49308,N_48874,N_48490);
xnor U49309 (N_49309,N_48833,N_48632);
nand U49310 (N_49310,N_48699,N_48660);
xnor U49311 (N_49311,N_48506,N_48748);
or U49312 (N_49312,N_48239,N_48161);
or U49313 (N_49313,N_48362,N_48905);
nand U49314 (N_49314,N_48821,N_48311);
nand U49315 (N_49315,N_48582,N_48220);
nor U49316 (N_49316,N_48407,N_48711);
xor U49317 (N_49317,N_48011,N_48250);
nand U49318 (N_49318,N_48240,N_48472);
and U49319 (N_49319,N_48283,N_48871);
nor U49320 (N_49320,N_48382,N_48086);
nand U49321 (N_49321,N_48166,N_48155);
nand U49322 (N_49322,N_48625,N_48686);
nand U49323 (N_49323,N_48545,N_48028);
and U49324 (N_49324,N_48433,N_48951);
or U49325 (N_49325,N_48500,N_48404);
nand U49326 (N_49326,N_48520,N_48071);
xnor U49327 (N_49327,N_48112,N_48093);
or U49328 (N_49328,N_48073,N_48730);
xnor U49329 (N_49329,N_48752,N_48916);
and U49330 (N_49330,N_48290,N_48183);
or U49331 (N_49331,N_48903,N_48955);
or U49332 (N_49332,N_48791,N_48478);
xor U49333 (N_49333,N_48154,N_48120);
or U49334 (N_49334,N_48055,N_48318);
and U49335 (N_49335,N_48529,N_48383);
or U49336 (N_49336,N_48214,N_48235);
and U49337 (N_49337,N_48749,N_48327);
and U49338 (N_49338,N_48109,N_48343);
nand U49339 (N_49339,N_48098,N_48554);
nor U49340 (N_49340,N_48794,N_48128);
nor U49341 (N_49341,N_48111,N_48961);
xor U49342 (N_49342,N_48344,N_48289);
xnor U49343 (N_49343,N_48495,N_48022);
nand U49344 (N_49344,N_48338,N_48844);
or U49345 (N_49345,N_48182,N_48522);
and U49346 (N_49346,N_48296,N_48016);
nor U49347 (N_49347,N_48746,N_48705);
or U49348 (N_49348,N_48925,N_48102);
nor U49349 (N_49349,N_48261,N_48836);
nor U49350 (N_49350,N_48249,N_48974);
nand U49351 (N_49351,N_48041,N_48443);
nor U49352 (N_49352,N_48979,N_48211);
nor U49353 (N_49353,N_48650,N_48911);
nand U49354 (N_49354,N_48770,N_48800);
xor U49355 (N_49355,N_48441,N_48896);
or U49356 (N_49356,N_48551,N_48807);
and U49357 (N_49357,N_48883,N_48256);
nand U49358 (N_49358,N_48826,N_48865);
or U49359 (N_49359,N_48168,N_48100);
nor U49360 (N_49360,N_48608,N_48619);
nand U49361 (N_49361,N_48635,N_48025);
nand U49362 (N_49362,N_48185,N_48479);
and U49363 (N_49363,N_48303,N_48208);
nor U49364 (N_49364,N_48306,N_48014);
xnor U49365 (N_49365,N_48592,N_48340);
nor U49366 (N_49366,N_48143,N_48788);
or U49367 (N_49367,N_48387,N_48805);
or U49368 (N_49368,N_48885,N_48975);
or U49369 (N_49369,N_48688,N_48540);
and U49370 (N_49370,N_48265,N_48347);
nor U49371 (N_49371,N_48541,N_48684);
nand U49372 (N_49372,N_48204,N_48271);
and U49373 (N_49373,N_48237,N_48001);
and U49374 (N_49374,N_48033,N_48546);
or U49375 (N_49375,N_48499,N_48819);
xnor U49376 (N_49376,N_48921,N_48898);
xor U49377 (N_49377,N_48654,N_48771);
and U49378 (N_49378,N_48083,N_48357);
and U49379 (N_49379,N_48444,N_48355);
or U49380 (N_49380,N_48848,N_48897);
nand U49381 (N_49381,N_48255,N_48262);
xor U49382 (N_49382,N_48119,N_48687);
nor U49383 (N_49383,N_48037,N_48427);
nor U49384 (N_49384,N_48206,N_48910);
and U49385 (N_49385,N_48457,N_48426);
and U49386 (N_49386,N_48813,N_48868);
xor U49387 (N_49387,N_48454,N_48315);
and U49388 (N_49388,N_48192,N_48491);
nor U49389 (N_49389,N_48328,N_48873);
or U49390 (N_49390,N_48297,N_48837);
xnor U49391 (N_49391,N_48458,N_48999);
or U49392 (N_49392,N_48411,N_48860);
nor U49393 (N_49393,N_48275,N_48468);
nor U49394 (N_49394,N_48982,N_48069);
nand U49395 (N_49395,N_48976,N_48922);
nor U49396 (N_49396,N_48095,N_48003);
nor U49397 (N_49397,N_48051,N_48157);
xnor U49398 (N_49398,N_48649,N_48779);
nand U49399 (N_49399,N_48307,N_48203);
or U49400 (N_49400,N_48448,N_48633);
and U49401 (N_49401,N_48040,N_48706);
xor U49402 (N_49402,N_48153,N_48417);
nor U49403 (N_49403,N_48931,N_48581);
nand U49404 (N_49404,N_48144,N_48070);
xnor U49405 (N_49405,N_48721,N_48267);
nand U49406 (N_49406,N_48053,N_48377);
and U49407 (N_49407,N_48614,N_48869);
nand U49408 (N_49408,N_48079,N_48562);
and U49409 (N_49409,N_48538,N_48489);
nor U49410 (N_49410,N_48831,N_48317);
nor U49411 (N_49411,N_48123,N_48442);
nand U49412 (N_49412,N_48943,N_48009);
or U49413 (N_49413,N_48075,N_48533);
nor U49414 (N_49414,N_48689,N_48946);
xor U49415 (N_49415,N_48030,N_48544);
or U49416 (N_49416,N_48223,N_48575);
and U49417 (N_49417,N_48179,N_48172);
nor U49418 (N_49418,N_48277,N_48810);
nor U49419 (N_49419,N_48944,N_48725);
nor U49420 (N_49420,N_48132,N_48469);
nor U49421 (N_49421,N_48854,N_48209);
and U49422 (N_49422,N_48298,N_48336);
nand U49423 (N_49423,N_48859,N_48062);
nand U49424 (N_49424,N_48021,N_48205);
and U49425 (N_49425,N_48439,N_48829);
xor U49426 (N_49426,N_48878,N_48659);
nor U49427 (N_49427,N_48937,N_48270);
nor U49428 (N_49428,N_48316,N_48636);
nor U49429 (N_49429,N_48515,N_48967);
and U49430 (N_49430,N_48254,N_48782);
xnor U49431 (N_49431,N_48384,N_48164);
and U49432 (N_49432,N_48723,N_48139);
nor U49433 (N_49433,N_48739,N_48348);
nor U49434 (N_49434,N_48933,N_48484);
or U49435 (N_49435,N_48222,N_48783);
nand U49436 (N_49436,N_48558,N_48219);
and U49437 (N_49437,N_48605,N_48076);
or U49438 (N_49438,N_48882,N_48744);
nand U49439 (N_49439,N_48017,N_48867);
nand U49440 (N_49440,N_48504,N_48876);
xor U49441 (N_49441,N_48906,N_48189);
nand U49442 (N_49442,N_48645,N_48754);
or U49443 (N_49443,N_48305,N_48956);
nand U49444 (N_49444,N_48201,N_48294);
xor U49445 (N_49445,N_48847,N_48396);
nor U49446 (N_49446,N_48412,N_48360);
nor U49447 (N_49447,N_48708,N_48333);
nand U49448 (N_49448,N_48085,N_48657);
xnor U49449 (N_49449,N_48712,N_48757);
xnor U49450 (N_49450,N_48138,N_48938);
nand U49451 (N_49451,N_48827,N_48480);
xnor U49452 (N_49452,N_48787,N_48511);
xnor U49453 (N_49453,N_48552,N_48423);
nand U49454 (N_49454,N_48043,N_48110);
or U49455 (N_49455,N_48631,N_48107);
nor U49456 (N_49456,N_48584,N_48919);
or U49457 (N_49457,N_48475,N_48186);
nor U49458 (N_49458,N_48253,N_48815);
and U49459 (N_49459,N_48509,N_48090);
xnor U49460 (N_49460,N_48866,N_48492);
nor U49461 (N_49461,N_48774,N_48061);
nand U49462 (N_49462,N_48672,N_48620);
xor U49463 (N_49463,N_48236,N_48229);
nand U49464 (N_49464,N_48187,N_48923);
or U49465 (N_49465,N_48399,N_48548);
nand U49466 (N_49466,N_48414,N_48719);
or U49467 (N_49467,N_48986,N_48745);
nand U49468 (N_49468,N_48637,N_48613);
nand U49469 (N_49469,N_48212,N_48301);
or U49470 (N_49470,N_48852,N_48543);
or U49471 (N_49471,N_48715,N_48451);
nand U49472 (N_49472,N_48162,N_48685);
xnor U49473 (N_49473,N_48936,N_48924);
and U49474 (N_49474,N_48323,N_48408);
and U49475 (N_49475,N_48374,N_48435);
and U49476 (N_49476,N_48567,N_48050);
xnor U49477 (N_49477,N_48517,N_48512);
nand U49478 (N_49478,N_48004,N_48226);
and U49479 (N_49479,N_48940,N_48731);
xnor U49480 (N_49480,N_48600,N_48560);
xor U49481 (N_49481,N_48365,N_48453);
or U49482 (N_49482,N_48855,N_48949);
nor U49483 (N_49483,N_48308,N_48048);
xor U49484 (N_49484,N_48590,N_48539);
nand U49485 (N_49485,N_48234,N_48269);
xor U49486 (N_49486,N_48364,N_48588);
nor U49487 (N_49487,N_48035,N_48568);
xnor U49488 (N_49488,N_48525,N_48796);
nand U49489 (N_49489,N_48702,N_48881);
nand U49490 (N_49490,N_48996,N_48493);
or U49491 (N_49491,N_48345,N_48218);
and U49492 (N_49492,N_48150,N_48935);
and U49493 (N_49493,N_48952,N_48170);
nor U49494 (N_49494,N_48369,N_48785);
nor U49495 (N_49495,N_48742,N_48918);
nor U49496 (N_49496,N_48096,N_48401);
and U49497 (N_49497,N_48467,N_48354);
or U49498 (N_49498,N_48734,N_48171);
or U49499 (N_49499,N_48681,N_48091);
xnor U49500 (N_49500,N_48269,N_48350);
nand U49501 (N_49501,N_48311,N_48235);
nor U49502 (N_49502,N_48014,N_48743);
nor U49503 (N_49503,N_48238,N_48903);
nand U49504 (N_49504,N_48364,N_48908);
nand U49505 (N_49505,N_48973,N_48070);
xor U49506 (N_49506,N_48920,N_48658);
or U49507 (N_49507,N_48028,N_48504);
nor U49508 (N_49508,N_48087,N_48571);
nand U49509 (N_49509,N_48610,N_48606);
or U49510 (N_49510,N_48001,N_48876);
xnor U49511 (N_49511,N_48892,N_48772);
xnor U49512 (N_49512,N_48059,N_48787);
or U49513 (N_49513,N_48629,N_48171);
or U49514 (N_49514,N_48193,N_48473);
nor U49515 (N_49515,N_48462,N_48933);
xor U49516 (N_49516,N_48607,N_48466);
or U49517 (N_49517,N_48715,N_48520);
xor U49518 (N_49518,N_48094,N_48526);
nor U49519 (N_49519,N_48815,N_48595);
nand U49520 (N_49520,N_48051,N_48980);
or U49521 (N_49521,N_48729,N_48655);
xnor U49522 (N_49522,N_48812,N_48740);
nor U49523 (N_49523,N_48423,N_48600);
or U49524 (N_49524,N_48707,N_48368);
nor U49525 (N_49525,N_48823,N_48618);
or U49526 (N_49526,N_48553,N_48153);
xnor U49527 (N_49527,N_48057,N_48718);
xor U49528 (N_49528,N_48527,N_48066);
or U49529 (N_49529,N_48347,N_48149);
nor U49530 (N_49530,N_48271,N_48128);
nand U49531 (N_49531,N_48325,N_48844);
xnor U49532 (N_49532,N_48750,N_48216);
or U49533 (N_49533,N_48290,N_48314);
xnor U49534 (N_49534,N_48820,N_48775);
and U49535 (N_49535,N_48324,N_48439);
or U49536 (N_49536,N_48144,N_48523);
nor U49537 (N_49537,N_48109,N_48216);
xor U49538 (N_49538,N_48266,N_48988);
nor U49539 (N_49539,N_48540,N_48190);
and U49540 (N_49540,N_48885,N_48487);
or U49541 (N_49541,N_48502,N_48699);
xor U49542 (N_49542,N_48423,N_48037);
nand U49543 (N_49543,N_48104,N_48400);
or U49544 (N_49544,N_48884,N_48071);
nand U49545 (N_49545,N_48870,N_48529);
xnor U49546 (N_49546,N_48617,N_48542);
nand U49547 (N_49547,N_48987,N_48415);
or U49548 (N_49548,N_48536,N_48152);
xnor U49549 (N_49549,N_48663,N_48591);
and U49550 (N_49550,N_48414,N_48468);
xnor U49551 (N_49551,N_48749,N_48461);
xnor U49552 (N_49552,N_48576,N_48125);
nor U49553 (N_49553,N_48245,N_48248);
nor U49554 (N_49554,N_48491,N_48646);
xor U49555 (N_49555,N_48536,N_48764);
xor U49556 (N_49556,N_48754,N_48530);
or U49557 (N_49557,N_48402,N_48166);
xor U49558 (N_49558,N_48977,N_48506);
nand U49559 (N_49559,N_48312,N_48309);
or U49560 (N_49560,N_48554,N_48819);
and U49561 (N_49561,N_48348,N_48735);
and U49562 (N_49562,N_48738,N_48141);
xor U49563 (N_49563,N_48413,N_48792);
xor U49564 (N_49564,N_48932,N_48944);
xnor U49565 (N_49565,N_48585,N_48136);
nand U49566 (N_49566,N_48118,N_48561);
nand U49567 (N_49567,N_48242,N_48220);
nand U49568 (N_49568,N_48031,N_48709);
or U49569 (N_49569,N_48534,N_48195);
nand U49570 (N_49570,N_48567,N_48773);
nand U49571 (N_49571,N_48236,N_48472);
xnor U49572 (N_49572,N_48699,N_48896);
or U49573 (N_49573,N_48467,N_48837);
and U49574 (N_49574,N_48619,N_48660);
or U49575 (N_49575,N_48372,N_48767);
xor U49576 (N_49576,N_48295,N_48326);
nor U49577 (N_49577,N_48095,N_48790);
and U49578 (N_49578,N_48049,N_48200);
xnor U49579 (N_49579,N_48127,N_48050);
or U49580 (N_49580,N_48253,N_48178);
nor U49581 (N_49581,N_48151,N_48313);
or U49582 (N_49582,N_48259,N_48726);
or U49583 (N_49583,N_48960,N_48223);
or U49584 (N_49584,N_48671,N_48738);
nor U49585 (N_49585,N_48233,N_48882);
xnor U49586 (N_49586,N_48255,N_48887);
nor U49587 (N_49587,N_48445,N_48463);
and U49588 (N_49588,N_48865,N_48625);
nand U49589 (N_49589,N_48387,N_48710);
nor U49590 (N_49590,N_48073,N_48490);
xnor U49591 (N_49591,N_48047,N_48615);
nand U49592 (N_49592,N_48666,N_48138);
xnor U49593 (N_49593,N_48678,N_48073);
or U49594 (N_49594,N_48116,N_48757);
xor U49595 (N_49595,N_48716,N_48365);
xnor U49596 (N_49596,N_48642,N_48124);
nand U49597 (N_49597,N_48433,N_48151);
or U49598 (N_49598,N_48111,N_48519);
or U49599 (N_49599,N_48937,N_48339);
xor U49600 (N_49600,N_48875,N_48869);
nand U49601 (N_49601,N_48023,N_48026);
xor U49602 (N_49602,N_48815,N_48534);
and U49603 (N_49603,N_48383,N_48163);
or U49604 (N_49604,N_48154,N_48528);
nand U49605 (N_49605,N_48543,N_48122);
nor U49606 (N_49606,N_48174,N_48134);
or U49607 (N_49607,N_48397,N_48499);
nand U49608 (N_49608,N_48317,N_48105);
or U49609 (N_49609,N_48771,N_48898);
and U49610 (N_49610,N_48343,N_48119);
or U49611 (N_49611,N_48260,N_48920);
nor U49612 (N_49612,N_48012,N_48446);
nand U49613 (N_49613,N_48267,N_48490);
nand U49614 (N_49614,N_48201,N_48036);
and U49615 (N_49615,N_48413,N_48257);
nand U49616 (N_49616,N_48200,N_48306);
and U49617 (N_49617,N_48474,N_48563);
or U49618 (N_49618,N_48191,N_48620);
or U49619 (N_49619,N_48062,N_48396);
nand U49620 (N_49620,N_48184,N_48285);
or U49621 (N_49621,N_48747,N_48424);
and U49622 (N_49622,N_48197,N_48257);
nor U49623 (N_49623,N_48094,N_48292);
and U49624 (N_49624,N_48650,N_48224);
or U49625 (N_49625,N_48116,N_48598);
and U49626 (N_49626,N_48333,N_48194);
or U49627 (N_49627,N_48312,N_48489);
nor U49628 (N_49628,N_48258,N_48368);
and U49629 (N_49629,N_48640,N_48726);
nand U49630 (N_49630,N_48047,N_48667);
xnor U49631 (N_49631,N_48034,N_48748);
and U49632 (N_49632,N_48062,N_48808);
nand U49633 (N_49633,N_48016,N_48627);
or U49634 (N_49634,N_48033,N_48058);
xnor U49635 (N_49635,N_48161,N_48503);
xnor U49636 (N_49636,N_48154,N_48444);
nand U49637 (N_49637,N_48614,N_48332);
or U49638 (N_49638,N_48663,N_48777);
nor U49639 (N_49639,N_48392,N_48774);
or U49640 (N_49640,N_48789,N_48934);
and U49641 (N_49641,N_48347,N_48585);
xnor U49642 (N_49642,N_48537,N_48327);
nor U49643 (N_49643,N_48520,N_48539);
or U49644 (N_49644,N_48228,N_48802);
and U49645 (N_49645,N_48452,N_48593);
nor U49646 (N_49646,N_48972,N_48262);
and U49647 (N_49647,N_48762,N_48196);
or U49648 (N_49648,N_48959,N_48011);
and U49649 (N_49649,N_48806,N_48246);
xor U49650 (N_49650,N_48398,N_48102);
xor U49651 (N_49651,N_48254,N_48936);
nor U49652 (N_49652,N_48275,N_48312);
nand U49653 (N_49653,N_48488,N_48798);
xor U49654 (N_49654,N_48155,N_48950);
nor U49655 (N_49655,N_48270,N_48237);
and U49656 (N_49656,N_48426,N_48564);
nor U49657 (N_49657,N_48195,N_48357);
and U49658 (N_49658,N_48166,N_48465);
nand U49659 (N_49659,N_48527,N_48585);
nand U49660 (N_49660,N_48820,N_48349);
or U49661 (N_49661,N_48888,N_48393);
nand U49662 (N_49662,N_48983,N_48204);
or U49663 (N_49663,N_48499,N_48740);
nor U49664 (N_49664,N_48473,N_48569);
or U49665 (N_49665,N_48078,N_48787);
and U49666 (N_49666,N_48936,N_48528);
nor U49667 (N_49667,N_48991,N_48335);
and U49668 (N_49668,N_48853,N_48907);
nor U49669 (N_49669,N_48565,N_48483);
and U49670 (N_49670,N_48188,N_48110);
xnor U49671 (N_49671,N_48138,N_48637);
nand U49672 (N_49672,N_48980,N_48034);
and U49673 (N_49673,N_48361,N_48175);
or U49674 (N_49674,N_48918,N_48740);
and U49675 (N_49675,N_48547,N_48162);
nand U49676 (N_49676,N_48574,N_48360);
xor U49677 (N_49677,N_48697,N_48117);
nor U49678 (N_49678,N_48059,N_48652);
xnor U49679 (N_49679,N_48282,N_48291);
or U49680 (N_49680,N_48023,N_48733);
nor U49681 (N_49681,N_48756,N_48496);
or U49682 (N_49682,N_48262,N_48375);
nand U49683 (N_49683,N_48776,N_48654);
xor U49684 (N_49684,N_48251,N_48562);
and U49685 (N_49685,N_48897,N_48716);
and U49686 (N_49686,N_48668,N_48709);
xnor U49687 (N_49687,N_48772,N_48462);
nor U49688 (N_49688,N_48527,N_48187);
nand U49689 (N_49689,N_48495,N_48603);
xor U49690 (N_49690,N_48891,N_48501);
nor U49691 (N_49691,N_48706,N_48612);
or U49692 (N_49692,N_48525,N_48343);
xor U49693 (N_49693,N_48400,N_48607);
nand U49694 (N_49694,N_48829,N_48458);
and U49695 (N_49695,N_48305,N_48588);
and U49696 (N_49696,N_48915,N_48146);
or U49697 (N_49697,N_48989,N_48909);
and U49698 (N_49698,N_48493,N_48710);
nor U49699 (N_49699,N_48079,N_48295);
and U49700 (N_49700,N_48014,N_48777);
and U49701 (N_49701,N_48462,N_48466);
or U49702 (N_49702,N_48587,N_48690);
nand U49703 (N_49703,N_48471,N_48313);
nor U49704 (N_49704,N_48800,N_48992);
nor U49705 (N_49705,N_48142,N_48365);
xor U49706 (N_49706,N_48611,N_48150);
nand U49707 (N_49707,N_48402,N_48008);
and U49708 (N_49708,N_48310,N_48952);
xor U49709 (N_49709,N_48472,N_48097);
xnor U49710 (N_49710,N_48880,N_48013);
nor U49711 (N_49711,N_48437,N_48603);
and U49712 (N_49712,N_48632,N_48409);
nor U49713 (N_49713,N_48242,N_48520);
xnor U49714 (N_49714,N_48465,N_48595);
nand U49715 (N_49715,N_48129,N_48397);
nand U49716 (N_49716,N_48895,N_48117);
xnor U49717 (N_49717,N_48451,N_48655);
nor U49718 (N_49718,N_48267,N_48673);
or U49719 (N_49719,N_48096,N_48571);
or U49720 (N_49720,N_48801,N_48773);
xnor U49721 (N_49721,N_48640,N_48846);
or U49722 (N_49722,N_48208,N_48600);
xnor U49723 (N_49723,N_48823,N_48481);
or U49724 (N_49724,N_48425,N_48832);
nor U49725 (N_49725,N_48354,N_48419);
and U49726 (N_49726,N_48320,N_48313);
and U49727 (N_49727,N_48729,N_48124);
xnor U49728 (N_49728,N_48558,N_48346);
xnor U49729 (N_49729,N_48115,N_48733);
or U49730 (N_49730,N_48843,N_48242);
and U49731 (N_49731,N_48141,N_48495);
nor U49732 (N_49732,N_48300,N_48415);
nand U49733 (N_49733,N_48372,N_48313);
or U49734 (N_49734,N_48056,N_48662);
nand U49735 (N_49735,N_48125,N_48468);
nand U49736 (N_49736,N_48563,N_48398);
xor U49737 (N_49737,N_48131,N_48077);
or U49738 (N_49738,N_48499,N_48714);
nand U49739 (N_49739,N_48819,N_48532);
or U49740 (N_49740,N_48524,N_48405);
xnor U49741 (N_49741,N_48591,N_48890);
and U49742 (N_49742,N_48411,N_48454);
xor U49743 (N_49743,N_48454,N_48946);
nand U49744 (N_49744,N_48399,N_48217);
nand U49745 (N_49745,N_48588,N_48095);
and U49746 (N_49746,N_48585,N_48540);
and U49747 (N_49747,N_48851,N_48089);
nor U49748 (N_49748,N_48661,N_48832);
nor U49749 (N_49749,N_48937,N_48735);
and U49750 (N_49750,N_48035,N_48065);
and U49751 (N_49751,N_48322,N_48987);
xnor U49752 (N_49752,N_48985,N_48386);
nor U49753 (N_49753,N_48017,N_48670);
and U49754 (N_49754,N_48729,N_48714);
nor U49755 (N_49755,N_48766,N_48786);
xor U49756 (N_49756,N_48346,N_48527);
or U49757 (N_49757,N_48308,N_48060);
or U49758 (N_49758,N_48934,N_48087);
or U49759 (N_49759,N_48000,N_48150);
nand U49760 (N_49760,N_48029,N_48752);
or U49761 (N_49761,N_48985,N_48509);
or U49762 (N_49762,N_48586,N_48229);
nor U49763 (N_49763,N_48794,N_48381);
and U49764 (N_49764,N_48834,N_48769);
xor U49765 (N_49765,N_48264,N_48515);
or U49766 (N_49766,N_48308,N_48093);
and U49767 (N_49767,N_48677,N_48978);
xor U49768 (N_49768,N_48933,N_48675);
or U49769 (N_49769,N_48458,N_48844);
nor U49770 (N_49770,N_48813,N_48566);
nand U49771 (N_49771,N_48429,N_48176);
xnor U49772 (N_49772,N_48018,N_48774);
or U49773 (N_49773,N_48938,N_48153);
or U49774 (N_49774,N_48543,N_48051);
xnor U49775 (N_49775,N_48796,N_48337);
or U49776 (N_49776,N_48820,N_48362);
nand U49777 (N_49777,N_48764,N_48174);
or U49778 (N_49778,N_48034,N_48418);
nand U49779 (N_49779,N_48976,N_48831);
xor U49780 (N_49780,N_48767,N_48184);
nor U49781 (N_49781,N_48661,N_48422);
nand U49782 (N_49782,N_48486,N_48255);
nand U49783 (N_49783,N_48501,N_48907);
nor U49784 (N_49784,N_48964,N_48654);
or U49785 (N_49785,N_48859,N_48236);
nand U49786 (N_49786,N_48337,N_48052);
nand U49787 (N_49787,N_48502,N_48139);
and U49788 (N_49788,N_48696,N_48462);
or U49789 (N_49789,N_48374,N_48197);
nand U49790 (N_49790,N_48470,N_48612);
nor U49791 (N_49791,N_48064,N_48242);
nor U49792 (N_49792,N_48513,N_48474);
nor U49793 (N_49793,N_48862,N_48286);
nor U49794 (N_49794,N_48397,N_48005);
nor U49795 (N_49795,N_48141,N_48263);
and U49796 (N_49796,N_48117,N_48719);
nand U49797 (N_49797,N_48991,N_48397);
xnor U49798 (N_49798,N_48895,N_48542);
nor U49799 (N_49799,N_48982,N_48502);
and U49800 (N_49800,N_48835,N_48744);
and U49801 (N_49801,N_48978,N_48432);
or U49802 (N_49802,N_48507,N_48572);
nand U49803 (N_49803,N_48751,N_48694);
and U49804 (N_49804,N_48562,N_48739);
nand U49805 (N_49805,N_48414,N_48363);
and U49806 (N_49806,N_48586,N_48792);
or U49807 (N_49807,N_48779,N_48119);
or U49808 (N_49808,N_48716,N_48973);
nor U49809 (N_49809,N_48564,N_48868);
nor U49810 (N_49810,N_48706,N_48879);
nand U49811 (N_49811,N_48797,N_48832);
or U49812 (N_49812,N_48813,N_48784);
nand U49813 (N_49813,N_48005,N_48909);
nand U49814 (N_49814,N_48750,N_48647);
nor U49815 (N_49815,N_48854,N_48947);
and U49816 (N_49816,N_48884,N_48937);
nand U49817 (N_49817,N_48861,N_48924);
or U49818 (N_49818,N_48125,N_48087);
or U49819 (N_49819,N_48381,N_48249);
or U49820 (N_49820,N_48046,N_48992);
and U49821 (N_49821,N_48160,N_48086);
nor U49822 (N_49822,N_48104,N_48634);
nor U49823 (N_49823,N_48444,N_48842);
nor U49824 (N_49824,N_48646,N_48638);
nor U49825 (N_49825,N_48894,N_48529);
or U49826 (N_49826,N_48635,N_48140);
or U49827 (N_49827,N_48377,N_48230);
nand U49828 (N_49828,N_48787,N_48908);
nor U49829 (N_49829,N_48619,N_48130);
nand U49830 (N_49830,N_48399,N_48737);
and U49831 (N_49831,N_48558,N_48325);
and U49832 (N_49832,N_48929,N_48186);
nand U49833 (N_49833,N_48817,N_48404);
xor U49834 (N_49834,N_48345,N_48212);
nand U49835 (N_49835,N_48444,N_48122);
or U49836 (N_49836,N_48743,N_48620);
nand U49837 (N_49837,N_48436,N_48534);
xor U49838 (N_49838,N_48398,N_48735);
and U49839 (N_49839,N_48946,N_48187);
nand U49840 (N_49840,N_48850,N_48021);
and U49841 (N_49841,N_48503,N_48740);
nor U49842 (N_49842,N_48108,N_48269);
and U49843 (N_49843,N_48164,N_48021);
nor U49844 (N_49844,N_48972,N_48145);
nor U49845 (N_49845,N_48705,N_48875);
and U49846 (N_49846,N_48531,N_48847);
and U49847 (N_49847,N_48287,N_48094);
and U49848 (N_49848,N_48290,N_48341);
or U49849 (N_49849,N_48888,N_48915);
nor U49850 (N_49850,N_48134,N_48581);
nand U49851 (N_49851,N_48049,N_48920);
xnor U49852 (N_49852,N_48181,N_48751);
xor U49853 (N_49853,N_48034,N_48093);
xor U49854 (N_49854,N_48486,N_48864);
and U49855 (N_49855,N_48379,N_48865);
nor U49856 (N_49856,N_48650,N_48169);
nor U49857 (N_49857,N_48665,N_48498);
and U49858 (N_49858,N_48985,N_48829);
nor U49859 (N_49859,N_48451,N_48487);
nand U49860 (N_49860,N_48236,N_48215);
nand U49861 (N_49861,N_48046,N_48900);
nor U49862 (N_49862,N_48378,N_48942);
and U49863 (N_49863,N_48496,N_48978);
xor U49864 (N_49864,N_48180,N_48765);
or U49865 (N_49865,N_48757,N_48627);
nor U49866 (N_49866,N_48136,N_48357);
nand U49867 (N_49867,N_48876,N_48097);
and U49868 (N_49868,N_48394,N_48693);
nor U49869 (N_49869,N_48637,N_48925);
nand U49870 (N_49870,N_48393,N_48822);
nor U49871 (N_49871,N_48550,N_48476);
nand U49872 (N_49872,N_48108,N_48906);
nor U49873 (N_49873,N_48189,N_48735);
xor U49874 (N_49874,N_48850,N_48633);
and U49875 (N_49875,N_48134,N_48047);
nand U49876 (N_49876,N_48383,N_48791);
nor U49877 (N_49877,N_48555,N_48515);
and U49878 (N_49878,N_48462,N_48962);
and U49879 (N_49879,N_48664,N_48145);
or U49880 (N_49880,N_48624,N_48660);
xor U49881 (N_49881,N_48821,N_48153);
and U49882 (N_49882,N_48971,N_48921);
or U49883 (N_49883,N_48480,N_48781);
nor U49884 (N_49884,N_48654,N_48590);
nor U49885 (N_49885,N_48123,N_48184);
xnor U49886 (N_49886,N_48788,N_48021);
nand U49887 (N_49887,N_48403,N_48689);
nand U49888 (N_49888,N_48165,N_48629);
nor U49889 (N_49889,N_48335,N_48750);
or U49890 (N_49890,N_48200,N_48360);
nand U49891 (N_49891,N_48351,N_48793);
or U49892 (N_49892,N_48354,N_48671);
or U49893 (N_49893,N_48451,N_48772);
nand U49894 (N_49894,N_48276,N_48473);
xnor U49895 (N_49895,N_48729,N_48266);
nand U49896 (N_49896,N_48359,N_48791);
or U49897 (N_49897,N_48691,N_48927);
and U49898 (N_49898,N_48819,N_48980);
xnor U49899 (N_49899,N_48053,N_48130);
or U49900 (N_49900,N_48214,N_48252);
and U49901 (N_49901,N_48940,N_48387);
nor U49902 (N_49902,N_48351,N_48228);
xor U49903 (N_49903,N_48740,N_48771);
nor U49904 (N_49904,N_48445,N_48535);
or U49905 (N_49905,N_48965,N_48006);
nand U49906 (N_49906,N_48748,N_48989);
xor U49907 (N_49907,N_48753,N_48225);
xor U49908 (N_49908,N_48631,N_48083);
and U49909 (N_49909,N_48644,N_48117);
and U49910 (N_49910,N_48202,N_48738);
xor U49911 (N_49911,N_48405,N_48442);
xnor U49912 (N_49912,N_48792,N_48386);
xnor U49913 (N_49913,N_48636,N_48014);
nand U49914 (N_49914,N_48615,N_48136);
and U49915 (N_49915,N_48710,N_48758);
or U49916 (N_49916,N_48489,N_48154);
or U49917 (N_49917,N_48031,N_48624);
nand U49918 (N_49918,N_48842,N_48300);
and U49919 (N_49919,N_48144,N_48156);
nor U49920 (N_49920,N_48380,N_48351);
or U49921 (N_49921,N_48961,N_48783);
nand U49922 (N_49922,N_48180,N_48182);
nor U49923 (N_49923,N_48124,N_48593);
xor U49924 (N_49924,N_48799,N_48294);
and U49925 (N_49925,N_48418,N_48232);
or U49926 (N_49926,N_48851,N_48395);
or U49927 (N_49927,N_48840,N_48666);
nor U49928 (N_49928,N_48122,N_48892);
or U49929 (N_49929,N_48355,N_48897);
or U49930 (N_49930,N_48419,N_48047);
nand U49931 (N_49931,N_48036,N_48408);
nor U49932 (N_49932,N_48337,N_48151);
xnor U49933 (N_49933,N_48352,N_48109);
and U49934 (N_49934,N_48785,N_48547);
and U49935 (N_49935,N_48667,N_48456);
and U49936 (N_49936,N_48918,N_48555);
and U49937 (N_49937,N_48033,N_48541);
nor U49938 (N_49938,N_48778,N_48962);
nand U49939 (N_49939,N_48770,N_48634);
xor U49940 (N_49940,N_48734,N_48696);
nand U49941 (N_49941,N_48113,N_48279);
xnor U49942 (N_49942,N_48148,N_48018);
nand U49943 (N_49943,N_48715,N_48146);
nor U49944 (N_49944,N_48789,N_48924);
xnor U49945 (N_49945,N_48017,N_48328);
and U49946 (N_49946,N_48987,N_48852);
nor U49947 (N_49947,N_48622,N_48767);
and U49948 (N_49948,N_48978,N_48457);
nor U49949 (N_49949,N_48303,N_48999);
xor U49950 (N_49950,N_48362,N_48605);
or U49951 (N_49951,N_48969,N_48577);
nand U49952 (N_49952,N_48861,N_48502);
and U49953 (N_49953,N_48396,N_48115);
or U49954 (N_49954,N_48778,N_48170);
or U49955 (N_49955,N_48860,N_48391);
and U49956 (N_49956,N_48054,N_48851);
nor U49957 (N_49957,N_48414,N_48520);
or U49958 (N_49958,N_48833,N_48331);
and U49959 (N_49959,N_48248,N_48836);
and U49960 (N_49960,N_48545,N_48847);
nor U49961 (N_49961,N_48476,N_48109);
xnor U49962 (N_49962,N_48113,N_48440);
and U49963 (N_49963,N_48240,N_48356);
and U49964 (N_49964,N_48827,N_48646);
xor U49965 (N_49965,N_48697,N_48903);
or U49966 (N_49966,N_48852,N_48801);
nand U49967 (N_49967,N_48092,N_48025);
or U49968 (N_49968,N_48607,N_48450);
nor U49969 (N_49969,N_48544,N_48450);
xnor U49970 (N_49970,N_48494,N_48172);
nand U49971 (N_49971,N_48717,N_48298);
or U49972 (N_49972,N_48100,N_48449);
xnor U49973 (N_49973,N_48652,N_48431);
nor U49974 (N_49974,N_48086,N_48291);
or U49975 (N_49975,N_48607,N_48494);
nand U49976 (N_49976,N_48034,N_48215);
nor U49977 (N_49977,N_48198,N_48962);
or U49978 (N_49978,N_48961,N_48437);
nand U49979 (N_49979,N_48954,N_48107);
and U49980 (N_49980,N_48828,N_48317);
xor U49981 (N_49981,N_48350,N_48367);
and U49982 (N_49982,N_48031,N_48748);
nor U49983 (N_49983,N_48736,N_48697);
xnor U49984 (N_49984,N_48224,N_48154);
xnor U49985 (N_49985,N_48168,N_48781);
xor U49986 (N_49986,N_48454,N_48027);
nand U49987 (N_49987,N_48256,N_48127);
and U49988 (N_49988,N_48259,N_48418);
and U49989 (N_49989,N_48068,N_48178);
nor U49990 (N_49990,N_48506,N_48807);
nand U49991 (N_49991,N_48729,N_48304);
and U49992 (N_49992,N_48785,N_48259);
nand U49993 (N_49993,N_48543,N_48367);
nand U49994 (N_49994,N_48757,N_48121);
nor U49995 (N_49995,N_48709,N_48593);
nand U49996 (N_49996,N_48861,N_48434);
xor U49997 (N_49997,N_48411,N_48251);
nor U49998 (N_49998,N_48349,N_48754);
nor U49999 (N_49999,N_48243,N_48735);
or UO_0 (O_0,N_49810,N_49160);
nor UO_1 (O_1,N_49667,N_49754);
nand UO_2 (O_2,N_49429,N_49078);
and UO_3 (O_3,N_49280,N_49194);
nor UO_4 (O_4,N_49283,N_49446);
xor UO_5 (O_5,N_49290,N_49248);
and UO_6 (O_6,N_49615,N_49686);
and UO_7 (O_7,N_49588,N_49554);
nand UO_8 (O_8,N_49816,N_49985);
nor UO_9 (O_9,N_49865,N_49025);
and UO_10 (O_10,N_49513,N_49591);
nor UO_11 (O_11,N_49433,N_49483);
and UO_12 (O_12,N_49219,N_49037);
xnor UO_13 (O_13,N_49300,N_49647);
nand UO_14 (O_14,N_49868,N_49352);
xnor UO_15 (O_15,N_49547,N_49031);
or UO_16 (O_16,N_49200,N_49074);
nor UO_17 (O_17,N_49691,N_49537);
xor UO_18 (O_18,N_49976,N_49975);
nand UO_19 (O_19,N_49286,N_49343);
nand UO_20 (O_20,N_49385,N_49707);
xnor UO_21 (O_21,N_49578,N_49313);
nand UO_22 (O_22,N_49546,N_49413);
nand UO_23 (O_23,N_49706,N_49632);
nand UO_24 (O_24,N_49684,N_49141);
and UO_25 (O_25,N_49581,N_49837);
and UO_26 (O_26,N_49409,N_49961);
nor UO_27 (O_27,N_49799,N_49240);
nor UO_28 (O_28,N_49963,N_49403);
nand UO_29 (O_29,N_49759,N_49855);
nand UO_30 (O_30,N_49238,N_49811);
xor UO_31 (O_31,N_49079,N_49293);
or UO_32 (O_32,N_49188,N_49830);
and UO_33 (O_33,N_49815,N_49666);
nor UO_34 (O_34,N_49886,N_49577);
and UO_35 (O_35,N_49199,N_49717);
and UO_36 (O_36,N_49368,N_49172);
nor UO_37 (O_37,N_49258,N_49121);
and UO_38 (O_38,N_49384,N_49391);
nand UO_39 (O_39,N_49056,N_49072);
and UO_40 (O_40,N_49872,N_49016);
nor UO_41 (O_41,N_49856,N_49840);
or UO_42 (O_42,N_49273,N_49355);
xnor UO_43 (O_43,N_49967,N_49347);
xnor UO_44 (O_44,N_49968,N_49875);
nor UO_45 (O_45,N_49338,N_49242);
nor UO_46 (O_46,N_49812,N_49898);
nand UO_47 (O_47,N_49998,N_49923);
nand UO_48 (O_48,N_49097,N_49251);
or UO_49 (O_49,N_49645,N_49274);
xnor UO_50 (O_50,N_49824,N_49900);
and UO_51 (O_51,N_49491,N_49128);
xnor UO_52 (O_52,N_49676,N_49992);
nor UO_53 (O_53,N_49096,N_49540);
xnor UO_54 (O_54,N_49979,N_49575);
nand UO_55 (O_55,N_49741,N_49517);
or UO_56 (O_56,N_49146,N_49880);
nand UO_57 (O_57,N_49606,N_49438);
nand UO_58 (O_58,N_49610,N_49425);
and UO_59 (O_59,N_49109,N_49298);
nor UO_60 (O_60,N_49076,N_49589);
or UO_61 (O_61,N_49253,N_49068);
nor UO_62 (O_62,N_49538,N_49829);
and UO_63 (O_63,N_49607,N_49753);
or UO_64 (O_64,N_49584,N_49044);
or UO_65 (O_65,N_49966,N_49239);
xnor UO_66 (O_66,N_49738,N_49652);
xor UO_67 (O_67,N_49921,N_49677);
or UO_68 (O_68,N_49322,N_49646);
nand UO_69 (O_69,N_49545,N_49291);
xor UO_70 (O_70,N_49061,N_49552);
nor UO_71 (O_71,N_49447,N_49709);
or UO_72 (O_72,N_49245,N_49374);
and UO_73 (O_73,N_49122,N_49278);
nor UO_74 (O_74,N_49225,N_49972);
xor UO_75 (O_75,N_49850,N_49416);
or UO_76 (O_76,N_49271,N_49507);
nor UO_77 (O_77,N_49262,N_49136);
and UO_78 (O_78,N_49372,N_49482);
or UO_79 (O_79,N_49550,N_49426);
nand UO_80 (O_80,N_49959,N_49530);
xor UO_81 (O_81,N_49612,N_49264);
nand UO_82 (O_82,N_49474,N_49272);
nand UO_83 (O_83,N_49557,N_49441);
and UO_84 (O_84,N_49783,N_49820);
nand UO_85 (O_85,N_49876,N_49023);
nor UO_86 (O_86,N_49523,N_49869);
nor UO_87 (O_87,N_49281,N_49462);
or UO_88 (O_88,N_49574,N_49616);
xor UO_89 (O_89,N_49542,N_49247);
nand UO_90 (O_90,N_49326,N_49341);
xor UO_91 (O_91,N_49693,N_49442);
or UO_92 (O_92,N_49661,N_49116);
nor UO_93 (O_93,N_49604,N_49756);
or UO_94 (O_94,N_49674,N_49903);
xor UO_95 (O_95,N_49479,N_49157);
nand UO_96 (O_96,N_49080,N_49318);
or UO_97 (O_97,N_49214,N_49135);
nand UO_98 (O_98,N_49496,N_49252);
or UO_99 (O_99,N_49763,N_49493);
nor UO_100 (O_100,N_49534,N_49489);
or UO_101 (O_101,N_49611,N_49703);
nand UO_102 (O_102,N_49958,N_49301);
or UO_103 (O_103,N_49087,N_49508);
or UO_104 (O_104,N_49001,N_49977);
xnor UO_105 (O_105,N_49360,N_49719);
nor UO_106 (O_106,N_49656,N_49487);
nand UO_107 (O_107,N_49231,N_49805);
nand UO_108 (O_108,N_49051,N_49039);
or UO_109 (O_109,N_49622,N_49062);
xor UO_110 (O_110,N_49004,N_49728);
nor UO_111 (O_111,N_49393,N_49465);
xor UO_112 (O_112,N_49701,N_49910);
or UO_113 (O_113,N_49295,N_49407);
nor UO_114 (O_114,N_49367,N_49924);
nor UO_115 (O_115,N_49395,N_49739);
and UO_116 (O_116,N_49640,N_49359);
xnor UO_117 (O_117,N_49038,N_49218);
and UO_118 (O_118,N_49234,N_49593);
xnor UO_119 (O_119,N_49100,N_49908);
and UO_120 (O_120,N_49854,N_49406);
nor UO_121 (O_121,N_49134,N_49637);
and UO_122 (O_122,N_49635,N_49381);
or UO_123 (O_123,N_49941,N_49323);
nand UO_124 (O_124,N_49651,N_49777);
and UO_125 (O_125,N_49965,N_49269);
xnor UO_126 (O_126,N_49205,N_49166);
xor UO_127 (O_127,N_49949,N_49867);
nor UO_128 (O_128,N_49931,N_49729);
nor UO_129 (O_129,N_49369,N_49005);
or UO_130 (O_130,N_49821,N_49354);
or UO_131 (O_131,N_49551,N_49505);
xor UO_132 (O_132,N_49871,N_49432);
or UO_133 (O_133,N_49766,N_49436);
and UO_134 (O_134,N_49158,N_49527);
xor UO_135 (O_135,N_49337,N_49119);
nand UO_136 (O_136,N_49771,N_49504);
nand UO_137 (O_137,N_49881,N_49373);
and UO_138 (O_138,N_49555,N_49917);
nand UO_139 (O_139,N_49843,N_49093);
and UO_140 (O_140,N_49882,N_49046);
and UO_141 (O_141,N_49648,N_49309);
xor UO_142 (O_142,N_49042,N_49101);
nand UO_143 (O_143,N_49411,N_49311);
or UO_144 (O_144,N_49579,N_49452);
nor UO_145 (O_145,N_49649,N_49712);
nand UO_146 (O_146,N_49492,N_49605);
nand UO_147 (O_147,N_49644,N_49981);
nor UO_148 (O_148,N_49720,N_49013);
and UO_149 (O_149,N_49866,N_49642);
and UO_150 (O_150,N_49069,N_49573);
nand UO_151 (O_151,N_49502,N_49559);
xor UO_152 (O_152,N_49246,N_49950);
nor UO_153 (O_153,N_49680,N_49027);
and UO_154 (O_154,N_49340,N_49156);
nor UO_155 (O_155,N_49665,N_49112);
xnor UO_156 (O_156,N_49955,N_49249);
nand UO_157 (O_157,N_49159,N_49212);
xor UO_158 (O_158,N_49501,N_49528);
nand UO_159 (O_159,N_49702,N_49202);
nand UO_160 (O_160,N_49105,N_49726);
xor UO_161 (O_161,N_49472,N_49983);
and UO_162 (O_162,N_49437,N_49599);
nand UO_163 (O_163,N_49724,N_49427);
and UO_164 (O_164,N_49678,N_49774);
nand UO_165 (O_165,N_49388,N_49223);
nand UO_166 (O_166,N_49449,N_49028);
or UO_167 (O_167,N_49948,N_49475);
or UO_168 (O_168,N_49690,N_49842);
or UO_169 (O_169,N_49417,N_49077);
nor UO_170 (O_170,N_49365,N_49107);
and UO_171 (O_171,N_49458,N_49618);
nor UO_172 (O_172,N_49879,N_49292);
xor UO_173 (O_173,N_49276,N_49902);
nor UO_174 (O_174,N_49735,N_49544);
or UO_175 (O_175,N_49059,N_49627);
xnor UO_176 (O_176,N_49435,N_49997);
and UO_177 (O_177,N_49410,N_49319);
or UO_178 (O_178,N_49220,N_49541);
nand UO_179 (O_179,N_49344,N_49423);
nand UO_180 (O_180,N_49021,N_49746);
xor UO_181 (O_181,N_49711,N_49945);
nand UO_182 (O_182,N_49813,N_49114);
xor UO_183 (O_183,N_49184,N_49800);
nand UO_184 (O_184,N_49768,N_49994);
nor UO_185 (O_185,N_49636,N_49339);
or UO_186 (O_186,N_49934,N_49520);
xnor UO_187 (O_187,N_49486,N_49329);
xor UO_188 (O_188,N_49216,N_49152);
nor UO_189 (O_189,N_49382,N_49862);
or UO_190 (O_190,N_49174,N_49564);
and UO_191 (O_191,N_49583,N_49792);
xor UO_192 (O_192,N_49823,N_49990);
nand UO_193 (O_193,N_49526,N_49034);
or UO_194 (O_194,N_49130,N_49495);
xnor UO_195 (O_195,N_49461,N_49560);
nand UO_196 (O_196,N_49129,N_49757);
xnor UO_197 (O_197,N_49389,N_49094);
xnor UO_198 (O_198,N_49919,N_49162);
xor UO_199 (O_199,N_49991,N_49722);
nor UO_200 (O_200,N_49418,N_49650);
nand UO_201 (O_201,N_49818,N_49918);
xor UO_202 (O_202,N_49566,N_49464);
nor UO_203 (O_203,N_49896,N_49822);
and UO_204 (O_204,N_49628,N_49890);
xor UO_205 (O_205,N_49089,N_49851);
nor UO_206 (O_206,N_49834,N_49082);
nor UO_207 (O_207,N_49529,N_49222);
or UO_208 (O_208,N_49254,N_49209);
nor UO_209 (O_209,N_49603,N_49192);
nor UO_210 (O_210,N_49884,N_49548);
or UO_211 (O_211,N_49699,N_49933);
nand UO_212 (O_212,N_49509,N_49095);
xor UO_213 (O_213,N_49852,N_49971);
nand UO_214 (O_214,N_49030,N_49161);
and UO_215 (O_215,N_49196,N_49050);
nand UO_216 (O_216,N_49450,N_49781);
xnor UO_217 (O_217,N_49600,N_49704);
nand UO_218 (O_218,N_49000,N_49210);
or UO_219 (O_219,N_49443,N_49939);
nor UO_220 (O_220,N_49909,N_49839);
xnor UO_221 (O_221,N_49477,N_49999);
and UO_222 (O_222,N_49685,N_49904);
and UO_223 (O_223,N_49658,N_49831);
and UO_224 (O_224,N_49110,N_49170);
and UO_225 (O_225,N_49598,N_49629);
or UO_226 (O_226,N_49467,N_49791);
or UO_227 (O_227,N_49190,N_49569);
xor UO_228 (O_228,N_49106,N_49532);
or UO_229 (O_229,N_49412,N_49498);
nor UO_230 (O_230,N_49476,N_49421);
or UO_231 (O_231,N_49480,N_49673);
nand UO_232 (O_232,N_49115,N_49187);
nand UO_233 (O_233,N_49775,N_49186);
nand UO_234 (O_234,N_49207,N_49178);
nand UO_235 (O_235,N_49349,N_49585);
or UO_236 (O_236,N_49989,N_49285);
xor UO_237 (O_237,N_49376,N_49597);
nand UO_238 (O_238,N_49624,N_49960);
xor UO_239 (O_239,N_49883,N_49377);
nand UO_240 (O_240,N_49232,N_49053);
nor UO_241 (O_241,N_49683,N_49054);
nand UO_242 (O_242,N_49996,N_49609);
nor UO_243 (O_243,N_49478,N_49952);
or UO_244 (O_244,N_49448,N_49362);
and UO_245 (O_245,N_49916,N_49206);
and UO_246 (O_246,N_49663,N_49075);
xnor UO_247 (O_247,N_49328,N_49317);
and UO_248 (O_248,N_49802,N_49613);
or UO_249 (O_249,N_49179,N_49858);
nor UO_250 (O_250,N_49090,N_49085);
or UO_251 (O_251,N_49133,N_49695);
or UO_252 (O_252,N_49149,N_49586);
and UO_253 (O_253,N_49197,N_49655);
or UO_254 (O_254,N_49743,N_49727);
xnor UO_255 (O_255,N_49137,N_49055);
or UO_256 (O_256,N_49964,N_49060);
xor UO_257 (O_257,N_49092,N_49497);
xor UO_258 (O_258,N_49164,N_49342);
nand UO_259 (O_259,N_49838,N_49926);
nor UO_260 (O_260,N_49229,N_49751);
and UO_261 (O_261,N_49671,N_49500);
or UO_262 (O_262,N_49696,N_49103);
xor UO_263 (O_263,N_49870,N_49601);
nand UO_264 (O_264,N_49543,N_49081);
or UO_265 (O_265,N_49859,N_49316);
nand UO_266 (O_266,N_49940,N_49399);
nor UO_267 (O_267,N_49324,N_49424);
xor UO_268 (O_268,N_49143,N_49330);
or UO_269 (O_269,N_49083,N_49067);
nor UO_270 (O_270,N_49463,N_49947);
or UO_271 (O_271,N_49063,N_49386);
or UO_272 (O_272,N_49198,N_49742);
or UO_273 (O_273,N_49394,N_49911);
nand UO_274 (O_274,N_49848,N_49953);
and UO_275 (O_275,N_49014,N_49236);
xor UO_276 (O_276,N_49710,N_49969);
nor UO_277 (O_277,N_49088,N_49980);
xor UO_278 (O_278,N_49086,N_49894);
or UO_279 (O_279,N_49936,N_49571);
xor UO_280 (O_280,N_49163,N_49761);
xor UO_281 (O_281,N_49444,N_49721);
and UO_282 (O_282,N_49503,N_49333);
or UO_283 (O_283,N_49414,N_49750);
nor UO_284 (O_284,N_49937,N_49327);
or UO_285 (O_285,N_49193,N_49131);
or UO_286 (O_286,N_49221,N_49572);
nor UO_287 (O_287,N_49380,N_49925);
nand UO_288 (O_288,N_49378,N_49630);
and UO_289 (O_289,N_49139,N_49984);
xor UO_290 (O_290,N_49621,N_49836);
xnor UO_291 (O_291,N_49625,N_49951);
and UO_292 (O_292,N_49405,N_49468);
nand UO_293 (O_293,N_49796,N_49906);
or UO_294 (O_294,N_49734,N_49008);
and UO_295 (O_295,N_49058,N_49889);
xor UO_296 (O_296,N_49689,N_49263);
nand UO_297 (O_297,N_49522,N_49594);
and UO_298 (O_298,N_49383,N_49457);
and UO_299 (O_299,N_49634,N_49453);
or UO_300 (O_300,N_49809,N_49512);
or UO_301 (O_301,N_49244,N_49404);
or UO_302 (O_302,N_49731,N_49325);
xor UO_303 (O_303,N_49203,N_49670);
and UO_304 (O_304,N_49901,N_49032);
nand UO_305 (O_305,N_49180,N_49120);
xnor UO_306 (O_306,N_49827,N_49456);
nor UO_307 (O_307,N_49790,N_49626);
nand UO_308 (O_308,N_49877,N_49752);
nor UO_309 (O_309,N_49714,N_49392);
nand UO_310 (O_310,N_49803,N_49697);
nor UO_311 (O_311,N_49125,N_49215);
nand UO_312 (O_312,N_49778,N_49978);
nor UO_313 (O_313,N_49204,N_49779);
nor UO_314 (O_314,N_49304,N_49619);
and UO_315 (O_315,N_49036,N_49428);
nor UO_316 (O_316,N_49108,N_49314);
and UO_317 (O_317,N_49142,N_49835);
xor UO_318 (O_318,N_49794,N_49460);
and UO_319 (O_319,N_49905,N_49357);
and UO_320 (O_320,N_49104,N_49124);
and UO_321 (O_321,N_49145,N_49113);
or UO_322 (O_322,N_49929,N_49439);
or UO_323 (O_323,N_49208,N_49748);
xor UO_324 (O_324,N_49725,N_49688);
xnor UO_325 (O_325,N_49175,N_49844);
and UO_326 (O_326,N_49847,N_49167);
nor UO_327 (O_327,N_49846,N_49303);
and UO_328 (O_328,N_49375,N_49587);
nand UO_329 (O_329,N_49144,N_49970);
and UO_330 (O_330,N_49899,N_49070);
xor UO_331 (O_331,N_49713,N_49806);
nor UO_332 (O_332,N_49195,N_49845);
and UO_333 (O_333,N_49266,N_49776);
or UO_334 (O_334,N_49469,N_49988);
xor UO_335 (O_335,N_49828,N_49857);
nor UO_336 (O_336,N_49277,N_49066);
xor UO_337 (O_337,N_49024,N_49211);
nor UO_338 (O_338,N_49260,N_49825);
or UO_339 (O_339,N_49226,N_49256);
nand UO_340 (O_340,N_49641,N_49073);
and UO_341 (O_341,N_49138,N_49568);
nand UO_342 (O_342,N_49602,N_49762);
xor UO_343 (O_343,N_49895,N_49864);
or UO_344 (O_344,N_49228,N_49631);
nor UO_345 (O_345,N_49071,N_49654);
nand UO_346 (O_346,N_49020,N_49912);
or UO_347 (O_347,N_49241,N_49506);
nor UO_348 (O_348,N_49396,N_49250);
nor UO_349 (O_349,N_49336,N_49307);
and UO_350 (O_350,N_49804,N_49785);
and UO_351 (O_351,N_49230,N_49282);
xor UO_352 (O_352,N_49920,N_49484);
or UO_353 (O_353,N_49420,N_49817);
nand UO_354 (O_354,N_49312,N_49265);
xor UO_355 (O_355,N_49043,N_49401);
or UO_356 (O_356,N_49029,N_49191);
or UO_357 (O_357,N_49118,N_49596);
xor UO_358 (O_358,N_49536,N_49350);
xor UO_359 (O_359,N_49363,N_49732);
nand UO_360 (O_360,N_49946,N_49764);
and UO_361 (O_361,N_49470,N_49102);
xnor UO_362 (O_362,N_49539,N_49772);
or UO_363 (O_363,N_49140,N_49927);
xor UO_364 (O_364,N_49694,N_49454);
nor UO_365 (O_365,N_49049,N_49795);
nand UO_366 (O_366,N_49730,N_49797);
nand UO_367 (O_367,N_49255,N_49715);
nand UO_368 (O_368,N_49954,N_49891);
nand UO_369 (O_369,N_49227,N_49408);
xnor UO_370 (O_370,N_49798,N_49814);
xor UO_371 (O_371,N_49773,N_49887);
xor UO_372 (O_372,N_49897,N_49692);
or UO_373 (O_373,N_49576,N_49047);
xor UO_374 (O_374,N_49788,N_49657);
xnor UO_375 (O_375,N_49767,N_49893);
and UO_376 (O_376,N_49494,N_49957);
xor UO_377 (O_377,N_49320,N_49789);
xor UO_378 (O_378,N_49525,N_49863);
nand UO_379 (O_379,N_49315,N_49306);
nand UO_380 (O_380,N_49348,N_49786);
nor UO_381 (O_381,N_49201,N_49679);
or UO_382 (O_382,N_49123,N_49758);
and UO_383 (O_383,N_49169,N_49760);
nand UO_384 (O_384,N_49052,N_49928);
nor UO_385 (O_385,N_49155,N_49451);
or UO_386 (O_386,N_49669,N_49364);
xnor UO_387 (O_387,N_49833,N_49787);
and UO_388 (O_388,N_49716,N_49708);
xnor UO_389 (O_389,N_49668,N_49807);
nand UO_390 (O_390,N_49973,N_49769);
and UO_391 (O_391,N_49065,N_49639);
or UO_392 (O_392,N_49400,N_49723);
and UO_393 (O_393,N_49740,N_49361);
nand UO_394 (O_394,N_49565,N_49993);
xnor UO_395 (O_395,N_49173,N_49653);
xnor UO_396 (O_396,N_49562,N_49595);
and UO_397 (O_397,N_49099,N_49022);
and UO_398 (O_398,N_49390,N_49516);
or UO_399 (O_399,N_49308,N_49006);
nor UO_400 (O_400,N_49705,N_49358);
or UO_401 (O_401,N_49018,N_49398);
and UO_402 (O_402,N_49268,N_49370);
nand UO_403 (O_403,N_49091,N_49681);
and UO_404 (O_404,N_49826,N_49459);
and UO_405 (O_405,N_49275,N_49419);
nand UO_406 (O_406,N_49356,N_49853);
or UO_407 (O_407,N_49302,N_49235);
or UO_408 (O_408,N_49287,N_49415);
and UO_409 (O_409,N_49007,N_49183);
nand UO_410 (O_410,N_49182,N_49284);
or UO_411 (O_411,N_49907,N_49176);
nand UO_412 (O_412,N_49533,N_49177);
and UO_413 (O_413,N_49440,N_49379);
xor UO_414 (O_414,N_49745,N_49288);
xnor UO_415 (O_415,N_49638,N_49995);
or UO_416 (O_416,N_49561,N_49366);
and UO_417 (O_417,N_49553,N_49535);
nand UO_418 (O_418,N_49267,N_49549);
nand UO_419 (O_419,N_49832,N_49132);
or UO_420 (O_420,N_49942,N_49003);
nor UO_421 (O_421,N_49747,N_49922);
nor UO_422 (O_422,N_49213,N_49387);
nand UO_423 (O_423,N_49422,N_49026);
nor UO_424 (O_424,N_49165,N_49986);
nand UO_425 (O_425,N_49321,N_49310);
and UO_426 (O_426,N_49057,N_49662);
nor UO_427 (O_427,N_49033,N_49473);
and UO_428 (O_428,N_49168,N_49860);
nand UO_429 (O_429,N_49181,N_49643);
nor UO_430 (O_430,N_49299,N_49956);
nand UO_431 (O_431,N_49892,N_49017);
nand UO_432 (O_432,N_49488,N_49010);
nor UO_433 (O_433,N_49117,N_49471);
or UO_434 (O_434,N_49913,N_49185);
and UO_435 (O_435,N_49617,N_49620);
nor UO_436 (O_436,N_49808,N_49098);
nand UO_437 (O_437,N_49127,N_49296);
nor UO_438 (O_438,N_49153,N_49445);
nand UO_439 (O_439,N_49888,N_49567);
xnor UO_440 (O_440,N_49664,N_49455);
and UO_441 (O_441,N_49755,N_49431);
nand UO_442 (O_442,N_49434,N_49885);
and UO_443 (O_443,N_49718,N_49733);
nor UO_444 (O_444,N_49521,N_49749);
and UO_445 (O_445,N_49849,N_49861);
or UO_446 (O_446,N_49556,N_49930);
nor UO_447 (O_447,N_49590,N_49744);
and UO_448 (O_448,N_49736,N_49700);
and UO_449 (O_449,N_49563,N_49259);
xor UO_450 (O_450,N_49040,N_49233);
or UO_451 (O_451,N_49841,N_49289);
nor UO_452 (O_452,N_49801,N_49614);
xnor UO_453 (O_453,N_49943,N_49334);
or UO_454 (O_454,N_49932,N_49148);
or UO_455 (O_455,N_49938,N_49793);
or UO_456 (O_456,N_49064,N_49397);
xnor UO_457 (O_457,N_49481,N_49765);
and UO_458 (O_458,N_49675,N_49009);
nor UO_459 (O_459,N_49257,N_49698);
or UO_460 (O_460,N_49171,N_49878);
nand UO_461 (O_461,N_49623,N_49819);
nor UO_462 (O_462,N_49045,N_49608);
or UO_463 (O_463,N_49002,N_49154);
or UO_464 (O_464,N_49935,N_49019);
and UO_465 (O_465,N_49294,N_49770);
xor UO_466 (O_466,N_49974,N_49873);
and UO_467 (O_467,N_49279,N_49633);
nor UO_468 (O_468,N_49237,N_49150);
and UO_469 (O_469,N_49660,N_49570);
and UO_470 (O_470,N_49147,N_49297);
and UO_471 (O_471,N_49331,N_49687);
nor UO_472 (O_472,N_49243,N_49682);
and UO_473 (O_473,N_49151,N_49982);
xor UO_474 (O_474,N_49041,N_49987);
nor UO_475 (O_475,N_49780,N_49874);
xnor UO_476 (O_476,N_49531,N_49012);
nand UO_477 (O_477,N_49672,N_49224);
or UO_478 (O_478,N_49962,N_49335);
xor UO_479 (O_479,N_49011,N_49084);
and UO_480 (O_480,N_49582,N_49485);
xor UO_481 (O_481,N_49189,N_49332);
nor UO_482 (O_482,N_49035,N_49048);
xnor UO_483 (O_483,N_49261,N_49270);
nand UO_484 (O_484,N_49346,N_49514);
and UO_485 (O_485,N_49737,N_49305);
xnor UO_486 (O_486,N_49914,N_49944);
or UO_487 (O_487,N_49402,N_49430);
nor UO_488 (O_488,N_49782,N_49490);
nand UO_489 (O_489,N_49353,N_49580);
or UO_490 (O_490,N_49345,N_49466);
xnor UO_491 (O_491,N_49518,N_49510);
nand UO_492 (O_492,N_49126,N_49524);
and UO_493 (O_493,N_49592,N_49015);
and UO_494 (O_494,N_49351,N_49558);
and UO_495 (O_495,N_49511,N_49111);
or UO_496 (O_496,N_49519,N_49784);
and UO_497 (O_497,N_49217,N_49499);
or UO_498 (O_498,N_49659,N_49371);
xor UO_499 (O_499,N_49915,N_49515);
nor UO_500 (O_500,N_49457,N_49407);
nor UO_501 (O_501,N_49994,N_49962);
and UO_502 (O_502,N_49183,N_49152);
nand UO_503 (O_503,N_49579,N_49234);
and UO_504 (O_504,N_49250,N_49324);
or UO_505 (O_505,N_49208,N_49953);
or UO_506 (O_506,N_49554,N_49147);
and UO_507 (O_507,N_49187,N_49164);
and UO_508 (O_508,N_49959,N_49687);
nand UO_509 (O_509,N_49976,N_49058);
xor UO_510 (O_510,N_49507,N_49677);
nor UO_511 (O_511,N_49376,N_49711);
nand UO_512 (O_512,N_49482,N_49031);
nand UO_513 (O_513,N_49158,N_49509);
and UO_514 (O_514,N_49581,N_49805);
nor UO_515 (O_515,N_49474,N_49074);
nor UO_516 (O_516,N_49961,N_49885);
and UO_517 (O_517,N_49101,N_49177);
nand UO_518 (O_518,N_49846,N_49202);
and UO_519 (O_519,N_49989,N_49316);
or UO_520 (O_520,N_49320,N_49728);
and UO_521 (O_521,N_49803,N_49655);
nand UO_522 (O_522,N_49626,N_49075);
and UO_523 (O_523,N_49515,N_49076);
nand UO_524 (O_524,N_49723,N_49360);
or UO_525 (O_525,N_49730,N_49101);
or UO_526 (O_526,N_49558,N_49836);
nor UO_527 (O_527,N_49806,N_49318);
or UO_528 (O_528,N_49694,N_49355);
nor UO_529 (O_529,N_49310,N_49115);
nand UO_530 (O_530,N_49829,N_49997);
xor UO_531 (O_531,N_49114,N_49575);
xnor UO_532 (O_532,N_49498,N_49434);
nor UO_533 (O_533,N_49145,N_49069);
and UO_534 (O_534,N_49184,N_49928);
nor UO_535 (O_535,N_49476,N_49825);
and UO_536 (O_536,N_49462,N_49643);
nor UO_537 (O_537,N_49626,N_49738);
nor UO_538 (O_538,N_49669,N_49774);
and UO_539 (O_539,N_49784,N_49577);
or UO_540 (O_540,N_49877,N_49389);
and UO_541 (O_541,N_49222,N_49551);
nor UO_542 (O_542,N_49239,N_49853);
and UO_543 (O_543,N_49412,N_49987);
xnor UO_544 (O_544,N_49047,N_49823);
xor UO_545 (O_545,N_49258,N_49584);
nor UO_546 (O_546,N_49253,N_49516);
or UO_547 (O_547,N_49203,N_49824);
and UO_548 (O_548,N_49990,N_49719);
and UO_549 (O_549,N_49740,N_49988);
nor UO_550 (O_550,N_49551,N_49861);
and UO_551 (O_551,N_49297,N_49451);
and UO_552 (O_552,N_49176,N_49573);
or UO_553 (O_553,N_49494,N_49531);
and UO_554 (O_554,N_49063,N_49280);
nand UO_555 (O_555,N_49784,N_49044);
or UO_556 (O_556,N_49589,N_49086);
xnor UO_557 (O_557,N_49888,N_49719);
or UO_558 (O_558,N_49806,N_49662);
or UO_559 (O_559,N_49164,N_49947);
nand UO_560 (O_560,N_49356,N_49607);
nand UO_561 (O_561,N_49754,N_49998);
nand UO_562 (O_562,N_49400,N_49526);
nand UO_563 (O_563,N_49003,N_49557);
xnor UO_564 (O_564,N_49062,N_49185);
xor UO_565 (O_565,N_49685,N_49357);
nand UO_566 (O_566,N_49203,N_49911);
nor UO_567 (O_567,N_49888,N_49734);
nand UO_568 (O_568,N_49554,N_49640);
xor UO_569 (O_569,N_49244,N_49558);
or UO_570 (O_570,N_49385,N_49527);
nand UO_571 (O_571,N_49696,N_49674);
xor UO_572 (O_572,N_49188,N_49736);
or UO_573 (O_573,N_49652,N_49535);
nor UO_574 (O_574,N_49979,N_49176);
or UO_575 (O_575,N_49257,N_49636);
nor UO_576 (O_576,N_49858,N_49145);
xnor UO_577 (O_577,N_49337,N_49699);
and UO_578 (O_578,N_49750,N_49947);
nor UO_579 (O_579,N_49365,N_49140);
xnor UO_580 (O_580,N_49363,N_49807);
xor UO_581 (O_581,N_49895,N_49079);
nor UO_582 (O_582,N_49396,N_49643);
and UO_583 (O_583,N_49723,N_49250);
xor UO_584 (O_584,N_49606,N_49250);
or UO_585 (O_585,N_49001,N_49745);
or UO_586 (O_586,N_49912,N_49082);
nor UO_587 (O_587,N_49798,N_49925);
xor UO_588 (O_588,N_49459,N_49266);
nor UO_589 (O_589,N_49234,N_49939);
and UO_590 (O_590,N_49805,N_49332);
nor UO_591 (O_591,N_49181,N_49108);
nand UO_592 (O_592,N_49044,N_49347);
nand UO_593 (O_593,N_49214,N_49585);
xor UO_594 (O_594,N_49686,N_49790);
nor UO_595 (O_595,N_49741,N_49804);
xor UO_596 (O_596,N_49357,N_49112);
or UO_597 (O_597,N_49458,N_49310);
nand UO_598 (O_598,N_49792,N_49107);
xnor UO_599 (O_599,N_49190,N_49330);
and UO_600 (O_600,N_49097,N_49612);
xnor UO_601 (O_601,N_49130,N_49298);
or UO_602 (O_602,N_49246,N_49702);
and UO_603 (O_603,N_49895,N_49070);
and UO_604 (O_604,N_49509,N_49376);
nand UO_605 (O_605,N_49266,N_49237);
nand UO_606 (O_606,N_49228,N_49928);
nor UO_607 (O_607,N_49782,N_49153);
xor UO_608 (O_608,N_49821,N_49647);
and UO_609 (O_609,N_49744,N_49889);
and UO_610 (O_610,N_49439,N_49086);
and UO_611 (O_611,N_49022,N_49671);
and UO_612 (O_612,N_49830,N_49888);
and UO_613 (O_613,N_49725,N_49268);
or UO_614 (O_614,N_49637,N_49093);
or UO_615 (O_615,N_49499,N_49922);
xor UO_616 (O_616,N_49447,N_49570);
or UO_617 (O_617,N_49373,N_49966);
and UO_618 (O_618,N_49144,N_49094);
xnor UO_619 (O_619,N_49368,N_49327);
xor UO_620 (O_620,N_49112,N_49732);
nand UO_621 (O_621,N_49293,N_49587);
and UO_622 (O_622,N_49394,N_49184);
nand UO_623 (O_623,N_49014,N_49934);
or UO_624 (O_624,N_49452,N_49127);
nand UO_625 (O_625,N_49305,N_49955);
xor UO_626 (O_626,N_49611,N_49704);
or UO_627 (O_627,N_49892,N_49832);
and UO_628 (O_628,N_49125,N_49051);
xnor UO_629 (O_629,N_49802,N_49745);
nand UO_630 (O_630,N_49351,N_49987);
and UO_631 (O_631,N_49911,N_49711);
and UO_632 (O_632,N_49174,N_49472);
and UO_633 (O_633,N_49850,N_49585);
nand UO_634 (O_634,N_49698,N_49347);
and UO_635 (O_635,N_49993,N_49552);
and UO_636 (O_636,N_49147,N_49235);
or UO_637 (O_637,N_49910,N_49696);
nand UO_638 (O_638,N_49074,N_49080);
or UO_639 (O_639,N_49021,N_49582);
or UO_640 (O_640,N_49283,N_49795);
xor UO_641 (O_641,N_49991,N_49281);
nand UO_642 (O_642,N_49798,N_49638);
nand UO_643 (O_643,N_49646,N_49383);
and UO_644 (O_644,N_49627,N_49904);
and UO_645 (O_645,N_49229,N_49573);
nor UO_646 (O_646,N_49388,N_49131);
xor UO_647 (O_647,N_49811,N_49322);
or UO_648 (O_648,N_49086,N_49729);
and UO_649 (O_649,N_49471,N_49816);
and UO_650 (O_650,N_49181,N_49578);
nor UO_651 (O_651,N_49551,N_49558);
xor UO_652 (O_652,N_49043,N_49994);
and UO_653 (O_653,N_49927,N_49523);
or UO_654 (O_654,N_49593,N_49663);
nor UO_655 (O_655,N_49868,N_49198);
xor UO_656 (O_656,N_49492,N_49650);
or UO_657 (O_657,N_49718,N_49488);
and UO_658 (O_658,N_49803,N_49217);
nor UO_659 (O_659,N_49582,N_49626);
and UO_660 (O_660,N_49860,N_49088);
and UO_661 (O_661,N_49082,N_49188);
and UO_662 (O_662,N_49109,N_49628);
or UO_663 (O_663,N_49946,N_49810);
nor UO_664 (O_664,N_49269,N_49725);
nand UO_665 (O_665,N_49336,N_49333);
or UO_666 (O_666,N_49258,N_49084);
or UO_667 (O_667,N_49944,N_49979);
nor UO_668 (O_668,N_49320,N_49588);
and UO_669 (O_669,N_49717,N_49362);
nor UO_670 (O_670,N_49978,N_49619);
and UO_671 (O_671,N_49471,N_49838);
xnor UO_672 (O_672,N_49259,N_49574);
xor UO_673 (O_673,N_49630,N_49519);
nand UO_674 (O_674,N_49212,N_49602);
and UO_675 (O_675,N_49344,N_49449);
or UO_676 (O_676,N_49614,N_49166);
or UO_677 (O_677,N_49118,N_49934);
xnor UO_678 (O_678,N_49416,N_49890);
or UO_679 (O_679,N_49001,N_49348);
xor UO_680 (O_680,N_49361,N_49953);
and UO_681 (O_681,N_49122,N_49032);
and UO_682 (O_682,N_49365,N_49777);
nand UO_683 (O_683,N_49060,N_49503);
xnor UO_684 (O_684,N_49780,N_49035);
nand UO_685 (O_685,N_49271,N_49464);
xor UO_686 (O_686,N_49419,N_49434);
xor UO_687 (O_687,N_49136,N_49590);
nand UO_688 (O_688,N_49232,N_49076);
nor UO_689 (O_689,N_49399,N_49827);
and UO_690 (O_690,N_49059,N_49526);
and UO_691 (O_691,N_49764,N_49262);
nor UO_692 (O_692,N_49213,N_49883);
xnor UO_693 (O_693,N_49057,N_49992);
or UO_694 (O_694,N_49330,N_49448);
and UO_695 (O_695,N_49998,N_49820);
xnor UO_696 (O_696,N_49322,N_49984);
nand UO_697 (O_697,N_49457,N_49829);
and UO_698 (O_698,N_49970,N_49538);
nand UO_699 (O_699,N_49691,N_49062);
xnor UO_700 (O_700,N_49245,N_49888);
or UO_701 (O_701,N_49728,N_49109);
nor UO_702 (O_702,N_49324,N_49248);
nand UO_703 (O_703,N_49075,N_49598);
nand UO_704 (O_704,N_49959,N_49458);
and UO_705 (O_705,N_49432,N_49183);
xnor UO_706 (O_706,N_49955,N_49245);
xnor UO_707 (O_707,N_49113,N_49853);
xnor UO_708 (O_708,N_49337,N_49318);
or UO_709 (O_709,N_49310,N_49067);
or UO_710 (O_710,N_49401,N_49526);
or UO_711 (O_711,N_49340,N_49382);
and UO_712 (O_712,N_49381,N_49674);
nor UO_713 (O_713,N_49292,N_49443);
xnor UO_714 (O_714,N_49852,N_49698);
xnor UO_715 (O_715,N_49868,N_49818);
and UO_716 (O_716,N_49622,N_49399);
xnor UO_717 (O_717,N_49183,N_49402);
or UO_718 (O_718,N_49514,N_49368);
nor UO_719 (O_719,N_49104,N_49812);
nor UO_720 (O_720,N_49880,N_49737);
nor UO_721 (O_721,N_49320,N_49591);
and UO_722 (O_722,N_49763,N_49096);
nand UO_723 (O_723,N_49884,N_49679);
nand UO_724 (O_724,N_49402,N_49936);
xnor UO_725 (O_725,N_49893,N_49195);
and UO_726 (O_726,N_49164,N_49611);
xnor UO_727 (O_727,N_49486,N_49791);
and UO_728 (O_728,N_49287,N_49588);
nor UO_729 (O_729,N_49445,N_49265);
and UO_730 (O_730,N_49618,N_49195);
nor UO_731 (O_731,N_49646,N_49870);
and UO_732 (O_732,N_49713,N_49885);
or UO_733 (O_733,N_49704,N_49553);
or UO_734 (O_734,N_49121,N_49234);
nor UO_735 (O_735,N_49248,N_49445);
nor UO_736 (O_736,N_49575,N_49472);
and UO_737 (O_737,N_49352,N_49125);
or UO_738 (O_738,N_49628,N_49142);
nor UO_739 (O_739,N_49796,N_49712);
or UO_740 (O_740,N_49150,N_49970);
nor UO_741 (O_741,N_49646,N_49303);
nand UO_742 (O_742,N_49359,N_49285);
or UO_743 (O_743,N_49799,N_49857);
and UO_744 (O_744,N_49794,N_49260);
and UO_745 (O_745,N_49979,N_49163);
and UO_746 (O_746,N_49982,N_49015);
or UO_747 (O_747,N_49626,N_49523);
nand UO_748 (O_748,N_49519,N_49492);
nor UO_749 (O_749,N_49203,N_49331);
xor UO_750 (O_750,N_49704,N_49905);
and UO_751 (O_751,N_49100,N_49509);
and UO_752 (O_752,N_49957,N_49363);
and UO_753 (O_753,N_49420,N_49398);
nand UO_754 (O_754,N_49204,N_49983);
xnor UO_755 (O_755,N_49421,N_49045);
xor UO_756 (O_756,N_49764,N_49544);
xnor UO_757 (O_757,N_49369,N_49722);
or UO_758 (O_758,N_49569,N_49957);
nand UO_759 (O_759,N_49256,N_49813);
and UO_760 (O_760,N_49677,N_49970);
xnor UO_761 (O_761,N_49799,N_49920);
or UO_762 (O_762,N_49465,N_49738);
and UO_763 (O_763,N_49921,N_49845);
and UO_764 (O_764,N_49589,N_49375);
xor UO_765 (O_765,N_49734,N_49434);
nor UO_766 (O_766,N_49110,N_49238);
and UO_767 (O_767,N_49098,N_49831);
or UO_768 (O_768,N_49738,N_49093);
xnor UO_769 (O_769,N_49168,N_49574);
xor UO_770 (O_770,N_49714,N_49529);
nor UO_771 (O_771,N_49763,N_49149);
xor UO_772 (O_772,N_49791,N_49188);
and UO_773 (O_773,N_49189,N_49351);
or UO_774 (O_774,N_49989,N_49804);
and UO_775 (O_775,N_49094,N_49071);
and UO_776 (O_776,N_49736,N_49020);
nand UO_777 (O_777,N_49540,N_49734);
xor UO_778 (O_778,N_49002,N_49943);
and UO_779 (O_779,N_49373,N_49593);
or UO_780 (O_780,N_49635,N_49855);
or UO_781 (O_781,N_49255,N_49040);
and UO_782 (O_782,N_49048,N_49032);
or UO_783 (O_783,N_49654,N_49404);
nand UO_784 (O_784,N_49078,N_49204);
and UO_785 (O_785,N_49144,N_49288);
xnor UO_786 (O_786,N_49226,N_49510);
and UO_787 (O_787,N_49333,N_49694);
and UO_788 (O_788,N_49492,N_49777);
or UO_789 (O_789,N_49183,N_49165);
and UO_790 (O_790,N_49130,N_49701);
xnor UO_791 (O_791,N_49136,N_49859);
nor UO_792 (O_792,N_49008,N_49356);
xor UO_793 (O_793,N_49194,N_49005);
and UO_794 (O_794,N_49839,N_49577);
nor UO_795 (O_795,N_49429,N_49558);
nor UO_796 (O_796,N_49872,N_49919);
or UO_797 (O_797,N_49814,N_49101);
and UO_798 (O_798,N_49774,N_49523);
nor UO_799 (O_799,N_49040,N_49364);
or UO_800 (O_800,N_49517,N_49656);
or UO_801 (O_801,N_49534,N_49506);
and UO_802 (O_802,N_49270,N_49826);
and UO_803 (O_803,N_49551,N_49866);
nor UO_804 (O_804,N_49231,N_49781);
and UO_805 (O_805,N_49973,N_49590);
xnor UO_806 (O_806,N_49431,N_49014);
xnor UO_807 (O_807,N_49126,N_49410);
nand UO_808 (O_808,N_49333,N_49506);
nor UO_809 (O_809,N_49508,N_49298);
nor UO_810 (O_810,N_49377,N_49444);
nor UO_811 (O_811,N_49057,N_49364);
or UO_812 (O_812,N_49701,N_49589);
and UO_813 (O_813,N_49449,N_49598);
nor UO_814 (O_814,N_49181,N_49236);
xor UO_815 (O_815,N_49608,N_49722);
nor UO_816 (O_816,N_49055,N_49559);
or UO_817 (O_817,N_49595,N_49756);
xnor UO_818 (O_818,N_49373,N_49675);
or UO_819 (O_819,N_49267,N_49829);
or UO_820 (O_820,N_49717,N_49591);
nand UO_821 (O_821,N_49941,N_49008);
xor UO_822 (O_822,N_49430,N_49949);
nand UO_823 (O_823,N_49976,N_49803);
xor UO_824 (O_824,N_49988,N_49706);
and UO_825 (O_825,N_49433,N_49053);
and UO_826 (O_826,N_49689,N_49597);
or UO_827 (O_827,N_49310,N_49483);
nand UO_828 (O_828,N_49134,N_49396);
xnor UO_829 (O_829,N_49949,N_49201);
xnor UO_830 (O_830,N_49021,N_49944);
xnor UO_831 (O_831,N_49491,N_49354);
nand UO_832 (O_832,N_49187,N_49972);
or UO_833 (O_833,N_49432,N_49491);
nand UO_834 (O_834,N_49710,N_49245);
nand UO_835 (O_835,N_49186,N_49343);
nand UO_836 (O_836,N_49650,N_49051);
xnor UO_837 (O_837,N_49226,N_49330);
xor UO_838 (O_838,N_49873,N_49034);
and UO_839 (O_839,N_49332,N_49375);
or UO_840 (O_840,N_49874,N_49640);
nand UO_841 (O_841,N_49951,N_49245);
nor UO_842 (O_842,N_49890,N_49430);
nand UO_843 (O_843,N_49557,N_49808);
nand UO_844 (O_844,N_49141,N_49233);
xnor UO_845 (O_845,N_49023,N_49460);
or UO_846 (O_846,N_49496,N_49096);
or UO_847 (O_847,N_49708,N_49676);
or UO_848 (O_848,N_49059,N_49154);
and UO_849 (O_849,N_49458,N_49243);
or UO_850 (O_850,N_49043,N_49701);
xor UO_851 (O_851,N_49907,N_49882);
and UO_852 (O_852,N_49242,N_49312);
and UO_853 (O_853,N_49970,N_49338);
nor UO_854 (O_854,N_49974,N_49626);
or UO_855 (O_855,N_49828,N_49724);
or UO_856 (O_856,N_49889,N_49291);
or UO_857 (O_857,N_49607,N_49833);
and UO_858 (O_858,N_49765,N_49294);
nor UO_859 (O_859,N_49250,N_49456);
nor UO_860 (O_860,N_49197,N_49716);
and UO_861 (O_861,N_49453,N_49257);
or UO_862 (O_862,N_49404,N_49014);
and UO_863 (O_863,N_49238,N_49292);
and UO_864 (O_864,N_49864,N_49521);
and UO_865 (O_865,N_49515,N_49785);
and UO_866 (O_866,N_49525,N_49068);
and UO_867 (O_867,N_49043,N_49757);
nand UO_868 (O_868,N_49739,N_49399);
nor UO_869 (O_869,N_49589,N_49552);
and UO_870 (O_870,N_49298,N_49585);
nand UO_871 (O_871,N_49015,N_49250);
nor UO_872 (O_872,N_49882,N_49573);
xnor UO_873 (O_873,N_49166,N_49878);
xnor UO_874 (O_874,N_49646,N_49064);
and UO_875 (O_875,N_49448,N_49261);
and UO_876 (O_876,N_49587,N_49496);
nand UO_877 (O_877,N_49230,N_49179);
nor UO_878 (O_878,N_49242,N_49853);
nand UO_879 (O_879,N_49947,N_49393);
xnor UO_880 (O_880,N_49822,N_49039);
or UO_881 (O_881,N_49179,N_49155);
and UO_882 (O_882,N_49668,N_49835);
and UO_883 (O_883,N_49393,N_49043);
and UO_884 (O_884,N_49550,N_49774);
nor UO_885 (O_885,N_49837,N_49329);
xnor UO_886 (O_886,N_49546,N_49163);
and UO_887 (O_887,N_49669,N_49219);
xor UO_888 (O_888,N_49147,N_49201);
nand UO_889 (O_889,N_49650,N_49657);
nor UO_890 (O_890,N_49427,N_49165);
or UO_891 (O_891,N_49417,N_49977);
and UO_892 (O_892,N_49069,N_49097);
or UO_893 (O_893,N_49528,N_49224);
nand UO_894 (O_894,N_49141,N_49083);
xor UO_895 (O_895,N_49840,N_49229);
nand UO_896 (O_896,N_49990,N_49290);
nor UO_897 (O_897,N_49902,N_49494);
and UO_898 (O_898,N_49786,N_49699);
or UO_899 (O_899,N_49292,N_49471);
or UO_900 (O_900,N_49651,N_49171);
xor UO_901 (O_901,N_49578,N_49997);
nand UO_902 (O_902,N_49156,N_49905);
or UO_903 (O_903,N_49867,N_49495);
xnor UO_904 (O_904,N_49097,N_49618);
and UO_905 (O_905,N_49403,N_49842);
or UO_906 (O_906,N_49689,N_49562);
nor UO_907 (O_907,N_49771,N_49537);
nand UO_908 (O_908,N_49850,N_49488);
and UO_909 (O_909,N_49285,N_49461);
xor UO_910 (O_910,N_49770,N_49478);
nor UO_911 (O_911,N_49805,N_49168);
or UO_912 (O_912,N_49333,N_49905);
or UO_913 (O_913,N_49816,N_49673);
nor UO_914 (O_914,N_49187,N_49847);
and UO_915 (O_915,N_49910,N_49098);
or UO_916 (O_916,N_49521,N_49036);
and UO_917 (O_917,N_49533,N_49326);
and UO_918 (O_918,N_49993,N_49636);
and UO_919 (O_919,N_49365,N_49023);
xnor UO_920 (O_920,N_49343,N_49765);
nand UO_921 (O_921,N_49436,N_49234);
and UO_922 (O_922,N_49233,N_49258);
or UO_923 (O_923,N_49695,N_49310);
nand UO_924 (O_924,N_49554,N_49771);
or UO_925 (O_925,N_49753,N_49611);
or UO_926 (O_926,N_49000,N_49603);
xnor UO_927 (O_927,N_49027,N_49117);
or UO_928 (O_928,N_49650,N_49448);
or UO_929 (O_929,N_49858,N_49421);
or UO_930 (O_930,N_49095,N_49199);
nor UO_931 (O_931,N_49209,N_49608);
nand UO_932 (O_932,N_49881,N_49874);
nor UO_933 (O_933,N_49945,N_49868);
and UO_934 (O_934,N_49961,N_49976);
nand UO_935 (O_935,N_49943,N_49925);
nand UO_936 (O_936,N_49859,N_49234);
nand UO_937 (O_937,N_49609,N_49248);
nand UO_938 (O_938,N_49268,N_49891);
nand UO_939 (O_939,N_49602,N_49721);
xnor UO_940 (O_940,N_49912,N_49092);
xor UO_941 (O_941,N_49323,N_49148);
nor UO_942 (O_942,N_49854,N_49983);
xnor UO_943 (O_943,N_49140,N_49154);
or UO_944 (O_944,N_49299,N_49740);
and UO_945 (O_945,N_49674,N_49852);
or UO_946 (O_946,N_49004,N_49572);
nand UO_947 (O_947,N_49720,N_49638);
nor UO_948 (O_948,N_49349,N_49937);
and UO_949 (O_949,N_49872,N_49651);
xor UO_950 (O_950,N_49095,N_49206);
nor UO_951 (O_951,N_49626,N_49289);
and UO_952 (O_952,N_49344,N_49124);
or UO_953 (O_953,N_49610,N_49671);
and UO_954 (O_954,N_49171,N_49644);
nand UO_955 (O_955,N_49947,N_49223);
nand UO_956 (O_956,N_49582,N_49340);
xnor UO_957 (O_957,N_49140,N_49620);
and UO_958 (O_958,N_49125,N_49123);
xnor UO_959 (O_959,N_49897,N_49465);
or UO_960 (O_960,N_49359,N_49021);
and UO_961 (O_961,N_49996,N_49972);
nor UO_962 (O_962,N_49601,N_49799);
nand UO_963 (O_963,N_49557,N_49209);
and UO_964 (O_964,N_49925,N_49677);
nor UO_965 (O_965,N_49298,N_49354);
xor UO_966 (O_966,N_49090,N_49098);
nor UO_967 (O_967,N_49300,N_49219);
nor UO_968 (O_968,N_49850,N_49242);
and UO_969 (O_969,N_49344,N_49463);
and UO_970 (O_970,N_49532,N_49726);
nor UO_971 (O_971,N_49887,N_49757);
and UO_972 (O_972,N_49370,N_49553);
nand UO_973 (O_973,N_49763,N_49328);
xor UO_974 (O_974,N_49906,N_49933);
nor UO_975 (O_975,N_49412,N_49586);
and UO_976 (O_976,N_49129,N_49366);
xor UO_977 (O_977,N_49009,N_49073);
xor UO_978 (O_978,N_49719,N_49035);
and UO_979 (O_979,N_49319,N_49189);
and UO_980 (O_980,N_49990,N_49171);
and UO_981 (O_981,N_49188,N_49060);
xor UO_982 (O_982,N_49895,N_49291);
nor UO_983 (O_983,N_49105,N_49605);
nand UO_984 (O_984,N_49966,N_49828);
or UO_985 (O_985,N_49868,N_49211);
xnor UO_986 (O_986,N_49749,N_49993);
xnor UO_987 (O_987,N_49281,N_49109);
or UO_988 (O_988,N_49835,N_49285);
and UO_989 (O_989,N_49235,N_49762);
nor UO_990 (O_990,N_49899,N_49912);
nand UO_991 (O_991,N_49120,N_49735);
nand UO_992 (O_992,N_49960,N_49471);
xor UO_993 (O_993,N_49487,N_49390);
and UO_994 (O_994,N_49935,N_49069);
nand UO_995 (O_995,N_49096,N_49388);
nand UO_996 (O_996,N_49467,N_49147);
nand UO_997 (O_997,N_49774,N_49797);
nor UO_998 (O_998,N_49515,N_49017);
and UO_999 (O_999,N_49903,N_49304);
nor UO_1000 (O_1000,N_49537,N_49363);
nand UO_1001 (O_1001,N_49757,N_49955);
or UO_1002 (O_1002,N_49529,N_49023);
xor UO_1003 (O_1003,N_49674,N_49720);
nand UO_1004 (O_1004,N_49998,N_49286);
nand UO_1005 (O_1005,N_49777,N_49503);
nand UO_1006 (O_1006,N_49540,N_49262);
nand UO_1007 (O_1007,N_49680,N_49831);
or UO_1008 (O_1008,N_49705,N_49561);
nand UO_1009 (O_1009,N_49614,N_49935);
xnor UO_1010 (O_1010,N_49918,N_49508);
nand UO_1011 (O_1011,N_49879,N_49322);
nand UO_1012 (O_1012,N_49124,N_49665);
xnor UO_1013 (O_1013,N_49495,N_49730);
and UO_1014 (O_1014,N_49956,N_49678);
nor UO_1015 (O_1015,N_49779,N_49434);
nand UO_1016 (O_1016,N_49688,N_49518);
nand UO_1017 (O_1017,N_49899,N_49746);
nand UO_1018 (O_1018,N_49745,N_49656);
xnor UO_1019 (O_1019,N_49339,N_49952);
or UO_1020 (O_1020,N_49896,N_49713);
or UO_1021 (O_1021,N_49185,N_49768);
nand UO_1022 (O_1022,N_49359,N_49394);
and UO_1023 (O_1023,N_49158,N_49519);
or UO_1024 (O_1024,N_49979,N_49389);
and UO_1025 (O_1025,N_49202,N_49348);
and UO_1026 (O_1026,N_49741,N_49708);
and UO_1027 (O_1027,N_49226,N_49351);
and UO_1028 (O_1028,N_49751,N_49075);
xnor UO_1029 (O_1029,N_49389,N_49613);
and UO_1030 (O_1030,N_49939,N_49460);
nor UO_1031 (O_1031,N_49868,N_49795);
and UO_1032 (O_1032,N_49645,N_49319);
or UO_1033 (O_1033,N_49551,N_49938);
xnor UO_1034 (O_1034,N_49171,N_49970);
nand UO_1035 (O_1035,N_49792,N_49102);
nand UO_1036 (O_1036,N_49785,N_49661);
nand UO_1037 (O_1037,N_49314,N_49747);
nand UO_1038 (O_1038,N_49992,N_49906);
xnor UO_1039 (O_1039,N_49473,N_49182);
and UO_1040 (O_1040,N_49712,N_49646);
or UO_1041 (O_1041,N_49792,N_49985);
xor UO_1042 (O_1042,N_49027,N_49423);
xor UO_1043 (O_1043,N_49234,N_49576);
xor UO_1044 (O_1044,N_49675,N_49215);
and UO_1045 (O_1045,N_49019,N_49715);
xnor UO_1046 (O_1046,N_49311,N_49143);
xor UO_1047 (O_1047,N_49631,N_49300);
and UO_1048 (O_1048,N_49162,N_49821);
xnor UO_1049 (O_1049,N_49892,N_49813);
xor UO_1050 (O_1050,N_49332,N_49950);
nor UO_1051 (O_1051,N_49571,N_49291);
or UO_1052 (O_1052,N_49537,N_49318);
and UO_1053 (O_1053,N_49518,N_49998);
xnor UO_1054 (O_1054,N_49825,N_49048);
xor UO_1055 (O_1055,N_49437,N_49385);
and UO_1056 (O_1056,N_49187,N_49112);
or UO_1057 (O_1057,N_49052,N_49321);
or UO_1058 (O_1058,N_49882,N_49660);
and UO_1059 (O_1059,N_49483,N_49588);
nor UO_1060 (O_1060,N_49054,N_49715);
or UO_1061 (O_1061,N_49478,N_49985);
xor UO_1062 (O_1062,N_49470,N_49165);
and UO_1063 (O_1063,N_49058,N_49065);
and UO_1064 (O_1064,N_49826,N_49711);
nor UO_1065 (O_1065,N_49349,N_49545);
and UO_1066 (O_1066,N_49974,N_49014);
or UO_1067 (O_1067,N_49698,N_49990);
nor UO_1068 (O_1068,N_49058,N_49115);
or UO_1069 (O_1069,N_49047,N_49995);
nor UO_1070 (O_1070,N_49320,N_49128);
nand UO_1071 (O_1071,N_49030,N_49843);
or UO_1072 (O_1072,N_49873,N_49308);
nor UO_1073 (O_1073,N_49291,N_49584);
nand UO_1074 (O_1074,N_49162,N_49331);
nand UO_1075 (O_1075,N_49725,N_49867);
xor UO_1076 (O_1076,N_49480,N_49933);
nor UO_1077 (O_1077,N_49280,N_49589);
nand UO_1078 (O_1078,N_49478,N_49071);
nand UO_1079 (O_1079,N_49655,N_49941);
xnor UO_1080 (O_1080,N_49683,N_49420);
and UO_1081 (O_1081,N_49496,N_49492);
nor UO_1082 (O_1082,N_49710,N_49811);
or UO_1083 (O_1083,N_49746,N_49897);
or UO_1084 (O_1084,N_49814,N_49793);
and UO_1085 (O_1085,N_49526,N_49554);
and UO_1086 (O_1086,N_49358,N_49656);
nand UO_1087 (O_1087,N_49878,N_49094);
nor UO_1088 (O_1088,N_49470,N_49041);
and UO_1089 (O_1089,N_49948,N_49770);
nor UO_1090 (O_1090,N_49460,N_49919);
xor UO_1091 (O_1091,N_49124,N_49916);
nand UO_1092 (O_1092,N_49321,N_49941);
xor UO_1093 (O_1093,N_49564,N_49562);
and UO_1094 (O_1094,N_49635,N_49571);
and UO_1095 (O_1095,N_49038,N_49807);
nand UO_1096 (O_1096,N_49179,N_49461);
nor UO_1097 (O_1097,N_49608,N_49496);
nand UO_1098 (O_1098,N_49422,N_49292);
nor UO_1099 (O_1099,N_49556,N_49384);
and UO_1100 (O_1100,N_49345,N_49214);
or UO_1101 (O_1101,N_49916,N_49490);
nand UO_1102 (O_1102,N_49572,N_49349);
nand UO_1103 (O_1103,N_49754,N_49645);
nand UO_1104 (O_1104,N_49318,N_49991);
nand UO_1105 (O_1105,N_49971,N_49470);
nor UO_1106 (O_1106,N_49444,N_49612);
and UO_1107 (O_1107,N_49951,N_49710);
nand UO_1108 (O_1108,N_49114,N_49083);
nand UO_1109 (O_1109,N_49161,N_49714);
or UO_1110 (O_1110,N_49723,N_49926);
and UO_1111 (O_1111,N_49807,N_49934);
nand UO_1112 (O_1112,N_49366,N_49657);
or UO_1113 (O_1113,N_49825,N_49468);
or UO_1114 (O_1114,N_49088,N_49183);
or UO_1115 (O_1115,N_49402,N_49756);
xor UO_1116 (O_1116,N_49531,N_49978);
xor UO_1117 (O_1117,N_49124,N_49237);
and UO_1118 (O_1118,N_49632,N_49921);
or UO_1119 (O_1119,N_49486,N_49723);
nand UO_1120 (O_1120,N_49924,N_49380);
nor UO_1121 (O_1121,N_49631,N_49183);
xor UO_1122 (O_1122,N_49293,N_49198);
xnor UO_1123 (O_1123,N_49247,N_49807);
nand UO_1124 (O_1124,N_49833,N_49528);
or UO_1125 (O_1125,N_49723,N_49613);
xnor UO_1126 (O_1126,N_49314,N_49499);
and UO_1127 (O_1127,N_49433,N_49700);
or UO_1128 (O_1128,N_49888,N_49709);
nand UO_1129 (O_1129,N_49912,N_49528);
and UO_1130 (O_1130,N_49591,N_49437);
or UO_1131 (O_1131,N_49711,N_49098);
or UO_1132 (O_1132,N_49731,N_49484);
nor UO_1133 (O_1133,N_49121,N_49054);
or UO_1134 (O_1134,N_49778,N_49337);
and UO_1135 (O_1135,N_49423,N_49110);
or UO_1136 (O_1136,N_49968,N_49719);
nor UO_1137 (O_1137,N_49435,N_49206);
nor UO_1138 (O_1138,N_49411,N_49987);
and UO_1139 (O_1139,N_49250,N_49331);
nand UO_1140 (O_1140,N_49839,N_49616);
xor UO_1141 (O_1141,N_49521,N_49292);
nor UO_1142 (O_1142,N_49662,N_49709);
nor UO_1143 (O_1143,N_49103,N_49697);
and UO_1144 (O_1144,N_49171,N_49385);
nor UO_1145 (O_1145,N_49262,N_49191);
and UO_1146 (O_1146,N_49488,N_49846);
and UO_1147 (O_1147,N_49895,N_49844);
or UO_1148 (O_1148,N_49144,N_49307);
xor UO_1149 (O_1149,N_49507,N_49264);
and UO_1150 (O_1150,N_49787,N_49468);
nor UO_1151 (O_1151,N_49514,N_49104);
or UO_1152 (O_1152,N_49875,N_49567);
nand UO_1153 (O_1153,N_49677,N_49937);
and UO_1154 (O_1154,N_49329,N_49401);
xor UO_1155 (O_1155,N_49284,N_49043);
and UO_1156 (O_1156,N_49502,N_49102);
or UO_1157 (O_1157,N_49812,N_49901);
nand UO_1158 (O_1158,N_49458,N_49476);
nand UO_1159 (O_1159,N_49975,N_49992);
and UO_1160 (O_1160,N_49816,N_49589);
nand UO_1161 (O_1161,N_49496,N_49796);
and UO_1162 (O_1162,N_49167,N_49060);
nand UO_1163 (O_1163,N_49813,N_49107);
nor UO_1164 (O_1164,N_49656,N_49648);
nor UO_1165 (O_1165,N_49273,N_49364);
nand UO_1166 (O_1166,N_49671,N_49009);
or UO_1167 (O_1167,N_49968,N_49585);
and UO_1168 (O_1168,N_49054,N_49700);
nand UO_1169 (O_1169,N_49961,N_49817);
nor UO_1170 (O_1170,N_49892,N_49478);
nor UO_1171 (O_1171,N_49013,N_49674);
xnor UO_1172 (O_1172,N_49546,N_49274);
nand UO_1173 (O_1173,N_49271,N_49261);
xor UO_1174 (O_1174,N_49924,N_49413);
nand UO_1175 (O_1175,N_49782,N_49245);
xor UO_1176 (O_1176,N_49140,N_49905);
or UO_1177 (O_1177,N_49703,N_49972);
and UO_1178 (O_1178,N_49121,N_49597);
xor UO_1179 (O_1179,N_49144,N_49599);
xnor UO_1180 (O_1180,N_49209,N_49794);
nand UO_1181 (O_1181,N_49890,N_49279);
or UO_1182 (O_1182,N_49366,N_49740);
or UO_1183 (O_1183,N_49401,N_49825);
or UO_1184 (O_1184,N_49644,N_49258);
nor UO_1185 (O_1185,N_49678,N_49421);
nor UO_1186 (O_1186,N_49918,N_49930);
and UO_1187 (O_1187,N_49769,N_49985);
or UO_1188 (O_1188,N_49613,N_49105);
xnor UO_1189 (O_1189,N_49782,N_49320);
nor UO_1190 (O_1190,N_49827,N_49001);
nand UO_1191 (O_1191,N_49926,N_49355);
nor UO_1192 (O_1192,N_49005,N_49362);
and UO_1193 (O_1193,N_49162,N_49539);
or UO_1194 (O_1194,N_49604,N_49116);
nor UO_1195 (O_1195,N_49803,N_49869);
nor UO_1196 (O_1196,N_49906,N_49032);
nand UO_1197 (O_1197,N_49085,N_49858);
and UO_1198 (O_1198,N_49713,N_49882);
nor UO_1199 (O_1199,N_49827,N_49707);
xor UO_1200 (O_1200,N_49455,N_49267);
and UO_1201 (O_1201,N_49464,N_49684);
and UO_1202 (O_1202,N_49961,N_49627);
xnor UO_1203 (O_1203,N_49236,N_49453);
or UO_1204 (O_1204,N_49148,N_49129);
and UO_1205 (O_1205,N_49603,N_49944);
nor UO_1206 (O_1206,N_49956,N_49784);
and UO_1207 (O_1207,N_49915,N_49340);
xnor UO_1208 (O_1208,N_49584,N_49969);
nand UO_1209 (O_1209,N_49534,N_49077);
and UO_1210 (O_1210,N_49537,N_49391);
nor UO_1211 (O_1211,N_49152,N_49062);
nand UO_1212 (O_1212,N_49265,N_49638);
or UO_1213 (O_1213,N_49268,N_49158);
nand UO_1214 (O_1214,N_49905,N_49370);
and UO_1215 (O_1215,N_49122,N_49937);
xnor UO_1216 (O_1216,N_49537,N_49070);
nor UO_1217 (O_1217,N_49678,N_49448);
and UO_1218 (O_1218,N_49303,N_49744);
xor UO_1219 (O_1219,N_49422,N_49150);
or UO_1220 (O_1220,N_49042,N_49665);
xnor UO_1221 (O_1221,N_49670,N_49985);
nor UO_1222 (O_1222,N_49712,N_49150);
xnor UO_1223 (O_1223,N_49407,N_49207);
and UO_1224 (O_1224,N_49728,N_49554);
nor UO_1225 (O_1225,N_49497,N_49507);
nand UO_1226 (O_1226,N_49377,N_49003);
xnor UO_1227 (O_1227,N_49212,N_49454);
and UO_1228 (O_1228,N_49376,N_49359);
and UO_1229 (O_1229,N_49427,N_49457);
nand UO_1230 (O_1230,N_49968,N_49679);
xor UO_1231 (O_1231,N_49346,N_49356);
and UO_1232 (O_1232,N_49302,N_49180);
nor UO_1233 (O_1233,N_49299,N_49640);
or UO_1234 (O_1234,N_49418,N_49658);
nand UO_1235 (O_1235,N_49734,N_49806);
nor UO_1236 (O_1236,N_49907,N_49799);
xor UO_1237 (O_1237,N_49233,N_49343);
nor UO_1238 (O_1238,N_49743,N_49931);
or UO_1239 (O_1239,N_49129,N_49822);
and UO_1240 (O_1240,N_49621,N_49642);
and UO_1241 (O_1241,N_49049,N_49679);
xor UO_1242 (O_1242,N_49872,N_49315);
nand UO_1243 (O_1243,N_49501,N_49537);
or UO_1244 (O_1244,N_49914,N_49725);
and UO_1245 (O_1245,N_49168,N_49551);
or UO_1246 (O_1246,N_49976,N_49875);
nand UO_1247 (O_1247,N_49948,N_49363);
nor UO_1248 (O_1248,N_49462,N_49638);
or UO_1249 (O_1249,N_49658,N_49184);
and UO_1250 (O_1250,N_49520,N_49371);
nor UO_1251 (O_1251,N_49629,N_49748);
nand UO_1252 (O_1252,N_49991,N_49017);
and UO_1253 (O_1253,N_49125,N_49951);
xnor UO_1254 (O_1254,N_49453,N_49185);
nor UO_1255 (O_1255,N_49312,N_49992);
or UO_1256 (O_1256,N_49782,N_49957);
or UO_1257 (O_1257,N_49970,N_49601);
and UO_1258 (O_1258,N_49278,N_49177);
and UO_1259 (O_1259,N_49868,N_49232);
or UO_1260 (O_1260,N_49230,N_49378);
and UO_1261 (O_1261,N_49258,N_49651);
xnor UO_1262 (O_1262,N_49879,N_49442);
xor UO_1263 (O_1263,N_49827,N_49619);
nor UO_1264 (O_1264,N_49701,N_49386);
or UO_1265 (O_1265,N_49352,N_49414);
or UO_1266 (O_1266,N_49311,N_49405);
or UO_1267 (O_1267,N_49170,N_49861);
nor UO_1268 (O_1268,N_49656,N_49625);
or UO_1269 (O_1269,N_49216,N_49206);
xor UO_1270 (O_1270,N_49275,N_49938);
nor UO_1271 (O_1271,N_49042,N_49585);
xnor UO_1272 (O_1272,N_49672,N_49899);
or UO_1273 (O_1273,N_49287,N_49932);
nand UO_1274 (O_1274,N_49141,N_49055);
xnor UO_1275 (O_1275,N_49025,N_49844);
xor UO_1276 (O_1276,N_49672,N_49190);
nand UO_1277 (O_1277,N_49132,N_49572);
or UO_1278 (O_1278,N_49757,N_49683);
nor UO_1279 (O_1279,N_49110,N_49112);
or UO_1280 (O_1280,N_49218,N_49534);
xor UO_1281 (O_1281,N_49393,N_49312);
or UO_1282 (O_1282,N_49855,N_49999);
xnor UO_1283 (O_1283,N_49300,N_49263);
nand UO_1284 (O_1284,N_49855,N_49576);
xnor UO_1285 (O_1285,N_49029,N_49185);
nand UO_1286 (O_1286,N_49985,N_49341);
nand UO_1287 (O_1287,N_49711,N_49472);
and UO_1288 (O_1288,N_49187,N_49827);
or UO_1289 (O_1289,N_49879,N_49768);
nand UO_1290 (O_1290,N_49734,N_49295);
nand UO_1291 (O_1291,N_49521,N_49246);
xnor UO_1292 (O_1292,N_49836,N_49920);
nand UO_1293 (O_1293,N_49646,N_49883);
nor UO_1294 (O_1294,N_49694,N_49875);
nor UO_1295 (O_1295,N_49779,N_49457);
and UO_1296 (O_1296,N_49780,N_49964);
and UO_1297 (O_1297,N_49408,N_49836);
nand UO_1298 (O_1298,N_49613,N_49092);
xor UO_1299 (O_1299,N_49659,N_49406);
or UO_1300 (O_1300,N_49077,N_49952);
nor UO_1301 (O_1301,N_49338,N_49518);
and UO_1302 (O_1302,N_49905,N_49736);
and UO_1303 (O_1303,N_49628,N_49160);
and UO_1304 (O_1304,N_49250,N_49227);
or UO_1305 (O_1305,N_49125,N_49553);
and UO_1306 (O_1306,N_49296,N_49325);
nor UO_1307 (O_1307,N_49701,N_49258);
nor UO_1308 (O_1308,N_49284,N_49132);
nand UO_1309 (O_1309,N_49165,N_49747);
or UO_1310 (O_1310,N_49040,N_49814);
nor UO_1311 (O_1311,N_49282,N_49871);
xnor UO_1312 (O_1312,N_49952,N_49545);
and UO_1313 (O_1313,N_49245,N_49342);
nand UO_1314 (O_1314,N_49261,N_49467);
and UO_1315 (O_1315,N_49033,N_49849);
or UO_1316 (O_1316,N_49189,N_49958);
nor UO_1317 (O_1317,N_49099,N_49787);
and UO_1318 (O_1318,N_49846,N_49801);
or UO_1319 (O_1319,N_49259,N_49521);
and UO_1320 (O_1320,N_49885,N_49414);
or UO_1321 (O_1321,N_49323,N_49418);
nand UO_1322 (O_1322,N_49602,N_49215);
nor UO_1323 (O_1323,N_49378,N_49844);
or UO_1324 (O_1324,N_49905,N_49092);
and UO_1325 (O_1325,N_49037,N_49921);
or UO_1326 (O_1326,N_49600,N_49260);
nand UO_1327 (O_1327,N_49789,N_49903);
and UO_1328 (O_1328,N_49465,N_49086);
and UO_1329 (O_1329,N_49849,N_49843);
and UO_1330 (O_1330,N_49924,N_49334);
and UO_1331 (O_1331,N_49575,N_49714);
or UO_1332 (O_1332,N_49409,N_49454);
and UO_1333 (O_1333,N_49738,N_49163);
and UO_1334 (O_1334,N_49588,N_49053);
xnor UO_1335 (O_1335,N_49565,N_49304);
and UO_1336 (O_1336,N_49670,N_49581);
xor UO_1337 (O_1337,N_49700,N_49110);
xnor UO_1338 (O_1338,N_49977,N_49503);
nor UO_1339 (O_1339,N_49553,N_49170);
nor UO_1340 (O_1340,N_49912,N_49473);
xor UO_1341 (O_1341,N_49634,N_49659);
and UO_1342 (O_1342,N_49524,N_49695);
nor UO_1343 (O_1343,N_49747,N_49646);
nand UO_1344 (O_1344,N_49472,N_49204);
and UO_1345 (O_1345,N_49088,N_49722);
and UO_1346 (O_1346,N_49377,N_49178);
or UO_1347 (O_1347,N_49080,N_49337);
and UO_1348 (O_1348,N_49433,N_49034);
or UO_1349 (O_1349,N_49668,N_49317);
nor UO_1350 (O_1350,N_49359,N_49527);
or UO_1351 (O_1351,N_49627,N_49168);
xor UO_1352 (O_1352,N_49261,N_49661);
xor UO_1353 (O_1353,N_49467,N_49400);
nand UO_1354 (O_1354,N_49136,N_49881);
xnor UO_1355 (O_1355,N_49277,N_49680);
and UO_1356 (O_1356,N_49950,N_49224);
or UO_1357 (O_1357,N_49701,N_49132);
or UO_1358 (O_1358,N_49797,N_49849);
or UO_1359 (O_1359,N_49502,N_49084);
and UO_1360 (O_1360,N_49241,N_49305);
or UO_1361 (O_1361,N_49420,N_49693);
xor UO_1362 (O_1362,N_49673,N_49315);
and UO_1363 (O_1363,N_49248,N_49109);
or UO_1364 (O_1364,N_49709,N_49498);
nor UO_1365 (O_1365,N_49713,N_49316);
xnor UO_1366 (O_1366,N_49593,N_49950);
or UO_1367 (O_1367,N_49202,N_49908);
nand UO_1368 (O_1368,N_49961,N_49070);
nand UO_1369 (O_1369,N_49090,N_49203);
nor UO_1370 (O_1370,N_49301,N_49610);
and UO_1371 (O_1371,N_49841,N_49676);
and UO_1372 (O_1372,N_49698,N_49819);
xor UO_1373 (O_1373,N_49677,N_49248);
xnor UO_1374 (O_1374,N_49598,N_49939);
nor UO_1375 (O_1375,N_49816,N_49402);
and UO_1376 (O_1376,N_49328,N_49006);
nor UO_1377 (O_1377,N_49443,N_49576);
or UO_1378 (O_1378,N_49600,N_49684);
and UO_1379 (O_1379,N_49244,N_49173);
or UO_1380 (O_1380,N_49905,N_49383);
xor UO_1381 (O_1381,N_49208,N_49474);
nor UO_1382 (O_1382,N_49925,N_49547);
nor UO_1383 (O_1383,N_49277,N_49111);
nor UO_1384 (O_1384,N_49464,N_49312);
nor UO_1385 (O_1385,N_49572,N_49146);
or UO_1386 (O_1386,N_49461,N_49729);
nand UO_1387 (O_1387,N_49445,N_49212);
nand UO_1388 (O_1388,N_49015,N_49574);
or UO_1389 (O_1389,N_49103,N_49110);
xor UO_1390 (O_1390,N_49392,N_49580);
or UO_1391 (O_1391,N_49964,N_49587);
nand UO_1392 (O_1392,N_49481,N_49335);
nand UO_1393 (O_1393,N_49930,N_49216);
nand UO_1394 (O_1394,N_49430,N_49871);
nand UO_1395 (O_1395,N_49901,N_49516);
nand UO_1396 (O_1396,N_49062,N_49596);
and UO_1397 (O_1397,N_49472,N_49262);
xor UO_1398 (O_1398,N_49897,N_49596);
or UO_1399 (O_1399,N_49597,N_49996);
or UO_1400 (O_1400,N_49926,N_49717);
and UO_1401 (O_1401,N_49477,N_49942);
or UO_1402 (O_1402,N_49887,N_49680);
xnor UO_1403 (O_1403,N_49743,N_49042);
xnor UO_1404 (O_1404,N_49561,N_49122);
or UO_1405 (O_1405,N_49694,N_49645);
nand UO_1406 (O_1406,N_49229,N_49401);
or UO_1407 (O_1407,N_49343,N_49080);
xnor UO_1408 (O_1408,N_49593,N_49875);
nand UO_1409 (O_1409,N_49916,N_49652);
or UO_1410 (O_1410,N_49059,N_49765);
or UO_1411 (O_1411,N_49517,N_49357);
xnor UO_1412 (O_1412,N_49263,N_49087);
or UO_1413 (O_1413,N_49562,N_49980);
or UO_1414 (O_1414,N_49311,N_49381);
xor UO_1415 (O_1415,N_49019,N_49879);
nor UO_1416 (O_1416,N_49858,N_49362);
nor UO_1417 (O_1417,N_49796,N_49689);
xnor UO_1418 (O_1418,N_49178,N_49640);
nor UO_1419 (O_1419,N_49142,N_49233);
or UO_1420 (O_1420,N_49184,N_49067);
and UO_1421 (O_1421,N_49720,N_49642);
nor UO_1422 (O_1422,N_49449,N_49712);
nand UO_1423 (O_1423,N_49693,N_49413);
nand UO_1424 (O_1424,N_49413,N_49406);
nand UO_1425 (O_1425,N_49146,N_49314);
and UO_1426 (O_1426,N_49862,N_49587);
nor UO_1427 (O_1427,N_49679,N_49328);
and UO_1428 (O_1428,N_49265,N_49014);
nor UO_1429 (O_1429,N_49420,N_49908);
nand UO_1430 (O_1430,N_49592,N_49674);
or UO_1431 (O_1431,N_49057,N_49378);
and UO_1432 (O_1432,N_49226,N_49534);
nor UO_1433 (O_1433,N_49110,N_49980);
or UO_1434 (O_1434,N_49147,N_49193);
nand UO_1435 (O_1435,N_49671,N_49795);
nand UO_1436 (O_1436,N_49709,N_49969);
xor UO_1437 (O_1437,N_49143,N_49402);
xnor UO_1438 (O_1438,N_49699,N_49408);
or UO_1439 (O_1439,N_49672,N_49083);
or UO_1440 (O_1440,N_49940,N_49858);
and UO_1441 (O_1441,N_49976,N_49884);
or UO_1442 (O_1442,N_49106,N_49291);
xnor UO_1443 (O_1443,N_49676,N_49978);
xor UO_1444 (O_1444,N_49441,N_49465);
nor UO_1445 (O_1445,N_49788,N_49520);
or UO_1446 (O_1446,N_49789,N_49248);
nor UO_1447 (O_1447,N_49897,N_49315);
or UO_1448 (O_1448,N_49056,N_49683);
nor UO_1449 (O_1449,N_49987,N_49824);
nor UO_1450 (O_1450,N_49037,N_49083);
or UO_1451 (O_1451,N_49806,N_49419);
nor UO_1452 (O_1452,N_49842,N_49542);
and UO_1453 (O_1453,N_49170,N_49885);
nand UO_1454 (O_1454,N_49402,N_49372);
xnor UO_1455 (O_1455,N_49121,N_49236);
nor UO_1456 (O_1456,N_49401,N_49836);
and UO_1457 (O_1457,N_49088,N_49158);
nor UO_1458 (O_1458,N_49138,N_49312);
nor UO_1459 (O_1459,N_49522,N_49591);
nand UO_1460 (O_1460,N_49067,N_49629);
nand UO_1461 (O_1461,N_49545,N_49350);
and UO_1462 (O_1462,N_49778,N_49299);
xor UO_1463 (O_1463,N_49742,N_49481);
xnor UO_1464 (O_1464,N_49279,N_49968);
and UO_1465 (O_1465,N_49732,N_49168);
or UO_1466 (O_1466,N_49625,N_49060);
nor UO_1467 (O_1467,N_49037,N_49739);
or UO_1468 (O_1468,N_49777,N_49550);
nor UO_1469 (O_1469,N_49175,N_49379);
nand UO_1470 (O_1470,N_49958,N_49237);
or UO_1471 (O_1471,N_49524,N_49645);
and UO_1472 (O_1472,N_49919,N_49602);
xnor UO_1473 (O_1473,N_49301,N_49313);
and UO_1474 (O_1474,N_49440,N_49272);
and UO_1475 (O_1475,N_49532,N_49599);
or UO_1476 (O_1476,N_49977,N_49422);
nor UO_1477 (O_1477,N_49215,N_49870);
nand UO_1478 (O_1478,N_49897,N_49679);
or UO_1479 (O_1479,N_49573,N_49134);
and UO_1480 (O_1480,N_49019,N_49283);
nand UO_1481 (O_1481,N_49557,N_49904);
and UO_1482 (O_1482,N_49865,N_49450);
or UO_1483 (O_1483,N_49542,N_49722);
nand UO_1484 (O_1484,N_49280,N_49990);
xor UO_1485 (O_1485,N_49105,N_49725);
and UO_1486 (O_1486,N_49866,N_49405);
or UO_1487 (O_1487,N_49176,N_49733);
and UO_1488 (O_1488,N_49855,N_49585);
xnor UO_1489 (O_1489,N_49237,N_49475);
nor UO_1490 (O_1490,N_49939,N_49250);
nand UO_1491 (O_1491,N_49321,N_49427);
nand UO_1492 (O_1492,N_49187,N_49854);
nand UO_1493 (O_1493,N_49958,N_49355);
and UO_1494 (O_1494,N_49519,N_49971);
xnor UO_1495 (O_1495,N_49775,N_49767);
nor UO_1496 (O_1496,N_49210,N_49096);
nor UO_1497 (O_1497,N_49804,N_49731);
or UO_1498 (O_1498,N_49686,N_49013);
nor UO_1499 (O_1499,N_49984,N_49619);
xor UO_1500 (O_1500,N_49258,N_49252);
nand UO_1501 (O_1501,N_49950,N_49633);
and UO_1502 (O_1502,N_49832,N_49310);
nor UO_1503 (O_1503,N_49158,N_49892);
or UO_1504 (O_1504,N_49284,N_49172);
and UO_1505 (O_1505,N_49268,N_49422);
and UO_1506 (O_1506,N_49551,N_49536);
nand UO_1507 (O_1507,N_49217,N_49030);
nor UO_1508 (O_1508,N_49712,N_49724);
xor UO_1509 (O_1509,N_49436,N_49127);
and UO_1510 (O_1510,N_49085,N_49366);
nor UO_1511 (O_1511,N_49792,N_49372);
xnor UO_1512 (O_1512,N_49766,N_49126);
nor UO_1513 (O_1513,N_49817,N_49774);
and UO_1514 (O_1514,N_49078,N_49762);
and UO_1515 (O_1515,N_49321,N_49383);
nand UO_1516 (O_1516,N_49505,N_49868);
nand UO_1517 (O_1517,N_49721,N_49447);
nand UO_1518 (O_1518,N_49166,N_49414);
nor UO_1519 (O_1519,N_49997,N_49082);
and UO_1520 (O_1520,N_49202,N_49033);
nor UO_1521 (O_1521,N_49156,N_49759);
nand UO_1522 (O_1522,N_49314,N_49851);
or UO_1523 (O_1523,N_49377,N_49865);
nand UO_1524 (O_1524,N_49869,N_49680);
and UO_1525 (O_1525,N_49535,N_49458);
or UO_1526 (O_1526,N_49533,N_49902);
xor UO_1527 (O_1527,N_49650,N_49653);
xor UO_1528 (O_1528,N_49925,N_49073);
nand UO_1529 (O_1529,N_49416,N_49634);
xnor UO_1530 (O_1530,N_49421,N_49328);
nor UO_1531 (O_1531,N_49768,N_49951);
nand UO_1532 (O_1532,N_49719,N_49251);
or UO_1533 (O_1533,N_49835,N_49972);
nor UO_1534 (O_1534,N_49537,N_49065);
and UO_1535 (O_1535,N_49056,N_49575);
xnor UO_1536 (O_1536,N_49743,N_49052);
nand UO_1537 (O_1537,N_49192,N_49985);
nor UO_1538 (O_1538,N_49258,N_49529);
nor UO_1539 (O_1539,N_49550,N_49020);
nor UO_1540 (O_1540,N_49357,N_49733);
nor UO_1541 (O_1541,N_49556,N_49982);
and UO_1542 (O_1542,N_49804,N_49517);
nand UO_1543 (O_1543,N_49011,N_49498);
and UO_1544 (O_1544,N_49305,N_49411);
nor UO_1545 (O_1545,N_49270,N_49053);
xor UO_1546 (O_1546,N_49037,N_49487);
nand UO_1547 (O_1547,N_49019,N_49575);
xor UO_1548 (O_1548,N_49159,N_49986);
nand UO_1549 (O_1549,N_49333,N_49126);
and UO_1550 (O_1550,N_49656,N_49200);
nand UO_1551 (O_1551,N_49106,N_49993);
xnor UO_1552 (O_1552,N_49720,N_49670);
xnor UO_1553 (O_1553,N_49393,N_49555);
or UO_1554 (O_1554,N_49019,N_49406);
nor UO_1555 (O_1555,N_49268,N_49686);
or UO_1556 (O_1556,N_49485,N_49695);
xnor UO_1557 (O_1557,N_49220,N_49077);
or UO_1558 (O_1558,N_49340,N_49848);
nor UO_1559 (O_1559,N_49287,N_49798);
nor UO_1560 (O_1560,N_49175,N_49673);
xor UO_1561 (O_1561,N_49868,N_49574);
or UO_1562 (O_1562,N_49470,N_49533);
nor UO_1563 (O_1563,N_49683,N_49595);
or UO_1564 (O_1564,N_49803,N_49075);
nor UO_1565 (O_1565,N_49300,N_49324);
nand UO_1566 (O_1566,N_49761,N_49545);
nand UO_1567 (O_1567,N_49912,N_49894);
nor UO_1568 (O_1568,N_49669,N_49294);
and UO_1569 (O_1569,N_49781,N_49091);
or UO_1570 (O_1570,N_49276,N_49656);
or UO_1571 (O_1571,N_49403,N_49206);
xor UO_1572 (O_1572,N_49748,N_49724);
xnor UO_1573 (O_1573,N_49689,N_49410);
xnor UO_1574 (O_1574,N_49261,N_49764);
xnor UO_1575 (O_1575,N_49634,N_49708);
xor UO_1576 (O_1576,N_49166,N_49902);
xor UO_1577 (O_1577,N_49702,N_49252);
nor UO_1578 (O_1578,N_49701,N_49887);
and UO_1579 (O_1579,N_49711,N_49873);
or UO_1580 (O_1580,N_49059,N_49494);
nor UO_1581 (O_1581,N_49959,N_49086);
nor UO_1582 (O_1582,N_49133,N_49267);
or UO_1583 (O_1583,N_49691,N_49221);
nor UO_1584 (O_1584,N_49067,N_49881);
nor UO_1585 (O_1585,N_49787,N_49250);
xor UO_1586 (O_1586,N_49447,N_49083);
nor UO_1587 (O_1587,N_49129,N_49723);
and UO_1588 (O_1588,N_49393,N_49357);
nor UO_1589 (O_1589,N_49883,N_49108);
xor UO_1590 (O_1590,N_49921,N_49272);
nor UO_1591 (O_1591,N_49333,N_49717);
and UO_1592 (O_1592,N_49663,N_49636);
nor UO_1593 (O_1593,N_49343,N_49407);
or UO_1594 (O_1594,N_49278,N_49031);
xor UO_1595 (O_1595,N_49865,N_49640);
xnor UO_1596 (O_1596,N_49019,N_49682);
nand UO_1597 (O_1597,N_49459,N_49201);
and UO_1598 (O_1598,N_49774,N_49065);
and UO_1599 (O_1599,N_49886,N_49020);
xnor UO_1600 (O_1600,N_49101,N_49245);
nor UO_1601 (O_1601,N_49850,N_49325);
and UO_1602 (O_1602,N_49662,N_49553);
or UO_1603 (O_1603,N_49090,N_49773);
xnor UO_1604 (O_1604,N_49757,N_49928);
nor UO_1605 (O_1605,N_49741,N_49021);
xor UO_1606 (O_1606,N_49984,N_49588);
or UO_1607 (O_1607,N_49560,N_49998);
nor UO_1608 (O_1608,N_49424,N_49851);
nand UO_1609 (O_1609,N_49626,N_49013);
or UO_1610 (O_1610,N_49881,N_49248);
nor UO_1611 (O_1611,N_49736,N_49055);
xor UO_1612 (O_1612,N_49464,N_49723);
xnor UO_1613 (O_1613,N_49079,N_49388);
nor UO_1614 (O_1614,N_49508,N_49880);
or UO_1615 (O_1615,N_49964,N_49692);
nand UO_1616 (O_1616,N_49201,N_49975);
nand UO_1617 (O_1617,N_49132,N_49114);
and UO_1618 (O_1618,N_49281,N_49721);
or UO_1619 (O_1619,N_49958,N_49557);
or UO_1620 (O_1620,N_49610,N_49790);
xnor UO_1621 (O_1621,N_49437,N_49539);
and UO_1622 (O_1622,N_49203,N_49601);
xor UO_1623 (O_1623,N_49568,N_49823);
nor UO_1624 (O_1624,N_49364,N_49578);
and UO_1625 (O_1625,N_49437,N_49187);
and UO_1626 (O_1626,N_49273,N_49211);
or UO_1627 (O_1627,N_49386,N_49844);
and UO_1628 (O_1628,N_49022,N_49845);
or UO_1629 (O_1629,N_49257,N_49829);
or UO_1630 (O_1630,N_49140,N_49911);
or UO_1631 (O_1631,N_49909,N_49929);
and UO_1632 (O_1632,N_49610,N_49984);
xnor UO_1633 (O_1633,N_49638,N_49687);
xor UO_1634 (O_1634,N_49597,N_49788);
and UO_1635 (O_1635,N_49837,N_49346);
or UO_1636 (O_1636,N_49178,N_49039);
or UO_1637 (O_1637,N_49648,N_49239);
and UO_1638 (O_1638,N_49471,N_49876);
and UO_1639 (O_1639,N_49855,N_49562);
nor UO_1640 (O_1640,N_49656,N_49790);
and UO_1641 (O_1641,N_49355,N_49004);
nor UO_1642 (O_1642,N_49801,N_49486);
or UO_1643 (O_1643,N_49208,N_49514);
xor UO_1644 (O_1644,N_49173,N_49631);
or UO_1645 (O_1645,N_49905,N_49138);
nor UO_1646 (O_1646,N_49265,N_49453);
and UO_1647 (O_1647,N_49572,N_49284);
and UO_1648 (O_1648,N_49756,N_49459);
or UO_1649 (O_1649,N_49113,N_49593);
nor UO_1650 (O_1650,N_49272,N_49116);
nand UO_1651 (O_1651,N_49692,N_49725);
xor UO_1652 (O_1652,N_49622,N_49995);
and UO_1653 (O_1653,N_49707,N_49039);
and UO_1654 (O_1654,N_49044,N_49718);
xnor UO_1655 (O_1655,N_49052,N_49223);
nor UO_1656 (O_1656,N_49665,N_49539);
nand UO_1657 (O_1657,N_49669,N_49877);
nor UO_1658 (O_1658,N_49950,N_49976);
xor UO_1659 (O_1659,N_49959,N_49500);
nand UO_1660 (O_1660,N_49247,N_49610);
and UO_1661 (O_1661,N_49044,N_49147);
nor UO_1662 (O_1662,N_49207,N_49648);
xor UO_1663 (O_1663,N_49383,N_49753);
nor UO_1664 (O_1664,N_49992,N_49744);
nor UO_1665 (O_1665,N_49099,N_49311);
or UO_1666 (O_1666,N_49485,N_49680);
and UO_1667 (O_1667,N_49963,N_49432);
nand UO_1668 (O_1668,N_49521,N_49127);
xnor UO_1669 (O_1669,N_49765,N_49416);
xnor UO_1670 (O_1670,N_49482,N_49803);
nand UO_1671 (O_1671,N_49743,N_49001);
nand UO_1672 (O_1672,N_49171,N_49423);
xor UO_1673 (O_1673,N_49460,N_49680);
nand UO_1674 (O_1674,N_49487,N_49322);
xnor UO_1675 (O_1675,N_49009,N_49577);
xnor UO_1676 (O_1676,N_49114,N_49674);
nor UO_1677 (O_1677,N_49251,N_49098);
or UO_1678 (O_1678,N_49098,N_49477);
or UO_1679 (O_1679,N_49231,N_49442);
and UO_1680 (O_1680,N_49882,N_49517);
or UO_1681 (O_1681,N_49020,N_49524);
or UO_1682 (O_1682,N_49018,N_49678);
xnor UO_1683 (O_1683,N_49095,N_49063);
xnor UO_1684 (O_1684,N_49958,N_49491);
and UO_1685 (O_1685,N_49756,N_49023);
nor UO_1686 (O_1686,N_49636,N_49208);
nand UO_1687 (O_1687,N_49289,N_49758);
nand UO_1688 (O_1688,N_49454,N_49509);
nor UO_1689 (O_1689,N_49008,N_49297);
nor UO_1690 (O_1690,N_49625,N_49655);
nor UO_1691 (O_1691,N_49106,N_49242);
nor UO_1692 (O_1692,N_49102,N_49056);
nor UO_1693 (O_1693,N_49697,N_49902);
xor UO_1694 (O_1694,N_49153,N_49427);
or UO_1695 (O_1695,N_49201,N_49029);
nor UO_1696 (O_1696,N_49193,N_49358);
xor UO_1697 (O_1697,N_49840,N_49332);
nand UO_1698 (O_1698,N_49111,N_49734);
nand UO_1699 (O_1699,N_49070,N_49597);
or UO_1700 (O_1700,N_49561,N_49074);
and UO_1701 (O_1701,N_49495,N_49348);
nand UO_1702 (O_1702,N_49306,N_49281);
nor UO_1703 (O_1703,N_49981,N_49008);
and UO_1704 (O_1704,N_49296,N_49021);
nand UO_1705 (O_1705,N_49224,N_49561);
and UO_1706 (O_1706,N_49452,N_49955);
and UO_1707 (O_1707,N_49430,N_49798);
xor UO_1708 (O_1708,N_49815,N_49120);
xnor UO_1709 (O_1709,N_49217,N_49986);
nor UO_1710 (O_1710,N_49874,N_49897);
or UO_1711 (O_1711,N_49815,N_49476);
nand UO_1712 (O_1712,N_49650,N_49207);
nand UO_1713 (O_1713,N_49835,N_49819);
nor UO_1714 (O_1714,N_49558,N_49206);
nor UO_1715 (O_1715,N_49366,N_49535);
and UO_1716 (O_1716,N_49586,N_49718);
and UO_1717 (O_1717,N_49077,N_49848);
xor UO_1718 (O_1718,N_49951,N_49260);
or UO_1719 (O_1719,N_49623,N_49909);
and UO_1720 (O_1720,N_49895,N_49065);
and UO_1721 (O_1721,N_49535,N_49330);
xor UO_1722 (O_1722,N_49839,N_49874);
or UO_1723 (O_1723,N_49764,N_49178);
nor UO_1724 (O_1724,N_49790,N_49812);
nand UO_1725 (O_1725,N_49837,N_49630);
or UO_1726 (O_1726,N_49932,N_49469);
and UO_1727 (O_1727,N_49383,N_49730);
or UO_1728 (O_1728,N_49941,N_49259);
and UO_1729 (O_1729,N_49479,N_49142);
nor UO_1730 (O_1730,N_49978,N_49595);
xnor UO_1731 (O_1731,N_49852,N_49954);
xnor UO_1732 (O_1732,N_49318,N_49036);
nand UO_1733 (O_1733,N_49686,N_49887);
nand UO_1734 (O_1734,N_49244,N_49207);
and UO_1735 (O_1735,N_49037,N_49466);
and UO_1736 (O_1736,N_49188,N_49875);
xor UO_1737 (O_1737,N_49433,N_49557);
and UO_1738 (O_1738,N_49346,N_49641);
nand UO_1739 (O_1739,N_49190,N_49872);
nor UO_1740 (O_1740,N_49993,N_49870);
nand UO_1741 (O_1741,N_49181,N_49429);
or UO_1742 (O_1742,N_49406,N_49633);
or UO_1743 (O_1743,N_49510,N_49190);
nor UO_1744 (O_1744,N_49725,N_49846);
nand UO_1745 (O_1745,N_49758,N_49867);
xnor UO_1746 (O_1746,N_49787,N_49781);
and UO_1747 (O_1747,N_49293,N_49616);
nand UO_1748 (O_1748,N_49786,N_49872);
nor UO_1749 (O_1749,N_49605,N_49266);
and UO_1750 (O_1750,N_49360,N_49025);
and UO_1751 (O_1751,N_49420,N_49776);
nand UO_1752 (O_1752,N_49500,N_49371);
and UO_1753 (O_1753,N_49549,N_49299);
or UO_1754 (O_1754,N_49881,N_49261);
and UO_1755 (O_1755,N_49624,N_49226);
xor UO_1756 (O_1756,N_49609,N_49828);
xor UO_1757 (O_1757,N_49879,N_49224);
xor UO_1758 (O_1758,N_49218,N_49331);
or UO_1759 (O_1759,N_49661,N_49403);
nand UO_1760 (O_1760,N_49120,N_49149);
nand UO_1761 (O_1761,N_49828,N_49007);
nand UO_1762 (O_1762,N_49695,N_49777);
and UO_1763 (O_1763,N_49141,N_49693);
and UO_1764 (O_1764,N_49348,N_49329);
nand UO_1765 (O_1765,N_49334,N_49014);
or UO_1766 (O_1766,N_49249,N_49889);
and UO_1767 (O_1767,N_49175,N_49622);
nand UO_1768 (O_1768,N_49329,N_49573);
or UO_1769 (O_1769,N_49243,N_49365);
xor UO_1770 (O_1770,N_49231,N_49925);
nand UO_1771 (O_1771,N_49917,N_49559);
or UO_1772 (O_1772,N_49572,N_49075);
nor UO_1773 (O_1773,N_49861,N_49572);
nand UO_1774 (O_1774,N_49632,N_49488);
nand UO_1775 (O_1775,N_49637,N_49514);
nor UO_1776 (O_1776,N_49845,N_49410);
nor UO_1777 (O_1777,N_49506,N_49801);
and UO_1778 (O_1778,N_49675,N_49666);
xnor UO_1779 (O_1779,N_49201,N_49999);
nor UO_1780 (O_1780,N_49951,N_49381);
xnor UO_1781 (O_1781,N_49639,N_49188);
nand UO_1782 (O_1782,N_49326,N_49265);
nand UO_1783 (O_1783,N_49719,N_49655);
or UO_1784 (O_1784,N_49071,N_49318);
nor UO_1785 (O_1785,N_49745,N_49803);
nand UO_1786 (O_1786,N_49088,N_49846);
nand UO_1787 (O_1787,N_49263,N_49544);
and UO_1788 (O_1788,N_49451,N_49740);
or UO_1789 (O_1789,N_49581,N_49313);
or UO_1790 (O_1790,N_49296,N_49365);
nor UO_1791 (O_1791,N_49156,N_49963);
nor UO_1792 (O_1792,N_49817,N_49014);
and UO_1793 (O_1793,N_49019,N_49610);
nand UO_1794 (O_1794,N_49260,N_49134);
or UO_1795 (O_1795,N_49861,N_49561);
nand UO_1796 (O_1796,N_49330,N_49611);
xor UO_1797 (O_1797,N_49632,N_49766);
and UO_1798 (O_1798,N_49718,N_49030);
xnor UO_1799 (O_1799,N_49741,N_49270);
and UO_1800 (O_1800,N_49534,N_49225);
or UO_1801 (O_1801,N_49942,N_49379);
nor UO_1802 (O_1802,N_49614,N_49162);
nor UO_1803 (O_1803,N_49213,N_49261);
or UO_1804 (O_1804,N_49706,N_49975);
nand UO_1805 (O_1805,N_49849,N_49425);
and UO_1806 (O_1806,N_49762,N_49111);
nand UO_1807 (O_1807,N_49851,N_49649);
xor UO_1808 (O_1808,N_49250,N_49851);
and UO_1809 (O_1809,N_49991,N_49011);
and UO_1810 (O_1810,N_49659,N_49745);
or UO_1811 (O_1811,N_49945,N_49500);
nor UO_1812 (O_1812,N_49105,N_49511);
or UO_1813 (O_1813,N_49700,N_49995);
xnor UO_1814 (O_1814,N_49353,N_49116);
xnor UO_1815 (O_1815,N_49854,N_49668);
xnor UO_1816 (O_1816,N_49385,N_49516);
nand UO_1817 (O_1817,N_49208,N_49732);
or UO_1818 (O_1818,N_49203,N_49821);
xnor UO_1819 (O_1819,N_49342,N_49887);
nand UO_1820 (O_1820,N_49414,N_49163);
nor UO_1821 (O_1821,N_49908,N_49323);
xnor UO_1822 (O_1822,N_49414,N_49186);
nand UO_1823 (O_1823,N_49915,N_49319);
and UO_1824 (O_1824,N_49855,N_49243);
nand UO_1825 (O_1825,N_49634,N_49459);
nor UO_1826 (O_1826,N_49287,N_49114);
nand UO_1827 (O_1827,N_49244,N_49586);
or UO_1828 (O_1828,N_49448,N_49051);
and UO_1829 (O_1829,N_49676,N_49964);
and UO_1830 (O_1830,N_49094,N_49315);
xor UO_1831 (O_1831,N_49214,N_49396);
and UO_1832 (O_1832,N_49117,N_49666);
and UO_1833 (O_1833,N_49296,N_49371);
nand UO_1834 (O_1834,N_49637,N_49465);
nor UO_1835 (O_1835,N_49526,N_49751);
and UO_1836 (O_1836,N_49035,N_49313);
nor UO_1837 (O_1837,N_49141,N_49558);
xor UO_1838 (O_1838,N_49860,N_49450);
and UO_1839 (O_1839,N_49911,N_49648);
or UO_1840 (O_1840,N_49591,N_49746);
nand UO_1841 (O_1841,N_49404,N_49737);
or UO_1842 (O_1842,N_49522,N_49066);
nor UO_1843 (O_1843,N_49627,N_49978);
or UO_1844 (O_1844,N_49828,N_49498);
xnor UO_1845 (O_1845,N_49273,N_49315);
and UO_1846 (O_1846,N_49809,N_49352);
nand UO_1847 (O_1847,N_49307,N_49383);
and UO_1848 (O_1848,N_49977,N_49458);
xor UO_1849 (O_1849,N_49877,N_49908);
or UO_1850 (O_1850,N_49167,N_49873);
nor UO_1851 (O_1851,N_49927,N_49535);
nand UO_1852 (O_1852,N_49082,N_49774);
nor UO_1853 (O_1853,N_49061,N_49147);
xor UO_1854 (O_1854,N_49353,N_49609);
nor UO_1855 (O_1855,N_49522,N_49410);
and UO_1856 (O_1856,N_49108,N_49017);
nor UO_1857 (O_1857,N_49846,N_49963);
or UO_1858 (O_1858,N_49864,N_49420);
nor UO_1859 (O_1859,N_49962,N_49343);
and UO_1860 (O_1860,N_49115,N_49526);
nand UO_1861 (O_1861,N_49038,N_49317);
or UO_1862 (O_1862,N_49520,N_49955);
nand UO_1863 (O_1863,N_49285,N_49952);
nor UO_1864 (O_1864,N_49372,N_49424);
nand UO_1865 (O_1865,N_49346,N_49245);
xnor UO_1866 (O_1866,N_49565,N_49445);
nand UO_1867 (O_1867,N_49829,N_49270);
or UO_1868 (O_1868,N_49600,N_49873);
xor UO_1869 (O_1869,N_49405,N_49957);
xor UO_1870 (O_1870,N_49924,N_49292);
xnor UO_1871 (O_1871,N_49587,N_49731);
xnor UO_1872 (O_1872,N_49934,N_49575);
and UO_1873 (O_1873,N_49325,N_49547);
xnor UO_1874 (O_1874,N_49534,N_49694);
nand UO_1875 (O_1875,N_49770,N_49730);
nand UO_1876 (O_1876,N_49929,N_49348);
xor UO_1877 (O_1877,N_49847,N_49362);
or UO_1878 (O_1878,N_49290,N_49239);
xnor UO_1879 (O_1879,N_49115,N_49190);
nor UO_1880 (O_1880,N_49335,N_49093);
or UO_1881 (O_1881,N_49865,N_49255);
nand UO_1882 (O_1882,N_49484,N_49282);
nand UO_1883 (O_1883,N_49838,N_49567);
and UO_1884 (O_1884,N_49507,N_49874);
nand UO_1885 (O_1885,N_49357,N_49919);
nand UO_1886 (O_1886,N_49770,N_49257);
nand UO_1887 (O_1887,N_49287,N_49339);
and UO_1888 (O_1888,N_49306,N_49098);
and UO_1889 (O_1889,N_49453,N_49808);
xor UO_1890 (O_1890,N_49057,N_49377);
xor UO_1891 (O_1891,N_49862,N_49176);
or UO_1892 (O_1892,N_49771,N_49193);
xnor UO_1893 (O_1893,N_49448,N_49739);
nor UO_1894 (O_1894,N_49042,N_49183);
nor UO_1895 (O_1895,N_49825,N_49524);
or UO_1896 (O_1896,N_49934,N_49130);
or UO_1897 (O_1897,N_49840,N_49031);
or UO_1898 (O_1898,N_49640,N_49149);
or UO_1899 (O_1899,N_49365,N_49268);
or UO_1900 (O_1900,N_49394,N_49173);
xnor UO_1901 (O_1901,N_49977,N_49016);
xnor UO_1902 (O_1902,N_49621,N_49438);
or UO_1903 (O_1903,N_49616,N_49420);
xor UO_1904 (O_1904,N_49031,N_49579);
nor UO_1905 (O_1905,N_49643,N_49004);
and UO_1906 (O_1906,N_49258,N_49897);
nand UO_1907 (O_1907,N_49302,N_49785);
nor UO_1908 (O_1908,N_49641,N_49564);
nor UO_1909 (O_1909,N_49435,N_49903);
and UO_1910 (O_1910,N_49053,N_49517);
xor UO_1911 (O_1911,N_49740,N_49907);
and UO_1912 (O_1912,N_49387,N_49564);
and UO_1913 (O_1913,N_49409,N_49688);
nand UO_1914 (O_1914,N_49760,N_49956);
or UO_1915 (O_1915,N_49362,N_49003);
or UO_1916 (O_1916,N_49199,N_49659);
and UO_1917 (O_1917,N_49373,N_49776);
nor UO_1918 (O_1918,N_49149,N_49237);
xor UO_1919 (O_1919,N_49964,N_49562);
and UO_1920 (O_1920,N_49910,N_49190);
nor UO_1921 (O_1921,N_49170,N_49968);
xnor UO_1922 (O_1922,N_49628,N_49266);
and UO_1923 (O_1923,N_49212,N_49447);
and UO_1924 (O_1924,N_49237,N_49326);
nand UO_1925 (O_1925,N_49103,N_49273);
and UO_1926 (O_1926,N_49579,N_49934);
nor UO_1927 (O_1927,N_49774,N_49683);
nand UO_1928 (O_1928,N_49560,N_49367);
nand UO_1929 (O_1929,N_49560,N_49407);
or UO_1930 (O_1930,N_49363,N_49285);
or UO_1931 (O_1931,N_49380,N_49193);
xor UO_1932 (O_1932,N_49698,N_49593);
nor UO_1933 (O_1933,N_49091,N_49468);
or UO_1934 (O_1934,N_49235,N_49595);
nor UO_1935 (O_1935,N_49315,N_49002);
xnor UO_1936 (O_1936,N_49640,N_49589);
nor UO_1937 (O_1937,N_49560,N_49607);
nor UO_1938 (O_1938,N_49390,N_49762);
nand UO_1939 (O_1939,N_49764,N_49322);
nor UO_1940 (O_1940,N_49850,N_49188);
xor UO_1941 (O_1941,N_49524,N_49476);
xor UO_1942 (O_1942,N_49056,N_49173);
nand UO_1943 (O_1943,N_49826,N_49483);
xor UO_1944 (O_1944,N_49108,N_49744);
nand UO_1945 (O_1945,N_49043,N_49587);
or UO_1946 (O_1946,N_49306,N_49773);
nand UO_1947 (O_1947,N_49756,N_49279);
xor UO_1948 (O_1948,N_49001,N_49831);
and UO_1949 (O_1949,N_49250,N_49376);
nor UO_1950 (O_1950,N_49441,N_49861);
and UO_1951 (O_1951,N_49487,N_49833);
and UO_1952 (O_1952,N_49501,N_49695);
nand UO_1953 (O_1953,N_49940,N_49808);
nand UO_1954 (O_1954,N_49508,N_49018);
nor UO_1955 (O_1955,N_49186,N_49908);
nand UO_1956 (O_1956,N_49146,N_49569);
xnor UO_1957 (O_1957,N_49476,N_49901);
nand UO_1958 (O_1958,N_49765,N_49956);
nand UO_1959 (O_1959,N_49607,N_49975);
nand UO_1960 (O_1960,N_49298,N_49408);
and UO_1961 (O_1961,N_49692,N_49018);
nand UO_1962 (O_1962,N_49913,N_49648);
nand UO_1963 (O_1963,N_49992,N_49201);
or UO_1964 (O_1964,N_49896,N_49740);
xnor UO_1965 (O_1965,N_49124,N_49099);
and UO_1966 (O_1966,N_49994,N_49065);
or UO_1967 (O_1967,N_49966,N_49457);
nor UO_1968 (O_1968,N_49129,N_49771);
or UO_1969 (O_1969,N_49514,N_49911);
nand UO_1970 (O_1970,N_49625,N_49459);
nor UO_1971 (O_1971,N_49347,N_49688);
xnor UO_1972 (O_1972,N_49037,N_49293);
nor UO_1973 (O_1973,N_49557,N_49821);
nand UO_1974 (O_1974,N_49649,N_49516);
nand UO_1975 (O_1975,N_49901,N_49308);
xor UO_1976 (O_1976,N_49008,N_49682);
and UO_1977 (O_1977,N_49935,N_49319);
nor UO_1978 (O_1978,N_49811,N_49963);
nor UO_1979 (O_1979,N_49897,N_49715);
xnor UO_1980 (O_1980,N_49308,N_49252);
nor UO_1981 (O_1981,N_49864,N_49192);
and UO_1982 (O_1982,N_49453,N_49833);
nor UO_1983 (O_1983,N_49609,N_49672);
and UO_1984 (O_1984,N_49825,N_49183);
or UO_1985 (O_1985,N_49468,N_49214);
and UO_1986 (O_1986,N_49606,N_49933);
xnor UO_1987 (O_1987,N_49425,N_49850);
nand UO_1988 (O_1988,N_49931,N_49177);
and UO_1989 (O_1989,N_49243,N_49788);
and UO_1990 (O_1990,N_49003,N_49282);
nand UO_1991 (O_1991,N_49106,N_49576);
or UO_1992 (O_1992,N_49622,N_49222);
xor UO_1993 (O_1993,N_49678,N_49424);
nor UO_1994 (O_1994,N_49144,N_49664);
or UO_1995 (O_1995,N_49024,N_49853);
nor UO_1996 (O_1996,N_49123,N_49063);
and UO_1997 (O_1997,N_49883,N_49917);
and UO_1998 (O_1998,N_49907,N_49287);
and UO_1999 (O_1999,N_49006,N_49966);
xnor UO_2000 (O_2000,N_49729,N_49172);
nor UO_2001 (O_2001,N_49136,N_49899);
or UO_2002 (O_2002,N_49973,N_49149);
or UO_2003 (O_2003,N_49474,N_49389);
nor UO_2004 (O_2004,N_49907,N_49881);
nand UO_2005 (O_2005,N_49374,N_49920);
or UO_2006 (O_2006,N_49057,N_49313);
and UO_2007 (O_2007,N_49498,N_49541);
nor UO_2008 (O_2008,N_49181,N_49192);
nand UO_2009 (O_2009,N_49863,N_49656);
and UO_2010 (O_2010,N_49078,N_49751);
or UO_2011 (O_2011,N_49109,N_49289);
and UO_2012 (O_2012,N_49869,N_49287);
xnor UO_2013 (O_2013,N_49134,N_49435);
xnor UO_2014 (O_2014,N_49018,N_49006);
or UO_2015 (O_2015,N_49781,N_49582);
nand UO_2016 (O_2016,N_49184,N_49753);
and UO_2017 (O_2017,N_49026,N_49803);
nand UO_2018 (O_2018,N_49581,N_49991);
or UO_2019 (O_2019,N_49364,N_49604);
nand UO_2020 (O_2020,N_49247,N_49763);
or UO_2021 (O_2021,N_49854,N_49968);
or UO_2022 (O_2022,N_49652,N_49607);
or UO_2023 (O_2023,N_49552,N_49108);
nor UO_2024 (O_2024,N_49780,N_49830);
nor UO_2025 (O_2025,N_49994,N_49987);
or UO_2026 (O_2026,N_49379,N_49787);
or UO_2027 (O_2027,N_49962,N_49978);
and UO_2028 (O_2028,N_49222,N_49037);
or UO_2029 (O_2029,N_49391,N_49748);
nor UO_2030 (O_2030,N_49836,N_49131);
xnor UO_2031 (O_2031,N_49177,N_49126);
xnor UO_2032 (O_2032,N_49087,N_49965);
nand UO_2033 (O_2033,N_49477,N_49195);
xnor UO_2034 (O_2034,N_49421,N_49604);
nand UO_2035 (O_2035,N_49432,N_49500);
or UO_2036 (O_2036,N_49390,N_49625);
or UO_2037 (O_2037,N_49636,N_49613);
nand UO_2038 (O_2038,N_49018,N_49867);
nor UO_2039 (O_2039,N_49217,N_49038);
xor UO_2040 (O_2040,N_49229,N_49459);
nand UO_2041 (O_2041,N_49780,N_49219);
xnor UO_2042 (O_2042,N_49742,N_49596);
xor UO_2043 (O_2043,N_49925,N_49386);
nor UO_2044 (O_2044,N_49041,N_49208);
xnor UO_2045 (O_2045,N_49465,N_49402);
nor UO_2046 (O_2046,N_49525,N_49297);
or UO_2047 (O_2047,N_49962,N_49043);
xor UO_2048 (O_2048,N_49817,N_49999);
xor UO_2049 (O_2049,N_49312,N_49243);
xnor UO_2050 (O_2050,N_49615,N_49092);
and UO_2051 (O_2051,N_49262,N_49202);
and UO_2052 (O_2052,N_49449,N_49555);
nand UO_2053 (O_2053,N_49573,N_49248);
or UO_2054 (O_2054,N_49356,N_49577);
xnor UO_2055 (O_2055,N_49322,N_49375);
nand UO_2056 (O_2056,N_49710,N_49177);
nand UO_2057 (O_2057,N_49674,N_49993);
xor UO_2058 (O_2058,N_49776,N_49241);
and UO_2059 (O_2059,N_49999,N_49161);
and UO_2060 (O_2060,N_49732,N_49565);
nand UO_2061 (O_2061,N_49814,N_49102);
nand UO_2062 (O_2062,N_49275,N_49947);
nor UO_2063 (O_2063,N_49726,N_49211);
xor UO_2064 (O_2064,N_49582,N_49785);
nand UO_2065 (O_2065,N_49998,N_49075);
nand UO_2066 (O_2066,N_49782,N_49950);
xor UO_2067 (O_2067,N_49749,N_49450);
or UO_2068 (O_2068,N_49087,N_49398);
or UO_2069 (O_2069,N_49912,N_49383);
or UO_2070 (O_2070,N_49426,N_49823);
nand UO_2071 (O_2071,N_49710,N_49864);
xnor UO_2072 (O_2072,N_49989,N_49762);
or UO_2073 (O_2073,N_49429,N_49265);
nor UO_2074 (O_2074,N_49271,N_49466);
nor UO_2075 (O_2075,N_49707,N_49139);
xor UO_2076 (O_2076,N_49134,N_49058);
xor UO_2077 (O_2077,N_49674,N_49161);
and UO_2078 (O_2078,N_49985,N_49632);
or UO_2079 (O_2079,N_49813,N_49916);
nand UO_2080 (O_2080,N_49810,N_49375);
or UO_2081 (O_2081,N_49212,N_49711);
xor UO_2082 (O_2082,N_49717,N_49823);
xor UO_2083 (O_2083,N_49526,N_49006);
nand UO_2084 (O_2084,N_49823,N_49783);
nor UO_2085 (O_2085,N_49907,N_49856);
xnor UO_2086 (O_2086,N_49593,N_49792);
nor UO_2087 (O_2087,N_49470,N_49126);
nor UO_2088 (O_2088,N_49383,N_49889);
xor UO_2089 (O_2089,N_49459,N_49664);
nor UO_2090 (O_2090,N_49307,N_49481);
or UO_2091 (O_2091,N_49764,N_49664);
nand UO_2092 (O_2092,N_49931,N_49672);
nand UO_2093 (O_2093,N_49964,N_49541);
and UO_2094 (O_2094,N_49420,N_49754);
nand UO_2095 (O_2095,N_49270,N_49586);
nand UO_2096 (O_2096,N_49055,N_49123);
nand UO_2097 (O_2097,N_49321,N_49167);
or UO_2098 (O_2098,N_49023,N_49669);
and UO_2099 (O_2099,N_49085,N_49486);
nand UO_2100 (O_2100,N_49592,N_49395);
nand UO_2101 (O_2101,N_49784,N_49913);
nor UO_2102 (O_2102,N_49902,N_49374);
nand UO_2103 (O_2103,N_49398,N_49509);
nor UO_2104 (O_2104,N_49293,N_49887);
nor UO_2105 (O_2105,N_49529,N_49921);
xor UO_2106 (O_2106,N_49284,N_49806);
xor UO_2107 (O_2107,N_49459,N_49470);
or UO_2108 (O_2108,N_49279,N_49162);
xor UO_2109 (O_2109,N_49123,N_49030);
and UO_2110 (O_2110,N_49978,N_49502);
and UO_2111 (O_2111,N_49452,N_49530);
xnor UO_2112 (O_2112,N_49623,N_49070);
and UO_2113 (O_2113,N_49431,N_49852);
xnor UO_2114 (O_2114,N_49894,N_49169);
xnor UO_2115 (O_2115,N_49604,N_49674);
xnor UO_2116 (O_2116,N_49145,N_49124);
xnor UO_2117 (O_2117,N_49536,N_49604);
or UO_2118 (O_2118,N_49865,N_49005);
or UO_2119 (O_2119,N_49433,N_49186);
and UO_2120 (O_2120,N_49490,N_49531);
xnor UO_2121 (O_2121,N_49080,N_49014);
xor UO_2122 (O_2122,N_49121,N_49336);
and UO_2123 (O_2123,N_49290,N_49178);
and UO_2124 (O_2124,N_49035,N_49393);
nand UO_2125 (O_2125,N_49030,N_49367);
and UO_2126 (O_2126,N_49253,N_49320);
nor UO_2127 (O_2127,N_49981,N_49698);
xnor UO_2128 (O_2128,N_49877,N_49432);
xor UO_2129 (O_2129,N_49825,N_49398);
or UO_2130 (O_2130,N_49196,N_49765);
nor UO_2131 (O_2131,N_49651,N_49294);
and UO_2132 (O_2132,N_49344,N_49000);
or UO_2133 (O_2133,N_49094,N_49221);
xor UO_2134 (O_2134,N_49985,N_49874);
nand UO_2135 (O_2135,N_49525,N_49568);
xnor UO_2136 (O_2136,N_49139,N_49401);
nand UO_2137 (O_2137,N_49758,N_49742);
xnor UO_2138 (O_2138,N_49318,N_49517);
or UO_2139 (O_2139,N_49857,N_49648);
or UO_2140 (O_2140,N_49846,N_49981);
nand UO_2141 (O_2141,N_49801,N_49298);
nand UO_2142 (O_2142,N_49178,N_49551);
nor UO_2143 (O_2143,N_49671,N_49328);
nor UO_2144 (O_2144,N_49897,N_49367);
nor UO_2145 (O_2145,N_49487,N_49387);
xnor UO_2146 (O_2146,N_49905,N_49386);
nand UO_2147 (O_2147,N_49735,N_49005);
and UO_2148 (O_2148,N_49027,N_49110);
and UO_2149 (O_2149,N_49551,N_49335);
nand UO_2150 (O_2150,N_49821,N_49762);
xnor UO_2151 (O_2151,N_49109,N_49901);
and UO_2152 (O_2152,N_49986,N_49498);
and UO_2153 (O_2153,N_49900,N_49208);
nand UO_2154 (O_2154,N_49186,N_49721);
xor UO_2155 (O_2155,N_49089,N_49930);
xor UO_2156 (O_2156,N_49822,N_49742);
and UO_2157 (O_2157,N_49904,N_49952);
nand UO_2158 (O_2158,N_49406,N_49160);
xnor UO_2159 (O_2159,N_49404,N_49848);
xor UO_2160 (O_2160,N_49019,N_49138);
nor UO_2161 (O_2161,N_49228,N_49449);
nor UO_2162 (O_2162,N_49940,N_49710);
nand UO_2163 (O_2163,N_49529,N_49329);
or UO_2164 (O_2164,N_49107,N_49340);
or UO_2165 (O_2165,N_49088,N_49878);
nor UO_2166 (O_2166,N_49892,N_49420);
or UO_2167 (O_2167,N_49418,N_49952);
or UO_2168 (O_2168,N_49109,N_49827);
and UO_2169 (O_2169,N_49420,N_49258);
or UO_2170 (O_2170,N_49767,N_49182);
xor UO_2171 (O_2171,N_49627,N_49271);
xor UO_2172 (O_2172,N_49746,N_49228);
nor UO_2173 (O_2173,N_49751,N_49205);
xor UO_2174 (O_2174,N_49356,N_49022);
nor UO_2175 (O_2175,N_49838,N_49468);
and UO_2176 (O_2176,N_49166,N_49495);
or UO_2177 (O_2177,N_49497,N_49387);
nand UO_2178 (O_2178,N_49562,N_49716);
and UO_2179 (O_2179,N_49632,N_49417);
or UO_2180 (O_2180,N_49930,N_49584);
nand UO_2181 (O_2181,N_49158,N_49690);
and UO_2182 (O_2182,N_49900,N_49571);
or UO_2183 (O_2183,N_49647,N_49063);
and UO_2184 (O_2184,N_49468,N_49792);
or UO_2185 (O_2185,N_49525,N_49564);
and UO_2186 (O_2186,N_49127,N_49973);
and UO_2187 (O_2187,N_49925,N_49257);
and UO_2188 (O_2188,N_49208,N_49206);
xnor UO_2189 (O_2189,N_49002,N_49538);
nor UO_2190 (O_2190,N_49731,N_49989);
or UO_2191 (O_2191,N_49250,N_49532);
and UO_2192 (O_2192,N_49311,N_49195);
xnor UO_2193 (O_2193,N_49048,N_49547);
nand UO_2194 (O_2194,N_49203,N_49659);
nor UO_2195 (O_2195,N_49400,N_49754);
nor UO_2196 (O_2196,N_49676,N_49726);
xor UO_2197 (O_2197,N_49145,N_49635);
nor UO_2198 (O_2198,N_49861,N_49005);
nor UO_2199 (O_2199,N_49467,N_49609);
and UO_2200 (O_2200,N_49122,N_49464);
or UO_2201 (O_2201,N_49495,N_49511);
or UO_2202 (O_2202,N_49551,N_49399);
and UO_2203 (O_2203,N_49905,N_49547);
nand UO_2204 (O_2204,N_49904,N_49225);
nand UO_2205 (O_2205,N_49756,N_49585);
and UO_2206 (O_2206,N_49075,N_49143);
xnor UO_2207 (O_2207,N_49693,N_49760);
xnor UO_2208 (O_2208,N_49285,N_49925);
xnor UO_2209 (O_2209,N_49691,N_49511);
and UO_2210 (O_2210,N_49647,N_49869);
or UO_2211 (O_2211,N_49596,N_49638);
or UO_2212 (O_2212,N_49395,N_49215);
and UO_2213 (O_2213,N_49427,N_49937);
and UO_2214 (O_2214,N_49555,N_49413);
or UO_2215 (O_2215,N_49827,N_49481);
xor UO_2216 (O_2216,N_49772,N_49022);
and UO_2217 (O_2217,N_49110,N_49370);
or UO_2218 (O_2218,N_49066,N_49696);
and UO_2219 (O_2219,N_49874,N_49138);
nor UO_2220 (O_2220,N_49080,N_49598);
nor UO_2221 (O_2221,N_49141,N_49267);
nor UO_2222 (O_2222,N_49729,N_49937);
and UO_2223 (O_2223,N_49500,N_49823);
nor UO_2224 (O_2224,N_49351,N_49474);
or UO_2225 (O_2225,N_49813,N_49772);
nand UO_2226 (O_2226,N_49454,N_49193);
xor UO_2227 (O_2227,N_49587,N_49798);
nand UO_2228 (O_2228,N_49605,N_49878);
xnor UO_2229 (O_2229,N_49335,N_49989);
nand UO_2230 (O_2230,N_49853,N_49465);
nand UO_2231 (O_2231,N_49138,N_49981);
or UO_2232 (O_2232,N_49672,N_49736);
xnor UO_2233 (O_2233,N_49523,N_49147);
or UO_2234 (O_2234,N_49788,N_49791);
or UO_2235 (O_2235,N_49911,N_49162);
xor UO_2236 (O_2236,N_49476,N_49355);
or UO_2237 (O_2237,N_49805,N_49506);
and UO_2238 (O_2238,N_49777,N_49279);
and UO_2239 (O_2239,N_49981,N_49343);
nand UO_2240 (O_2240,N_49568,N_49174);
xnor UO_2241 (O_2241,N_49119,N_49445);
nor UO_2242 (O_2242,N_49738,N_49840);
nand UO_2243 (O_2243,N_49877,N_49354);
xnor UO_2244 (O_2244,N_49683,N_49133);
nor UO_2245 (O_2245,N_49533,N_49053);
or UO_2246 (O_2246,N_49331,N_49913);
and UO_2247 (O_2247,N_49967,N_49466);
and UO_2248 (O_2248,N_49921,N_49857);
xor UO_2249 (O_2249,N_49879,N_49803);
xor UO_2250 (O_2250,N_49527,N_49554);
or UO_2251 (O_2251,N_49440,N_49837);
nand UO_2252 (O_2252,N_49212,N_49703);
xnor UO_2253 (O_2253,N_49582,N_49048);
nand UO_2254 (O_2254,N_49868,N_49910);
and UO_2255 (O_2255,N_49038,N_49741);
xnor UO_2256 (O_2256,N_49528,N_49347);
or UO_2257 (O_2257,N_49815,N_49759);
or UO_2258 (O_2258,N_49156,N_49799);
nand UO_2259 (O_2259,N_49129,N_49097);
or UO_2260 (O_2260,N_49149,N_49831);
xor UO_2261 (O_2261,N_49189,N_49826);
xnor UO_2262 (O_2262,N_49235,N_49331);
nand UO_2263 (O_2263,N_49523,N_49545);
nor UO_2264 (O_2264,N_49659,N_49210);
xnor UO_2265 (O_2265,N_49696,N_49257);
and UO_2266 (O_2266,N_49398,N_49158);
nor UO_2267 (O_2267,N_49031,N_49461);
and UO_2268 (O_2268,N_49466,N_49410);
nor UO_2269 (O_2269,N_49141,N_49238);
xnor UO_2270 (O_2270,N_49230,N_49579);
nand UO_2271 (O_2271,N_49174,N_49250);
nor UO_2272 (O_2272,N_49726,N_49132);
or UO_2273 (O_2273,N_49590,N_49215);
and UO_2274 (O_2274,N_49830,N_49078);
and UO_2275 (O_2275,N_49425,N_49846);
xnor UO_2276 (O_2276,N_49388,N_49179);
and UO_2277 (O_2277,N_49537,N_49396);
nor UO_2278 (O_2278,N_49569,N_49480);
or UO_2279 (O_2279,N_49889,N_49197);
nand UO_2280 (O_2280,N_49756,N_49807);
or UO_2281 (O_2281,N_49242,N_49354);
and UO_2282 (O_2282,N_49386,N_49442);
xor UO_2283 (O_2283,N_49507,N_49709);
and UO_2284 (O_2284,N_49046,N_49257);
xnor UO_2285 (O_2285,N_49961,N_49722);
nor UO_2286 (O_2286,N_49635,N_49829);
nor UO_2287 (O_2287,N_49818,N_49256);
nand UO_2288 (O_2288,N_49359,N_49425);
nor UO_2289 (O_2289,N_49006,N_49007);
or UO_2290 (O_2290,N_49892,N_49771);
and UO_2291 (O_2291,N_49012,N_49542);
and UO_2292 (O_2292,N_49868,N_49257);
xor UO_2293 (O_2293,N_49232,N_49894);
nand UO_2294 (O_2294,N_49201,N_49786);
nor UO_2295 (O_2295,N_49459,N_49839);
nor UO_2296 (O_2296,N_49224,N_49340);
and UO_2297 (O_2297,N_49381,N_49213);
xor UO_2298 (O_2298,N_49040,N_49515);
or UO_2299 (O_2299,N_49542,N_49255);
and UO_2300 (O_2300,N_49865,N_49039);
nand UO_2301 (O_2301,N_49066,N_49753);
and UO_2302 (O_2302,N_49691,N_49842);
xnor UO_2303 (O_2303,N_49192,N_49034);
nor UO_2304 (O_2304,N_49350,N_49394);
nor UO_2305 (O_2305,N_49683,N_49996);
nand UO_2306 (O_2306,N_49793,N_49945);
and UO_2307 (O_2307,N_49387,N_49227);
nand UO_2308 (O_2308,N_49365,N_49443);
nor UO_2309 (O_2309,N_49773,N_49408);
nor UO_2310 (O_2310,N_49408,N_49951);
or UO_2311 (O_2311,N_49046,N_49623);
and UO_2312 (O_2312,N_49566,N_49509);
or UO_2313 (O_2313,N_49522,N_49204);
or UO_2314 (O_2314,N_49051,N_49032);
or UO_2315 (O_2315,N_49305,N_49749);
or UO_2316 (O_2316,N_49848,N_49407);
or UO_2317 (O_2317,N_49230,N_49247);
nor UO_2318 (O_2318,N_49579,N_49734);
nor UO_2319 (O_2319,N_49831,N_49570);
xor UO_2320 (O_2320,N_49524,N_49647);
or UO_2321 (O_2321,N_49596,N_49200);
nand UO_2322 (O_2322,N_49310,N_49926);
nand UO_2323 (O_2323,N_49472,N_49341);
nor UO_2324 (O_2324,N_49772,N_49426);
or UO_2325 (O_2325,N_49856,N_49060);
xor UO_2326 (O_2326,N_49622,N_49655);
and UO_2327 (O_2327,N_49528,N_49572);
nand UO_2328 (O_2328,N_49170,N_49447);
nand UO_2329 (O_2329,N_49371,N_49693);
nor UO_2330 (O_2330,N_49025,N_49474);
nor UO_2331 (O_2331,N_49469,N_49016);
and UO_2332 (O_2332,N_49860,N_49987);
and UO_2333 (O_2333,N_49179,N_49548);
nor UO_2334 (O_2334,N_49752,N_49497);
nand UO_2335 (O_2335,N_49066,N_49774);
and UO_2336 (O_2336,N_49427,N_49357);
and UO_2337 (O_2337,N_49292,N_49922);
and UO_2338 (O_2338,N_49225,N_49183);
nand UO_2339 (O_2339,N_49342,N_49972);
and UO_2340 (O_2340,N_49480,N_49952);
and UO_2341 (O_2341,N_49950,N_49147);
xnor UO_2342 (O_2342,N_49644,N_49612);
nand UO_2343 (O_2343,N_49293,N_49435);
nand UO_2344 (O_2344,N_49404,N_49422);
xor UO_2345 (O_2345,N_49540,N_49923);
nor UO_2346 (O_2346,N_49847,N_49684);
and UO_2347 (O_2347,N_49580,N_49826);
nor UO_2348 (O_2348,N_49769,N_49477);
nor UO_2349 (O_2349,N_49242,N_49576);
and UO_2350 (O_2350,N_49682,N_49095);
nor UO_2351 (O_2351,N_49077,N_49826);
and UO_2352 (O_2352,N_49678,N_49305);
and UO_2353 (O_2353,N_49256,N_49548);
nor UO_2354 (O_2354,N_49587,N_49061);
xnor UO_2355 (O_2355,N_49368,N_49698);
xnor UO_2356 (O_2356,N_49863,N_49725);
xor UO_2357 (O_2357,N_49331,N_49883);
xnor UO_2358 (O_2358,N_49039,N_49668);
xnor UO_2359 (O_2359,N_49660,N_49951);
or UO_2360 (O_2360,N_49257,N_49071);
or UO_2361 (O_2361,N_49682,N_49502);
or UO_2362 (O_2362,N_49395,N_49722);
nand UO_2363 (O_2363,N_49087,N_49994);
xor UO_2364 (O_2364,N_49107,N_49467);
or UO_2365 (O_2365,N_49916,N_49275);
and UO_2366 (O_2366,N_49493,N_49636);
and UO_2367 (O_2367,N_49393,N_49325);
and UO_2368 (O_2368,N_49658,N_49328);
nor UO_2369 (O_2369,N_49854,N_49120);
nor UO_2370 (O_2370,N_49944,N_49867);
nand UO_2371 (O_2371,N_49984,N_49101);
nand UO_2372 (O_2372,N_49699,N_49868);
nand UO_2373 (O_2373,N_49355,N_49388);
nor UO_2374 (O_2374,N_49142,N_49629);
or UO_2375 (O_2375,N_49720,N_49781);
xor UO_2376 (O_2376,N_49742,N_49006);
nor UO_2377 (O_2377,N_49513,N_49019);
or UO_2378 (O_2378,N_49715,N_49991);
or UO_2379 (O_2379,N_49425,N_49119);
xor UO_2380 (O_2380,N_49133,N_49012);
or UO_2381 (O_2381,N_49265,N_49435);
nor UO_2382 (O_2382,N_49122,N_49428);
and UO_2383 (O_2383,N_49507,N_49575);
and UO_2384 (O_2384,N_49058,N_49679);
and UO_2385 (O_2385,N_49606,N_49730);
xor UO_2386 (O_2386,N_49961,N_49531);
or UO_2387 (O_2387,N_49090,N_49372);
or UO_2388 (O_2388,N_49299,N_49658);
xor UO_2389 (O_2389,N_49754,N_49295);
and UO_2390 (O_2390,N_49419,N_49580);
xnor UO_2391 (O_2391,N_49312,N_49695);
nor UO_2392 (O_2392,N_49050,N_49996);
xor UO_2393 (O_2393,N_49533,N_49770);
xor UO_2394 (O_2394,N_49745,N_49333);
and UO_2395 (O_2395,N_49048,N_49965);
nor UO_2396 (O_2396,N_49309,N_49427);
xnor UO_2397 (O_2397,N_49150,N_49277);
nor UO_2398 (O_2398,N_49980,N_49818);
and UO_2399 (O_2399,N_49756,N_49509);
nand UO_2400 (O_2400,N_49912,N_49805);
nand UO_2401 (O_2401,N_49254,N_49448);
or UO_2402 (O_2402,N_49565,N_49143);
xor UO_2403 (O_2403,N_49194,N_49630);
or UO_2404 (O_2404,N_49032,N_49466);
nor UO_2405 (O_2405,N_49765,N_49134);
nor UO_2406 (O_2406,N_49966,N_49745);
nand UO_2407 (O_2407,N_49761,N_49583);
xor UO_2408 (O_2408,N_49602,N_49477);
xor UO_2409 (O_2409,N_49814,N_49191);
nor UO_2410 (O_2410,N_49898,N_49483);
and UO_2411 (O_2411,N_49514,N_49869);
nand UO_2412 (O_2412,N_49092,N_49641);
xnor UO_2413 (O_2413,N_49345,N_49183);
or UO_2414 (O_2414,N_49014,N_49681);
nor UO_2415 (O_2415,N_49960,N_49241);
xor UO_2416 (O_2416,N_49304,N_49784);
nor UO_2417 (O_2417,N_49787,N_49252);
or UO_2418 (O_2418,N_49539,N_49681);
or UO_2419 (O_2419,N_49665,N_49995);
xor UO_2420 (O_2420,N_49311,N_49359);
xor UO_2421 (O_2421,N_49327,N_49141);
or UO_2422 (O_2422,N_49627,N_49630);
and UO_2423 (O_2423,N_49032,N_49409);
and UO_2424 (O_2424,N_49602,N_49456);
nor UO_2425 (O_2425,N_49820,N_49357);
nor UO_2426 (O_2426,N_49935,N_49249);
nor UO_2427 (O_2427,N_49295,N_49566);
nor UO_2428 (O_2428,N_49186,N_49871);
nand UO_2429 (O_2429,N_49156,N_49378);
nor UO_2430 (O_2430,N_49202,N_49379);
or UO_2431 (O_2431,N_49519,N_49913);
xor UO_2432 (O_2432,N_49109,N_49158);
and UO_2433 (O_2433,N_49808,N_49244);
nand UO_2434 (O_2434,N_49881,N_49821);
nor UO_2435 (O_2435,N_49556,N_49030);
and UO_2436 (O_2436,N_49235,N_49832);
nor UO_2437 (O_2437,N_49993,N_49003);
and UO_2438 (O_2438,N_49138,N_49898);
and UO_2439 (O_2439,N_49652,N_49165);
nor UO_2440 (O_2440,N_49577,N_49748);
nor UO_2441 (O_2441,N_49939,N_49418);
or UO_2442 (O_2442,N_49774,N_49737);
or UO_2443 (O_2443,N_49375,N_49057);
nand UO_2444 (O_2444,N_49566,N_49626);
xor UO_2445 (O_2445,N_49800,N_49214);
xor UO_2446 (O_2446,N_49416,N_49698);
or UO_2447 (O_2447,N_49272,N_49432);
or UO_2448 (O_2448,N_49331,N_49568);
nor UO_2449 (O_2449,N_49234,N_49765);
and UO_2450 (O_2450,N_49125,N_49217);
and UO_2451 (O_2451,N_49782,N_49308);
nor UO_2452 (O_2452,N_49166,N_49685);
nor UO_2453 (O_2453,N_49064,N_49707);
nand UO_2454 (O_2454,N_49630,N_49033);
nand UO_2455 (O_2455,N_49718,N_49901);
xor UO_2456 (O_2456,N_49010,N_49618);
or UO_2457 (O_2457,N_49058,N_49931);
nand UO_2458 (O_2458,N_49934,N_49044);
and UO_2459 (O_2459,N_49256,N_49037);
nand UO_2460 (O_2460,N_49349,N_49747);
xor UO_2461 (O_2461,N_49038,N_49385);
nand UO_2462 (O_2462,N_49126,N_49180);
and UO_2463 (O_2463,N_49918,N_49047);
nor UO_2464 (O_2464,N_49298,N_49089);
nor UO_2465 (O_2465,N_49850,N_49180);
nor UO_2466 (O_2466,N_49633,N_49557);
xnor UO_2467 (O_2467,N_49178,N_49904);
nor UO_2468 (O_2468,N_49517,N_49431);
xnor UO_2469 (O_2469,N_49007,N_49472);
nand UO_2470 (O_2470,N_49540,N_49680);
nor UO_2471 (O_2471,N_49772,N_49028);
nor UO_2472 (O_2472,N_49440,N_49259);
nor UO_2473 (O_2473,N_49788,N_49371);
and UO_2474 (O_2474,N_49652,N_49601);
xnor UO_2475 (O_2475,N_49945,N_49475);
xnor UO_2476 (O_2476,N_49193,N_49190);
nor UO_2477 (O_2477,N_49712,N_49226);
xor UO_2478 (O_2478,N_49326,N_49346);
xnor UO_2479 (O_2479,N_49520,N_49962);
nor UO_2480 (O_2480,N_49000,N_49734);
or UO_2481 (O_2481,N_49726,N_49704);
nand UO_2482 (O_2482,N_49480,N_49497);
and UO_2483 (O_2483,N_49648,N_49403);
nor UO_2484 (O_2484,N_49040,N_49050);
and UO_2485 (O_2485,N_49946,N_49918);
nand UO_2486 (O_2486,N_49517,N_49025);
xor UO_2487 (O_2487,N_49464,N_49650);
or UO_2488 (O_2488,N_49152,N_49550);
and UO_2489 (O_2489,N_49316,N_49306);
nor UO_2490 (O_2490,N_49726,N_49789);
nor UO_2491 (O_2491,N_49112,N_49499);
and UO_2492 (O_2492,N_49544,N_49067);
nor UO_2493 (O_2493,N_49059,N_49573);
nor UO_2494 (O_2494,N_49494,N_49550);
xor UO_2495 (O_2495,N_49568,N_49391);
nor UO_2496 (O_2496,N_49125,N_49820);
and UO_2497 (O_2497,N_49950,N_49046);
nand UO_2498 (O_2498,N_49300,N_49268);
nor UO_2499 (O_2499,N_49141,N_49833);
and UO_2500 (O_2500,N_49669,N_49867);
nor UO_2501 (O_2501,N_49438,N_49184);
nor UO_2502 (O_2502,N_49553,N_49999);
xor UO_2503 (O_2503,N_49561,N_49657);
xnor UO_2504 (O_2504,N_49462,N_49959);
xor UO_2505 (O_2505,N_49638,N_49342);
and UO_2506 (O_2506,N_49882,N_49130);
nand UO_2507 (O_2507,N_49233,N_49639);
and UO_2508 (O_2508,N_49794,N_49189);
and UO_2509 (O_2509,N_49119,N_49663);
and UO_2510 (O_2510,N_49587,N_49542);
nand UO_2511 (O_2511,N_49548,N_49282);
or UO_2512 (O_2512,N_49728,N_49833);
nor UO_2513 (O_2513,N_49984,N_49975);
or UO_2514 (O_2514,N_49749,N_49998);
nor UO_2515 (O_2515,N_49322,N_49351);
or UO_2516 (O_2516,N_49176,N_49848);
or UO_2517 (O_2517,N_49548,N_49911);
and UO_2518 (O_2518,N_49569,N_49965);
and UO_2519 (O_2519,N_49892,N_49665);
nor UO_2520 (O_2520,N_49912,N_49362);
nor UO_2521 (O_2521,N_49896,N_49677);
nand UO_2522 (O_2522,N_49554,N_49323);
or UO_2523 (O_2523,N_49542,N_49300);
xnor UO_2524 (O_2524,N_49542,N_49761);
or UO_2525 (O_2525,N_49134,N_49700);
and UO_2526 (O_2526,N_49655,N_49171);
xnor UO_2527 (O_2527,N_49624,N_49657);
or UO_2528 (O_2528,N_49994,N_49826);
xnor UO_2529 (O_2529,N_49466,N_49419);
or UO_2530 (O_2530,N_49861,N_49844);
xnor UO_2531 (O_2531,N_49616,N_49457);
or UO_2532 (O_2532,N_49702,N_49378);
and UO_2533 (O_2533,N_49015,N_49558);
nand UO_2534 (O_2534,N_49640,N_49387);
xnor UO_2535 (O_2535,N_49460,N_49275);
nor UO_2536 (O_2536,N_49777,N_49522);
nor UO_2537 (O_2537,N_49645,N_49380);
xnor UO_2538 (O_2538,N_49227,N_49528);
xnor UO_2539 (O_2539,N_49426,N_49526);
nor UO_2540 (O_2540,N_49910,N_49155);
and UO_2541 (O_2541,N_49280,N_49603);
nor UO_2542 (O_2542,N_49610,N_49130);
and UO_2543 (O_2543,N_49026,N_49129);
or UO_2544 (O_2544,N_49390,N_49978);
or UO_2545 (O_2545,N_49216,N_49362);
nand UO_2546 (O_2546,N_49653,N_49344);
and UO_2547 (O_2547,N_49775,N_49357);
xor UO_2548 (O_2548,N_49222,N_49477);
nor UO_2549 (O_2549,N_49133,N_49316);
nand UO_2550 (O_2550,N_49115,N_49282);
or UO_2551 (O_2551,N_49925,N_49087);
or UO_2552 (O_2552,N_49244,N_49018);
nand UO_2553 (O_2553,N_49377,N_49481);
nand UO_2554 (O_2554,N_49923,N_49644);
and UO_2555 (O_2555,N_49360,N_49504);
nand UO_2556 (O_2556,N_49498,N_49106);
nand UO_2557 (O_2557,N_49494,N_49132);
nor UO_2558 (O_2558,N_49206,N_49655);
and UO_2559 (O_2559,N_49445,N_49672);
nand UO_2560 (O_2560,N_49831,N_49356);
xor UO_2561 (O_2561,N_49228,N_49068);
and UO_2562 (O_2562,N_49758,N_49302);
or UO_2563 (O_2563,N_49340,N_49204);
nand UO_2564 (O_2564,N_49636,N_49533);
xnor UO_2565 (O_2565,N_49466,N_49238);
and UO_2566 (O_2566,N_49249,N_49120);
nor UO_2567 (O_2567,N_49782,N_49177);
xor UO_2568 (O_2568,N_49268,N_49944);
and UO_2569 (O_2569,N_49651,N_49678);
nand UO_2570 (O_2570,N_49168,N_49799);
xor UO_2571 (O_2571,N_49385,N_49826);
nand UO_2572 (O_2572,N_49421,N_49186);
and UO_2573 (O_2573,N_49484,N_49744);
nand UO_2574 (O_2574,N_49366,N_49608);
or UO_2575 (O_2575,N_49301,N_49614);
or UO_2576 (O_2576,N_49342,N_49899);
or UO_2577 (O_2577,N_49741,N_49637);
nand UO_2578 (O_2578,N_49571,N_49307);
xor UO_2579 (O_2579,N_49449,N_49129);
nor UO_2580 (O_2580,N_49048,N_49823);
and UO_2581 (O_2581,N_49927,N_49349);
nor UO_2582 (O_2582,N_49780,N_49727);
nand UO_2583 (O_2583,N_49667,N_49651);
nand UO_2584 (O_2584,N_49948,N_49972);
nand UO_2585 (O_2585,N_49288,N_49783);
nand UO_2586 (O_2586,N_49523,N_49895);
or UO_2587 (O_2587,N_49015,N_49426);
nor UO_2588 (O_2588,N_49690,N_49798);
nand UO_2589 (O_2589,N_49489,N_49843);
or UO_2590 (O_2590,N_49003,N_49322);
nor UO_2591 (O_2591,N_49628,N_49927);
nor UO_2592 (O_2592,N_49128,N_49979);
nand UO_2593 (O_2593,N_49406,N_49004);
xnor UO_2594 (O_2594,N_49166,N_49940);
nand UO_2595 (O_2595,N_49329,N_49551);
xor UO_2596 (O_2596,N_49302,N_49442);
nand UO_2597 (O_2597,N_49605,N_49813);
nand UO_2598 (O_2598,N_49488,N_49943);
or UO_2599 (O_2599,N_49977,N_49591);
nor UO_2600 (O_2600,N_49988,N_49825);
and UO_2601 (O_2601,N_49279,N_49471);
nand UO_2602 (O_2602,N_49119,N_49300);
and UO_2603 (O_2603,N_49583,N_49939);
or UO_2604 (O_2604,N_49916,N_49282);
and UO_2605 (O_2605,N_49074,N_49935);
xnor UO_2606 (O_2606,N_49899,N_49626);
nor UO_2607 (O_2607,N_49226,N_49688);
nor UO_2608 (O_2608,N_49045,N_49297);
and UO_2609 (O_2609,N_49669,N_49099);
nor UO_2610 (O_2610,N_49043,N_49404);
or UO_2611 (O_2611,N_49908,N_49592);
nand UO_2612 (O_2612,N_49359,N_49062);
and UO_2613 (O_2613,N_49735,N_49854);
xnor UO_2614 (O_2614,N_49711,N_49048);
nor UO_2615 (O_2615,N_49688,N_49477);
nand UO_2616 (O_2616,N_49744,N_49306);
nand UO_2617 (O_2617,N_49637,N_49189);
nor UO_2618 (O_2618,N_49118,N_49936);
or UO_2619 (O_2619,N_49130,N_49836);
nor UO_2620 (O_2620,N_49985,N_49971);
or UO_2621 (O_2621,N_49670,N_49736);
and UO_2622 (O_2622,N_49441,N_49739);
nand UO_2623 (O_2623,N_49640,N_49284);
xor UO_2624 (O_2624,N_49546,N_49915);
nor UO_2625 (O_2625,N_49648,N_49153);
or UO_2626 (O_2626,N_49004,N_49009);
nor UO_2627 (O_2627,N_49003,N_49563);
or UO_2628 (O_2628,N_49979,N_49225);
and UO_2629 (O_2629,N_49345,N_49533);
nor UO_2630 (O_2630,N_49337,N_49710);
or UO_2631 (O_2631,N_49312,N_49988);
nor UO_2632 (O_2632,N_49445,N_49463);
xor UO_2633 (O_2633,N_49537,N_49756);
nor UO_2634 (O_2634,N_49322,N_49512);
xor UO_2635 (O_2635,N_49528,N_49802);
nand UO_2636 (O_2636,N_49984,N_49120);
xnor UO_2637 (O_2637,N_49799,N_49574);
xor UO_2638 (O_2638,N_49053,N_49139);
xor UO_2639 (O_2639,N_49450,N_49061);
xnor UO_2640 (O_2640,N_49760,N_49742);
and UO_2641 (O_2641,N_49361,N_49111);
or UO_2642 (O_2642,N_49837,N_49847);
xor UO_2643 (O_2643,N_49391,N_49938);
nand UO_2644 (O_2644,N_49522,N_49833);
nand UO_2645 (O_2645,N_49510,N_49344);
nor UO_2646 (O_2646,N_49758,N_49975);
and UO_2647 (O_2647,N_49004,N_49992);
or UO_2648 (O_2648,N_49024,N_49845);
nor UO_2649 (O_2649,N_49825,N_49842);
xor UO_2650 (O_2650,N_49207,N_49563);
nor UO_2651 (O_2651,N_49770,N_49708);
xor UO_2652 (O_2652,N_49959,N_49397);
nand UO_2653 (O_2653,N_49918,N_49577);
nand UO_2654 (O_2654,N_49493,N_49390);
and UO_2655 (O_2655,N_49637,N_49015);
or UO_2656 (O_2656,N_49080,N_49868);
nor UO_2657 (O_2657,N_49810,N_49698);
and UO_2658 (O_2658,N_49176,N_49244);
xor UO_2659 (O_2659,N_49524,N_49307);
nand UO_2660 (O_2660,N_49888,N_49867);
nor UO_2661 (O_2661,N_49076,N_49268);
xnor UO_2662 (O_2662,N_49004,N_49868);
nor UO_2663 (O_2663,N_49260,N_49090);
xor UO_2664 (O_2664,N_49440,N_49694);
or UO_2665 (O_2665,N_49412,N_49825);
xnor UO_2666 (O_2666,N_49709,N_49011);
nand UO_2667 (O_2667,N_49774,N_49427);
nor UO_2668 (O_2668,N_49574,N_49589);
nor UO_2669 (O_2669,N_49986,N_49782);
nand UO_2670 (O_2670,N_49152,N_49297);
or UO_2671 (O_2671,N_49310,N_49364);
nor UO_2672 (O_2672,N_49805,N_49363);
or UO_2673 (O_2673,N_49555,N_49210);
nor UO_2674 (O_2674,N_49040,N_49995);
nand UO_2675 (O_2675,N_49418,N_49395);
nand UO_2676 (O_2676,N_49840,N_49328);
xor UO_2677 (O_2677,N_49142,N_49508);
xor UO_2678 (O_2678,N_49500,N_49672);
nand UO_2679 (O_2679,N_49704,N_49657);
or UO_2680 (O_2680,N_49189,N_49198);
nor UO_2681 (O_2681,N_49562,N_49182);
xnor UO_2682 (O_2682,N_49842,N_49175);
nand UO_2683 (O_2683,N_49094,N_49143);
or UO_2684 (O_2684,N_49812,N_49506);
or UO_2685 (O_2685,N_49897,N_49661);
nor UO_2686 (O_2686,N_49781,N_49499);
and UO_2687 (O_2687,N_49056,N_49862);
nor UO_2688 (O_2688,N_49276,N_49314);
or UO_2689 (O_2689,N_49759,N_49392);
nand UO_2690 (O_2690,N_49983,N_49501);
nor UO_2691 (O_2691,N_49898,N_49781);
nand UO_2692 (O_2692,N_49716,N_49622);
xor UO_2693 (O_2693,N_49477,N_49298);
or UO_2694 (O_2694,N_49524,N_49489);
and UO_2695 (O_2695,N_49265,N_49977);
xnor UO_2696 (O_2696,N_49245,N_49418);
and UO_2697 (O_2697,N_49687,N_49008);
nor UO_2698 (O_2698,N_49684,N_49366);
nor UO_2699 (O_2699,N_49483,N_49085);
nand UO_2700 (O_2700,N_49077,N_49928);
nor UO_2701 (O_2701,N_49173,N_49651);
xnor UO_2702 (O_2702,N_49960,N_49254);
nor UO_2703 (O_2703,N_49116,N_49741);
or UO_2704 (O_2704,N_49927,N_49669);
nand UO_2705 (O_2705,N_49979,N_49482);
and UO_2706 (O_2706,N_49165,N_49293);
and UO_2707 (O_2707,N_49563,N_49976);
or UO_2708 (O_2708,N_49216,N_49261);
or UO_2709 (O_2709,N_49551,N_49954);
xor UO_2710 (O_2710,N_49082,N_49011);
nor UO_2711 (O_2711,N_49799,N_49349);
nand UO_2712 (O_2712,N_49951,N_49539);
xnor UO_2713 (O_2713,N_49271,N_49837);
nor UO_2714 (O_2714,N_49740,N_49807);
nand UO_2715 (O_2715,N_49720,N_49681);
nor UO_2716 (O_2716,N_49876,N_49290);
nand UO_2717 (O_2717,N_49771,N_49733);
and UO_2718 (O_2718,N_49351,N_49427);
nand UO_2719 (O_2719,N_49373,N_49862);
xnor UO_2720 (O_2720,N_49695,N_49137);
xor UO_2721 (O_2721,N_49101,N_49295);
xor UO_2722 (O_2722,N_49048,N_49081);
xor UO_2723 (O_2723,N_49172,N_49067);
nor UO_2724 (O_2724,N_49936,N_49607);
or UO_2725 (O_2725,N_49381,N_49651);
xnor UO_2726 (O_2726,N_49939,N_49547);
or UO_2727 (O_2727,N_49514,N_49579);
and UO_2728 (O_2728,N_49288,N_49482);
nor UO_2729 (O_2729,N_49595,N_49989);
xor UO_2730 (O_2730,N_49190,N_49715);
nand UO_2731 (O_2731,N_49204,N_49220);
nor UO_2732 (O_2732,N_49596,N_49139);
or UO_2733 (O_2733,N_49395,N_49306);
xor UO_2734 (O_2734,N_49715,N_49113);
or UO_2735 (O_2735,N_49671,N_49303);
xor UO_2736 (O_2736,N_49643,N_49001);
xor UO_2737 (O_2737,N_49988,N_49346);
nand UO_2738 (O_2738,N_49472,N_49790);
nand UO_2739 (O_2739,N_49349,N_49078);
nand UO_2740 (O_2740,N_49035,N_49619);
and UO_2741 (O_2741,N_49993,N_49375);
xnor UO_2742 (O_2742,N_49676,N_49402);
nor UO_2743 (O_2743,N_49329,N_49188);
nor UO_2744 (O_2744,N_49658,N_49399);
nand UO_2745 (O_2745,N_49682,N_49047);
nand UO_2746 (O_2746,N_49399,N_49225);
nor UO_2747 (O_2747,N_49740,N_49084);
or UO_2748 (O_2748,N_49531,N_49897);
or UO_2749 (O_2749,N_49935,N_49117);
nand UO_2750 (O_2750,N_49324,N_49712);
xnor UO_2751 (O_2751,N_49226,N_49128);
and UO_2752 (O_2752,N_49800,N_49458);
and UO_2753 (O_2753,N_49002,N_49332);
xnor UO_2754 (O_2754,N_49421,N_49770);
xnor UO_2755 (O_2755,N_49786,N_49117);
nor UO_2756 (O_2756,N_49689,N_49781);
nand UO_2757 (O_2757,N_49469,N_49874);
or UO_2758 (O_2758,N_49224,N_49307);
nor UO_2759 (O_2759,N_49151,N_49571);
and UO_2760 (O_2760,N_49988,N_49642);
nor UO_2761 (O_2761,N_49909,N_49207);
nand UO_2762 (O_2762,N_49167,N_49824);
xnor UO_2763 (O_2763,N_49268,N_49869);
and UO_2764 (O_2764,N_49507,N_49975);
nand UO_2765 (O_2765,N_49417,N_49192);
or UO_2766 (O_2766,N_49051,N_49031);
nand UO_2767 (O_2767,N_49410,N_49267);
xnor UO_2768 (O_2768,N_49587,N_49298);
or UO_2769 (O_2769,N_49545,N_49209);
and UO_2770 (O_2770,N_49935,N_49569);
nor UO_2771 (O_2771,N_49950,N_49902);
nand UO_2772 (O_2772,N_49812,N_49632);
and UO_2773 (O_2773,N_49035,N_49550);
or UO_2774 (O_2774,N_49928,N_49006);
and UO_2775 (O_2775,N_49560,N_49271);
nand UO_2776 (O_2776,N_49689,N_49279);
nor UO_2777 (O_2777,N_49969,N_49806);
nand UO_2778 (O_2778,N_49161,N_49304);
nand UO_2779 (O_2779,N_49758,N_49069);
nand UO_2780 (O_2780,N_49826,N_49702);
xnor UO_2781 (O_2781,N_49821,N_49148);
or UO_2782 (O_2782,N_49092,N_49674);
xnor UO_2783 (O_2783,N_49157,N_49469);
nor UO_2784 (O_2784,N_49110,N_49944);
xnor UO_2785 (O_2785,N_49106,N_49905);
nor UO_2786 (O_2786,N_49863,N_49937);
xor UO_2787 (O_2787,N_49172,N_49179);
and UO_2788 (O_2788,N_49336,N_49213);
nor UO_2789 (O_2789,N_49770,N_49439);
nand UO_2790 (O_2790,N_49022,N_49630);
xor UO_2791 (O_2791,N_49444,N_49614);
nand UO_2792 (O_2792,N_49606,N_49271);
nand UO_2793 (O_2793,N_49035,N_49839);
xor UO_2794 (O_2794,N_49747,N_49578);
or UO_2795 (O_2795,N_49802,N_49405);
nand UO_2796 (O_2796,N_49972,N_49280);
nand UO_2797 (O_2797,N_49374,N_49452);
nor UO_2798 (O_2798,N_49772,N_49742);
and UO_2799 (O_2799,N_49130,N_49571);
nand UO_2800 (O_2800,N_49979,N_49916);
xor UO_2801 (O_2801,N_49672,N_49213);
nor UO_2802 (O_2802,N_49261,N_49361);
or UO_2803 (O_2803,N_49381,N_49565);
nand UO_2804 (O_2804,N_49782,N_49789);
and UO_2805 (O_2805,N_49751,N_49428);
xnor UO_2806 (O_2806,N_49908,N_49473);
or UO_2807 (O_2807,N_49434,N_49392);
or UO_2808 (O_2808,N_49096,N_49778);
nand UO_2809 (O_2809,N_49980,N_49733);
nor UO_2810 (O_2810,N_49333,N_49290);
nor UO_2811 (O_2811,N_49878,N_49594);
or UO_2812 (O_2812,N_49854,N_49927);
nand UO_2813 (O_2813,N_49051,N_49528);
and UO_2814 (O_2814,N_49677,N_49553);
nor UO_2815 (O_2815,N_49504,N_49932);
xor UO_2816 (O_2816,N_49152,N_49492);
and UO_2817 (O_2817,N_49117,N_49460);
nor UO_2818 (O_2818,N_49847,N_49289);
and UO_2819 (O_2819,N_49308,N_49331);
nor UO_2820 (O_2820,N_49750,N_49409);
nor UO_2821 (O_2821,N_49897,N_49828);
or UO_2822 (O_2822,N_49329,N_49456);
nor UO_2823 (O_2823,N_49267,N_49034);
and UO_2824 (O_2824,N_49786,N_49199);
nor UO_2825 (O_2825,N_49272,N_49237);
nor UO_2826 (O_2826,N_49714,N_49469);
nand UO_2827 (O_2827,N_49834,N_49664);
xor UO_2828 (O_2828,N_49673,N_49370);
or UO_2829 (O_2829,N_49166,N_49458);
nor UO_2830 (O_2830,N_49711,N_49097);
or UO_2831 (O_2831,N_49817,N_49536);
or UO_2832 (O_2832,N_49666,N_49204);
and UO_2833 (O_2833,N_49773,N_49080);
nor UO_2834 (O_2834,N_49393,N_49517);
nand UO_2835 (O_2835,N_49926,N_49613);
nor UO_2836 (O_2836,N_49731,N_49472);
xnor UO_2837 (O_2837,N_49549,N_49151);
nand UO_2838 (O_2838,N_49233,N_49457);
nand UO_2839 (O_2839,N_49278,N_49764);
nand UO_2840 (O_2840,N_49730,N_49325);
or UO_2841 (O_2841,N_49883,N_49628);
xnor UO_2842 (O_2842,N_49816,N_49562);
or UO_2843 (O_2843,N_49125,N_49042);
nand UO_2844 (O_2844,N_49609,N_49860);
xnor UO_2845 (O_2845,N_49917,N_49322);
xor UO_2846 (O_2846,N_49393,N_49353);
nand UO_2847 (O_2847,N_49824,N_49801);
xnor UO_2848 (O_2848,N_49961,N_49156);
nand UO_2849 (O_2849,N_49725,N_49288);
nand UO_2850 (O_2850,N_49597,N_49565);
and UO_2851 (O_2851,N_49259,N_49254);
nor UO_2852 (O_2852,N_49602,N_49199);
xnor UO_2853 (O_2853,N_49108,N_49587);
xor UO_2854 (O_2854,N_49784,N_49802);
xnor UO_2855 (O_2855,N_49419,N_49120);
nor UO_2856 (O_2856,N_49165,N_49478);
nand UO_2857 (O_2857,N_49716,N_49324);
or UO_2858 (O_2858,N_49670,N_49367);
xor UO_2859 (O_2859,N_49896,N_49420);
nor UO_2860 (O_2860,N_49708,N_49781);
xor UO_2861 (O_2861,N_49413,N_49619);
xor UO_2862 (O_2862,N_49156,N_49405);
and UO_2863 (O_2863,N_49273,N_49347);
or UO_2864 (O_2864,N_49408,N_49816);
and UO_2865 (O_2865,N_49688,N_49023);
nand UO_2866 (O_2866,N_49768,N_49593);
and UO_2867 (O_2867,N_49065,N_49956);
nand UO_2868 (O_2868,N_49137,N_49383);
nand UO_2869 (O_2869,N_49176,N_49557);
and UO_2870 (O_2870,N_49856,N_49467);
xor UO_2871 (O_2871,N_49257,N_49975);
or UO_2872 (O_2872,N_49465,N_49665);
or UO_2873 (O_2873,N_49213,N_49344);
xor UO_2874 (O_2874,N_49532,N_49215);
xnor UO_2875 (O_2875,N_49050,N_49364);
or UO_2876 (O_2876,N_49639,N_49421);
or UO_2877 (O_2877,N_49673,N_49229);
nand UO_2878 (O_2878,N_49241,N_49161);
nand UO_2879 (O_2879,N_49159,N_49370);
or UO_2880 (O_2880,N_49201,N_49116);
xnor UO_2881 (O_2881,N_49191,N_49749);
nand UO_2882 (O_2882,N_49749,N_49912);
nand UO_2883 (O_2883,N_49417,N_49516);
and UO_2884 (O_2884,N_49760,N_49246);
and UO_2885 (O_2885,N_49678,N_49963);
nor UO_2886 (O_2886,N_49192,N_49152);
nor UO_2887 (O_2887,N_49403,N_49201);
and UO_2888 (O_2888,N_49109,N_49366);
nand UO_2889 (O_2889,N_49718,N_49881);
or UO_2890 (O_2890,N_49367,N_49527);
nor UO_2891 (O_2891,N_49641,N_49965);
nor UO_2892 (O_2892,N_49767,N_49667);
nor UO_2893 (O_2893,N_49898,N_49044);
or UO_2894 (O_2894,N_49060,N_49034);
or UO_2895 (O_2895,N_49066,N_49644);
or UO_2896 (O_2896,N_49102,N_49095);
nor UO_2897 (O_2897,N_49901,N_49224);
xor UO_2898 (O_2898,N_49865,N_49410);
nand UO_2899 (O_2899,N_49144,N_49768);
and UO_2900 (O_2900,N_49211,N_49645);
nor UO_2901 (O_2901,N_49429,N_49426);
nor UO_2902 (O_2902,N_49947,N_49583);
xnor UO_2903 (O_2903,N_49849,N_49907);
xnor UO_2904 (O_2904,N_49410,N_49699);
nand UO_2905 (O_2905,N_49918,N_49253);
xor UO_2906 (O_2906,N_49560,N_49582);
or UO_2907 (O_2907,N_49932,N_49878);
and UO_2908 (O_2908,N_49526,N_49179);
or UO_2909 (O_2909,N_49998,N_49434);
and UO_2910 (O_2910,N_49599,N_49687);
nor UO_2911 (O_2911,N_49666,N_49813);
nand UO_2912 (O_2912,N_49993,N_49864);
or UO_2913 (O_2913,N_49862,N_49988);
nor UO_2914 (O_2914,N_49431,N_49370);
nand UO_2915 (O_2915,N_49859,N_49983);
nor UO_2916 (O_2916,N_49902,N_49207);
and UO_2917 (O_2917,N_49059,N_49096);
and UO_2918 (O_2918,N_49143,N_49877);
and UO_2919 (O_2919,N_49129,N_49756);
nor UO_2920 (O_2920,N_49348,N_49337);
or UO_2921 (O_2921,N_49416,N_49168);
nand UO_2922 (O_2922,N_49412,N_49127);
nand UO_2923 (O_2923,N_49462,N_49647);
xnor UO_2924 (O_2924,N_49023,N_49768);
xor UO_2925 (O_2925,N_49398,N_49898);
nand UO_2926 (O_2926,N_49672,N_49888);
and UO_2927 (O_2927,N_49395,N_49756);
xor UO_2928 (O_2928,N_49070,N_49696);
nor UO_2929 (O_2929,N_49775,N_49220);
or UO_2930 (O_2930,N_49876,N_49726);
nand UO_2931 (O_2931,N_49019,N_49933);
or UO_2932 (O_2932,N_49698,N_49332);
nor UO_2933 (O_2933,N_49681,N_49877);
or UO_2934 (O_2934,N_49820,N_49520);
and UO_2935 (O_2935,N_49347,N_49342);
nor UO_2936 (O_2936,N_49872,N_49555);
nand UO_2937 (O_2937,N_49297,N_49781);
or UO_2938 (O_2938,N_49492,N_49018);
or UO_2939 (O_2939,N_49587,N_49057);
and UO_2940 (O_2940,N_49452,N_49092);
nand UO_2941 (O_2941,N_49758,N_49079);
nand UO_2942 (O_2942,N_49884,N_49465);
or UO_2943 (O_2943,N_49318,N_49754);
and UO_2944 (O_2944,N_49599,N_49367);
nor UO_2945 (O_2945,N_49016,N_49570);
nor UO_2946 (O_2946,N_49403,N_49954);
and UO_2947 (O_2947,N_49837,N_49380);
xor UO_2948 (O_2948,N_49723,N_49047);
nor UO_2949 (O_2949,N_49328,N_49237);
xor UO_2950 (O_2950,N_49110,N_49940);
nor UO_2951 (O_2951,N_49112,N_49037);
and UO_2952 (O_2952,N_49997,N_49005);
nor UO_2953 (O_2953,N_49947,N_49499);
nor UO_2954 (O_2954,N_49799,N_49919);
nand UO_2955 (O_2955,N_49117,N_49703);
nor UO_2956 (O_2956,N_49935,N_49067);
and UO_2957 (O_2957,N_49404,N_49481);
or UO_2958 (O_2958,N_49047,N_49870);
and UO_2959 (O_2959,N_49809,N_49749);
nand UO_2960 (O_2960,N_49082,N_49184);
nor UO_2961 (O_2961,N_49076,N_49634);
xnor UO_2962 (O_2962,N_49830,N_49855);
nor UO_2963 (O_2963,N_49990,N_49650);
and UO_2964 (O_2964,N_49169,N_49162);
and UO_2965 (O_2965,N_49254,N_49513);
nor UO_2966 (O_2966,N_49881,N_49833);
and UO_2967 (O_2967,N_49569,N_49061);
nand UO_2968 (O_2968,N_49699,N_49878);
nand UO_2969 (O_2969,N_49370,N_49426);
and UO_2970 (O_2970,N_49653,N_49476);
and UO_2971 (O_2971,N_49377,N_49398);
nor UO_2972 (O_2972,N_49348,N_49927);
and UO_2973 (O_2973,N_49490,N_49236);
nor UO_2974 (O_2974,N_49177,N_49868);
nor UO_2975 (O_2975,N_49408,N_49213);
xor UO_2976 (O_2976,N_49821,N_49382);
xnor UO_2977 (O_2977,N_49383,N_49537);
nor UO_2978 (O_2978,N_49336,N_49841);
and UO_2979 (O_2979,N_49620,N_49455);
and UO_2980 (O_2980,N_49400,N_49933);
nand UO_2981 (O_2981,N_49783,N_49120);
or UO_2982 (O_2982,N_49859,N_49322);
nor UO_2983 (O_2983,N_49281,N_49537);
or UO_2984 (O_2984,N_49154,N_49716);
nand UO_2985 (O_2985,N_49637,N_49810);
nand UO_2986 (O_2986,N_49847,N_49012);
xor UO_2987 (O_2987,N_49813,N_49032);
xor UO_2988 (O_2988,N_49849,N_49514);
and UO_2989 (O_2989,N_49420,N_49795);
xnor UO_2990 (O_2990,N_49658,N_49983);
and UO_2991 (O_2991,N_49414,N_49422);
nor UO_2992 (O_2992,N_49759,N_49925);
xnor UO_2993 (O_2993,N_49829,N_49446);
and UO_2994 (O_2994,N_49053,N_49477);
xor UO_2995 (O_2995,N_49878,N_49161);
nor UO_2996 (O_2996,N_49026,N_49458);
xnor UO_2997 (O_2997,N_49909,N_49872);
or UO_2998 (O_2998,N_49114,N_49628);
and UO_2999 (O_2999,N_49093,N_49322);
and UO_3000 (O_3000,N_49486,N_49476);
nand UO_3001 (O_3001,N_49242,N_49631);
nor UO_3002 (O_3002,N_49433,N_49272);
and UO_3003 (O_3003,N_49776,N_49363);
nand UO_3004 (O_3004,N_49787,N_49080);
nor UO_3005 (O_3005,N_49428,N_49203);
or UO_3006 (O_3006,N_49007,N_49422);
and UO_3007 (O_3007,N_49668,N_49576);
and UO_3008 (O_3008,N_49251,N_49171);
or UO_3009 (O_3009,N_49357,N_49634);
or UO_3010 (O_3010,N_49818,N_49646);
nand UO_3011 (O_3011,N_49712,N_49012);
and UO_3012 (O_3012,N_49615,N_49471);
nand UO_3013 (O_3013,N_49799,N_49662);
and UO_3014 (O_3014,N_49058,N_49834);
and UO_3015 (O_3015,N_49961,N_49579);
or UO_3016 (O_3016,N_49109,N_49421);
nand UO_3017 (O_3017,N_49424,N_49928);
nand UO_3018 (O_3018,N_49128,N_49119);
nand UO_3019 (O_3019,N_49069,N_49371);
nor UO_3020 (O_3020,N_49316,N_49803);
xnor UO_3021 (O_3021,N_49024,N_49589);
and UO_3022 (O_3022,N_49266,N_49233);
xnor UO_3023 (O_3023,N_49766,N_49943);
xor UO_3024 (O_3024,N_49300,N_49391);
nand UO_3025 (O_3025,N_49386,N_49158);
nand UO_3026 (O_3026,N_49458,N_49763);
nand UO_3027 (O_3027,N_49199,N_49856);
nor UO_3028 (O_3028,N_49966,N_49170);
nand UO_3029 (O_3029,N_49756,N_49933);
xnor UO_3030 (O_3030,N_49795,N_49287);
or UO_3031 (O_3031,N_49445,N_49787);
xor UO_3032 (O_3032,N_49183,N_49241);
and UO_3033 (O_3033,N_49055,N_49109);
nor UO_3034 (O_3034,N_49902,N_49942);
xnor UO_3035 (O_3035,N_49668,N_49316);
nand UO_3036 (O_3036,N_49311,N_49765);
and UO_3037 (O_3037,N_49018,N_49343);
or UO_3038 (O_3038,N_49914,N_49172);
nor UO_3039 (O_3039,N_49823,N_49409);
xor UO_3040 (O_3040,N_49843,N_49384);
and UO_3041 (O_3041,N_49744,N_49831);
nor UO_3042 (O_3042,N_49320,N_49887);
and UO_3043 (O_3043,N_49225,N_49993);
and UO_3044 (O_3044,N_49349,N_49547);
xor UO_3045 (O_3045,N_49646,N_49337);
xor UO_3046 (O_3046,N_49868,N_49046);
nor UO_3047 (O_3047,N_49147,N_49477);
or UO_3048 (O_3048,N_49055,N_49314);
nand UO_3049 (O_3049,N_49694,N_49999);
nand UO_3050 (O_3050,N_49252,N_49754);
and UO_3051 (O_3051,N_49651,N_49746);
or UO_3052 (O_3052,N_49946,N_49559);
xnor UO_3053 (O_3053,N_49291,N_49880);
and UO_3054 (O_3054,N_49662,N_49835);
or UO_3055 (O_3055,N_49028,N_49900);
xor UO_3056 (O_3056,N_49938,N_49504);
or UO_3057 (O_3057,N_49222,N_49302);
nand UO_3058 (O_3058,N_49044,N_49915);
or UO_3059 (O_3059,N_49762,N_49784);
xnor UO_3060 (O_3060,N_49381,N_49613);
nand UO_3061 (O_3061,N_49740,N_49701);
xnor UO_3062 (O_3062,N_49453,N_49831);
or UO_3063 (O_3063,N_49375,N_49814);
nor UO_3064 (O_3064,N_49566,N_49573);
or UO_3065 (O_3065,N_49539,N_49271);
or UO_3066 (O_3066,N_49500,N_49089);
nand UO_3067 (O_3067,N_49495,N_49788);
and UO_3068 (O_3068,N_49908,N_49507);
xor UO_3069 (O_3069,N_49512,N_49897);
or UO_3070 (O_3070,N_49220,N_49673);
nand UO_3071 (O_3071,N_49084,N_49501);
and UO_3072 (O_3072,N_49243,N_49138);
and UO_3073 (O_3073,N_49890,N_49716);
nor UO_3074 (O_3074,N_49820,N_49492);
nand UO_3075 (O_3075,N_49120,N_49541);
xor UO_3076 (O_3076,N_49106,N_49799);
and UO_3077 (O_3077,N_49956,N_49411);
nor UO_3078 (O_3078,N_49486,N_49815);
and UO_3079 (O_3079,N_49727,N_49073);
nor UO_3080 (O_3080,N_49976,N_49395);
and UO_3081 (O_3081,N_49992,N_49577);
and UO_3082 (O_3082,N_49419,N_49047);
or UO_3083 (O_3083,N_49762,N_49369);
xor UO_3084 (O_3084,N_49087,N_49034);
or UO_3085 (O_3085,N_49740,N_49195);
xnor UO_3086 (O_3086,N_49879,N_49258);
or UO_3087 (O_3087,N_49773,N_49506);
or UO_3088 (O_3088,N_49322,N_49951);
nand UO_3089 (O_3089,N_49581,N_49853);
xor UO_3090 (O_3090,N_49870,N_49082);
xor UO_3091 (O_3091,N_49880,N_49787);
xnor UO_3092 (O_3092,N_49806,N_49516);
or UO_3093 (O_3093,N_49561,N_49907);
or UO_3094 (O_3094,N_49036,N_49791);
xor UO_3095 (O_3095,N_49906,N_49570);
or UO_3096 (O_3096,N_49112,N_49135);
and UO_3097 (O_3097,N_49733,N_49010);
xor UO_3098 (O_3098,N_49311,N_49982);
or UO_3099 (O_3099,N_49377,N_49490);
or UO_3100 (O_3100,N_49661,N_49250);
xor UO_3101 (O_3101,N_49996,N_49711);
nor UO_3102 (O_3102,N_49842,N_49770);
and UO_3103 (O_3103,N_49416,N_49993);
xor UO_3104 (O_3104,N_49703,N_49767);
and UO_3105 (O_3105,N_49153,N_49549);
and UO_3106 (O_3106,N_49922,N_49350);
nand UO_3107 (O_3107,N_49425,N_49636);
and UO_3108 (O_3108,N_49848,N_49741);
nor UO_3109 (O_3109,N_49512,N_49820);
and UO_3110 (O_3110,N_49833,N_49114);
nor UO_3111 (O_3111,N_49565,N_49795);
nand UO_3112 (O_3112,N_49085,N_49444);
xor UO_3113 (O_3113,N_49943,N_49773);
nor UO_3114 (O_3114,N_49977,N_49383);
xor UO_3115 (O_3115,N_49862,N_49163);
nor UO_3116 (O_3116,N_49470,N_49555);
nor UO_3117 (O_3117,N_49165,N_49959);
and UO_3118 (O_3118,N_49577,N_49523);
xor UO_3119 (O_3119,N_49154,N_49322);
xnor UO_3120 (O_3120,N_49929,N_49795);
nand UO_3121 (O_3121,N_49186,N_49002);
or UO_3122 (O_3122,N_49341,N_49357);
and UO_3123 (O_3123,N_49374,N_49461);
xor UO_3124 (O_3124,N_49143,N_49035);
nor UO_3125 (O_3125,N_49825,N_49307);
or UO_3126 (O_3126,N_49194,N_49953);
nor UO_3127 (O_3127,N_49771,N_49102);
nor UO_3128 (O_3128,N_49141,N_49882);
and UO_3129 (O_3129,N_49693,N_49375);
nand UO_3130 (O_3130,N_49018,N_49072);
nand UO_3131 (O_3131,N_49292,N_49729);
nor UO_3132 (O_3132,N_49971,N_49430);
and UO_3133 (O_3133,N_49490,N_49605);
or UO_3134 (O_3134,N_49486,N_49997);
and UO_3135 (O_3135,N_49073,N_49138);
nand UO_3136 (O_3136,N_49419,N_49508);
or UO_3137 (O_3137,N_49768,N_49109);
nor UO_3138 (O_3138,N_49559,N_49270);
or UO_3139 (O_3139,N_49507,N_49124);
nand UO_3140 (O_3140,N_49552,N_49165);
nor UO_3141 (O_3141,N_49908,N_49290);
nor UO_3142 (O_3142,N_49891,N_49973);
or UO_3143 (O_3143,N_49329,N_49544);
or UO_3144 (O_3144,N_49726,N_49005);
or UO_3145 (O_3145,N_49452,N_49422);
nand UO_3146 (O_3146,N_49753,N_49514);
nand UO_3147 (O_3147,N_49048,N_49659);
nand UO_3148 (O_3148,N_49993,N_49753);
nor UO_3149 (O_3149,N_49223,N_49393);
xor UO_3150 (O_3150,N_49446,N_49543);
or UO_3151 (O_3151,N_49857,N_49670);
or UO_3152 (O_3152,N_49604,N_49047);
xor UO_3153 (O_3153,N_49824,N_49732);
nand UO_3154 (O_3154,N_49839,N_49045);
or UO_3155 (O_3155,N_49526,N_49749);
and UO_3156 (O_3156,N_49173,N_49263);
and UO_3157 (O_3157,N_49219,N_49809);
nand UO_3158 (O_3158,N_49156,N_49779);
nor UO_3159 (O_3159,N_49414,N_49814);
xor UO_3160 (O_3160,N_49076,N_49691);
or UO_3161 (O_3161,N_49897,N_49179);
nor UO_3162 (O_3162,N_49564,N_49324);
and UO_3163 (O_3163,N_49954,N_49845);
nor UO_3164 (O_3164,N_49820,N_49579);
nand UO_3165 (O_3165,N_49416,N_49219);
and UO_3166 (O_3166,N_49506,N_49412);
nor UO_3167 (O_3167,N_49395,N_49461);
xor UO_3168 (O_3168,N_49474,N_49769);
or UO_3169 (O_3169,N_49551,N_49590);
and UO_3170 (O_3170,N_49536,N_49974);
or UO_3171 (O_3171,N_49113,N_49280);
or UO_3172 (O_3172,N_49570,N_49352);
xor UO_3173 (O_3173,N_49946,N_49728);
xor UO_3174 (O_3174,N_49182,N_49652);
xnor UO_3175 (O_3175,N_49038,N_49873);
and UO_3176 (O_3176,N_49422,N_49804);
nor UO_3177 (O_3177,N_49730,N_49904);
nor UO_3178 (O_3178,N_49221,N_49292);
or UO_3179 (O_3179,N_49912,N_49343);
and UO_3180 (O_3180,N_49709,N_49413);
or UO_3181 (O_3181,N_49721,N_49532);
nor UO_3182 (O_3182,N_49397,N_49513);
xnor UO_3183 (O_3183,N_49044,N_49704);
and UO_3184 (O_3184,N_49614,N_49536);
xor UO_3185 (O_3185,N_49307,N_49270);
or UO_3186 (O_3186,N_49855,N_49109);
and UO_3187 (O_3187,N_49182,N_49078);
or UO_3188 (O_3188,N_49038,N_49737);
xnor UO_3189 (O_3189,N_49344,N_49169);
nand UO_3190 (O_3190,N_49536,N_49637);
nand UO_3191 (O_3191,N_49256,N_49602);
or UO_3192 (O_3192,N_49891,N_49445);
or UO_3193 (O_3193,N_49509,N_49740);
nand UO_3194 (O_3194,N_49945,N_49422);
nor UO_3195 (O_3195,N_49467,N_49477);
or UO_3196 (O_3196,N_49637,N_49520);
xnor UO_3197 (O_3197,N_49004,N_49909);
nor UO_3198 (O_3198,N_49413,N_49040);
and UO_3199 (O_3199,N_49676,N_49530);
or UO_3200 (O_3200,N_49925,N_49519);
and UO_3201 (O_3201,N_49462,N_49563);
and UO_3202 (O_3202,N_49329,N_49309);
or UO_3203 (O_3203,N_49861,N_49956);
nand UO_3204 (O_3204,N_49091,N_49267);
nand UO_3205 (O_3205,N_49650,N_49524);
nand UO_3206 (O_3206,N_49743,N_49827);
xor UO_3207 (O_3207,N_49318,N_49032);
nand UO_3208 (O_3208,N_49950,N_49199);
xor UO_3209 (O_3209,N_49066,N_49001);
or UO_3210 (O_3210,N_49592,N_49494);
xnor UO_3211 (O_3211,N_49490,N_49466);
nor UO_3212 (O_3212,N_49127,N_49803);
nand UO_3213 (O_3213,N_49784,N_49937);
nor UO_3214 (O_3214,N_49694,N_49341);
xor UO_3215 (O_3215,N_49523,N_49848);
xnor UO_3216 (O_3216,N_49228,N_49640);
xor UO_3217 (O_3217,N_49378,N_49122);
nor UO_3218 (O_3218,N_49596,N_49680);
xnor UO_3219 (O_3219,N_49986,N_49883);
xor UO_3220 (O_3220,N_49055,N_49579);
or UO_3221 (O_3221,N_49326,N_49279);
nor UO_3222 (O_3222,N_49078,N_49403);
xor UO_3223 (O_3223,N_49788,N_49817);
nor UO_3224 (O_3224,N_49553,N_49719);
xnor UO_3225 (O_3225,N_49335,N_49115);
or UO_3226 (O_3226,N_49338,N_49159);
and UO_3227 (O_3227,N_49019,N_49839);
xnor UO_3228 (O_3228,N_49596,N_49410);
nand UO_3229 (O_3229,N_49515,N_49178);
nand UO_3230 (O_3230,N_49229,N_49829);
xnor UO_3231 (O_3231,N_49646,N_49066);
nor UO_3232 (O_3232,N_49902,N_49569);
nor UO_3233 (O_3233,N_49392,N_49750);
or UO_3234 (O_3234,N_49662,N_49506);
nor UO_3235 (O_3235,N_49033,N_49894);
nor UO_3236 (O_3236,N_49408,N_49171);
or UO_3237 (O_3237,N_49749,N_49800);
nor UO_3238 (O_3238,N_49911,N_49617);
and UO_3239 (O_3239,N_49186,N_49169);
nand UO_3240 (O_3240,N_49395,N_49331);
xnor UO_3241 (O_3241,N_49885,N_49453);
and UO_3242 (O_3242,N_49360,N_49724);
or UO_3243 (O_3243,N_49692,N_49599);
or UO_3244 (O_3244,N_49064,N_49880);
or UO_3245 (O_3245,N_49102,N_49258);
xor UO_3246 (O_3246,N_49629,N_49852);
and UO_3247 (O_3247,N_49239,N_49602);
nand UO_3248 (O_3248,N_49713,N_49595);
nor UO_3249 (O_3249,N_49059,N_49662);
nor UO_3250 (O_3250,N_49570,N_49914);
nand UO_3251 (O_3251,N_49503,N_49545);
and UO_3252 (O_3252,N_49195,N_49471);
and UO_3253 (O_3253,N_49579,N_49095);
and UO_3254 (O_3254,N_49424,N_49420);
nand UO_3255 (O_3255,N_49967,N_49688);
nor UO_3256 (O_3256,N_49514,N_49327);
nand UO_3257 (O_3257,N_49689,N_49932);
xnor UO_3258 (O_3258,N_49679,N_49353);
nand UO_3259 (O_3259,N_49010,N_49011);
and UO_3260 (O_3260,N_49716,N_49942);
nor UO_3261 (O_3261,N_49206,N_49891);
or UO_3262 (O_3262,N_49931,N_49924);
nand UO_3263 (O_3263,N_49102,N_49526);
or UO_3264 (O_3264,N_49956,N_49682);
nand UO_3265 (O_3265,N_49318,N_49941);
xnor UO_3266 (O_3266,N_49423,N_49261);
or UO_3267 (O_3267,N_49094,N_49474);
and UO_3268 (O_3268,N_49505,N_49720);
and UO_3269 (O_3269,N_49808,N_49828);
nand UO_3270 (O_3270,N_49402,N_49947);
xor UO_3271 (O_3271,N_49510,N_49102);
or UO_3272 (O_3272,N_49215,N_49292);
xor UO_3273 (O_3273,N_49147,N_49232);
and UO_3274 (O_3274,N_49449,N_49522);
nor UO_3275 (O_3275,N_49009,N_49903);
nor UO_3276 (O_3276,N_49163,N_49779);
nand UO_3277 (O_3277,N_49181,N_49022);
or UO_3278 (O_3278,N_49218,N_49016);
xnor UO_3279 (O_3279,N_49006,N_49498);
xor UO_3280 (O_3280,N_49020,N_49443);
nor UO_3281 (O_3281,N_49887,N_49075);
xor UO_3282 (O_3282,N_49266,N_49351);
nor UO_3283 (O_3283,N_49579,N_49902);
xnor UO_3284 (O_3284,N_49944,N_49938);
and UO_3285 (O_3285,N_49216,N_49283);
xor UO_3286 (O_3286,N_49121,N_49464);
xor UO_3287 (O_3287,N_49838,N_49365);
nand UO_3288 (O_3288,N_49497,N_49737);
xnor UO_3289 (O_3289,N_49404,N_49583);
and UO_3290 (O_3290,N_49047,N_49329);
and UO_3291 (O_3291,N_49313,N_49167);
or UO_3292 (O_3292,N_49357,N_49735);
and UO_3293 (O_3293,N_49644,N_49860);
xor UO_3294 (O_3294,N_49049,N_49145);
xor UO_3295 (O_3295,N_49782,N_49761);
and UO_3296 (O_3296,N_49670,N_49003);
nand UO_3297 (O_3297,N_49369,N_49953);
nor UO_3298 (O_3298,N_49864,N_49609);
nor UO_3299 (O_3299,N_49883,N_49826);
and UO_3300 (O_3300,N_49464,N_49481);
and UO_3301 (O_3301,N_49320,N_49563);
and UO_3302 (O_3302,N_49337,N_49062);
xnor UO_3303 (O_3303,N_49182,N_49423);
or UO_3304 (O_3304,N_49035,N_49145);
xnor UO_3305 (O_3305,N_49083,N_49265);
xnor UO_3306 (O_3306,N_49205,N_49780);
and UO_3307 (O_3307,N_49457,N_49458);
or UO_3308 (O_3308,N_49095,N_49905);
xnor UO_3309 (O_3309,N_49263,N_49519);
and UO_3310 (O_3310,N_49388,N_49683);
nand UO_3311 (O_3311,N_49447,N_49227);
nor UO_3312 (O_3312,N_49663,N_49906);
or UO_3313 (O_3313,N_49881,N_49470);
xor UO_3314 (O_3314,N_49064,N_49534);
and UO_3315 (O_3315,N_49017,N_49798);
or UO_3316 (O_3316,N_49280,N_49397);
nand UO_3317 (O_3317,N_49055,N_49666);
and UO_3318 (O_3318,N_49413,N_49541);
or UO_3319 (O_3319,N_49597,N_49485);
nor UO_3320 (O_3320,N_49937,N_49340);
nand UO_3321 (O_3321,N_49421,N_49592);
and UO_3322 (O_3322,N_49215,N_49325);
and UO_3323 (O_3323,N_49814,N_49895);
xor UO_3324 (O_3324,N_49690,N_49062);
nor UO_3325 (O_3325,N_49386,N_49983);
and UO_3326 (O_3326,N_49494,N_49620);
xnor UO_3327 (O_3327,N_49932,N_49229);
xnor UO_3328 (O_3328,N_49285,N_49805);
nand UO_3329 (O_3329,N_49932,N_49370);
nor UO_3330 (O_3330,N_49988,N_49015);
and UO_3331 (O_3331,N_49244,N_49578);
and UO_3332 (O_3332,N_49126,N_49010);
xnor UO_3333 (O_3333,N_49172,N_49431);
or UO_3334 (O_3334,N_49588,N_49585);
nor UO_3335 (O_3335,N_49002,N_49375);
nand UO_3336 (O_3336,N_49039,N_49792);
or UO_3337 (O_3337,N_49660,N_49538);
nand UO_3338 (O_3338,N_49487,N_49299);
nand UO_3339 (O_3339,N_49503,N_49355);
nand UO_3340 (O_3340,N_49552,N_49154);
xor UO_3341 (O_3341,N_49324,N_49782);
nand UO_3342 (O_3342,N_49391,N_49926);
and UO_3343 (O_3343,N_49440,N_49589);
nand UO_3344 (O_3344,N_49992,N_49411);
and UO_3345 (O_3345,N_49646,N_49817);
and UO_3346 (O_3346,N_49885,N_49361);
nand UO_3347 (O_3347,N_49202,N_49059);
or UO_3348 (O_3348,N_49992,N_49099);
or UO_3349 (O_3349,N_49076,N_49257);
and UO_3350 (O_3350,N_49653,N_49432);
or UO_3351 (O_3351,N_49777,N_49076);
xnor UO_3352 (O_3352,N_49014,N_49669);
xnor UO_3353 (O_3353,N_49063,N_49221);
xor UO_3354 (O_3354,N_49952,N_49764);
nand UO_3355 (O_3355,N_49366,N_49607);
nand UO_3356 (O_3356,N_49824,N_49050);
and UO_3357 (O_3357,N_49981,N_49074);
and UO_3358 (O_3358,N_49979,N_49993);
nand UO_3359 (O_3359,N_49209,N_49836);
and UO_3360 (O_3360,N_49022,N_49174);
and UO_3361 (O_3361,N_49241,N_49333);
or UO_3362 (O_3362,N_49303,N_49757);
xor UO_3363 (O_3363,N_49465,N_49337);
or UO_3364 (O_3364,N_49080,N_49392);
nor UO_3365 (O_3365,N_49372,N_49606);
nand UO_3366 (O_3366,N_49989,N_49099);
nand UO_3367 (O_3367,N_49888,N_49600);
nor UO_3368 (O_3368,N_49813,N_49315);
nand UO_3369 (O_3369,N_49518,N_49178);
xor UO_3370 (O_3370,N_49333,N_49793);
or UO_3371 (O_3371,N_49564,N_49274);
nand UO_3372 (O_3372,N_49861,N_49428);
xnor UO_3373 (O_3373,N_49041,N_49561);
nor UO_3374 (O_3374,N_49523,N_49442);
or UO_3375 (O_3375,N_49836,N_49503);
and UO_3376 (O_3376,N_49565,N_49038);
xor UO_3377 (O_3377,N_49768,N_49335);
nor UO_3378 (O_3378,N_49145,N_49936);
nand UO_3379 (O_3379,N_49641,N_49604);
and UO_3380 (O_3380,N_49733,N_49291);
nand UO_3381 (O_3381,N_49058,N_49458);
xnor UO_3382 (O_3382,N_49131,N_49632);
nand UO_3383 (O_3383,N_49966,N_49622);
nor UO_3384 (O_3384,N_49719,N_49537);
xor UO_3385 (O_3385,N_49297,N_49257);
or UO_3386 (O_3386,N_49849,N_49290);
and UO_3387 (O_3387,N_49966,N_49986);
nand UO_3388 (O_3388,N_49162,N_49235);
and UO_3389 (O_3389,N_49706,N_49927);
nor UO_3390 (O_3390,N_49578,N_49798);
nand UO_3391 (O_3391,N_49771,N_49413);
and UO_3392 (O_3392,N_49968,N_49241);
or UO_3393 (O_3393,N_49950,N_49929);
nor UO_3394 (O_3394,N_49588,N_49778);
xor UO_3395 (O_3395,N_49895,N_49936);
nor UO_3396 (O_3396,N_49545,N_49362);
or UO_3397 (O_3397,N_49375,N_49995);
or UO_3398 (O_3398,N_49934,N_49468);
and UO_3399 (O_3399,N_49811,N_49570);
nand UO_3400 (O_3400,N_49125,N_49080);
nor UO_3401 (O_3401,N_49230,N_49014);
and UO_3402 (O_3402,N_49785,N_49356);
nor UO_3403 (O_3403,N_49461,N_49637);
or UO_3404 (O_3404,N_49669,N_49070);
nor UO_3405 (O_3405,N_49120,N_49169);
nor UO_3406 (O_3406,N_49636,N_49804);
and UO_3407 (O_3407,N_49429,N_49738);
or UO_3408 (O_3408,N_49011,N_49352);
nor UO_3409 (O_3409,N_49170,N_49504);
nor UO_3410 (O_3410,N_49973,N_49770);
and UO_3411 (O_3411,N_49116,N_49915);
or UO_3412 (O_3412,N_49345,N_49580);
nor UO_3413 (O_3413,N_49185,N_49700);
xnor UO_3414 (O_3414,N_49410,N_49858);
nand UO_3415 (O_3415,N_49535,N_49865);
nor UO_3416 (O_3416,N_49876,N_49428);
xor UO_3417 (O_3417,N_49784,N_49433);
or UO_3418 (O_3418,N_49593,N_49802);
or UO_3419 (O_3419,N_49366,N_49126);
nor UO_3420 (O_3420,N_49312,N_49416);
and UO_3421 (O_3421,N_49269,N_49577);
nor UO_3422 (O_3422,N_49192,N_49312);
and UO_3423 (O_3423,N_49415,N_49047);
nor UO_3424 (O_3424,N_49851,N_49757);
xnor UO_3425 (O_3425,N_49441,N_49235);
nor UO_3426 (O_3426,N_49872,N_49354);
or UO_3427 (O_3427,N_49875,N_49121);
nor UO_3428 (O_3428,N_49851,N_49149);
nor UO_3429 (O_3429,N_49893,N_49781);
nor UO_3430 (O_3430,N_49374,N_49031);
nor UO_3431 (O_3431,N_49729,N_49793);
xnor UO_3432 (O_3432,N_49103,N_49417);
nand UO_3433 (O_3433,N_49884,N_49754);
xnor UO_3434 (O_3434,N_49887,N_49545);
nand UO_3435 (O_3435,N_49387,N_49468);
nand UO_3436 (O_3436,N_49986,N_49340);
xnor UO_3437 (O_3437,N_49177,N_49112);
nor UO_3438 (O_3438,N_49257,N_49865);
nand UO_3439 (O_3439,N_49250,N_49726);
or UO_3440 (O_3440,N_49051,N_49736);
and UO_3441 (O_3441,N_49460,N_49303);
nand UO_3442 (O_3442,N_49480,N_49917);
and UO_3443 (O_3443,N_49520,N_49025);
xnor UO_3444 (O_3444,N_49363,N_49078);
or UO_3445 (O_3445,N_49076,N_49306);
or UO_3446 (O_3446,N_49561,N_49684);
xnor UO_3447 (O_3447,N_49214,N_49626);
or UO_3448 (O_3448,N_49047,N_49947);
or UO_3449 (O_3449,N_49809,N_49135);
and UO_3450 (O_3450,N_49506,N_49578);
nor UO_3451 (O_3451,N_49454,N_49517);
nand UO_3452 (O_3452,N_49956,N_49804);
xor UO_3453 (O_3453,N_49371,N_49110);
xor UO_3454 (O_3454,N_49979,N_49918);
nor UO_3455 (O_3455,N_49125,N_49267);
nand UO_3456 (O_3456,N_49990,N_49126);
xor UO_3457 (O_3457,N_49068,N_49357);
or UO_3458 (O_3458,N_49564,N_49029);
or UO_3459 (O_3459,N_49794,N_49448);
xnor UO_3460 (O_3460,N_49408,N_49311);
or UO_3461 (O_3461,N_49497,N_49353);
nand UO_3462 (O_3462,N_49845,N_49762);
and UO_3463 (O_3463,N_49079,N_49043);
or UO_3464 (O_3464,N_49446,N_49164);
or UO_3465 (O_3465,N_49422,N_49898);
nor UO_3466 (O_3466,N_49196,N_49024);
nand UO_3467 (O_3467,N_49304,N_49347);
and UO_3468 (O_3468,N_49630,N_49319);
or UO_3469 (O_3469,N_49432,N_49563);
xor UO_3470 (O_3470,N_49523,N_49976);
nor UO_3471 (O_3471,N_49634,N_49118);
nor UO_3472 (O_3472,N_49537,N_49242);
or UO_3473 (O_3473,N_49928,N_49687);
nor UO_3474 (O_3474,N_49184,N_49806);
nor UO_3475 (O_3475,N_49299,N_49900);
nand UO_3476 (O_3476,N_49651,N_49750);
and UO_3477 (O_3477,N_49688,N_49133);
xnor UO_3478 (O_3478,N_49386,N_49749);
and UO_3479 (O_3479,N_49635,N_49206);
and UO_3480 (O_3480,N_49187,N_49763);
and UO_3481 (O_3481,N_49082,N_49490);
nand UO_3482 (O_3482,N_49485,N_49199);
and UO_3483 (O_3483,N_49828,N_49271);
and UO_3484 (O_3484,N_49695,N_49590);
xnor UO_3485 (O_3485,N_49778,N_49575);
and UO_3486 (O_3486,N_49232,N_49062);
or UO_3487 (O_3487,N_49738,N_49222);
or UO_3488 (O_3488,N_49000,N_49430);
nor UO_3489 (O_3489,N_49183,N_49504);
nand UO_3490 (O_3490,N_49956,N_49374);
nand UO_3491 (O_3491,N_49273,N_49069);
and UO_3492 (O_3492,N_49126,N_49506);
xnor UO_3493 (O_3493,N_49296,N_49918);
and UO_3494 (O_3494,N_49688,N_49893);
xor UO_3495 (O_3495,N_49397,N_49605);
nand UO_3496 (O_3496,N_49952,N_49799);
xor UO_3497 (O_3497,N_49525,N_49670);
nand UO_3498 (O_3498,N_49519,N_49137);
xor UO_3499 (O_3499,N_49481,N_49963);
nand UO_3500 (O_3500,N_49741,N_49002);
and UO_3501 (O_3501,N_49449,N_49211);
or UO_3502 (O_3502,N_49975,N_49048);
or UO_3503 (O_3503,N_49111,N_49965);
nor UO_3504 (O_3504,N_49358,N_49126);
nand UO_3505 (O_3505,N_49513,N_49455);
nand UO_3506 (O_3506,N_49605,N_49095);
or UO_3507 (O_3507,N_49712,N_49228);
nor UO_3508 (O_3508,N_49766,N_49130);
nand UO_3509 (O_3509,N_49734,N_49697);
or UO_3510 (O_3510,N_49213,N_49610);
xnor UO_3511 (O_3511,N_49171,N_49147);
or UO_3512 (O_3512,N_49012,N_49046);
or UO_3513 (O_3513,N_49214,N_49271);
nand UO_3514 (O_3514,N_49361,N_49692);
and UO_3515 (O_3515,N_49147,N_49078);
nand UO_3516 (O_3516,N_49422,N_49059);
xor UO_3517 (O_3517,N_49896,N_49887);
or UO_3518 (O_3518,N_49967,N_49432);
nand UO_3519 (O_3519,N_49395,N_49450);
or UO_3520 (O_3520,N_49560,N_49248);
or UO_3521 (O_3521,N_49804,N_49649);
and UO_3522 (O_3522,N_49969,N_49685);
nand UO_3523 (O_3523,N_49962,N_49199);
xor UO_3524 (O_3524,N_49816,N_49778);
nand UO_3525 (O_3525,N_49933,N_49398);
or UO_3526 (O_3526,N_49154,N_49253);
or UO_3527 (O_3527,N_49282,N_49578);
and UO_3528 (O_3528,N_49053,N_49599);
and UO_3529 (O_3529,N_49635,N_49706);
nand UO_3530 (O_3530,N_49464,N_49053);
and UO_3531 (O_3531,N_49715,N_49852);
nor UO_3532 (O_3532,N_49008,N_49608);
nor UO_3533 (O_3533,N_49016,N_49813);
xnor UO_3534 (O_3534,N_49362,N_49759);
xor UO_3535 (O_3535,N_49341,N_49388);
and UO_3536 (O_3536,N_49551,N_49022);
and UO_3537 (O_3537,N_49713,N_49200);
and UO_3538 (O_3538,N_49370,N_49861);
or UO_3539 (O_3539,N_49603,N_49506);
nor UO_3540 (O_3540,N_49638,N_49039);
and UO_3541 (O_3541,N_49295,N_49258);
nand UO_3542 (O_3542,N_49215,N_49464);
xor UO_3543 (O_3543,N_49584,N_49202);
xor UO_3544 (O_3544,N_49216,N_49757);
xor UO_3545 (O_3545,N_49184,N_49988);
or UO_3546 (O_3546,N_49330,N_49994);
or UO_3547 (O_3547,N_49173,N_49552);
nand UO_3548 (O_3548,N_49113,N_49044);
nor UO_3549 (O_3549,N_49172,N_49894);
xnor UO_3550 (O_3550,N_49401,N_49941);
nand UO_3551 (O_3551,N_49447,N_49051);
or UO_3552 (O_3552,N_49456,N_49306);
and UO_3553 (O_3553,N_49322,N_49220);
and UO_3554 (O_3554,N_49968,N_49663);
nor UO_3555 (O_3555,N_49094,N_49955);
nand UO_3556 (O_3556,N_49696,N_49508);
and UO_3557 (O_3557,N_49432,N_49584);
nand UO_3558 (O_3558,N_49809,N_49955);
nor UO_3559 (O_3559,N_49380,N_49303);
or UO_3560 (O_3560,N_49786,N_49487);
xor UO_3561 (O_3561,N_49861,N_49638);
xnor UO_3562 (O_3562,N_49940,N_49320);
xnor UO_3563 (O_3563,N_49765,N_49532);
nor UO_3564 (O_3564,N_49973,N_49324);
xor UO_3565 (O_3565,N_49100,N_49009);
nor UO_3566 (O_3566,N_49766,N_49747);
xnor UO_3567 (O_3567,N_49685,N_49830);
nand UO_3568 (O_3568,N_49635,N_49491);
or UO_3569 (O_3569,N_49225,N_49408);
nor UO_3570 (O_3570,N_49814,N_49691);
or UO_3571 (O_3571,N_49945,N_49472);
xor UO_3572 (O_3572,N_49661,N_49723);
and UO_3573 (O_3573,N_49180,N_49287);
and UO_3574 (O_3574,N_49094,N_49434);
nor UO_3575 (O_3575,N_49223,N_49672);
nand UO_3576 (O_3576,N_49060,N_49971);
and UO_3577 (O_3577,N_49606,N_49268);
nand UO_3578 (O_3578,N_49313,N_49126);
or UO_3579 (O_3579,N_49812,N_49285);
xor UO_3580 (O_3580,N_49982,N_49827);
nor UO_3581 (O_3581,N_49038,N_49714);
nand UO_3582 (O_3582,N_49040,N_49009);
xor UO_3583 (O_3583,N_49597,N_49052);
xnor UO_3584 (O_3584,N_49139,N_49143);
nand UO_3585 (O_3585,N_49985,N_49026);
nor UO_3586 (O_3586,N_49216,N_49563);
and UO_3587 (O_3587,N_49764,N_49557);
xor UO_3588 (O_3588,N_49165,N_49818);
nor UO_3589 (O_3589,N_49114,N_49007);
and UO_3590 (O_3590,N_49443,N_49722);
xnor UO_3591 (O_3591,N_49875,N_49389);
nor UO_3592 (O_3592,N_49975,N_49628);
and UO_3593 (O_3593,N_49616,N_49335);
xor UO_3594 (O_3594,N_49128,N_49203);
or UO_3595 (O_3595,N_49412,N_49601);
and UO_3596 (O_3596,N_49083,N_49997);
xor UO_3597 (O_3597,N_49671,N_49921);
nor UO_3598 (O_3598,N_49942,N_49230);
and UO_3599 (O_3599,N_49704,N_49194);
nand UO_3600 (O_3600,N_49649,N_49988);
nor UO_3601 (O_3601,N_49333,N_49098);
and UO_3602 (O_3602,N_49576,N_49484);
or UO_3603 (O_3603,N_49004,N_49709);
or UO_3604 (O_3604,N_49684,N_49011);
and UO_3605 (O_3605,N_49409,N_49257);
and UO_3606 (O_3606,N_49614,N_49112);
nor UO_3607 (O_3607,N_49992,N_49176);
and UO_3608 (O_3608,N_49626,N_49709);
and UO_3609 (O_3609,N_49652,N_49504);
or UO_3610 (O_3610,N_49082,N_49010);
nor UO_3611 (O_3611,N_49126,N_49248);
or UO_3612 (O_3612,N_49218,N_49938);
or UO_3613 (O_3613,N_49083,N_49082);
or UO_3614 (O_3614,N_49724,N_49238);
nand UO_3615 (O_3615,N_49733,N_49075);
or UO_3616 (O_3616,N_49560,N_49110);
or UO_3617 (O_3617,N_49455,N_49831);
or UO_3618 (O_3618,N_49962,N_49053);
nand UO_3619 (O_3619,N_49649,N_49659);
nand UO_3620 (O_3620,N_49653,N_49213);
nand UO_3621 (O_3621,N_49947,N_49324);
xnor UO_3622 (O_3622,N_49345,N_49009);
xor UO_3623 (O_3623,N_49083,N_49440);
or UO_3624 (O_3624,N_49498,N_49911);
xnor UO_3625 (O_3625,N_49655,N_49820);
or UO_3626 (O_3626,N_49366,N_49399);
or UO_3627 (O_3627,N_49643,N_49222);
nor UO_3628 (O_3628,N_49523,N_49133);
nor UO_3629 (O_3629,N_49007,N_49428);
xor UO_3630 (O_3630,N_49894,N_49808);
and UO_3631 (O_3631,N_49653,N_49981);
nor UO_3632 (O_3632,N_49908,N_49311);
and UO_3633 (O_3633,N_49025,N_49097);
xnor UO_3634 (O_3634,N_49757,N_49232);
or UO_3635 (O_3635,N_49847,N_49291);
or UO_3636 (O_3636,N_49047,N_49839);
xnor UO_3637 (O_3637,N_49661,N_49645);
or UO_3638 (O_3638,N_49568,N_49611);
nor UO_3639 (O_3639,N_49903,N_49626);
xnor UO_3640 (O_3640,N_49336,N_49088);
nand UO_3641 (O_3641,N_49612,N_49378);
and UO_3642 (O_3642,N_49719,N_49050);
nor UO_3643 (O_3643,N_49524,N_49405);
or UO_3644 (O_3644,N_49635,N_49259);
nand UO_3645 (O_3645,N_49228,N_49423);
nor UO_3646 (O_3646,N_49336,N_49461);
nor UO_3647 (O_3647,N_49447,N_49135);
nor UO_3648 (O_3648,N_49684,N_49718);
nand UO_3649 (O_3649,N_49283,N_49269);
nand UO_3650 (O_3650,N_49351,N_49800);
nor UO_3651 (O_3651,N_49153,N_49542);
and UO_3652 (O_3652,N_49004,N_49589);
nor UO_3653 (O_3653,N_49019,N_49770);
or UO_3654 (O_3654,N_49432,N_49834);
and UO_3655 (O_3655,N_49005,N_49491);
or UO_3656 (O_3656,N_49489,N_49375);
nand UO_3657 (O_3657,N_49814,N_49132);
xor UO_3658 (O_3658,N_49448,N_49311);
xor UO_3659 (O_3659,N_49607,N_49729);
or UO_3660 (O_3660,N_49496,N_49267);
xnor UO_3661 (O_3661,N_49318,N_49582);
nand UO_3662 (O_3662,N_49071,N_49254);
nor UO_3663 (O_3663,N_49328,N_49081);
nor UO_3664 (O_3664,N_49009,N_49210);
nand UO_3665 (O_3665,N_49256,N_49828);
nor UO_3666 (O_3666,N_49773,N_49212);
nor UO_3667 (O_3667,N_49624,N_49019);
and UO_3668 (O_3668,N_49103,N_49462);
xor UO_3669 (O_3669,N_49231,N_49674);
nor UO_3670 (O_3670,N_49791,N_49343);
xnor UO_3671 (O_3671,N_49197,N_49602);
or UO_3672 (O_3672,N_49486,N_49104);
nand UO_3673 (O_3673,N_49908,N_49440);
and UO_3674 (O_3674,N_49237,N_49052);
or UO_3675 (O_3675,N_49163,N_49257);
xor UO_3676 (O_3676,N_49583,N_49504);
xor UO_3677 (O_3677,N_49554,N_49207);
nor UO_3678 (O_3678,N_49620,N_49579);
or UO_3679 (O_3679,N_49723,N_49058);
nand UO_3680 (O_3680,N_49068,N_49468);
nand UO_3681 (O_3681,N_49275,N_49962);
or UO_3682 (O_3682,N_49258,N_49912);
nor UO_3683 (O_3683,N_49465,N_49371);
or UO_3684 (O_3684,N_49193,N_49660);
nor UO_3685 (O_3685,N_49626,N_49658);
xor UO_3686 (O_3686,N_49490,N_49805);
nor UO_3687 (O_3687,N_49022,N_49412);
xnor UO_3688 (O_3688,N_49501,N_49578);
nor UO_3689 (O_3689,N_49721,N_49007);
xnor UO_3690 (O_3690,N_49801,N_49786);
nand UO_3691 (O_3691,N_49837,N_49890);
or UO_3692 (O_3692,N_49118,N_49245);
nand UO_3693 (O_3693,N_49931,N_49927);
or UO_3694 (O_3694,N_49330,N_49100);
or UO_3695 (O_3695,N_49208,N_49753);
xnor UO_3696 (O_3696,N_49197,N_49282);
and UO_3697 (O_3697,N_49008,N_49252);
xnor UO_3698 (O_3698,N_49705,N_49212);
and UO_3699 (O_3699,N_49624,N_49119);
and UO_3700 (O_3700,N_49541,N_49486);
nand UO_3701 (O_3701,N_49219,N_49482);
nor UO_3702 (O_3702,N_49361,N_49204);
nand UO_3703 (O_3703,N_49544,N_49950);
nand UO_3704 (O_3704,N_49294,N_49191);
or UO_3705 (O_3705,N_49651,N_49683);
xor UO_3706 (O_3706,N_49519,N_49997);
xnor UO_3707 (O_3707,N_49261,N_49709);
nor UO_3708 (O_3708,N_49941,N_49800);
nor UO_3709 (O_3709,N_49870,N_49027);
nand UO_3710 (O_3710,N_49741,N_49853);
nor UO_3711 (O_3711,N_49539,N_49253);
or UO_3712 (O_3712,N_49368,N_49044);
xnor UO_3713 (O_3713,N_49614,N_49629);
nor UO_3714 (O_3714,N_49563,N_49306);
nand UO_3715 (O_3715,N_49381,N_49856);
nand UO_3716 (O_3716,N_49148,N_49803);
nor UO_3717 (O_3717,N_49694,N_49339);
or UO_3718 (O_3718,N_49019,N_49222);
nand UO_3719 (O_3719,N_49801,N_49255);
or UO_3720 (O_3720,N_49728,N_49827);
xnor UO_3721 (O_3721,N_49673,N_49451);
nor UO_3722 (O_3722,N_49938,N_49873);
nand UO_3723 (O_3723,N_49094,N_49564);
nor UO_3724 (O_3724,N_49531,N_49165);
nand UO_3725 (O_3725,N_49623,N_49083);
or UO_3726 (O_3726,N_49494,N_49087);
xor UO_3727 (O_3727,N_49182,N_49240);
nand UO_3728 (O_3728,N_49393,N_49145);
and UO_3729 (O_3729,N_49955,N_49646);
or UO_3730 (O_3730,N_49188,N_49743);
xnor UO_3731 (O_3731,N_49340,N_49104);
and UO_3732 (O_3732,N_49890,N_49372);
nand UO_3733 (O_3733,N_49900,N_49666);
xnor UO_3734 (O_3734,N_49892,N_49636);
and UO_3735 (O_3735,N_49547,N_49289);
or UO_3736 (O_3736,N_49872,N_49109);
nor UO_3737 (O_3737,N_49891,N_49439);
or UO_3738 (O_3738,N_49028,N_49896);
nand UO_3739 (O_3739,N_49034,N_49746);
or UO_3740 (O_3740,N_49765,N_49824);
nor UO_3741 (O_3741,N_49469,N_49409);
or UO_3742 (O_3742,N_49877,N_49037);
nand UO_3743 (O_3743,N_49598,N_49567);
and UO_3744 (O_3744,N_49968,N_49266);
xor UO_3745 (O_3745,N_49593,N_49549);
and UO_3746 (O_3746,N_49880,N_49017);
or UO_3747 (O_3747,N_49533,N_49410);
xnor UO_3748 (O_3748,N_49403,N_49277);
xnor UO_3749 (O_3749,N_49811,N_49198);
xor UO_3750 (O_3750,N_49984,N_49606);
or UO_3751 (O_3751,N_49280,N_49035);
nor UO_3752 (O_3752,N_49668,N_49503);
nand UO_3753 (O_3753,N_49824,N_49078);
and UO_3754 (O_3754,N_49904,N_49624);
nor UO_3755 (O_3755,N_49979,N_49656);
nand UO_3756 (O_3756,N_49758,N_49220);
or UO_3757 (O_3757,N_49084,N_49971);
xnor UO_3758 (O_3758,N_49619,N_49788);
xor UO_3759 (O_3759,N_49159,N_49046);
or UO_3760 (O_3760,N_49231,N_49715);
nor UO_3761 (O_3761,N_49754,N_49408);
xor UO_3762 (O_3762,N_49420,N_49212);
and UO_3763 (O_3763,N_49422,N_49077);
nand UO_3764 (O_3764,N_49903,N_49733);
nand UO_3765 (O_3765,N_49044,N_49750);
xnor UO_3766 (O_3766,N_49734,N_49477);
nand UO_3767 (O_3767,N_49354,N_49127);
xnor UO_3768 (O_3768,N_49134,N_49560);
nor UO_3769 (O_3769,N_49221,N_49272);
nand UO_3770 (O_3770,N_49316,N_49545);
and UO_3771 (O_3771,N_49289,N_49831);
and UO_3772 (O_3772,N_49314,N_49807);
xor UO_3773 (O_3773,N_49961,N_49321);
nor UO_3774 (O_3774,N_49678,N_49757);
and UO_3775 (O_3775,N_49576,N_49591);
nand UO_3776 (O_3776,N_49081,N_49982);
nor UO_3777 (O_3777,N_49423,N_49578);
or UO_3778 (O_3778,N_49328,N_49474);
nor UO_3779 (O_3779,N_49671,N_49455);
nand UO_3780 (O_3780,N_49443,N_49817);
xnor UO_3781 (O_3781,N_49599,N_49311);
and UO_3782 (O_3782,N_49777,N_49364);
nor UO_3783 (O_3783,N_49763,N_49121);
nand UO_3784 (O_3784,N_49507,N_49291);
or UO_3785 (O_3785,N_49058,N_49518);
and UO_3786 (O_3786,N_49431,N_49038);
nand UO_3787 (O_3787,N_49604,N_49504);
nor UO_3788 (O_3788,N_49742,N_49027);
nand UO_3789 (O_3789,N_49754,N_49170);
xnor UO_3790 (O_3790,N_49762,N_49136);
nand UO_3791 (O_3791,N_49095,N_49505);
or UO_3792 (O_3792,N_49723,N_49034);
and UO_3793 (O_3793,N_49188,N_49118);
or UO_3794 (O_3794,N_49446,N_49515);
nand UO_3795 (O_3795,N_49790,N_49910);
or UO_3796 (O_3796,N_49809,N_49010);
nor UO_3797 (O_3797,N_49686,N_49529);
xnor UO_3798 (O_3798,N_49543,N_49883);
nand UO_3799 (O_3799,N_49192,N_49777);
and UO_3800 (O_3800,N_49180,N_49405);
and UO_3801 (O_3801,N_49692,N_49689);
nor UO_3802 (O_3802,N_49501,N_49751);
xor UO_3803 (O_3803,N_49512,N_49459);
xnor UO_3804 (O_3804,N_49298,N_49182);
nor UO_3805 (O_3805,N_49849,N_49516);
nor UO_3806 (O_3806,N_49723,N_49302);
xnor UO_3807 (O_3807,N_49596,N_49146);
nand UO_3808 (O_3808,N_49009,N_49023);
xor UO_3809 (O_3809,N_49793,N_49703);
xnor UO_3810 (O_3810,N_49889,N_49707);
and UO_3811 (O_3811,N_49562,N_49776);
or UO_3812 (O_3812,N_49796,N_49913);
and UO_3813 (O_3813,N_49360,N_49017);
nand UO_3814 (O_3814,N_49042,N_49288);
xnor UO_3815 (O_3815,N_49740,N_49468);
and UO_3816 (O_3816,N_49787,N_49059);
nor UO_3817 (O_3817,N_49907,N_49330);
and UO_3818 (O_3818,N_49208,N_49812);
or UO_3819 (O_3819,N_49211,N_49093);
and UO_3820 (O_3820,N_49185,N_49508);
nand UO_3821 (O_3821,N_49224,N_49815);
and UO_3822 (O_3822,N_49625,N_49308);
nand UO_3823 (O_3823,N_49475,N_49092);
nand UO_3824 (O_3824,N_49230,N_49594);
and UO_3825 (O_3825,N_49077,N_49693);
or UO_3826 (O_3826,N_49074,N_49274);
nor UO_3827 (O_3827,N_49062,N_49693);
xor UO_3828 (O_3828,N_49111,N_49177);
nand UO_3829 (O_3829,N_49164,N_49619);
or UO_3830 (O_3830,N_49558,N_49025);
and UO_3831 (O_3831,N_49239,N_49627);
nor UO_3832 (O_3832,N_49681,N_49812);
or UO_3833 (O_3833,N_49630,N_49055);
nand UO_3834 (O_3834,N_49465,N_49901);
or UO_3835 (O_3835,N_49943,N_49083);
nor UO_3836 (O_3836,N_49463,N_49159);
or UO_3837 (O_3837,N_49057,N_49249);
xor UO_3838 (O_3838,N_49609,N_49460);
xnor UO_3839 (O_3839,N_49446,N_49549);
nor UO_3840 (O_3840,N_49090,N_49855);
or UO_3841 (O_3841,N_49996,N_49540);
xor UO_3842 (O_3842,N_49338,N_49953);
or UO_3843 (O_3843,N_49779,N_49334);
nand UO_3844 (O_3844,N_49850,N_49720);
or UO_3845 (O_3845,N_49549,N_49631);
nand UO_3846 (O_3846,N_49956,N_49092);
or UO_3847 (O_3847,N_49191,N_49145);
and UO_3848 (O_3848,N_49733,N_49813);
nor UO_3849 (O_3849,N_49176,N_49570);
and UO_3850 (O_3850,N_49667,N_49682);
xnor UO_3851 (O_3851,N_49851,N_49662);
or UO_3852 (O_3852,N_49093,N_49920);
or UO_3853 (O_3853,N_49041,N_49124);
or UO_3854 (O_3854,N_49700,N_49398);
xor UO_3855 (O_3855,N_49950,N_49234);
and UO_3856 (O_3856,N_49341,N_49126);
or UO_3857 (O_3857,N_49070,N_49858);
xnor UO_3858 (O_3858,N_49671,N_49652);
nor UO_3859 (O_3859,N_49902,N_49332);
nand UO_3860 (O_3860,N_49944,N_49702);
nand UO_3861 (O_3861,N_49924,N_49068);
nor UO_3862 (O_3862,N_49295,N_49563);
and UO_3863 (O_3863,N_49695,N_49328);
nand UO_3864 (O_3864,N_49365,N_49933);
nand UO_3865 (O_3865,N_49988,N_49018);
xor UO_3866 (O_3866,N_49502,N_49898);
or UO_3867 (O_3867,N_49502,N_49831);
nor UO_3868 (O_3868,N_49486,N_49309);
xnor UO_3869 (O_3869,N_49171,N_49448);
and UO_3870 (O_3870,N_49061,N_49959);
and UO_3871 (O_3871,N_49057,N_49972);
and UO_3872 (O_3872,N_49345,N_49218);
xnor UO_3873 (O_3873,N_49859,N_49199);
nor UO_3874 (O_3874,N_49233,N_49013);
nand UO_3875 (O_3875,N_49072,N_49008);
and UO_3876 (O_3876,N_49848,N_49493);
xnor UO_3877 (O_3877,N_49789,N_49839);
nor UO_3878 (O_3878,N_49513,N_49667);
nor UO_3879 (O_3879,N_49963,N_49091);
nor UO_3880 (O_3880,N_49821,N_49543);
and UO_3881 (O_3881,N_49414,N_49569);
xor UO_3882 (O_3882,N_49551,N_49519);
xnor UO_3883 (O_3883,N_49093,N_49921);
xor UO_3884 (O_3884,N_49919,N_49791);
nor UO_3885 (O_3885,N_49395,N_49881);
nor UO_3886 (O_3886,N_49671,N_49292);
nor UO_3887 (O_3887,N_49151,N_49462);
xor UO_3888 (O_3888,N_49343,N_49037);
xnor UO_3889 (O_3889,N_49940,N_49933);
and UO_3890 (O_3890,N_49330,N_49367);
nand UO_3891 (O_3891,N_49736,N_49594);
xor UO_3892 (O_3892,N_49251,N_49634);
xnor UO_3893 (O_3893,N_49519,N_49087);
and UO_3894 (O_3894,N_49793,N_49207);
nand UO_3895 (O_3895,N_49901,N_49857);
or UO_3896 (O_3896,N_49298,N_49223);
nor UO_3897 (O_3897,N_49154,N_49035);
xor UO_3898 (O_3898,N_49639,N_49363);
or UO_3899 (O_3899,N_49622,N_49710);
xnor UO_3900 (O_3900,N_49932,N_49653);
nor UO_3901 (O_3901,N_49713,N_49024);
xnor UO_3902 (O_3902,N_49224,N_49742);
nor UO_3903 (O_3903,N_49539,N_49763);
or UO_3904 (O_3904,N_49477,N_49590);
or UO_3905 (O_3905,N_49551,N_49490);
xnor UO_3906 (O_3906,N_49856,N_49476);
or UO_3907 (O_3907,N_49258,N_49107);
or UO_3908 (O_3908,N_49133,N_49788);
or UO_3909 (O_3909,N_49805,N_49891);
and UO_3910 (O_3910,N_49447,N_49799);
or UO_3911 (O_3911,N_49003,N_49859);
and UO_3912 (O_3912,N_49141,N_49259);
nor UO_3913 (O_3913,N_49613,N_49516);
nand UO_3914 (O_3914,N_49109,N_49818);
and UO_3915 (O_3915,N_49761,N_49507);
xnor UO_3916 (O_3916,N_49087,N_49835);
nor UO_3917 (O_3917,N_49372,N_49751);
xor UO_3918 (O_3918,N_49264,N_49160);
xnor UO_3919 (O_3919,N_49254,N_49124);
and UO_3920 (O_3920,N_49642,N_49390);
or UO_3921 (O_3921,N_49949,N_49805);
or UO_3922 (O_3922,N_49717,N_49603);
and UO_3923 (O_3923,N_49212,N_49337);
xor UO_3924 (O_3924,N_49425,N_49847);
nor UO_3925 (O_3925,N_49562,N_49524);
nor UO_3926 (O_3926,N_49450,N_49004);
nand UO_3927 (O_3927,N_49174,N_49565);
xnor UO_3928 (O_3928,N_49741,N_49909);
or UO_3929 (O_3929,N_49377,N_49256);
nor UO_3930 (O_3930,N_49903,N_49654);
nor UO_3931 (O_3931,N_49705,N_49424);
xnor UO_3932 (O_3932,N_49347,N_49314);
and UO_3933 (O_3933,N_49963,N_49349);
nand UO_3934 (O_3934,N_49366,N_49717);
and UO_3935 (O_3935,N_49783,N_49946);
and UO_3936 (O_3936,N_49541,N_49712);
nor UO_3937 (O_3937,N_49872,N_49081);
or UO_3938 (O_3938,N_49671,N_49410);
nand UO_3939 (O_3939,N_49594,N_49364);
or UO_3940 (O_3940,N_49350,N_49332);
or UO_3941 (O_3941,N_49700,N_49475);
nand UO_3942 (O_3942,N_49595,N_49312);
nand UO_3943 (O_3943,N_49348,N_49700);
xnor UO_3944 (O_3944,N_49857,N_49382);
nor UO_3945 (O_3945,N_49821,N_49293);
xnor UO_3946 (O_3946,N_49793,N_49504);
xnor UO_3947 (O_3947,N_49834,N_49381);
and UO_3948 (O_3948,N_49538,N_49965);
nor UO_3949 (O_3949,N_49583,N_49722);
nor UO_3950 (O_3950,N_49650,N_49333);
and UO_3951 (O_3951,N_49161,N_49668);
xor UO_3952 (O_3952,N_49227,N_49384);
nor UO_3953 (O_3953,N_49629,N_49273);
xnor UO_3954 (O_3954,N_49812,N_49058);
nor UO_3955 (O_3955,N_49017,N_49791);
or UO_3956 (O_3956,N_49411,N_49861);
xor UO_3957 (O_3957,N_49083,N_49897);
nor UO_3958 (O_3958,N_49554,N_49685);
nor UO_3959 (O_3959,N_49140,N_49896);
nor UO_3960 (O_3960,N_49415,N_49019);
or UO_3961 (O_3961,N_49697,N_49285);
and UO_3962 (O_3962,N_49484,N_49952);
nor UO_3963 (O_3963,N_49131,N_49092);
xnor UO_3964 (O_3964,N_49982,N_49273);
xor UO_3965 (O_3965,N_49256,N_49941);
or UO_3966 (O_3966,N_49851,N_49346);
and UO_3967 (O_3967,N_49762,N_49969);
xor UO_3968 (O_3968,N_49964,N_49776);
xnor UO_3969 (O_3969,N_49275,N_49893);
or UO_3970 (O_3970,N_49419,N_49174);
or UO_3971 (O_3971,N_49311,N_49391);
nor UO_3972 (O_3972,N_49677,N_49701);
nor UO_3973 (O_3973,N_49230,N_49108);
and UO_3974 (O_3974,N_49068,N_49654);
xor UO_3975 (O_3975,N_49814,N_49730);
nand UO_3976 (O_3976,N_49536,N_49244);
xor UO_3977 (O_3977,N_49849,N_49299);
xor UO_3978 (O_3978,N_49691,N_49945);
nor UO_3979 (O_3979,N_49382,N_49327);
and UO_3980 (O_3980,N_49690,N_49987);
nand UO_3981 (O_3981,N_49782,N_49705);
nand UO_3982 (O_3982,N_49346,N_49332);
xor UO_3983 (O_3983,N_49257,N_49365);
and UO_3984 (O_3984,N_49764,N_49653);
nor UO_3985 (O_3985,N_49871,N_49737);
or UO_3986 (O_3986,N_49597,N_49673);
nor UO_3987 (O_3987,N_49158,N_49948);
nand UO_3988 (O_3988,N_49246,N_49044);
nor UO_3989 (O_3989,N_49539,N_49919);
xnor UO_3990 (O_3990,N_49137,N_49579);
nand UO_3991 (O_3991,N_49276,N_49934);
and UO_3992 (O_3992,N_49060,N_49084);
or UO_3993 (O_3993,N_49273,N_49215);
xor UO_3994 (O_3994,N_49745,N_49501);
nor UO_3995 (O_3995,N_49753,N_49419);
or UO_3996 (O_3996,N_49476,N_49767);
nor UO_3997 (O_3997,N_49626,N_49357);
and UO_3998 (O_3998,N_49794,N_49924);
nor UO_3999 (O_3999,N_49644,N_49332);
xor UO_4000 (O_4000,N_49863,N_49827);
or UO_4001 (O_4001,N_49059,N_49314);
nand UO_4002 (O_4002,N_49226,N_49067);
nor UO_4003 (O_4003,N_49254,N_49088);
or UO_4004 (O_4004,N_49180,N_49209);
nor UO_4005 (O_4005,N_49216,N_49758);
xor UO_4006 (O_4006,N_49863,N_49009);
nor UO_4007 (O_4007,N_49519,N_49870);
nand UO_4008 (O_4008,N_49338,N_49849);
xor UO_4009 (O_4009,N_49740,N_49199);
nor UO_4010 (O_4010,N_49942,N_49184);
and UO_4011 (O_4011,N_49350,N_49477);
xnor UO_4012 (O_4012,N_49825,N_49939);
nor UO_4013 (O_4013,N_49726,N_49716);
or UO_4014 (O_4014,N_49163,N_49208);
and UO_4015 (O_4015,N_49597,N_49963);
nor UO_4016 (O_4016,N_49459,N_49047);
xor UO_4017 (O_4017,N_49536,N_49593);
xor UO_4018 (O_4018,N_49482,N_49029);
nand UO_4019 (O_4019,N_49798,N_49302);
nand UO_4020 (O_4020,N_49334,N_49040);
nor UO_4021 (O_4021,N_49386,N_49070);
or UO_4022 (O_4022,N_49230,N_49252);
nand UO_4023 (O_4023,N_49737,N_49612);
or UO_4024 (O_4024,N_49311,N_49746);
and UO_4025 (O_4025,N_49365,N_49246);
and UO_4026 (O_4026,N_49019,N_49787);
xnor UO_4027 (O_4027,N_49073,N_49607);
nor UO_4028 (O_4028,N_49480,N_49437);
or UO_4029 (O_4029,N_49117,N_49825);
and UO_4030 (O_4030,N_49515,N_49460);
nand UO_4031 (O_4031,N_49735,N_49632);
and UO_4032 (O_4032,N_49253,N_49920);
or UO_4033 (O_4033,N_49784,N_49983);
or UO_4034 (O_4034,N_49363,N_49520);
and UO_4035 (O_4035,N_49922,N_49638);
xnor UO_4036 (O_4036,N_49685,N_49370);
or UO_4037 (O_4037,N_49614,N_49399);
nand UO_4038 (O_4038,N_49002,N_49579);
nor UO_4039 (O_4039,N_49511,N_49288);
and UO_4040 (O_4040,N_49035,N_49338);
or UO_4041 (O_4041,N_49164,N_49105);
or UO_4042 (O_4042,N_49624,N_49163);
or UO_4043 (O_4043,N_49881,N_49234);
or UO_4044 (O_4044,N_49281,N_49244);
nand UO_4045 (O_4045,N_49675,N_49255);
xnor UO_4046 (O_4046,N_49856,N_49138);
nand UO_4047 (O_4047,N_49265,N_49049);
and UO_4048 (O_4048,N_49326,N_49446);
xnor UO_4049 (O_4049,N_49395,N_49412);
nand UO_4050 (O_4050,N_49564,N_49474);
nand UO_4051 (O_4051,N_49306,N_49340);
nor UO_4052 (O_4052,N_49206,N_49239);
xor UO_4053 (O_4053,N_49751,N_49061);
and UO_4054 (O_4054,N_49747,N_49288);
or UO_4055 (O_4055,N_49218,N_49567);
nand UO_4056 (O_4056,N_49695,N_49550);
and UO_4057 (O_4057,N_49357,N_49505);
nor UO_4058 (O_4058,N_49328,N_49492);
and UO_4059 (O_4059,N_49650,N_49096);
xnor UO_4060 (O_4060,N_49901,N_49871);
and UO_4061 (O_4061,N_49390,N_49608);
or UO_4062 (O_4062,N_49192,N_49604);
nor UO_4063 (O_4063,N_49823,N_49499);
or UO_4064 (O_4064,N_49784,N_49174);
and UO_4065 (O_4065,N_49047,N_49596);
nand UO_4066 (O_4066,N_49128,N_49529);
nor UO_4067 (O_4067,N_49619,N_49186);
nor UO_4068 (O_4068,N_49141,N_49242);
nor UO_4069 (O_4069,N_49477,N_49712);
xnor UO_4070 (O_4070,N_49275,N_49680);
nand UO_4071 (O_4071,N_49438,N_49783);
nor UO_4072 (O_4072,N_49394,N_49071);
and UO_4073 (O_4073,N_49363,N_49374);
nand UO_4074 (O_4074,N_49523,N_49909);
nand UO_4075 (O_4075,N_49937,N_49795);
xnor UO_4076 (O_4076,N_49570,N_49319);
or UO_4077 (O_4077,N_49622,N_49343);
nand UO_4078 (O_4078,N_49841,N_49955);
and UO_4079 (O_4079,N_49247,N_49288);
nand UO_4080 (O_4080,N_49152,N_49251);
or UO_4081 (O_4081,N_49951,N_49862);
or UO_4082 (O_4082,N_49829,N_49919);
nand UO_4083 (O_4083,N_49974,N_49242);
and UO_4084 (O_4084,N_49642,N_49909);
and UO_4085 (O_4085,N_49828,N_49711);
and UO_4086 (O_4086,N_49212,N_49881);
or UO_4087 (O_4087,N_49678,N_49010);
and UO_4088 (O_4088,N_49133,N_49569);
nor UO_4089 (O_4089,N_49259,N_49077);
xor UO_4090 (O_4090,N_49086,N_49227);
nand UO_4091 (O_4091,N_49897,N_49901);
xor UO_4092 (O_4092,N_49925,N_49995);
xnor UO_4093 (O_4093,N_49759,N_49143);
or UO_4094 (O_4094,N_49898,N_49287);
nand UO_4095 (O_4095,N_49058,N_49623);
and UO_4096 (O_4096,N_49073,N_49558);
nor UO_4097 (O_4097,N_49336,N_49061);
and UO_4098 (O_4098,N_49371,N_49766);
nand UO_4099 (O_4099,N_49546,N_49515);
nand UO_4100 (O_4100,N_49072,N_49343);
nand UO_4101 (O_4101,N_49623,N_49621);
nor UO_4102 (O_4102,N_49265,N_49962);
and UO_4103 (O_4103,N_49205,N_49142);
and UO_4104 (O_4104,N_49528,N_49891);
or UO_4105 (O_4105,N_49981,N_49411);
or UO_4106 (O_4106,N_49348,N_49016);
or UO_4107 (O_4107,N_49048,N_49879);
nor UO_4108 (O_4108,N_49081,N_49140);
nor UO_4109 (O_4109,N_49949,N_49483);
nor UO_4110 (O_4110,N_49404,N_49670);
nor UO_4111 (O_4111,N_49282,N_49885);
and UO_4112 (O_4112,N_49535,N_49436);
nor UO_4113 (O_4113,N_49574,N_49430);
nand UO_4114 (O_4114,N_49777,N_49215);
or UO_4115 (O_4115,N_49163,N_49300);
and UO_4116 (O_4116,N_49175,N_49952);
nor UO_4117 (O_4117,N_49539,N_49458);
nor UO_4118 (O_4118,N_49885,N_49259);
xor UO_4119 (O_4119,N_49311,N_49712);
nor UO_4120 (O_4120,N_49735,N_49974);
xnor UO_4121 (O_4121,N_49663,N_49813);
and UO_4122 (O_4122,N_49474,N_49148);
nor UO_4123 (O_4123,N_49335,N_49745);
nand UO_4124 (O_4124,N_49438,N_49046);
and UO_4125 (O_4125,N_49796,N_49699);
nand UO_4126 (O_4126,N_49783,N_49265);
nor UO_4127 (O_4127,N_49576,N_49946);
nand UO_4128 (O_4128,N_49411,N_49998);
xnor UO_4129 (O_4129,N_49678,N_49337);
or UO_4130 (O_4130,N_49485,N_49440);
or UO_4131 (O_4131,N_49695,N_49252);
xnor UO_4132 (O_4132,N_49360,N_49768);
nand UO_4133 (O_4133,N_49473,N_49204);
or UO_4134 (O_4134,N_49171,N_49117);
nor UO_4135 (O_4135,N_49566,N_49013);
nor UO_4136 (O_4136,N_49089,N_49139);
nor UO_4137 (O_4137,N_49296,N_49938);
and UO_4138 (O_4138,N_49541,N_49642);
or UO_4139 (O_4139,N_49592,N_49211);
nor UO_4140 (O_4140,N_49456,N_49243);
nor UO_4141 (O_4141,N_49953,N_49430);
nand UO_4142 (O_4142,N_49827,N_49644);
and UO_4143 (O_4143,N_49628,N_49354);
xnor UO_4144 (O_4144,N_49806,N_49655);
and UO_4145 (O_4145,N_49139,N_49852);
nand UO_4146 (O_4146,N_49545,N_49344);
and UO_4147 (O_4147,N_49839,N_49931);
nand UO_4148 (O_4148,N_49692,N_49959);
or UO_4149 (O_4149,N_49428,N_49091);
nor UO_4150 (O_4150,N_49486,N_49600);
or UO_4151 (O_4151,N_49362,N_49091);
or UO_4152 (O_4152,N_49660,N_49955);
nor UO_4153 (O_4153,N_49177,N_49327);
or UO_4154 (O_4154,N_49703,N_49864);
and UO_4155 (O_4155,N_49645,N_49471);
xnor UO_4156 (O_4156,N_49469,N_49470);
xor UO_4157 (O_4157,N_49685,N_49819);
or UO_4158 (O_4158,N_49338,N_49326);
xor UO_4159 (O_4159,N_49196,N_49867);
or UO_4160 (O_4160,N_49583,N_49533);
nand UO_4161 (O_4161,N_49617,N_49983);
nand UO_4162 (O_4162,N_49922,N_49539);
or UO_4163 (O_4163,N_49483,N_49894);
nand UO_4164 (O_4164,N_49187,N_49095);
and UO_4165 (O_4165,N_49256,N_49499);
nor UO_4166 (O_4166,N_49259,N_49204);
nand UO_4167 (O_4167,N_49003,N_49948);
nand UO_4168 (O_4168,N_49903,N_49627);
or UO_4169 (O_4169,N_49310,N_49577);
or UO_4170 (O_4170,N_49079,N_49438);
nand UO_4171 (O_4171,N_49606,N_49577);
or UO_4172 (O_4172,N_49022,N_49031);
or UO_4173 (O_4173,N_49912,N_49756);
nor UO_4174 (O_4174,N_49669,N_49011);
xnor UO_4175 (O_4175,N_49988,N_49843);
xnor UO_4176 (O_4176,N_49972,N_49447);
and UO_4177 (O_4177,N_49516,N_49302);
xnor UO_4178 (O_4178,N_49996,N_49871);
nor UO_4179 (O_4179,N_49522,N_49622);
and UO_4180 (O_4180,N_49716,N_49287);
or UO_4181 (O_4181,N_49023,N_49371);
and UO_4182 (O_4182,N_49381,N_49733);
xor UO_4183 (O_4183,N_49135,N_49068);
and UO_4184 (O_4184,N_49852,N_49965);
and UO_4185 (O_4185,N_49199,N_49540);
nand UO_4186 (O_4186,N_49931,N_49410);
nor UO_4187 (O_4187,N_49988,N_49904);
nand UO_4188 (O_4188,N_49742,N_49061);
and UO_4189 (O_4189,N_49702,N_49300);
and UO_4190 (O_4190,N_49161,N_49593);
xnor UO_4191 (O_4191,N_49381,N_49868);
xor UO_4192 (O_4192,N_49181,N_49905);
and UO_4193 (O_4193,N_49312,N_49380);
nand UO_4194 (O_4194,N_49637,N_49964);
nand UO_4195 (O_4195,N_49234,N_49956);
and UO_4196 (O_4196,N_49966,N_49198);
or UO_4197 (O_4197,N_49260,N_49987);
or UO_4198 (O_4198,N_49286,N_49452);
nand UO_4199 (O_4199,N_49367,N_49004);
or UO_4200 (O_4200,N_49026,N_49941);
nor UO_4201 (O_4201,N_49219,N_49289);
nor UO_4202 (O_4202,N_49294,N_49633);
or UO_4203 (O_4203,N_49081,N_49307);
and UO_4204 (O_4204,N_49640,N_49294);
nand UO_4205 (O_4205,N_49545,N_49836);
and UO_4206 (O_4206,N_49140,N_49131);
and UO_4207 (O_4207,N_49141,N_49903);
or UO_4208 (O_4208,N_49009,N_49790);
and UO_4209 (O_4209,N_49406,N_49618);
nor UO_4210 (O_4210,N_49860,N_49580);
nor UO_4211 (O_4211,N_49911,N_49708);
or UO_4212 (O_4212,N_49142,N_49402);
or UO_4213 (O_4213,N_49264,N_49809);
or UO_4214 (O_4214,N_49861,N_49347);
nor UO_4215 (O_4215,N_49658,N_49089);
nand UO_4216 (O_4216,N_49897,N_49976);
xnor UO_4217 (O_4217,N_49951,N_49462);
and UO_4218 (O_4218,N_49299,N_49288);
and UO_4219 (O_4219,N_49375,N_49360);
xor UO_4220 (O_4220,N_49367,N_49258);
xor UO_4221 (O_4221,N_49908,N_49207);
and UO_4222 (O_4222,N_49307,N_49544);
xnor UO_4223 (O_4223,N_49487,N_49022);
nand UO_4224 (O_4224,N_49203,N_49906);
and UO_4225 (O_4225,N_49157,N_49089);
nor UO_4226 (O_4226,N_49731,N_49451);
nand UO_4227 (O_4227,N_49943,N_49310);
or UO_4228 (O_4228,N_49278,N_49794);
nand UO_4229 (O_4229,N_49095,N_49668);
or UO_4230 (O_4230,N_49395,N_49178);
and UO_4231 (O_4231,N_49804,N_49025);
nor UO_4232 (O_4232,N_49267,N_49555);
and UO_4233 (O_4233,N_49531,N_49462);
and UO_4234 (O_4234,N_49833,N_49252);
or UO_4235 (O_4235,N_49622,N_49624);
nor UO_4236 (O_4236,N_49884,N_49368);
or UO_4237 (O_4237,N_49305,N_49807);
xor UO_4238 (O_4238,N_49107,N_49880);
or UO_4239 (O_4239,N_49720,N_49105);
nor UO_4240 (O_4240,N_49600,N_49277);
nand UO_4241 (O_4241,N_49636,N_49475);
nand UO_4242 (O_4242,N_49511,N_49393);
nor UO_4243 (O_4243,N_49093,N_49173);
and UO_4244 (O_4244,N_49560,N_49699);
or UO_4245 (O_4245,N_49316,N_49893);
nand UO_4246 (O_4246,N_49776,N_49522);
nor UO_4247 (O_4247,N_49577,N_49105);
and UO_4248 (O_4248,N_49750,N_49509);
or UO_4249 (O_4249,N_49869,N_49319);
nand UO_4250 (O_4250,N_49703,N_49041);
xor UO_4251 (O_4251,N_49038,N_49791);
or UO_4252 (O_4252,N_49234,N_49416);
or UO_4253 (O_4253,N_49184,N_49397);
xnor UO_4254 (O_4254,N_49877,N_49299);
or UO_4255 (O_4255,N_49296,N_49065);
and UO_4256 (O_4256,N_49532,N_49123);
nand UO_4257 (O_4257,N_49906,N_49097);
xor UO_4258 (O_4258,N_49482,N_49502);
nand UO_4259 (O_4259,N_49585,N_49068);
nor UO_4260 (O_4260,N_49969,N_49439);
or UO_4261 (O_4261,N_49537,N_49209);
nor UO_4262 (O_4262,N_49918,N_49309);
nor UO_4263 (O_4263,N_49545,N_49957);
nand UO_4264 (O_4264,N_49011,N_49095);
nand UO_4265 (O_4265,N_49746,N_49483);
xnor UO_4266 (O_4266,N_49909,N_49303);
nor UO_4267 (O_4267,N_49373,N_49115);
and UO_4268 (O_4268,N_49358,N_49922);
or UO_4269 (O_4269,N_49068,N_49399);
xor UO_4270 (O_4270,N_49995,N_49163);
nand UO_4271 (O_4271,N_49125,N_49817);
or UO_4272 (O_4272,N_49405,N_49657);
and UO_4273 (O_4273,N_49478,N_49899);
or UO_4274 (O_4274,N_49482,N_49887);
xnor UO_4275 (O_4275,N_49919,N_49147);
xor UO_4276 (O_4276,N_49421,N_49361);
and UO_4277 (O_4277,N_49788,N_49768);
and UO_4278 (O_4278,N_49947,N_49222);
nand UO_4279 (O_4279,N_49879,N_49530);
nor UO_4280 (O_4280,N_49922,N_49955);
or UO_4281 (O_4281,N_49812,N_49957);
nor UO_4282 (O_4282,N_49902,N_49355);
xor UO_4283 (O_4283,N_49478,N_49126);
nand UO_4284 (O_4284,N_49556,N_49458);
xnor UO_4285 (O_4285,N_49789,N_49817);
or UO_4286 (O_4286,N_49892,N_49291);
xor UO_4287 (O_4287,N_49476,N_49076);
or UO_4288 (O_4288,N_49484,N_49530);
or UO_4289 (O_4289,N_49168,N_49623);
nor UO_4290 (O_4290,N_49976,N_49182);
or UO_4291 (O_4291,N_49761,N_49344);
or UO_4292 (O_4292,N_49141,N_49587);
nand UO_4293 (O_4293,N_49413,N_49308);
nor UO_4294 (O_4294,N_49917,N_49995);
and UO_4295 (O_4295,N_49190,N_49906);
nor UO_4296 (O_4296,N_49933,N_49745);
and UO_4297 (O_4297,N_49136,N_49113);
nor UO_4298 (O_4298,N_49792,N_49089);
or UO_4299 (O_4299,N_49493,N_49106);
nor UO_4300 (O_4300,N_49513,N_49597);
xor UO_4301 (O_4301,N_49680,N_49169);
xnor UO_4302 (O_4302,N_49392,N_49787);
xor UO_4303 (O_4303,N_49584,N_49571);
nor UO_4304 (O_4304,N_49656,N_49742);
nand UO_4305 (O_4305,N_49654,N_49583);
and UO_4306 (O_4306,N_49761,N_49321);
xnor UO_4307 (O_4307,N_49473,N_49382);
nor UO_4308 (O_4308,N_49756,N_49257);
or UO_4309 (O_4309,N_49554,N_49952);
or UO_4310 (O_4310,N_49454,N_49497);
and UO_4311 (O_4311,N_49725,N_49583);
or UO_4312 (O_4312,N_49731,N_49116);
nor UO_4313 (O_4313,N_49587,N_49291);
nand UO_4314 (O_4314,N_49148,N_49790);
and UO_4315 (O_4315,N_49171,N_49872);
or UO_4316 (O_4316,N_49980,N_49062);
and UO_4317 (O_4317,N_49157,N_49743);
or UO_4318 (O_4318,N_49026,N_49138);
and UO_4319 (O_4319,N_49591,N_49368);
xnor UO_4320 (O_4320,N_49726,N_49488);
or UO_4321 (O_4321,N_49897,N_49927);
nor UO_4322 (O_4322,N_49769,N_49901);
or UO_4323 (O_4323,N_49977,N_49445);
or UO_4324 (O_4324,N_49738,N_49920);
or UO_4325 (O_4325,N_49168,N_49267);
xnor UO_4326 (O_4326,N_49041,N_49655);
or UO_4327 (O_4327,N_49013,N_49642);
nor UO_4328 (O_4328,N_49458,N_49991);
xor UO_4329 (O_4329,N_49731,N_49322);
nand UO_4330 (O_4330,N_49530,N_49308);
or UO_4331 (O_4331,N_49568,N_49062);
or UO_4332 (O_4332,N_49090,N_49813);
xnor UO_4333 (O_4333,N_49728,N_49001);
nand UO_4334 (O_4334,N_49581,N_49180);
xor UO_4335 (O_4335,N_49077,N_49011);
or UO_4336 (O_4336,N_49070,N_49519);
nor UO_4337 (O_4337,N_49241,N_49949);
nor UO_4338 (O_4338,N_49062,N_49131);
nand UO_4339 (O_4339,N_49899,N_49896);
nand UO_4340 (O_4340,N_49331,N_49572);
or UO_4341 (O_4341,N_49534,N_49483);
xnor UO_4342 (O_4342,N_49262,N_49739);
or UO_4343 (O_4343,N_49131,N_49158);
xor UO_4344 (O_4344,N_49755,N_49592);
or UO_4345 (O_4345,N_49506,N_49131);
nand UO_4346 (O_4346,N_49520,N_49347);
nand UO_4347 (O_4347,N_49436,N_49152);
or UO_4348 (O_4348,N_49596,N_49316);
and UO_4349 (O_4349,N_49673,N_49017);
nor UO_4350 (O_4350,N_49278,N_49741);
or UO_4351 (O_4351,N_49495,N_49629);
and UO_4352 (O_4352,N_49947,N_49819);
or UO_4353 (O_4353,N_49449,N_49224);
nand UO_4354 (O_4354,N_49547,N_49208);
nor UO_4355 (O_4355,N_49407,N_49196);
nor UO_4356 (O_4356,N_49419,N_49809);
xor UO_4357 (O_4357,N_49083,N_49838);
and UO_4358 (O_4358,N_49498,N_49784);
xor UO_4359 (O_4359,N_49367,N_49347);
nand UO_4360 (O_4360,N_49569,N_49714);
nor UO_4361 (O_4361,N_49560,N_49107);
xor UO_4362 (O_4362,N_49489,N_49959);
or UO_4363 (O_4363,N_49400,N_49186);
or UO_4364 (O_4364,N_49903,N_49727);
and UO_4365 (O_4365,N_49968,N_49648);
or UO_4366 (O_4366,N_49279,N_49525);
xnor UO_4367 (O_4367,N_49631,N_49348);
and UO_4368 (O_4368,N_49777,N_49804);
xor UO_4369 (O_4369,N_49582,N_49732);
and UO_4370 (O_4370,N_49767,N_49127);
and UO_4371 (O_4371,N_49833,N_49968);
and UO_4372 (O_4372,N_49644,N_49673);
nand UO_4373 (O_4373,N_49571,N_49636);
or UO_4374 (O_4374,N_49692,N_49756);
nor UO_4375 (O_4375,N_49403,N_49499);
nor UO_4376 (O_4376,N_49745,N_49138);
nor UO_4377 (O_4377,N_49497,N_49791);
xnor UO_4378 (O_4378,N_49527,N_49395);
or UO_4379 (O_4379,N_49333,N_49131);
nor UO_4380 (O_4380,N_49243,N_49701);
xnor UO_4381 (O_4381,N_49286,N_49687);
xnor UO_4382 (O_4382,N_49828,N_49876);
nor UO_4383 (O_4383,N_49828,N_49812);
nor UO_4384 (O_4384,N_49511,N_49530);
and UO_4385 (O_4385,N_49278,N_49083);
and UO_4386 (O_4386,N_49188,N_49368);
and UO_4387 (O_4387,N_49124,N_49932);
nand UO_4388 (O_4388,N_49634,N_49129);
nand UO_4389 (O_4389,N_49573,N_49043);
nand UO_4390 (O_4390,N_49415,N_49493);
and UO_4391 (O_4391,N_49654,N_49383);
and UO_4392 (O_4392,N_49195,N_49239);
nand UO_4393 (O_4393,N_49950,N_49011);
and UO_4394 (O_4394,N_49106,N_49779);
nor UO_4395 (O_4395,N_49834,N_49227);
and UO_4396 (O_4396,N_49362,N_49587);
xnor UO_4397 (O_4397,N_49414,N_49223);
nand UO_4398 (O_4398,N_49046,N_49506);
and UO_4399 (O_4399,N_49729,N_49741);
nand UO_4400 (O_4400,N_49015,N_49429);
or UO_4401 (O_4401,N_49449,N_49130);
and UO_4402 (O_4402,N_49448,N_49219);
nand UO_4403 (O_4403,N_49003,N_49389);
nand UO_4404 (O_4404,N_49705,N_49299);
nor UO_4405 (O_4405,N_49377,N_49159);
or UO_4406 (O_4406,N_49876,N_49055);
and UO_4407 (O_4407,N_49064,N_49134);
or UO_4408 (O_4408,N_49963,N_49590);
nor UO_4409 (O_4409,N_49975,N_49847);
nand UO_4410 (O_4410,N_49994,N_49921);
xnor UO_4411 (O_4411,N_49355,N_49447);
nand UO_4412 (O_4412,N_49424,N_49901);
or UO_4413 (O_4413,N_49797,N_49385);
nand UO_4414 (O_4414,N_49379,N_49644);
nor UO_4415 (O_4415,N_49754,N_49957);
nand UO_4416 (O_4416,N_49120,N_49266);
or UO_4417 (O_4417,N_49875,N_49788);
xor UO_4418 (O_4418,N_49495,N_49055);
nor UO_4419 (O_4419,N_49185,N_49914);
xor UO_4420 (O_4420,N_49823,N_49294);
nor UO_4421 (O_4421,N_49945,N_49308);
nand UO_4422 (O_4422,N_49532,N_49662);
nand UO_4423 (O_4423,N_49650,N_49879);
xor UO_4424 (O_4424,N_49576,N_49845);
xnor UO_4425 (O_4425,N_49000,N_49189);
or UO_4426 (O_4426,N_49121,N_49888);
or UO_4427 (O_4427,N_49671,N_49044);
or UO_4428 (O_4428,N_49010,N_49393);
or UO_4429 (O_4429,N_49001,N_49670);
xor UO_4430 (O_4430,N_49743,N_49120);
nor UO_4431 (O_4431,N_49767,N_49611);
or UO_4432 (O_4432,N_49403,N_49990);
nor UO_4433 (O_4433,N_49204,N_49521);
and UO_4434 (O_4434,N_49758,N_49947);
xnor UO_4435 (O_4435,N_49138,N_49644);
nor UO_4436 (O_4436,N_49510,N_49763);
and UO_4437 (O_4437,N_49138,N_49146);
xor UO_4438 (O_4438,N_49189,N_49181);
and UO_4439 (O_4439,N_49360,N_49212);
xor UO_4440 (O_4440,N_49737,N_49319);
and UO_4441 (O_4441,N_49440,N_49806);
nor UO_4442 (O_4442,N_49638,N_49094);
or UO_4443 (O_4443,N_49649,N_49523);
xnor UO_4444 (O_4444,N_49272,N_49553);
or UO_4445 (O_4445,N_49152,N_49006);
xnor UO_4446 (O_4446,N_49671,N_49553);
xor UO_4447 (O_4447,N_49997,N_49956);
xnor UO_4448 (O_4448,N_49927,N_49924);
or UO_4449 (O_4449,N_49646,N_49539);
nor UO_4450 (O_4450,N_49607,N_49693);
xnor UO_4451 (O_4451,N_49417,N_49652);
nand UO_4452 (O_4452,N_49393,N_49368);
or UO_4453 (O_4453,N_49075,N_49972);
xnor UO_4454 (O_4454,N_49202,N_49713);
xnor UO_4455 (O_4455,N_49348,N_49404);
xor UO_4456 (O_4456,N_49518,N_49936);
or UO_4457 (O_4457,N_49699,N_49733);
or UO_4458 (O_4458,N_49970,N_49679);
nor UO_4459 (O_4459,N_49850,N_49248);
nor UO_4460 (O_4460,N_49657,N_49458);
nand UO_4461 (O_4461,N_49563,N_49061);
and UO_4462 (O_4462,N_49610,N_49378);
xor UO_4463 (O_4463,N_49051,N_49916);
or UO_4464 (O_4464,N_49651,N_49734);
nor UO_4465 (O_4465,N_49058,N_49190);
or UO_4466 (O_4466,N_49711,N_49551);
or UO_4467 (O_4467,N_49971,N_49876);
nand UO_4468 (O_4468,N_49980,N_49121);
nand UO_4469 (O_4469,N_49486,N_49161);
xor UO_4470 (O_4470,N_49236,N_49072);
and UO_4471 (O_4471,N_49161,N_49072);
and UO_4472 (O_4472,N_49263,N_49127);
nor UO_4473 (O_4473,N_49004,N_49517);
and UO_4474 (O_4474,N_49992,N_49565);
or UO_4475 (O_4475,N_49645,N_49693);
nand UO_4476 (O_4476,N_49742,N_49821);
nor UO_4477 (O_4477,N_49610,N_49217);
xnor UO_4478 (O_4478,N_49725,N_49990);
or UO_4479 (O_4479,N_49619,N_49163);
or UO_4480 (O_4480,N_49918,N_49664);
xnor UO_4481 (O_4481,N_49009,N_49760);
xnor UO_4482 (O_4482,N_49823,N_49431);
nand UO_4483 (O_4483,N_49147,N_49517);
nand UO_4484 (O_4484,N_49663,N_49014);
nand UO_4485 (O_4485,N_49259,N_49221);
nand UO_4486 (O_4486,N_49438,N_49380);
or UO_4487 (O_4487,N_49637,N_49407);
nand UO_4488 (O_4488,N_49241,N_49592);
and UO_4489 (O_4489,N_49535,N_49188);
nor UO_4490 (O_4490,N_49735,N_49220);
xor UO_4491 (O_4491,N_49743,N_49896);
xnor UO_4492 (O_4492,N_49066,N_49295);
nand UO_4493 (O_4493,N_49264,N_49613);
nand UO_4494 (O_4494,N_49979,N_49571);
and UO_4495 (O_4495,N_49728,N_49052);
and UO_4496 (O_4496,N_49592,N_49461);
xnor UO_4497 (O_4497,N_49936,N_49388);
and UO_4498 (O_4498,N_49681,N_49556);
or UO_4499 (O_4499,N_49386,N_49977);
nand UO_4500 (O_4500,N_49684,N_49495);
nand UO_4501 (O_4501,N_49969,N_49648);
xor UO_4502 (O_4502,N_49431,N_49295);
xnor UO_4503 (O_4503,N_49433,N_49399);
and UO_4504 (O_4504,N_49726,N_49577);
nand UO_4505 (O_4505,N_49719,N_49005);
and UO_4506 (O_4506,N_49392,N_49169);
and UO_4507 (O_4507,N_49102,N_49430);
nor UO_4508 (O_4508,N_49673,N_49040);
or UO_4509 (O_4509,N_49081,N_49373);
and UO_4510 (O_4510,N_49589,N_49377);
nor UO_4511 (O_4511,N_49901,N_49826);
xnor UO_4512 (O_4512,N_49879,N_49653);
or UO_4513 (O_4513,N_49597,N_49562);
xnor UO_4514 (O_4514,N_49422,N_49889);
xnor UO_4515 (O_4515,N_49976,N_49807);
nor UO_4516 (O_4516,N_49386,N_49044);
and UO_4517 (O_4517,N_49635,N_49264);
xnor UO_4518 (O_4518,N_49277,N_49497);
nand UO_4519 (O_4519,N_49625,N_49725);
and UO_4520 (O_4520,N_49248,N_49179);
and UO_4521 (O_4521,N_49759,N_49500);
nor UO_4522 (O_4522,N_49887,N_49977);
nand UO_4523 (O_4523,N_49599,N_49812);
and UO_4524 (O_4524,N_49914,N_49475);
nor UO_4525 (O_4525,N_49449,N_49865);
xnor UO_4526 (O_4526,N_49153,N_49347);
and UO_4527 (O_4527,N_49755,N_49744);
nor UO_4528 (O_4528,N_49590,N_49633);
nor UO_4529 (O_4529,N_49111,N_49798);
and UO_4530 (O_4530,N_49080,N_49848);
nor UO_4531 (O_4531,N_49329,N_49142);
and UO_4532 (O_4532,N_49407,N_49211);
xnor UO_4533 (O_4533,N_49530,N_49076);
or UO_4534 (O_4534,N_49196,N_49172);
nand UO_4535 (O_4535,N_49262,N_49497);
xor UO_4536 (O_4536,N_49929,N_49267);
or UO_4537 (O_4537,N_49815,N_49308);
or UO_4538 (O_4538,N_49554,N_49411);
nand UO_4539 (O_4539,N_49483,N_49220);
xor UO_4540 (O_4540,N_49051,N_49946);
nand UO_4541 (O_4541,N_49886,N_49801);
or UO_4542 (O_4542,N_49947,N_49411);
or UO_4543 (O_4543,N_49671,N_49478);
nand UO_4544 (O_4544,N_49900,N_49608);
nand UO_4545 (O_4545,N_49925,N_49857);
or UO_4546 (O_4546,N_49923,N_49010);
or UO_4547 (O_4547,N_49787,N_49607);
xnor UO_4548 (O_4548,N_49896,N_49306);
xor UO_4549 (O_4549,N_49525,N_49484);
nand UO_4550 (O_4550,N_49998,N_49095);
nand UO_4551 (O_4551,N_49868,N_49808);
nor UO_4552 (O_4552,N_49706,N_49357);
and UO_4553 (O_4553,N_49247,N_49309);
xnor UO_4554 (O_4554,N_49989,N_49940);
nor UO_4555 (O_4555,N_49609,N_49369);
nor UO_4556 (O_4556,N_49912,N_49035);
and UO_4557 (O_4557,N_49954,N_49225);
or UO_4558 (O_4558,N_49078,N_49530);
and UO_4559 (O_4559,N_49055,N_49256);
nor UO_4560 (O_4560,N_49020,N_49294);
xor UO_4561 (O_4561,N_49165,N_49628);
nor UO_4562 (O_4562,N_49637,N_49909);
and UO_4563 (O_4563,N_49792,N_49176);
nand UO_4564 (O_4564,N_49357,N_49674);
and UO_4565 (O_4565,N_49906,N_49831);
nor UO_4566 (O_4566,N_49839,N_49553);
nor UO_4567 (O_4567,N_49896,N_49219);
and UO_4568 (O_4568,N_49145,N_49491);
and UO_4569 (O_4569,N_49037,N_49763);
nor UO_4570 (O_4570,N_49531,N_49075);
or UO_4571 (O_4571,N_49825,N_49998);
nor UO_4572 (O_4572,N_49976,N_49302);
nor UO_4573 (O_4573,N_49157,N_49300);
or UO_4574 (O_4574,N_49774,N_49718);
or UO_4575 (O_4575,N_49624,N_49581);
and UO_4576 (O_4576,N_49988,N_49651);
xor UO_4577 (O_4577,N_49252,N_49620);
nor UO_4578 (O_4578,N_49403,N_49667);
nor UO_4579 (O_4579,N_49468,N_49094);
nand UO_4580 (O_4580,N_49207,N_49258);
and UO_4581 (O_4581,N_49463,N_49205);
nand UO_4582 (O_4582,N_49487,N_49126);
and UO_4583 (O_4583,N_49702,N_49112);
nor UO_4584 (O_4584,N_49370,N_49942);
nor UO_4585 (O_4585,N_49061,N_49104);
and UO_4586 (O_4586,N_49606,N_49889);
or UO_4587 (O_4587,N_49294,N_49812);
nor UO_4588 (O_4588,N_49664,N_49296);
nor UO_4589 (O_4589,N_49130,N_49779);
nand UO_4590 (O_4590,N_49460,N_49779);
nor UO_4591 (O_4591,N_49236,N_49174);
xnor UO_4592 (O_4592,N_49532,N_49145);
or UO_4593 (O_4593,N_49066,N_49615);
or UO_4594 (O_4594,N_49253,N_49263);
xnor UO_4595 (O_4595,N_49866,N_49146);
xor UO_4596 (O_4596,N_49424,N_49133);
nand UO_4597 (O_4597,N_49773,N_49108);
nor UO_4598 (O_4598,N_49021,N_49614);
nand UO_4599 (O_4599,N_49309,N_49155);
or UO_4600 (O_4600,N_49600,N_49833);
or UO_4601 (O_4601,N_49739,N_49818);
and UO_4602 (O_4602,N_49013,N_49993);
xnor UO_4603 (O_4603,N_49504,N_49462);
nand UO_4604 (O_4604,N_49749,N_49017);
and UO_4605 (O_4605,N_49065,N_49782);
or UO_4606 (O_4606,N_49823,N_49446);
xor UO_4607 (O_4607,N_49225,N_49388);
or UO_4608 (O_4608,N_49239,N_49168);
nand UO_4609 (O_4609,N_49900,N_49490);
nand UO_4610 (O_4610,N_49573,N_49230);
and UO_4611 (O_4611,N_49815,N_49916);
nand UO_4612 (O_4612,N_49507,N_49218);
xnor UO_4613 (O_4613,N_49161,N_49256);
nand UO_4614 (O_4614,N_49761,N_49812);
xor UO_4615 (O_4615,N_49365,N_49011);
xnor UO_4616 (O_4616,N_49834,N_49561);
or UO_4617 (O_4617,N_49177,N_49882);
xnor UO_4618 (O_4618,N_49222,N_49168);
and UO_4619 (O_4619,N_49574,N_49471);
xnor UO_4620 (O_4620,N_49128,N_49213);
nor UO_4621 (O_4621,N_49324,N_49930);
nand UO_4622 (O_4622,N_49667,N_49949);
nand UO_4623 (O_4623,N_49517,N_49272);
and UO_4624 (O_4624,N_49138,N_49386);
or UO_4625 (O_4625,N_49445,N_49436);
or UO_4626 (O_4626,N_49079,N_49810);
or UO_4627 (O_4627,N_49567,N_49548);
or UO_4628 (O_4628,N_49276,N_49836);
xnor UO_4629 (O_4629,N_49208,N_49930);
nand UO_4630 (O_4630,N_49796,N_49470);
nor UO_4631 (O_4631,N_49598,N_49816);
and UO_4632 (O_4632,N_49156,N_49233);
and UO_4633 (O_4633,N_49480,N_49107);
nand UO_4634 (O_4634,N_49882,N_49174);
or UO_4635 (O_4635,N_49801,N_49671);
and UO_4636 (O_4636,N_49109,N_49456);
xnor UO_4637 (O_4637,N_49134,N_49486);
nand UO_4638 (O_4638,N_49963,N_49543);
nor UO_4639 (O_4639,N_49612,N_49595);
or UO_4640 (O_4640,N_49871,N_49804);
and UO_4641 (O_4641,N_49183,N_49134);
nor UO_4642 (O_4642,N_49297,N_49108);
or UO_4643 (O_4643,N_49542,N_49584);
and UO_4644 (O_4644,N_49834,N_49963);
nand UO_4645 (O_4645,N_49810,N_49156);
or UO_4646 (O_4646,N_49158,N_49855);
or UO_4647 (O_4647,N_49270,N_49998);
or UO_4648 (O_4648,N_49472,N_49891);
and UO_4649 (O_4649,N_49754,N_49824);
nor UO_4650 (O_4650,N_49430,N_49826);
or UO_4651 (O_4651,N_49935,N_49108);
nor UO_4652 (O_4652,N_49112,N_49115);
or UO_4653 (O_4653,N_49554,N_49507);
nor UO_4654 (O_4654,N_49874,N_49236);
nor UO_4655 (O_4655,N_49949,N_49749);
nand UO_4656 (O_4656,N_49431,N_49089);
nand UO_4657 (O_4657,N_49132,N_49206);
nand UO_4658 (O_4658,N_49654,N_49891);
xor UO_4659 (O_4659,N_49886,N_49697);
nand UO_4660 (O_4660,N_49767,N_49737);
nand UO_4661 (O_4661,N_49788,N_49835);
and UO_4662 (O_4662,N_49915,N_49660);
nor UO_4663 (O_4663,N_49456,N_49418);
and UO_4664 (O_4664,N_49296,N_49243);
and UO_4665 (O_4665,N_49005,N_49651);
nand UO_4666 (O_4666,N_49235,N_49800);
xor UO_4667 (O_4667,N_49852,N_49670);
or UO_4668 (O_4668,N_49352,N_49866);
and UO_4669 (O_4669,N_49622,N_49523);
nand UO_4670 (O_4670,N_49662,N_49765);
or UO_4671 (O_4671,N_49758,N_49043);
nor UO_4672 (O_4672,N_49319,N_49760);
nand UO_4673 (O_4673,N_49981,N_49901);
nand UO_4674 (O_4674,N_49951,N_49145);
nor UO_4675 (O_4675,N_49656,N_49683);
nor UO_4676 (O_4676,N_49427,N_49584);
and UO_4677 (O_4677,N_49427,N_49098);
and UO_4678 (O_4678,N_49632,N_49679);
xor UO_4679 (O_4679,N_49342,N_49170);
nor UO_4680 (O_4680,N_49070,N_49614);
nand UO_4681 (O_4681,N_49054,N_49203);
xor UO_4682 (O_4682,N_49594,N_49816);
xnor UO_4683 (O_4683,N_49897,N_49712);
xnor UO_4684 (O_4684,N_49629,N_49204);
and UO_4685 (O_4685,N_49006,N_49692);
nor UO_4686 (O_4686,N_49774,N_49338);
nor UO_4687 (O_4687,N_49610,N_49160);
xnor UO_4688 (O_4688,N_49306,N_49726);
nor UO_4689 (O_4689,N_49075,N_49959);
xnor UO_4690 (O_4690,N_49283,N_49017);
xor UO_4691 (O_4691,N_49498,N_49320);
nand UO_4692 (O_4692,N_49741,N_49754);
xor UO_4693 (O_4693,N_49767,N_49583);
nand UO_4694 (O_4694,N_49932,N_49702);
nand UO_4695 (O_4695,N_49673,N_49936);
nor UO_4696 (O_4696,N_49214,N_49334);
or UO_4697 (O_4697,N_49461,N_49876);
nand UO_4698 (O_4698,N_49076,N_49738);
nor UO_4699 (O_4699,N_49374,N_49566);
nand UO_4700 (O_4700,N_49086,N_49420);
and UO_4701 (O_4701,N_49504,N_49804);
xor UO_4702 (O_4702,N_49334,N_49402);
nor UO_4703 (O_4703,N_49097,N_49260);
xnor UO_4704 (O_4704,N_49833,N_49042);
xnor UO_4705 (O_4705,N_49277,N_49987);
nand UO_4706 (O_4706,N_49088,N_49776);
xor UO_4707 (O_4707,N_49119,N_49902);
and UO_4708 (O_4708,N_49595,N_49871);
nor UO_4709 (O_4709,N_49173,N_49301);
and UO_4710 (O_4710,N_49836,N_49102);
nor UO_4711 (O_4711,N_49404,N_49940);
or UO_4712 (O_4712,N_49953,N_49013);
nor UO_4713 (O_4713,N_49917,N_49358);
xor UO_4714 (O_4714,N_49989,N_49943);
nand UO_4715 (O_4715,N_49083,N_49405);
nand UO_4716 (O_4716,N_49357,N_49163);
xnor UO_4717 (O_4717,N_49325,N_49854);
nand UO_4718 (O_4718,N_49423,N_49014);
and UO_4719 (O_4719,N_49233,N_49940);
or UO_4720 (O_4720,N_49553,N_49487);
nand UO_4721 (O_4721,N_49184,N_49779);
nor UO_4722 (O_4722,N_49549,N_49646);
nand UO_4723 (O_4723,N_49275,N_49163);
nand UO_4724 (O_4724,N_49385,N_49270);
or UO_4725 (O_4725,N_49444,N_49167);
nor UO_4726 (O_4726,N_49427,N_49400);
nor UO_4727 (O_4727,N_49735,N_49918);
xor UO_4728 (O_4728,N_49092,N_49859);
nor UO_4729 (O_4729,N_49897,N_49848);
nor UO_4730 (O_4730,N_49794,N_49014);
xnor UO_4731 (O_4731,N_49746,N_49929);
nor UO_4732 (O_4732,N_49994,N_49309);
nor UO_4733 (O_4733,N_49382,N_49540);
and UO_4734 (O_4734,N_49109,N_49826);
or UO_4735 (O_4735,N_49875,N_49619);
and UO_4736 (O_4736,N_49315,N_49269);
and UO_4737 (O_4737,N_49147,N_49663);
or UO_4738 (O_4738,N_49950,N_49917);
and UO_4739 (O_4739,N_49998,N_49738);
nand UO_4740 (O_4740,N_49067,N_49052);
nand UO_4741 (O_4741,N_49133,N_49732);
nand UO_4742 (O_4742,N_49247,N_49592);
or UO_4743 (O_4743,N_49983,N_49782);
xor UO_4744 (O_4744,N_49208,N_49269);
xor UO_4745 (O_4745,N_49966,N_49666);
or UO_4746 (O_4746,N_49362,N_49156);
nor UO_4747 (O_4747,N_49213,N_49137);
or UO_4748 (O_4748,N_49395,N_49373);
nor UO_4749 (O_4749,N_49608,N_49059);
and UO_4750 (O_4750,N_49463,N_49281);
xor UO_4751 (O_4751,N_49401,N_49751);
nand UO_4752 (O_4752,N_49846,N_49983);
nor UO_4753 (O_4753,N_49492,N_49408);
and UO_4754 (O_4754,N_49914,N_49890);
xnor UO_4755 (O_4755,N_49203,N_49439);
and UO_4756 (O_4756,N_49538,N_49913);
nand UO_4757 (O_4757,N_49242,N_49530);
nor UO_4758 (O_4758,N_49589,N_49724);
or UO_4759 (O_4759,N_49737,N_49277);
nand UO_4760 (O_4760,N_49950,N_49717);
xor UO_4761 (O_4761,N_49131,N_49484);
nand UO_4762 (O_4762,N_49925,N_49490);
xnor UO_4763 (O_4763,N_49919,N_49654);
and UO_4764 (O_4764,N_49812,N_49321);
nand UO_4765 (O_4765,N_49354,N_49841);
nand UO_4766 (O_4766,N_49770,N_49022);
or UO_4767 (O_4767,N_49131,N_49713);
nand UO_4768 (O_4768,N_49480,N_49871);
xor UO_4769 (O_4769,N_49338,N_49695);
xnor UO_4770 (O_4770,N_49941,N_49898);
or UO_4771 (O_4771,N_49674,N_49389);
xor UO_4772 (O_4772,N_49590,N_49723);
or UO_4773 (O_4773,N_49239,N_49201);
xor UO_4774 (O_4774,N_49979,N_49192);
nand UO_4775 (O_4775,N_49792,N_49242);
and UO_4776 (O_4776,N_49576,N_49044);
nand UO_4777 (O_4777,N_49254,N_49867);
nand UO_4778 (O_4778,N_49698,N_49666);
and UO_4779 (O_4779,N_49220,N_49973);
xnor UO_4780 (O_4780,N_49212,N_49457);
xnor UO_4781 (O_4781,N_49508,N_49059);
and UO_4782 (O_4782,N_49897,N_49862);
nor UO_4783 (O_4783,N_49099,N_49662);
nand UO_4784 (O_4784,N_49664,N_49019);
xnor UO_4785 (O_4785,N_49723,N_49503);
nor UO_4786 (O_4786,N_49312,N_49423);
xnor UO_4787 (O_4787,N_49607,N_49284);
or UO_4788 (O_4788,N_49068,N_49939);
or UO_4789 (O_4789,N_49130,N_49031);
and UO_4790 (O_4790,N_49191,N_49815);
nor UO_4791 (O_4791,N_49924,N_49688);
xor UO_4792 (O_4792,N_49987,N_49611);
nand UO_4793 (O_4793,N_49124,N_49816);
or UO_4794 (O_4794,N_49164,N_49679);
and UO_4795 (O_4795,N_49733,N_49956);
xnor UO_4796 (O_4796,N_49833,N_49666);
and UO_4797 (O_4797,N_49729,N_49728);
or UO_4798 (O_4798,N_49024,N_49454);
xor UO_4799 (O_4799,N_49144,N_49184);
or UO_4800 (O_4800,N_49227,N_49915);
and UO_4801 (O_4801,N_49327,N_49415);
and UO_4802 (O_4802,N_49154,N_49307);
xnor UO_4803 (O_4803,N_49131,N_49497);
or UO_4804 (O_4804,N_49017,N_49937);
nand UO_4805 (O_4805,N_49365,N_49008);
or UO_4806 (O_4806,N_49841,N_49595);
nand UO_4807 (O_4807,N_49034,N_49788);
nand UO_4808 (O_4808,N_49645,N_49169);
and UO_4809 (O_4809,N_49004,N_49625);
and UO_4810 (O_4810,N_49847,N_49773);
or UO_4811 (O_4811,N_49214,N_49467);
xor UO_4812 (O_4812,N_49914,N_49716);
xnor UO_4813 (O_4813,N_49190,N_49502);
or UO_4814 (O_4814,N_49611,N_49364);
or UO_4815 (O_4815,N_49315,N_49284);
nor UO_4816 (O_4816,N_49348,N_49963);
or UO_4817 (O_4817,N_49363,N_49505);
xnor UO_4818 (O_4818,N_49922,N_49281);
or UO_4819 (O_4819,N_49366,N_49024);
nand UO_4820 (O_4820,N_49330,N_49467);
or UO_4821 (O_4821,N_49050,N_49909);
or UO_4822 (O_4822,N_49356,N_49651);
xnor UO_4823 (O_4823,N_49199,N_49811);
or UO_4824 (O_4824,N_49725,N_49241);
or UO_4825 (O_4825,N_49546,N_49893);
xnor UO_4826 (O_4826,N_49435,N_49981);
nor UO_4827 (O_4827,N_49813,N_49711);
nor UO_4828 (O_4828,N_49635,N_49301);
nor UO_4829 (O_4829,N_49839,N_49656);
nor UO_4830 (O_4830,N_49754,N_49861);
nand UO_4831 (O_4831,N_49647,N_49449);
and UO_4832 (O_4832,N_49044,N_49369);
xnor UO_4833 (O_4833,N_49731,N_49084);
xnor UO_4834 (O_4834,N_49748,N_49251);
xor UO_4835 (O_4835,N_49817,N_49066);
nor UO_4836 (O_4836,N_49852,N_49570);
xnor UO_4837 (O_4837,N_49631,N_49519);
nor UO_4838 (O_4838,N_49171,N_49227);
xnor UO_4839 (O_4839,N_49116,N_49598);
nand UO_4840 (O_4840,N_49196,N_49038);
and UO_4841 (O_4841,N_49553,N_49757);
nor UO_4842 (O_4842,N_49098,N_49807);
nand UO_4843 (O_4843,N_49094,N_49795);
nand UO_4844 (O_4844,N_49437,N_49816);
or UO_4845 (O_4845,N_49285,N_49980);
or UO_4846 (O_4846,N_49060,N_49184);
nand UO_4847 (O_4847,N_49528,N_49593);
and UO_4848 (O_4848,N_49434,N_49054);
and UO_4849 (O_4849,N_49714,N_49033);
nand UO_4850 (O_4850,N_49021,N_49371);
nand UO_4851 (O_4851,N_49898,N_49412);
or UO_4852 (O_4852,N_49068,N_49061);
and UO_4853 (O_4853,N_49265,N_49143);
or UO_4854 (O_4854,N_49965,N_49437);
xnor UO_4855 (O_4855,N_49456,N_49000);
xor UO_4856 (O_4856,N_49721,N_49746);
xor UO_4857 (O_4857,N_49203,N_49127);
and UO_4858 (O_4858,N_49031,N_49524);
xor UO_4859 (O_4859,N_49812,N_49434);
nand UO_4860 (O_4860,N_49603,N_49735);
or UO_4861 (O_4861,N_49756,N_49731);
nor UO_4862 (O_4862,N_49657,N_49012);
nor UO_4863 (O_4863,N_49270,N_49159);
xor UO_4864 (O_4864,N_49423,N_49280);
and UO_4865 (O_4865,N_49314,N_49701);
nor UO_4866 (O_4866,N_49848,N_49835);
nand UO_4867 (O_4867,N_49221,N_49741);
nor UO_4868 (O_4868,N_49121,N_49371);
nand UO_4869 (O_4869,N_49708,N_49555);
nor UO_4870 (O_4870,N_49306,N_49833);
nand UO_4871 (O_4871,N_49119,N_49093);
and UO_4872 (O_4872,N_49446,N_49102);
nor UO_4873 (O_4873,N_49625,N_49074);
nand UO_4874 (O_4874,N_49150,N_49877);
or UO_4875 (O_4875,N_49539,N_49904);
and UO_4876 (O_4876,N_49758,N_49768);
nor UO_4877 (O_4877,N_49561,N_49099);
nand UO_4878 (O_4878,N_49108,N_49766);
xor UO_4879 (O_4879,N_49520,N_49438);
or UO_4880 (O_4880,N_49823,N_49964);
nor UO_4881 (O_4881,N_49748,N_49849);
nor UO_4882 (O_4882,N_49679,N_49475);
xnor UO_4883 (O_4883,N_49659,N_49843);
nor UO_4884 (O_4884,N_49991,N_49905);
nor UO_4885 (O_4885,N_49209,N_49438);
or UO_4886 (O_4886,N_49172,N_49296);
xor UO_4887 (O_4887,N_49851,N_49763);
nand UO_4888 (O_4888,N_49189,N_49528);
xnor UO_4889 (O_4889,N_49395,N_49874);
and UO_4890 (O_4890,N_49416,N_49944);
nand UO_4891 (O_4891,N_49067,N_49421);
xnor UO_4892 (O_4892,N_49090,N_49296);
or UO_4893 (O_4893,N_49428,N_49961);
nor UO_4894 (O_4894,N_49875,N_49300);
nor UO_4895 (O_4895,N_49895,N_49016);
nand UO_4896 (O_4896,N_49315,N_49103);
xor UO_4897 (O_4897,N_49123,N_49719);
or UO_4898 (O_4898,N_49985,N_49135);
or UO_4899 (O_4899,N_49122,N_49782);
or UO_4900 (O_4900,N_49710,N_49204);
or UO_4901 (O_4901,N_49690,N_49265);
nand UO_4902 (O_4902,N_49968,N_49638);
and UO_4903 (O_4903,N_49832,N_49628);
nand UO_4904 (O_4904,N_49418,N_49217);
and UO_4905 (O_4905,N_49003,N_49189);
or UO_4906 (O_4906,N_49385,N_49880);
nor UO_4907 (O_4907,N_49172,N_49625);
nand UO_4908 (O_4908,N_49126,N_49501);
nor UO_4909 (O_4909,N_49592,N_49300);
nand UO_4910 (O_4910,N_49061,N_49559);
nand UO_4911 (O_4911,N_49404,N_49692);
nand UO_4912 (O_4912,N_49047,N_49131);
xor UO_4913 (O_4913,N_49413,N_49963);
nor UO_4914 (O_4914,N_49012,N_49830);
and UO_4915 (O_4915,N_49703,N_49502);
xnor UO_4916 (O_4916,N_49756,N_49629);
or UO_4917 (O_4917,N_49030,N_49121);
and UO_4918 (O_4918,N_49175,N_49432);
and UO_4919 (O_4919,N_49599,N_49055);
nor UO_4920 (O_4920,N_49946,N_49612);
or UO_4921 (O_4921,N_49286,N_49341);
xor UO_4922 (O_4922,N_49748,N_49894);
or UO_4923 (O_4923,N_49371,N_49025);
nor UO_4924 (O_4924,N_49500,N_49966);
nor UO_4925 (O_4925,N_49989,N_49945);
and UO_4926 (O_4926,N_49244,N_49203);
xor UO_4927 (O_4927,N_49644,N_49102);
xor UO_4928 (O_4928,N_49148,N_49092);
or UO_4929 (O_4929,N_49190,N_49876);
nand UO_4930 (O_4930,N_49074,N_49222);
xnor UO_4931 (O_4931,N_49067,N_49633);
xor UO_4932 (O_4932,N_49395,N_49003);
xnor UO_4933 (O_4933,N_49206,N_49552);
nor UO_4934 (O_4934,N_49395,N_49135);
or UO_4935 (O_4935,N_49569,N_49582);
xor UO_4936 (O_4936,N_49848,N_49600);
xor UO_4937 (O_4937,N_49579,N_49487);
nor UO_4938 (O_4938,N_49281,N_49881);
and UO_4939 (O_4939,N_49286,N_49251);
nand UO_4940 (O_4940,N_49843,N_49944);
nor UO_4941 (O_4941,N_49476,N_49613);
or UO_4942 (O_4942,N_49717,N_49530);
xor UO_4943 (O_4943,N_49888,N_49855);
nor UO_4944 (O_4944,N_49134,N_49518);
or UO_4945 (O_4945,N_49466,N_49590);
xor UO_4946 (O_4946,N_49475,N_49923);
nor UO_4947 (O_4947,N_49337,N_49468);
and UO_4948 (O_4948,N_49614,N_49908);
nand UO_4949 (O_4949,N_49298,N_49004);
and UO_4950 (O_4950,N_49491,N_49879);
nand UO_4951 (O_4951,N_49916,N_49899);
xor UO_4952 (O_4952,N_49426,N_49964);
and UO_4953 (O_4953,N_49187,N_49256);
or UO_4954 (O_4954,N_49912,N_49615);
and UO_4955 (O_4955,N_49607,N_49856);
or UO_4956 (O_4956,N_49300,N_49842);
xnor UO_4957 (O_4957,N_49495,N_49147);
nor UO_4958 (O_4958,N_49850,N_49937);
and UO_4959 (O_4959,N_49127,N_49052);
and UO_4960 (O_4960,N_49972,N_49586);
or UO_4961 (O_4961,N_49363,N_49591);
and UO_4962 (O_4962,N_49107,N_49388);
or UO_4963 (O_4963,N_49429,N_49686);
xnor UO_4964 (O_4964,N_49694,N_49776);
or UO_4965 (O_4965,N_49655,N_49550);
nor UO_4966 (O_4966,N_49504,N_49043);
nor UO_4967 (O_4967,N_49700,N_49963);
xnor UO_4968 (O_4968,N_49414,N_49472);
or UO_4969 (O_4969,N_49876,N_49722);
nand UO_4970 (O_4970,N_49356,N_49537);
and UO_4971 (O_4971,N_49206,N_49571);
nor UO_4972 (O_4972,N_49118,N_49989);
xnor UO_4973 (O_4973,N_49356,N_49877);
or UO_4974 (O_4974,N_49088,N_49360);
nand UO_4975 (O_4975,N_49486,N_49269);
or UO_4976 (O_4976,N_49529,N_49378);
xor UO_4977 (O_4977,N_49503,N_49126);
xor UO_4978 (O_4978,N_49137,N_49801);
nor UO_4979 (O_4979,N_49520,N_49432);
and UO_4980 (O_4980,N_49122,N_49761);
and UO_4981 (O_4981,N_49469,N_49656);
nor UO_4982 (O_4982,N_49396,N_49203);
or UO_4983 (O_4983,N_49973,N_49288);
nand UO_4984 (O_4984,N_49975,N_49588);
xor UO_4985 (O_4985,N_49014,N_49844);
xnor UO_4986 (O_4986,N_49503,N_49794);
and UO_4987 (O_4987,N_49119,N_49183);
nor UO_4988 (O_4988,N_49338,N_49093);
and UO_4989 (O_4989,N_49135,N_49827);
or UO_4990 (O_4990,N_49111,N_49857);
and UO_4991 (O_4991,N_49788,N_49483);
or UO_4992 (O_4992,N_49697,N_49051);
xor UO_4993 (O_4993,N_49515,N_49894);
nor UO_4994 (O_4994,N_49358,N_49398);
nor UO_4995 (O_4995,N_49325,N_49495);
nor UO_4996 (O_4996,N_49951,N_49194);
or UO_4997 (O_4997,N_49076,N_49870);
or UO_4998 (O_4998,N_49660,N_49358);
or UO_4999 (O_4999,N_49969,N_49387);
endmodule