module basic_2000_20000_2500_25_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1861,In_1575);
and U1 (N_1,In_1703,In_686);
nor U2 (N_2,In_1490,In_1886);
or U3 (N_3,In_1618,In_1151);
or U4 (N_4,In_6,In_587);
nor U5 (N_5,In_821,In_890);
nor U6 (N_6,In_1790,In_981);
and U7 (N_7,In_184,In_1252);
and U8 (N_8,In_125,In_1200);
or U9 (N_9,In_1552,In_538);
nor U10 (N_10,In_1850,In_1075);
or U11 (N_11,In_1817,In_1671);
and U12 (N_12,In_1279,In_168);
and U13 (N_13,In_9,In_1158);
and U14 (N_14,In_1256,In_893);
or U15 (N_15,In_1557,In_1218);
and U16 (N_16,In_760,In_1129);
nand U17 (N_17,In_395,In_1686);
nor U18 (N_18,In_1479,In_471);
and U19 (N_19,In_1138,In_1794);
or U20 (N_20,In_1634,In_959);
xnor U21 (N_21,In_983,In_1410);
or U22 (N_22,In_273,In_1412);
nand U23 (N_23,In_951,In_551);
or U24 (N_24,In_444,In_1620);
and U25 (N_25,In_1989,In_1821);
nor U26 (N_26,In_1317,In_1147);
or U27 (N_27,In_1532,In_1026);
xnor U28 (N_28,In_1155,In_1705);
and U29 (N_29,In_1809,In_1675);
or U30 (N_30,In_371,In_952);
nand U31 (N_31,In_1053,In_1462);
xor U32 (N_32,In_7,In_896);
nor U33 (N_33,In_30,In_1952);
nor U34 (N_34,In_1550,In_1626);
and U35 (N_35,In_369,In_143);
nand U36 (N_36,In_1023,In_1382);
and U37 (N_37,In_1072,In_1760);
and U38 (N_38,In_693,In_1078);
or U39 (N_39,In_100,In_345);
nand U40 (N_40,In_1347,In_1609);
or U41 (N_41,In_401,In_1459);
or U42 (N_42,In_801,In_921);
and U43 (N_43,In_1638,In_436);
or U44 (N_44,In_1879,In_628);
and U45 (N_45,In_1493,In_192);
or U46 (N_46,In_1040,In_1236);
nor U47 (N_47,In_1646,In_1406);
nand U48 (N_48,In_789,In_1987);
nand U49 (N_49,In_1362,In_944);
or U50 (N_50,In_1178,In_35);
nor U51 (N_51,In_846,In_60);
or U52 (N_52,In_229,In_1536);
xor U53 (N_53,In_27,In_8);
nor U54 (N_54,In_1662,In_323);
xnor U55 (N_55,In_1453,In_694);
nand U56 (N_56,In_601,In_1699);
nor U57 (N_57,In_1170,In_1648);
nand U58 (N_58,In_1571,In_493);
nor U59 (N_59,In_1656,In_281);
nor U60 (N_60,In_1525,In_12);
xor U61 (N_61,In_1544,In_439);
nor U62 (N_62,In_1471,In_680);
and U63 (N_63,In_234,In_120);
nand U64 (N_64,In_1628,In_1878);
and U65 (N_65,In_1866,In_1402);
nand U66 (N_66,In_1566,In_230);
or U67 (N_67,In_1707,In_849);
nand U68 (N_68,In_931,In_1497);
nand U69 (N_69,In_726,In_1919);
nor U70 (N_70,In_332,In_909);
nand U71 (N_71,In_1297,In_594);
and U72 (N_72,In_999,In_966);
nand U73 (N_73,In_151,In_1177);
nor U74 (N_74,In_1610,In_520);
and U75 (N_75,In_813,In_1345);
or U76 (N_76,In_1344,In_270);
and U77 (N_77,In_1215,In_1841);
xor U78 (N_78,In_533,In_853);
nor U79 (N_79,In_415,In_465);
or U80 (N_80,In_1237,In_1341);
xor U81 (N_81,In_1086,In_1365);
xor U82 (N_82,In_1813,In_1063);
xor U83 (N_83,In_861,In_366);
and U84 (N_84,In_1833,In_832);
and U85 (N_85,In_1730,In_1804);
nand U86 (N_86,In_441,In_1971);
or U87 (N_87,In_1473,In_309);
nor U88 (N_88,In_827,In_68);
nor U89 (N_89,In_571,In_1499);
xnor U90 (N_90,In_246,In_497);
and U91 (N_91,In_1088,In_241);
and U92 (N_92,In_182,In_550);
xnor U93 (N_93,In_1176,In_1533);
nor U94 (N_94,In_1067,In_796);
nand U95 (N_95,In_1801,In_397);
xnor U96 (N_96,In_505,In_809);
and U97 (N_97,In_808,In_1383);
xnor U98 (N_98,In_166,In_1839);
xor U99 (N_99,In_1269,In_1732);
and U100 (N_100,In_895,In_231);
or U101 (N_101,In_902,In_637);
and U102 (N_102,In_1961,In_202);
nor U103 (N_103,In_1188,In_961);
xor U104 (N_104,In_1857,In_1426);
and U105 (N_105,In_1738,In_1911);
or U106 (N_106,In_36,In_354);
nand U107 (N_107,In_1593,In_287);
nand U108 (N_108,In_1685,In_1980);
or U109 (N_109,In_1585,In_512);
xor U110 (N_110,In_1411,In_263);
and U111 (N_111,In_1918,In_348);
or U112 (N_112,In_560,In_1856);
nor U113 (N_113,In_511,In_1951);
or U114 (N_114,In_266,In_347);
and U115 (N_115,In_1832,In_445);
or U116 (N_116,In_606,In_352);
and U117 (N_117,In_984,In_524);
xor U118 (N_118,In_1229,In_1294);
or U119 (N_119,In_559,In_1991);
or U120 (N_120,In_1372,In_150);
nor U121 (N_121,In_1051,In_1554);
or U122 (N_122,In_1842,In_1762);
nand U123 (N_123,In_1826,In_854);
and U124 (N_124,In_492,In_146);
and U125 (N_125,In_1590,In_179);
or U126 (N_126,In_1085,In_109);
nand U127 (N_127,In_1444,In_1767);
and U128 (N_128,In_1069,In_28);
and U129 (N_129,In_1538,In_1549);
or U130 (N_130,In_1454,In_1189);
nand U131 (N_131,In_357,In_1670);
nor U132 (N_132,In_19,In_1744);
nand U133 (N_133,In_887,In_1340);
xor U134 (N_134,In_80,In_1999);
or U135 (N_135,In_1579,In_632);
nor U136 (N_136,In_1859,In_545);
nor U137 (N_137,In_1400,In_189);
or U138 (N_138,In_90,In_1522);
or U139 (N_139,In_1721,In_647);
nand U140 (N_140,In_1715,In_1277);
and U141 (N_141,In_841,In_1969);
xor U142 (N_142,In_148,In_40);
and U143 (N_143,In_769,In_1587);
xnor U144 (N_144,In_312,In_670);
xnor U145 (N_145,In_763,In_479);
or U146 (N_146,In_617,In_719);
and U147 (N_147,In_448,In_1672);
nand U148 (N_148,In_1811,In_1131);
xor U149 (N_149,In_1925,In_768);
or U150 (N_150,In_1258,In_64);
or U151 (N_151,In_1021,In_1239);
xnor U152 (N_152,In_424,In_1097);
xor U153 (N_153,In_736,In_1786);
nor U154 (N_154,In_1759,In_970);
nor U155 (N_155,In_1581,In_703);
nor U156 (N_156,In_1805,In_502);
nor U157 (N_157,In_1301,In_836);
or U158 (N_158,In_254,In_1436);
xnor U159 (N_159,In_1933,In_1386);
xnor U160 (N_160,In_1642,In_1348);
or U161 (N_161,In_379,In_1379);
nor U162 (N_162,In_1116,In_177);
xor U163 (N_163,In_29,In_1184);
nor U164 (N_164,In_842,In_1289);
or U165 (N_165,In_522,In_679);
nand U166 (N_166,In_1776,In_925);
xor U167 (N_167,In_111,In_888);
xor U168 (N_168,In_1843,In_905);
nor U169 (N_169,In_1880,In_222);
nor U170 (N_170,In_1824,In_1173);
or U171 (N_171,In_765,In_593);
nand U172 (N_172,In_462,In_857);
xor U173 (N_173,In_1114,In_33);
nor U174 (N_174,In_1146,In_1064);
and U175 (N_175,In_728,In_1797);
nand U176 (N_176,In_1384,In_1673);
xor U177 (N_177,In_420,In_1862);
xor U178 (N_178,In_116,In_1113);
xor U179 (N_179,In_1038,In_608);
nor U180 (N_180,In_58,In_1746);
or U181 (N_181,In_558,In_1443);
xnor U182 (N_182,In_1576,In_130);
or U183 (N_183,In_47,In_882);
nor U184 (N_184,In_958,In_1773);
or U185 (N_185,In_1992,In_531);
and U186 (N_186,In_1586,In_1003);
or U187 (N_187,In_1710,In_877);
nand U188 (N_188,In_541,In_1244);
or U189 (N_189,In_567,In_1562);
nor U190 (N_190,In_1927,In_1511);
xnor U191 (N_191,In_71,In_1932);
or U192 (N_192,In_859,In_1181);
xor U193 (N_193,In_862,In_1713);
or U194 (N_194,In_1605,In_486);
nand U195 (N_195,In_1357,In_1165);
or U196 (N_196,In_1083,In_132);
nor U197 (N_197,In_1442,In_1748);
nor U198 (N_198,In_427,In_1104);
and U199 (N_199,In_387,In_1488);
and U200 (N_200,In_734,In_26);
nand U201 (N_201,In_1986,In_1392);
nor U202 (N_202,In_211,In_1601);
and U203 (N_203,In_405,In_432);
or U204 (N_204,In_76,In_1346);
nand U205 (N_205,In_20,In_139);
xnor U206 (N_206,In_880,In_307);
and U207 (N_207,In_1908,In_1280);
and U208 (N_208,In_1690,In_1355);
nand U209 (N_209,In_1988,In_1098);
nand U210 (N_210,In_1774,In_1700);
and U211 (N_211,In_217,In_1015);
nor U212 (N_212,In_55,In_1894);
nand U213 (N_213,In_583,In_363);
and U214 (N_214,In_1506,In_1373);
nor U215 (N_215,In_1860,In_554);
or U216 (N_216,In_1953,In_786);
nand U217 (N_217,In_1926,In_1807);
xnor U218 (N_218,In_1564,In_816);
nand U219 (N_219,In_1095,In_899);
xnor U220 (N_220,In_1413,In_1186);
nor U221 (N_221,In_1339,In_536);
and U222 (N_222,In_1045,In_322);
or U223 (N_223,In_106,In_337);
nand U224 (N_224,In_965,In_659);
and U225 (N_225,In_592,In_712);
and U226 (N_226,In_1769,In_1134);
nor U227 (N_227,In_602,In_1726);
and U228 (N_228,In_262,In_1046);
xnor U229 (N_229,In_579,In_1283);
or U230 (N_230,In_1791,In_1990);
or U231 (N_231,In_1474,In_500);
xnor U232 (N_232,In_1655,In_223);
and U233 (N_233,In_57,In_691);
and U234 (N_234,In_982,In_1888);
and U235 (N_235,In_1515,In_955);
xnor U236 (N_236,In_1460,In_510);
and U237 (N_237,In_1820,In_800);
nor U238 (N_238,In_919,In_1121);
nand U239 (N_239,In_1127,In_1500);
xnor U240 (N_240,In_581,In_1834);
nand U241 (N_241,In_1541,In_1304);
xnor U242 (N_242,In_1977,In_1111);
nor U243 (N_243,In_741,In_922);
xnor U244 (N_244,In_1916,In_985);
or U245 (N_245,In_742,In_580);
nor U246 (N_246,In_1900,In_450);
and U247 (N_247,In_360,In_1882);
xnor U248 (N_248,In_928,In_1041);
nor U249 (N_249,In_45,In_286);
nor U250 (N_250,In_936,In_1540);
and U251 (N_251,In_1145,In_577);
xor U252 (N_252,In_1750,In_1378);
nor U253 (N_253,In_1440,In_1260);
nand U254 (N_254,In_1368,In_240);
nand U255 (N_255,In_875,In_1309);
and U256 (N_256,In_960,In_710);
xor U257 (N_257,In_306,In_152);
xor U258 (N_258,In_1066,In_381);
xnor U259 (N_259,In_41,In_328);
or U260 (N_260,In_1679,In_613);
or U261 (N_261,In_1315,In_1293);
xor U262 (N_262,In_783,In_390);
or U263 (N_263,In_1125,In_947);
and U264 (N_264,In_1812,In_288);
nor U265 (N_265,In_1955,In_1463);
or U266 (N_266,In_1795,In_34);
and U267 (N_267,In_764,In_137);
xnor U268 (N_268,In_1616,In_95);
xnor U269 (N_269,In_514,In_1005);
nand U270 (N_270,In_1316,In_94);
or U271 (N_271,In_488,In_1603);
or U272 (N_272,In_320,In_1221);
and U273 (N_273,In_1354,In_761);
or U274 (N_274,In_225,In_1204);
or U275 (N_275,In_259,In_1207);
and U276 (N_276,In_651,In_249);
nor U277 (N_277,In_1028,In_353);
nor U278 (N_278,In_1580,In_1160);
xor U279 (N_279,In_785,In_1338);
xnor U280 (N_280,In_738,In_1464);
nand U281 (N_281,In_23,In_663);
and U282 (N_282,In_256,In_639);
or U283 (N_283,In_16,In_1012);
nand U284 (N_284,In_784,In_169);
nand U285 (N_285,In_1337,In_1222);
nor U286 (N_286,In_1684,In_667);
or U287 (N_287,In_812,In_1037);
nand U288 (N_288,In_410,In_452);
nand U289 (N_289,In_186,In_634);
xor U290 (N_290,In_1321,In_790);
and U291 (N_291,In_1192,In_355);
and U292 (N_292,In_671,In_546);
and U293 (N_293,In_375,In_1565);
xnor U294 (N_294,In_1892,In_992);
and U295 (N_295,In_469,In_25);
nor U296 (N_296,In_1897,In_1240);
nor U297 (N_297,In_731,In_1496);
nand U298 (N_298,In_1629,In_1470);
or U299 (N_299,In_838,In_829);
xnor U300 (N_300,In_1367,In_297);
nor U301 (N_301,In_1139,In_279);
nor U302 (N_302,In_508,In_1814);
xnor U303 (N_303,In_1122,In_277);
nor U304 (N_304,In_1042,In_403);
and U305 (N_305,In_190,In_692);
nand U306 (N_306,In_1872,In_336);
nand U307 (N_307,In_119,In_1819);
and U308 (N_308,In_1198,In_478);
and U309 (N_309,In_329,In_1984);
nor U310 (N_310,In_1483,In_1945);
xor U311 (N_311,In_388,In_1263);
xor U312 (N_312,In_14,In_54);
nor U313 (N_313,In_313,In_885);
and U314 (N_314,In_1806,In_860);
and U315 (N_315,In_1491,In_428);
nand U316 (N_316,In_1143,In_1723);
nor U317 (N_317,In_1858,In_1154);
nand U318 (N_318,In_187,In_1388);
or U319 (N_319,In_476,In_743);
or U320 (N_320,In_178,In_62);
nand U321 (N_321,In_1572,In_1545);
nand U322 (N_322,In_1534,In_2);
nor U323 (N_323,In_1976,In_1622);
nand U324 (N_324,In_1696,In_1115);
or U325 (N_325,In_561,In_1692);
nor U326 (N_326,In_117,In_1219);
xor U327 (N_327,In_1030,In_216);
and U328 (N_328,In_1680,In_1725);
nor U329 (N_329,In_721,In_674);
xor U330 (N_330,In_457,In_1663);
xor U331 (N_331,In_1787,In_1307);
nand U332 (N_332,In_614,In_1539);
or U333 (N_333,In_400,In_668);
nor U334 (N_334,In_1895,In_1871);
and U335 (N_335,In_748,In_1494);
nand U336 (N_336,In_707,In_0);
nand U337 (N_337,In_616,In_704);
nor U338 (N_338,In_384,In_1966);
nor U339 (N_339,In_1033,In_830);
nand U340 (N_340,In_1845,In_1006);
nor U341 (N_341,In_737,In_1017);
or U342 (N_342,In_876,In_113);
and U343 (N_343,In_1272,In_525);
and U344 (N_344,In_280,In_472);
nor U345 (N_345,In_455,In_1528);
nor U346 (N_346,In_641,In_310);
nand U347 (N_347,In_386,In_1695);
xnor U348 (N_348,In_688,In_781);
or U349 (N_349,In_562,In_1108);
xor U350 (N_350,In_1889,In_622);
nor U351 (N_351,In_1191,In_101);
and U352 (N_352,In_564,In_1654);
and U353 (N_353,In_1201,In_1978);
xnor U354 (N_354,In_269,In_973);
xnor U355 (N_355,In_891,In_1569);
xnor U356 (N_356,In_1573,In_1822);
and U357 (N_357,In_1251,In_702);
nand U358 (N_358,In_1553,In_200);
nand U359 (N_359,In_1329,In_526);
or U360 (N_360,In_1517,In_814);
xnor U361 (N_361,In_213,In_1687);
xnor U362 (N_362,In_595,In_1153);
or U363 (N_363,In_1310,In_969);
xor U364 (N_364,In_1446,In_53);
nand U365 (N_365,In_1632,In_1298);
xnor U366 (N_366,In_529,In_247);
and U367 (N_367,In_1941,In_547);
nor U368 (N_368,In_1323,In_1942);
nor U369 (N_369,In_250,In_1855);
and U370 (N_370,In_159,In_272);
nand U371 (N_371,In_1107,In_1816);
nand U372 (N_372,In_233,In_1333);
and U373 (N_373,In_1250,In_650);
and U374 (N_374,In_293,In_1351);
and U375 (N_375,In_46,In_276);
nand U376 (N_376,In_507,In_1885);
and U377 (N_377,In_1560,In_1602);
and U378 (N_378,In_1080,In_1688);
and U379 (N_379,In_638,In_1611);
or U380 (N_380,In_126,In_963);
and U381 (N_381,In_1405,In_610);
and U382 (N_382,In_603,In_372);
xor U383 (N_383,In_787,In_1981);
or U384 (N_384,In_170,In_807);
xnor U385 (N_385,In_1034,In_831);
or U386 (N_386,In_343,In_1306);
nor U387 (N_387,In_1391,In_1356);
or U388 (N_388,In_715,In_687);
nand U389 (N_389,In_604,In_833);
or U390 (N_390,In_1935,In_1360);
nand U391 (N_391,In_1947,In_349);
xor U392 (N_392,In_1166,In_308);
or U393 (N_393,In_335,In_624);
and U394 (N_394,In_39,In_156);
xor U395 (N_395,In_443,In_775);
nor U396 (N_396,In_660,In_1657);
xnor U397 (N_397,In_491,In_585);
nand U398 (N_398,In_883,In_1285);
and U399 (N_399,In_160,In_851);
or U400 (N_400,In_1445,In_1011);
or U401 (N_401,In_932,In_459);
xnor U402 (N_402,In_1768,In_1349);
nor U403 (N_403,In_867,In_794);
nor U404 (N_404,In_1708,In_141);
xnor U405 (N_405,In_38,In_93);
or U406 (N_406,In_10,In_1904);
or U407 (N_407,In_1905,In_221);
xnor U408 (N_408,In_723,In_147);
nand U409 (N_409,In_114,In_1543);
nor U410 (N_410,In_1796,In_986);
and U411 (N_411,In_138,In_1253);
or U412 (N_412,In_1979,In_563);
nor U413 (N_413,In_940,In_1148);
xnor U414 (N_414,In_1970,In_1387);
and U415 (N_415,In_154,In_578);
nand U416 (N_416,In_772,In_73);
nand U417 (N_417,In_664,In_1238);
nand U418 (N_418,In_1706,In_174);
nand U419 (N_419,In_1230,In_317);
nor U420 (N_420,In_1577,In_1948);
and U421 (N_421,In_1943,In_1183);
or U422 (N_422,In_753,In_1676);
and U423 (N_423,In_378,In_941);
or U424 (N_424,In_1765,In_1884);
xnor U425 (N_425,In_122,In_805);
nor U426 (N_426,In_980,In_1359);
nand U427 (N_427,In_1044,In_964);
xnor U428 (N_428,In_894,In_88);
and U429 (N_429,In_1752,In_662);
xor U430 (N_430,In_819,In_237);
nand U431 (N_431,In_1245,In_474);
xnor U432 (N_432,In_487,In_1142);
nand U433 (N_433,In_708,In_411);
and U434 (N_434,In_914,In_732);
xor U435 (N_435,In_18,In_66);
or U436 (N_436,In_180,In_584);
nand U437 (N_437,In_1788,In_1002);
xor U438 (N_438,In_1025,In_630);
xnor U439 (N_439,In_950,In_283);
and U440 (N_440,In_815,In_1290);
nor U441 (N_441,In_1082,In_1071);
and U442 (N_442,In_1920,In_1847);
nand U443 (N_443,In_1174,In_724);
xnor U444 (N_444,In_140,In_1852);
nor U445 (N_445,In_1241,In_224);
nor U446 (N_446,In_1950,In_1724);
and U447 (N_447,In_107,In_1612);
and U448 (N_448,In_793,In_540);
nand U449 (N_449,In_82,In_1849);
xor U450 (N_450,In_135,In_705);
and U451 (N_451,In_275,In_615);
and U452 (N_452,In_569,In_588);
or U453 (N_453,In_904,In_1190);
nor U454 (N_454,In_1325,In_1484);
or U455 (N_455,In_1608,In_22);
or U456 (N_456,In_1408,In_417);
or U457 (N_457,In_652,In_1492);
or U458 (N_458,In_866,In_677);
xor U459 (N_459,In_1930,In_195);
or U460 (N_460,In_1836,In_1717);
and U461 (N_461,In_1424,In_70);
nand U462 (N_462,In_239,In_549);
and U463 (N_463,In_466,In_542);
or U464 (N_464,In_3,In_1389);
and U465 (N_465,In_1175,In_431);
or U466 (N_466,In_1284,In_997);
and U467 (N_467,In_1014,In_1658);
nor U468 (N_468,In_191,In_1156);
nand U469 (N_469,In_1764,In_1875);
or U470 (N_470,In_356,In_1419);
nor U471 (N_471,In_1909,In_1777);
or U472 (N_472,In_1427,In_924);
nand U473 (N_473,In_1457,In_1428);
and U474 (N_474,In_1766,In_1783);
or U475 (N_475,In_665,In_1737);
nor U476 (N_476,In_1944,In_1763);
and U477 (N_477,In_52,In_1126);
xor U478 (N_478,In_108,In_1828);
and U479 (N_479,In_1314,In_1659);
or U480 (N_480,In_409,In_1974);
xnor U481 (N_481,In_1110,In_1595);
nand U482 (N_482,In_1194,In_1734);
or U483 (N_483,In_1224,In_494);
nand U484 (N_484,In_1225,In_157);
nand U485 (N_485,In_773,In_611);
nand U486 (N_486,In_797,In_657);
nor U487 (N_487,In_1827,In_1214);
nand U488 (N_488,In_1417,In_566);
nor U489 (N_489,In_1435,In_711);
and U490 (N_490,In_1683,In_817);
nand U491 (N_491,In_1815,In_1024);
nor U492 (N_492,In_1780,In_1397);
and U493 (N_493,In_454,In_302);
or U494 (N_494,In_1718,In_1458);
nor U495 (N_495,In_442,In_1331);
and U496 (N_496,In_1563,In_1906);
nand U497 (N_497,In_757,In_878);
nand U498 (N_498,In_1701,In_518);
nor U499 (N_499,In_1607,In_1267);
nand U500 (N_500,In_1376,In_480);
nor U501 (N_501,In_1010,In_1917);
xnor U502 (N_502,In_599,In_1693);
nor U503 (N_503,In_1433,In_1077);
or U504 (N_504,In_839,In_1936);
or U505 (N_505,In_1374,In_1639);
or U506 (N_506,In_527,In_1132);
or U507 (N_507,In_1048,In_464);
or U508 (N_508,In_218,In_1288);
or U509 (N_509,In_646,In_1519);
xnor U510 (N_510,In_1180,In_321);
nor U511 (N_511,In_72,In_949);
xor U512 (N_512,In_1722,In_1757);
or U513 (N_513,In_1883,In_725);
or U514 (N_514,In_1649,In_1447);
and U515 (N_515,In_1799,In_1669);
xnor U516 (N_516,In_210,In_1150);
xnor U517 (N_517,In_127,In_699);
nor U518 (N_518,In_1123,In_1016);
xor U519 (N_519,In_1808,In_391);
nand U520 (N_520,In_1914,In_1720);
or U521 (N_521,In_1202,In_4);
or U522 (N_522,In_1495,In_456);
or U523 (N_523,In_1223,In_730);
nor U524 (N_524,In_1472,In_700);
nor U525 (N_525,In_557,In_1630);
xnor U526 (N_526,In_1509,In_1516);
nand U527 (N_527,In_252,In_1208);
or U528 (N_528,In_1537,In_1963);
and U529 (N_529,In_110,In_684);
nand U530 (N_530,In_245,In_258);
nand U531 (N_531,In_1101,In_1217);
nand U532 (N_532,In_568,In_373);
or U533 (N_533,In_591,In_1268);
and U534 (N_534,In_235,In_1962);
xor U535 (N_535,In_869,In_1887);
nand U536 (N_536,In_714,In_49);
nor U537 (N_537,In_1964,In_864);
xnor U538 (N_538,In_1414,In_1136);
and U539 (N_539,In_848,In_1729);
and U540 (N_540,In_1060,In_83);
and U541 (N_541,In_1466,In_666);
and U542 (N_542,In_1983,In_449);
nand U543 (N_543,In_1865,In_1247);
xor U544 (N_544,In_1691,In_778);
xnor U545 (N_545,In_1117,In_1130);
nand U546 (N_546,In_318,In_1476);
or U547 (N_547,In_385,In_1869);
nor U548 (N_548,In_1548,In_818);
or U549 (N_549,In_1650,In_574);
or U550 (N_550,In_917,In_1698);
xnor U551 (N_551,In_284,In_621);
nand U552 (N_552,In_1508,In_1782);
nor U553 (N_553,In_382,In_1266);
nor U554 (N_554,In_828,In_257);
nand U555 (N_555,In_1570,In_50);
and U556 (N_556,In_327,In_1084);
or U557 (N_557,In_516,In_1598);
nand U558 (N_558,In_804,In_623);
xnor U559 (N_559,In_1838,In_17);
nor U560 (N_560,In_1281,In_1891);
xor U561 (N_561,In_460,In_75);
xnor U562 (N_562,In_196,In_346);
nor U563 (N_563,In_889,In_291);
or U564 (N_564,In_935,In_1956);
nor U565 (N_565,In_426,In_31);
xor U566 (N_566,In_1312,In_1793);
nor U567 (N_567,In_1418,In_1678);
xnor U568 (N_568,In_121,In_795);
or U569 (N_569,In_1264,In_1489);
nor U570 (N_570,In_1390,In_1430);
and U571 (N_571,In_755,In_521);
or U572 (N_572,In_482,In_331);
nor U573 (N_573,In_771,In_695);
or U574 (N_574,In_1328,In_642);
nand U575 (N_575,In_555,In_244);
xor U576 (N_576,In_1255,In_1985);
nor U577 (N_577,In_1369,In_393);
and U578 (N_578,In_1324,In_453);
or U579 (N_579,In_717,In_265);
or U580 (N_580,In_1363,In_655);
nor U581 (N_581,In_777,In_1651);
or U582 (N_582,In_946,In_1624);
and U583 (N_583,In_1756,In_1334);
xnor U584 (N_584,In_548,In_537);
xor U585 (N_585,In_1404,In_1596);
or U586 (N_586,In_1531,In_433);
and U587 (N_587,In_204,In_653);
and U588 (N_588,In_1800,In_1105);
and U589 (N_589,In_483,In_1332);
xor U590 (N_590,In_458,In_1275);
nor U591 (N_591,In_845,In_988);
nor U592 (N_592,In_1825,In_1873);
and U593 (N_593,In_1246,In_1931);
xor U594 (N_594,In_1530,In_1704);
xnor U595 (N_595,In_682,In_1870);
xor U596 (N_596,In_954,In_627);
xor U597 (N_597,In_1469,In_1232);
nor U598 (N_598,In_1997,In_576);
xnor U599 (N_599,In_501,In_1099);
and U600 (N_600,In_1343,In_1020);
nand U601 (N_601,In_1227,In_1004);
nor U602 (N_602,In_102,In_1381);
nor U603 (N_603,In_435,In_1439);
nand U604 (N_604,In_636,In_1273);
or U605 (N_605,In_1308,In_1637);
xor U606 (N_606,In_1036,In_1965);
nand U607 (N_607,In_798,In_897);
nor U608 (N_608,In_84,In_1396);
xnor U609 (N_609,In_1185,In_43);
xor U610 (N_610,In_163,In_1907);
xnor U611 (N_611,In_774,In_467);
nor U612 (N_612,In_1398,In_85);
and U613 (N_613,In_1226,In_1954);
xor U614 (N_614,In_1582,In_1823);
nand U615 (N_615,In_837,In_333);
xnor U616 (N_616,In_1874,In_945);
nand U617 (N_617,In_1923,In_1631);
nor U618 (N_618,In_468,In_722);
nand U619 (N_619,In_918,In_1877);
and U620 (N_620,In_656,In_1090);
or U621 (N_621,In_1592,In_900);
nor U622 (N_622,In_133,In_1830);
xnor U623 (N_623,In_1450,In_506);
nand U624 (N_624,In_1159,In_530);
nor U625 (N_625,In_1087,In_943);
xnor U626 (N_626,In_1162,In_871);
nand U627 (N_627,In_418,In_1504);
nor U628 (N_628,In_1556,In_1606);
and U629 (N_629,In_1001,In_906);
nand U630 (N_630,In_910,In_1054);
nand U631 (N_631,In_1623,In_609);
and U632 (N_632,In_172,In_776);
nor U633 (N_633,In_1633,In_1199);
nor U634 (N_634,In_131,In_972);
nand U635 (N_635,In_1371,In_1588);
and U636 (N_636,In_1432,In_1124);
nand U637 (N_637,In_1431,In_1102);
or U638 (N_638,In_134,In_251);
xor U639 (N_639,In_412,In_718);
or U640 (N_640,In_207,In_274);
or U641 (N_641,In_413,In_744);
xor U642 (N_642,In_938,In_359);
nand U643 (N_643,In_1061,In_1667);
xnor U644 (N_644,In_625,In_123);
or U645 (N_645,In_112,In_1149);
xor U646 (N_646,In_1228,In_1755);
or U647 (N_647,In_600,In_1336);
xnor U648 (N_648,In_1546,In_1772);
xor U649 (N_649,In_1674,In_463);
nor U650 (N_650,In_1621,In_77);
nor U651 (N_651,In_994,In_1851);
or U652 (N_652,In_1475,In_1320);
and U653 (N_653,In_672,In_69);
and U654 (N_654,In_1257,In_1558);
and U655 (N_655,In_1524,In_1899);
nor U656 (N_656,In_1555,In_619);
xnor U657 (N_657,In_873,In_739);
nand U658 (N_658,In_1278,In_1890);
or U659 (N_659,In_1771,In_908);
and U660 (N_660,In_37,In_698);
xor U661 (N_661,In_1465,In_304);
nor U662 (N_662,In_1599,In_1179);
and U663 (N_663,In_176,In_750);
xor U664 (N_664,In_1578,In_1167);
and U665 (N_665,In_886,In_669);
and U666 (N_666,In_242,In_1056);
xnor U667 (N_667,In_185,In_362);
nand U668 (N_668,In_629,In_389);
nor U669 (N_669,In_929,In_1395);
xor U670 (N_670,In_438,In_572);
nor U671 (N_671,In_1448,In_1993);
or U672 (N_672,In_78,In_1520);
and U673 (N_673,In_844,In_1209);
nand U674 (N_674,In_1144,In_67);
and U675 (N_675,In_1600,In_295);
xor U676 (N_676,In_74,In_879);
nand U677 (N_677,In_175,In_1318);
nor U678 (N_678,In_1503,In_142);
nor U679 (N_679,In_979,In_290);
xor U680 (N_680,In_1665,In_701);
or U681 (N_681,In_1422,In_1135);
nand U682 (N_682,In_1501,In_810);
nand U683 (N_683,In_340,In_1171);
xor U684 (N_684,In_749,In_1625);
xor U685 (N_685,In_1058,In_792);
and U686 (N_686,In_1982,In_490);
nor U687 (N_687,In_1094,In_1287);
nor U688 (N_688,In_1451,In_199);
nand U689 (N_689,In_298,In_597);
nor U690 (N_690,In_998,In_1478);
and U691 (N_691,In_1259,In_1079);
and U692 (N_692,In_746,In_1921);
or U693 (N_693,In_271,In_219);
or U694 (N_694,In_1770,In_1216);
nand U695 (N_695,In_1583,In_1254);
and U696 (N_696,In_872,In_1784);
and U697 (N_697,In_89,In_1584);
nand U698 (N_698,In_1893,In_1589);
and U699 (N_699,In_65,In_1898);
or U700 (N_700,In_1161,In_1480);
nand U701 (N_701,In_377,In_326);
or U702 (N_702,In_1792,In_1689);
xnor U703 (N_703,In_419,In_911);
nand U704 (N_704,In_1393,In_383);
or U705 (N_705,In_425,In_1712);
or U706 (N_706,In_380,In_1749);
xnor U707 (N_707,In_820,In_1643);
nand U708 (N_708,In_1910,In_1802);
nand U709 (N_709,In_953,In_1140);
and U710 (N_710,In_361,In_87);
or U711 (N_711,In_1487,In_865);
or U712 (N_712,In_1975,In_161);
nor U713 (N_713,In_1957,In_214);
xor U714 (N_714,In_1535,In_967);
nand U715 (N_715,In_118,In_181);
xnor U716 (N_716,In_440,In_232);
xor U717 (N_717,In_193,In_752);
nor U718 (N_718,In_1353,In_1653);
and U719 (N_719,In_676,In_1743);
and U720 (N_720,In_1913,In_1291);
and U721 (N_721,In_342,In_1903);
nand U722 (N_722,In_856,In_364);
nor U723 (N_723,In_1152,In_802);
or U724 (N_724,In_912,In_5);
nor U725 (N_725,In_1922,In_1868);
and U726 (N_726,In_556,In_1261);
nand U727 (N_727,In_430,In_689);
nand U728 (N_728,In_408,In_351);
or U729 (N_729,In_626,In_197);
nand U730 (N_730,In_1091,In_1437);
nand U731 (N_731,In_1747,In_292);
and U732 (N_732,In_446,In_1694);
nor U733 (N_733,In_640,In_201);
and U734 (N_734,In_780,In_956);
nand U735 (N_735,In_1853,In_303);
xor U736 (N_736,In_103,In_1840);
or U737 (N_737,In_1081,In_392);
nor U738 (N_738,In_1137,In_79);
nor U739 (N_739,In_1206,In_1785);
nor U740 (N_740,In_834,In_586);
or U741 (N_741,In_683,In_206);
nand U742 (N_742,In_962,In_539);
nor U743 (N_743,In_926,In_1881);
nand U744 (N_744,In_1361,In_1901);
xor U745 (N_745,In_1967,In_835);
xnor U746 (N_746,In_826,In_1709);
nor U747 (N_747,In_1468,In_1120);
or U748 (N_748,In_255,In_582);
nand U749 (N_749,In_164,In_1604);
nor U750 (N_750,In_1529,In_1798);
nor U751 (N_751,In_863,In_729);
and U752 (N_752,In_374,In_1661);
xor U753 (N_753,In_1292,In_1835);
xor U754 (N_754,In_673,In_1299);
nand U755 (N_755,In_1449,In_916);
and U756 (N_756,In_97,In_1375);
xor U757 (N_757,In_1594,In_937);
and U758 (N_758,In_1477,In_1711);
nor U759 (N_759,In_324,In_461);
nor U760 (N_760,In_759,In_1929);
and U761 (N_761,In_1031,In_260);
xor U762 (N_762,In_1635,In_1342);
nor U763 (N_763,In_1296,In_1716);
or U764 (N_764,In_1043,In_341);
nand U765 (N_765,In_733,In_330);
or U766 (N_766,In_898,In_643);
xnor U767 (N_767,In_1322,In_1641);
nor U768 (N_768,In_553,In_1065);
nand U769 (N_769,In_920,In_1093);
or U770 (N_770,In_220,In_1);
nor U771 (N_771,In_316,In_1335);
and U772 (N_772,In_1995,In_523);
xor U773 (N_773,In_86,In_1498);
xnor U774 (N_774,In_987,In_294);
nor U775 (N_775,In_1741,In_1364);
nor U776 (N_776,In_1282,In_188);
and U777 (N_777,In_1867,In_1568);
xor U778 (N_778,In_915,In_1193);
or U779 (N_779,In_503,In_1248);
nand U780 (N_780,In_416,In_1330);
or U781 (N_781,In_756,In_422);
xor U782 (N_782,In_1636,In_1169);
or U783 (N_783,In_870,In_645);
nor U784 (N_784,In_406,In_1262);
and U785 (N_785,In_15,In_365);
and U786 (N_786,In_319,In_565);
and U787 (N_787,In_414,In_1513);
nor U788 (N_788,In_1502,In_791);
nor U789 (N_789,In_824,In_1429);
nor U790 (N_790,In_1103,In_253);
nand U791 (N_791,In_811,In_1481);
and U792 (N_792,In_59,In_1863);
and U793 (N_793,In_1697,In_1810);
and U794 (N_794,In_515,In_99);
xnor U795 (N_795,In_823,In_1682);
nand U796 (N_796,In_1394,In_1265);
xor U797 (N_797,In_1055,In_1203);
nand U798 (N_798,In_1270,In_552);
nor U799 (N_799,In_128,In_261);
and U800 (N_800,N_52,In_1681);
or U801 (N_801,N_197,In_1505);
xnor U802 (N_802,In_939,N_313);
and U803 (N_803,N_70,In_149);
nand U804 (N_804,N_188,N_265);
xnor U805 (N_805,In_762,N_557);
xor U806 (N_806,N_493,In_1164);
nand U807 (N_807,N_650,N_798);
or U808 (N_808,In_368,N_494);
xor U809 (N_809,N_305,In_1702);
or U810 (N_810,N_60,N_225);
or U811 (N_811,N_463,N_440);
nand U812 (N_812,N_107,In_434);
xnor U813 (N_813,In_421,In_1271);
or U814 (N_814,N_680,In_98);
nand U815 (N_815,N_504,N_377);
xor U816 (N_816,N_785,N_284);
or U817 (N_817,N_664,In_1779);
or U818 (N_818,N_474,N_288);
xor U819 (N_819,In_1133,N_111);
or U820 (N_820,N_117,N_148);
and U821 (N_821,N_73,N_215);
xnor U822 (N_822,N_74,N_670);
xnor U823 (N_823,N_607,N_471);
or U824 (N_824,N_737,N_100);
and U825 (N_825,In_104,In_489);
nand U826 (N_826,N_676,N_481);
nand U827 (N_827,In_766,In_934);
nand U828 (N_828,N_24,N_280);
xnor U829 (N_829,In_770,N_383);
nand U830 (N_830,N_546,N_71);
nand U831 (N_831,N_310,N_297);
nand U832 (N_832,N_622,N_38);
or U833 (N_833,N_718,N_26);
and U834 (N_834,In_1049,N_139);
or U835 (N_835,In_598,N_793);
nand U836 (N_836,In_913,N_690);
nor U837 (N_837,In_1547,N_562);
xnor U838 (N_838,In_1829,N_610);
and U839 (N_839,N_693,In_1029);
and U840 (N_840,In_311,N_534);
or U841 (N_841,N_242,N_3);
nor U842 (N_842,N_9,N_287);
xor U843 (N_843,In_32,N_286);
nor U844 (N_844,In_1735,N_113);
or U845 (N_845,N_300,N_437);
and U846 (N_846,N_469,N_395);
or U847 (N_847,In_350,N_406);
and U848 (N_848,N_103,N_449);
nand U849 (N_849,N_775,In_1740);
nand U850 (N_850,N_204,N_203);
or U851 (N_851,In_658,N_116);
nor U852 (N_852,N_397,N_506);
nand U853 (N_853,In_226,N_551);
nor U854 (N_854,N_643,N_23);
xnor U855 (N_855,In_1380,N_735);
nand U856 (N_856,N_296,N_61);
or U857 (N_857,In_1172,N_638);
nand U858 (N_858,In_1854,N_446);
and U859 (N_859,N_704,N_637);
or U860 (N_860,N_387,N_672);
nor U861 (N_861,N_520,In_570);
xnor U862 (N_862,N_80,In_105);
nand U863 (N_863,N_128,N_279);
or U864 (N_864,N_571,In_315);
nor U865 (N_865,In_767,N_669);
or U866 (N_866,N_77,N_753);
or U867 (N_867,In_1486,N_220);
xor U868 (N_868,In_575,N_491);
nand U869 (N_869,In_519,In_1619);
nand U870 (N_870,N_129,In_825);
nand U871 (N_871,N_432,N_6);
and U872 (N_872,In_509,In_716);
and U873 (N_873,In_696,N_336);
or U874 (N_874,In_1666,N_332);
and U875 (N_875,N_325,N_516);
or U876 (N_876,N_114,N_715);
or U877 (N_877,N_316,N_210);
nand U878 (N_878,N_599,In_1100);
nand U879 (N_879,In_1719,In_1303);
nor U880 (N_880,N_264,In_806);
nand U881 (N_881,In_484,N_651);
nand U882 (N_882,In_990,N_528);
xnor U883 (N_883,N_403,In_1022);
nand U884 (N_884,N_307,In_51);
nand U885 (N_885,In_11,N_705);
nand U886 (N_886,N_450,N_88);
nand U887 (N_887,In_358,N_613);
xor U888 (N_888,N_617,In_243);
and U889 (N_889,N_298,N_467);
and U890 (N_890,N_726,N_179);
and U891 (N_891,N_368,N_164);
xor U892 (N_892,N_349,N_512);
or U893 (N_893,N_119,N_55);
and U894 (N_894,N_238,N_631);
nand U895 (N_895,In_923,N_646);
and U896 (N_896,N_40,N_748);
nor U897 (N_897,N_490,In_198);
nand U898 (N_898,In_1818,N_549);
or U899 (N_899,N_470,N_22);
or U900 (N_900,In_850,N_795);
or U901 (N_901,In_1319,N_400);
xnor U902 (N_902,N_369,N_663);
nor U903 (N_903,N_654,N_439);
or U904 (N_904,N_665,N_413);
and U905 (N_905,N_658,N_181);
and U906 (N_906,In_690,N_187);
xor U907 (N_907,In_1597,N_58);
nor U908 (N_908,N_792,N_96);
or U909 (N_909,N_333,N_515);
and U910 (N_910,N_579,In_1902);
xor U911 (N_911,N_683,N_707);
or U912 (N_912,N_206,N_157);
nor U913 (N_913,In_1407,N_177);
xnor U914 (N_914,N_418,N_623);
nor U915 (N_915,In_268,N_405);
xnor U916 (N_916,N_547,N_766);
or U917 (N_917,N_112,N_379);
nor U918 (N_918,In_596,In_404);
nor U919 (N_919,N_681,In_993);
or U920 (N_920,N_410,N_759);
xor U921 (N_921,N_222,In_451);
or U922 (N_922,N_521,N_110);
xor U923 (N_923,N_270,N_480);
nand U924 (N_924,N_322,In_285);
and U925 (N_925,N_248,In_1574);
nand U926 (N_926,N_739,N_442);
and U927 (N_927,N_559,N_271);
nand U928 (N_928,N_125,In_314);
nor U929 (N_929,N_628,N_656);
or U930 (N_930,N_170,In_649);
xor U931 (N_931,In_1467,N_736);
nand U932 (N_932,In_61,N_580);
nor U933 (N_933,N_427,N_302);
nand U934 (N_934,N_621,N_452);
nand U935 (N_935,In_754,N_543);
and U936 (N_936,N_741,In_1482);
xor U937 (N_937,N_374,N_201);
xnor U938 (N_938,N_575,N_538);
or U939 (N_939,In_685,In_1212);
or U940 (N_940,In_173,N_144);
nand U941 (N_941,N_722,N_772);
nand U942 (N_942,N_586,N_78);
xnor U943 (N_943,N_636,N_584);
and U944 (N_944,N_781,In_868);
nor U945 (N_945,In_1295,In_162);
nand U946 (N_946,N_102,In_1118);
nand U947 (N_947,In_971,In_654);
and U948 (N_948,In_532,N_511);
and U949 (N_949,N_412,N_232);
nor U950 (N_950,In_92,In_1736);
and U951 (N_951,In_399,N_535);
xnor U952 (N_952,In_1559,N_694);
and U953 (N_953,N_216,N_200);
nand U954 (N_954,N_142,In_1613);
nor U955 (N_955,N_505,N_193);
nor U956 (N_956,N_283,N_385);
or U957 (N_957,N_10,N_13);
and U958 (N_958,In_858,In_843);
nor U959 (N_959,N_790,N_484);
nor U960 (N_960,N_508,N_751);
xnor U961 (N_961,N_578,N_509);
or U962 (N_962,N_183,In_1062);
or U963 (N_963,In_1311,In_236);
and U964 (N_964,N_253,In_325);
nand U965 (N_965,N_198,N_97);
nand U966 (N_966,N_545,N_268);
nor U967 (N_967,N_237,N_411);
nand U968 (N_968,In_1848,N_353);
and U969 (N_969,In_822,In_1370);
and U970 (N_970,N_421,N_478);
xor U971 (N_971,N_438,In_678);
xor U972 (N_972,N_199,In_1837);
xor U973 (N_973,N_0,N_252);
xnor U974 (N_974,N_338,N_93);
nand U975 (N_975,In_423,N_539);
or U976 (N_976,N_79,In_1731);
and U977 (N_977,N_15,N_640);
nand U978 (N_978,N_419,In_398);
nor U979 (N_979,N_784,In_975);
nor U980 (N_980,In_589,In_499);
xnor U981 (N_981,N_346,N_647);
xor U982 (N_982,N_317,N_563);
nand U983 (N_983,In_544,N_277);
xor U984 (N_984,N_36,N_218);
nand U985 (N_985,In_644,N_12);
xor U986 (N_986,N_574,N_624);
and U987 (N_987,N_655,In_1235);
nor U988 (N_988,N_124,In_1000);
or U989 (N_989,In_24,In_1959);
or U990 (N_990,N_489,N_1);
and U991 (N_991,In_635,N_604);
or U992 (N_992,In_155,In_1327);
nand U993 (N_993,N_76,N_269);
nor U994 (N_994,N_230,N_716);
or U995 (N_995,N_255,N_141);
nand U996 (N_996,N_661,N_314);
or U997 (N_997,In_136,In_1019);
nor U998 (N_998,N_189,In_339);
nand U999 (N_999,N_330,In_927);
xor U1000 (N_1000,N_517,In_158);
nand U1001 (N_1001,In_1213,In_709);
and U1002 (N_1002,In_396,N_389);
nand U1003 (N_1003,N_339,N_703);
or U1004 (N_1004,N_91,N_319);
nand U1005 (N_1005,N_25,N_47);
nand U1006 (N_1006,N_444,N_33);
nor U1007 (N_1007,N_761,In_1455);
or U1008 (N_1008,In_376,N_526);
or U1009 (N_1009,In_194,N_48);
and U1010 (N_1010,N_137,In_1518);
nand U1011 (N_1011,N_644,N_530);
xnor U1012 (N_1012,N_262,N_20);
or U1013 (N_1013,N_371,N_361);
and U1014 (N_1014,In_475,N_57);
and U1015 (N_1015,In_1938,In_300);
nor U1016 (N_1016,N_659,N_660);
xnor U1017 (N_1017,N_696,N_618);
and U1018 (N_1018,N_619,N_35);
nor U1019 (N_1019,N_794,N_8);
nand U1020 (N_1020,N_393,N_261);
nand U1021 (N_1021,In_1243,In_1452);
xor U1022 (N_1022,N_99,In_1994);
xor U1023 (N_1023,In_1242,In_504);
xnor U1024 (N_1024,In_1934,N_104);
nand U1025 (N_1025,In_167,N_717);
nand U1026 (N_1026,N_308,In_513);
xnor U1027 (N_1027,N_367,N_246);
or U1028 (N_1028,In_1416,N_347);
nand U1029 (N_1029,N_692,N_777);
nand U1030 (N_1030,N_689,N_335);
nor U1031 (N_1031,In_989,N_165);
nand U1032 (N_1032,N_49,In_81);
and U1033 (N_1033,In_228,In_727);
xnor U1034 (N_1034,N_64,N_243);
or U1035 (N_1035,N_462,In_607);
and U1036 (N_1036,N_750,In_1423);
and U1037 (N_1037,N_634,N_732);
or U1038 (N_1038,N_351,N_459);
nand U1039 (N_1039,N_495,N_32);
xnor U1040 (N_1040,N_501,N_382);
and U1041 (N_1041,N_344,N_611);
xnor U1042 (N_1042,In_296,N_699);
or U1043 (N_1043,N_518,N_468);
and U1044 (N_1044,N_697,N_274);
nand U1045 (N_1045,In_1233,In_282);
nand U1046 (N_1046,N_106,N_662);
and U1047 (N_1047,N_725,In_933);
xnor U1048 (N_1048,N_453,In_437);
and U1049 (N_1049,N_84,N_227);
nand U1050 (N_1050,In_1514,N_90);
and U1051 (N_1051,N_756,In_1972);
and U1052 (N_1052,In_1420,N_388);
or U1053 (N_1053,N_479,In_1205);
and U1054 (N_1054,N_743,N_194);
nand U1055 (N_1055,In_1168,N_687);
or U1056 (N_1056,N_500,In_264);
xor U1057 (N_1057,N_711,In_205);
nand U1058 (N_1058,N_779,N_391);
nor U1059 (N_1059,In_124,N_649);
nand U1060 (N_1060,N_724,N_115);
nor U1061 (N_1061,In_1210,N_706);
nand U1062 (N_1062,In_407,N_208);
nor U1063 (N_1063,N_475,N_132);
xnor U1064 (N_1064,In_1109,N_303);
or U1065 (N_1065,N_272,N_763);
or U1066 (N_1066,In_1924,N_169);
or U1067 (N_1067,N_83,In_1647);
xnor U1068 (N_1068,N_54,N_552);
or U1069 (N_1069,N_18,In_535);
or U1070 (N_1070,N_529,N_577);
nand U1071 (N_1071,N_376,N_375);
xnor U1072 (N_1072,In_1074,N_561);
nor U1073 (N_1073,N_625,N_256);
nand U1074 (N_1074,N_487,In_1781);
xnor U1075 (N_1075,N_384,N_131);
and U1076 (N_1076,N_50,In_1434);
and U1077 (N_1077,N_629,N_92);
nor U1078 (N_1078,N_101,In_1660);
and U1079 (N_1079,N_714,N_380);
xnor U1080 (N_1080,In_713,N_87);
xnor U1081 (N_1081,N_68,In_1403);
nor U1082 (N_1082,N_686,N_461);
xor U1083 (N_1083,N_457,N_250);
nor U1084 (N_1084,N_642,In_402);
xor U1085 (N_1085,N_677,In_1352);
nor U1086 (N_1086,N_254,N_712);
xor U1087 (N_1087,In_758,N_721);
nand U1088 (N_1088,In_1300,In_1157);
and U1089 (N_1089,N_594,N_458);
nor U1090 (N_1090,N_630,In_1761);
nor U1091 (N_1091,In_706,N_752);
or U1092 (N_1092,N_757,N_331);
or U1093 (N_1093,In_1068,N_455);
nand U1094 (N_1094,N_143,In_1009);
and U1095 (N_1095,N_155,N_257);
xor U1096 (N_1096,N_45,In_44);
nand U1097 (N_1097,N_290,In_840);
or U1098 (N_1098,N_11,N_312);
xor U1099 (N_1099,N_598,N_345);
xnor U1100 (N_1100,N_560,In_1302);
xnor U1101 (N_1101,N_770,N_733);
or U1102 (N_1102,N_596,N_477);
nor U1103 (N_1103,In_976,N_259);
or U1104 (N_1104,In_968,In_1050);
nor U1105 (N_1105,N_229,In_907);
xnor U1106 (N_1106,In_996,In_1527);
nor U1107 (N_1107,N_217,N_558);
xor U1108 (N_1108,N_267,In_720);
and U1109 (N_1109,In_1076,N_791);
or U1110 (N_1110,In_1664,N_778);
xor U1111 (N_1111,N_612,N_565);
nand U1112 (N_1112,N_334,In_267);
nand U1113 (N_1113,In_1112,N_151);
xnor U1114 (N_1114,N_82,N_592);
nand U1115 (N_1115,In_1057,In_590);
and U1116 (N_1116,In_803,N_657);
or U1117 (N_1117,In_367,N_360);
and U1118 (N_1118,N_633,N_632);
nor U1119 (N_1119,In_1211,In_1141);
xor U1120 (N_1120,N_588,N_476);
nand U1121 (N_1121,N_202,N_328);
or U1122 (N_1122,N_460,N_409);
or U1123 (N_1123,N_178,N_240);
and U1124 (N_1124,N_548,N_429);
nor U1125 (N_1125,In_56,In_517);
xnor U1126 (N_1126,In_238,In_534);
or U1127 (N_1127,In_633,N_196);
nand U1128 (N_1128,N_760,N_674);
xnor U1129 (N_1129,N_394,N_441);
or U1130 (N_1130,N_709,N_42);
nand U1131 (N_1131,In_212,In_1274);
and U1132 (N_1132,N_700,N_289);
or U1133 (N_1133,In_1831,N_544);
and U1134 (N_1134,N_524,In_1441);
nor U1135 (N_1135,N_789,N_570);
and U1136 (N_1136,N_466,N_593);
xnor U1137 (N_1137,N_63,N_192);
or U1138 (N_1138,In_1092,In_1803);
xnor U1139 (N_1139,In_930,N_95);
nor U1140 (N_1140,N_498,N_402);
nand U1141 (N_1141,N_454,N_89);
or U1142 (N_1142,N_620,N_483);
nor U1143 (N_1143,In_481,In_1197);
nand U1144 (N_1144,N_684,N_627);
nand U1145 (N_1145,N_456,N_698);
nand U1146 (N_1146,N_329,N_171);
and U1147 (N_1147,N_738,N_597);
xnor U1148 (N_1148,In_1778,N_702);
or U1149 (N_1149,N_352,N_364);
nand U1150 (N_1150,In_1973,In_115);
nand U1151 (N_1151,N_86,N_266);
nor U1152 (N_1152,In_1542,N_315);
and U1153 (N_1153,N_464,N_31);
nor U1154 (N_1154,N_241,N_710);
or U1155 (N_1155,N_85,In_1521);
xor U1156 (N_1156,In_1615,N_430);
nor U1157 (N_1157,N_768,N_341);
or U1158 (N_1158,N_555,N_595);
xor U1159 (N_1159,In_153,N_723);
or U1160 (N_1160,In_884,N_354);
nand U1161 (N_1161,In_745,In_681);
nand U1162 (N_1162,N_731,N_497);
xnor U1163 (N_1163,N_231,In_1409);
nor U1164 (N_1164,N_499,N_235);
nor U1165 (N_1165,N_754,N_425);
or U1166 (N_1166,In_215,In_1939);
or U1167 (N_1167,N_742,N_435);
xor U1168 (N_1168,N_507,N_282);
nor U1169 (N_1169,In_248,In_1591);
or U1170 (N_1170,N_214,N_109);
nand U1171 (N_1171,N_140,N_416);
xnor U1172 (N_1172,In_1089,In_1996);
nand U1173 (N_1173,In_995,N_744);
xor U1174 (N_1174,N_569,N_306);
nor U1175 (N_1175,In_1640,N_730);
or U1176 (N_1176,In_874,N_372);
nor U1177 (N_1177,N_496,N_166);
and U1178 (N_1178,N_348,In_1182);
or U1179 (N_1179,In_1751,N_207);
or U1180 (N_1180,N_381,In_496);
nor U1181 (N_1181,In_1614,N_278);
and U1182 (N_1182,In_1896,In_1937);
nand U1183 (N_1183,N_436,N_136);
nor U1184 (N_1184,In_528,In_1128);
and U1185 (N_1185,N_773,N_399);
nor U1186 (N_1186,N_182,N_783);
and U1187 (N_1187,N_488,In_1286);
xnor U1188 (N_1188,N_675,In_370);
xnor U1189 (N_1189,N_75,N_566);
nor U1190 (N_1190,In_661,N_767);
and U1191 (N_1191,N_465,In_1946);
nand U1192 (N_1192,In_1617,N_127);
nand U1193 (N_1193,In_1512,N_244);
and U1194 (N_1194,In_477,N_350);
and U1195 (N_1195,N_108,N_156);
or U1196 (N_1196,N_685,N_734);
nor U1197 (N_1197,N_167,N_398);
and U1198 (N_1198,N_145,N_72);
and U1199 (N_1199,N_249,In_96);
nand U1200 (N_1200,N_98,In_799);
or U1201 (N_1201,N_787,N_679);
nand U1202 (N_1202,N_209,In_751);
nand U1203 (N_1203,N_130,N_219);
xnor U1204 (N_1204,N_682,N_713);
nor U1205 (N_1205,N_163,N_29);
and U1206 (N_1206,N_159,N_276);
nor U1207 (N_1207,N_46,N_424);
nand U1208 (N_1208,In_1627,N_190);
nor U1209 (N_1209,N_28,N_522);
nand U1210 (N_1210,In_1758,N_41);
nor U1211 (N_1211,N_285,N_135);
xnor U1212 (N_1212,N_745,N_447);
or U1213 (N_1213,In_1059,N_531);
nor U1214 (N_1214,N_691,In_892);
xor U1215 (N_1215,In_605,N_396);
and U1216 (N_1216,N_482,N_433);
nand U1217 (N_1217,N_275,N_585);
nand U1218 (N_1218,In_1035,N_688);
or U1219 (N_1219,In_1526,In_1510);
nor U1220 (N_1220,In_855,In_171);
and U1221 (N_1221,N_417,In_1377);
xnor U1222 (N_1222,N_523,In_1399);
nand U1223 (N_1223,In_1915,N_34);
nand U1224 (N_1224,N_324,In_1385);
nor U1225 (N_1225,In_344,N_525);
or U1226 (N_1226,N_451,N_755);
nor U1227 (N_1227,N_363,In_1106);
nand U1228 (N_1228,In_1008,N_609);
xnor U1229 (N_1229,N_527,In_21);
xor U1230 (N_1230,N_582,N_653);
nor U1231 (N_1231,N_581,In_1358);
nand U1232 (N_1232,N_408,N_774);
nand U1233 (N_1233,In_1928,N_386);
nor U1234 (N_1234,In_1039,N_590);
xnor U1235 (N_1235,In_747,In_278);
nor U1236 (N_1236,N_245,N_639);
and U1237 (N_1237,N_666,N_291);
nor U1238 (N_1238,In_1745,In_782);
nand U1239 (N_1239,N_294,N_94);
nand U1240 (N_1240,N_614,N_59);
and U1241 (N_1241,N_21,N_573);
or U1242 (N_1242,N_236,N_600);
nand U1243 (N_1243,N_161,N_556);
and U1244 (N_1244,In_1645,In_903);
xor U1245 (N_1245,In_1775,N_514);
nand U1246 (N_1246,N_186,N_564);
or U1247 (N_1247,N_486,In_1421);
nand U1248 (N_1248,In_447,N_281);
xor U1249 (N_1249,In_13,N_414);
and U1250 (N_1250,N_485,N_251);
nor U1251 (N_1251,In_1234,N_320);
nand U1252 (N_1252,N_769,N_519);
and U1253 (N_1253,In_299,N_572);
and U1254 (N_1254,N_635,N_138);
nand U1255 (N_1255,In_543,N_7);
nand U1256 (N_1256,N_796,In_1960);
nor U1257 (N_1257,In_1940,N_152);
and U1258 (N_1258,N_295,In_612);
and U1259 (N_1259,In_1507,N_671);
nand U1260 (N_1260,N_4,N_431);
xnor U1261 (N_1261,N_606,In_63);
xor U1262 (N_1262,In_618,N_765);
or U1263 (N_1263,N_780,N_358);
xnor U1264 (N_1264,N_583,N_788);
nand U1265 (N_1265,In_1864,In_470);
xnor U1266 (N_1266,N_589,In_1119);
or U1267 (N_1267,N_536,N_727);
nor U1268 (N_1268,N_258,N_318);
nor U1269 (N_1269,N_176,In_1677);
or U1270 (N_1270,N_782,N_5);
and U1271 (N_1271,In_305,In_1523);
nor U1272 (N_1272,N_420,N_407);
xor U1273 (N_1273,N_153,N_67);
nor U1274 (N_1274,In_473,In_1018);
nor U1275 (N_1275,In_740,In_779);
and U1276 (N_1276,N_292,In_485);
nor U1277 (N_1277,N_158,N_66);
or U1278 (N_1278,N_537,N_532);
or U1279 (N_1279,In_1366,N_357);
xor U1280 (N_1280,N_708,N_173);
nand U1281 (N_1281,N_401,N_701);
and U1282 (N_1282,In_1220,N_16);
xor U1283 (N_1283,N_602,N_641);
nor U1284 (N_1284,N_729,In_1231);
nor U1285 (N_1285,In_1567,In_183);
nor U1286 (N_1286,In_209,In_1350);
nor U1287 (N_1287,In_991,N_228);
or U1288 (N_1288,In_1733,In_1032);
nor U1289 (N_1289,N_567,In_1013);
xor U1290 (N_1290,N_513,N_764);
nor U1291 (N_1291,N_172,N_797);
nand U1292 (N_1292,In_495,N_191);
or U1293 (N_1293,N_150,N_645);
nor U1294 (N_1294,N_502,In_573);
or U1295 (N_1295,In_1652,N_184);
nand U1296 (N_1296,In_1195,In_1727);
nor U1297 (N_1297,In_1305,In_620);
xnor U1298 (N_1298,N_362,N_53);
xnor U1299 (N_1299,N_226,N_366);
or U1300 (N_1300,N_65,N_355);
and U1301 (N_1301,In_394,N_799);
or U1302 (N_1302,N_373,N_133);
and U1303 (N_1303,In_1876,In_1401);
xnor U1304 (N_1304,N_749,In_203);
xnor U1305 (N_1305,N_615,N_540);
nor U1306 (N_1306,In_1096,N_180);
and U1307 (N_1307,N_415,N_134);
nor U1308 (N_1308,N_472,N_154);
nor U1309 (N_1309,N_648,In_338);
and U1310 (N_1310,In_977,N_492);
or U1311 (N_1311,N_233,In_1163);
xnor U1312 (N_1312,N_510,N_122);
and U1313 (N_1313,N_323,N_747);
xnor U1314 (N_1314,N_601,N_603);
and U1315 (N_1315,N_62,In_1561);
and U1316 (N_1316,N_533,N_542);
xor U1317 (N_1317,N_626,In_1644);
nand U1318 (N_1318,In_847,In_48);
and U1319 (N_1319,N_160,In_735);
nor U1320 (N_1320,In_498,In_144);
xnor U1321 (N_1321,In_1326,N_426);
and U1322 (N_1322,N_776,N_678);
xnor U1323 (N_1323,In_301,N_205);
or U1324 (N_1324,N_342,N_56);
or U1325 (N_1325,N_223,N_118);
nor U1326 (N_1326,N_263,In_1415);
xnor U1327 (N_1327,N_359,N_321);
or U1328 (N_1328,N_673,N_221);
nor U1329 (N_1329,N_568,N_174);
xor U1330 (N_1330,In_881,In_1461);
or U1331 (N_1331,N_311,N_293);
nand U1332 (N_1332,N_81,N_356);
nand U1333 (N_1333,In_1844,N_162);
and U1334 (N_1334,N_126,N_443);
or U1335 (N_1335,N_239,N_175);
nor U1336 (N_1336,N_616,N_168);
xor U1337 (N_1337,N_550,In_948);
nor U1338 (N_1338,N_445,N_2);
and U1339 (N_1339,In_1551,N_327);
or U1340 (N_1340,In_1073,N_762);
or U1341 (N_1341,N_428,N_39);
nor U1342 (N_1342,In_1456,In_1753);
xor U1343 (N_1343,N_378,N_404);
and U1344 (N_1344,In_788,In_1668);
or U1345 (N_1345,N_473,In_42);
nor U1346 (N_1346,N_30,In_1070);
nor U1347 (N_1347,N_503,In_974);
nor U1348 (N_1348,N_309,In_1714);
nor U1349 (N_1349,In_1754,N_370);
xor U1350 (N_1350,N_51,In_227);
or U1351 (N_1351,In_145,N_123);
nor U1352 (N_1352,In_1052,N_304);
nor U1353 (N_1353,In_165,N_587);
or U1354 (N_1354,In_1438,N_608);
and U1355 (N_1355,N_247,N_299);
nand U1356 (N_1356,In_1047,N_337);
nor U1357 (N_1357,N_121,N_422);
or U1358 (N_1358,N_37,In_1425);
xor U1359 (N_1359,In_208,N_69);
and U1360 (N_1360,In_1742,N_541);
xnor U1361 (N_1361,N_758,In_648);
nand U1362 (N_1362,In_1949,N_234);
nand U1363 (N_1363,N_591,In_429);
and U1364 (N_1364,N_326,N_668);
nor U1365 (N_1365,In_1249,In_901);
and U1366 (N_1366,In_1998,In_942);
xor U1367 (N_1367,N_120,N_149);
or U1368 (N_1368,In_1276,N_448);
xnor U1369 (N_1369,N_43,N_740);
or U1370 (N_1370,N_719,N_19);
nor U1371 (N_1371,In_978,N_605);
and U1372 (N_1372,N_260,In_1313);
and U1373 (N_1373,N_423,In_289);
xnor U1374 (N_1374,N_211,N_27);
nor U1375 (N_1375,In_1728,N_554);
or U1376 (N_1376,In_852,N_720);
and U1377 (N_1377,N_195,In_1187);
xnor U1378 (N_1378,In_1739,In_697);
and U1379 (N_1379,In_129,In_334);
or U1380 (N_1380,In_957,N_390);
xnor U1381 (N_1381,N_273,N_553);
nor U1382 (N_1382,N_147,N_392);
or U1383 (N_1383,In_1958,N_14);
or U1384 (N_1384,N_212,N_576);
and U1385 (N_1385,In_1912,N_146);
nor U1386 (N_1386,In_91,N_695);
nor U1387 (N_1387,N_786,In_1027);
or U1388 (N_1388,N_213,N_44);
xnor U1389 (N_1389,N_365,N_434);
nor U1390 (N_1390,N_343,N_224);
nand U1391 (N_1391,In_1968,N_301);
nand U1392 (N_1392,N_728,In_675);
nor U1393 (N_1393,In_1789,N_105);
nand U1394 (N_1394,N_340,N_17);
nand U1395 (N_1395,N_771,N_667);
and U1396 (N_1396,In_1007,In_631);
nor U1397 (N_1397,N_652,N_746);
or U1398 (N_1398,In_1846,In_1485);
nor U1399 (N_1399,N_185,In_1196);
nor U1400 (N_1400,N_783,N_68);
or U1401 (N_1401,In_971,In_1210);
nor U1402 (N_1402,In_1057,N_480);
nor U1403 (N_1403,N_34,In_1187);
nand U1404 (N_1404,In_315,N_281);
or U1405 (N_1405,In_1195,In_991);
nand U1406 (N_1406,In_198,N_60);
nor U1407 (N_1407,N_662,N_467);
nand U1408 (N_1408,N_490,N_15);
nor U1409 (N_1409,N_313,In_243);
xor U1410 (N_1410,N_195,N_449);
nand U1411 (N_1411,N_471,N_476);
and U1412 (N_1412,In_1526,In_1949);
xor U1413 (N_1413,In_706,N_84);
and U1414 (N_1414,N_86,N_567);
and U1415 (N_1415,N_701,N_350);
nand U1416 (N_1416,N_200,N_150);
nor U1417 (N_1417,In_1233,N_42);
nand U1418 (N_1418,N_780,N_434);
and U1419 (N_1419,N_783,In_976);
xor U1420 (N_1420,In_799,N_435);
xnor U1421 (N_1421,N_349,In_1380);
and U1422 (N_1422,N_241,N_62);
nand U1423 (N_1423,N_246,In_1416);
xnor U1424 (N_1424,In_1960,In_504);
nand U1425 (N_1425,N_257,N_134);
nand U1426 (N_1426,In_1938,N_146);
and U1427 (N_1427,In_44,In_1727);
and U1428 (N_1428,In_1664,In_1619);
and U1429 (N_1429,N_351,N_799);
nand U1430 (N_1430,N_137,In_1702);
xnor U1431 (N_1431,N_725,N_765);
xnor U1432 (N_1432,In_1831,N_512);
or U1433 (N_1433,In_205,In_678);
xnor U1434 (N_1434,N_168,N_278);
xor U1435 (N_1435,N_774,N_751);
xnor U1436 (N_1436,In_44,In_1733);
nand U1437 (N_1437,N_312,In_1702);
nor U1438 (N_1438,N_220,N_15);
nor U1439 (N_1439,N_577,N_166);
nor U1440 (N_1440,In_806,N_707);
or U1441 (N_1441,N_576,N_104);
and U1442 (N_1442,N_49,N_180);
and U1443 (N_1443,In_788,In_212);
nor U1444 (N_1444,In_1781,N_480);
nand U1445 (N_1445,N_694,N_609);
nor U1446 (N_1446,N_456,N_540);
xnor U1447 (N_1447,N_467,N_732);
and U1448 (N_1448,In_155,In_1728);
and U1449 (N_1449,In_1829,N_180);
or U1450 (N_1450,N_318,N_784);
nand U1451 (N_1451,N_430,In_1938);
and U1452 (N_1452,N_554,N_360);
xnor U1453 (N_1453,N_303,In_300);
xor U1454 (N_1454,N_54,N_223);
nand U1455 (N_1455,N_743,N_687);
and U1456 (N_1456,In_1781,In_612);
and U1457 (N_1457,In_847,N_464);
nand U1458 (N_1458,N_726,N_785);
and U1459 (N_1459,N_448,N_473);
nand U1460 (N_1460,N_550,In_1182);
and U1461 (N_1461,In_124,N_674);
and U1462 (N_1462,N_478,N_220);
or U1463 (N_1463,N_611,N_5);
nand U1464 (N_1464,N_556,In_1567);
or U1465 (N_1465,In_1677,N_416);
and U1466 (N_1466,N_795,N_464);
nand U1467 (N_1467,N_748,In_1742);
nand U1468 (N_1468,N_631,N_748);
and U1469 (N_1469,N_189,In_1027);
nand U1470 (N_1470,In_948,N_224);
or U1471 (N_1471,In_91,N_607);
or U1472 (N_1472,N_177,N_173);
or U1473 (N_1473,N_156,N_501);
and U1474 (N_1474,N_366,N_521);
nand U1475 (N_1475,N_116,N_799);
and U1476 (N_1476,In_367,N_317);
nand U1477 (N_1477,In_1133,N_661);
or U1478 (N_1478,N_563,N_777);
nor U1479 (N_1479,In_1231,In_1243);
and U1480 (N_1480,N_646,In_1074);
nor U1481 (N_1481,In_63,In_1438);
nand U1482 (N_1482,N_414,N_620);
or U1483 (N_1483,N_182,N_115);
or U1484 (N_1484,N_354,N_591);
and U1485 (N_1485,In_1846,N_738);
or U1486 (N_1486,In_1425,In_1551);
nand U1487 (N_1487,N_594,N_563);
xor U1488 (N_1488,N_282,N_607);
and U1489 (N_1489,N_731,N_570);
xnor U1490 (N_1490,N_19,N_226);
nand U1491 (N_1491,N_785,N_564);
nand U1492 (N_1492,N_110,In_1973);
or U1493 (N_1493,N_768,N_567);
nor U1494 (N_1494,In_635,N_334);
or U1495 (N_1495,In_1049,In_1370);
and U1496 (N_1496,N_392,N_98);
nand U1497 (N_1497,N_614,In_991);
xor U1498 (N_1498,N_247,In_1505);
nor U1499 (N_1499,N_21,N_614);
and U1500 (N_1500,N_509,In_205);
or U1501 (N_1501,In_589,N_44);
xnor U1502 (N_1502,N_39,N_717);
or U1503 (N_1503,N_794,N_229);
nand U1504 (N_1504,In_475,In_1714);
nor U1505 (N_1505,In_1029,N_754);
xnor U1506 (N_1506,In_1456,N_373);
nand U1507 (N_1507,N_308,N_464);
and U1508 (N_1508,N_376,N_775);
nand U1509 (N_1509,N_30,In_1854);
nand U1510 (N_1510,N_679,In_1009);
nor U1511 (N_1511,N_193,N_745);
xnor U1512 (N_1512,N_141,N_696);
and U1513 (N_1513,N_794,N_620);
xor U1514 (N_1514,N_76,N_409);
and U1515 (N_1515,N_771,N_498);
and U1516 (N_1516,In_1052,In_1640);
xor U1517 (N_1517,N_767,N_660);
xnor U1518 (N_1518,N_594,N_211);
nor U1519 (N_1519,In_644,In_1022);
xnor U1520 (N_1520,N_0,N_632);
nor U1521 (N_1521,N_784,N_314);
nand U1522 (N_1522,In_98,In_314);
nor U1523 (N_1523,N_503,N_532);
xor U1524 (N_1524,N_75,N_105);
and U1525 (N_1525,N_688,N_651);
and U1526 (N_1526,N_322,N_139);
or U1527 (N_1527,In_56,In_825);
and U1528 (N_1528,N_639,In_1514);
xnor U1529 (N_1529,N_480,N_791);
xor U1530 (N_1530,In_1163,N_416);
nand U1531 (N_1531,N_476,N_20);
nand U1532 (N_1532,In_136,N_401);
nor U1533 (N_1533,In_81,In_1047);
and U1534 (N_1534,In_1753,N_677);
xnor U1535 (N_1535,N_471,In_1644);
and U1536 (N_1536,N_275,N_244);
and U1537 (N_1537,N_232,N_590);
xnor U1538 (N_1538,N_67,In_1547);
nor U1539 (N_1539,N_157,N_211);
and U1540 (N_1540,N_465,N_466);
and U1541 (N_1541,In_104,N_128);
and U1542 (N_1542,N_681,N_324);
xor U1543 (N_1543,N_405,N_169);
nand U1544 (N_1544,N_147,N_46);
and U1545 (N_1545,In_1614,N_548);
nand U1546 (N_1546,In_1409,In_1574);
nor U1547 (N_1547,N_533,N_527);
nand U1548 (N_1548,N_34,N_413);
and U1549 (N_1549,N_668,N_41);
nor U1550 (N_1550,In_1008,In_368);
nor U1551 (N_1551,In_519,In_658);
xnor U1552 (N_1552,N_721,In_884);
nor U1553 (N_1553,N_316,N_337);
nand U1554 (N_1554,N_138,In_504);
nand U1555 (N_1555,In_1109,N_70);
nand U1556 (N_1556,In_770,In_847);
and U1557 (N_1557,N_649,N_416);
and U1558 (N_1558,N_672,In_243);
nand U1559 (N_1559,N_789,N_337);
and U1560 (N_1560,N_649,N_466);
nand U1561 (N_1561,N_386,N_452);
or U1562 (N_1562,In_421,In_1163);
and U1563 (N_1563,In_1740,N_735);
xor U1564 (N_1564,N_309,N_273);
nand U1565 (N_1565,N_442,N_559);
nor U1566 (N_1566,N_106,N_195);
nor U1567 (N_1567,N_546,N_195);
or U1568 (N_1568,In_1946,N_578);
or U1569 (N_1569,In_1521,N_455);
and U1570 (N_1570,In_203,N_786);
nand U1571 (N_1571,In_429,N_79);
xor U1572 (N_1572,N_529,In_993);
or U1573 (N_1573,N_691,N_583);
and U1574 (N_1574,N_179,N_290);
xor U1575 (N_1575,N_249,N_15);
and U1576 (N_1576,N_338,In_504);
and U1577 (N_1577,N_278,N_756);
nand U1578 (N_1578,N_237,N_559);
nor U1579 (N_1579,N_144,In_285);
nor U1580 (N_1580,In_305,N_777);
or U1581 (N_1581,In_1018,In_1438);
or U1582 (N_1582,N_26,In_1740);
and U1583 (N_1583,N_496,N_135);
and U1584 (N_1584,N_355,In_977);
or U1585 (N_1585,N_98,In_1996);
nand U1586 (N_1586,N_183,In_1876);
nand U1587 (N_1587,N_698,N_87);
nand U1588 (N_1588,N_506,N_528);
nand U1589 (N_1589,N_696,N_630);
or U1590 (N_1590,In_165,N_789);
nand U1591 (N_1591,N_597,N_524);
and U1592 (N_1592,N_468,N_453);
and U1593 (N_1593,N_715,N_777);
nor U1594 (N_1594,N_484,N_383);
nand U1595 (N_1595,N_38,N_131);
and U1596 (N_1596,N_496,In_1949);
xnor U1597 (N_1597,N_419,N_246);
and U1598 (N_1598,In_923,N_377);
and U1599 (N_1599,In_394,In_1617);
or U1600 (N_1600,N_1205,N_982);
xor U1601 (N_1601,N_1544,N_835);
nor U1602 (N_1602,N_1407,N_1250);
or U1603 (N_1603,N_1060,N_815);
nor U1604 (N_1604,N_1420,N_1073);
and U1605 (N_1605,N_1516,N_1235);
and U1606 (N_1606,N_1416,N_1541);
or U1607 (N_1607,N_1281,N_1553);
nand U1608 (N_1608,N_1288,N_1154);
and U1609 (N_1609,N_1206,N_1198);
xnor U1610 (N_1610,N_947,N_1243);
or U1611 (N_1611,N_917,N_1080);
xor U1612 (N_1612,N_1443,N_1030);
xor U1613 (N_1613,N_979,N_1240);
and U1614 (N_1614,N_1364,N_1472);
or U1615 (N_1615,N_1279,N_969);
and U1616 (N_1616,N_1136,N_1134);
nand U1617 (N_1617,N_1565,N_858);
xnor U1618 (N_1618,N_1119,N_1261);
nand U1619 (N_1619,N_829,N_961);
xnor U1620 (N_1620,N_1519,N_1373);
and U1621 (N_1621,N_1524,N_1070);
or U1622 (N_1622,N_1582,N_970);
or U1623 (N_1623,N_1123,N_1085);
nor U1624 (N_1624,N_842,N_924);
nand U1625 (N_1625,N_1367,N_1483);
nand U1626 (N_1626,N_854,N_1444);
or U1627 (N_1627,N_1458,N_997);
or U1628 (N_1628,N_1034,N_1242);
or U1629 (N_1629,N_849,N_1266);
or U1630 (N_1630,N_888,N_1564);
nand U1631 (N_1631,N_1337,N_1551);
xor U1632 (N_1632,N_1233,N_1532);
and U1633 (N_1633,N_991,N_993);
or U1634 (N_1634,N_1267,N_956);
nor U1635 (N_1635,N_1446,N_1041);
nand U1636 (N_1636,N_1063,N_1538);
xnor U1637 (N_1637,N_1112,N_977);
nand U1638 (N_1638,N_1043,N_1179);
and U1639 (N_1639,N_939,N_1380);
xor U1640 (N_1640,N_1534,N_1211);
nand U1641 (N_1641,N_812,N_1548);
or U1642 (N_1642,N_1078,N_868);
xor U1643 (N_1643,N_1020,N_1419);
nor U1644 (N_1644,N_1236,N_1103);
and U1645 (N_1645,N_978,N_1405);
and U1646 (N_1646,N_1287,N_1230);
and U1647 (N_1647,N_1015,N_1357);
xor U1648 (N_1648,N_1479,N_1387);
or U1649 (N_1649,N_1258,N_1086);
nor U1650 (N_1650,N_1019,N_1385);
xor U1651 (N_1651,N_1332,N_954);
nor U1652 (N_1652,N_1098,N_1336);
or U1653 (N_1653,N_1576,N_1511);
nand U1654 (N_1654,N_1214,N_1167);
and U1655 (N_1655,N_1526,N_811);
xnor U1656 (N_1656,N_1115,N_1454);
nor U1657 (N_1657,N_1440,N_1504);
xnor U1658 (N_1658,N_846,N_822);
nor U1659 (N_1659,N_1118,N_1330);
and U1660 (N_1660,N_1442,N_1088);
and U1661 (N_1661,N_957,N_1408);
or U1662 (N_1662,N_1592,N_1459);
and U1663 (N_1663,N_874,N_872);
and U1664 (N_1664,N_1087,N_850);
and U1665 (N_1665,N_1315,N_1201);
and U1666 (N_1666,N_1004,N_1577);
nor U1667 (N_1667,N_995,N_1274);
nand U1668 (N_1668,N_820,N_813);
nor U1669 (N_1669,N_1424,N_1505);
xor U1670 (N_1670,N_1450,N_1377);
xor U1671 (N_1671,N_1521,N_1462);
xnor U1672 (N_1672,N_996,N_900);
xnor U1673 (N_1673,N_1559,N_1161);
xnor U1674 (N_1674,N_1506,N_1189);
xor U1675 (N_1675,N_1025,N_1224);
nand U1676 (N_1676,N_1393,N_843);
nor U1677 (N_1677,N_1291,N_1071);
nand U1678 (N_1678,N_1386,N_1554);
nor U1679 (N_1679,N_955,N_1418);
and U1680 (N_1680,N_1583,N_1094);
xnor U1681 (N_1681,N_832,N_892);
nand U1682 (N_1682,N_1221,N_1245);
nand U1683 (N_1683,N_1338,N_1091);
nor U1684 (N_1684,N_926,N_1121);
xnor U1685 (N_1685,N_834,N_1421);
nand U1686 (N_1686,N_1557,N_934);
or U1687 (N_1687,N_937,N_1570);
xnor U1688 (N_1688,N_895,N_1222);
and U1689 (N_1689,N_1100,N_1067);
and U1690 (N_1690,N_1264,N_1394);
nand U1691 (N_1691,N_1590,N_1263);
nor U1692 (N_1692,N_1057,N_1110);
nand U1693 (N_1693,N_1113,N_1006);
nand U1694 (N_1694,N_1515,N_1321);
nand U1695 (N_1695,N_1275,N_929);
and U1696 (N_1696,N_1477,N_810);
nand U1697 (N_1697,N_1077,N_851);
and U1698 (N_1698,N_804,N_1493);
xor U1699 (N_1699,N_1269,N_1456);
nand U1700 (N_1700,N_1111,N_1014);
or U1701 (N_1701,N_1035,N_1527);
or U1702 (N_1702,N_1202,N_1595);
nand U1703 (N_1703,N_1135,N_1573);
or U1704 (N_1704,N_1227,N_984);
and U1705 (N_1705,N_1413,N_1574);
and U1706 (N_1706,N_1069,N_1417);
nor U1707 (N_1707,N_1422,N_994);
and U1708 (N_1708,N_1023,N_1474);
nand U1709 (N_1709,N_831,N_1089);
nor U1710 (N_1710,N_884,N_837);
or U1711 (N_1711,N_1531,N_1383);
and U1712 (N_1712,N_1178,N_1426);
or U1713 (N_1713,N_1322,N_1029);
and U1714 (N_1714,N_1163,N_894);
nand U1715 (N_1715,N_886,N_1503);
xor U1716 (N_1716,N_1523,N_1193);
nor U1717 (N_1717,N_1475,N_1268);
nand U1718 (N_1718,N_1328,N_1009);
xor U1719 (N_1719,N_1372,N_800);
nor U1720 (N_1720,N_1545,N_953);
nor U1721 (N_1721,N_1585,N_1180);
and U1722 (N_1722,N_1125,N_838);
nor U1723 (N_1723,N_919,N_1355);
and U1724 (N_1724,N_1273,N_1358);
nand U1725 (N_1725,N_827,N_1507);
or U1726 (N_1726,N_1410,N_1105);
nand U1727 (N_1727,N_1171,N_1158);
nor U1728 (N_1728,N_1514,N_1285);
or U1729 (N_1729,N_908,N_1476);
nand U1730 (N_1730,N_1348,N_1294);
nand U1731 (N_1731,N_1396,N_1297);
or U1732 (N_1732,N_1276,N_1176);
nand U1733 (N_1733,N_1594,N_1292);
xnor U1734 (N_1734,N_897,N_967);
and U1735 (N_1735,N_861,N_1032);
nand U1736 (N_1736,N_1349,N_1109);
nand U1737 (N_1737,N_1464,N_1122);
or U1738 (N_1738,N_1492,N_1449);
or U1739 (N_1739,N_1239,N_1166);
nand U1740 (N_1740,N_1191,N_1064);
xor U1741 (N_1741,N_1461,N_1153);
nand U1742 (N_1742,N_1301,N_1156);
nand U1743 (N_1743,N_1402,N_881);
nor U1744 (N_1744,N_1046,N_841);
and U1745 (N_1745,N_1145,N_1249);
and U1746 (N_1746,N_1509,N_1302);
and U1747 (N_1747,N_1467,N_1003);
xor U1748 (N_1748,N_1142,N_1342);
nor U1749 (N_1749,N_1010,N_1399);
nand U1750 (N_1750,N_1339,N_1177);
and U1751 (N_1751,N_1307,N_945);
and U1752 (N_1752,N_1150,N_1560);
and U1753 (N_1753,N_988,N_1568);
xor U1754 (N_1754,N_1219,N_949);
nand U1755 (N_1755,N_935,N_1093);
nor U1756 (N_1756,N_1575,N_1423);
or U1757 (N_1757,N_941,N_903);
xor U1758 (N_1758,N_1262,N_959);
and U1759 (N_1759,N_1429,N_1151);
nand U1760 (N_1760,N_1351,N_1453);
xnor U1761 (N_1761,N_1598,N_1096);
nand U1762 (N_1762,N_1488,N_1354);
nand U1763 (N_1763,N_867,N_1562);
nand U1764 (N_1764,N_1382,N_928);
xnor U1765 (N_1765,N_1400,N_1072);
nor U1766 (N_1766,N_855,N_1343);
and U1767 (N_1767,N_1237,N_856);
and U1768 (N_1768,N_1244,N_816);
xor U1769 (N_1769,N_1414,N_860);
or U1770 (N_1770,N_1099,N_1437);
nand U1771 (N_1771,N_1141,N_818);
xor U1772 (N_1772,N_1137,N_942);
or U1773 (N_1773,N_1207,N_1327);
nor U1774 (N_1774,N_948,N_1578);
xor U1775 (N_1775,N_1572,N_1487);
or U1776 (N_1776,N_1320,N_866);
nor U1777 (N_1777,N_833,N_1140);
and U1778 (N_1778,N_1484,N_1186);
xor U1779 (N_1779,N_1203,N_859);
xnor U1780 (N_1780,N_1312,N_1473);
and U1781 (N_1781,N_1480,N_1303);
or U1782 (N_1782,N_1319,N_1370);
and U1783 (N_1783,N_1368,N_806);
and U1784 (N_1784,N_1300,N_890);
nor U1785 (N_1785,N_1478,N_938);
xor U1786 (N_1786,N_1491,N_1016);
nand U1787 (N_1787,N_1008,N_936);
xor U1788 (N_1788,N_1164,N_1425);
xor U1789 (N_1789,N_1028,N_925);
nand U1790 (N_1790,N_1107,N_1012);
or U1791 (N_1791,N_862,N_814);
and U1792 (N_1792,N_964,N_1048);
and U1793 (N_1793,N_1318,N_1563);
and U1794 (N_1794,N_933,N_1365);
xnor U1795 (N_1795,N_1469,N_1361);
nand U1796 (N_1796,N_1068,N_887);
nand U1797 (N_1797,N_1314,N_1044);
nand U1798 (N_1798,N_1584,N_1259);
nor U1799 (N_1799,N_1173,N_1079);
and U1800 (N_1800,N_1229,N_1238);
xnor U1801 (N_1801,N_1452,N_1520);
nand U1802 (N_1802,N_1495,N_1579);
and U1803 (N_1803,N_1065,N_1311);
xor U1804 (N_1804,N_1181,N_1502);
xor U1805 (N_1805,N_1432,N_1208);
and U1806 (N_1806,N_1038,N_1284);
xnor U1807 (N_1807,N_1175,N_871);
nand U1808 (N_1808,N_1468,N_1256);
xor U1809 (N_1809,N_1018,N_1522);
nand U1810 (N_1810,N_1066,N_1129);
nor U1811 (N_1811,N_1593,N_1097);
xor U1812 (N_1812,N_1143,N_1260);
and U1813 (N_1813,N_910,N_1340);
or U1814 (N_1814,N_1092,N_817);
and U1815 (N_1815,N_819,N_1194);
nor U1816 (N_1816,N_989,N_1147);
xnor U1817 (N_1817,N_1124,N_1324);
and U1818 (N_1818,N_1555,N_1546);
nand U1819 (N_1819,N_1535,N_1362);
nand U1820 (N_1820,N_808,N_1039);
xor U1821 (N_1821,N_962,N_857);
or U1822 (N_1822,N_976,N_1257);
and U1823 (N_1823,N_836,N_1530);
nand U1824 (N_1824,N_1310,N_1172);
nor U1825 (N_1825,N_1225,N_1436);
xor U1826 (N_1826,N_1196,N_906);
xnor U1827 (N_1827,N_1498,N_1588);
xnor U1828 (N_1828,N_1460,N_1308);
nand U1829 (N_1829,N_824,N_1499);
xor U1830 (N_1830,N_1031,N_1001);
nand U1831 (N_1831,N_1363,N_1309);
or U1832 (N_1832,N_1253,N_1518);
or U1833 (N_1833,N_1101,N_1567);
or U1834 (N_1834,N_1199,N_1286);
xor U1835 (N_1835,N_1333,N_1131);
xnor U1836 (N_1836,N_873,N_1599);
nand U1837 (N_1837,N_1430,N_1438);
nand U1838 (N_1838,N_882,N_1283);
nor U1839 (N_1839,N_1525,N_968);
nand U1840 (N_1840,N_1306,N_1427);
and U1841 (N_1841,N_1289,N_1226);
or U1842 (N_1842,N_1329,N_885);
xnor U1843 (N_1843,N_913,N_1051);
nor U1844 (N_1844,N_1090,N_1587);
or U1845 (N_1845,N_932,N_1549);
xor U1846 (N_1846,N_1130,N_877);
xnor U1847 (N_1847,N_958,N_1138);
nor U1848 (N_1848,N_1200,N_980);
and U1849 (N_1849,N_1036,N_1447);
nand U1850 (N_1850,N_1074,N_966);
nor U1851 (N_1851,N_848,N_1313);
nor U1852 (N_1852,N_1183,N_809);
or U1853 (N_1853,N_1389,N_911);
nand U1854 (N_1854,N_1448,N_1106);
nand U1855 (N_1855,N_922,N_907);
or U1856 (N_1856,N_1528,N_1013);
nand U1857 (N_1857,N_1049,N_1415);
and U1858 (N_1858,N_1580,N_1381);
nand U1859 (N_1859,N_1082,N_1581);
nand U1860 (N_1860,N_927,N_1344);
or U1861 (N_1861,N_1277,N_1465);
nor U1862 (N_1862,N_840,N_1547);
xnor U1863 (N_1863,N_1021,N_1455);
xor U1864 (N_1864,N_1350,N_1061);
and U1865 (N_1865,N_863,N_1037);
nor U1866 (N_1866,N_1508,N_1395);
nor U1867 (N_1867,N_1215,N_1494);
xnor U1868 (N_1868,N_1435,N_883);
xor U1869 (N_1869,N_865,N_1102);
and U1870 (N_1870,N_1558,N_807);
or U1871 (N_1871,N_904,N_1160);
nor U1872 (N_1872,N_1155,N_830);
or U1873 (N_1873,N_1146,N_802);
or U1874 (N_1874,N_1411,N_1406);
xor U1875 (N_1875,N_1187,N_821);
nand U1876 (N_1876,N_1352,N_1571);
or U1877 (N_1877,N_1500,N_912);
and U1878 (N_1878,N_1075,N_1597);
xnor U1879 (N_1879,N_1047,N_1084);
or U1880 (N_1880,N_1378,N_1190);
or U1881 (N_1881,N_1513,N_1133);
xnor U1882 (N_1882,N_1445,N_1293);
nand U1883 (N_1883,N_1347,N_1317);
or U1884 (N_1884,N_1392,N_1005);
nand U1885 (N_1885,N_1271,N_987);
nand U1886 (N_1886,N_915,N_1168);
nand U1887 (N_1887,N_847,N_896);
and U1888 (N_1888,N_1369,N_943);
nor U1889 (N_1889,N_1374,N_1120);
and U1890 (N_1890,N_1384,N_889);
nor U1891 (N_1891,N_1404,N_1550);
or U1892 (N_1892,N_1223,N_870);
and U1893 (N_1893,N_1296,N_1512);
nand U1894 (N_1894,N_1290,N_898);
or U1895 (N_1895,N_1024,N_1536);
or U1896 (N_1896,N_1356,N_844);
nor U1897 (N_1897,N_1255,N_920);
and U1898 (N_1898,N_1316,N_1589);
and U1899 (N_1899,N_1371,N_1326);
and U1900 (N_1900,N_1482,N_1045);
nor U1901 (N_1901,N_1148,N_1388);
nor U1902 (N_1902,N_1433,N_891);
nand U1903 (N_1903,N_1108,N_869);
and U1904 (N_1904,N_1184,N_902);
and U1905 (N_1905,N_963,N_986);
or U1906 (N_1906,N_1561,N_1050);
nor U1907 (N_1907,N_1359,N_1197);
and U1908 (N_1908,N_972,N_1055);
nand U1909 (N_1909,N_1052,N_1058);
or U1910 (N_1910,N_1159,N_1298);
nand U1911 (N_1911,N_852,N_1213);
xor U1912 (N_1912,N_801,N_946);
and U1913 (N_1913,N_1537,N_1490);
nand U1914 (N_1914,N_960,N_965);
or U1915 (N_1915,N_1027,N_1501);
or U1916 (N_1916,N_1056,N_909);
nor U1917 (N_1917,N_1231,N_951);
or U1918 (N_1918,N_1246,N_1441);
or U1919 (N_1919,N_1325,N_1366);
nor U1920 (N_1920,N_1489,N_1254);
or U1921 (N_1921,N_985,N_1210);
xor U1922 (N_1922,N_899,N_1596);
xnor U1923 (N_1923,N_1000,N_805);
xor U1924 (N_1924,N_1334,N_1081);
nor U1925 (N_1925,N_1282,N_1346);
nor U1926 (N_1926,N_1412,N_825);
and U1927 (N_1927,N_1062,N_1466);
and U1928 (N_1928,N_1566,N_1533);
nand U1929 (N_1929,N_1204,N_1451);
xnor U1930 (N_1930,N_853,N_823);
nor U1931 (N_1931,N_1539,N_1241);
nand U1932 (N_1932,N_1529,N_1152);
or U1933 (N_1933,N_1220,N_1463);
and U1934 (N_1934,N_1252,N_1496);
xnor U1935 (N_1935,N_1434,N_1182);
xor U1936 (N_1936,N_1439,N_1059);
xnor U1937 (N_1937,N_1591,N_1042);
or U1938 (N_1938,N_1095,N_875);
nand U1939 (N_1939,N_1510,N_1022);
or U1940 (N_1940,N_914,N_1403);
nor U1941 (N_1941,N_1323,N_1011);
and U1942 (N_1942,N_1248,N_1542);
nor U1943 (N_1943,N_1228,N_1033);
nand U1944 (N_1944,N_1185,N_1116);
xnor U1945 (N_1945,N_940,N_1517);
or U1946 (N_1946,N_1304,N_1169);
or U1947 (N_1947,N_1128,N_1391);
nor U1948 (N_1948,N_1569,N_1127);
nor U1949 (N_1949,N_880,N_1586);
xnor U1950 (N_1950,N_998,N_1295);
and U1951 (N_1951,N_1376,N_944);
nor U1952 (N_1952,N_1165,N_1212);
xnor U1953 (N_1953,N_983,N_1379);
nor U1954 (N_1954,N_1251,N_1188);
nor U1955 (N_1955,N_1247,N_1265);
xnor U1956 (N_1956,N_878,N_1126);
nor U1957 (N_1957,N_1232,N_1139);
and U1958 (N_1958,N_916,N_1457);
xor U1959 (N_1959,N_1054,N_1053);
nand U1960 (N_1960,N_1040,N_1390);
xnor U1961 (N_1961,N_1209,N_1162);
or U1962 (N_1962,N_1192,N_828);
and U1963 (N_1963,N_1397,N_1083);
nor U1964 (N_1964,N_923,N_1117);
or U1965 (N_1965,N_1017,N_990);
or U1966 (N_1966,N_1481,N_931);
xor U1967 (N_1967,N_826,N_1278);
nor U1968 (N_1968,N_1552,N_1007);
xor U1969 (N_1969,N_1217,N_1341);
nand U1970 (N_1970,N_1299,N_1218);
and U1971 (N_1971,N_1195,N_1104);
and U1972 (N_1972,N_1335,N_1132);
and U1973 (N_1973,N_1401,N_879);
and U1974 (N_1974,N_1353,N_1497);
xor U1975 (N_1975,N_1540,N_1485);
xor U1976 (N_1976,N_1149,N_901);
or U1977 (N_1977,N_952,N_1331);
and U1978 (N_1978,N_974,N_1556);
or U1979 (N_1979,N_971,N_999);
and U1980 (N_1980,N_921,N_973);
and U1981 (N_1981,N_1174,N_1375);
nand U1982 (N_1982,N_1026,N_864);
nand U1983 (N_1983,N_1234,N_992);
nor U1984 (N_1984,N_1360,N_1409);
nor U1985 (N_1985,N_1272,N_1470);
or U1986 (N_1986,N_803,N_1157);
xor U1987 (N_1987,N_1114,N_930);
and U1988 (N_1988,N_839,N_1076);
or U1989 (N_1989,N_1270,N_1144);
nor U1990 (N_1990,N_1305,N_1398);
nand U1991 (N_1991,N_981,N_1471);
xor U1992 (N_1992,N_1170,N_1280);
xor U1993 (N_1993,N_876,N_1345);
or U1994 (N_1994,N_1428,N_893);
or U1995 (N_1995,N_918,N_1002);
nor U1996 (N_1996,N_1216,N_950);
nor U1997 (N_1997,N_845,N_1431);
or U1998 (N_1998,N_905,N_1486);
nand U1999 (N_1999,N_975,N_1543);
nand U2000 (N_2000,N_809,N_1422);
nand U2001 (N_2001,N_1401,N_952);
xor U2002 (N_2002,N_998,N_1558);
or U2003 (N_2003,N_819,N_906);
or U2004 (N_2004,N_1182,N_872);
or U2005 (N_2005,N_1279,N_1455);
nor U2006 (N_2006,N_1422,N_1040);
xor U2007 (N_2007,N_1426,N_1341);
or U2008 (N_2008,N_852,N_1550);
nand U2009 (N_2009,N_1477,N_908);
and U2010 (N_2010,N_1137,N_1126);
and U2011 (N_2011,N_1594,N_1403);
and U2012 (N_2012,N_842,N_1022);
and U2013 (N_2013,N_938,N_1127);
and U2014 (N_2014,N_1332,N_1190);
xnor U2015 (N_2015,N_1083,N_974);
nor U2016 (N_2016,N_809,N_1061);
and U2017 (N_2017,N_822,N_1236);
nand U2018 (N_2018,N_1278,N_1422);
or U2019 (N_2019,N_1257,N_1195);
and U2020 (N_2020,N_1117,N_1218);
and U2021 (N_2021,N_1398,N_1562);
nand U2022 (N_2022,N_1594,N_1586);
and U2023 (N_2023,N_1428,N_1427);
xnor U2024 (N_2024,N_1502,N_1478);
or U2025 (N_2025,N_1354,N_1441);
or U2026 (N_2026,N_1400,N_803);
and U2027 (N_2027,N_1048,N_1498);
or U2028 (N_2028,N_1146,N_1492);
xnor U2029 (N_2029,N_1488,N_1215);
nand U2030 (N_2030,N_1193,N_1420);
xor U2031 (N_2031,N_820,N_1360);
or U2032 (N_2032,N_1042,N_1244);
or U2033 (N_2033,N_1593,N_1163);
xnor U2034 (N_2034,N_897,N_1000);
nand U2035 (N_2035,N_950,N_1471);
xor U2036 (N_2036,N_1567,N_1158);
nand U2037 (N_2037,N_922,N_1564);
nand U2038 (N_2038,N_1403,N_1230);
xor U2039 (N_2039,N_1069,N_1054);
nand U2040 (N_2040,N_1189,N_896);
nand U2041 (N_2041,N_1433,N_1105);
nand U2042 (N_2042,N_1512,N_1196);
nor U2043 (N_2043,N_1142,N_1438);
xor U2044 (N_2044,N_1359,N_860);
or U2045 (N_2045,N_976,N_955);
and U2046 (N_2046,N_1115,N_1190);
nand U2047 (N_2047,N_1311,N_1514);
nor U2048 (N_2048,N_1192,N_1250);
nor U2049 (N_2049,N_1097,N_1309);
nand U2050 (N_2050,N_998,N_1031);
xor U2051 (N_2051,N_1295,N_1341);
and U2052 (N_2052,N_1228,N_1588);
nand U2053 (N_2053,N_1599,N_1272);
or U2054 (N_2054,N_1185,N_932);
xnor U2055 (N_2055,N_1429,N_1469);
xor U2056 (N_2056,N_1063,N_1533);
nand U2057 (N_2057,N_1585,N_1029);
nor U2058 (N_2058,N_934,N_1554);
and U2059 (N_2059,N_1455,N_1050);
or U2060 (N_2060,N_1144,N_1494);
nor U2061 (N_2061,N_1462,N_987);
xnor U2062 (N_2062,N_1545,N_1180);
nor U2063 (N_2063,N_961,N_1246);
nor U2064 (N_2064,N_1322,N_1030);
or U2065 (N_2065,N_1353,N_1058);
nor U2066 (N_2066,N_1166,N_1443);
and U2067 (N_2067,N_883,N_1592);
nand U2068 (N_2068,N_1084,N_1323);
xnor U2069 (N_2069,N_1234,N_881);
or U2070 (N_2070,N_1572,N_1381);
nand U2071 (N_2071,N_1301,N_921);
and U2072 (N_2072,N_1410,N_1398);
nor U2073 (N_2073,N_1083,N_1366);
nor U2074 (N_2074,N_1242,N_1069);
and U2075 (N_2075,N_1322,N_1422);
nor U2076 (N_2076,N_1035,N_1414);
xnor U2077 (N_2077,N_1209,N_1546);
xor U2078 (N_2078,N_868,N_1317);
nor U2079 (N_2079,N_999,N_1266);
or U2080 (N_2080,N_1454,N_996);
or U2081 (N_2081,N_1568,N_1267);
nand U2082 (N_2082,N_1163,N_908);
or U2083 (N_2083,N_1343,N_1292);
xor U2084 (N_2084,N_1193,N_1301);
or U2085 (N_2085,N_1447,N_1084);
or U2086 (N_2086,N_877,N_977);
or U2087 (N_2087,N_1103,N_805);
xor U2088 (N_2088,N_1079,N_875);
nand U2089 (N_2089,N_945,N_1339);
nor U2090 (N_2090,N_1141,N_1487);
xor U2091 (N_2091,N_1566,N_1476);
xnor U2092 (N_2092,N_1003,N_1047);
nand U2093 (N_2093,N_1432,N_1317);
or U2094 (N_2094,N_1390,N_1302);
nor U2095 (N_2095,N_1294,N_1160);
or U2096 (N_2096,N_1492,N_1511);
or U2097 (N_2097,N_1577,N_1039);
and U2098 (N_2098,N_1567,N_1442);
xor U2099 (N_2099,N_1387,N_1453);
nand U2100 (N_2100,N_1180,N_877);
or U2101 (N_2101,N_1357,N_973);
and U2102 (N_2102,N_985,N_812);
nand U2103 (N_2103,N_1055,N_1181);
nand U2104 (N_2104,N_1598,N_1468);
and U2105 (N_2105,N_1048,N_1070);
and U2106 (N_2106,N_864,N_1536);
nand U2107 (N_2107,N_1312,N_1335);
or U2108 (N_2108,N_1471,N_1150);
nor U2109 (N_2109,N_1010,N_1185);
or U2110 (N_2110,N_1472,N_1333);
or U2111 (N_2111,N_1106,N_1152);
or U2112 (N_2112,N_1339,N_1410);
or U2113 (N_2113,N_1159,N_1161);
nand U2114 (N_2114,N_1291,N_1292);
and U2115 (N_2115,N_1539,N_1431);
and U2116 (N_2116,N_898,N_843);
nand U2117 (N_2117,N_896,N_1110);
xor U2118 (N_2118,N_1246,N_1147);
and U2119 (N_2119,N_1560,N_1490);
nor U2120 (N_2120,N_963,N_1083);
nand U2121 (N_2121,N_1368,N_1516);
or U2122 (N_2122,N_888,N_1042);
nand U2123 (N_2123,N_1201,N_905);
nor U2124 (N_2124,N_1240,N_1271);
nor U2125 (N_2125,N_1560,N_838);
or U2126 (N_2126,N_951,N_1274);
nand U2127 (N_2127,N_1426,N_1457);
or U2128 (N_2128,N_1183,N_1173);
and U2129 (N_2129,N_913,N_1527);
nand U2130 (N_2130,N_1562,N_979);
nor U2131 (N_2131,N_1588,N_1374);
nor U2132 (N_2132,N_1493,N_863);
or U2133 (N_2133,N_816,N_1538);
and U2134 (N_2134,N_1262,N_1460);
nand U2135 (N_2135,N_962,N_913);
nand U2136 (N_2136,N_890,N_951);
xor U2137 (N_2137,N_1065,N_882);
and U2138 (N_2138,N_1513,N_1174);
xor U2139 (N_2139,N_1484,N_842);
nand U2140 (N_2140,N_865,N_1331);
nand U2141 (N_2141,N_1445,N_852);
xor U2142 (N_2142,N_1463,N_829);
xnor U2143 (N_2143,N_1004,N_1515);
nor U2144 (N_2144,N_1147,N_1586);
and U2145 (N_2145,N_1484,N_1259);
or U2146 (N_2146,N_1253,N_1368);
nand U2147 (N_2147,N_1092,N_1312);
nor U2148 (N_2148,N_1253,N_1352);
nor U2149 (N_2149,N_1292,N_1366);
nand U2150 (N_2150,N_1416,N_1092);
xor U2151 (N_2151,N_911,N_1429);
and U2152 (N_2152,N_1188,N_911);
nand U2153 (N_2153,N_1420,N_1377);
nor U2154 (N_2154,N_1542,N_1363);
nand U2155 (N_2155,N_1582,N_1061);
or U2156 (N_2156,N_1014,N_936);
and U2157 (N_2157,N_1571,N_1232);
or U2158 (N_2158,N_833,N_863);
xor U2159 (N_2159,N_1398,N_1388);
nor U2160 (N_2160,N_1388,N_1201);
and U2161 (N_2161,N_1448,N_1453);
nand U2162 (N_2162,N_1592,N_1397);
nand U2163 (N_2163,N_1443,N_1471);
and U2164 (N_2164,N_1276,N_884);
or U2165 (N_2165,N_1452,N_861);
nor U2166 (N_2166,N_1140,N_877);
xor U2167 (N_2167,N_1500,N_951);
nand U2168 (N_2168,N_1077,N_1240);
and U2169 (N_2169,N_1153,N_1556);
or U2170 (N_2170,N_994,N_1035);
or U2171 (N_2171,N_1153,N_1408);
nand U2172 (N_2172,N_1590,N_1285);
nand U2173 (N_2173,N_1258,N_1214);
nand U2174 (N_2174,N_1115,N_900);
xor U2175 (N_2175,N_1301,N_1416);
nor U2176 (N_2176,N_1201,N_1102);
or U2177 (N_2177,N_1467,N_917);
nand U2178 (N_2178,N_1305,N_1445);
nand U2179 (N_2179,N_1150,N_1556);
nand U2180 (N_2180,N_1049,N_1462);
and U2181 (N_2181,N_920,N_1223);
nand U2182 (N_2182,N_1546,N_967);
xnor U2183 (N_2183,N_970,N_939);
and U2184 (N_2184,N_1342,N_1423);
or U2185 (N_2185,N_1185,N_1310);
nand U2186 (N_2186,N_1335,N_1292);
nor U2187 (N_2187,N_1309,N_1170);
nor U2188 (N_2188,N_1439,N_1477);
nor U2189 (N_2189,N_1390,N_1287);
nor U2190 (N_2190,N_1336,N_1248);
xnor U2191 (N_2191,N_1348,N_1305);
nand U2192 (N_2192,N_984,N_1385);
or U2193 (N_2193,N_1076,N_1046);
and U2194 (N_2194,N_1251,N_831);
nand U2195 (N_2195,N_1515,N_934);
or U2196 (N_2196,N_834,N_1486);
xor U2197 (N_2197,N_981,N_1533);
and U2198 (N_2198,N_1412,N_1210);
and U2199 (N_2199,N_1310,N_1222);
or U2200 (N_2200,N_1470,N_1595);
xor U2201 (N_2201,N_1094,N_1473);
xor U2202 (N_2202,N_903,N_919);
xnor U2203 (N_2203,N_1237,N_1358);
xor U2204 (N_2204,N_1496,N_1009);
nand U2205 (N_2205,N_1401,N_1520);
xor U2206 (N_2206,N_1296,N_1005);
and U2207 (N_2207,N_1137,N_1065);
or U2208 (N_2208,N_1229,N_883);
nor U2209 (N_2209,N_1370,N_876);
nor U2210 (N_2210,N_1058,N_1474);
and U2211 (N_2211,N_947,N_1139);
or U2212 (N_2212,N_942,N_946);
nor U2213 (N_2213,N_1377,N_876);
and U2214 (N_2214,N_1133,N_1435);
and U2215 (N_2215,N_1185,N_1009);
xor U2216 (N_2216,N_1538,N_1285);
or U2217 (N_2217,N_1203,N_1210);
nand U2218 (N_2218,N_1540,N_1144);
or U2219 (N_2219,N_1423,N_1059);
xor U2220 (N_2220,N_1492,N_1003);
nand U2221 (N_2221,N_1560,N_1555);
nor U2222 (N_2222,N_1536,N_803);
and U2223 (N_2223,N_1514,N_1323);
and U2224 (N_2224,N_1101,N_1193);
xnor U2225 (N_2225,N_1073,N_880);
xnor U2226 (N_2226,N_1591,N_1397);
and U2227 (N_2227,N_1062,N_1500);
xor U2228 (N_2228,N_1361,N_1373);
nor U2229 (N_2229,N_1584,N_1032);
nand U2230 (N_2230,N_1373,N_1475);
or U2231 (N_2231,N_1352,N_1102);
and U2232 (N_2232,N_1457,N_925);
or U2233 (N_2233,N_1369,N_1541);
nor U2234 (N_2234,N_801,N_1012);
nor U2235 (N_2235,N_1289,N_1490);
nor U2236 (N_2236,N_878,N_906);
or U2237 (N_2237,N_1021,N_935);
nand U2238 (N_2238,N_1294,N_943);
or U2239 (N_2239,N_1330,N_1002);
xnor U2240 (N_2240,N_1171,N_1008);
or U2241 (N_2241,N_1029,N_1168);
nor U2242 (N_2242,N_1334,N_1256);
nand U2243 (N_2243,N_1545,N_1279);
nor U2244 (N_2244,N_1101,N_865);
nor U2245 (N_2245,N_1167,N_990);
xnor U2246 (N_2246,N_1078,N_1366);
or U2247 (N_2247,N_1170,N_879);
or U2248 (N_2248,N_1113,N_1438);
and U2249 (N_2249,N_1266,N_1009);
xnor U2250 (N_2250,N_1231,N_1328);
or U2251 (N_2251,N_1148,N_1414);
or U2252 (N_2252,N_959,N_1142);
nand U2253 (N_2253,N_1221,N_1192);
nand U2254 (N_2254,N_1270,N_1313);
and U2255 (N_2255,N_1387,N_1018);
nand U2256 (N_2256,N_1034,N_953);
or U2257 (N_2257,N_1235,N_841);
xor U2258 (N_2258,N_1220,N_1420);
or U2259 (N_2259,N_876,N_1001);
nand U2260 (N_2260,N_1055,N_1072);
nor U2261 (N_2261,N_1515,N_1031);
xnor U2262 (N_2262,N_1215,N_1258);
and U2263 (N_2263,N_1350,N_1397);
and U2264 (N_2264,N_1261,N_1411);
nor U2265 (N_2265,N_1240,N_879);
and U2266 (N_2266,N_859,N_982);
or U2267 (N_2267,N_1033,N_1201);
nor U2268 (N_2268,N_912,N_1038);
or U2269 (N_2269,N_1568,N_1168);
nor U2270 (N_2270,N_1041,N_1165);
nand U2271 (N_2271,N_1443,N_1163);
and U2272 (N_2272,N_1192,N_1457);
nand U2273 (N_2273,N_949,N_1584);
and U2274 (N_2274,N_1379,N_1350);
xor U2275 (N_2275,N_1244,N_1153);
xnor U2276 (N_2276,N_1461,N_1538);
or U2277 (N_2277,N_1146,N_1316);
and U2278 (N_2278,N_1219,N_1077);
nand U2279 (N_2279,N_1169,N_1142);
nor U2280 (N_2280,N_929,N_1261);
xor U2281 (N_2281,N_1418,N_1478);
xor U2282 (N_2282,N_1247,N_1099);
or U2283 (N_2283,N_1378,N_1400);
nor U2284 (N_2284,N_1502,N_1361);
nand U2285 (N_2285,N_1483,N_944);
xor U2286 (N_2286,N_928,N_834);
xnor U2287 (N_2287,N_1015,N_1123);
or U2288 (N_2288,N_936,N_1350);
nand U2289 (N_2289,N_1036,N_1481);
nor U2290 (N_2290,N_1332,N_1280);
xor U2291 (N_2291,N_923,N_905);
nand U2292 (N_2292,N_1047,N_823);
nor U2293 (N_2293,N_986,N_943);
nor U2294 (N_2294,N_954,N_1074);
and U2295 (N_2295,N_899,N_1113);
and U2296 (N_2296,N_1360,N_877);
nor U2297 (N_2297,N_890,N_1072);
or U2298 (N_2298,N_1002,N_1346);
nor U2299 (N_2299,N_1192,N_1503);
and U2300 (N_2300,N_1254,N_958);
xor U2301 (N_2301,N_1525,N_1194);
or U2302 (N_2302,N_1261,N_887);
and U2303 (N_2303,N_1389,N_1341);
nor U2304 (N_2304,N_850,N_1005);
nor U2305 (N_2305,N_976,N_1411);
nand U2306 (N_2306,N_1288,N_1094);
or U2307 (N_2307,N_873,N_1011);
nor U2308 (N_2308,N_1246,N_1556);
xnor U2309 (N_2309,N_1403,N_945);
or U2310 (N_2310,N_1322,N_920);
and U2311 (N_2311,N_1038,N_1587);
and U2312 (N_2312,N_873,N_840);
nor U2313 (N_2313,N_824,N_1455);
and U2314 (N_2314,N_811,N_1080);
nor U2315 (N_2315,N_1123,N_857);
nand U2316 (N_2316,N_1586,N_1347);
and U2317 (N_2317,N_952,N_969);
xor U2318 (N_2318,N_1416,N_870);
nor U2319 (N_2319,N_1587,N_1356);
nor U2320 (N_2320,N_1270,N_1586);
and U2321 (N_2321,N_1332,N_1158);
xnor U2322 (N_2322,N_1148,N_1529);
xor U2323 (N_2323,N_888,N_1117);
nor U2324 (N_2324,N_1309,N_1438);
or U2325 (N_2325,N_1140,N_977);
nand U2326 (N_2326,N_1568,N_915);
xnor U2327 (N_2327,N_1357,N_1344);
or U2328 (N_2328,N_905,N_921);
and U2329 (N_2329,N_856,N_1034);
nor U2330 (N_2330,N_1205,N_1329);
nand U2331 (N_2331,N_952,N_957);
nor U2332 (N_2332,N_1198,N_922);
xor U2333 (N_2333,N_1362,N_1269);
nor U2334 (N_2334,N_985,N_1086);
xnor U2335 (N_2335,N_825,N_1572);
and U2336 (N_2336,N_849,N_938);
or U2337 (N_2337,N_1107,N_1580);
or U2338 (N_2338,N_855,N_1429);
xor U2339 (N_2339,N_1528,N_982);
and U2340 (N_2340,N_1078,N_1573);
nor U2341 (N_2341,N_975,N_1245);
nor U2342 (N_2342,N_1033,N_1265);
nor U2343 (N_2343,N_1273,N_1464);
nor U2344 (N_2344,N_865,N_1171);
or U2345 (N_2345,N_1177,N_1369);
or U2346 (N_2346,N_996,N_1261);
and U2347 (N_2347,N_945,N_1166);
and U2348 (N_2348,N_1480,N_1161);
and U2349 (N_2349,N_1460,N_949);
nand U2350 (N_2350,N_993,N_1079);
and U2351 (N_2351,N_1212,N_1008);
and U2352 (N_2352,N_986,N_906);
xor U2353 (N_2353,N_1386,N_1026);
nor U2354 (N_2354,N_1477,N_898);
nor U2355 (N_2355,N_1157,N_1532);
and U2356 (N_2356,N_1416,N_850);
nor U2357 (N_2357,N_978,N_1130);
xor U2358 (N_2358,N_1017,N_1541);
nand U2359 (N_2359,N_966,N_1497);
and U2360 (N_2360,N_1093,N_1463);
xor U2361 (N_2361,N_1135,N_1120);
or U2362 (N_2362,N_1048,N_1492);
and U2363 (N_2363,N_1381,N_1548);
and U2364 (N_2364,N_1102,N_1598);
nand U2365 (N_2365,N_1140,N_858);
or U2366 (N_2366,N_1436,N_1358);
nor U2367 (N_2367,N_1221,N_1051);
or U2368 (N_2368,N_1208,N_1199);
and U2369 (N_2369,N_1519,N_822);
nand U2370 (N_2370,N_977,N_1001);
and U2371 (N_2371,N_1589,N_1271);
xor U2372 (N_2372,N_1006,N_1091);
or U2373 (N_2373,N_1573,N_820);
xor U2374 (N_2374,N_1011,N_1186);
nor U2375 (N_2375,N_1529,N_1254);
or U2376 (N_2376,N_872,N_1037);
nor U2377 (N_2377,N_906,N_866);
xnor U2378 (N_2378,N_1588,N_943);
nor U2379 (N_2379,N_1223,N_1428);
or U2380 (N_2380,N_1247,N_1053);
and U2381 (N_2381,N_921,N_1366);
or U2382 (N_2382,N_1520,N_1218);
xor U2383 (N_2383,N_1504,N_1501);
xor U2384 (N_2384,N_1322,N_1032);
nand U2385 (N_2385,N_1052,N_977);
nand U2386 (N_2386,N_904,N_1574);
nand U2387 (N_2387,N_936,N_959);
and U2388 (N_2388,N_938,N_883);
nor U2389 (N_2389,N_1336,N_1362);
xor U2390 (N_2390,N_1015,N_1462);
or U2391 (N_2391,N_890,N_1366);
and U2392 (N_2392,N_1443,N_1044);
nand U2393 (N_2393,N_905,N_1270);
nand U2394 (N_2394,N_890,N_834);
xor U2395 (N_2395,N_852,N_846);
nor U2396 (N_2396,N_1519,N_1049);
or U2397 (N_2397,N_857,N_950);
nor U2398 (N_2398,N_1375,N_1356);
and U2399 (N_2399,N_1193,N_971);
nor U2400 (N_2400,N_1874,N_1643);
nor U2401 (N_2401,N_2119,N_2354);
or U2402 (N_2402,N_1891,N_2174);
and U2403 (N_2403,N_1910,N_2066);
nor U2404 (N_2404,N_2360,N_1777);
nor U2405 (N_2405,N_2065,N_1832);
or U2406 (N_2406,N_1716,N_2003);
nand U2407 (N_2407,N_2345,N_1636);
nand U2408 (N_2408,N_2233,N_2293);
nor U2409 (N_2409,N_2200,N_1807);
xor U2410 (N_2410,N_2133,N_2333);
xnor U2411 (N_2411,N_1884,N_2173);
xor U2412 (N_2412,N_1943,N_2347);
and U2413 (N_2413,N_1961,N_2241);
nand U2414 (N_2414,N_2036,N_1794);
or U2415 (N_2415,N_1619,N_2280);
nor U2416 (N_2416,N_1725,N_1847);
or U2417 (N_2417,N_2145,N_1821);
and U2418 (N_2418,N_1787,N_2004);
nand U2419 (N_2419,N_2160,N_2175);
and U2420 (N_2420,N_1786,N_2052);
and U2421 (N_2421,N_1728,N_1852);
and U2422 (N_2422,N_1880,N_1984);
nand U2423 (N_2423,N_2330,N_2054);
xor U2424 (N_2424,N_1705,N_1650);
and U2425 (N_2425,N_2159,N_1945);
and U2426 (N_2426,N_2262,N_1625);
and U2427 (N_2427,N_2236,N_1676);
and U2428 (N_2428,N_1780,N_2137);
or U2429 (N_2429,N_1604,N_1686);
nand U2430 (N_2430,N_1956,N_2032);
nand U2431 (N_2431,N_2186,N_2304);
or U2432 (N_2432,N_2088,N_1843);
nor U2433 (N_2433,N_2047,N_1666);
and U2434 (N_2434,N_2115,N_2316);
and U2435 (N_2435,N_1668,N_2273);
nor U2436 (N_2436,N_2076,N_1745);
nand U2437 (N_2437,N_2080,N_1765);
xor U2438 (N_2438,N_1730,N_1746);
nor U2439 (N_2439,N_1749,N_2015);
xor U2440 (N_2440,N_1875,N_1747);
nand U2441 (N_2441,N_1848,N_2090);
and U2442 (N_2442,N_2179,N_2290);
and U2443 (N_2443,N_2298,N_2049);
nand U2444 (N_2444,N_1656,N_1939);
or U2445 (N_2445,N_1944,N_1674);
and U2446 (N_2446,N_2107,N_2388);
or U2447 (N_2447,N_2079,N_1799);
or U2448 (N_2448,N_1975,N_1648);
or U2449 (N_2449,N_2399,N_1687);
xnor U2450 (N_2450,N_1906,N_2206);
or U2451 (N_2451,N_2037,N_2039);
or U2452 (N_2452,N_2104,N_2251);
nor U2453 (N_2453,N_1743,N_1667);
nor U2454 (N_2454,N_2222,N_2148);
nand U2455 (N_2455,N_1697,N_2342);
xnor U2456 (N_2456,N_1854,N_1673);
xnor U2457 (N_2457,N_1644,N_1958);
nand U2458 (N_2458,N_1758,N_2320);
and U2459 (N_2459,N_2365,N_1767);
nor U2460 (N_2460,N_1817,N_2092);
nor U2461 (N_2461,N_1803,N_1978);
xnor U2462 (N_2462,N_2265,N_1830);
and U2463 (N_2463,N_2276,N_2191);
and U2464 (N_2464,N_2257,N_2202);
or U2465 (N_2465,N_2196,N_2213);
nand U2466 (N_2466,N_1925,N_1957);
nor U2467 (N_2467,N_1935,N_1715);
nor U2468 (N_2468,N_1699,N_2042);
nor U2469 (N_2469,N_2268,N_2194);
or U2470 (N_2470,N_1896,N_2271);
nor U2471 (N_2471,N_2162,N_1970);
xnor U2472 (N_2472,N_1640,N_1851);
nor U2473 (N_2473,N_1694,N_2114);
nor U2474 (N_2474,N_1712,N_2180);
nor U2475 (N_2475,N_2182,N_1729);
xnor U2476 (N_2476,N_1811,N_2146);
nor U2477 (N_2477,N_2382,N_1647);
nor U2478 (N_2478,N_2131,N_2156);
xnor U2479 (N_2479,N_2163,N_2309);
and U2480 (N_2480,N_1708,N_1865);
or U2481 (N_2481,N_1655,N_1789);
nand U2482 (N_2482,N_1839,N_1998);
nor U2483 (N_2483,N_2331,N_1620);
or U2484 (N_2484,N_2256,N_2327);
nor U2485 (N_2485,N_1704,N_1654);
nor U2486 (N_2486,N_2324,N_2128);
xor U2487 (N_2487,N_2310,N_1714);
xnor U2488 (N_2488,N_1937,N_2009);
nor U2489 (N_2489,N_2329,N_1952);
nand U2490 (N_2490,N_1898,N_2120);
xor U2491 (N_2491,N_2249,N_1923);
nor U2492 (N_2492,N_2151,N_2288);
and U2493 (N_2493,N_1889,N_2081);
nor U2494 (N_2494,N_1846,N_2278);
xor U2495 (N_2495,N_2025,N_1915);
xor U2496 (N_2496,N_1792,N_2197);
nand U2497 (N_2497,N_2060,N_2044);
xnor U2498 (N_2498,N_1669,N_2281);
nor U2499 (N_2499,N_2117,N_2282);
nor U2500 (N_2500,N_1649,N_2011);
or U2501 (N_2501,N_1932,N_2127);
or U2502 (N_2502,N_1633,N_2006);
and U2503 (N_2503,N_1717,N_1624);
or U2504 (N_2504,N_2231,N_2379);
or U2505 (N_2505,N_2067,N_1709);
or U2506 (N_2506,N_2242,N_2377);
or U2507 (N_2507,N_1825,N_2002);
or U2508 (N_2508,N_1735,N_1740);
and U2509 (N_2509,N_1626,N_2207);
nor U2510 (N_2510,N_1713,N_2363);
or U2511 (N_2511,N_1679,N_2258);
nor U2512 (N_2512,N_2337,N_2362);
or U2513 (N_2513,N_1942,N_1914);
or U2514 (N_2514,N_2183,N_1778);
xor U2515 (N_2515,N_1738,N_2245);
or U2516 (N_2516,N_1718,N_1903);
xor U2517 (N_2517,N_1861,N_1742);
or U2518 (N_2518,N_2118,N_1834);
nor U2519 (N_2519,N_2043,N_1719);
xnor U2520 (N_2520,N_1610,N_1701);
xnor U2521 (N_2521,N_1707,N_1741);
xor U2522 (N_2522,N_1658,N_2390);
nor U2523 (N_2523,N_2246,N_1922);
and U2524 (N_2524,N_2392,N_2167);
xnor U2525 (N_2525,N_2108,N_1993);
and U2526 (N_2526,N_1841,N_2389);
and U2527 (N_2527,N_1917,N_1857);
and U2528 (N_2528,N_2286,N_2220);
nand U2529 (N_2529,N_1801,N_1813);
xnor U2530 (N_2530,N_2210,N_1685);
and U2531 (N_2531,N_2024,N_1788);
nor U2532 (N_2532,N_2026,N_2157);
and U2533 (N_2533,N_2299,N_2274);
and U2534 (N_2534,N_1710,N_1631);
nor U2535 (N_2535,N_2164,N_2319);
and U2536 (N_2536,N_2204,N_1876);
or U2537 (N_2537,N_2121,N_1815);
and U2538 (N_2538,N_1814,N_2355);
nand U2539 (N_2539,N_2021,N_1862);
nor U2540 (N_2540,N_1809,N_2239);
xor U2541 (N_2541,N_1907,N_1842);
and U2542 (N_2542,N_1632,N_1642);
nor U2543 (N_2543,N_2103,N_2102);
and U2544 (N_2544,N_1963,N_2357);
and U2545 (N_2545,N_1659,N_1868);
and U2546 (N_2546,N_1831,N_1757);
nor U2547 (N_2547,N_1913,N_2188);
nor U2548 (N_2548,N_2283,N_1911);
or U2549 (N_2549,N_1802,N_2353);
nand U2550 (N_2550,N_1791,N_2168);
nand U2551 (N_2551,N_1886,N_1635);
or U2552 (N_2552,N_1688,N_2126);
nand U2553 (N_2553,N_2247,N_1806);
nor U2554 (N_2554,N_1623,N_1946);
or U2555 (N_2555,N_2378,N_2031);
or U2556 (N_2556,N_1881,N_2014);
or U2557 (N_2557,N_1615,N_2209);
nor U2558 (N_2558,N_2335,N_2059);
nand U2559 (N_2559,N_1905,N_1819);
or U2560 (N_2560,N_1700,N_1721);
xnor U2561 (N_2561,N_2184,N_1951);
nor U2562 (N_2562,N_1948,N_1873);
and U2563 (N_2563,N_2050,N_2123);
nand U2564 (N_2564,N_2253,N_1657);
xnor U2565 (N_2565,N_1869,N_1790);
nand U2566 (N_2566,N_2072,N_2359);
and U2567 (N_2567,N_1926,N_2226);
nor U2568 (N_2568,N_2149,N_2139);
and U2569 (N_2569,N_2314,N_2346);
nand U2570 (N_2570,N_2007,N_1678);
and U2571 (N_2571,N_2113,N_2185);
xor U2572 (N_2572,N_1971,N_2035);
xnor U2573 (N_2573,N_2308,N_1870);
nand U2574 (N_2574,N_1726,N_2208);
xnor U2575 (N_2575,N_2195,N_1810);
nor U2576 (N_2576,N_2373,N_2270);
nand U2577 (N_2577,N_2394,N_1950);
xnor U2578 (N_2578,N_1894,N_2318);
xor U2579 (N_2579,N_1645,N_2013);
or U2580 (N_2580,N_2296,N_2395);
and U2581 (N_2581,N_1621,N_1822);
xnor U2582 (N_2582,N_2348,N_2228);
nand U2583 (N_2583,N_1637,N_2255);
and U2584 (N_2584,N_1611,N_2351);
nor U2585 (N_2585,N_1639,N_1613);
xor U2586 (N_2586,N_1867,N_2074);
and U2587 (N_2587,N_1979,N_1770);
or U2588 (N_2588,N_2303,N_1805);
or U2589 (N_2589,N_2093,N_1997);
nor U2590 (N_2590,N_2078,N_2312);
nor U2591 (N_2591,N_1689,N_2305);
nor U2592 (N_2592,N_1761,N_1967);
and U2593 (N_2593,N_2223,N_2307);
xor U2594 (N_2594,N_1955,N_2277);
or U2595 (N_2595,N_2234,N_1879);
or U2596 (N_2596,N_1773,N_1722);
nor U2597 (N_2597,N_1760,N_2306);
and U2598 (N_2598,N_1949,N_1996);
and U2599 (N_2599,N_2016,N_2215);
nor U2600 (N_2600,N_2192,N_2338);
xnor U2601 (N_2601,N_2366,N_1837);
and U2602 (N_2602,N_2010,N_2205);
nor U2603 (N_2603,N_2297,N_2235);
or U2604 (N_2604,N_1693,N_2325);
nor U2605 (N_2605,N_1804,N_1681);
xor U2606 (N_2606,N_2352,N_2254);
xnor U2607 (N_2607,N_1605,N_2266);
and U2608 (N_2608,N_2252,N_2141);
or U2609 (N_2609,N_1629,N_2361);
xor U2610 (N_2610,N_1748,N_2053);
nand U2611 (N_2611,N_2100,N_2387);
and U2612 (N_2612,N_1703,N_1828);
nor U2613 (N_2613,N_2248,N_2000);
nor U2614 (N_2614,N_1606,N_2165);
nor U2615 (N_2615,N_1859,N_2094);
nor U2616 (N_2616,N_1912,N_1981);
and U2617 (N_2617,N_2048,N_2240);
nor U2618 (N_2618,N_2087,N_2029);
or U2619 (N_2619,N_2144,N_2218);
xnor U2620 (N_2620,N_1882,N_2358);
xor U2621 (N_2621,N_2155,N_2367);
or U2622 (N_2622,N_1601,N_1856);
nor U2623 (N_2623,N_2101,N_1927);
xnor U2624 (N_2624,N_1877,N_2135);
nor U2625 (N_2625,N_2030,N_2370);
xnor U2626 (N_2626,N_2152,N_2105);
nand U2627 (N_2627,N_1883,N_2012);
nand U2628 (N_2628,N_2170,N_2001);
nand U2629 (N_2629,N_1887,N_1969);
or U2630 (N_2630,N_2193,N_2064);
nand U2631 (N_2631,N_2368,N_1820);
or U2632 (N_2632,N_1863,N_2166);
xnor U2633 (N_2633,N_2109,N_2129);
xnor U2634 (N_2634,N_1994,N_1779);
and U2635 (N_2635,N_2322,N_2040);
or U2636 (N_2636,N_2301,N_1989);
or U2637 (N_2637,N_2364,N_2203);
nor U2638 (N_2638,N_2190,N_2089);
nand U2639 (N_2639,N_2311,N_2153);
or U2640 (N_2640,N_2381,N_1731);
nand U2641 (N_2641,N_1764,N_1671);
nor U2642 (N_2642,N_2398,N_2323);
nor U2643 (N_2643,N_1796,N_1824);
or U2644 (N_2644,N_2058,N_1684);
and U2645 (N_2645,N_1691,N_2350);
nand U2646 (N_2646,N_2122,N_1964);
nor U2647 (N_2647,N_1782,N_1628);
or U2648 (N_2648,N_1924,N_1720);
and U2649 (N_2649,N_1918,N_1634);
or U2650 (N_2650,N_1853,N_1763);
nor U2651 (N_2651,N_1766,N_2136);
xnor U2652 (N_2652,N_1756,N_2020);
nand U2653 (N_2653,N_1968,N_1617);
nand U2654 (N_2654,N_2385,N_1878);
and U2655 (N_2655,N_1744,N_1630);
or U2656 (N_2656,N_1947,N_2380);
xor U2657 (N_2657,N_1638,N_1808);
nor U2658 (N_2658,N_1823,N_1662);
nand U2659 (N_2659,N_2349,N_2284);
nor U2660 (N_2660,N_2275,N_1783);
or U2661 (N_2661,N_1953,N_2384);
nor U2662 (N_2662,N_1690,N_1737);
xor U2663 (N_2663,N_1973,N_1835);
xnor U2664 (N_2664,N_2272,N_2169);
and U2665 (N_2665,N_1954,N_1724);
and U2666 (N_2666,N_2369,N_2112);
and U2667 (N_2667,N_1618,N_2219);
xnor U2668 (N_2668,N_2396,N_2022);
nand U2669 (N_2669,N_2041,N_1732);
and U2670 (N_2670,N_1609,N_2143);
xnor U2671 (N_2671,N_2198,N_2383);
or U2672 (N_2672,N_2317,N_1774);
nand U2673 (N_2673,N_2097,N_1871);
nand U2674 (N_2674,N_2110,N_2372);
nand U2675 (N_2675,N_2336,N_1602);
and U2676 (N_2676,N_2328,N_2264);
and U2677 (N_2677,N_1696,N_1931);
or U2678 (N_2678,N_1739,N_1976);
and U2679 (N_2679,N_1733,N_1983);
or U2680 (N_2680,N_1916,N_2028);
xor U2681 (N_2681,N_2334,N_1921);
nor U2682 (N_2682,N_1646,N_1972);
xnor U2683 (N_2683,N_2051,N_2287);
xnor U2684 (N_2684,N_2393,N_1986);
or U2685 (N_2685,N_1776,N_1838);
nand U2686 (N_2686,N_1988,N_1670);
or U2687 (N_2687,N_2285,N_1759);
or U2688 (N_2688,N_1762,N_2138);
nand U2689 (N_2689,N_2023,N_1892);
xnor U2690 (N_2690,N_1754,N_2201);
nand U2691 (N_2691,N_2142,N_1855);
or U2692 (N_2692,N_1850,N_1622);
or U2693 (N_2693,N_2056,N_1781);
nand U2694 (N_2694,N_2294,N_1798);
xnor U2695 (N_2695,N_1600,N_1734);
nor U2696 (N_2696,N_2034,N_2147);
and U2697 (N_2697,N_1919,N_2315);
nor U2698 (N_2698,N_2181,N_1872);
or U2699 (N_2699,N_2176,N_1797);
and U2700 (N_2700,N_2085,N_2057);
xnor U2701 (N_2701,N_1885,N_2211);
xnor U2702 (N_2702,N_1812,N_2177);
and U2703 (N_2703,N_2232,N_1959);
and U2704 (N_2704,N_2106,N_2229);
nand U2705 (N_2705,N_2260,N_1936);
nor U2706 (N_2706,N_1829,N_1826);
or U2707 (N_2707,N_2221,N_2017);
and U2708 (N_2708,N_1995,N_1866);
nor U2709 (N_2709,N_2095,N_1840);
nor U2710 (N_2710,N_2062,N_1895);
or U2711 (N_2711,N_1677,N_1608);
or U2712 (N_2712,N_2096,N_1934);
and U2713 (N_2713,N_2386,N_1663);
xnor U2714 (N_2714,N_2124,N_2259);
nor U2715 (N_2715,N_1795,N_1753);
nor U2716 (N_2716,N_1752,N_1771);
and U2717 (N_2717,N_1706,N_1750);
nor U2718 (N_2718,N_2134,N_1664);
and U2719 (N_2719,N_2238,N_1900);
xor U2720 (N_2720,N_1965,N_1672);
or U2721 (N_2721,N_2140,N_1682);
or U2722 (N_2722,N_2225,N_1698);
nand U2723 (N_2723,N_2199,N_2116);
xor U2724 (N_2724,N_1768,N_1928);
nand U2725 (N_2725,N_2313,N_1616);
xor U2726 (N_2726,N_2230,N_1940);
xnor U2727 (N_2727,N_1612,N_2237);
xnor U2728 (N_2728,N_2339,N_2243);
or U2729 (N_2729,N_1897,N_2341);
nor U2730 (N_2730,N_1784,N_2130);
or U2731 (N_2731,N_2289,N_2295);
nor U2732 (N_2732,N_1818,N_1909);
xnor U2733 (N_2733,N_2045,N_2321);
nand U2734 (N_2734,N_1893,N_1941);
nand U2735 (N_2735,N_1977,N_2227);
nand U2736 (N_2736,N_2217,N_1723);
or U2737 (N_2737,N_2397,N_2077);
nor U2738 (N_2738,N_2005,N_1827);
and U2739 (N_2739,N_2158,N_1653);
nor U2740 (N_2740,N_2046,N_1962);
or U2741 (N_2741,N_2267,N_1680);
and U2742 (N_2742,N_1607,N_2292);
nand U2743 (N_2743,N_2212,N_2083);
nand U2744 (N_2744,N_1785,N_1751);
and U2745 (N_2745,N_2027,N_1683);
or U2746 (N_2746,N_1966,N_2178);
or U2747 (N_2747,N_2189,N_1816);
nand U2748 (N_2748,N_2154,N_1845);
xor U2749 (N_2749,N_2018,N_1902);
nor U2750 (N_2750,N_2068,N_2033);
xnor U2751 (N_2751,N_1920,N_2063);
nand U2752 (N_2752,N_1711,N_1769);
or U2753 (N_2753,N_2061,N_2172);
xnor U2754 (N_2754,N_1938,N_2038);
or U2755 (N_2755,N_2326,N_1836);
or U2756 (N_2756,N_2391,N_2125);
or U2757 (N_2757,N_1849,N_2376);
or U2758 (N_2758,N_2214,N_2091);
xor U2759 (N_2759,N_1641,N_1844);
or U2760 (N_2760,N_1800,N_2084);
or U2761 (N_2761,N_2344,N_1929);
or U2762 (N_2762,N_1675,N_1695);
nand U2763 (N_2763,N_1614,N_1736);
xor U2764 (N_2764,N_1858,N_1772);
or U2765 (N_2765,N_2300,N_1901);
nand U2766 (N_2766,N_2086,N_2069);
or U2767 (N_2767,N_2019,N_1930);
nand U2768 (N_2768,N_2261,N_2150);
or U2769 (N_2769,N_2099,N_1651);
nor U2770 (N_2770,N_1992,N_2356);
nor U2771 (N_2771,N_1692,N_2375);
nand U2772 (N_2772,N_2171,N_2250);
xor U2773 (N_2773,N_2302,N_1987);
nand U2774 (N_2774,N_1864,N_1985);
and U2775 (N_2775,N_2263,N_1980);
nor U2776 (N_2776,N_2279,N_2075);
xor U2777 (N_2777,N_2343,N_1793);
or U2778 (N_2778,N_2071,N_2332);
nor U2779 (N_2779,N_2291,N_2055);
xor U2780 (N_2780,N_1999,N_2371);
xor U2781 (N_2781,N_1899,N_1933);
nand U2782 (N_2782,N_2269,N_1991);
or U2783 (N_2783,N_1755,N_2070);
xor U2784 (N_2784,N_2224,N_1652);
or U2785 (N_2785,N_1860,N_1888);
and U2786 (N_2786,N_1603,N_2098);
xor U2787 (N_2787,N_2008,N_1702);
or U2788 (N_2788,N_2073,N_1660);
and U2789 (N_2789,N_1727,N_1833);
xnor U2790 (N_2790,N_1661,N_2082);
nor U2791 (N_2791,N_1775,N_1974);
or U2792 (N_2792,N_2111,N_2216);
and U2793 (N_2793,N_2374,N_1982);
xnor U2794 (N_2794,N_2132,N_2340);
and U2795 (N_2795,N_1890,N_1665);
nor U2796 (N_2796,N_1990,N_2187);
or U2797 (N_2797,N_1960,N_2161);
and U2798 (N_2798,N_1904,N_1908);
xnor U2799 (N_2799,N_1627,N_2244);
nand U2800 (N_2800,N_2175,N_1722);
and U2801 (N_2801,N_2079,N_1686);
nor U2802 (N_2802,N_2244,N_1869);
or U2803 (N_2803,N_2394,N_2291);
xnor U2804 (N_2804,N_2084,N_2376);
or U2805 (N_2805,N_2242,N_1683);
xnor U2806 (N_2806,N_2124,N_1829);
and U2807 (N_2807,N_2218,N_1978);
nand U2808 (N_2808,N_2045,N_1692);
and U2809 (N_2809,N_1958,N_2000);
or U2810 (N_2810,N_2331,N_2230);
nor U2811 (N_2811,N_1641,N_1942);
nand U2812 (N_2812,N_2335,N_2145);
and U2813 (N_2813,N_1973,N_2332);
and U2814 (N_2814,N_1705,N_1734);
xor U2815 (N_2815,N_1671,N_1745);
nand U2816 (N_2816,N_1642,N_1824);
xor U2817 (N_2817,N_1943,N_2096);
xor U2818 (N_2818,N_1977,N_1725);
xor U2819 (N_2819,N_2227,N_1924);
nand U2820 (N_2820,N_2290,N_1692);
nand U2821 (N_2821,N_2225,N_1759);
and U2822 (N_2822,N_1764,N_2220);
or U2823 (N_2823,N_2127,N_2281);
nor U2824 (N_2824,N_1864,N_1635);
nor U2825 (N_2825,N_2258,N_2232);
and U2826 (N_2826,N_2380,N_1912);
xor U2827 (N_2827,N_1728,N_2335);
nand U2828 (N_2828,N_2244,N_1619);
or U2829 (N_2829,N_2054,N_1741);
and U2830 (N_2830,N_2157,N_1881);
and U2831 (N_2831,N_1877,N_2187);
or U2832 (N_2832,N_1821,N_2227);
or U2833 (N_2833,N_2174,N_2334);
nor U2834 (N_2834,N_2068,N_1959);
and U2835 (N_2835,N_1764,N_2061);
nor U2836 (N_2836,N_1729,N_1730);
and U2837 (N_2837,N_2087,N_2387);
nand U2838 (N_2838,N_1765,N_1997);
nand U2839 (N_2839,N_2391,N_2384);
or U2840 (N_2840,N_1788,N_2373);
xor U2841 (N_2841,N_2068,N_1794);
or U2842 (N_2842,N_1728,N_1636);
nor U2843 (N_2843,N_2269,N_2306);
xnor U2844 (N_2844,N_1682,N_1851);
and U2845 (N_2845,N_1656,N_1993);
or U2846 (N_2846,N_2159,N_2076);
nand U2847 (N_2847,N_2386,N_2162);
xor U2848 (N_2848,N_1967,N_2217);
nand U2849 (N_2849,N_2182,N_1957);
nor U2850 (N_2850,N_2398,N_1939);
and U2851 (N_2851,N_2249,N_1825);
and U2852 (N_2852,N_2190,N_1999);
nor U2853 (N_2853,N_1674,N_1661);
and U2854 (N_2854,N_1610,N_2029);
nand U2855 (N_2855,N_2297,N_2063);
and U2856 (N_2856,N_1897,N_1603);
nor U2857 (N_2857,N_1765,N_2036);
or U2858 (N_2858,N_1808,N_2273);
nor U2859 (N_2859,N_2392,N_2302);
and U2860 (N_2860,N_2003,N_1904);
or U2861 (N_2861,N_1911,N_2169);
xor U2862 (N_2862,N_1861,N_2281);
nand U2863 (N_2863,N_1914,N_2304);
or U2864 (N_2864,N_1979,N_2377);
and U2865 (N_2865,N_2307,N_2362);
nor U2866 (N_2866,N_2382,N_1720);
or U2867 (N_2867,N_1804,N_2110);
nand U2868 (N_2868,N_2029,N_2184);
nor U2869 (N_2869,N_1673,N_1813);
xor U2870 (N_2870,N_2057,N_1922);
xor U2871 (N_2871,N_2005,N_2361);
or U2872 (N_2872,N_2240,N_1661);
nor U2873 (N_2873,N_1725,N_2296);
and U2874 (N_2874,N_1691,N_1736);
xnor U2875 (N_2875,N_2022,N_2200);
and U2876 (N_2876,N_2097,N_1885);
xnor U2877 (N_2877,N_1881,N_1609);
or U2878 (N_2878,N_1944,N_1636);
or U2879 (N_2879,N_2346,N_2114);
or U2880 (N_2880,N_2202,N_2029);
nor U2881 (N_2881,N_1614,N_2113);
or U2882 (N_2882,N_2103,N_2203);
nand U2883 (N_2883,N_1996,N_1881);
nor U2884 (N_2884,N_2244,N_2148);
or U2885 (N_2885,N_2035,N_1892);
nor U2886 (N_2886,N_2301,N_2030);
nor U2887 (N_2887,N_2301,N_2078);
nor U2888 (N_2888,N_2183,N_1837);
nand U2889 (N_2889,N_1653,N_1615);
nor U2890 (N_2890,N_2078,N_1874);
or U2891 (N_2891,N_1807,N_1658);
nor U2892 (N_2892,N_1786,N_1693);
or U2893 (N_2893,N_2051,N_1631);
xor U2894 (N_2894,N_1620,N_2376);
or U2895 (N_2895,N_2184,N_1943);
nand U2896 (N_2896,N_1829,N_2092);
nor U2897 (N_2897,N_1703,N_1914);
xnor U2898 (N_2898,N_1902,N_1766);
nand U2899 (N_2899,N_2027,N_2225);
nor U2900 (N_2900,N_2041,N_1829);
and U2901 (N_2901,N_2345,N_1684);
or U2902 (N_2902,N_2397,N_2141);
or U2903 (N_2903,N_1885,N_1983);
xnor U2904 (N_2904,N_1694,N_2061);
nor U2905 (N_2905,N_2258,N_1978);
xor U2906 (N_2906,N_1972,N_1758);
xor U2907 (N_2907,N_1973,N_2352);
nor U2908 (N_2908,N_2374,N_1753);
and U2909 (N_2909,N_2163,N_2036);
and U2910 (N_2910,N_1658,N_1973);
and U2911 (N_2911,N_1808,N_1668);
or U2912 (N_2912,N_1937,N_2361);
or U2913 (N_2913,N_1715,N_1966);
or U2914 (N_2914,N_1703,N_1843);
nand U2915 (N_2915,N_1738,N_2034);
and U2916 (N_2916,N_2196,N_1836);
or U2917 (N_2917,N_2051,N_2161);
or U2918 (N_2918,N_1856,N_2265);
or U2919 (N_2919,N_1660,N_2212);
xor U2920 (N_2920,N_2230,N_1709);
nor U2921 (N_2921,N_1917,N_2023);
or U2922 (N_2922,N_2156,N_2371);
xnor U2923 (N_2923,N_2071,N_2078);
nand U2924 (N_2924,N_1919,N_1817);
xor U2925 (N_2925,N_2184,N_1972);
nor U2926 (N_2926,N_2060,N_1973);
xor U2927 (N_2927,N_1614,N_1660);
or U2928 (N_2928,N_1664,N_2075);
or U2929 (N_2929,N_2125,N_2030);
nand U2930 (N_2930,N_1760,N_1833);
and U2931 (N_2931,N_2399,N_2075);
nand U2932 (N_2932,N_1631,N_1904);
or U2933 (N_2933,N_2138,N_2381);
nor U2934 (N_2934,N_2162,N_1611);
nor U2935 (N_2935,N_2193,N_1815);
nand U2936 (N_2936,N_1834,N_1909);
nor U2937 (N_2937,N_2186,N_1951);
nand U2938 (N_2938,N_2380,N_1759);
and U2939 (N_2939,N_1840,N_2270);
nand U2940 (N_2940,N_2372,N_1610);
or U2941 (N_2941,N_2211,N_1972);
nor U2942 (N_2942,N_1863,N_2033);
nor U2943 (N_2943,N_2201,N_2139);
xnor U2944 (N_2944,N_2024,N_1861);
and U2945 (N_2945,N_1911,N_2361);
or U2946 (N_2946,N_2235,N_1862);
and U2947 (N_2947,N_1939,N_1728);
xnor U2948 (N_2948,N_1865,N_1952);
xor U2949 (N_2949,N_2311,N_1741);
nor U2950 (N_2950,N_2173,N_1796);
and U2951 (N_2951,N_2242,N_2206);
nor U2952 (N_2952,N_1770,N_2329);
or U2953 (N_2953,N_2285,N_1716);
and U2954 (N_2954,N_1760,N_2294);
nor U2955 (N_2955,N_2129,N_2225);
nand U2956 (N_2956,N_1854,N_1876);
xor U2957 (N_2957,N_2228,N_2023);
nand U2958 (N_2958,N_1909,N_2187);
nand U2959 (N_2959,N_1647,N_2128);
and U2960 (N_2960,N_2219,N_1761);
xor U2961 (N_2961,N_2287,N_2223);
and U2962 (N_2962,N_2293,N_2332);
xor U2963 (N_2963,N_2016,N_1828);
nor U2964 (N_2964,N_2010,N_2333);
nor U2965 (N_2965,N_2095,N_2001);
and U2966 (N_2966,N_1921,N_2394);
nand U2967 (N_2967,N_2059,N_1640);
xnor U2968 (N_2968,N_1918,N_2201);
and U2969 (N_2969,N_2295,N_2327);
and U2970 (N_2970,N_1987,N_1671);
and U2971 (N_2971,N_2057,N_1666);
or U2972 (N_2972,N_1794,N_2136);
xor U2973 (N_2973,N_2222,N_2080);
nor U2974 (N_2974,N_1663,N_2326);
xor U2975 (N_2975,N_1882,N_2364);
nand U2976 (N_2976,N_2196,N_2125);
nand U2977 (N_2977,N_1651,N_1726);
xor U2978 (N_2978,N_1831,N_1866);
or U2979 (N_2979,N_2201,N_2376);
and U2980 (N_2980,N_2079,N_1700);
or U2981 (N_2981,N_2038,N_1958);
nand U2982 (N_2982,N_1778,N_2042);
or U2983 (N_2983,N_2344,N_2246);
and U2984 (N_2984,N_2349,N_1640);
or U2985 (N_2985,N_1849,N_2267);
xor U2986 (N_2986,N_1920,N_2312);
or U2987 (N_2987,N_1700,N_2254);
xnor U2988 (N_2988,N_1698,N_1741);
or U2989 (N_2989,N_2079,N_1864);
nor U2990 (N_2990,N_2353,N_1726);
or U2991 (N_2991,N_2134,N_2072);
nand U2992 (N_2992,N_2149,N_1851);
xnor U2993 (N_2993,N_1693,N_1750);
and U2994 (N_2994,N_2023,N_1637);
or U2995 (N_2995,N_1925,N_1768);
nand U2996 (N_2996,N_2321,N_1750);
nand U2997 (N_2997,N_2376,N_1875);
nand U2998 (N_2998,N_1692,N_1711);
nor U2999 (N_2999,N_2066,N_2021);
nand U3000 (N_3000,N_2091,N_1662);
nand U3001 (N_3001,N_1874,N_1860);
nor U3002 (N_3002,N_2050,N_1934);
or U3003 (N_3003,N_1720,N_2392);
or U3004 (N_3004,N_2003,N_1905);
and U3005 (N_3005,N_1895,N_1957);
xor U3006 (N_3006,N_1964,N_1846);
nand U3007 (N_3007,N_2038,N_1912);
xnor U3008 (N_3008,N_2357,N_1727);
and U3009 (N_3009,N_2086,N_1725);
and U3010 (N_3010,N_1812,N_2225);
nor U3011 (N_3011,N_2020,N_1694);
xor U3012 (N_3012,N_1796,N_2212);
nor U3013 (N_3013,N_2382,N_1652);
nor U3014 (N_3014,N_1795,N_1944);
nand U3015 (N_3015,N_1702,N_2014);
xor U3016 (N_3016,N_1619,N_1956);
or U3017 (N_3017,N_2142,N_1823);
nor U3018 (N_3018,N_2038,N_2043);
nand U3019 (N_3019,N_2185,N_2143);
or U3020 (N_3020,N_1749,N_1616);
or U3021 (N_3021,N_1668,N_2278);
or U3022 (N_3022,N_1729,N_2044);
or U3023 (N_3023,N_1607,N_1758);
or U3024 (N_3024,N_1807,N_1860);
or U3025 (N_3025,N_2364,N_2220);
nand U3026 (N_3026,N_1874,N_2120);
nor U3027 (N_3027,N_2252,N_2122);
xnor U3028 (N_3028,N_2204,N_2085);
or U3029 (N_3029,N_1863,N_1911);
or U3030 (N_3030,N_2355,N_2168);
nor U3031 (N_3031,N_1743,N_1765);
nor U3032 (N_3032,N_1614,N_2317);
and U3033 (N_3033,N_2000,N_1911);
xnor U3034 (N_3034,N_1901,N_2037);
nor U3035 (N_3035,N_2116,N_1951);
or U3036 (N_3036,N_1958,N_1797);
or U3037 (N_3037,N_1821,N_2031);
or U3038 (N_3038,N_1626,N_1691);
or U3039 (N_3039,N_1697,N_1894);
or U3040 (N_3040,N_2316,N_1906);
nor U3041 (N_3041,N_1775,N_1742);
nand U3042 (N_3042,N_1615,N_1744);
nor U3043 (N_3043,N_2076,N_2239);
xnor U3044 (N_3044,N_1947,N_2339);
or U3045 (N_3045,N_1925,N_1645);
nand U3046 (N_3046,N_2373,N_1971);
xor U3047 (N_3047,N_1901,N_1992);
or U3048 (N_3048,N_1932,N_1816);
xor U3049 (N_3049,N_1977,N_2284);
and U3050 (N_3050,N_2385,N_2361);
or U3051 (N_3051,N_2068,N_1939);
nor U3052 (N_3052,N_2176,N_2292);
and U3053 (N_3053,N_1894,N_2322);
nor U3054 (N_3054,N_1667,N_1725);
or U3055 (N_3055,N_1762,N_1664);
xnor U3056 (N_3056,N_2219,N_1887);
xnor U3057 (N_3057,N_1870,N_1945);
and U3058 (N_3058,N_2057,N_2326);
and U3059 (N_3059,N_1938,N_2144);
or U3060 (N_3060,N_2328,N_2043);
nor U3061 (N_3061,N_1834,N_1992);
nand U3062 (N_3062,N_1985,N_2381);
xnor U3063 (N_3063,N_2118,N_1809);
nor U3064 (N_3064,N_2011,N_1812);
xor U3065 (N_3065,N_2197,N_1832);
nand U3066 (N_3066,N_2266,N_1842);
or U3067 (N_3067,N_2006,N_1941);
or U3068 (N_3068,N_1733,N_1685);
xnor U3069 (N_3069,N_1994,N_1809);
xnor U3070 (N_3070,N_1664,N_2307);
xor U3071 (N_3071,N_2171,N_2174);
nor U3072 (N_3072,N_2006,N_2073);
xnor U3073 (N_3073,N_2359,N_2234);
nor U3074 (N_3074,N_1914,N_1854);
nor U3075 (N_3075,N_2277,N_2023);
or U3076 (N_3076,N_1929,N_1671);
nand U3077 (N_3077,N_1863,N_1714);
and U3078 (N_3078,N_2123,N_2306);
and U3079 (N_3079,N_1650,N_1723);
xor U3080 (N_3080,N_2109,N_2144);
nand U3081 (N_3081,N_1968,N_2011);
xor U3082 (N_3082,N_2143,N_1627);
nand U3083 (N_3083,N_2136,N_2133);
or U3084 (N_3084,N_1960,N_2377);
and U3085 (N_3085,N_1708,N_2147);
nand U3086 (N_3086,N_2084,N_1898);
and U3087 (N_3087,N_1886,N_2157);
and U3088 (N_3088,N_1866,N_2256);
nor U3089 (N_3089,N_2238,N_2314);
and U3090 (N_3090,N_2262,N_1678);
nor U3091 (N_3091,N_1912,N_1782);
and U3092 (N_3092,N_2354,N_1720);
xnor U3093 (N_3093,N_1697,N_1800);
xnor U3094 (N_3094,N_2184,N_2001);
nor U3095 (N_3095,N_1776,N_1928);
xor U3096 (N_3096,N_2062,N_2262);
and U3097 (N_3097,N_1780,N_2093);
nand U3098 (N_3098,N_1906,N_1903);
xnor U3099 (N_3099,N_1782,N_1687);
nor U3100 (N_3100,N_2029,N_2290);
nand U3101 (N_3101,N_1711,N_1938);
or U3102 (N_3102,N_2193,N_1947);
and U3103 (N_3103,N_1935,N_2238);
nor U3104 (N_3104,N_2370,N_2351);
and U3105 (N_3105,N_1945,N_1812);
nor U3106 (N_3106,N_1706,N_1960);
xor U3107 (N_3107,N_1733,N_2217);
and U3108 (N_3108,N_1726,N_1656);
nand U3109 (N_3109,N_1849,N_1994);
nor U3110 (N_3110,N_1966,N_2304);
nand U3111 (N_3111,N_2212,N_1881);
xnor U3112 (N_3112,N_1778,N_1637);
nand U3113 (N_3113,N_2310,N_1629);
xnor U3114 (N_3114,N_2369,N_2203);
and U3115 (N_3115,N_2380,N_1737);
and U3116 (N_3116,N_1629,N_2249);
nor U3117 (N_3117,N_2128,N_2203);
and U3118 (N_3118,N_1656,N_2132);
nand U3119 (N_3119,N_2354,N_2366);
nand U3120 (N_3120,N_1784,N_2084);
nor U3121 (N_3121,N_1968,N_1952);
nand U3122 (N_3122,N_2117,N_1600);
nor U3123 (N_3123,N_1962,N_2321);
and U3124 (N_3124,N_2341,N_1657);
nand U3125 (N_3125,N_2129,N_1937);
and U3126 (N_3126,N_1755,N_2273);
or U3127 (N_3127,N_2202,N_2393);
and U3128 (N_3128,N_2310,N_1670);
xor U3129 (N_3129,N_1626,N_1753);
nor U3130 (N_3130,N_2302,N_2170);
xor U3131 (N_3131,N_2335,N_1661);
nand U3132 (N_3132,N_2048,N_1742);
or U3133 (N_3133,N_1792,N_2106);
and U3134 (N_3134,N_2170,N_1801);
or U3135 (N_3135,N_2223,N_1654);
xor U3136 (N_3136,N_1965,N_2344);
or U3137 (N_3137,N_2352,N_1677);
xor U3138 (N_3138,N_2361,N_1969);
and U3139 (N_3139,N_1772,N_1959);
xnor U3140 (N_3140,N_2282,N_1890);
xor U3141 (N_3141,N_1744,N_1967);
nand U3142 (N_3142,N_2210,N_1620);
nand U3143 (N_3143,N_1721,N_1977);
or U3144 (N_3144,N_2187,N_2132);
xor U3145 (N_3145,N_2205,N_1805);
or U3146 (N_3146,N_1929,N_2227);
and U3147 (N_3147,N_2115,N_1766);
nor U3148 (N_3148,N_2162,N_2012);
nand U3149 (N_3149,N_2173,N_2039);
nor U3150 (N_3150,N_2392,N_2007);
xor U3151 (N_3151,N_2226,N_1888);
and U3152 (N_3152,N_2338,N_2037);
or U3153 (N_3153,N_1896,N_2103);
xnor U3154 (N_3154,N_1961,N_2144);
nor U3155 (N_3155,N_1718,N_1951);
or U3156 (N_3156,N_1915,N_2376);
xnor U3157 (N_3157,N_2268,N_1906);
and U3158 (N_3158,N_2230,N_2142);
nand U3159 (N_3159,N_2027,N_2144);
xnor U3160 (N_3160,N_2170,N_1666);
xor U3161 (N_3161,N_2141,N_2237);
nand U3162 (N_3162,N_1734,N_2105);
nor U3163 (N_3163,N_2034,N_1974);
xnor U3164 (N_3164,N_2102,N_2307);
xor U3165 (N_3165,N_2346,N_2348);
nor U3166 (N_3166,N_1899,N_1609);
or U3167 (N_3167,N_1861,N_2231);
or U3168 (N_3168,N_2275,N_2267);
xor U3169 (N_3169,N_1996,N_2000);
xnor U3170 (N_3170,N_1968,N_1897);
nor U3171 (N_3171,N_1747,N_2061);
and U3172 (N_3172,N_2280,N_2285);
nor U3173 (N_3173,N_2285,N_2172);
nand U3174 (N_3174,N_2181,N_1774);
nor U3175 (N_3175,N_2179,N_2273);
xor U3176 (N_3176,N_1942,N_2220);
nor U3177 (N_3177,N_1957,N_1911);
or U3178 (N_3178,N_1874,N_2162);
or U3179 (N_3179,N_2283,N_1862);
xnor U3180 (N_3180,N_2158,N_1943);
nor U3181 (N_3181,N_2255,N_1937);
and U3182 (N_3182,N_2021,N_1947);
or U3183 (N_3183,N_2394,N_2390);
and U3184 (N_3184,N_2256,N_1837);
and U3185 (N_3185,N_1638,N_1748);
or U3186 (N_3186,N_1671,N_1625);
xnor U3187 (N_3187,N_2273,N_1778);
nor U3188 (N_3188,N_1889,N_2180);
nand U3189 (N_3189,N_1715,N_1973);
xor U3190 (N_3190,N_2276,N_1990);
xor U3191 (N_3191,N_1786,N_1636);
xor U3192 (N_3192,N_1689,N_2323);
or U3193 (N_3193,N_1601,N_1634);
or U3194 (N_3194,N_2258,N_2171);
nor U3195 (N_3195,N_2074,N_1667);
xor U3196 (N_3196,N_2140,N_2183);
nand U3197 (N_3197,N_2342,N_2139);
and U3198 (N_3198,N_2181,N_1771);
nand U3199 (N_3199,N_1776,N_2355);
nand U3200 (N_3200,N_3120,N_2722);
or U3201 (N_3201,N_2806,N_3197);
xor U3202 (N_3202,N_2919,N_2863);
or U3203 (N_3203,N_2442,N_3144);
or U3204 (N_3204,N_2676,N_2778);
or U3205 (N_3205,N_3132,N_2413);
or U3206 (N_3206,N_3115,N_2881);
nor U3207 (N_3207,N_2695,N_2664);
and U3208 (N_3208,N_3175,N_2440);
xnor U3209 (N_3209,N_2864,N_2999);
or U3210 (N_3210,N_2993,N_2738);
xor U3211 (N_3211,N_2846,N_2563);
nand U3212 (N_3212,N_2815,N_2894);
and U3213 (N_3213,N_2735,N_2980);
and U3214 (N_3214,N_2946,N_3033);
nand U3215 (N_3215,N_2656,N_3008);
or U3216 (N_3216,N_2781,N_2857);
xnor U3217 (N_3217,N_3028,N_2928);
nand U3218 (N_3218,N_2851,N_2924);
nand U3219 (N_3219,N_3140,N_2541);
xnor U3220 (N_3220,N_3081,N_2711);
and U3221 (N_3221,N_2400,N_2606);
and U3222 (N_3222,N_2609,N_3089);
nor U3223 (N_3223,N_3125,N_3088);
nor U3224 (N_3224,N_2945,N_2532);
nor U3225 (N_3225,N_2504,N_2639);
nand U3226 (N_3226,N_3025,N_2876);
and U3227 (N_3227,N_2691,N_2506);
and U3228 (N_3228,N_3065,N_2731);
nand U3229 (N_3229,N_2721,N_2410);
xnor U3230 (N_3230,N_3138,N_2840);
nor U3231 (N_3231,N_2904,N_2907);
or U3232 (N_3232,N_2688,N_2645);
xnor U3233 (N_3233,N_2890,N_3164);
or U3234 (N_3234,N_2984,N_2720);
or U3235 (N_3235,N_2622,N_2540);
xor U3236 (N_3236,N_3075,N_2730);
or U3237 (N_3237,N_2481,N_2581);
nor U3238 (N_3238,N_2987,N_2430);
xor U3239 (N_3239,N_2403,N_3002);
xnor U3240 (N_3240,N_3198,N_2421);
nand U3241 (N_3241,N_2514,N_2478);
and U3242 (N_3242,N_2602,N_2658);
xnor U3243 (N_3243,N_3005,N_3113);
or U3244 (N_3244,N_2967,N_2424);
nand U3245 (N_3245,N_2627,N_2800);
nor U3246 (N_3246,N_3090,N_3013);
xor U3247 (N_3247,N_2943,N_2592);
nor U3248 (N_3248,N_2550,N_3024);
nand U3249 (N_3249,N_2740,N_2921);
or U3250 (N_3250,N_2401,N_2949);
and U3251 (N_3251,N_3043,N_3052);
nor U3252 (N_3252,N_2427,N_2978);
and U3253 (N_3253,N_2564,N_3072);
nor U3254 (N_3254,N_3034,N_2476);
xnor U3255 (N_3255,N_2742,N_3030);
nor U3256 (N_3256,N_2870,N_2957);
nand U3257 (N_3257,N_2775,N_3101);
or U3258 (N_3258,N_2681,N_3128);
nand U3259 (N_3259,N_2646,N_3064);
nand U3260 (N_3260,N_3083,N_2728);
xnor U3261 (N_3261,N_2764,N_2968);
nor U3262 (N_3262,N_3050,N_2958);
xor U3263 (N_3263,N_2460,N_2719);
and U3264 (N_3264,N_3047,N_2404);
nand U3265 (N_3265,N_3068,N_3119);
or U3266 (N_3266,N_2888,N_2752);
nand U3267 (N_3267,N_2572,N_2704);
and U3268 (N_3268,N_3170,N_2917);
nor U3269 (N_3269,N_2623,N_2603);
nor U3270 (N_3270,N_2573,N_2866);
or U3271 (N_3271,N_3186,N_3106);
xnor U3272 (N_3272,N_2829,N_2548);
or U3273 (N_3273,N_3146,N_3029);
and U3274 (N_3274,N_2831,N_3108);
or U3275 (N_3275,N_2977,N_3179);
or U3276 (N_3276,N_2755,N_3185);
nand U3277 (N_3277,N_2419,N_2961);
nor U3278 (N_3278,N_2845,N_2576);
and U3279 (N_3279,N_3009,N_2626);
and U3280 (N_3280,N_2791,N_3134);
nand U3281 (N_3281,N_2685,N_2471);
xnor U3282 (N_3282,N_2694,N_2431);
nand U3283 (N_3283,N_2543,N_2933);
or U3284 (N_3284,N_2426,N_2874);
and U3285 (N_3285,N_2853,N_2582);
xnor U3286 (N_3286,N_2597,N_3014);
nor U3287 (N_3287,N_2748,N_2480);
xnor U3288 (N_3288,N_3161,N_2774);
or U3289 (N_3289,N_3006,N_2590);
xor U3290 (N_3290,N_2779,N_2882);
nor U3291 (N_3291,N_3011,N_2792);
or U3292 (N_3292,N_2766,N_3093);
nor U3293 (N_3293,N_2935,N_2951);
and U3294 (N_3294,N_3103,N_2428);
nor U3295 (N_3295,N_2584,N_2544);
nor U3296 (N_3296,N_2445,N_3171);
and U3297 (N_3297,N_2560,N_2641);
nand U3298 (N_3298,N_2594,N_2830);
and U3299 (N_3299,N_2724,N_2542);
or U3300 (N_3300,N_2484,N_3145);
and U3301 (N_3301,N_2895,N_2529);
and U3302 (N_3302,N_3032,N_2652);
and U3303 (N_3303,N_2710,N_2802);
and U3304 (N_3304,N_2633,N_2976);
and U3305 (N_3305,N_2632,N_3177);
and U3306 (N_3306,N_3078,N_2556);
and U3307 (N_3307,N_2953,N_2897);
nand U3308 (N_3308,N_2447,N_2975);
nand U3309 (N_3309,N_2482,N_2679);
xnor U3310 (N_3310,N_3196,N_3135);
nor U3311 (N_3311,N_2486,N_2608);
and U3312 (N_3312,N_2959,N_2408);
or U3313 (N_3313,N_2657,N_2827);
nor U3314 (N_3314,N_2545,N_3122);
and U3315 (N_3315,N_2983,N_3053);
nor U3316 (N_3316,N_2725,N_3085);
and U3317 (N_3317,N_2449,N_3069);
nor U3318 (N_3318,N_3046,N_2687);
nand U3319 (N_3319,N_2616,N_2803);
nand U3320 (N_3320,N_2925,N_3073);
nor U3321 (N_3321,N_2816,N_2457);
or U3322 (N_3322,N_2972,N_2871);
and U3323 (N_3323,N_3184,N_2988);
xor U3324 (N_3324,N_3100,N_2726);
and U3325 (N_3325,N_3129,N_2415);
nand U3326 (N_3326,N_2466,N_2769);
nand U3327 (N_3327,N_3131,N_3157);
nand U3328 (N_3328,N_2732,N_2526);
nor U3329 (N_3329,N_2589,N_2610);
and U3330 (N_3330,N_2879,N_3151);
nor U3331 (N_3331,N_3044,N_2587);
or U3332 (N_3332,N_2452,N_3174);
nand U3333 (N_3333,N_3097,N_2750);
xnor U3334 (N_3334,N_3137,N_2528);
xnor U3335 (N_3335,N_3155,N_2865);
nand U3336 (N_3336,N_2655,N_2867);
or U3337 (N_3337,N_2797,N_2799);
nor U3338 (N_3338,N_2861,N_3020);
xnor U3339 (N_3339,N_2434,N_2783);
xnor U3340 (N_3340,N_2989,N_3082);
or U3341 (N_3341,N_3169,N_2926);
and U3342 (N_3342,N_3124,N_3036);
nand U3343 (N_3343,N_2636,N_2425);
nor U3344 (N_3344,N_2821,N_2672);
nor U3345 (N_3345,N_2841,N_3118);
and U3346 (N_3346,N_2509,N_2647);
and U3347 (N_3347,N_2765,N_3133);
xnor U3348 (N_3348,N_2673,N_2565);
and U3349 (N_3349,N_2574,N_2474);
xnor U3350 (N_3350,N_2937,N_2810);
nand U3351 (N_3351,N_3143,N_2693);
nor U3352 (N_3352,N_2773,N_2599);
nand U3353 (N_3353,N_2835,N_3156);
or U3354 (N_3354,N_2985,N_2884);
nand U3355 (N_3355,N_3192,N_2598);
nor U3356 (N_3356,N_3079,N_2669);
and U3357 (N_3357,N_2960,N_3139);
nand U3358 (N_3358,N_2561,N_3112);
or U3359 (N_3359,N_2577,N_2690);
xnor U3360 (N_3360,N_2575,N_3195);
nand U3361 (N_3361,N_2630,N_2931);
nand U3362 (N_3362,N_2838,N_3153);
xor U3363 (N_3363,N_2499,N_3194);
or U3364 (N_3364,N_2448,N_2770);
nor U3365 (N_3365,N_2796,N_2635);
and U3366 (N_3366,N_2644,N_2507);
or U3367 (N_3367,N_2776,N_2618);
nor U3368 (N_3368,N_2578,N_2569);
or U3369 (N_3369,N_3084,N_2708);
nor U3370 (N_3370,N_2600,N_2444);
or U3371 (N_3371,N_2746,N_3162);
or U3372 (N_3372,N_2734,N_3126);
and U3373 (N_3373,N_2813,N_2727);
nand U3374 (N_3374,N_2579,N_2642);
xnor U3375 (N_3375,N_2787,N_3057);
xor U3376 (N_3376,N_2903,N_2820);
nand U3377 (N_3377,N_2511,N_2786);
nand U3378 (N_3378,N_2612,N_2458);
nor U3379 (N_3379,N_2941,N_2790);
or U3380 (N_3380,N_2872,N_2530);
and U3381 (N_3381,N_3023,N_2950);
nand U3382 (N_3382,N_2498,N_3091);
and U3383 (N_3383,N_2510,N_2625);
nor U3384 (N_3384,N_2889,N_3176);
or U3385 (N_3385,N_3038,N_2605);
nand U3386 (N_3386,N_3076,N_2745);
and U3387 (N_3387,N_2604,N_2947);
and U3388 (N_3388,N_2557,N_2854);
and U3389 (N_3389,N_3042,N_2615);
and U3390 (N_3390,N_3172,N_2661);
or U3391 (N_3391,N_2450,N_2583);
or U3392 (N_3392,N_2849,N_2414);
and U3393 (N_3393,N_2753,N_2817);
and U3394 (N_3394,N_3107,N_2407);
xor U3395 (N_3395,N_2539,N_3021);
nand U3396 (N_3396,N_3063,N_3040);
nand U3397 (N_3397,N_2964,N_2525);
nor U3398 (N_3398,N_3018,N_2715);
or U3399 (N_3399,N_3074,N_2523);
or U3400 (N_3400,N_2944,N_2438);
or U3401 (N_3401,N_2472,N_2670);
or U3402 (N_3402,N_2621,N_2505);
nand U3403 (N_3403,N_2536,N_2675);
nand U3404 (N_3404,N_2789,N_2684);
and U3405 (N_3405,N_2737,N_2782);
and U3406 (N_3406,N_2952,N_2654);
and U3407 (N_3407,N_2883,N_3109);
nor U3408 (N_3408,N_2619,N_2429);
nor U3409 (N_3409,N_2887,N_2878);
or U3410 (N_3410,N_2814,N_2409);
or U3411 (N_3411,N_2828,N_2974);
and U3412 (N_3412,N_2743,N_2862);
nand U3413 (N_3413,N_3062,N_2631);
nor U3414 (N_3414,N_2520,N_2558);
nor U3415 (N_3415,N_2634,N_2406);
nor U3416 (N_3416,N_2749,N_2446);
nand U3417 (N_3417,N_2512,N_2467);
nor U3418 (N_3418,N_2848,N_2825);
or U3419 (N_3419,N_2553,N_3019);
and U3420 (N_3420,N_2809,N_2515);
or U3421 (N_3421,N_2456,N_2491);
nor U3422 (N_3422,N_2439,N_2649);
and U3423 (N_3423,N_2847,N_2703);
nand U3424 (N_3424,N_2464,N_2920);
nor U3425 (N_3425,N_3149,N_2699);
or U3426 (N_3426,N_2593,N_2822);
or U3427 (N_3427,N_2868,N_3015);
nand U3428 (N_3428,N_2683,N_2503);
nand U3429 (N_3429,N_3001,N_2762);
and U3430 (N_3430,N_2826,N_2899);
and U3431 (N_3431,N_2707,N_2911);
nor U3432 (N_3432,N_2842,N_2905);
nor U3433 (N_3433,N_3056,N_2757);
nor U3434 (N_3434,N_3022,N_2468);
nor U3435 (N_3435,N_2954,N_2873);
xor U3436 (N_3436,N_3080,N_2844);
or U3437 (N_3437,N_2858,N_3193);
xor U3438 (N_3438,N_2698,N_2518);
nor U3439 (N_3439,N_2678,N_2677);
and U3440 (N_3440,N_2516,N_3114);
xor U3441 (N_3441,N_2701,N_3182);
or U3442 (N_3442,N_2712,N_2836);
and U3443 (N_3443,N_2990,N_3105);
nand U3444 (N_3444,N_2461,N_3048);
nor U3445 (N_3445,N_3000,N_2566);
or U3446 (N_3446,N_3190,N_2758);
nor U3447 (N_3447,N_3099,N_3027);
xor U3448 (N_3448,N_2936,N_3049);
or U3449 (N_3449,N_2547,N_2521);
xnor U3450 (N_3450,N_2912,N_3154);
nand U3451 (N_3451,N_3148,N_3168);
xnor U3452 (N_3452,N_2892,N_2497);
xor U3453 (N_3453,N_2741,N_2706);
xnor U3454 (N_3454,N_2519,N_2979);
and U3455 (N_3455,N_2948,N_2513);
xor U3456 (N_3456,N_2856,N_2896);
and U3457 (N_3457,N_2549,N_2479);
xor U3458 (N_3458,N_2686,N_2780);
and U3459 (N_3459,N_3158,N_2487);
or U3460 (N_3460,N_3007,N_2568);
nor U3461 (N_3461,N_2423,N_2852);
nor U3462 (N_3462,N_2767,N_2875);
xnor U3463 (N_3463,N_2996,N_2995);
or U3464 (N_3464,N_2405,N_3180);
xor U3465 (N_3465,N_2729,N_3191);
or U3466 (N_3466,N_2420,N_2723);
nor U3467 (N_3467,N_2788,N_2805);
xor U3468 (N_3468,N_3031,N_2963);
nand U3469 (N_3469,N_2462,N_2965);
and U3470 (N_3470,N_2777,N_2760);
and U3471 (N_3471,N_3178,N_2939);
and U3472 (N_3472,N_2966,N_3167);
xor U3473 (N_3473,N_2585,N_2812);
nor U3474 (N_3474,N_2808,N_2908);
xnor U3475 (N_3475,N_2885,N_2411);
xnor U3476 (N_3476,N_2538,N_2611);
xor U3477 (N_3477,N_2763,N_3121);
nor U3478 (N_3478,N_3054,N_2860);
or U3479 (N_3479,N_3166,N_2671);
and U3480 (N_3480,N_2485,N_2682);
nor U3481 (N_3481,N_2929,N_2470);
nor U3482 (N_3482,N_2417,N_2807);
xnor U3483 (N_3483,N_2489,N_2588);
or U3484 (N_3484,N_2886,N_2665);
or U3485 (N_3485,N_2914,N_2473);
xnor U3486 (N_3486,N_2927,N_3136);
or U3487 (N_3487,N_2488,N_3039);
nor U3488 (N_3488,N_2663,N_2463);
nand U3489 (N_3489,N_3183,N_2716);
xor U3490 (N_3490,N_2620,N_2697);
nand U3491 (N_3491,N_3037,N_2680);
nand U3492 (N_3492,N_2567,N_2637);
nand U3493 (N_3493,N_3150,N_2465);
and U3494 (N_3494,N_2795,N_2591);
and U3495 (N_3495,N_2923,N_2839);
nor U3496 (N_3496,N_2955,N_2794);
xnor U3497 (N_3497,N_2824,N_3116);
nor U3498 (N_3498,N_3017,N_2898);
or U3499 (N_3499,N_2416,N_2982);
and U3500 (N_3500,N_3189,N_3117);
nor U3501 (N_3501,N_2801,N_3070);
and U3502 (N_3502,N_2934,N_2973);
and U3503 (N_3503,N_2700,N_2859);
nor U3504 (N_3504,N_2662,N_3092);
xor U3505 (N_3505,N_2546,N_2902);
or U3506 (N_3506,N_2475,N_3104);
nand U3507 (N_3507,N_3058,N_2940);
xor U3508 (N_3508,N_2648,N_3041);
xor U3509 (N_3509,N_2880,N_2580);
xor U3510 (N_3510,N_2453,N_3160);
and U3511 (N_3511,N_2768,N_2855);
nor U3512 (N_3512,N_2833,N_2651);
nor U3513 (N_3513,N_3060,N_2667);
xnor U3514 (N_3514,N_2624,N_2502);
nor U3515 (N_3515,N_2596,N_2942);
nand U3516 (N_3516,N_2744,N_3123);
or U3517 (N_3517,N_2932,N_3012);
nand U3518 (N_3518,N_2714,N_2869);
xor U3519 (N_3519,N_2494,N_2692);
or U3520 (N_3520,N_2702,N_3071);
or U3521 (N_3521,N_3066,N_3188);
or U3522 (N_3522,N_2436,N_2522);
xor U3523 (N_3523,N_2555,N_2922);
nand U3524 (N_3524,N_2994,N_2531);
nand U3525 (N_3525,N_3163,N_3004);
nor U3526 (N_3526,N_2811,N_2653);
or U3527 (N_3527,N_2422,N_2524);
nor U3528 (N_3528,N_2918,N_3045);
and U3529 (N_3529,N_2628,N_2909);
nand U3530 (N_3530,N_2747,N_3067);
nor U3531 (N_3531,N_3111,N_2517);
nand U3532 (N_3532,N_2818,N_2477);
and U3533 (N_3533,N_2804,N_2640);
nand U3534 (N_3534,N_2607,N_2493);
and U3535 (N_3535,N_3096,N_2772);
and U3536 (N_3536,N_2938,N_3181);
nor U3537 (N_3537,N_2643,N_2490);
and U3538 (N_3538,N_2877,N_2850);
nand U3539 (N_3539,N_2412,N_3051);
and U3540 (N_3540,N_2891,N_3086);
and U3541 (N_3541,N_3199,N_3102);
and U3542 (N_3542,N_2617,N_2571);
or U3543 (N_3543,N_2916,N_2534);
xnor U3544 (N_3544,N_2689,N_3055);
xor U3545 (N_3545,N_2906,N_2674);
nand U3546 (N_3546,N_2508,N_2736);
or U3547 (N_3547,N_3147,N_3016);
and U3548 (N_3548,N_3127,N_3095);
nor U3549 (N_3549,N_2696,N_2454);
and U3550 (N_3550,N_2991,N_2900);
nand U3551 (N_3551,N_2443,N_3141);
xnor U3552 (N_3552,N_2659,N_3187);
xor U3553 (N_3553,N_2533,N_2459);
and U3554 (N_3554,N_2718,N_2638);
and U3555 (N_3555,N_2650,N_2660);
nor U3556 (N_3556,N_2913,N_2793);
xor U3557 (N_3557,N_2551,N_2717);
xnor U3558 (N_3558,N_3110,N_2559);
or U3559 (N_3559,N_3026,N_2962);
or U3560 (N_3560,N_2451,N_2971);
xor U3561 (N_3561,N_2441,N_2761);
or U3562 (N_3562,N_2537,N_2562);
xor U3563 (N_3563,N_2601,N_2969);
or U3564 (N_3564,N_2586,N_2666);
and U3565 (N_3565,N_3142,N_2756);
xor U3566 (N_3566,N_3010,N_2733);
and U3567 (N_3567,N_2910,N_2798);
or U3568 (N_3568,N_2437,N_2402);
and U3569 (N_3569,N_2552,N_2501);
or U3570 (N_3570,N_3094,N_2705);
xnor U3571 (N_3571,N_2970,N_2992);
xnor U3572 (N_3572,N_2784,N_2435);
xor U3573 (N_3573,N_2713,N_3152);
xnor U3574 (N_3574,N_3061,N_2901);
xnor U3575 (N_3575,N_2455,N_2432);
nor U3576 (N_3576,N_3098,N_2893);
nor U3577 (N_3577,N_2823,N_2739);
and U3578 (N_3578,N_2930,N_2595);
nor U3579 (N_3579,N_2570,N_2956);
xor U3580 (N_3580,N_2629,N_2843);
or U3581 (N_3581,N_2483,N_2759);
and U3582 (N_3582,N_3130,N_2469);
xnor U3583 (N_3583,N_3059,N_2915);
nor U3584 (N_3584,N_3003,N_2418);
nor U3585 (N_3585,N_2785,N_3077);
and U3586 (N_3586,N_3035,N_3087);
or U3587 (N_3587,N_2535,N_2754);
nand U3588 (N_3588,N_2819,N_2709);
xor U3589 (N_3589,N_2613,N_3159);
xor U3590 (N_3590,N_2981,N_2500);
nor U3591 (N_3591,N_3165,N_2527);
nand U3592 (N_3592,N_2751,N_2496);
xor U3593 (N_3593,N_2837,N_2997);
nor U3594 (N_3594,N_2495,N_3173);
nand U3595 (N_3595,N_2771,N_2554);
or U3596 (N_3596,N_2492,N_2614);
nor U3597 (N_3597,N_2834,N_2668);
nor U3598 (N_3598,N_2986,N_2832);
xnor U3599 (N_3599,N_2998,N_2433);
and U3600 (N_3600,N_3110,N_2897);
or U3601 (N_3601,N_2638,N_2560);
or U3602 (N_3602,N_3071,N_2620);
and U3603 (N_3603,N_3100,N_2892);
and U3604 (N_3604,N_3032,N_2784);
nand U3605 (N_3605,N_2964,N_2918);
xnor U3606 (N_3606,N_2757,N_2410);
or U3607 (N_3607,N_3111,N_3056);
or U3608 (N_3608,N_2440,N_2898);
nor U3609 (N_3609,N_3059,N_2455);
and U3610 (N_3610,N_2849,N_3014);
nor U3611 (N_3611,N_2476,N_2463);
nand U3612 (N_3612,N_3071,N_3103);
or U3613 (N_3613,N_3052,N_2930);
xnor U3614 (N_3614,N_2803,N_2623);
and U3615 (N_3615,N_2994,N_2758);
nor U3616 (N_3616,N_2656,N_2702);
xor U3617 (N_3617,N_2979,N_2454);
or U3618 (N_3618,N_3148,N_2853);
xor U3619 (N_3619,N_2985,N_2581);
nor U3620 (N_3620,N_2663,N_2597);
nand U3621 (N_3621,N_2602,N_3109);
nand U3622 (N_3622,N_2441,N_2851);
nand U3623 (N_3623,N_2527,N_2448);
nand U3624 (N_3624,N_2960,N_2973);
nand U3625 (N_3625,N_3154,N_2686);
and U3626 (N_3626,N_2934,N_2454);
nor U3627 (N_3627,N_2596,N_2626);
and U3628 (N_3628,N_2885,N_2930);
xnor U3629 (N_3629,N_2996,N_2857);
xnor U3630 (N_3630,N_2817,N_2541);
nor U3631 (N_3631,N_2600,N_2510);
nand U3632 (N_3632,N_3025,N_2954);
nand U3633 (N_3633,N_3014,N_3147);
or U3634 (N_3634,N_2597,N_2695);
nor U3635 (N_3635,N_2966,N_2569);
or U3636 (N_3636,N_2428,N_2886);
nor U3637 (N_3637,N_3153,N_2798);
nor U3638 (N_3638,N_3051,N_3144);
or U3639 (N_3639,N_2978,N_2958);
nor U3640 (N_3640,N_2950,N_2614);
nand U3641 (N_3641,N_2473,N_2881);
nand U3642 (N_3642,N_3101,N_2561);
xor U3643 (N_3643,N_2990,N_2613);
or U3644 (N_3644,N_3199,N_3151);
and U3645 (N_3645,N_2744,N_2512);
or U3646 (N_3646,N_2607,N_2904);
or U3647 (N_3647,N_3085,N_2794);
and U3648 (N_3648,N_2933,N_3062);
xnor U3649 (N_3649,N_2430,N_3133);
and U3650 (N_3650,N_2917,N_3144);
nor U3651 (N_3651,N_2893,N_3046);
and U3652 (N_3652,N_2611,N_2922);
and U3653 (N_3653,N_2559,N_2829);
nand U3654 (N_3654,N_2989,N_2777);
and U3655 (N_3655,N_2525,N_3060);
or U3656 (N_3656,N_2457,N_2894);
nor U3657 (N_3657,N_3043,N_2414);
and U3658 (N_3658,N_2764,N_2639);
nor U3659 (N_3659,N_2760,N_2885);
nor U3660 (N_3660,N_2944,N_2792);
and U3661 (N_3661,N_2431,N_2837);
or U3662 (N_3662,N_2597,N_2630);
and U3663 (N_3663,N_2766,N_2885);
xnor U3664 (N_3664,N_3073,N_2603);
xnor U3665 (N_3665,N_2554,N_2667);
or U3666 (N_3666,N_2496,N_2890);
or U3667 (N_3667,N_3180,N_3111);
and U3668 (N_3668,N_2763,N_2735);
or U3669 (N_3669,N_2737,N_2456);
nand U3670 (N_3670,N_2878,N_2483);
and U3671 (N_3671,N_2434,N_2960);
and U3672 (N_3672,N_3134,N_2737);
nor U3673 (N_3673,N_2532,N_2826);
or U3674 (N_3674,N_2508,N_2777);
and U3675 (N_3675,N_2839,N_2718);
or U3676 (N_3676,N_2559,N_3153);
or U3677 (N_3677,N_2737,N_2764);
xor U3678 (N_3678,N_2931,N_2906);
or U3679 (N_3679,N_2951,N_3135);
and U3680 (N_3680,N_3184,N_2908);
or U3681 (N_3681,N_3163,N_2408);
nand U3682 (N_3682,N_3015,N_2529);
xnor U3683 (N_3683,N_3162,N_2705);
nand U3684 (N_3684,N_2494,N_2928);
or U3685 (N_3685,N_2447,N_3195);
xor U3686 (N_3686,N_2827,N_3075);
nor U3687 (N_3687,N_2998,N_3137);
nand U3688 (N_3688,N_2879,N_2470);
and U3689 (N_3689,N_3038,N_2575);
xor U3690 (N_3690,N_2739,N_2490);
nand U3691 (N_3691,N_2674,N_2464);
xor U3692 (N_3692,N_3141,N_2849);
and U3693 (N_3693,N_3099,N_2624);
nor U3694 (N_3694,N_2977,N_2900);
and U3695 (N_3695,N_3177,N_2874);
nand U3696 (N_3696,N_2873,N_2655);
and U3697 (N_3697,N_3111,N_2633);
or U3698 (N_3698,N_2509,N_2957);
xnor U3699 (N_3699,N_2832,N_2438);
or U3700 (N_3700,N_3061,N_2715);
nand U3701 (N_3701,N_2983,N_2497);
or U3702 (N_3702,N_2733,N_2592);
or U3703 (N_3703,N_2659,N_2809);
nand U3704 (N_3704,N_2600,N_2861);
or U3705 (N_3705,N_3125,N_2639);
xnor U3706 (N_3706,N_2564,N_2776);
nand U3707 (N_3707,N_2855,N_3155);
and U3708 (N_3708,N_2703,N_3034);
nor U3709 (N_3709,N_2975,N_2469);
nand U3710 (N_3710,N_3187,N_2946);
and U3711 (N_3711,N_2693,N_3085);
nand U3712 (N_3712,N_3058,N_2580);
nor U3713 (N_3713,N_2891,N_2669);
xor U3714 (N_3714,N_3145,N_2676);
xor U3715 (N_3715,N_2439,N_2692);
xor U3716 (N_3716,N_2744,N_2940);
or U3717 (N_3717,N_3142,N_2445);
xnor U3718 (N_3718,N_2672,N_2733);
nor U3719 (N_3719,N_2947,N_2550);
xor U3720 (N_3720,N_2415,N_3059);
or U3721 (N_3721,N_3166,N_3031);
nand U3722 (N_3722,N_2992,N_2665);
and U3723 (N_3723,N_2976,N_3190);
or U3724 (N_3724,N_3178,N_2676);
nand U3725 (N_3725,N_2567,N_2752);
nand U3726 (N_3726,N_2917,N_2672);
xor U3727 (N_3727,N_2425,N_3179);
xnor U3728 (N_3728,N_2479,N_2593);
and U3729 (N_3729,N_2531,N_2890);
or U3730 (N_3730,N_2623,N_2721);
xnor U3731 (N_3731,N_2951,N_2667);
and U3732 (N_3732,N_2998,N_2990);
or U3733 (N_3733,N_2426,N_3180);
nand U3734 (N_3734,N_2850,N_2665);
or U3735 (N_3735,N_2624,N_2933);
and U3736 (N_3736,N_2883,N_3143);
nor U3737 (N_3737,N_3139,N_2847);
or U3738 (N_3738,N_2836,N_3148);
nor U3739 (N_3739,N_3089,N_2906);
and U3740 (N_3740,N_2966,N_2601);
and U3741 (N_3741,N_3035,N_3054);
or U3742 (N_3742,N_2508,N_2410);
and U3743 (N_3743,N_2847,N_2782);
xnor U3744 (N_3744,N_2505,N_2614);
nand U3745 (N_3745,N_3140,N_2794);
xor U3746 (N_3746,N_3124,N_2493);
or U3747 (N_3747,N_2981,N_2426);
and U3748 (N_3748,N_2563,N_3015);
and U3749 (N_3749,N_2688,N_2844);
xor U3750 (N_3750,N_2546,N_2660);
or U3751 (N_3751,N_2564,N_3138);
xnor U3752 (N_3752,N_2783,N_2869);
xnor U3753 (N_3753,N_3056,N_3070);
nor U3754 (N_3754,N_3053,N_2872);
nand U3755 (N_3755,N_2440,N_2809);
and U3756 (N_3756,N_2993,N_2811);
and U3757 (N_3757,N_2596,N_2825);
and U3758 (N_3758,N_2733,N_2679);
and U3759 (N_3759,N_3106,N_2896);
nor U3760 (N_3760,N_2604,N_2521);
nand U3761 (N_3761,N_2758,N_2995);
nor U3762 (N_3762,N_3163,N_2811);
and U3763 (N_3763,N_2573,N_2479);
nor U3764 (N_3764,N_2723,N_3182);
nor U3765 (N_3765,N_2987,N_2686);
nand U3766 (N_3766,N_2770,N_2722);
nor U3767 (N_3767,N_2554,N_2894);
nor U3768 (N_3768,N_2998,N_2441);
nor U3769 (N_3769,N_2975,N_3026);
nand U3770 (N_3770,N_3050,N_2852);
nand U3771 (N_3771,N_2516,N_3013);
nand U3772 (N_3772,N_2539,N_2778);
or U3773 (N_3773,N_2951,N_2955);
nor U3774 (N_3774,N_2431,N_2516);
xnor U3775 (N_3775,N_3052,N_2567);
nor U3776 (N_3776,N_3179,N_2560);
nand U3777 (N_3777,N_2570,N_3101);
nor U3778 (N_3778,N_2809,N_3150);
nor U3779 (N_3779,N_2993,N_2878);
and U3780 (N_3780,N_2908,N_2762);
nor U3781 (N_3781,N_2525,N_2578);
nor U3782 (N_3782,N_2898,N_2654);
or U3783 (N_3783,N_2583,N_2912);
and U3784 (N_3784,N_2680,N_2884);
nor U3785 (N_3785,N_3046,N_2453);
and U3786 (N_3786,N_3154,N_3183);
nor U3787 (N_3787,N_2591,N_3053);
and U3788 (N_3788,N_2906,N_2583);
and U3789 (N_3789,N_2993,N_2474);
xor U3790 (N_3790,N_3127,N_2412);
and U3791 (N_3791,N_2886,N_2644);
or U3792 (N_3792,N_2822,N_2710);
or U3793 (N_3793,N_2492,N_3073);
nor U3794 (N_3794,N_2595,N_2607);
xor U3795 (N_3795,N_3170,N_2922);
and U3796 (N_3796,N_2977,N_2710);
and U3797 (N_3797,N_2711,N_2787);
or U3798 (N_3798,N_3117,N_2512);
and U3799 (N_3799,N_2835,N_3005);
and U3800 (N_3800,N_2765,N_2939);
and U3801 (N_3801,N_3119,N_3092);
nand U3802 (N_3802,N_2645,N_2915);
and U3803 (N_3803,N_2828,N_2576);
nand U3804 (N_3804,N_2653,N_3007);
or U3805 (N_3805,N_2409,N_3160);
xnor U3806 (N_3806,N_2454,N_2701);
nand U3807 (N_3807,N_2527,N_2561);
xor U3808 (N_3808,N_2794,N_2640);
nand U3809 (N_3809,N_2653,N_3100);
or U3810 (N_3810,N_3199,N_2705);
nor U3811 (N_3811,N_2861,N_2710);
or U3812 (N_3812,N_2737,N_2514);
or U3813 (N_3813,N_2942,N_3089);
nand U3814 (N_3814,N_2916,N_3156);
and U3815 (N_3815,N_3029,N_2532);
and U3816 (N_3816,N_2411,N_2514);
and U3817 (N_3817,N_3100,N_3119);
xnor U3818 (N_3818,N_2739,N_2654);
xnor U3819 (N_3819,N_3098,N_2489);
nor U3820 (N_3820,N_2728,N_2939);
nor U3821 (N_3821,N_2997,N_2720);
or U3822 (N_3822,N_2577,N_2816);
xnor U3823 (N_3823,N_2414,N_2745);
and U3824 (N_3824,N_2924,N_2490);
nor U3825 (N_3825,N_2457,N_2590);
and U3826 (N_3826,N_2630,N_2532);
nor U3827 (N_3827,N_2434,N_3184);
xor U3828 (N_3828,N_2859,N_2931);
xor U3829 (N_3829,N_3040,N_2462);
nor U3830 (N_3830,N_3089,N_3087);
nor U3831 (N_3831,N_2685,N_3065);
nand U3832 (N_3832,N_2466,N_2794);
and U3833 (N_3833,N_2815,N_2574);
nor U3834 (N_3834,N_2453,N_2765);
xor U3835 (N_3835,N_2784,N_3055);
nand U3836 (N_3836,N_2874,N_2765);
or U3837 (N_3837,N_2755,N_2599);
xor U3838 (N_3838,N_3026,N_2907);
nor U3839 (N_3839,N_3149,N_2737);
or U3840 (N_3840,N_2542,N_2974);
nor U3841 (N_3841,N_3026,N_3141);
nand U3842 (N_3842,N_2719,N_3087);
xnor U3843 (N_3843,N_3049,N_3056);
and U3844 (N_3844,N_3028,N_2467);
and U3845 (N_3845,N_3133,N_2819);
nand U3846 (N_3846,N_3156,N_2679);
xnor U3847 (N_3847,N_2718,N_3070);
xnor U3848 (N_3848,N_3164,N_3172);
and U3849 (N_3849,N_3196,N_3038);
and U3850 (N_3850,N_2478,N_2715);
nand U3851 (N_3851,N_2986,N_2627);
xnor U3852 (N_3852,N_2439,N_3145);
xnor U3853 (N_3853,N_2676,N_2543);
or U3854 (N_3854,N_2922,N_2714);
and U3855 (N_3855,N_2885,N_2814);
nor U3856 (N_3856,N_2815,N_2784);
nor U3857 (N_3857,N_3178,N_3050);
nand U3858 (N_3858,N_3115,N_2582);
and U3859 (N_3859,N_3041,N_2715);
or U3860 (N_3860,N_2466,N_2726);
xnor U3861 (N_3861,N_2981,N_3105);
xor U3862 (N_3862,N_3033,N_2907);
nor U3863 (N_3863,N_2873,N_3000);
xnor U3864 (N_3864,N_3181,N_3146);
and U3865 (N_3865,N_2728,N_2784);
and U3866 (N_3866,N_3045,N_2737);
and U3867 (N_3867,N_3057,N_2530);
and U3868 (N_3868,N_2677,N_3087);
nand U3869 (N_3869,N_2554,N_3106);
and U3870 (N_3870,N_2769,N_3150);
or U3871 (N_3871,N_2607,N_2987);
xor U3872 (N_3872,N_2531,N_3076);
nor U3873 (N_3873,N_2665,N_2899);
or U3874 (N_3874,N_2957,N_2553);
nand U3875 (N_3875,N_3109,N_2900);
nand U3876 (N_3876,N_2415,N_2804);
and U3877 (N_3877,N_3192,N_2770);
nand U3878 (N_3878,N_3075,N_3114);
nand U3879 (N_3879,N_3029,N_2749);
xnor U3880 (N_3880,N_2815,N_2831);
and U3881 (N_3881,N_3017,N_2864);
nor U3882 (N_3882,N_2801,N_3147);
xor U3883 (N_3883,N_2712,N_3029);
xor U3884 (N_3884,N_3014,N_2862);
and U3885 (N_3885,N_2678,N_2735);
or U3886 (N_3886,N_2700,N_2899);
nand U3887 (N_3887,N_3185,N_3091);
nor U3888 (N_3888,N_2950,N_3174);
nor U3889 (N_3889,N_2580,N_2506);
nand U3890 (N_3890,N_2880,N_2402);
and U3891 (N_3891,N_2724,N_2983);
or U3892 (N_3892,N_2753,N_2813);
or U3893 (N_3893,N_2859,N_3106);
xnor U3894 (N_3894,N_2420,N_2499);
and U3895 (N_3895,N_3160,N_2822);
or U3896 (N_3896,N_2923,N_2773);
or U3897 (N_3897,N_2502,N_2475);
nand U3898 (N_3898,N_2633,N_2815);
and U3899 (N_3899,N_2593,N_2431);
xor U3900 (N_3900,N_2626,N_3182);
xor U3901 (N_3901,N_3175,N_2781);
nand U3902 (N_3902,N_2712,N_3102);
or U3903 (N_3903,N_3000,N_2458);
nand U3904 (N_3904,N_2619,N_2729);
and U3905 (N_3905,N_2712,N_2926);
and U3906 (N_3906,N_2506,N_2919);
or U3907 (N_3907,N_2561,N_3066);
or U3908 (N_3908,N_2739,N_2716);
and U3909 (N_3909,N_2625,N_2439);
and U3910 (N_3910,N_2915,N_2411);
xor U3911 (N_3911,N_2756,N_2875);
and U3912 (N_3912,N_2651,N_2436);
and U3913 (N_3913,N_2589,N_3167);
or U3914 (N_3914,N_3121,N_3041);
nor U3915 (N_3915,N_2706,N_2964);
or U3916 (N_3916,N_3095,N_2891);
nand U3917 (N_3917,N_2584,N_2474);
nand U3918 (N_3918,N_2888,N_2518);
and U3919 (N_3919,N_2454,N_3112);
nor U3920 (N_3920,N_2455,N_2879);
xor U3921 (N_3921,N_3164,N_3045);
nand U3922 (N_3922,N_2826,N_2409);
and U3923 (N_3923,N_2668,N_2706);
nand U3924 (N_3924,N_3039,N_2587);
and U3925 (N_3925,N_2554,N_2715);
nor U3926 (N_3926,N_3135,N_2787);
and U3927 (N_3927,N_2739,N_2759);
nand U3928 (N_3928,N_2579,N_2708);
or U3929 (N_3929,N_3037,N_3065);
and U3930 (N_3930,N_2873,N_2838);
and U3931 (N_3931,N_2767,N_2671);
or U3932 (N_3932,N_2549,N_2568);
or U3933 (N_3933,N_2617,N_2913);
and U3934 (N_3934,N_2528,N_2915);
or U3935 (N_3935,N_3119,N_2977);
nor U3936 (N_3936,N_2517,N_2908);
xnor U3937 (N_3937,N_2965,N_2797);
nand U3938 (N_3938,N_2672,N_2497);
xnor U3939 (N_3939,N_2744,N_3013);
nand U3940 (N_3940,N_2916,N_2704);
xor U3941 (N_3941,N_2575,N_2775);
or U3942 (N_3942,N_3158,N_2781);
nor U3943 (N_3943,N_2501,N_3053);
nand U3944 (N_3944,N_2619,N_2762);
nor U3945 (N_3945,N_3103,N_2872);
and U3946 (N_3946,N_2443,N_2760);
nor U3947 (N_3947,N_2652,N_3197);
xor U3948 (N_3948,N_2909,N_3108);
or U3949 (N_3949,N_2797,N_3007);
and U3950 (N_3950,N_2690,N_2628);
or U3951 (N_3951,N_3146,N_2863);
or U3952 (N_3952,N_2428,N_3126);
nand U3953 (N_3953,N_2871,N_2729);
or U3954 (N_3954,N_2995,N_3132);
nand U3955 (N_3955,N_2500,N_2455);
nor U3956 (N_3956,N_2990,N_2403);
xnor U3957 (N_3957,N_2969,N_3083);
or U3958 (N_3958,N_3070,N_2600);
xor U3959 (N_3959,N_2782,N_2585);
and U3960 (N_3960,N_2998,N_2655);
xnor U3961 (N_3961,N_2803,N_2849);
xor U3962 (N_3962,N_2422,N_3066);
nor U3963 (N_3963,N_2540,N_2759);
or U3964 (N_3964,N_2538,N_3088);
or U3965 (N_3965,N_2729,N_3165);
nor U3966 (N_3966,N_2909,N_3054);
nand U3967 (N_3967,N_2905,N_3138);
and U3968 (N_3968,N_2746,N_3035);
xor U3969 (N_3969,N_3098,N_2459);
xnor U3970 (N_3970,N_2759,N_2588);
and U3971 (N_3971,N_2937,N_2576);
nor U3972 (N_3972,N_2500,N_2646);
nor U3973 (N_3973,N_2999,N_3169);
xnor U3974 (N_3974,N_2811,N_2912);
xnor U3975 (N_3975,N_2846,N_2825);
xnor U3976 (N_3976,N_3125,N_2728);
nor U3977 (N_3977,N_2570,N_3048);
nor U3978 (N_3978,N_3014,N_2987);
or U3979 (N_3979,N_3199,N_2808);
and U3980 (N_3980,N_2876,N_2412);
nand U3981 (N_3981,N_2839,N_2968);
or U3982 (N_3982,N_2423,N_3163);
nand U3983 (N_3983,N_3041,N_2464);
or U3984 (N_3984,N_2609,N_2665);
xor U3985 (N_3985,N_2592,N_2577);
xnor U3986 (N_3986,N_2408,N_2945);
and U3987 (N_3987,N_2524,N_2811);
xor U3988 (N_3988,N_2913,N_2418);
nand U3989 (N_3989,N_2942,N_2514);
nor U3990 (N_3990,N_2564,N_3129);
or U3991 (N_3991,N_2474,N_2463);
xor U3992 (N_3992,N_2400,N_2743);
nand U3993 (N_3993,N_3102,N_2849);
xor U3994 (N_3994,N_2402,N_2519);
nand U3995 (N_3995,N_2961,N_3050);
xor U3996 (N_3996,N_3117,N_2802);
or U3997 (N_3997,N_3075,N_3158);
or U3998 (N_3998,N_2975,N_2938);
nand U3999 (N_3999,N_3148,N_2859);
or U4000 (N_4000,N_3688,N_3339);
or U4001 (N_4001,N_3643,N_3969);
xnor U4002 (N_4002,N_3592,N_3202);
nor U4003 (N_4003,N_3956,N_3576);
nor U4004 (N_4004,N_3776,N_3857);
nand U4005 (N_4005,N_3500,N_3660);
or U4006 (N_4006,N_3303,N_3779);
and U4007 (N_4007,N_3685,N_3760);
xor U4008 (N_4008,N_3567,N_3447);
or U4009 (N_4009,N_3542,N_3423);
xor U4010 (N_4010,N_3644,N_3413);
xor U4011 (N_4011,N_3568,N_3613);
and U4012 (N_4012,N_3392,N_3931);
nand U4013 (N_4013,N_3754,N_3965);
and U4014 (N_4014,N_3970,N_3813);
nand U4015 (N_4015,N_3269,N_3878);
or U4016 (N_4016,N_3256,N_3564);
nor U4017 (N_4017,N_3422,N_3680);
nand U4018 (N_4018,N_3234,N_3980);
and U4019 (N_4019,N_3571,N_3844);
or U4020 (N_4020,N_3839,N_3597);
nand U4021 (N_4021,N_3694,N_3595);
and U4022 (N_4022,N_3549,N_3376);
and U4023 (N_4023,N_3848,N_3274);
nand U4024 (N_4024,N_3212,N_3792);
nor U4025 (N_4025,N_3273,N_3229);
and U4026 (N_4026,N_3559,N_3448);
and U4027 (N_4027,N_3768,N_3890);
nor U4028 (N_4028,N_3535,N_3762);
nand U4029 (N_4029,N_3979,N_3245);
and U4030 (N_4030,N_3489,N_3582);
xnor U4031 (N_4031,N_3652,N_3203);
nand U4032 (N_4032,N_3615,N_3524);
xor U4033 (N_4033,N_3424,N_3835);
nor U4034 (N_4034,N_3976,N_3278);
nand U4035 (N_4035,N_3536,N_3991);
and U4036 (N_4036,N_3646,N_3640);
nand U4037 (N_4037,N_3497,N_3521);
nand U4038 (N_4038,N_3636,N_3238);
or U4039 (N_4039,N_3719,N_3226);
and U4040 (N_4040,N_3317,N_3602);
nor U4041 (N_4041,N_3657,N_3903);
or U4042 (N_4042,N_3958,N_3594);
xor U4043 (N_4043,N_3604,N_3606);
xnor U4044 (N_4044,N_3275,N_3201);
nor U4045 (N_4045,N_3838,N_3850);
nand U4046 (N_4046,N_3810,N_3340);
and U4047 (N_4047,N_3794,N_3881);
or U4048 (N_4048,N_3742,N_3371);
nand U4049 (N_4049,N_3369,N_3593);
xnor U4050 (N_4050,N_3924,N_3656);
xor U4051 (N_4051,N_3842,N_3578);
xnor U4052 (N_4052,N_3739,N_3654);
xnor U4053 (N_4053,N_3458,N_3411);
nand U4054 (N_4054,N_3298,N_3505);
nand U4055 (N_4055,N_3953,N_3311);
nor U4056 (N_4056,N_3287,N_3437);
nand U4057 (N_4057,N_3612,N_3486);
or U4058 (N_4058,N_3778,N_3570);
xor U4059 (N_4059,N_3673,N_3892);
nor U4060 (N_4060,N_3511,N_3206);
or U4061 (N_4061,N_3599,N_3966);
nor U4062 (N_4062,N_3459,N_3292);
and U4063 (N_4063,N_3992,N_3475);
and U4064 (N_4064,N_3806,N_3558);
nor U4065 (N_4065,N_3815,N_3331);
and U4066 (N_4066,N_3337,N_3359);
and U4067 (N_4067,N_3638,N_3309);
and U4068 (N_4068,N_3435,N_3253);
and U4069 (N_4069,N_3741,N_3279);
or U4070 (N_4070,N_3932,N_3951);
and U4071 (N_4071,N_3299,N_3283);
xor U4072 (N_4072,N_3420,N_3560);
nor U4073 (N_4073,N_3682,N_3710);
nor U4074 (N_4074,N_3323,N_3538);
or U4075 (N_4075,N_3978,N_3734);
or U4076 (N_4076,N_3623,N_3733);
xor U4077 (N_4077,N_3215,N_3313);
nand U4078 (N_4078,N_3277,N_3596);
xnor U4079 (N_4079,N_3616,N_3817);
nor U4080 (N_4080,N_3907,N_3666);
xnor U4081 (N_4081,N_3709,N_3508);
and U4082 (N_4082,N_3282,N_3659);
and U4083 (N_4083,N_3669,N_3391);
or U4084 (N_4084,N_3429,N_3876);
xor U4085 (N_4085,N_3946,N_3672);
nand U4086 (N_4086,N_3565,N_3374);
nor U4087 (N_4087,N_3355,N_3952);
xor U4088 (N_4088,N_3987,N_3745);
nand U4089 (N_4089,N_3783,N_3889);
nand U4090 (N_4090,N_3626,N_3860);
and U4091 (N_4091,N_3761,N_3703);
nor U4092 (N_4092,N_3380,N_3388);
nor U4093 (N_4093,N_3352,N_3863);
and U4094 (N_4094,N_3994,N_3950);
xnor U4095 (N_4095,N_3771,N_3905);
and U4096 (N_4096,N_3985,N_3763);
or U4097 (N_4097,N_3796,N_3875);
xor U4098 (N_4098,N_3302,N_3457);
xor U4099 (N_4099,N_3552,N_3822);
nand U4100 (N_4100,N_3514,N_3324);
nand U4101 (N_4101,N_3642,N_3715);
nor U4102 (N_4102,N_3605,N_3533);
and U4103 (N_4103,N_3264,N_3356);
or U4104 (N_4104,N_3713,N_3653);
nor U4105 (N_4105,N_3820,N_3327);
xor U4106 (N_4106,N_3921,N_3743);
nand U4107 (N_4107,N_3845,N_3320);
nand U4108 (N_4108,N_3444,N_3364);
and U4109 (N_4109,N_3419,N_3989);
and U4110 (N_4110,N_3827,N_3479);
xnor U4111 (N_4111,N_3284,N_3528);
nand U4112 (N_4112,N_3716,N_3230);
xnor U4113 (N_4113,N_3569,N_3221);
nand U4114 (N_4114,N_3865,N_3790);
and U4115 (N_4115,N_3481,N_3516);
xor U4116 (N_4116,N_3214,N_3466);
nand U4117 (N_4117,N_3454,N_3488);
xor U4118 (N_4118,N_3579,N_3756);
or U4119 (N_4119,N_3498,N_3543);
or U4120 (N_4120,N_3793,N_3891);
or U4121 (N_4121,N_3825,N_3333);
xnor U4122 (N_4122,N_3919,N_3577);
nor U4123 (N_4123,N_3607,N_3834);
and U4124 (N_4124,N_3740,N_3681);
xor U4125 (N_4125,N_3859,N_3861);
xnor U4126 (N_4126,N_3831,N_3665);
nor U4127 (N_4127,N_3765,N_3699);
or U4128 (N_4128,N_3233,N_3769);
nand U4129 (N_4129,N_3809,N_3248);
or U4130 (N_4130,N_3799,N_3310);
or U4131 (N_4131,N_3651,N_3718);
or U4132 (N_4132,N_3684,N_3727);
nand U4133 (N_4133,N_3780,N_3237);
nand U4134 (N_4134,N_3294,N_3295);
and U4135 (N_4135,N_3400,N_3736);
nor U4136 (N_4136,N_3496,N_3749);
or U4137 (N_4137,N_3353,N_3583);
xor U4138 (N_4138,N_3971,N_3276);
nand U4139 (N_4139,N_3668,N_3322);
nor U4140 (N_4140,N_3770,N_3618);
nor U4141 (N_4141,N_3897,N_3895);
nor U4142 (N_4142,N_3686,N_3735);
nand U4143 (N_4143,N_3480,N_3963);
nor U4144 (N_4144,N_3416,N_3955);
or U4145 (N_4145,N_3633,N_3883);
xnor U4146 (N_4146,N_3463,N_3590);
or U4147 (N_4147,N_3401,N_3887);
xor U4148 (N_4148,N_3625,N_3574);
nor U4149 (N_4149,N_3246,N_3397);
and U4150 (N_4150,N_3909,N_3812);
nand U4151 (N_4151,N_3724,N_3344);
nor U4152 (N_4152,N_3412,N_3960);
nor U4153 (N_4153,N_3720,N_3922);
and U4154 (N_4154,N_3798,N_3531);
nor U4155 (N_4155,N_3473,N_3414);
nand U4156 (N_4156,N_3930,N_3873);
xnor U4157 (N_4157,N_3433,N_3336);
and U4158 (N_4158,N_3872,N_3707);
nor U4159 (N_4159,N_3689,N_3774);
or U4160 (N_4160,N_3426,N_3787);
nor U4161 (N_4161,N_3959,N_3649);
and U4162 (N_4162,N_3477,N_3772);
nand U4163 (N_4163,N_3990,N_3485);
xor U4164 (N_4164,N_3676,N_3841);
xor U4165 (N_4165,N_3675,N_3914);
xor U4166 (N_4166,N_3972,N_3587);
nand U4167 (N_4167,N_3510,N_3241);
xor U4168 (N_4168,N_3418,N_3512);
and U4169 (N_4169,N_3244,N_3807);
or U4170 (N_4170,N_3301,N_3691);
or U4171 (N_4171,N_3445,N_3517);
and U4172 (N_4172,N_3847,N_3572);
xnor U4173 (N_4173,N_3884,N_3777);
nand U4174 (N_4174,N_3826,N_3236);
or U4175 (N_4175,N_3375,N_3213);
nand U4176 (N_4176,N_3291,N_3258);
or U4177 (N_4177,N_3630,N_3679);
xor U4178 (N_4178,N_3254,N_3462);
or U4179 (N_4179,N_3453,N_3266);
nand U4180 (N_4180,N_3701,N_3757);
nor U4181 (N_4181,N_3526,N_3286);
xor U4182 (N_4182,N_3967,N_3728);
nand U4183 (N_4183,N_3936,N_3923);
and U4184 (N_4184,N_3281,N_3853);
nor U4185 (N_4185,N_3747,N_3677);
and U4186 (N_4186,N_3372,N_3941);
nor U4187 (N_4187,N_3641,N_3661);
nand U4188 (N_4188,N_3219,N_3854);
or U4189 (N_4189,N_3732,N_3316);
and U4190 (N_4190,N_3986,N_3947);
nand U4191 (N_4191,N_3797,N_3671);
xnor U4192 (N_4192,N_3746,N_3483);
nor U4193 (N_4193,N_3363,N_3598);
nor U4194 (N_4194,N_3289,N_3998);
xnor U4195 (N_4195,N_3628,N_3823);
nor U4196 (N_4196,N_3920,N_3490);
nor U4197 (N_4197,N_3252,N_3929);
or U4198 (N_4198,N_3288,N_3280);
nor U4199 (N_4199,N_3441,N_3629);
or U4200 (N_4200,N_3655,N_3984);
xnor U4201 (N_4201,N_3900,N_3525);
or U4202 (N_4202,N_3545,N_3390);
xor U4203 (N_4203,N_3999,N_3725);
or U4204 (N_4204,N_3243,N_3239);
xnor U4205 (N_4205,N_3753,N_3621);
xnor U4206 (N_4206,N_3700,N_3619);
nand U4207 (N_4207,N_3635,N_3415);
nand U4208 (N_4208,N_3381,N_3436);
xor U4209 (N_4209,N_3405,N_3886);
nand U4210 (N_4210,N_3818,N_3804);
or U4211 (N_4211,N_3370,N_3648);
and U4212 (N_4212,N_3235,N_3620);
nor U4213 (N_4213,N_3232,N_3901);
or U4214 (N_4214,N_3529,N_3982);
nor U4215 (N_4215,N_3730,N_3431);
and U4216 (N_4216,N_3404,N_3696);
nand U4217 (N_4217,N_3764,N_3326);
xnor U4218 (N_4218,N_3911,N_3870);
xnor U4219 (N_4219,N_3662,N_3819);
nor U4220 (N_4220,N_3711,N_3358);
xor U4221 (N_4221,N_3474,N_3603);
xnor U4222 (N_4222,N_3383,N_3968);
nand U4223 (N_4223,N_3240,N_3801);
and U4224 (N_4224,N_3504,N_3609);
and U4225 (N_4225,N_3446,N_3611);
xnor U4226 (N_4226,N_3908,N_3544);
nand U4227 (N_4227,N_3365,N_3726);
xnor U4228 (N_4228,N_3904,N_3555);
nand U4229 (N_4229,N_3785,N_3428);
or U4230 (N_4230,N_3268,N_3407);
or U4231 (N_4231,N_3906,N_3974);
nand U4232 (N_4232,N_3962,N_3335);
or U4233 (N_4233,N_3341,N_3805);
or U4234 (N_4234,N_3403,N_3692);
or U4235 (N_4235,N_3250,N_3846);
nand U4236 (N_4236,N_3537,N_3231);
nand U4237 (N_4237,N_3386,N_3518);
or U4238 (N_4238,N_3200,N_3484);
or U4239 (N_4239,N_3639,N_3396);
nor U4240 (N_4240,N_3981,N_3836);
and U4241 (N_4241,N_3265,N_3223);
xor U4242 (N_4242,N_3803,N_3634);
nor U4243 (N_4243,N_3297,N_3750);
nand U4244 (N_4244,N_3402,N_3464);
xor U4245 (N_4245,N_3362,N_3357);
nor U4246 (N_4246,N_3430,N_3210);
and U4247 (N_4247,N_3385,N_3589);
nor U4248 (N_4248,N_3548,N_3561);
xor U4249 (N_4249,N_3434,N_3714);
nand U4250 (N_4250,N_3880,N_3964);
or U4251 (N_4251,N_3751,N_3328);
nor U4252 (N_4252,N_3916,N_3285);
or U4253 (N_4253,N_3368,N_3949);
nor U4254 (N_4254,N_3584,N_3491);
or U4255 (N_4255,N_3408,N_3262);
nor U4256 (N_4256,N_3759,N_3722);
nand U4257 (N_4257,N_3993,N_3670);
xor U4258 (N_4258,N_3678,N_3440);
nand U4259 (N_4259,N_3821,N_3476);
nor U4260 (N_4260,N_3926,N_3373);
and U4261 (N_4261,N_3915,N_3347);
or U4262 (N_4262,N_3314,N_3553);
or U4263 (N_4263,N_3389,N_3443);
nand U4264 (N_4264,N_3896,N_3781);
nand U4265 (N_4265,N_3351,N_3933);
nand U4266 (N_4266,N_3290,N_3866);
nor U4267 (N_4267,N_3910,N_3871);
and U4268 (N_4268,N_3755,N_3855);
nor U4269 (N_4269,N_3867,N_3257);
xor U4270 (N_4270,N_3329,N_3338);
nor U4271 (N_4271,N_3957,N_3717);
or U4272 (N_4272,N_3575,N_3918);
or U4273 (N_4273,N_3708,N_3706);
xnor U4274 (N_4274,N_3468,N_3631);
nor U4275 (N_4275,N_3218,N_3997);
and U4276 (N_4276,N_3507,N_3346);
nand U4277 (N_4277,N_3767,N_3738);
nor U4278 (N_4278,N_3697,N_3208);
and U4279 (N_4279,N_3687,N_3852);
or U4280 (N_4280,N_3869,N_3795);
xor U4281 (N_4281,N_3387,N_3345);
nand U4282 (N_4282,N_3472,N_3800);
xnor U4283 (N_4283,N_3948,N_3913);
nor U4284 (N_4284,N_3541,N_3493);
xnor U4285 (N_4285,N_3249,N_3349);
or U4286 (N_4286,N_3379,N_3455);
nor U4287 (N_4287,N_3554,N_3220);
nand U4288 (N_4288,N_3406,N_3366);
nand U4289 (N_4289,N_3945,N_3829);
or U4290 (N_4290,N_3306,N_3450);
or U4291 (N_4291,N_3704,N_3944);
and U4292 (N_4292,N_3874,N_3608);
xnor U4293 (N_4293,N_3752,N_3983);
nand U4294 (N_4294,N_3293,N_3833);
xor U4295 (N_4295,N_3766,N_3384);
nand U4296 (N_4296,N_3942,N_3432);
and U4297 (N_4297,N_3744,N_3674);
or U4298 (N_4298,N_3858,N_3530);
xnor U4299 (N_4299,N_3225,N_3478);
and U4300 (N_4300,N_3995,N_3438);
and U4301 (N_4301,N_3784,N_3624);
nand U4302 (N_4302,N_3361,N_3378);
nor U4303 (N_4303,N_3562,N_3399);
nor U4304 (N_4304,N_3690,N_3503);
and U4305 (N_4305,N_3263,N_3988);
or U4306 (N_4306,N_3260,N_3614);
nand U4307 (N_4307,N_3216,N_3856);
nor U4308 (N_4308,N_3885,N_3843);
nor U4309 (N_4309,N_3494,N_3581);
xor U4310 (N_4310,N_3786,N_3532);
nor U4311 (N_4311,N_3695,N_3601);
nand U4312 (N_4312,N_3712,N_3811);
nand U4313 (N_4313,N_3318,N_3556);
nand U4314 (N_4314,N_3664,N_3927);
or U4315 (N_4315,N_3591,N_3632);
nor U4316 (N_4316,N_3830,N_3802);
nand U4317 (N_4317,N_3622,N_3702);
xnor U4318 (N_4318,N_3460,N_3224);
nand U4319 (N_4319,N_3663,N_3816);
or U4320 (N_4320,N_3205,N_3315);
nor U4321 (N_4321,N_3456,N_3247);
or U4322 (N_4322,N_3814,N_3513);
xor U4323 (N_4323,N_3394,N_3502);
nand U4324 (N_4324,N_3271,N_3332);
or U4325 (N_4325,N_3954,N_3585);
nor U4326 (N_4326,N_3996,N_3395);
nand U4327 (N_4327,N_3773,N_3312);
and U4328 (N_4328,N_3627,N_3840);
nand U4329 (N_4329,N_3207,N_3851);
or U4330 (N_4330,N_3228,N_3360);
xnor U4331 (N_4331,N_3350,N_3849);
xor U4332 (N_4332,N_3393,N_3487);
and U4333 (N_4333,N_3540,N_3705);
or U4334 (N_4334,N_3442,N_3547);
nor U4335 (N_4335,N_3469,N_3586);
nor U4336 (N_4336,N_3367,N_3398);
and U4337 (N_4337,N_3471,N_3452);
and U4338 (N_4338,N_3534,N_3617);
xnor U4339 (N_4339,N_3334,N_3520);
xor U4340 (N_4340,N_3917,N_3894);
and U4341 (N_4341,N_3343,N_3975);
or U4342 (N_4342,N_3600,N_3551);
nand U4343 (N_4343,N_3898,N_3828);
nor U4344 (N_4344,N_3864,N_3211);
and U4345 (N_4345,N_3300,N_3934);
and U4346 (N_4346,N_3566,N_3342);
nand U4347 (N_4347,N_3482,N_3698);
xnor U4348 (N_4348,N_3637,N_3527);
nor U4349 (N_4349,N_3449,N_3425);
xnor U4350 (N_4350,N_3251,N_3515);
xnor U4351 (N_4351,N_3647,N_3325);
xnor U4352 (N_4352,N_3204,N_3775);
nand U4353 (N_4353,N_3658,N_3499);
or U4354 (N_4354,N_3808,N_3588);
or U4355 (N_4355,N_3506,N_3902);
xnor U4356 (N_4356,N_3409,N_3882);
or U4357 (N_4357,N_3563,N_3261);
nor U4358 (N_4358,N_3888,N_3550);
xnor U4359 (N_4359,N_3935,N_3321);
xnor U4360 (N_4360,N_3267,N_3937);
nand U4361 (N_4361,N_3421,N_3319);
and U4362 (N_4362,N_3573,N_3862);
or U4363 (N_4363,N_3305,N_3308);
xnor U4364 (N_4364,N_3439,N_3354);
nor U4365 (N_4365,N_3721,N_3522);
and U4366 (N_4366,N_3645,N_3961);
nand U4367 (N_4367,N_3973,N_3417);
nand U4368 (N_4368,N_3451,N_3272);
or U4369 (N_4369,N_3899,N_3255);
and U4370 (N_4370,N_3693,N_3877);
nand U4371 (N_4371,N_3667,N_3940);
nand U4372 (N_4372,N_3879,N_3467);
or U4373 (N_4373,N_3546,N_3330);
and U4374 (N_4374,N_3791,N_3461);
nand U4375 (N_4375,N_3509,N_3209);
xor U4376 (N_4376,N_3492,N_3242);
or U4377 (N_4377,N_3382,N_3683);
and U4378 (N_4378,N_3729,N_3938);
nor U4379 (N_4379,N_3939,N_3304);
and U4380 (N_4380,N_3788,N_3580);
nand U4381 (N_4381,N_3610,N_3377);
and U4382 (N_4382,N_3758,N_3470);
xnor U4383 (N_4383,N_3523,N_3893);
nor U4384 (N_4384,N_3227,N_3465);
nand U4385 (N_4385,N_3737,N_3519);
nand U4386 (N_4386,N_3259,N_3943);
xor U4387 (N_4387,N_3539,N_3868);
xnor U4388 (N_4388,N_3650,N_3270);
nor U4389 (N_4389,N_3217,N_3222);
or U4390 (N_4390,N_3348,N_3789);
nand U4391 (N_4391,N_3495,N_3912);
nor U4392 (N_4392,N_3501,N_3782);
or U4393 (N_4393,N_3824,N_3832);
and U4394 (N_4394,N_3557,N_3925);
nand U4395 (N_4395,N_3723,N_3837);
xnor U4396 (N_4396,N_3427,N_3410);
xor U4397 (N_4397,N_3296,N_3307);
nor U4398 (N_4398,N_3748,N_3731);
xnor U4399 (N_4399,N_3977,N_3928);
or U4400 (N_4400,N_3787,N_3880);
nand U4401 (N_4401,N_3926,N_3299);
xnor U4402 (N_4402,N_3588,N_3269);
nor U4403 (N_4403,N_3568,N_3793);
and U4404 (N_4404,N_3828,N_3958);
and U4405 (N_4405,N_3330,N_3998);
or U4406 (N_4406,N_3374,N_3516);
nand U4407 (N_4407,N_3935,N_3748);
or U4408 (N_4408,N_3672,N_3488);
xnor U4409 (N_4409,N_3322,N_3333);
xor U4410 (N_4410,N_3256,N_3442);
nor U4411 (N_4411,N_3236,N_3370);
and U4412 (N_4412,N_3569,N_3917);
or U4413 (N_4413,N_3783,N_3240);
and U4414 (N_4414,N_3228,N_3258);
nand U4415 (N_4415,N_3448,N_3567);
or U4416 (N_4416,N_3567,N_3568);
xnor U4417 (N_4417,N_3868,N_3824);
nand U4418 (N_4418,N_3430,N_3768);
nand U4419 (N_4419,N_3822,N_3848);
xor U4420 (N_4420,N_3758,N_3330);
nor U4421 (N_4421,N_3974,N_3304);
nor U4422 (N_4422,N_3946,N_3548);
nor U4423 (N_4423,N_3288,N_3835);
and U4424 (N_4424,N_3331,N_3258);
or U4425 (N_4425,N_3302,N_3856);
or U4426 (N_4426,N_3536,N_3667);
nor U4427 (N_4427,N_3249,N_3696);
or U4428 (N_4428,N_3831,N_3443);
and U4429 (N_4429,N_3374,N_3809);
and U4430 (N_4430,N_3866,N_3757);
nor U4431 (N_4431,N_3778,N_3647);
nand U4432 (N_4432,N_3457,N_3815);
and U4433 (N_4433,N_3359,N_3322);
nand U4434 (N_4434,N_3381,N_3404);
nand U4435 (N_4435,N_3952,N_3878);
nor U4436 (N_4436,N_3678,N_3340);
or U4437 (N_4437,N_3952,N_3472);
nand U4438 (N_4438,N_3331,N_3431);
xnor U4439 (N_4439,N_3915,N_3264);
nand U4440 (N_4440,N_3251,N_3979);
and U4441 (N_4441,N_3823,N_3436);
or U4442 (N_4442,N_3599,N_3961);
and U4443 (N_4443,N_3611,N_3779);
nor U4444 (N_4444,N_3447,N_3471);
xnor U4445 (N_4445,N_3715,N_3947);
xnor U4446 (N_4446,N_3427,N_3399);
or U4447 (N_4447,N_3890,N_3910);
nand U4448 (N_4448,N_3608,N_3797);
nand U4449 (N_4449,N_3343,N_3520);
and U4450 (N_4450,N_3266,N_3350);
nor U4451 (N_4451,N_3638,N_3468);
nand U4452 (N_4452,N_3354,N_3935);
and U4453 (N_4453,N_3218,N_3695);
xnor U4454 (N_4454,N_3500,N_3525);
xnor U4455 (N_4455,N_3485,N_3282);
or U4456 (N_4456,N_3462,N_3267);
nand U4457 (N_4457,N_3785,N_3304);
and U4458 (N_4458,N_3204,N_3934);
xnor U4459 (N_4459,N_3338,N_3775);
and U4460 (N_4460,N_3551,N_3589);
or U4461 (N_4461,N_3945,N_3549);
nand U4462 (N_4462,N_3754,N_3495);
and U4463 (N_4463,N_3510,N_3529);
and U4464 (N_4464,N_3324,N_3850);
nor U4465 (N_4465,N_3372,N_3978);
nor U4466 (N_4466,N_3354,N_3874);
nor U4467 (N_4467,N_3572,N_3410);
or U4468 (N_4468,N_3790,N_3289);
and U4469 (N_4469,N_3368,N_3841);
and U4470 (N_4470,N_3376,N_3701);
xnor U4471 (N_4471,N_3745,N_3224);
or U4472 (N_4472,N_3826,N_3334);
xor U4473 (N_4473,N_3924,N_3227);
xor U4474 (N_4474,N_3433,N_3706);
nor U4475 (N_4475,N_3341,N_3477);
nor U4476 (N_4476,N_3943,N_3918);
and U4477 (N_4477,N_3530,N_3517);
or U4478 (N_4478,N_3820,N_3365);
and U4479 (N_4479,N_3449,N_3740);
xnor U4480 (N_4480,N_3964,N_3706);
and U4481 (N_4481,N_3217,N_3635);
xor U4482 (N_4482,N_3328,N_3274);
or U4483 (N_4483,N_3813,N_3994);
xor U4484 (N_4484,N_3413,N_3460);
nand U4485 (N_4485,N_3475,N_3808);
and U4486 (N_4486,N_3832,N_3810);
and U4487 (N_4487,N_3265,N_3950);
and U4488 (N_4488,N_3905,N_3871);
and U4489 (N_4489,N_3525,N_3340);
nand U4490 (N_4490,N_3654,N_3706);
or U4491 (N_4491,N_3569,N_3417);
nand U4492 (N_4492,N_3268,N_3961);
xor U4493 (N_4493,N_3421,N_3271);
xor U4494 (N_4494,N_3568,N_3609);
xnor U4495 (N_4495,N_3934,N_3799);
and U4496 (N_4496,N_3966,N_3622);
and U4497 (N_4497,N_3688,N_3247);
or U4498 (N_4498,N_3237,N_3226);
xor U4499 (N_4499,N_3608,N_3514);
or U4500 (N_4500,N_3901,N_3569);
nand U4501 (N_4501,N_3871,N_3606);
nor U4502 (N_4502,N_3722,N_3326);
and U4503 (N_4503,N_3742,N_3609);
or U4504 (N_4504,N_3803,N_3243);
nand U4505 (N_4505,N_3887,N_3236);
or U4506 (N_4506,N_3293,N_3914);
and U4507 (N_4507,N_3544,N_3206);
nor U4508 (N_4508,N_3666,N_3680);
nand U4509 (N_4509,N_3640,N_3441);
nor U4510 (N_4510,N_3778,N_3410);
xor U4511 (N_4511,N_3605,N_3489);
xnor U4512 (N_4512,N_3836,N_3300);
and U4513 (N_4513,N_3817,N_3454);
or U4514 (N_4514,N_3761,N_3478);
and U4515 (N_4515,N_3468,N_3683);
and U4516 (N_4516,N_3572,N_3921);
or U4517 (N_4517,N_3979,N_3339);
or U4518 (N_4518,N_3860,N_3508);
nor U4519 (N_4519,N_3459,N_3320);
nor U4520 (N_4520,N_3258,N_3693);
or U4521 (N_4521,N_3501,N_3491);
and U4522 (N_4522,N_3657,N_3856);
nand U4523 (N_4523,N_3826,N_3206);
nand U4524 (N_4524,N_3958,N_3546);
xnor U4525 (N_4525,N_3303,N_3940);
or U4526 (N_4526,N_3561,N_3733);
xnor U4527 (N_4527,N_3507,N_3254);
xnor U4528 (N_4528,N_3252,N_3766);
xor U4529 (N_4529,N_3554,N_3687);
xor U4530 (N_4530,N_3960,N_3918);
and U4531 (N_4531,N_3206,N_3727);
and U4532 (N_4532,N_3847,N_3442);
nor U4533 (N_4533,N_3689,N_3659);
xor U4534 (N_4534,N_3957,N_3405);
and U4535 (N_4535,N_3882,N_3755);
or U4536 (N_4536,N_3760,N_3345);
nor U4537 (N_4537,N_3234,N_3274);
and U4538 (N_4538,N_3488,N_3752);
nand U4539 (N_4539,N_3543,N_3856);
and U4540 (N_4540,N_3792,N_3608);
xor U4541 (N_4541,N_3938,N_3941);
or U4542 (N_4542,N_3421,N_3600);
or U4543 (N_4543,N_3723,N_3224);
nor U4544 (N_4544,N_3716,N_3488);
nand U4545 (N_4545,N_3655,N_3795);
nor U4546 (N_4546,N_3413,N_3726);
and U4547 (N_4547,N_3626,N_3504);
and U4548 (N_4548,N_3689,N_3390);
nand U4549 (N_4549,N_3971,N_3668);
or U4550 (N_4550,N_3769,N_3901);
or U4551 (N_4551,N_3222,N_3494);
and U4552 (N_4552,N_3639,N_3844);
xnor U4553 (N_4553,N_3255,N_3908);
nor U4554 (N_4554,N_3438,N_3307);
xor U4555 (N_4555,N_3787,N_3219);
nand U4556 (N_4556,N_3207,N_3843);
and U4557 (N_4557,N_3887,N_3716);
xor U4558 (N_4558,N_3223,N_3429);
nor U4559 (N_4559,N_3996,N_3400);
xnor U4560 (N_4560,N_3678,N_3586);
and U4561 (N_4561,N_3615,N_3328);
or U4562 (N_4562,N_3477,N_3729);
and U4563 (N_4563,N_3836,N_3459);
xnor U4564 (N_4564,N_3943,N_3544);
or U4565 (N_4565,N_3456,N_3860);
nand U4566 (N_4566,N_3923,N_3515);
nor U4567 (N_4567,N_3304,N_3617);
nor U4568 (N_4568,N_3571,N_3757);
nand U4569 (N_4569,N_3829,N_3921);
and U4570 (N_4570,N_3497,N_3239);
and U4571 (N_4571,N_3851,N_3891);
nor U4572 (N_4572,N_3381,N_3204);
and U4573 (N_4573,N_3237,N_3473);
nand U4574 (N_4574,N_3763,N_3650);
or U4575 (N_4575,N_3506,N_3454);
and U4576 (N_4576,N_3633,N_3682);
or U4577 (N_4577,N_3636,N_3976);
xnor U4578 (N_4578,N_3598,N_3237);
or U4579 (N_4579,N_3444,N_3525);
xor U4580 (N_4580,N_3707,N_3257);
nor U4581 (N_4581,N_3370,N_3993);
nand U4582 (N_4582,N_3920,N_3552);
or U4583 (N_4583,N_3849,N_3700);
nor U4584 (N_4584,N_3919,N_3688);
nor U4585 (N_4585,N_3635,N_3766);
or U4586 (N_4586,N_3617,N_3332);
or U4587 (N_4587,N_3841,N_3310);
nand U4588 (N_4588,N_3577,N_3725);
and U4589 (N_4589,N_3899,N_3749);
nand U4590 (N_4590,N_3439,N_3916);
nor U4591 (N_4591,N_3970,N_3538);
and U4592 (N_4592,N_3351,N_3346);
or U4593 (N_4593,N_3202,N_3432);
and U4594 (N_4594,N_3428,N_3730);
and U4595 (N_4595,N_3914,N_3959);
nor U4596 (N_4596,N_3444,N_3441);
nand U4597 (N_4597,N_3549,N_3921);
xnor U4598 (N_4598,N_3774,N_3990);
xnor U4599 (N_4599,N_3426,N_3644);
and U4600 (N_4600,N_3494,N_3455);
or U4601 (N_4601,N_3412,N_3885);
nor U4602 (N_4602,N_3366,N_3253);
nand U4603 (N_4603,N_3548,N_3666);
or U4604 (N_4604,N_3927,N_3875);
nor U4605 (N_4605,N_3474,N_3444);
and U4606 (N_4606,N_3890,N_3335);
nor U4607 (N_4607,N_3691,N_3491);
xnor U4608 (N_4608,N_3968,N_3830);
or U4609 (N_4609,N_3305,N_3414);
or U4610 (N_4610,N_3954,N_3511);
nor U4611 (N_4611,N_3654,N_3993);
xnor U4612 (N_4612,N_3432,N_3693);
nor U4613 (N_4613,N_3226,N_3629);
nor U4614 (N_4614,N_3877,N_3686);
nand U4615 (N_4615,N_3783,N_3325);
and U4616 (N_4616,N_3754,N_3562);
xnor U4617 (N_4617,N_3786,N_3456);
xnor U4618 (N_4618,N_3800,N_3810);
nor U4619 (N_4619,N_3225,N_3230);
xnor U4620 (N_4620,N_3282,N_3846);
and U4621 (N_4621,N_3594,N_3803);
or U4622 (N_4622,N_3913,N_3955);
nand U4623 (N_4623,N_3883,N_3643);
nand U4624 (N_4624,N_3972,N_3481);
xor U4625 (N_4625,N_3916,N_3751);
nand U4626 (N_4626,N_3893,N_3966);
or U4627 (N_4627,N_3232,N_3737);
or U4628 (N_4628,N_3295,N_3268);
nand U4629 (N_4629,N_3252,N_3943);
or U4630 (N_4630,N_3585,N_3499);
and U4631 (N_4631,N_3995,N_3367);
xor U4632 (N_4632,N_3353,N_3682);
xnor U4633 (N_4633,N_3610,N_3412);
nand U4634 (N_4634,N_3967,N_3769);
nand U4635 (N_4635,N_3982,N_3682);
and U4636 (N_4636,N_3477,N_3938);
and U4637 (N_4637,N_3226,N_3951);
nand U4638 (N_4638,N_3482,N_3859);
nor U4639 (N_4639,N_3252,N_3700);
xor U4640 (N_4640,N_3434,N_3692);
nand U4641 (N_4641,N_3947,N_3924);
or U4642 (N_4642,N_3930,N_3452);
or U4643 (N_4643,N_3281,N_3576);
xnor U4644 (N_4644,N_3636,N_3231);
and U4645 (N_4645,N_3571,N_3405);
nor U4646 (N_4646,N_3222,N_3735);
nand U4647 (N_4647,N_3679,N_3351);
nor U4648 (N_4648,N_3302,N_3644);
and U4649 (N_4649,N_3950,N_3295);
nor U4650 (N_4650,N_3271,N_3269);
nor U4651 (N_4651,N_3692,N_3763);
nor U4652 (N_4652,N_3877,N_3792);
nor U4653 (N_4653,N_3908,N_3729);
or U4654 (N_4654,N_3439,N_3587);
or U4655 (N_4655,N_3441,N_3881);
or U4656 (N_4656,N_3820,N_3407);
nor U4657 (N_4657,N_3677,N_3678);
nor U4658 (N_4658,N_3521,N_3501);
and U4659 (N_4659,N_3230,N_3552);
nand U4660 (N_4660,N_3469,N_3861);
nor U4661 (N_4661,N_3424,N_3271);
or U4662 (N_4662,N_3575,N_3812);
nand U4663 (N_4663,N_3937,N_3660);
nand U4664 (N_4664,N_3574,N_3337);
and U4665 (N_4665,N_3842,N_3548);
xor U4666 (N_4666,N_3240,N_3241);
nand U4667 (N_4667,N_3363,N_3911);
or U4668 (N_4668,N_3716,N_3574);
nor U4669 (N_4669,N_3977,N_3761);
xnor U4670 (N_4670,N_3420,N_3357);
nand U4671 (N_4671,N_3367,N_3361);
xnor U4672 (N_4672,N_3538,N_3348);
nand U4673 (N_4673,N_3318,N_3814);
or U4674 (N_4674,N_3655,N_3809);
or U4675 (N_4675,N_3763,N_3368);
and U4676 (N_4676,N_3961,N_3721);
or U4677 (N_4677,N_3220,N_3510);
or U4678 (N_4678,N_3433,N_3733);
xor U4679 (N_4679,N_3245,N_3668);
or U4680 (N_4680,N_3303,N_3615);
xnor U4681 (N_4681,N_3722,N_3563);
and U4682 (N_4682,N_3803,N_3343);
xor U4683 (N_4683,N_3758,N_3380);
nand U4684 (N_4684,N_3347,N_3984);
xor U4685 (N_4685,N_3673,N_3493);
and U4686 (N_4686,N_3720,N_3666);
nand U4687 (N_4687,N_3886,N_3258);
xor U4688 (N_4688,N_3605,N_3743);
nand U4689 (N_4689,N_3379,N_3705);
nand U4690 (N_4690,N_3871,N_3634);
and U4691 (N_4691,N_3367,N_3754);
xor U4692 (N_4692,N_3684,N_3586);
and U4693 (N_4693,N_3889,N_3672);
and U4694 (N_4694,N_3832,N_3856);
and U4695 (N_4695,N_3924,N_3380);
nor U4696 (N_4696,N_3734,N_3403);
nand U4697 (N_4697,N_3609,N_3343);
xor U4698 (N_4698,N_3594,N_3325);
or U4699 (N_4699,N_3626,N_3503);
nor U4700 (N_4700,N_3857,N_3624);
and U4701 (N_4701,N_3574,N_3909);
nor U4702 (N_4702,N_3399,N_3715);
or U4703 (N_4703,N_3672,N_3841);
and U4704 (N_4704,N_3403,N_3662);
or U4705 (N_4705,N_3778,N_3425);
and U4706 (N_4706,N_3595,N_3888);
xnor U4707 (N_4707,N_3734,N_3228);
xnor U4708 (N_4708,N_3425,N_3538);
and U4709 (N_4709,N_3508,N_3711);
or U4710 (N_4710,N_3754,N_3269);
nor U4711 (N_4711,N_3359,N_3663);
nand U4712 (N_4712,N_3801,N_3489);
xnor U4713 (N_4713,N_3232,N_3729);
nand U4714 (N_4714,N_3626,N_3209);
and U4715 (N_4715,N_3865,N_3423);
or U4716 (N_4716,N_3459,N_3383);
and U4717 (N_4717,N_3698,N_3938);
xor U4718 (N_4718,N_3605,N_3313);
nor U4719 (N_4719,N_3491,N_3468);
xor U4720 (N_4720,N_3841,N_3207);
or U4721 (N_4721,N_3980,N_3809);
and U4722 (N_4722,N_3898,N_3707);
and U4723 (N_4723,N_3648,N_3769);
nor U4724 (N_4724,N_3894,N_3278);
xnor U4725 (N_4725,N_3890,N_3338);
and U4726 (N_4726,N_3220,N_3271);
nand U4727 (N_4727,N_3404,N_3532);
nor U4728 (N_4728,N_3636,N_3705);
or U4729 (N_4729,N_3383,N_3687);
and U4730 (N_4730,N_3526,N_3681);
nor U4731 (N_4731,N_3461,N_3538);
nand U4732 (N_4732,N_3708,N_3912);
xor U4733 (N_4733,N_3263,N_3361);
xnor U4734 (N_4734,N_3833,N_3837);
or U4735 (N_4735,N_3751,N_3695);
nand U4736 (N_4736,N_3353,N_3846);
or U4737 (N_4737,N_3202,N_3351);
and U4738 (N_4738,N_3429,N_3462);
nor U4739 (N_4739,N_3521,N_3998);
nand U4740 (N_4740,N_3776,N_3356);
nor U4741 (N_4741,N_3769,N_3930);
nand U4742 (N_4742,N_3276,N_3660);
nand U4743 (N_4743,N_3555,N_3356);
nand U4744 (N_4744,N_3831,N_3932);
or U4745 (N_4745,N_3555,N_3612);
or U4746 (N_4746,N_3565,N_3609);
or U4747 (N_4747,N_3425,N_3455);
or U4748 (N_4748,N_3209,N_3387);
nand U4749 (N_4749,N_3867,N_3226);
nor U4750 (N_4750,N_3600,N_3406);
nor U4751 (N_4751,N_3977,N_3934);
and U4752 (N_4752,N_3847,N_3840);
nand U4753 (N_4753,N_3907,N_3978);
nor U4754 (N_4754,N_3530,N_3450);
nor U4755 (N_4755,N_3281,N_3396);
or U4756 (N_4756,N_3276,N_3746);
and U4757 (N_4757,N_3668,N_3562);
xor U4758 (N_4758,N_3463,N_3406);
nand U4759 (N_4759,N_3749,N_3350);
xor U4760 (N_4760,N_3427,N_3491);
nand U4761 (N_4761,N_3465,N_3598);
and U4762 (N_4762,N_3895,N_3549);
nor U4763 (N_4763,N_3387,N_3455);
xnor U4764 (N_4764,N_3532,N_3392);
and U4765 (N_4765,N_3912,N_3798);
nor U4766 (N_4766,N_3438,N_3991);
nor U4767 (N_4767,N_3583,N_3524);
nand U4768 (N_4768,N_3747,N_3915);
xnor U4769 (N_4769,N_3705,N_3702);
or U4770 (N_4770,N_3904,N_3852);
nor U4771 (N_4771,N_3825,N_3634);
or U4772 (N_4772,N_3489,N_3867);
nand U4773 (N_4773,N_3983,N_3744);
or U4774 (N_4774,N_3586,N_3430);
xnor U4775 (N_4775,N_3787,N_3608);
or U4776 (N_4776,N_3729,N_3441);
or U4777 (N_4777,N_3891,N_3828);
nand U4778 (N_4778,N_3239,N_3232);
nor U4779 (N_4779,N_3889,N_3846);
nor U4780 (N_4780,N_3250,N_3556);
and U4781 (N_4781,N_3818,N_3671);
xnor U4782 (N_4782,N_3672,N_3735);
nand U4783 (N_4783,N_3771,N_3236);
or U4784 (N_4784,N_3905,N_3417);
and U4785 (N_4785,N_3801,N_3669);
xnor U4786 (N_4786,N_3788,N_3377);
and U4787 (N_4787,N_3262,N_3412);
nand U4788 (N_4788,N_3953,N_3214);
or U4789 (N_4789,N_3450,N_3430);
or U4790 (N_4790,N_3851,N_3876);
nor U4791 (N_4791,N_3953,N_3207);
xor U4792 (N_4792,N_3991,N_3392);
nor U4793 (N_4793,N_3753,N_3516);
xnor U4794 (N_4794,N_3964,N_3607);
and U4795 (N_4795,N_3594,N_3622);
xnor U4796 (N_4796,N_3896,N_3702);
nor U4797 (N_4797,N_3868,N_3503);
nand U4798 (N_4798,N_3257,N_3768);
or U4799 (N_4799,N_3979,N_3680);
xnor U4800 (N_4800,N_4080,N_4263);
and U4801 (N_4801,N_4567,N_4769);
and U4802 (N_4802,N_4173,N_4762);
nand U4803 (N_4803,N_4752,N_4755);
xnor U4804 (N_4804,N_4469,N_4262);
or U4805 (N_4805,N_4373,N_4783);
nor U4806 (N_4806,N_4682,N_4181);
xor U4807 (N_4807,N_4668,N_4000);
nand U4808 (N_4808,N_4369,N_4447);
or U4809 (N_4809,N_4104,N_4127);
nor U4810 (N_4810,N_4652,N_4163);
nor U4811 (N_4811,N_4098,N_4674);
nand U4812 (N_4812,N_4568,N_4406);
or U4813 (N_4813,N_4093,N_4663);
nand U4814 (N_4814,N_4362,N_4525);
and U4815 (N_4815,N_4251,N_4595);
or U4816 (N_4816,N_4268,N_4639);
nand U4817 (N_4817,N_4150,N_4267);
nor U4818 (N_4818,N_4110,N_4403);
and U4819 (N_4819,N_4074,N_4596);
nand U4820 (N_4820,N_4059,N_4272);
nand U4821 (N_4821,N_4332,N_4113);
and U4822 (N_4822,N_4408,N_4587);
or U4823 (N_4823,N_4258,N_4256);
nand U4824 (N_4824,N_4294,N_4685);
nand U4825 (N_4825,N_4271,N_4358);
nand U4826 (N_4826,N_4288,N_4348);
and U4827 (N_4827,N_4095,N_4419);
and U4828 (N_4828,N_4243,N_4437);
xor U4829 (N_4829,N_4515,N_4784);
xor U4830 (N_4830,N_4052,N_4002);
or U4831 (N_4831,N_4790,N_4625);
and U4832 (N_4832,N_4201,N_4139);
and U4833 (N_4833,N_4751,N_4363);
nor U4834 (N_4834,N_4791,N_4314);
and U4835 (N_4835,N_4505,N_4149);
or U4836 (N_4836,N_4577,N_4609);
and U4837 (N_4837,N_4213,N_4431);
nand U4838 (N_4838,N_4073,N_4022);
or U4839 (N_4839,N_4683,N_4313);
or U4840 (N_4840,N_4510,N_4232);
nor U4841 (N_4841,N_4013,N_4071);
xnor U4842 (N_4842,N_4130,N_4455);
nor U4843 (N_4843,N_4266,N_4666);
or U4844 (N_4844,N_4100,N_4675);
nand U4845 (N_4845,N_4659,N_4296);
and U4846 (N_4846,N_4055,N_4318);
nor U4847 (N_4847,N_4005,N_4562);
or U4848 (N_4848,N_4028,N_4215);
xor U4849 (N_4849,N_4295,N_4043);
nand U4850 (N_4850,N_4621,N_4643);
nand U4851 (N_4851,N_4153,N_4338);
xor U4852 (N_4852,N_4383,N_4731);
and U4853 (N_4853,N_4223,N_4696);
or U4854 (N_4854,N_4786,N_4399);
or U4855 (N_4855,N_4367,N_4698);
and U4856 (N_4856,N_4216,N_4617);
nand U4857 (N_4857,N_4774,N_4514);
nand U4858 (N_4858,N_4671,N_4670);
or U4859 (N_4859,N_4361,N_4550);
or U4860 (N_4860,N_4404,N_4753);
xor U4861 (N_4861,N_4046,N_4465);
or U4862 (N_4862,N_4270,N_4307);
and U4863 (N_4863,N_4390,N_4584);
or U4864 (N_4864,N_4261,N_4182);
or U4865 (N_4865,N_4311,N_4166);
nand U4866 (N_4866,N_4082,N_4772);
nand U4867 (N_4867,N_4773,N_4047);
xor U4868 (N_4868,N_4351,N_4021);
xnor U4869 (N_4869,N_4661,N_4347);
nand U4870 (N_4870,N_4344,N_4102);
or U4871 (N_4871,N_4247,N_4170);
and U4872 (N_4872,N_4077,N_4282);
and U4873 (N_4873,N_4560,N_4426);
nand U4874 (N_4874,N_4320,N_4044);
and U4875 (N_4875,N_4356,N_4045);
or U4876 (N_4876,N_4602,N_4694);
and U4877 (N_4877,N_4716,N_4407);
nand U4878 (N_4878,N_4205,N_4548);
or U4879 (N_4879,N_4741,N_4248);
or U4880 (N_4880,N_4544,N_4711);
nor U4881 (N_4881,N_4039,N_4765);
nor U4882 (N_4882,N_4474,N_4192);
or U4883 (N_4883,N_4637,N_4485);
and U4884 (N_4884,N_4576,N_4687);
or U4885 (N_4885,N_4375,N_4580);
nor U4886 (N_4886,N_4276,N_4143);
or U4887 (N_4887,N_4635,N_4309);
nor U4888 (N_4888,N_4597,N_4789);
nand U4889 (N_4889,N_4012,N_4357);
or U4890 (N_4890,N_4747,N_4487);
or U4891 (N_4891,N_4412,N_4532);
nand U4892 (N_4892,N_4334,N_4520);
nand U4893 (N_4893,N_4224,N_4122);
or U4894 (N_4894,N_4345,N_4691);
xor U4895 (N_4895,N_4323,N_4036);
and U4896 (N_4896,N_4700,N_4780);
nor U4897 (N_4897,N_4148,N_4193);
and U4898 (N_4898,N_4027,N_4582);
nor U4899 (N_4899,N_4537,N_4647);
or U4900 (N_4900,N_4624,N_4417);
nor U4901 (N_4901,N_4655,N_4759);
or U4902 (N_4902,N_4316,N_4608);
nor U4903 (N_4903,N_4079,N_4340);
or U4904 (N_4904,N_4421,N_4598);
or U4905 (N_4905,N_4535,N_4391);
or U4906 (N_4906,N_4226,N_4440);
xor U4907 (N_4907,N_4008,N_4425);
xor U4908 (N_4908,N_4023,N_4557);
nand U4909 (N_4909,N_4007,N_4057);
nor U4910 (N_4910,N_4255,N_4086);
nand U4911 (N_4911,N_4128,N_4191);
nor U4912 (N_4912,N_4650,N_4371);
or U4913 (N_4913,N_4135,N_4385);
or U4914 (N_4914,N_4556,N_4062);
or U4915 (N_4915,N_4709,N_4402);
nand U4916 (N_4916,N_4350,N_4764);
nand U4917 (N_4917,N_4105,N_4214);
xnor U4918 (N_4918,N_4676,N_4010);
nor U4919 (N_4919,N_4502,N_4614);
and U4920 (N_4920,N_4491,N_4626);
and U4921 (N_4921,N_4378,N_4591);
and U4922 (N_4922,N_4152,N_4068);
or U4923 (N_4923,N_4097,N_4689);
and U4924 (N_4924,N_4497,N_4114);
or U4925 (N_4925,N_4111,N_4604);
and U4926 (N_4926,N_4457,N_4481);
xnor U4927 (N_4927,N_4254,N_4636);
nor U4928 (N_4928,N_4257,N_4706);
nor U4929 (N_4929,N_4241,N_4631);
xnor U4930 (N_4930,N_4720,N_4579);
or U4931 (N_4931,N_4681,N_4620);
and U4932 (N_4932,N_4667,N_4501);
nor U4933 (N_4933,N_4467,N_4763);
nand U4934 (N_4934,N_4503,N_4066);
or U4935 (N_4935,N_4429,N_4777);
and U4936 (N_4936,N_4418,N_4287);
and U4937 (N_4937,N_4336,N_4414);
nor U4938 (N_4938,N_4710,N_4119);
nor U4939 (N_4939,N_4168,N_4436);
nand U4940 (N_4940,N_4496,N_4517);
or U4941 (N_4941,N_4328,N_4554);
or U4942 (N_4942,N_4209,N_4411);
xnor U4943 (N_4943,N_4032,N_4211);
xnor U4944 (N_4944,N_4592,N_4240);
nand U4945 (N_4945,N_4787,N_4275);
or U4946 (N_4946,N_4398,N_4291);
and U4947 (N_4947,N_4613,N_4743);
or U4948 (N_4948,N_4322,N_4641);
nand U4949 (N_4949,N_4518,N_4574);
nor U4950 (N_4950,N_4793,N_4234);
nand U4951 (N_4951,N_4733,N_4669);
xor U4952 (N_4952,N_4125,N_4569);
or U4953 (N_4953,N_4714,N_4285);
nand U4954 (N_4954,N_4194,N_4078);
or U4955 (N_4955,N_4151,N_4376);
nand U4956 (N_4956,N_4394,N_4767);
and U4957 (N_4957,N_4482,N_4651);
nand U4958 (N_4958,N_4473,N_4237);
nand U4959 (N_4959,N_4730,N_4735);
nor U4960 (N_4960,N_4088,N_4183);
and U4961 (N_4961,N_4728,N_4349);
xnor U4962 (N_4962,N_4795,N_4570);
and U4963 (N_4963,N_4396,N_4754);
nand U4964 (N_4964,N_4472,N_4739);
or U4965 (N_4965,N_4176,N_4297);
and U4966 (N_4966,N_4054,N_4470);
nor U4967 (N_4967,N_4660,N_4638);
or U4968 (N_4968,N_4204,N_4360);
nor U4969 (N_4969,N_4154,N_4413);
xor U4970 (N_4970,N_4600,N_4703);
xor U4971 (N_4971,N_4132,N_4433);
and U4972 (N_4972,N_4265,N_4603);
and U4973 (N_4973,N_4004,N_4409);
nor U4974 (N_4974,N_4033,N_4432);
xnor U4975 (N_4975,N_4372,N_4384);
and U4976 (N_4976,N_4718,N_4355);
and U4977 (N_4977,N_4180,N_4219);
and U4978 (N_4978,N_4280,N_4281);
xnor U4979 (N_4979,N_4623,N_4165);
or U4980 (N_4980,N_4559,N_4513);
and U4981 (N_4981,N_4756,N_4038);
and U4982 (N_4982,N_4476,N_4393);
and U4983 (N_4983,N_4448,N_4317);
or U4984 (N_4984,N_4352,N_4123);
and U4985 (N_4985,N_4616,N_4064);
and U4986 (N_4986,N_4627,N_4222);
xnor U4987 (N_4987,N_4069,N_4306);
nor U4988 (N_4988,N_4583,N_4178);
or U4989 (N_4989,N_4549,N_4329);
nand U4990 (N_4990,N_4003,N_4722);
or U4991 (N_4991,N_4619,N_4680);
nand U4992 (N_4992,N_4654,N_4422);
and U4993 (N_4993,N_4343,N_4662);
or U4994 (N_4994,N_4321,N_4236);
nor U4995 (N_4995,N_4758,N_4277);
nand U4996 (N_4996,N_4504,N_4686);
nand U4997 (N_4997,N_4133,N_4284);
nor U4998 (N_4998,N_4508,N_4629);
and U4999 (N_4999,N_4701,N_4319);
and U5000 (N_5000,N_4239,N_4566);
nand U5001 (N_5001,N_4792,N_4389);
xor U5002 (N_5002,N_4737,N_4342);
nand U5003 (N_5003,N_4492,N_4206);
and U5004 (N_5004,N_4212,N_4512);
nand U5005 (N_5005,N_4415,N_4458);
nor U5006 (N_5006,N_4245,N_4196);
nand U5007 (N_5007,N_4697,N_4279);
nand U5008 (N_5008,N_4386,N_4649);
or U5009 (N_5009,N_4264,N_4161);
nor U5010 (N_5010,N_4142,N_4452);
xnor U5011 (N_5011,N_4109,N_4278);
nand U5012 (N_5012,N_4766,N_4060);
nand U5013 (N_5013,N_4558,N_4541);
nor U5014 (N_5014,N_4781,N_4511);
nand U5015 (N_5015,N_4561,N_4089);
nand U5016 (N_5016,N_4341,N_4692);
nor U5017 (N_5017,N_4218,N_4456);
and U5018 (N_5018,N_4230,N_4203);
nor U5019 (N_5019,N_4157,N_4075);
nand U5020 (N_5020,N_4745,N_4175);
and U5021 (N_5021,N_4030,N_4500);
or U5022 (N_5022,N_4087,N_4040);
nand U5023 (N_5023,N_4308,N_4594);
xnor U5024 (N_5024,N_4672,N_4794);
nand U5025 (N_5025,N_4374,N_4640);
and U5026 (N_5026,N_4782,N_4269);
xor U5027 (N_5027,N_4494,N_4746);
xnor U5028 (N_5028,N_4227,N_4736);
nand U5029 (N_5029,N_4312,N_4395);
and U5030 (N_5030,N_4634,N_4303);
nand U5031 (N_5031,N_4498,N_4615);
nor U5032 (N_5032,N_4612,N_4019);
xnor U5033 (N_5033,N_4785,N_4648);
xnor U5034 (N_5034,N_4656,N_4664);
nand U5035 (N_5035,N_4118,N_4590);
nor U5036 (N_5036,N_4547,N_4162);
nand U5037 (N_5037,N_4174,N_4050);
nor U5038 (N_5038,N_4477,N_4124);
xnor U5039 (N_5039,N_4586,N_4724);
or U5040 (N_5040,N_4092,N_4042);
nor U5041 (N_5041,N_4188,N_4011);
or U5042 (N_5042,N_4381,N_4147);
and U5043 (N_5043,N_4072,N_4770);
xor U5044 (N_5044,N_4081,N_4145);
xnor U5045 (N_5045,N_4428,N_4335);
nor U5046 (N_5046,N_4026,N_4677);
and U5047 (N_5047,N_4799,N_4293);
or U5048 (N_5048,N_4665,N_4533);
nand U5049 (N_5049,N_4695,N_4366);
and U5050 (N_5050,N_4434,N_4489);
xnor U5051 (N_5051,N_4144,N_4090);
nand U5052 (N_5052,N_4025,N_4707);
and U5053 (N_5053,N_4259,N_4723);
xor U5054 (N_5054,N_4460,N_4136);
xnor U5055 (N_5055,N_4464,N_4540);
and U5056 (N_5056,N_4037,N_4543);
nand U5057 (N_5057,N_4400,N_4289);
nor U5058 (N_5058,N_4326,N_4775);
nand U5059 (N_5059,N_4286,N_4459);
xnor U5060 (N_5060,N_4009,N_4463);
xor U5061 (N_5061,N_4325,N_4169);
xnor U5062 (N_5062,N_4712,N_4776);
and U5063 (N_5063,N_4014,N_4611);
or U5064 (N_5064,N_4601,N_4717);
nand U5065 (N_5065,N_4462,N_4186);
nand U5066 (N_5066,N_4380,N_4475);
or U5067 (N_5067,N_4779,N_4172);
and U5068 (N_5068,N_4370,N_4461);
nor U5069 (N_5069,N_4006,N_4159);
xor U5070 (N_5070,N_4471,N_4177);
nand U5071 (N_5071,N_4108,N_4673);
and U5072 (N_5072,N_4713,N_4653);
nor U5073 (N_5073,N_4138,N_4112);
or U5074 (N_5074,N_4439,N_4020);
or U5075 (N_5075,N_4091,N_4190);
nor U5076 (N_5076,N_4427,N_4024);
nand U5077 (N_5077,N_4704,N_4410);
or U5078 (N_5078,N_4688,N_4725);
and U5079 (N_5079,N_4690,N_4017);
or U5080 (N_5080,N_4575,N_4678);
or U5081 (N_5081,N_4446,N_4632);
nand U5082 (N_5082,N_4260,N_4484);
nor U5083 (N_5083,N_4238,N_4197);
nand U5084 (N_5084,N_4379,N_4368);
or U5085 (N_5085,N_4516,N_4435);
xor U5086 (N_5086,N_4524,N_4451);
and U5087 (N_5087,N_4480,N_4571);
nor U5088 (N_5088,N_4644,N_4760);
nand U5089 (N_5089,N_4438,N_4750);
nand U5090 (N_5090,N_4063,N_4117);
xor U5091 (N_5091,N_4630,N_4015);
nand U5092 (N_5092,N_4483,N_4140);
or U5093 (N_5093,N_4231,N_4699);
nand U5094 (N_5094,N_4274,N_4053);
xnor U5095 (N_5095,N_4049,N_4103);
nand U5096 (N_5096,N_4198,N_4423);
or U5097 (N_5097,N_4397,N_4096);
and U5098 (N_5098,N_4658,N_4099);
nor U5099 (N_5099,N_4581,N_4522);
or U5100 (N_5100,N_4708,N_4466);
or U5101 (N_5101,N_4521,N_4539);
nor U5102 (N_5102,N_4454,N_4134);
nor U5103 (N_5103,N_4495,N_4573);
and U5104 (N_5104,N_4158,N_4749);
or U5105 (N_5105,N_4221,N_4083);
or U5106 (N_5106,N_4126,N_4300);
or U5107 (N_5107,N_4246,N_4486);
xnor U5108 (N_5108,N_4382,N_4121);
and U5109 (N_5109,N_4061,N_4189);
or U5110 (N_5110,N_4748,N_4195);
or U5111 (N_5111,N_4365,N_4208);
nand U5112 (N_5112,N_4405,N_4304);
xor U5113 (N_5113,N_4578,N_4273);
nand U5114 (N_5114,N_4084,N_4633);
nand U5115 (N_5115,N_4029,N_4353);
and U5116 (N_5116,N_4354,N_4200);
nand U5117 (N_5117,N_4129,N_4622);
xnor U5118 (N_5118,N_4478,N_4684);
and U5119 (N_5119,N_4058,N_4606);
and U5120 (N_5120,N_4771,N_4065);
nand U5121 (N_5121,N_4016,N_4164);
or U5122 (N_5122,N_4035,N_4424);
nor U5123 (N_5123,N_4018,N_4001);
or U5124 (N_5124,N_4796,N_4416);
and U5125 (N_5125,N_4387,N_4337);
nand U5126 (N_5126,N_4283,N_4377);
nand U5127 (N_5127,N_4202,N_4726);
nand U5128 (N_5128,N_4499,N_4588);
nor U5129 (N_5129,N_4538,N_4116);
xor U5130 (N_5130,N_4715,N_4242);
nor U5131 (N_5131,N_4645,N_4070);
nor U5132 (N_5132,N_4607,N_4553);
xnor U5133 (N_5133,N_4101,N_4563);
nand U5134 (N_5134,N_4401,N_4493);
nand U5135 (N_5135,N_4507,N_4527);
and U5136 (N_5136,N_4229,N_4757);
or U5137 (N_5137,N_4642,N_4220);
xor U5138 (N_5138,N_4721,N_4551);
xor U5139 (N_5139,N_4778,N_4528);
xor U5140 (N_5140,N_4346,N_4331);
or U5141 (N_5141,N_4107,N_4572);
nor U5142 (N_5142,N_4420,N_4761);
nor U5143 (N_5143,N_4235,N_4727);
nor U5144 (N_5144,N_4490,N_4290);
xor U5145 (N_5145,N_4217,N_4253);
or U5146 (N_5146,N_4788,N_4299);
and U5147 (N_5147,N_4453,N_4339);
xnor U5148 (N_5148,N_4732,N_4509);
or U5149 (N_5149,N_4131,N_4610);
xor U5150 (N_5150,N_4228,N_4184);
and U5151 (N_5151,N_4449,N_4301);
xnor U5152 (N_5152,N_4564,N_4094);
nor U5153 (N_5153,N_4744,N_4392);
xnor U5154 (N_5154,N_4244,N_4450);
or U5155 (N_5155,N_4167,N_4479);
and U5156 (N_5156,N_4534,N_4705);
and U5157 (N_5157,N_4798,N_4679);
nor U5158 (N_5158,N_4628,N_4048);
nand U5159 (N_5159,N_4041,N_4364);
xnor U5160 (N_5160,N_4742,N_4179);
and U5161 (N_5161,N_4187,N_4442);
nand U5162 (N_5162,N_4441,N_4618);
xor U5163 (N_5163,N_4031,N_4555);
xor U5164 (N_5164,N_4388,N_4106);
nor U5165 (N_5165,N_4305,N_4137);
nor U5166 (N_5166,N_4529,N_4207);
or U5167 (N_5167,N_4359,N_4199);
and U5168 (N_5168,N_4250,N_4249);
or U5169 (N_5169,N_4646,N_4605);
nor U5170 (N_5170,N_4141,N_4797);
and U5171 (N_5171,N_4599,N_4430);
or U5172 (N_5172,N_4067,N_4120);
xnor U5173 (N_5173,N_4506,N_4155);
or U5174 (N_5174,N_4526,N_4443);
and U5175 (N_5175,N_4546,N_4702);
or U5176 (N_5176,N_4589,N_4468);
or U5177 (N_5177,N_4768,N_4298);
nor U5178 (N_5178,N_4536,N_4738);
xnor U5179 (N_5179,N_4523,N_4657);
nor U5180 (N_5180,N_4530,N_4333);
xor U5181 (N_5181,N_4488,N_4160);
nor U5182 (N_5182,N_4056,N_4585);
nor U5183 (N_5183,N_4171,N_4315);
and U5184 (N_5184,N_4034,N_4445);
nand U5185 (N_5185,N_4085,N_4542);
nor U5186 (N_5186,N_4327,N_4156);
nor U5187 (N_5187,N_4225,N_4310);
nand U5188 (N_5188,N_4210,N_4740);
or U5189 (N_5189,N_4115,N_4444);
or U5190 (N_5190,N_4302,N_4292);
and U5191 (N_5191,N_4051,N_4233);
nand U5192 (N_5192,N_4593,N_4076);
xor U5193 (N_5193,N_4729,N_4185);
xnor U5194 (N_5194,N_4719,N_4693);
nor U5195 (N_5195,N_4146,N_4252);
xor U5196 (N_5196,N_4545,N_4734);
or U5197 (N_5197,N_4565,N_4531);
nand U5198 (N_5198,N_4330,N_4519);
or U5199 (N_5199,N_4324,N_4552);
or U5200 (N_5200,N_4254,N_4749);
nand U5201 (N_5201,N_4538,N_4381);
or U5202 (N_5202,N_4702,N_4107);
xnor U5203 (N_5203,N_4733,N_4167);
xnor U5204 (N_5204,N_4520,N_4417);
and U5205 (N_5205,N_4539,N_4072);
nor U5206 (N_5206,N_4426,N_4670);
nand U5207 (N_5207,N_4642,N_4177);
nor U5208 (N_5208,N_4205,N_4438);
and U5209 (N_5209,N_4412,N_4300);
and U5210 (N_5210,N_4331,N_4047);
nor U5211 (N_5211,N_4104,N_4339);
nor U5212 (N_5212,N_4755,N_4568);
xnor U5213 (N_5213,N_4438,N_4023);
xnor U5214 (N_5214,N_4141,N_4530);
and U5215 (N_5215,N_4128,N_4086);
nor U5216 (N_5216,N_4330,N_4462);
or U5217 (N_5217,N_4124,N_4127);
nor U5218 (N_5218,N_4152,N_4131);
xor U5219 (N_5219,N_4375,N_4536);
xnor U5220 (N_5220,N_4065,N_4433);
xnor U5221 (N_5221,N_4504,N_4285);
nand U5222 (N_5222,N_4288,N_4529);
and U5223 (N_5223,N_4740,N_4797);
nand U5224 (N_5224,N_4221,N_4618);
and U5225 (N_5225,N_4645,N_4482);
nor U5226 (N_5226,N_4304,N_4390);
and U5227 (N_5227,N_4568,N_4549);
or U5228 (N_5228,N_4512,N_4505);
and U5229 (N_5229,N_4060,N_4461);
nand U5230 (N_5230,N_4416,N_4434);
and U5231 (N_5231,N_4274,N_4128);
nand U5232 (N_5232,N_4339,N_4645);
xnor U5233 (N_5233,N_4526,N_4730);
and U5234 (N_5234,N_4196,N_4607);
or U5235 (N_5235,N_4369,N_4631);
nand U5236 (N_5236,N_4518,N_4333);
or U5237 (N_5237,N_4315,N_4532);
nor U5238 (N_5238,N_4447,N_4164);
or U5239 (N_5239,N_4313,N_4367);
nand U5240 (N_5240,N_4555,N_4079);
or U5241 (N_5241,N_4366,N_4023);
xor U5242 (N_5242,N_4349,N_4201);
nand U5243 (N_5243,N_4001,N_4656);
nor U5244 (N_5244,N_4168,N_4537);
xnor U5245 (N_5245,N_4579,N_4046);
or U5246 (N_5246,N_4435,N_4662);
xor U5247 (N_5247,N_4497,N_4640);
and U5248 (N_5248,N_4232,N_4130);
xor U5249 (N_5249,N_4324,N_4123);
xor U5250 (N_5250,N_4219,N_4393);
nor U5251 (N_5251,N_4011,N_4177);
and U5252 (N_5252,N_4433,N_4194);
nor U5253 (N_5253,N_4549,N_4212);
nor U5254 (N_5254,N_4082,N_4733);
nand U5255 (N_5255,N_4390,N_4502);
and U5256 (N_5256,N_4343,N_4024);
and U5257 (N_5257,N_4721,N_4688);
or U5258 (N_5258,N_4705,N_4181);
nand U5259 (N_5259,N_4447,N_4491);
nor U5260 (N_5260,N_4327,N_4666);
nor U5261 (N_5261,N_4600,N_4298);
xor U5262 (N_5262,N_4219,N_4751);
nor U5263 (N_5263,N_4593,N_4214);
nand U5264 (N_5264,N_4122,N_4652);
xnor U5265 (N_5265,N_4643,N_4026);
nor U5266 (N_5266,N_4559,N_4469);
nand U5267 (N_5267,N_4081,N_4560);
nor U5268 (N_5268,N_4761,N_4597);
nand U5269 (N_5269,N_4749,N_4673);
or U5270 (N_5270,N_4064,N_4307);
nor U5271 (N_5271,N_4499,N_4740);
xnor U5272 (N_5272,N_4305,N_4240);
nor U5273 (N_5273,N_4713,N_4425);
xor U5274 (N_5274,N_4709,N_4188);
or U5275 (N_5275,N_4006,N_4038);
xor U5276 (N_5276,N_4374,N_4495);
nor U5277 (N_5277,N_4026,N_4342);
xor U5278 (N_5278,N_4054,N_4024);
nor U5279 (N_5279,N_4166,N_4054);
xor U5280 (N_5280,N_4034,N_4104);
nor U5281 (N_5281,N_4040,N_4191);
nand U5282 (N_5282,N_4434,N_4322);
nand U5283 (N_5283,N_4278,N_4269);
or U5284 (N_5284,N_4394,N_4352);
nand U5285 (N_5285,N_4499,N_4450);
and U5286 (N_5286,N_4586,N_4026);
and U5287 (N_5287,N_4567,N_4597);
xnor U5288 (N_5288,N_4039,N_4428);
nand U5289 (N_5289,N_4232,N_4133);
nor U5290 (N_5290,N_4646,N_4490);
or U5291 (N_5291,N_4449,N_4540);
or U5292 (N_5292,N_4436,N_4536);
nand U5293 (N_5293,N_4302,N_4187);
or U5294 (N_5294,N_4153,N_4618);
or U5295 (N_5295,N_4788,N_4392);
xor U5296 (N_5296,N_4460,N_4020);
nand U5297 (N_5297,N_4744,N_4270);
and U5298 (N_5298,N_4393,N_4144);
or U5299 (N_5299,N_4672,N_4503);
nand U5300 (N_5300,N_4646,N_4219);
nand U5301 (N_5301,N_4650,N_4150);
and U5302 (N_5302,N_4590,N_4172);
xor U5303 (N_5303,N_4469,N_4252);
xor U5304 (N_5304,N_4209,N_4199);
or U5305 (N_5305,N_4487,N_4563);
nor U5306 (N_5306,N_4405,N_4061);
nand U5307 (N_5307,N_4407,N_4422);
or U5308 (N_5308,N_4133,N_4499);
and U5309 (N_5309,N_4702,N_4453);
and U5310 (N_5310,N_4567,N_4434);
nand U5311 (N_5311,N_4698,N_4649);
and U5312 (N_5312,N_4321,N_4384);
and U5313 (N_5313,N_4008,N_4124);
nand U5314 (N_5314,N_4351,N_4510);
nor U5315 (N_5315,N_4151,N_4111);
nand U5316 (N_5316,N_4140,N_4321);
and U5317 (N_5317,N_4399,N_4790);
nor U5318 (N_5318,N_4745,N_4009);
xnor U5319 (N_5319,N_4334,N_4534);
and U5320 (N_5320,N_4281,N_4096);
nand U5321 (N_5321,N_4241,N_4115);
nor U5322 (N_5322,N_4472,N_4621);
and U5323 (N_5323,N_4259,N_4516);
or U5324 (N_5324,N_4101,N_4278);
nor U5325 (N_5325,N_4646,N_4489);
and U5326 (N_5326,N_4516,N_4646);
and U5327 (N_5327,N_4504,N_4468);
nor U5328 (N_5328,N_4321,N_4357);
xor U5329 (N_5329,N_4699,N_4439);
xor U5330 (N_5330,N_4166,N_4118);
or U5331 (N_5331,N_4032,N_4202);
and U5332 (N_5332,N_4204,N_4337);
nor U5333 (N_5333,N_4195,N_4580);
xor U5334 (N_5334,N_4764,N_4795);
xor U5335 (N_5335,N_4785,N_4573);
or U5336 (N_5336,N_4576,N_4572);
and U5337 (N_5337,N_4699,N_4259);
nor U5338 (N_5338,N_4369,N_4466);
nand U5339 (N_5339,N_4487,N_4723);
nor U5340 (N_5340,N_4049,N_4706);
or U5341 (N_5341,N_4540,N_4287);
xor U5342 (N_5342,N_4386,N_4396);
xnor U5343 (N_5343,N_4050,N_4099);
nand U5344 (N_5344,N_4436,N_4690);
or U5345 (N_5345,N_4647,N_4069);
nand U5346 (N_5346,N_4141,N_4659);
nor U5347 (N_5347,N_4344,N_4161);
xnor U5348 (N_5348,N_4413,N_4650);
or U5349 (N_5349,N_4081,N_4619);
and U5350 (N_5350,N_4132,N_4232);
nand U5351 (N_5351,N_4735,N_4042);
xnor U5352 (N_5352,N_4477,N_4751);
nor U5353 (N_5353,N_4542,N_4450);
nand U5354 (N_5354,N_4378,N_4561);
nor U5355 (N_5355,N_4443,N_4281);
nand U5356 (N_5356,N_4177,N_4348);
xor U5357 (N_5357,N_4639,N_4041);
nand U5358 (N_5358,N_4018,N_4656);
nor U5359 (N_5359,N_4593,N_4476);
or U5360 (N_5360,N_4263,N_4149);
and U5361 (N_5361,N_4716,N_4244);
nor U5362 (N_5362,N_4095,N_4323);
nor U5363 (N_5363,N_4353,N_4552);
or U5364 (N_5364,N_4387,N_4716);
nor U5365 (N_5365,N_4694,N_4381);
nor U5366 (N_5366,N_4653,N_4258);
or U5367 (N_5367,N_4779,N_4092);
or U5368 (N_5368,N_4300,N_4438);
or U5369 (N_5369,N_4157,N_4693);
and U5370 (N_5370,N_4360,N_4658);
and U5371 (N_5371,N_4614,N_4517);
nor U5372 (N_5372,N_4551,N_4378);
and U5373 (N_5373,N_4201,N_4543);
or U5374 (N_5374,N_4317,N_4316);
xnor U5375 (N_5375,N_4456,N_4751);
or U5376 (N_5376,N_4038,N_4518);
nor U5377 (N_5377,N_4660,N_4306);
xor U5378 (N_5378,N_4553,N_4670);
xnor U5379 (N_5379,N_4020,N_4455);
and U5380 (N_5380,N_4782,N_4157);
xnor U5381 (N_5381,N_4439,N_4137);
nand U5382 (N_5382,N_4382,N_4246);
xor U5383 (N_5383,N_4297,N_4088);
nand U5384 (N_5384,N_4083,N_4685);
or U5385 (N_5385,N_4002,N_4005);
xor U5386 (N_5386,N_4677,N_4063);
xor U5387 (N_5387,N_4544,N_4124);
nor U5388 (N_5388,N_4107,N_4073);
and U5389 (N_5389,N_4392,N_4172);
or U5390 (N_5390,N_4603,N_4085);
nor U5391 (N_5391,N_4262,N_4789);
or U5392 (N_5392,N_4199,N_4250);
xnor U5393 (N_5393,N_4443,N_4114);
xnor U5394 (N_5394,N_4148,N_4262);
or U5395 (N_5395,N_4619,N_4284);
or U5396 (N_5396,N_4174,N_4513);
xnor U5397 (N_5397,N_4318,N_4590);
nor U5398 (N_5398,N_4712,N_4265);
nand U5399 (N_5399,N_4702,N_4588);
nand U5400 (N_5400,N_4224,N_4220);
nor U5401 (N_5401,N_4104,N_4750);
and U5402 (N_5402,N_4018,N_4556);
xnor U5403 (N_5403,N_4463,N_4539);
or U5404 (N_5404,N_4497,N_4744);
or U5405 (N_5405,N_4796,N_4210);
nor U5406 (N_5406,N_4765,N_4361);
nor U5407 (N_5407,N_4460,N_4331);
nand U5408 (N_5408,N_4769,N_4427);
or U5409 (N_5409,N_4707,N_4747);
nor U5410 (N_5410,N_4218,N_4242);
nor U5411 (N_5411,N_4641,N_4310);
xnor U5412 (N_5412,N_4275,N_4541);
or U5413 (N_5413,N_4472,N_4612);
xnor U5414 (N_5414,N_4774,N_4435);
xor U5415 (N_5415,N_4610,N_4178);
and U5416 (N_5416,N_4665,N_4271);
nand U5417 (N_5417,N_4176,N_4559);
or U5418 (N_5418,N_4292,N_4225);
nor U5419 (N_5419,N_4439,N_4523);
nand U5420 (N_5420,N_4271,N_4794);
nor U5421 (N_5421,N_4590,N_4092);
nand U5422 (N_5422,N_4597,N_4346);
nand U5423 (N_5423,N_4122,N_4048);
or U5424 (N_5424,N_4204,N_4296);
and U5425 (N_5425,N_4495,N_4041);
xnor U5426 (N_5426,N_4612,N_4148);
and U5427 (N_5427,N_4345,N_4675);
and U5428 (N_5428,N_4173,N_4286);
nand U5429 (N_5429,N_4716,N_4145);
and U5430 (N_5430,N_4652,N_4708);
or U5431 (N_5431,N_4767,N_4310);
nor U5432 (N_5432,N_4647,N_4314);
or U5433 (N_5433,N_4069,N_4369);
nand U5434 (N_5434,N_4188,N_4659);
and U5435 (N_5435,N_4170,N_4136);
and U5436 (N_5436,N_4696,N_4243);
xnor U5437 (N_5437,N_4360,N_4491);
or U5438 (N_5438,N_4389,N_4751);
nor U5439 (N_5439,N_4017,N_4257);
and U5440 (N_5440,N_4274,N_4777);
xnor U5441 (N_5441,N_4178,N_4448);
nand U5442 (N_5442,N_4762,N_4406);
or U5443 (N_5443,N_4462,N_4786);
and U5444 (N_5444,N_4378,N_4328);
or U5445 (N_5445,N_4043,N_4473);
nand U5446 (N_5446,N_4511,N_4179);
and U5447 (N_5447,N_4271,N_4383);
and U5448 (N_5448,N_4645,N_4086);
nor U5449 (N_5449,N_4358,N_4033);
or U5450 (N_5450,N_4624,N_4765);
or U5451 (N_5451,N_4651,N_4242);
nor U5452 (N_5452,N_4530,N_4059);
and U5453 (N_5453,N_4465,N_4785);
or U5454 (N_5454,N_4684,N_4456);
nor U5455 (N_5455,N_4012,N_4755);
nand U5456 (N_5456,N_4471,N_4319);
and U5457 (N_5457,N_4297,N_4254);
or U5458 (N_5458,N_4234,N_4587);
nand U5459 (N_5459,N_4427,N_4595);
or U5460 (N_5460,N_4475,N_4747);
nand U5461 (N_5461,N_4394,N_4341);
or U5462 (N_5462,N_4634,N_4077);
xor U5463 (N_5463,N_4395,N_4393);
nor U5464 (N_5464,N_4557,N_4421);
or U5465 (N_5465,N_4475,N_4294);
nor U5466 (N_5466,N_4439,N_4729);
xor U5467 (N_5467,N_4421,N_4685);
xor U5468 (N_5468,N_4746,N_4125);
or U5469 (N_5469,N_4014,N_4517);
xnor U5470 (N_5470,N_4561,N_4787);
xnor U5471 (N_5471,N_4380,N_4009);
or U5472 (N_5472,N_4610,N_4005);
xor U5473 (N_5473,N_4132,N_4423);
and U5474 (N_5474,N_4345,N_4595);
and U5475 (N_5475,N_4044,N_4492);
nand U5476 (N_5476,N_4375,N_4234);
or U5477 (N_5477,N_4242,N_4356);
xnor U5478 (N_5478,N_4416,N_4283);
nand U5479 (N_5479,N_4121,N_4477);
and U5480 (N_5480,N_4638,N_4305);
xnor U5481 (N_5481,N_4427,N_4460);
or U5482 (N_5482,N_4324,N_4611);
nor U5483 (N_5483,N_4664,N_4743);
xor U5484 (N_5484,N_4269,N_4218);
and U5485 (N_5485,N_4701,N_4322);
or U5486 (N_5486,N_4276,N_4636);
or U5487 (N_5487,N_4052,N_4575);
xor U5488 (N_5488,N_4326,N_4433);
and U5489 (N_5489,N_4217,N_4785);
and U5490 (N_5490,N_4487,N_4134);
and U5491 (N_5491,N_4406,N_4516);
xnor U5492 (N_5492,N_4751,N_4005);
and U5493 (N_5493,N_4446,N_4201);
xnor U5494 (N_5494,N_4553,N_4783);
nand U5495 (N_5495,N_4105,N_4172);
or U5496 (N_5496,N_4631,N_4438);
xor U5497 (N_5497,N_4671,N_4061);
nand U5498 (N_5498,N_4434,N_4667);
and U5499 (N_5499,N_4136,N_4620);
nor U5500 (N_5500,N_4052,N_4296);
and U5501 (N_5501,N_4593,N_4655);
xor U5502 (N_5502,N_4321,N_4666);
and U5503 (N_5503,N_4297,N_4134);
xor U5504 (N_5504,N_4433,N_4346);
nor U5505 (N_5505,N_4227,N_4569);
nor U5506 (N_5506,N_4385,N_4176);
or U5507 (N_5507,N_4640,N_4729);
nand U5508 (N_5508,N_4487,N_4229);
nand U5509 (N_5509,N_4586,N_4078);
or U5510 (N_5510,N_4034,N_4142);
xnor U5511 (N_5511,N_4394,N_4303);
and U5512 (N_5512,N_4641,N_4138);
and U5513 (N_5513,N_4416,N_4066);
nand U5514 (N_5514,N_4721,N_4144);
or U5515 (N_5515,N_4261,N_4319);
nand U5516 (N_5516,N_4723,N_4474);
nor U5517 (N_5517,N_4686,N_4032);
and U5518 (N_5518,N_4460,N_4772);
or U5519 (N_5519,N_4183,N_4108);
xor U5520 (N_5520,N_4602,N_4508);
and U5521 (N_5521,N_4469,N_4090);
xor U5522 (N_5522,N_4741,N_4642);
or U5523 (N_5523,N_4632,N_4191);
and U5524 (N_5524,N_4243,N_4380);
nor U5525 (N_5525,N_4590,N_4040);
nand U5526 (N_5526,N_4184,N_4689);
xnor U5527 (N_5527,N_4171,N_4466);
nand U5528 (N_5528,N_4015,N_4659);
and U5529 (N_5529,N_4655,N_4332);
or U5530 (N_5530,N_4645,N_4123);
nor U5531 (N_5531,N_4112,N_4698);
xnor U5532 (N_5532,N_4469,N_4538);
and U5533 (N_5533,N_4516,N_4493);
and U5534 (N_5534,N_4577,N_4527);
and U5535 (N_5535,N_4047,N_4281);
xor U5536 (N_5536,N_4760,N_4566);
or U5537 (N_5537,N_4034,N_4045);
xnor U5538 (N_5538,N_4278,N_4774);
nand U5539 (N_5539,N_4353,N_4491);
xor U5540 (N_5540,N_4394,N_4099);
or U5541 (N_5541,N_4071,N_4536);
nor U5542 (N_5542,N_4302,N_4681);
nor U5543 (N_5543,N_4085,N_4166);
xor U5544 (N_5544,N_4552,N_4611);
nand U5545 (N_5545,N_4665,N_4364);
and U5546 (N_5546,N_4708,N_4254);
or U5547 (N_5547,N_4495,N_4665);
nand U5548 (N_5548,N_4036,N_4407);
nand U5549 (N_5549,N_4410,N_4273);
xnor U5550 (N_5550,N_4324,N_4554);
nor U5551 (N_5551,N_4288,N_4272);
and U5552 (N_5552,N_4190,N_4511);
or U5553 (N_5553,N_4283,N_4400);
nor U5554 (N_5554,N_4635,N_4494);
or U5555 (N_5555,N_4238,N_4515);
and U5556 (N_5556,N_4245,N_4581);
or U5557 (N_5557,N_4082,N_4623);
xor U5558 (N_5558,N_4107,N_4408);
or U5559 (N_5559,N_4248,N_4769);
or U5560 (N_5560,N_4590,N_4055);
and U5561 (N_5561,N_4539,N_4471);
xor U5562 (N_5562,N_4032,N_4301);
xnor U5563 (N_5563,N_4220,N_4451);
nor U5564 (N_5564,N_4559,N_4242);
nand U5565 (N_5565,N_4114,N_4310);
xnor U5566 (N_5566,N_4746,N_4061);
and U5567 (N_5567,N_4105,N_4672);
nand U5568 (N_5568,N_4229,N_4614);
or U5569 (N_5569,N_4074,N_4135);
or U5570 (N_5570,N_4039,N_4479);
or U5571 (N_5571,N_4033,N_4734);
or U5572 (N_5572,N_4455,N_4516);
or U5573 (N_5573,N_4065,N_4768);
nor U5574 (N_5574,N_4265,N_4238);
nor U5575 (N_5575,N_4709,N_4730);
or U5576 (N_5576,N_4247,N_4144);
nor U5577 (N_5577,N_4391,N_4484);
or U5578 (N_5578,N_4601,N_4283);
nand U5579 (N_5579,N_4756,N_4471);
xnor U5580 (N_5580,N_4645,N_4489);
xor U5581 (N_5581,N_4453,N_4154);
and U5582 (N_5582,N_4313,N_4777);
nor U5583 (N_5583,N_4427,N_4333);
xor U5584 (N_5584,N_4656,N_4208);
nor U5585 (N_5585,N_4099,N_4304);
and U5586 (N_5586,N_4653,N_4200);
nand U5587 (N_5587,N_4760,N_4274);
and U5588 (N_5588,N_4560,N_4105);
nor U5589 (N_5589,N_4529,N_4186);
xor U5590 (N_5590,N_4645,N_4792);
xor U5591 (N_5591,N_4643,N_4144);
and U5592 (N_5592,N_4298,N_4589);
and U5593 (N_5593,N_4525,N_4423);
or U5594 (N_5594,N_4316,N_4367);
nor U5595 (N_5595,N_4414,N_4594);
nand U5596 (N_5596,N_4016,N_4369);
nor U5597 (N_5597,N_4298,N_4280);
xor U5598 (N_5598,N_4143,N_4331);
or U5599 (N_5599,N_4080,N_4594);
or U5600 (N_5600,N_5079,N_5581);
xnor U5601 (N_5601,N_5372,N_5162);
and U5602 (N_5602,N_5554,N_5595);
nor U5603 (N_5603,N_5267,N_5117);
and U5604 (N_5604,N_5473,N_5413);
nand U5605 (N_5605,N_5199,N_5388);
or U5606 (N_5606,N_4826,N_5052);
xor U5607 (N_5607,N_5095,N_4984);
or U5608 (N_5608,N_5013,N_5328);
nand U5609 (N_5609,N_4943,N_5431);
or U5610 (N_5610,N_4901,N_5030);
and U5611 (N_5611,N_4992,N_5424);
or U5612 (N_5612,N_5190,N_4962);
xor U5613 (N_5613,N_5081,N_5035);
and U5614 (N_5614,N_5029,N_5256);
xor U5615 (N_5615,N_4838,N_5153);
and U5616 (N_5616,N_5545,N_5332);
nor U5617 (N_5617,N_5341,N_4823);
xnor U5618 (N_5618,N_5155,N_5154);
nor U5619 (N_5619,N_5495,N_5563);
or U5620 (N_5620,N_4946,N_5214);
and U5621 (N_5621,N_4923,N_5592);
nand U5622 (N_5622,N_4812,N_5116);
or U5623 (N_5623,N_5259,N_5324);
xnor U5624 (N_5624,N_5167,N_5419);
nand U5625 (N_5625,N_5379,N_5232);
xnor U5626 (N_5626,N_5446,N_5350);
and U5627 (N_5627,N_5498,N_5156);
xnor U5628 (N_5628,N_5230,N_5089);
or U5629 (N_5629,N_4819,N_4836);
nand U5630 (N_5630,N_5058,N_5489);
and U5631 (N_5631,N_5285,N_5150);
xnor U5632 (N_5632,N_5304,N_4816);
xor U5633 (N_5633,N_5134,N_5497);
nor U5634 (N_5634,N_5564,N_5309);
nand U5635 (N_5635,N_4869,N_5492);
and U5636 (N_5636,N_5011,N_5096);
or U5637 (N_5637,N_5201,N_5051);
nand U5638 (N_5638,N_5480,N_5010);
nor U5639 (N_5639,N_5394,N_5503);
xnor U5640 (N_5640,N_5561,N_5351);
and U5641 (N_5641,N_4807,N_4861);
nor U5642 (N_5642,N_4999,N_5093);
nand U5643 (N_5643,N_4871,N_5042);
and U5644 (N_5644,N_5044,N_5175);
xor U5645 (N_5645,N_5061,N_5034);
nor U5646 (N_5646,N_5063,N_5123);
or U5647 (N_5647,N_5120,N_4817);
nor U5648 (N_5648,N_5420,N_5477);
or U5649 (N_5649,N_4844,N_5091);
or U5650 (N_5650,N_5435,N_5414);
or U5651 (N_5651,N_5223,N_5550);
xor U5652 (N_5652,N_4841,N_4857);
xnor U5653 (N_5653,N_4976,N_5344);
xor U5654 (N_5654,N_5457,N_5205);
and U5655 (N_5655,N_5004,N_5121);
nor U5656 (N_5656,N_4971,N_5142);
or U5657 (N_5657,N_5478,N_5407);
and U5658 (N_5658,N_4828,N_5272);
and U5659 (N_5659,N_5448,N_5415);
nand U5660 (N_5660,N_5118,N_4883);
and U5661 (N_5661,N_5085,N_5196);
xnor U5662 (N_5662,N_5166,N_5247);
nor U5663 (N_5663,N_4804,N_5390);
nand U5664 (N_5664,N_5026,N_5322);
and U5665 (N_5665,N_4960,N_4919);
and U5666 (N_5666,N_5455,N_5306);
nor U5667 (N_5667,N_5077,N_4998);
and U5668 (N_5668,N_5228,N_5231);
nand U5669 (N_5669,N_4986,N_4996);
xnor U5670 (N_5670,N_5193,N_5406);
and U5671 (N_5671,N_5486,N_5296);
or U5672 (N_5672,N_5366,N_5585);
and U5673 (N_5673,N_5298,N_5182);
and U5674 (N_5674,N_5207,N_5050);
nor U5675 (N_5675,N_4865,N_5377);
xor U5676 (N_5676,N_5084,N_5482);
nand U5677 (N_5677,N_5066,N_4941);
xnor U5678 (N_5678,N_5152,N_5009);
nor U5679 (N_5679,N_4965,N_5151);
xnor U5680 (N_5680,N_5251,N_5395);
and U5681 (N_5681,N_4940,N_4934);
or U5682 (N_5682,N_5040,N_5500);
and U5683 (N_5683,N_5534,N_5293);
or U5684 (N_5684,N_4955,N_5580);
nand U5685 (N_5685,N_4933,N_5147);
nor U5686 (N_5686,N_5039,N_5253);
nand U5687 (N_5687,N_5336,N_4967);
nand U5688 (N_5688,N_5551,N_4852);
or U5689 (N_5689,N_5496,N_5168);
nor U5690 (N_5690,N_5276,N_5481);
nand U5691 (N_5691,N_5467,N_4886);
nand U5692 (N_5692,N_5518,N_5082);
xor U5693 (N_5693,N_5227,N_5140);
nor U5694 (N_5694,N_5280,N_5187);
xor U5695 (N_5695,N_4927,N_5454);
xor U5696 (N_5696,N_5593,N_5434);
xor U5697 (N_5697,N_4859,N_4954);
nand U5698 (N_5698,N_5249,N_5098);
xnor U5699 (N_5699,N_5074,N_5261);
and U5700 (N_5700,N_4888,N_5427);
xor U5701 (N_5701,N_5437,N_4881);
xnor U5702 (N_5702,N_5114,N_4851);
nor U5703 (N_5703,N_5240,N_5024);
or U5704 (N_5704,N_5472,N_5343);
nor U5705 (N_5705,N_5352,N_5381);
xnor U5706 (N_5706,N_4931,N_5226);
xnor U5707 (N_5707,N_4825,N_5036);
or U5708 (N_5708,N_5290,N_4890);
nand U5709 (N_5709,N_5549,N_5405);
and U5710 (N_5710,N_5105,N_5456);
or U5711 (N_5711,N_4832,N_5255);
nor U5712 (N_5712,N_5522,N_5520);
nor U5713 (N_5713,N_5109,N_5436);
nand U5714 (N_5714,N_5005,N_4977);
nand U5715 (N_5715,N_4800,N_5502);
xor U5716 (N_5716,N_5494,N_5062);
nand U5717 (N_5717,N_4952,N_4806);
xnor U5718 (N_5718,N_5440,N_5542);
and U5719 (N_5719,N_5501,N_5311);
xnor U5720 (N_5720,N_5566,N_5138);
xnor U5721 (N_5721,N_4975,N_5452);
nor U5722 (N_5722,N_4875,N_5568);
or U5723 (N_5723,N_4930,N_5465);
or U5724 (N_5724,N_5099,N_5334);
and U5725 (N_5725,N_5001,N_5519);
xor U5726 (N_5726,N_5560,N_5169);
nand U5727 (N_5727,N_5521,N_5313);
nand U5728 (N_5728,N_4897,N_5006);
nor U5729 (N_5729,N_5347,N_5179);
xnor U5730 (N_5730,N_5181,N_5003);
nand U5731 (N_5731,N_4981,N_5428);
nor U5732 (N_5732,N_5357,N_4829);
nor U5733 (N_5733,N_5335,N_4892);
xnor U5734 (N_5734,N_5246,N_5163);
xnor U5735 (N_5735,N_4922,N_4866);
xor U5736 (N_5736,N_5224,N_4863);
and U5737 (N_5737,N_5137,N_5198);
xnor U5738 (N_5738,N_4903,N_5443);
nand U5739 (N_5739,N_4902,N_5479);
nor U5740 (N_5740,N_4877,N_4963);
and U5741 (N_5741,N_5469,N_5191);
or U5742 (N_5742,N_4970,N_4924);
nor U5743 (N_5743,N_5080,N_5587);
and U5744 (N_5744,N_4891,N_5028);
nand U5745 (N_5745,N_5361,N_5514);
nand U5746 (N_5746,N_5476,N_5386);
and U5747 (N_5747,N_5189,N_5139);
or U5748 (N_5748,N_5057,N_5043);
and U5749 (N_5749,N_5283,N_5583);
nor U5750 (N_5750,N_5556,N_5576);
xor U5751 (N_5751,N_5316,N_5348);
xor U5752 (N_5752,N_5515,N_5056);
or U5753 (N_5753,N_5369,N_5220);
and U5754 (N_5754,N_5252,N_5289);
nor U5755 (N_5755,N_5119,N_5070);
nand U5756 (N_5756,N_5216,N_5046);
nor U5757 (N_5757,N_5064,N_5398);
nor U5758 (N_5758,N_5229,N_5543);
nor U5759 (N_5759,N_5364,N_5371);
nand U5760 (N_5760,N_5149,N_4935);
or U5761 (N_5761,N_5233,N_4928);
nor U5762 (N_5762,N_5319,N_5483);
nand U5763 (N_5763,N_5559,N_5279);
or U5764 (N_5764,N_5132,N_5432);
nor U5765 (N_5765,N_4853,N_4840);
and U5766 (N_5766,N_5106,N_4951);
nor U5767 (N_5767,N_4969,N_5088);
xor U5768 (N_5768,N_5254,N_5411);
and U5769 (N_5769,N_5594,N_4990);
nand U5770 (N_5770,N_5392,N_5072);
or U5771 (N_5771,N_5192,N_5530);
nand U5772 (N_5772,N_4856,N_5499);
xnor U5773 (N_5773,N_5389,N_5177);
or U5774 (N_5774,N_5451,N_5111);
nor U5775 (N_5775,N_4839,N_5470);
nand U5776 (N_5776,N_4989,N_5474);
and U5777 (N_5777,N_5374,N_5108);
nand U5778 (N_5778,N_5023,N_5217);
or U5779 (N_5779,N_5490,N_5596);
or U5780 (N_5780,N_4994,N_5513);
nor U5781 (N_5781,N_5429,N_5218);
nor U5782 (N_5782,N_5421,N_4810);
or U5783 (N_5783,N_5048,N_4909);
or U5784 (N_5784,N_5222,N_4818);
xnor U5785 (N_5785,N_4862,N_5213);
nor U5786 (N_5786,N_5022,N_5508);
or U5787 (N_5787,N_4926,N_4929);
nand U5788 (N_5788,N_4980,N_5572);
or U5789 (N_5789,N_5487,N_5025);
xor U5790 (N_5790,N_5209,N_5412);
nand U5791 (N_5791,N_4815,N_5104);
xnor U5792 (N_5792,N_5321,N_5200);
nor U5793 (N_5793,N_5598,N_5271);
nor U5794 (N_5794,N_5297,N_5397);
nand U5795 (N_5795,N_5387,N_5577);
nor U5796 (N_5796,N_4887,N_5422);
or U5797 (N_5797,N_5288,N_5242);
and U5798 (N_5798,N_5076,N_5349);
nand U5799 (N_5799,N_4958,N_5273);
nor U5800 (N_5800,N_5017,N_5423);
and U5801 (N_5801,N_5346,N_5071);
nand U5802 (N_5802,N_5176,N_5538);
nand U5803 (N_5803,N_5541,N_5342);
nand U5804 (N_5804,N_4956,N_5575);
xnor U5805 (N_5805,N_5203,N_4824);
and U5806 (N_5806,N_5110,N_5202);
nor U5807 (N_5807,N_4864,N_4830);
xnor U5808 (N_5808,N_5212,N_4837);
and U5809 (N_5809,N_5065,N_5250);
and U5810 (N_5810,N_4882,N_5416);
xnor U5811 (N_5811,N_5512,N_4845);
and U5812 (N_5812,N_5268,N_4885);
or U5813 (N_5813,N_4936,N_5532);
and U5814 (N_5814,N_4915,N_5488);
nor U5815 (N_5815,N_5525,N_5015);
xor U5816 (N_5816,N_5225,N_5102);
or U5817 (N_5817,N_4910,N_5567);
nand U5818 (N_5818,N_5409,N_5008);
or U5819 (N_5819,N_4985,N_5314);
xor U5820 (N_5820,N_4854,N_4966);
and U5821 (N_5821,N_5449,N_4833);
or U5822 (N_5822,N_5358,N_5399);
xnor U5823 (N_5823,N_5517,N_4821);
nor U5824 (N_5824,N_5305,N_5281);
nand U5825 (N_5825,N_5330,N_5107);
nor U5826 (N_5826,N_5590,N_5439);
nand U5827 (N_5827,N_5403,N_5337);
nand U5828 (N_5828,N_4893,N_5049);
nand U5829 (N_5829,N_5248,N_5383);
xnor U5830 (N_5830,N_5582,N_5258);
or U5831 (N_5831,N_5329,N_5385);
nand U5832 (N_5832,N_4831,N_4917);
and U5833 (N_5833,N_4911,N_5204);
xnor U5834 (N_5834,N_4995,N_5353);
and U5835 (N_5835,N_5012,N_4843);
and U5836 (N_5836,N_5073,N_5000);
or U5837 (N_5837,N_5069,N_5165);
xnor U5838 (N_5838,N_5462,N_5112);
nor U5839 (N_5839,N_5055,N_5245);
or U5840 (N_5840,N_5509,N_5404);
nand U5841 (N_5841,N_4988,N_5131);
or U5842 (N_5842,N_5236,N_5333);
xor U5843 (N_5843,N_5370,N_5453);
and U5844 (N_5844,N_4849,N_4874);
nor U5845 (N_5845,N_4913,N_4900);
or U5846 (N_5846,N_4822,N_5274);
or U5847 (N_5847,N_5378,N_5527);
or U5848 (N_5848,N_5038,N_5505);
and U5849 (N_5849,N_4899,N_5468);
or U5850 (N_5850,N_5363,N_4964);
and U5851 (N_5851,N_5345,N_5243);
nand U5852 (N_5852,N_4942,N_5375);
xor U5853 (N_5853,N_5368,N_5463);
or U5854 (N_5854,N_5135,N_5053);
or U5855 (N_5855,N_5555,N_4925);
and U5856 (N_5856,N_5067,N_5360);
or U5857 (N_5857,N_5277,N_5103);
nor U5858 (N_5858,N_5186,N_5506);
xnor U5859 (N_5859,N_5339,N_5211);
xor U5860 (N_5860,N_5376,N_5571);
nand U5861 (N_5861,N_4809,N_4855);
nor U5862 (N_5862,N_5417,N_5578);
xor U5863 (N_5863,N_5589,N_5031);
nand U5864 (N_5864,N_5591,N_5291);
nand U5865 (N_5865,N_5020,N_5239);
and U5866 (N_5866,N_4820,N_5524);
nand U5867 (N_5867,N_5340,N_5302);
nand U5868 (N_5868,N_4937,N_4914);
or U5869 (N_5869,N_4906,N_5599);
nor U5870 (N_5870,N_5529,N_4932);
or U5871 (N_5871,N_5060,N_5426);
xnor U5872 (N_5872,N_4827,N_5402);
nor U5873 (N_5873,N_5188,N_5059);
xor U5874 (N_5874,N_4896,N_5126);
nand U5875 (N_5875,N_5143,N_5170);
nand U5876 (N_5876,N_5068,N_4895);
nor U5877 (N_5877,N_5160,N_5400);
xor U5878 (N_5878,N_5410,N_4868);
nor U5879 (N_5879,N_4873,N_5552);
and U5880 (N_5880,N_4944,N_4879);
or U5881 (N_5881,N_5194,N_5299);
and U5882 (N_5882,N_5037,N_5215);
xor U5883 (N_5883,N_5384,N_5331);
nor U5884 (N_5884,N_5128,N_5325);
xor U5885 (N_5885,N_5235,N_5546);
nand U5886 (N_5886,N_5544,N_4987);
nand U5887 (N_5887,N_5450,N_4950);
and U5888 (N_5888,N_5558,N_4948);
or U5889 (N_5889,N_5401,N_5338);
and U5890 (N_5890,N_5312,N_5101);
and U5891 (N_5891,N_5493,N_4846);
and U5892 (N_5892,N_5445,N_4921);
nor U5893 (N_5893,N_4894,N_5282);
xnor U5894 (N_5894,N_5159,N_5206);
nor U5895 (N_5895,N_5300,N_5584);
nor U5896 (N_5896,N_5510,N_5172);
and U5897 (N_5897,N_5127,N_4858);
and U5898 (N_5898,N_4912,N_5210);
xnor U5899 (N_5899,N_5540,N_5511);
nor U5900 (N_5900,N_5113,N_4860);
or U5901 (N_5901,N_4939,N_5533);
nand U5902 (N_5902,N_5396,N_5491);
or U5903 (N_5903,N_5174,N_4880);
or U5904 (N_5904,N_5086,N_5234);
nor U5905 (N_5905,N_5588,N_5125);
and U5906 (N_5906,N_5425,N_4938);
nor U5907 (N_5907,N_4918,N_5535);
and U5908 (N_5908,N_5041,N_4907);
nor U5909 (N_5909,N_5260,N_5531);
xnor U5910 (N_5910,N_5016,N_5145);
and U5911 (N_5911,N_5327,N_5092);
xnor U5912 (N_5912,N_5507,N_4993);
xnor U5913 (N_5913,N_5265,N_5365);
nand U5914 (N_5914,N_4808,N_5569);
nor U5915 (N_5915,N_5574,N_5553);
and U5916 (N_5916,N_5317,N_5315);
or U5917 (N_5917,N_5078,N_5565);
xor U5918 (N_5918,N_5045,N_5178);
and U5919 (N_5919,N_5320,N_5144);
and U5920 (N_5920,N_5307,N_5461);
xor U5921 (N_5921,N_5278,N_5504);
or U5922 (N_5922,N_5238,N_5286);
xnor U5923 (N_5923,N_5019,N_5244);
xor U5924 (N_5924,N_5141,N_5146);
xnor U5925 (N_5925,N_5275,N_4889);
xor U5926 (N_5926,N_5097,N_4813);
nor U5927 (N_5927,N_5464,N_5441);
or U5928 (N_5928,N_5184,N_4884);
or U5929 (N_5929,N_4848,N_5014);
or U5930 (N_5930,N_4972,N_5570);
or U5931 (N_5931,N_4876,N_5367);
nand U5932 (N_5932,N_4945,N_5197);
or U5933 (N_5933,N_4878,N_4847);
or U5934 (N_5934,N_4947,N_5292);
xor U5935 (N_5935,N_5266,N_4904);
xor U5936 (N_5936,N_5054,N_5460);
or U5937 (N_5937,N_5354,N_5148);
nor U5938 (N_5938,N_5484,N_5183);
or U5939 (N_5939,N_5310,N_5459);
xnor U5940 (N_5940,N_5438,N_5359);
and U5941 (N_5941,N_5241,N_5161);
xnor U5942 (N_5942,N_5075,N_5393);
nor U5943 (N_5943,N_5308,N_4905);
nor U5944 (N_5944,N_4961,N_5158);
xor U5945 (N_5945,N_5180,N_5548);
or U5946 (N_5946,N_5356,N_5264);
or U5947 (N_5947,N_5408,N_4867);
nand U5948 (N_5948,N_5094,N_5418);
xor U5949 (N_5949,N_5547,N_5130);
xor U5950 (N_5950,N_5516,N_5326);
xnor U5951 (N_5951,N_5129,N_4973);
and U5952 (N_5952,N_5269,N_5018);
nor U5953 (N_5953,N_4842,N_4802);
nor U5954 (N_5954,N_5033,N_5391);
nor U5955 (N_5955,N_4814,N_5318);
and U5956 (N_5956,N_5442,N_5171);
xnor U5957 (N_5957,N_5485,N_5164);
nor U5958 (N_5958,N_5475,N_5573);
nor U5959 (N_5959,N_5083,N_5047);
or U5960 (N_5960,N_4957,N_4997);
xnor U5961 (N_5961,N_5087,N_5557);
or U5962 (N_5962,N_5221,N_4979);
or U5963 (N_5963,N_5007,N_5526);
and U5964 (N_5964,N_4974,N_5597);
and U5965 (N_5965,N_5430,N_4991);
or U5966 (N_5966,N_5157,N_4811);
xor U5967 (N_5967,N_5032,N_5380);
nor U5968 (N_5968,N_5536,N_4949);
nand U5969 (N_5969,N_5301,N_5444);
and U5970 (N_5970,N_4953,N_5284);
nor U5971 (N_5971,N_5124,N_5122);
xor U5972 (N_5972,N_5090,N_4978);
or U5973 (N_5973,N_5185,N_5466);
nor U5974 (N_5974,N_5027,N_4959);
or U5975 (N_5975,N_5382,N_5539);
xor U5976 (N_5976,N_4834,N_5471);
or U5977 (N_5977,N_4803,N_4805);
xor U5978 (N_5978,N_4872,N_5447);
or U5979 (N_5979,N_5100,N_5173);
nor U5980 (N_5980,N_4850,N_5195);
nor U5981 (N_5981,N_5262,N_5362);
or U5982 (N_5982,N_5433,N_5323);
nand U5983 (N_5983,N_5208,N_5586);
xor U5984 (N_5984,N_5237,N_4916);
nand U5985 (N_5985,N_5263,N_5355);
or U5986 (N_5986,N_4835,N_5373);
nand U5987 (N_5987,N_5537,N_5136);
or U5988 (N_5988,N_5270,N_4983);
and U5989 (N_5989,N_4968,N_5295);
nor U5990 (N_5990,N_5523,N_5219);
nand U5991 (N_5991,N_5458,N_5002);
nand U5992 (N_5992,N_5528,N_5294);
nand U5993 (N_5993,N_5133,N_4898);
and U5994 (N_5994,N_5303,N_4908);
nor U5995 (N_5995,N_4801,N_5257);
nor U5996 (N_5996,N_5287,N_5579);
xor U5997 (N_5997,N_4920,N_4982);
nand U5998 (N_5998,N_5562,N_5115);
xor U5999 (N_5999,N_4870,N_5021);
or U6000 (N_6000,N_5285,N_5466);
xnor U6001 (N_6001,N_4836,N_4995);
nor U6002 (N_6002,N_5169,N_4823);
nor U6003 (N_6003,N_5489,N_5297);
nand U6004 (N_6004,N_4807,N_5486);
and U6005 (N_6005,N_4982,N_4980);
nand U6006 (N_6006,N_4981,N_5196);
xor U6007 (N_6007,N_5146,N_5218);
or U6008 (N_6008,N_5327,N_4981);
nor U6009 (N_6009,N_5439,N_5397);
nand U6010 (N_6010,N_5062,N_4872);
or U6011 (N_6011,N_5467,N_5098);
nand U6012 (N_6012,N_5574,N_4868);
nor U6013 (N_6013,N_5546,N_4931);
and U6014 (N_6014,N_5458,N_5084);
xor U6015 (N_6015,N_5464,N_5034);
or U6016 (N_6016,N_5482,N_5279);
or U6017 (N_6017,N_5018,N_5365);
nand U6018 (N_6018,N_5123,N_5599);
or U6019 (N_6019,N_5361,N_5286);
nor U6020 (N_6020,N_4995,N_4984);
nand U6021 (N_6021,N_5222,N_5172);
nor U6022 (N_6022,N_4963,N_5039);
or U6023 (N_6023,N_5368,N_5531);
xor U6024 (N_6024,N_4914,N_5164);
nand U6025 (N_6025,N_4959,N_5461);
or U6026 (N_6026,N_4952,N_5022);
and U6027 (N_6027,N_5117,N_4996);
and U6028 (N_6028,N_5355,N_5149);
or U6029 (N_6029,N_5007,N_4958);
or U6030 (N_6030,N_5154,N_5070);
xnor U6031 (N_6031,N_5045,N_5398);
xor U6032 (N_6032,N_4814,N_5290);
or U6033 (N_6033,N_5162,N_5274);
nand U6034 (N_6034,N_4846,N_5430);
nand U6035 (N_6035,N_5389,N_4900);
and U6036 (N_6036,N_4883,N_5502);
and U6037 (N_6037,N_5594,N_5059);
nor U6038 (N_6038,N_5576,N_4850);
or U6039 (N_6039,N_4848,N_5330);
nand U6040 (N_6040,N_5493,N_5343);
and U6041 (N_6041,N_4839,N_5555);
and U6042 (N_6042,N_5044,N_5053);
nor U6043 (N_6043,N_5368,N_5553);
nand U6044 (N_6044,N_5068,N_5064);
xnor U6045 (N_6045,N_5301,N_5196);
and U6046 (N_6046,N_5182,N_5546);
or U6047 (N_6047,N_4837,N_5398);
nand U6048 (N_6048,N_5538,N_5504);
xnor U6049 (N_6049,N_5410,N_5558);
xor U6050 (N_6050,N_4825,N_4808);
and U6051 (N_6051,N_4876,N_5110);
nor U6052 (N_6052,N_5564,N_5537);
and U6053 (N_6053,N_5324,N_5331);
xor U6054 (N_6054,N_5262,N_5043);
and U6055 (N_6055,N_5224,N_5506);
xnor U6056 (N_6056,N_4851,N_5457);
nand U6057 (N_6057,N_5325,N_4954);
or U6058 (N_6058,N_5293,N_4919);
and U6059 (N_6059,N_5506,N_5200);
nand U6060 (N_6060,N_5125,N_5063);
xor U6061 (N_6061,N_5328,N_4868);
or U6062 (N_6062,N_4812,N_4950);
xor U6063 (N_6063,N_5139,N_4899);
nor U6064 (N_6064,N_5381,N_5203);
and U6065 (N_6065,N_5521,N_5497);
xor U6066 (N_6066,N_5073,N_5449);
nand U6067 (N_6067,N_4977,N_4964);
xor U6068 (N_6068,N_4867,N_5263);
nand U6069 (N_6069,N_5013,N_5569);
nand U6070 (N_6070,N_4995,N_5145);
nor U6071 (N_6071,N_5409,N_5493);
nor U6072 (N_6072,N_5219,N_5213);
or U6073 (N_6073,N_5172,N_5452);
xnor U6074 (N_6074,N_5587,N_5373);
nor U6075 (N_6075,N_4900,N_5180);
nor U6076 (N_6076,N_4958,N_5567);
and U6077 (N_6077,N_4913,N_5586);
xnor U6078 (N_6078,N_4900,N_5007);
or U6079 (N_6079,N_5302,N_5287);
xnor U6080 (N_6080,N_4991,N_4871);
nor U6081 (N_6081,N_4992,N_5181);
nor U6082 (N_6082,N_4972,N_5552);
nand U6083 (N_6083,N_5585,N_5163);
xor U6084 (N_6084,N_5524,N_4819);
nor U6085 (N_6085,N_4966,N_4932);
and U6086 (N_6086,N_5360,N_5423);
nand U6087 (N_6087,N_5398,N_4834);
and U6088 (N_6088,N_5252,N_5420);
or U6089 (N_6089,N_4889,N_5264);
nand U6090 (N_6090,N_5395,N_4850);
nand U6091 (N_6091,N_5534,N_5289);
xor U6092 (N_6092,N_5027,N_5343);
or U6093 (N_6093,N_4928,N_5146);
xor U6094 (N_6094,N_5032,N_5035);
and U6095 (N_6095,N_5404,N_5362);
and U6096 (N_6096,N_4869,N_4945);
and U6097 (N_6097,N_5565,N_4800);
nor U6098 (N_6098,N_5557,N_5385);
nand U6099 (N_6099,N_5274,N_5529);
xnor U6100 (N_6100,N_4879,N_5569);
nor U6101 (N_6101,N_4838,N_5027);
nand U6102 (N_6102,N_5340,N_5097);
nor U6103 (N_6103,N_5493,N_4983);
or U6104 (N_6104,N_5518,N_5370);
nand U6105 (N_6105,N_5275,N_4969);
nor U6106 (N_6106,N_4932,N_4844);
nand U6107 (N_6107,N_5472,N_5573);
nand U6108 (N_6108,N_5139,N_4814);
xnor U6109 (N_6109,N_5313,N_5214);
and U6110 (N_6110,N_5082,N_5185);
nor U6111 (N_6111,N_4845,N_5360);
xnor U6112 (N_6112,N_5598,N_5387);
xnor U6113 (N_6113,N_4876,N_5511);
nor U6114 (N_6114,N_4983,N_5549);
and U6115 (N_6115,N_5361,N_5104);
or U6116 (N_6116,N_5504,N_5204);
xnor U6117 (N_6117,N_5060,N_4801);
and U6118 (N_6118,N_4922,N_5342);
and U6119 (N_6119,N_4990,N_5045);
nand U6120 (N_6120,N_5080,N_4949);
nor U6121 (N_6121,N_4819,N_5560);
nand U6122 (N_6122,N_4934,N_5445);
nand U6123 (N_6123,N_4838,N_5531);
nand U6124 (N_6124,N_4847,N_5577);
xor U6125 (N_6125,N_5073,N_5017);
nor U6126 (N_6126,N_5258,N_4803);
xor U6127 (N_6127,N_5308,N_4903);
or U6128 (N_6128,N_5521,N_5319);
nor U6129 (N_6129,N_5237,N_4892);
nand U6130 (N_6130,N_5552,N_4989);
and U6131 (N_6131,N_5563,N_4831);
or U6132 (N_6132,N_5358,N_4812);
or U6133 (N_6133,N_4894,N_5041);
nor U6134 (N_6134,N_5140,N_5160);
xnor U6135 (N_6135,N_5135,N_5021);
nor U6136 (N_6136,N_4838,N_5030);
nand U6137 (N_6137,N_5251,N_4910);
and U6138 (N_6138,N_5151,N_5227);
nand U6139 (N_6139,N_5414,N_5098);
and U6140 (N_6140,N_5569,N_5067);
nor U6141 (N_6141,N_5339,N_5457);
and U6142 (N_6142,N_5445,N_4944);
xor U6143 (N_6143,N_4938,N_4929);
nand U6144 (N_6144,N_4833,N_5270);
or U6145 (N_6145,N_4851,N_4985);
and U6146 (N_6146,N_4890,N_5474);
xnor U6147 (N_6147,N_5276,N_5277);
nor U6148 (N_6148,N_4890,N_5015);
xor U6149 (N_6149,N_5094,N_4921);
and U6150 (N_6150,N_5237,N_5459);
nand U6151 (N_6151,N_5089,N_5109);
nor U6152 (N_6152,N_5084,N_4890);
and U6153 (N_6153,N_5111,N_5101);
nand U6154 (N_6154,N_5516,N_5337);
or U6155 (N_6155,N_5441,N_5492);
xnor U6156 (N_6156,N_5505,N_4823);
or U6157 (N_6157,N_5375,N_5054);
or U6158 (N_6158,N_5257,N_5178);
and U6159 (N_6159,N_5581,N_5455);
xnor U6160 (N_6160,N_5106,N_5355);
or U6161 (N_6161,N_5181,N_5155);
or U6162 (N_6162,N_4911,N_4815);
xnor U6163 (N_6163,N_4931,N_5385);
and U6164 (N_6164,N_5567,N_5170);
nor U6165 (N_6165,N_5501,N_5386);
nand U6166 (N_6166,N_4916,N_5279);
or U6167 (N_6167,N_5018,N_5201);
nor U6168 (N_6168,N_5578,N_5266);
or U6169 (N_6169,N_5349,N_5220);
or U6170 (N_6170,N_5086,N_4966);
nor U6171 (N_6171,N_5358,N_5423);
nor U6172 (N_6172,N_5393,N_5349);
nor U6173 (N_6173,N_5251,N_5479);
nand U6174 (N_6174,N_4963,N_5206);
nand U6175 (N_6175,N_5320,N_5074);
xor U6176 (N_6176,N_4817,N_5519);
and U6177 (N_6177,N_4884,N_5288);
or U6178 (N_6178,N_5439,N_5145);
and U6179 (N_6179,N_4935,N_5231);
xor U6180 (N_6180,N_5279,N_5316);
nor U6181 (N_6181,N_5075,N_4879);
or U6182 (N_6182,N_4846,N_5299);
or U6183 (N_6183,N_5364,N_5484);
and U6184 (N_6184,N_5445,N_5181);
xnor U6185 (N_6185,N_5299,N_5451);
nor U6186 (N_6186,N_4935,N_4866);
nand U6187 (N_6187,N_5291,N_5269);
nand U6188 (N_6188,N_5468,N_4927);
or U6189 (N_6189,N_5422,N_5515);
xnor U6190 (N_6190,N_5465,N_5329);
and U6191 (N_6191,N_5533,N_5022);
nor U6192 (N_6192,N_5332,N_5085);
or U6193 (N_6193,N_5352,N_5228);
nor U6194 (N_6194,N_5444,N_5150);
or U6195 (N_6195,N_5472,N_5034);
nand U6196 (N_6196,N_4927,N_5452);
xnor U6197 (N_6197,N_5029,N_5199);
and U6198 (N_6198,N_5062,N_4990);
nand U6199 (N_6199,N_5188,N_5148);
and U6200 (N_6200,N_5063,N_4931);
and U6201 (N_6201,N_4999,N_5250);
nand U6202 (N_6202,N_5355,N_4980);
nor U6203 (N_6203,N_5372,N_5081);
and U6204 (N_6204,N_4925,N_5548);
nand U6205 (N_6205,N_4957,N_5017);
nand U6206 (N_6206,N_5412,N_4985);
xnor U6207 (N_6207,N_4982,N_5266);
or U6208 (N_6208,N_5033,N_5502);
and U6209 (N_6209,N_5050,N_5560);
nor U6210 (N_6210,N_5020,N_5351);
xnor U6211 (N_6211,N_4816,N_5123);
xnor U6212 (N_6212,N_4866,N_5233);
nand U6213 (N_6213,N_5594,N_5364);
xor U6214 (N_6214,N_5200,N_5271);
nor U6215 (N_6215,N_5439,N_5429);
nor U6216 (N_6216,N_5190,N_5418);
nand U6217 (N_6217,N_4900,N_4840);
nand U6218 (N_6218,N_5393,N_5479);
or U6219 (N_6219,N_4866,N_5370);
or U6220 (N_6220,N_5412,N_4918);
nand U6221 (N_6221,N_5347,N_5517);
xor U6222 (N_6222,N_5475,N_4925);
nor U6223 (N_6223,N_5450,N_5096);
or U6224 (N_6224,N_5235,N_4871);
and U6225 (N_6225,N_5075,N_4924);
nor U6226 (N_6226,N_5014,N_4912);
and U6227 (N_6227,N_4979,N_5155);
nor U6228 (N_6228,N_5596,N_5132);
nand U6229 (N_6229,N_4871,N_4806);
xnor U6230 (N_6230,N_5065,N_5408);
nand U6231 (N_6231,N_4874,N_5402);
xnor U6232 (N_6232,N_5103,N_5123);
and U6233 (N_6233,N_5425,N_5540);
xor U6234 (N_6234,N_5583,N_4988);
nand U6235 (N_6235,N_5366,N_5471);
or U6236 (N_6236,N_5127,N_5555);
and U6237 (N_6237,N_4901,N_4846);
and U6238 (N_6238,N_5550,N_5188);
and U6239 (N_6239,N_5472,N_5075);
and U6240 (N_6240,N_5311,N_4922);
xor U6241 (N_6241,N_5289,N_5227);
nand U6242 (N_6242,N_5201,N_4929);
nand U6243 (N_6243,N_4909,N_5478);
and U6244 (N_6244,N_5084,N_5230);
nand U6245 (N_6245,N_4858,N_5232);
nand U6246 (N_6246,N_5052,N_5470);
nor U6247 (N_6247,N_4895,N_5096);
nand U6248 (N_6248,N_4935,N_5122);
or U6249 (N_6249,N_5210,N_5212);
nor U6250 (N_6250,N_4985,N_5358);
xor U6251 (N_6251,N_5255,N_5029);
nand U6252 (N_6252,N_5110,N_5003);
nand U6253 (N_6253,N_5588,N_5398);
nor U6254 (N_6254,N_5144,N_5001);
xnor U6255 (N_6255,N_4801,N_5238);
nand U6256 (N_6256,N_5365,N_4838);
and U6257 (N_6257,N_5155,N_5056);
or U6258 (N_6258,N_4973,N_5355);
nor U6259 (N_6259,N_4818,N_5038);
and U6260 (N_6260,N_4949,N_5293);
xnor U6261 (N_6261,N_4898,N_4940);
or U6262 (N_6262,N_5527,N_5061);
nor U6263 (N_6263,N_5518,N_5190);
or U6264 (N_6264,N_5478,N_5075);
nor U6265 (N_6265,N_5508,N_4855);
nor U6266 (N_6266,N_5562,N_5446);
or U6267 (N_6267,N_4891,N_5056);
nand U6268 (N_6268,N_5029,N_5031);
and U6269 (N_6269,N_5191,N_4901);
nand U6270 (N_6270,N_5428,N_4918);
and U6271 (N_6271,N_5424,N_4840);
or U6272 (N_6272,N_5490,N_5141);
or U6273 (N_6273,N_5126,N_5429);
xor U6274 (N_6274,N_5057,N_4877);
nand U6275 (N_6275,N_5369,N_5088);
nand U6276 (N_6276,N_5175,N_4874);
xnor U6277 (N_6277,N_5037,N_5459);
or U6278 (N_6278,N_5252,N_5539);
nor U6279 (N_6279,N_5489,N_5341);
and U6280 (N_6280,N_5225,N_5317);
and U6281 (N_6281,N_4829,N_4801);
or U6282 (N_6282,N_4910,N_5587);
nand U6283 (N_6283,N_5593,N_5154);
and U6284 (N_6284,N_5404,N_5168);
or U6285 (N_6285,N_5258,N_5262);
and U6286 (N_6286,N_5414,N_5183);
or U6287 (N_6287,N_5432,N_5091);
xor U6288 (N_6288,N_5389,N_4808);
nor U6289 (N_6289,N_4963,N_5555);
nor U6290 (N_6290,N_5325,N_5489);
or U6291 (N_6291,N_5111,N_4923);
and U6292 (N_6292,N_5115,N_5167);
nor U6293 (N_6293,N_4828,N_5211);
or U6294 (N_6294,N_5187,N_4890);
nor U6295 (N_6295,N_5185,N_5021);
xor U6296 (N_6296,N_5256,N_5442);
or U6297 (N_6297,N_5291,N_4855);
or U6298 (N_6298,N_5076,N_5000);
xor U6299 (N_6299,N_4859,N_5226);
xor U6300 (N_6300,N_5073,N_4819);
and U6301 (N_6301,N_5512,N_5393);
or U6302 (N_6302,N_5215,N_5237);
and U6303 (N_6303,N_5370,N_5475);
xnor U6304 (N_6304,N_5061,N_5412);
nor U6305 (N_6305,N_5053,N_5183);
or U6306 (N_6306,N_4849,N_5169);
and U6307 (N_6307,N_4856,N_4887);
nand U6308 (N_6308,N_5076,N_5110);
nand U6309 (N_6309,N_5438,N_5239);
nand U6310 (N_6310,N_5501,N_5037);
and U6311 (N_6311,N_4921,N_5194);
or U6312 (N_6312,N_5222,N_5418);
or U6313 (N_6313,N_5284,N_5168);
xor U6314 (N_6314,N_5312,N_5519);
nand U6315 (N_6315,N_5016,N_4806);
nor U6316 (N_6316,N_5498,N_5038);
and U6317 (N_6317,N_4899,N_5013);
nand U6318 (N_6318,N_5146,N_4829);
and U6319 (N_6319,N_5317,N_4834);
nand U6320 (N_6320,N_5081,N_5336);
nor U6321 (N_6321,N_5453,N_5193);
nor U6322 (N_6322,N_5371,N_5313);
nor U6323 (N_6323,N_5160,N_5352);
nand U6324 (N_6324,N_4875,N_4820);
nand U6325 (N_6325,N_4856,N_5454);
nor U6326 (N_6326,N_5101,N_4945);
nand U6327 (N_6327,N_4964,N_5340);
or U6328 (N_6328,N_5291,N_5123);
xnor U6329 (N_6329,N_4910,N_5241);
or U6330 (N_6330,N_5488,N_5424);
xor U6331 (N_6331,N_4832,N_5402);
and U6332 (N_6332,N_4980,N_4931);
or U6333 (N_6333,N_4975,N_4973);
nand U6334 (N_6334,N_4827,N_5103);
nor U6335 (N_6335,N_5468,N_5037);
nor U6336 (N_6336,N_5495,N_5130);
nand U6337 (N_6337,N_5197,N_5468);
nor U6338 (N_6338,N_5001,N_4974);
and U6339 (N_6339,N_5023,N_5309);
nor U6340 (N_6340,N_4841,N_5070);
and U6341 (N_6341,N_5415,N_5441);
xor U6342 (N_6342,N_5083,N_5448);
nand U6343 (N_6343,N_5518,N_4846);
nor U6344 (N_6344,N_5097,N_5392);
and U6345 (N_6345,N_4962,N_5465);
nand U6346 (N_6346,N_5553,N_5006);
nor U6347 (N_6347,N_5583,N_4929);
nand U6348 (N_6348,N_5035,N_5306);
nor U6349 (N_6349,N_5263,N_5497);
nor U6350 (N_6350,N_5210,N_5436);
or U6351 (N_6351,N_5376,N_4887);
nor U6352 (N_6352,N_5534,N_4946);
nand U6353 (N_6353,N_5043,N_5317);
nor U6354 (N_6354,N_4814,N_5246);
nor U6355 (N_6355,N_5290,N_4888);
or U6356 (N_6356,N_5335,N_5374);
nand U6357 (N_6357,N_5124,N_4961);
or U6358 (N_6358,N_4965,N_5010);
nand U6359 (N_6359,N_4985,N_5507);
or U6360 (N_6360,N_4860,N_5365);
or U6361 (N_6361,N_5466,N_5424);
or U6362 (N_6362,N_4879,N_5336);
nand U6363 (N_6363,N_4896,N_5305);
nand U6364 (N_6364,N_4875,N_4834);
or U6365 (N_6365,N_5072,N_5384);
nand U6366 (N_6366,N_5587,N_4916);
xor U6367 (N_6367,N_5231,N_5111);
xnor U6368 (N_6368,N_4872,N_5206);
xor U6369 (N_6369,N_5381,N_5537);
nor U6370 (N_6370,N_4828,N_4845);
xor U6371 (N_6371,N_5314,N_5220);
nor U6372 (N_6372,N_5172,N_5292);
xor U6373 (N_6373,N_5361,N_5154);
and U6374 (N_6374,N_5517,N_4883);
or U6375 (N_6375,N_5057,N_5411);
nor U6376 (N_6376,N_4866,N_5398);
and U6377 (N_6377,N_4984,N_4912);
nand U6378 (N_6378,N_4815,N_4979);
or U6379 (N_6379,N_4983,N_5423);
and U6380 (N_6380,N_5274,N_4845);
xor U6381 (N_6381,N_5349,N_5258);
xor U6382 (N_6382,N_5196,N_5310);
nand U6383 (N_6383,N_5472,N_5190);
nand U6384 (N_6384,N_4883,N_4814);
nor U6385 (N_6385,N_4801,N_5484);
xnor U6386 (N_6386,N_4918,N_5171);
nor U6387 (N_6387,N_5513,N_4832);
or U6388 (N_6388,N_5109,N_5029);
or U6389 (N_6389,N_5307,N_5341);
xnor U6390 (N_6390,N_5270,N_4935);
nand U6391 (N_6391,N_5167,N_5378);
nand U6392 (N_6392,N_5251,N_5325);
and U6393 (N_6393,N_4801,N_4840);
nor U6394 (N_6394,N_5130,N_4905);
xor U6395 (N_6395,N_5149,N_5542);
nor U6396 (N_6396,N_5410,N_5488);
xnor U6397 (N_6397,N_5120,N_4969);
or U6398 (N_6398,N_5168,N_4908);
nor U6399 (N_6399,N_5595,N_5325);
xor U6400 (N_6400,N_6068,N_5650);
or U6401 (N_6401,N_6010,N_5920);
nor U6402 (N_6402,N_5791,N_6289);
nand U6403 (N_6403,N_6374,N_6067);
nand U6404 (N_6404,N_6369,N_6000);
xnor U6405 (N_6405,N_6300,N_6230);
and U6406 (N_6406,N_6207,N_6310);
xnor U6407 (N_6407,N_6364,N_6034);
nand U6408 (N_6408,N_5667,N_6383);
nand U6409 (N_6409,N_6328,N_6027);
or U6410 (N_6410,N_5632,N_5910);
or U6411 (N_6411,N_6016,N_5918);
or U6412 (N_6412,N_6317,N_6339);
xnor U6413 (N_6413,N_5831,N_5890);
nand U6414 (N_6414,N_6201,N_5685);
and U6415 (N_6415,N_6170,N_5848);
xor U6416 (N_6416,N_6345,N_6274);
nand U6417 (N_6417,N_6244,N_6265);
or U6418 (N_6418,N_5929,N_5767);
and U6419 (N_6419,N_6280,N_6299);
xor U6420 (N_6420,N_5675,N_5949);
and U6421 (N_6421,N_5972,N_6281);
nand U6422 (N_6422,N_5859,N_5936);
nand U6423 (N_6423,N_6053,N_6368);
and U6424 (N_6424,N_5677,N_6162);
xor U6425 (N_6425,N_5905,N_6298);
nand U6426 (N_6426,N_6312,N_5790);
nand U6427 (N_6427,N_6257,N_5997);
or U6428 (N_6428,N_6022,N_6371);
xnor U6429 (N_6429,N_5935,N_6071);
nand U6430 (N_6430,N_5840,N_5817);
nand U6431 (N_6431,N_5656,N_5653);
nor U6432 (N_6432,N_6247,N_6321);
xor U6433 (N_6433,N_6182,N_6133);
nand U6434 (N_6434,N_6065,N_5953);
nand U6435 (N_6435,N_6164,N_5960);
and U6436 (N_6436,N_6059,N_5721);
and U6437 (N_6437,N_5925,N_5627);
xnor U6438 (N_6438,N_5928,N_5658);
or U6439 (N_6439,N_6212,N_5850);
nand U6440 (N_6440,N_6017,N_5891);
xor U6441 (N_6441,N_6268,N_6101);
nand U6442 (N_6442,N_5605,N_5993);
or U6443 (N_6443,N_5815,N_5734);
nand U6444 (N_6444,N_5630,N_6040);
nor U6445 (N_6445,N_6278,N_6066);
nor U6446 (N_6446,N_6200,N_6116);
nor U6447 (N_6447,N_5718,N_5603);
xor U6448 (N_6448,N_6377,N_6325);
nand U6449 (N_6449,N_5607,N_6052);
nor U6450 (N_6450,N_5780,N_6018);
nor U6451 (N_6451,N_6287,N_6106);
and U6452 (N_6452,N_6097,N_6256);
nor U6453 (N_6453,N_5646,N_6284);
and U6454 (N_6454,N_5865,N_5713);
nor U6455 (N_6455,N_6114,N_6081);
nor U6456 (N_6456,N_5720,N_5678);
nand U6457 (N_6457,N_6211,N_6054);
nor U6458 (N_6458,N_6096,N_5893);
nor U6459 (N_6459,N_6141,N_5947);
or U6460 (N_6460,N_6179,N_5971);
or U6461 (N_6461,N_6224,N_5946);
and U6462 (N_6462,N_6183,N_6095);
or U6463 (N_6463,N_5937,N_5857);
nor U6464 (N_6464,N_5714,N_5979);
nand U6465 (N_6465,N_6286,N_6142);
xor U6466 (N_6466,N_5619,N_5730);
xor U6467 (N_6467,N_6235,N_5797);
xnor U6468 (N_6468,N_6214,N_5670);
nor U6469 (N_6469,N_5832,N_6005);
or U6470 (N_6470,N_5680,N_5862);
xnor U6471 (N_6471,N_6050,N_6174);
nand U6472 (N_6472,N_5980,N_5965);
nor U6473 (N_6473,N_6329,N_5833);
and U6474 (N_6474,N_5834,N_5793);
xnor U6475 (N_6475,N_6283,N_6367);
nor U6476 (N_6476,N_5835,N_6159);
and U6477 (N_6477,N_5940,N_6226);
xor U6478 (N_6478,N_6213,N_5813);
or U6479 (N_6479,N_6245,N_6242);
nand U6480 (N_6480,N_6015,N_5736);
nor U6481 (N_6481,N_6083,N_5768);
nor U6482 (N_6482,N_5753,N_5687);
or U6483 (N_6483,N_6397,N_5784);
and U6484 (N_6484,N_6236,N_6243);
and U6485 (N_6485,N_6175,N_6026);
or U6486 (N_6486,N_6234,N_6056);
nand U6487 (N_6487,N_6176,N_5970);
and U6488 (N_6488,N_6398,N_6252);
nor U6489 (N_6489,N_6172,N_5717);
nand U6490 (N_6490,N_5846,N_6294);
and U6491 (N_6491,N_5877,N_5726);
nand U6492 (N_6492,N_6125,N_5967);
or U6493 (N_6493,N_5629,N_6119);
xnor U6494 (N_6494,N_5623,N_5694);
xnor U6495 (N_6495,N_5864,N_5727);
or U6496 (N_6496,N_6131,N_5858);
nor U6497 (N_6497,N_6113,N_5961);
nand U6498 (N_6498,N_6382,N_6057);
xor U6499 (N_6499,N_6137,N_6269);
xnor U6500 (N_6500,N_5991,N_5776);
xnor U6501 (N_6501,N_5917,N_6177);
nand U6502 (N_6502,N_6145,N_6228);
xor U6503 (N_6503,N_5869,N_5651);
xnor U6504 (N_6504,N_6266,N_6080);
nand U6505 (N_6505,N_5686,N_5769);
or U6506 (N_6506,N_6277,N_5710);
xnor U6507 (N_6507,N_6203,N_6042);
and U6508 (N_6508,N_6324,N_5676);
nand U6509 (N_6509,N_6044,N_6102);
xnor U6510 (N_6510,N_6360,N_5824);
nor U6511 (N_6511,N_6115,N_6033);
and U6512 (N_6512,N_6253,N_5954);
and U6513 (N_6513,N_5948,N_6046);
and U6514 (N_6514,N_5887,N_5661);
and U6515 (N_6515,N_5735,N_5889);
or U6516 (N_6516,N_6394,N_5693);
and U6517 (N_6517,N_6273,N_6149);
xor U6518 (N_6518,N_6351,N_5707);
and U6519 (N_6519,N_5702,N_5963);
or U6520 (N_6520,N_5641,N_5919);
and U6521 (N_6521,N_5986,N_6297);
or U6522 (N_6522,N_5748,N_5913);
or U6523 (N_6523,N_6388,N_6144);
nor U6524 (N_6524,N_6334,N_6396);
nor U6525 (N_6525,N_5803,N_5932);
nor U6526 (N_6526,N_5825,N_6169);
xnor U6527 (N_6527,N_5900,N_5778);
or U6528 (N_6528,N_6073,N_6121);
or U6529 (N_6529,N_6094,N_5912);
xor U6530 (N_6530,N_5634,N_5657);
nor U6531 (N_6531,N_5942,N_5615);
and U6532 (N_6532,N_5655,N_5724);
nand U6533 (N_6533,N_6237,N_5620);
and U6534 (N_6534,N_6204,N_6304);
xnor U6535 (N_6535,N_6129,N_6028);
or U6536 (N_6536,N_5716,N_6276);
nor U6537 (N_6537,N_5841,N_5959);
nor U6538 (N_6538,N_6373,N_5851);
nand U6539 (N_6539,N_6032,N_6258);
nand U6540 (N_6540,N_5943,N_5847);
xnor U6541 (N_6541,N_6002,N_6075);
nand U6542 (N_6542,N_6047,N_6140);
xor U6543 (N_6543,N_5766,N_5795);
nor U6544 (N_6544,N_5617,N_5941);
and U6545 (N_6545,N_5985,N_6039);
nor U6546 (N_6546,N_6215,N_5772);
and U6547 (N_6547,N_5637,N_5894);
nand U6548 (N_6548,N_5749,N_5806);
nor U6549 (N_6549,N_6348,N_5888);
and U6550 (N_6550,N_5875,N_5868);
nor U6551 (N_6551,N_5944,N_6126);
or U6552 (N_6552,N_5808,N_6156);
or U6553 (N_6553,N_5684,N_6217);
nand U6554 (N_6554,N_6337,N_5699);
or U6555 (N_6555,N_5951,N_5731);
xor U6556 (N_6556,N_5878,N_5810);
nand U6557 (N_6557,N_5628,N_5647);
nor U6558 (N_6558,N_5799,N_5770);
and U6559 (N_6559,N_5861,N_5642);
or U6560 (N_6560,N_6161,N_5897);
or U6561 (N_6561,N_6363,N_5981);
xor U6562 (N_6562,N_6086,N_5988);
xnor U6563 (N_6563,N_6338,N_5994);
or U6564 (N_6564,N_5837,N_6282);
or U6565 (N_6565,N_6138,N_5649);
nor U6566 (N_6566,N_5669,N_5785);
xor U6567 (N_6567,N_5755,N_6271);
and U6568 (N_6568,N_5990,N_6134);
and U6569 (N_6569,N_5921,N_5923);
xor U6570 (N_6570,N_6186,N_6238);
nand U6571 (N_6571,N_6158,N_5672);
or U6572 (N_6572,N_6370,N_5836);
nor U6573 (N_6573,N_6255,N_6185);
or U6574 (N_6574,N_6036,N_5924);
nand U6575 (N_6575,N_6232,N_6350);
xnor U6576 (N_6576,N_5758,N_6030);
nor U6577 (N_6577,N_5922,N_6381);
and U6578 (N_6578,N_6108,N_6051);
xnor U6579 (N_6579,N_6320,N_5608);
or U6580 (N_6580,N_6199,N_6390);
or U6581 (N_6581,N_6393,N_6288);
and U6582 (N_6582,N_5728,N_5779);
nor U6583 (N_6583,N_5674,N_5800);
nor U6584 (N_6584,N_5783,N_5622);
xnor U6585 (N_6585,N_5618,N_5606);
or U6586 (N_6586,N_5939,N_5759);
xor U6587 (N_6587,N_6391,N_5855);
and U6588 (N_6588,N_6260,N_5998);
nor U6589 (N_6589,N_5660,N_5663);
and U6590 (N_6590,N_5955,N_6181);
xnor U6591 (N_6591,N_6089,N_5640);
xor U6592 (N_6592,N_5654,N_6092);
nor U6593 (N_6593,N_5982,N_5635);
nor U6594 (N_6594,N_6303,N_5743);
or U6595 (N_6595,N_6352,N_5867);
xnor U6596 (N_6596,N_5816,N_5818);
xnor U6597 (N_6597,N_5984,N_5931);
xor U6598 (N_6598,N_5908,N_6006);
or U6599 (N_6599,N_5911,N_6385);
and U6600 (N_6600,N_6190,N_5898);
and U6601 (N_6601,N_5754,N_5819);
and U6602 (N_6602,N_6103,N_5631);
nand U6603 (N_6603,N_6167,N_5742);
and U6604 (N_6604,N_6384,N_6130);
or U6605 (N_6605,N_5788,N_6091);
or U6606 (N_6606,N_5609,N_5823);
nand U6607 (N_6607,N_6291,N_6305);
xnor U6608 (N_6608,N_5652,N_5828);
or U6609 (N_6609,N_6014,N_5934);
and U6610 (N_6610,N_5762,N_5659);
nor U6611 (N_6611,N_6151,N_6392);
xnor U6612 (N_6612,N_6023,N_5916);
nor U6613 (N_6613,N_5826,N_6219);
nand U6614 (N_6614,N_6187,N_5977);
nand U6615 (N_6615,N_6117,N_5611);
nand U6616 (N_6616,N_6254,N_6275);
nand U6617 (N_6617,N_6031,N_6038);
nor U6618 (N_6618,N_6229,N_6007);
xor U6619 (N_6619,N_6074,N_6262);
and U6620 (N_6620,N_5668,N_5950);
nor U6621 (N_6621,N_6314,N_6165);
nor U6622 (N_6622,N_5610,N_6353);
nor U6623 (N_6623,N_5625,N_6222);
or U6624 (N_6624,N_5933,N_6020);
nand U6625 (N_6625,N_5761,N_5787);
or U6626 (N_6626,N_6099,N_6296);
or U6627 (N_6627,N_5899,N_6013);
nand U6628 (N_6628,N_5976,N_6209);
nand U6629 (N_6629,N_6048,N_5804);
or U6630 (N_6630,N_5673,N_5792);
nand U6631 (N_6631,N_6315,N_6198);
xnor U6632 (N_6632,N_5771,N_5822);
xnor U6633 (N_6633,N_6154,N_5821);
and U6634 (N_6634,N_6062,N_5741);
nor U6635 (N_6635,N_5626,N_6316);
nor U6636 (N_6636,N_6399,N_5740);
and U6637 (N_6637,N_6358,N_6157);
xor U6638 (N_6638,N_6021,N_5705);
nor U6639 (N_6639,N_6330,N_6264);
and U6640 (N_6640,N_6221,N_6009);
nand U6641 (N_6641,N_6064,N_6387);
or U6642 (N_6642,N_5969,N_5706);
and U6643 (N_6643,N_5958,N_6136);
nand U6644 (N_6644,N_5957,N_6123);
xor U6645 (N_6645,N_5695,N_5895);
xor U6646 (N_6646,N_6118,N_5689);
and U6647 (N_6647,N_6347,N_6318);
and U6648 (N_6648,N_6069,N_6376);
nand U6649 (N_6649,N_5722,N_5995);
nor U6650 (N_6650,N_6354,N_6272);
xor U6651 (N_6651,N_6061,N_5633);
nand U6652 (N_6652,N_6340,N_6146);
and U6653 (N_6653,N_5830,N_6076);
and U6654 (N_6654,N_5756,N_6223);
nand U6655 (N_6655,N_6210,N_6389);
nor U6656 (N_6656,N_6292,N_6395);
xnor U6657 (N_6657,N_5664,N_6218);
nand U6658 (N_6658,N_6202,N_5812);
and U6659 (N_6659,N_6361,N_5719);
and U6660 (N_6660,N_6105,N_5885);
nor U6661 (N_6661,N_5996,N_5600);
and U6662 (N_6662,N_6220,N_5765);
xnor U6663 (N_6663,N_6309,N_5733);
xnor U6664 (N_6664,N_5854,N_6122);
nand U6665 (N_6665,N_5945,N_6196);
and U6666 (N_6666,N_6035,N_5901);
xor U6667 (N_6667,N_5704,N_5691);
and U6668 (N_6668,N_6319,N_5644);
or U6669 (N_6669,N_5802,N_6155);
nor U6670 (N_6670,N_5681,N_6152);
or U6671 (N_6671,N_6285,N_5809);
and U6672 (N_6672,N_6024,N_6343);
nor U6673 (N_6673,N_6093,N_6249);
or U6674 (N_6674,N_5956,N_5838);
or U6675 (N_6675,N_5968,N_5729);
nand U6676 (N_6676,N_6111,N_6060);
nor U6677 (N_6677,N_5915,N_6263);
or U6678 (N_6678,N_6072,N_5866);
xor U6679 (N_6679,N_6191,N_6104);
or U6680 (N_6680,N_6380,N_6239);
xnor U6681 (N_6681,N_5786,N_5973);
nand U6682 (N_6682,N_6331,N_6100);
nand U6683 (N_6683,N_5870,N_5814);
and U6684 (N_6684,N_5930,N_6045);
nor U6685 (N_6685,N_6098,N_5872);
nand U6686 (N_6686,N_6189,N_6326);
or U6687 (N_6687,N_6128,N_5764);
or U6688 (N_6688,N_6240,N_5839);
or U6689 (N_6689,N_6019,N_5671);
xor U6690 (N_6690,N_6206,N_6349);
and U6691 (N_6691,N_5688,N_5796);
xor U6692 (N_6692,N_6084,N_5751);
nor U6693 (N_6693,N_6193,N_5801);
or U6694 (N_6694,N_6077,N_6279);
or U6695 (N_6695,N_5983,N_5978);
or U6696 (N_6696,N_6088,N_5966);
nor U6697 (N_6697,N_6173,N_5880);
nand U6698 (N_6698,N_5781,N_5992);
or U6699 (N_6699,N_6003,N_5698);
nand U6700 (N_6700,N_5909,N_6184);
xnor U6701 (N_6701,N_5974,N_5665);
xor U6702 (N_6702,N_6306,N_5709);
and U6703 (N_6703,N_5914,N_6078);
xor U6704 (N_6704,N_6188,N_6087);
xnor U6705 (N_6705,N_5636,N_5737);
or U6706 (N_6706,N_6225,N_5777);
or U6707 (N_6707,N_6082,N_5679);
nor U6708 (N_6708,N_5849,N_6148);
nand U6709 (N_6709,N_6029,N_5807);
and U6710 (N_6710,N_6063,N_6366);
nand U6711 (N_6711,N_6379,N_6043);
xnor U6712 (N_6712,N_5738,N_6335);
and U6713 (N_6713,N_5752,N_5638);
xnor U6714 (N_6714,N_5906,N_5811);
and U6715 (N_6715,N_6070,N_5798);
and U6716 (N_6716,N_6233,N_6344);
nor U6717 (N_6717,N_5747,N_5842);
xnor U6718 (N_6718,N_5662,N_6313);
or U6719 (N_6719,N_6001,N_5884);
xor U6720 (N_6720,N_5711,N_6246);
xor U6721 (N_6721,N_6375,N_5999);
nor U6722 (N_6722,N_5703,N_5975);
nor U6723 (N_6723,N_6160,N_5856);
xor U6724 (N_6724,N_6251,N_5601);
or U6725 (N_6725,N_5863,N_5883);
xor U6726 (N_6726,N_6341,N_6227);
and U6727 (N_6727,N_5604,N_6132);
nand U6728 (N_6728,N_6012,N_5612);
xor U6729 (N_6729,N_5964,N_5852);
nor U6730 (N_6730,N_6290,N_6205);
xor U6731 (N_6731,N_5682,N_6166);
or U6732 (N_6732,N_5789,N_6308);
and U6733 (N_6733,N_5774,N_6180);
nor U6734 (N_6734,N_6085,N_6231);
nand U6735 (N_6735,N_6124,N_5902);
nor U6736 (N_6736,N_5860,N_6372);
nor U6737 (N_6737,N_5683,N_5645);
nand U6738 (N_6738,N_6386,N_5732);
xnor U6739 (N_6739,N_5746,N_6107);
and U6740 (N_6740,N_5794,N_6311);
or U6741 (N_6741,N_5763,N_5696);
or U6742 (N_6742,N_5614,N_6109);
or U6743 (N_6743,N_5697,N_6295);
nand U6744 (N_6744,N_6362,N_6139);
or U6745 (N_6745,N_5962,N_6127);
nand U6746 (N_6746,N_5775,N_6216);
nor U6747 (N_6747,N_6004,N_6342);
or U6748 (N_6748,N_6110,N_6267);
or U6749 (N_6749,N_6378,N_5616);
xor U6750 (N_6750,N_6336,N_5757);
nor U6751 (N_6751,N_6147,N_5853);
or U6752 (N_6752,N_6049,N_5725);
and U6753 (N_6753,N_6168,N_6055);
nor U6754 (N_6754,N_6143,N_5739);
nand U6755 (N_6755,N_5879,N_6357);
or U6756 (N_6756,N_5701,N_5896);
xor U6757 (N_6757,N_6359,N_5750);
and U6758 (N_6758,N_5648,N_5876);
nand U6759 (N_6759,N_5700,N_5745);
and U6760 (N_6760,N_5874,N_5892);
or U6761 (N_6761,N_5989,N_5666);
xor U6762 (N_6762,N_6355,N_5613);
nand U6763 (N_6763,N_6293,N_6195);
and U6764 (N_6764,N_5882,N_6079);
and U6765 (N_6765,N_6241,N_5871);
or U6766 (N_6766,N_5643,N_5621);
or U6767 (N_6767,N_6356,N_6323);
or U6768 (N_6768,N_5712,N_6041);
and U6769 (N_6769,N_5715,N_5926);
xnor U6770 (N_6770,N_6194,N_6332);
nand U6771 (N_6771,N_5723,N_6192);
xnor U6772 (N_6772,N_6011,N_5881);
and U6773 (N_6773,N_5624,N_6163);
nand U6774 (N_6774,N_6365,N_6025);
and U6775 (N_6775,N_6259,N_6346);
nor U6776 (N_6776,N_6171,N_5903);
and U6777 (N_6777,N_5844,N_5952);
nor U6778 (N_6778,N_5829,N_5845);
and U6779 (N_6779,N_5987,N_6250);
xnor U6780 (N_6780,N_5782,N_5927);
or U6781 (N_6781,N_5744,N_6322);
or U6782 (N_6782,N_5907,N_5805);
nor U6783 (N_6783,N_5639,N_5760);
nand U6784 (N_6784,N_6197,N_5904);
nand U6785 (N_6785,N_6301,N_6037);
xor U6786 (N_6786,N_6120,N_5773);
or U6787 (N_6787,N_6150,N_6058);
xor U6788 (N_6788,N_6248,N_6327);
nand U6789 (N_6789,N_6270,N_5938);
nand U6790 (N_6790,N_6112,N_5690);
xnor U6791 (N_6791,N_5708,N_6261);
nor U6792 (N_6792,N_5820,N_6208);
xnor U6793 (N_6793,N_5827,N_6178);
or U6794 (N_6794,N_6008,N_5886);
nand U6795 (N_6795,N_5873,N_5692);
nand U6796 (N_6796,N_6307,N_6135);
or U6797 (N_6797,N_5602,N_6153);
nor U6798 (N_6798,N_6302,N_6090);
nand U6799 (N_6799,N_6333,N_5843);
or U6800 (N_6800,N_5738,N_6265);
or U6801 (N_6801,N_5747,N_6097);
nand U6802 (N_6802,N_5700,N_5826);
or U6803 (N_6803,N_5964,N_5832);
and U6804 (N_6804,N_6010,N_6189);
nand U6805 (N_6805,N_5997,N_6365);
nor U6806 (N_6806,N_5688,N_6077);
and U6807 (N_6807,N_5759,N_5738);
nor U6808 (N_6808,N_6168,N_6233);
nand U6809 (N_6809,N_5980,N_5889);
or U6810 (N_6810,N_5622,N_5607);
or U6811 (N_6811,N_5949,N_5648);
nor U6812 (N_6812,N_5633,N_6330);
nand U6813 (N_6813,N_6071,N_6063);
nor U6814 (N_6814,N_6317,N_6003);
nand U6815 (N_6815,N_5890,N_5832);
xor U6816 (N_6816,N_6153,N_6013);
or U6817 (N_6817,N_5937,N_6381);
nand U6818 (N_6818,N_6036,N_6178);
and U6819 (N_6819,N_5607,N_5690);
nor U6820 (N_6820,N_5769,N_6334);
nand U6821 (N_6821,N_5748,N_5881);
nand U6822 (N_6822,N_5644,N_5911);
nand U6823 (N_6823,N_6274,N_6367);
or U6824 (N_6824,N_5724,N_5890);
and U6825 (N_6825,N_6124,N_6364);
nand U6826 (N_6826,N_5763,N_6115);
xor U6827 (N_6827,N_5841,N_6021);
and U6828 (N_6828,N_6263,N_6363);
nand U6829 (N_6829,N_5661,N_5679);
and U6830 (N_6830,N_5745,N_5957);
and U6831 (N_6831,N_5713,N_6168);
nor U6832 (N_6832,N_6296,N_6121);
xnor U6833 (N_6833,N_6211,N_5825);
and U6834 (N_6834,N_5860,N_5869);
and U6835 (N_6835,N_6026,N_5858);
nor U6836 (N_6836,N_5819,N_6242);
and U6837 (N_6837,N_6020,N_6039);
xor U6838 (N_6838,N_5948,N_5914);
nand U6839 (N_6839,N_5765,N_5808);
nor U6840 (N_6840,N_6233,N_6297);
xnor U6841 (N_6841,N_5685,N_5627);
or U6842 (N_6842,N_5694,N_6330);
and U6843 (N_6843,N_5648,N_6004);
or U6844 (N_6844,N_5990,N_5973);
nand U6845 (N_6845,N_5826,N_5891);
nor U6846 (N_6846,N_6046,N_6074);
nand U6847 (N_6847,N_5610,N_6135);
xor U6848 (N_6848,N_6087,N_5785);
and U6849 (N_6849,N_5726,N_6312);
and U6850 (N_6850,N_6155,N_5685);
nor U6851 (N_6851,N_5966,N_5601);
nor U6852 (N_6852,N_5732,N_6032);
nand U6853 (N_6853,N_5605,N_5780);
nand U6854 (N_6854,N_6388,N_5902);
nor U6855 (N_6855,N_5757,N_6322);
and U6856 (N_6856,N_6222,N_6190);
xnor U6857 (N_6857,N_6275,N_6026);
xor U6858 (N_6858,N_6280,N_5900);
and U6859 (N_6859,N_6024,N_6359);
or U6860 (N_6860,N_5890,N_6195);
nand U6861 (N_6861,N_6069,N_6324);
nand U6862 (N_6862,N_6144,N_5755);
or U6863 (N_6863,N_6059,N_5984);
nand U6864 (N_6864,N_6312,N_5762);
nor U6865 (N_6865,N_5802,N_5789);
nor U6866 (N_6866,N_6009,N_5956);
nor U6867 (N_6867,N_5796,N_6244);
and U6868 (N_6868,N_6287,N_6163);
and U6869 (N_6869,N_6263,N_6144);
xor U6870 (N_6870,N_6378,N_6318);
nor U6871 (N_6871,N_6172,N_5691);
nand U6872 (N_6872,N_5825,N_6157);
or U6873 (N_6873,N_5912,N_6147);
nor U6874 (N_6874,N_5668,N_5797);
and U6875 (N_6875,N_6022,N_5738);
nor U6876 (N_6876,N_5882,N_6183);
nor U6877 (N_6877,N_5679,N_6095);
nand U6878 (N_6878,N_5769,N_5632);
xor U6879 (N_6879,N_5781,N_5760);
nor U6880 (N_6880,N_6330,N_5666);
nand U6881 (N_6881,N_6083,N_6239);
nor U6882 (N_6882,N_6280,N_5904);
nor U6883 (N_6883,N_6051,N_6163);
nor U6884 (N_6884,N_5897,N_5797);
xor U6885 (N_6885,N_6165,N_6283);
xnor U6886 (N_6886,N_6088,N_6032);
or U6887 (N_6887,N_5733,N_5895);
and U6888 (N_6888,N_5660,N_5892);
or U6889 (N_6889,N_5722,N_5609);
nor U6890 (N_6890,N_5882,N_6366);
xor U6891 (N_6891,N_6392,N_6238);
nor U6892 (N_6892,N_5720,N_5929);
and U6893 (N_6893,N_6235,N_5810);
and U6894 (N_6894,N_5625,N_6262);
and U6895 (N_6895,N_6054,N_6108);
and U6896 (N_6896,N_5781,N_6355);
nand U6897 (N_6897,N_6246,N_6258);
nor U6898 (N_6898,N_6210,N_5722);
nand U6899 (N_6899,N_6112,N_6188);
nand U6900 (N_6900,N_6019,N_6263);
nor U6901 (N_6901,N_6385,N_5618);
nand U6902 (N_6902,N_5978,N_5803);
xnor U6903 (N_6903,N_6022,N_5869);
xnor U6904 (N_6904,N_5867,N_6165);
or U6905 (N_6905,N_5836,N_5704);
nor U6906 (N_6906,N_5895,N_6269);
nor U6907 (N_6907,N_6318,N_5605);
xnor U6908 (N_6908,N_6206,N_6134);
and U6909 (N_6909,N_6162,N_6149);
nand U6910 (N_6910,N_6288,N_6299);
or U6911 (N_6911,N_6231,N_6131);
or U6912 (N_6912,N_5607,N_5632);
or U6913 (N_6913,N_6087,N_6214);
nand U6914 (N_6914,N_6001,N_6299);
or U6915 (N_6915,N_5798,N_5874);
nor U6916 (N_6916,N_6255,N_5745);
and U6917 (N_6917,N_6102,N_6303);
xor U6918 (N_6918,N_6223,N_6068);
xor U6919 (N_6919,N_5684,N_5617);
xnor U6920 (N_6920,N_6079,N_5943);
nor U6921 (N_6921,N_5913,N_5722);
nor U6922 (N_6922,N_6267,N_5853);
nand U6923 (N_6923,N_5828,N_5867);
xor U6924 (N_6924,N_6220,N_5699);
or U6925 (N_6925,N_5815,N_6333);
nor U6926 (N_6926,N_6087,N_6303);
and U6927 (N_6927,N_6127,N_6221);
nor U6928 (N_6928,N_5865,N_5928);
and U6929 (N_6929,N_6033,N_5606);
or U6930 (N_6930,N_5725,N_6076);
or U6931 (N_6931,N_5968,N_5874);
and U6932 (N_6932,N_5995,N_5839);
nor U6933 (N_6933,N_5804,N_6035);
nand U6934 (N_6934,N_5718,N_6385);
xor U6935 (N_6935,N_5691,N_6338);
xor U6936 (N_6936,N_5795,N_6113);
nand U6937 (N_6937,N_5986,N_6052);
and U6938 (N_6938,N_5806,N_6027);
nand U6939 (N_6939,N_6087,N_5714);
nand U6940 (N_6940,N_6347,N_5841);
nor U6941 (N_6941,N_5745,N_5814);
nor U6942 (N_6942,N_5900,N_5838);
nor U6943 (N_6943,N_5922,N_6353);
nand U6944 (N_6944,N_5966,N_6258);
nor U6945 (N_6945,N_5725,N_5777);
and U6946 (N_6946,N_6161,N_5928);
nor U6947 (N_6947,N_5942,N_5871);
and U6948 (N_6948,N_6096,N_5751);
nor U6949 (N_6949,N_5656,N_6314);
nor U6950 (N_6950,N_6036,N_6114);
nand U6951 (N_6951,N_5638,N_6288);
and U6952 (N_6952,N_6351,N_5730);
xnor U6953 (N_6953,N_5786,N_6030);
nand U6954 (N_6954,N_6108,N_5837);
xor U6955 (N_6955,N_6358,N_5976);
nand U6956 (N_6956,N_6204,N_6081);
nand U6957 (N_6957,N_5848,N_6250);
nor U6958 (N_6958,N_6162,N_5785);
and U6959 (N_6959,N_6054,N_5643);
and U6960 (N_6960,N_5703,N_6100);
nor U6961 (N_6961,N_5921,N_6372);
xnor U6962 (N_6962,N_5697,N_5635);
nor U6963 (N_6963,N_6339,N_5913);
and U6964 (N_6964,N_6103,N_6233);
and U6965 (N_6965,N_5831,N_5705);
xor U6966 (N_6966,N_6200,N_5766);
xor U6967 (N_6967,N_6344,N_5847);
nand U6968 (N_6968,N_5681,N_6124);
xnor U6969 (N_6969,N_6107,N_6055);
xor U6970 (N_6970,N_5887,N_5867);
and U6971 (N_6971,N_5743,N_6090);
xor U6972 (N_6972,N_5967,N_5893);
or U6973 (N_6973,N_6306,N_5922);
nand U6974 (N_6974,N_5875,N_6295);
and U6975 (N_6975,N_6073,N_6098);
and U6976 (N_6976,N_5990,N_5600);
or U6977 (N_6977,N_6242,N_5644);
and U6978 (N_6978,N_5958,N_5697);
or U6979 (N_6979,N_5707,N_6122);
or U6980 (N_6980,N_6302,N_6245);
nand U6981 (N_6981,N_5977,N_6077);
or U6982 (N_6982,N_6080,N_6328);
xor U6983 (N_6983,N_6027,N_6197);
xor U6984 (N_6984,N_6103,N_6118);
and U6985 (N_6985,N_5718,N_6341);
and U6986 (N_6986,N_6398,N_5910);
or U6987 (N_6987,N_5857,N_6031);
nor U6988 (N_6988,N_6062,N_5784);
xnor U6989 (N_6989,N_6178,N_5738);
nor U6990 (N_6990,N_5968,N_5911);
nor U6991 (N_6991,N_5927,N_5895);
nor U6992 (N_6992,N_6344,N_5651);
or U6993 (N_6993,N_5630,N_6160);
and U6994 (N_6994,N_6186,N_5627);
xor U6995 (N_6995,N_5985,N_6382);
xnor U6996 (N_6996,N_5969,N_6060);
or U6997 (N_6997,N_5620,N_6293);
nor U6998 (N_6998,N_6121,N_5885);
xnor U6999 (N_6999,N_6137,N_5850);
or U7000 (N_7000,N_5875,N_5624);
xor U7001 (N_7001,N_6164,N_5768);
and U7002 (N_7002,N_5644,N_5701);
or U7003 (N_7003,N_5846,N_5766);
and U7004 (N_7004,N_5920,N_6094);
xnor U7005 (N_7005,N_6350,N_6205);
nor U7006 (N_7006,N_6146,N_5938);
nand U7007 (N_7007,N_5838,N_5682);
xor U7008 (N_7008,N_6393,N_6070);
and U7009 (N_7009,N_6363,N_5715);
and U7010 (N_7010,N_6090,N_5826);
nor U7011 (N_7011,N_5886,N_5921);
nand U7012 (N_7012,N_5983,N_6160);
or U7013 (N_7013,N_6211,N_5625);
xnor U7014 (N_7014,N_5849,N_5749);
nor U7015 (N_7015,N_5916,N_6243);
xnor U7016 (N_7016,N_5955,N_6381);
and U7017 (N_7017,N_5789,N_5739);
xnor U7018 (N_7018,N_5844,N_5757);
nand U7019 (N_7019,N_6172,N_5904);
or U7020 (N_7020,N_6222,N_6343);
nor U7021 (N_7021,N_5612,N_5912);
nor U7022 (N_7022,N_5886,N_5823);
nor U7023 (N_7023,N_5864,N_5866);
nand U7024 (N_7024,N_6350,N_5917);
xnor U7025 (N_7025,N_6201,N_5606);
and U7026 (N_7026,N_6388,N_5843);
xnor U7027 (N_7027,N_5767,N_5702);
and U7028 (N_7028,N_5754,N_5845);
and U7029 (N_7029,N_5682,N_5977);
nand U7030 (N_7030,N_5882,N_6280);
and U7031 (N_7031,N_6381,N_5773);
and U7032 (N_7032,N_6316,N_6309);
or U7033 (N_7033,N_5722,N_5721);
or U7034 (N_7034,N_6042,N_5718);
nand U7035 (N_7035,N_5734,N_5788);
and U7036 (N_7036,N_6298,N_6304);
or U7037 (N_7037,N_5757,N_6085);
nor U7038 (N_7038,N_5977,N_6161);
xnor U7039 (N_7039,N_5860,N_5742);
nand U7040 (N_7040,N_5759,N_6329);
nor U7041 (N_7041,N_6132,N_5881);
nor U7042 (N_7042,N_6037,N_6354);
and U7043 (N_7043,N_6196,N_6125);
or U7044 (N_7044,N_5727,N_5792);
and U7045 (N_7045,N_5672,N_5684);
and U7046 (N_7046,N_5852,N_5923);
xnor U7047 (N_7047,N_5882,N_6208);
or U7048 (N_7048,N_5999,N_6362);
nand U7049 (N_7049,N_5691,N_6040);
xnor U7050 (N_7050,N_6342,N_6271);
nand U7051 (N_7051,N_6376,N_6388);
nand U7052 (N_7052,N_6097,N_5667);
xor U7053 (N_7053,N_5959,N_6262);
nor U7054 (N_7054,N_6014,N_5870);
and U7055 (N_7055,N_6136,N_6121);
nand U7056 (N_7056,N_5914,N_5943);
xor U7057 (N_7057,N_6117,N_6115);
nand U7058 (N_7058,N_6221,N_5650);
and U7059 (N_7059,N_6397,N_6077);
nand U7060 (N_7060,N_5705,N_6310);
or U7061 (N_7061,N_6276,N_6073);
or U7062 (N_7062,N_5724,N_6043);
or U7063 (N_7063,N_5754,N_6034);
nor U7064 (N_7064,N_5886,N_5982);
and U7065 (N_7065,N_5718,N_5766);
xnor U7066 (N_7066,N_5878,N_5637);
or U7067 (N_7067,N_6300,N_5754);
xor U7068 (N_7068,N_5730,N_6280);
nand U7069 (N_7069,N_6333,N_6249);
nand U7070 (N_7070,N_5995,N_5693);
and U7071 (N_7071,N_5878,N_5785);
nor U7072 (N_7072,N_5911,N_6045);
nand U7073 (N_7073,N_5859,N_5739);
nor U7074 (N_7074,N_6356,N_5733);
nor U7075 (N_7075,N_5839,N_6232);
nand U7076 (N_7076,N_5965,N_6097);
xor U7077 (N_7077,N_5734,N_5783);
nand U7078 (N_7078,N_6193,N_5721);
nor U7079 (N_7079,N_6080,N_6399);
nand U7080 (N_7080,N_6383,N_5853);
xnor U7081 (N_7081,N_5731,N_5928);
or U7082 (N_7082,N_5948,N_5669);
xnor U7083 (N_7083,N_6073,N_6035);
and U7084 (N_7084,N_6085,N_6202);
xnor U7085 (N_7085,N_5903,N_6304);
xor U7086 (N_7086,N_6393,N_5867);
xor U7087 (N_7087,N_5714,N_6100);
or U7088 (N_7088,N_5827,N_6262);
nor U7089 (N_7089,N_6182,N_6000);
nand U7090 (N_7090,N_5966,N_5603);
xor U7091 (N_7091,N_6271,N_5700);
xnor U7092 (N_7092,N_6165,N_5729);
or U7093 (N_7093,N_5692,N_6032);
nand U7094 (N_7094,N_5963,N_5962);
and U7095 (N_7095,N_5602,N_5726);
nand U7096 (N_7096,N_5767,N_6085);
xnor U7097 (N_7097,N_5729,N_6209);
and U7098 (N_7098,N_6392,N_5866);
nand U7099 (N_7099,N_6102,N_6133);
nand U7100 (N_7100,N_6350,N_6155);
xnor U7101 (N_7101,N_6389,N_6187);
xor U7102 (N_7102,N_6287,N_5709);
nand U7103 (N_7103,N_5956,N_6265);
nand U7104 (N_7104,N_5615,N_5906);
or U7105 (N_7105,N_6311,N_5812);
xnor U7106 (N_7106,N_6272,N_5801);
nand U7107 (N_7107,N_5993,N_6222);
and U7108 (N_7108,N_6146,N_5846);
or U7109 (N_7109,N_6391,N_6286);
or U7110 (N_7110,N_6017,N_5975);
nor U7111 (N_7111,N_5915,N_5887);
xnor U7112 (N_7112,N_6053,N_6086);
xor U7113 (N_7113,N_6169,N_5718);
or U7114 (N_7114,N_5896,N_6166);
nand U7115 (N_7115,N_5722,N_5627);
or U7116 (N_7116,N_5705,N_6300);
and U7117 (N_7117,N_6364,N_6200);
nand U7118 (N_7118,N_6308,N_6159);
nor U7119 (N_7119,N_5821,N_6347);
nor U7120 (N_7120,N_6189,N_5668);
or U7121 (N_7121,N_6286,N_5973);
nor U7122 (N_7122,N_6125,N_5931);
or U7123 (N_7123,N_5886,N_5826);
nand U7124 (N_7124,N_5617,N_6382);
xnor U7125 (N_7125,N_5761,N_6133);
or U7126 (N_7126,N_5783,N_6020);
nand U7127 (N_7127,N_5639,N_6024);
or U7128 (N_7128,N_6385,N_6026);
and U7129 (N_7129,N_5980,N_6294);
nand U7130 (N_7130,N_5626,N_5947);
nor U7131 (N_7131,N_6205,N_5736);
xor U7132 (N_7132,N_6133,N_6143);
or U7133 (N_7133,N_5903,N_5987);
xnor U7134 (N_7134,N_5830,N_6163);
or U7135 (N_7135,N_5689,N_6054);
xnor U7136 (N_7136,N_5776,N_6077);
nand U7137 (N_7137,N_6244,N_6090);
or U7138 (N_7138,N_6028,N_5644);
nand U7139 (N_7139,N_5943,N_5878);
xor U7140 (N_7140,N_5749,N_6394);
nor U7141 (N_7141,N_6241,N_5842);
and U7142 (N_7142,N_6016,N_5792);
nor U7143 (N_7143,N_5904,N_5966);
nand U7144 (N_7144,N_6204,N_6385);
nand U7145 (N_7145,N_5774,N_6248);
nand U7146 (N_7146,N_5671,N_5751);
xnor U7147 (N_7147,N_6373,N_5618);
xnor U7148 (N_7148,N_5832,N_5859);
xor U7149 (N_7149,N_6241,N_6137);
nor U7150 (N_7150,N_6205,N_6119);
xor U7151 (N_7151,N_6352,N_6365);
or U7152 (N_7152,N_6233,N_6241);
nand U7153 (N_7153,N_5602,N_6336);
nor U7154 (N_7154,N_5871,N_5969);
nor U7155 (N_7155,N_5725,N_5895);
nand U7156 (N_7156,N_6193,N_5931);
or U7157 (N_7157,N_6359,N_5856);
and U7158 (N_7158,N_6111,N_6108);
nor U7159 (N_7159,N_5624,N_5632);
nand U7160 (N_7160,N_6327,N_6074);
or U7161 (N_7161,N_5698,N_5687);
xor U7162 (N_7162,N_5723,N_6262);
nor U7163 (N_7163,N_5999,N_6354);
or U7164 (N_7164,N_5863,N_6299);
and U7165 (N_7165,N_5766,N_6126);
nor U7166 (N_7166,N_5668,N_6239);
nor U7167 (N_7167,N_5711,N_5799);
xnor U7168 (N_7168,N_5776,N_5825);
xnor U7169 (N_7169,N_6119,N_6174);
nor U7170 (N_7170,N_5738,N_6393);
xnor U7171 (N_7171,N_5959,N_6175);
or U7172 (N_7172,N_5856,N_6029);
and U7173 (N_7173,N_5753,N_5723);
and U7174 (N_7174,N_5633,N_5693);
xnor U7175 (N_7175,N_6298,N_6305);
or U7176 (N_7176,N_5836,N_5937);
nand U7177 (N_7177,N_5667,N_5717);
nor U7178 (N_7178,N_5950,N_5702);
or U7179 (N_7179,N_5691,N_6179);
xnor U7180 (N_7180,N_6120,N_5766);
or U7181 (N_7181,N_6038,N_5830);
nand U7182 (N_7182,N_5974,N_5674);
or U7183 (N_7183,N_6347,N_5832);
or U7184 (N_7184,N_6192,N_6386);
xnor U7185 (N_7185,N_6137,N_6300);
or U7186 (N_7186,N_6007,N_6091);
nor U7187 (N_7187,N_6079,N_6013);
or U7188 (N_7188,N_5747,N_6046);
nor U7189 (N_7189,N_5949,N_5984);
or U7190 (N_7190,N_6097,N_5699);
or U7191 (N_7191,N_6193,N_5949);
and U7192 (N_7192,N_6264,N_5927);
and U7193 (N_7193,N_6335,N_6076);
nand U7194 (N_7194,N_5628,N_6105);
nor U7195 (N_7195,N_5898,N_5974);
and U7196 (N_7196,N_6034,N_6226);
and U7197 (N_7197,N_6255,N_5958);
nor U7198 (N_7198,N_6211,N_5851);
or U7199 (N_7199,N_5997,N_5828);
or U7200 (N_7200,N_7148,N_6524);
and U7201 (N_7201,N_7155,N_7153);
or U7202 (N_7202,N_6584,N_6432);
nand U7203 (N_7203,N_6558,N_6709);
xnor U7204 (N_7204,N_6540,N_6454);
nand U7205 (N_7205,N_6693,N_6724);
and U7206 (N_7206,N_6997,N_6784);
and U7207 (N_7207,N_6975,N_6671);
nor U7208 (N_7208,N_6758,N_6768);
nand U7209 (N_7209,N_7106,N_6409);
or U7210 (N_7210,N_6920,N_6806);
nor U7211 (N_7211,N_7126,N_6469);
or U7212 (N_7212,N_6562,N_7011);
and U7213 (N_7213,N_6501,N_6559);
nand U7214 (N_7214,N_6579,N_6948);
or U7215 (N_7215,N_7117,N_6917);
xor U7216 (N_7216,N_6848,N_7170);
xnor U7217 (N_7217,N_6926,N_7040);
nor U7218 (N_7218,N_6809,N_6872);
and U7219 (N_7219,N_6860,N_7099);
nand U7220 (N_7220,N_6849,N_7116);
and U7221 (N_7221,N_6545,N_6827);
xor U7222 (N_7222,N_6633,N_6852);
or U7223 (N_7223,N_6624,N_6581);
and U7224 (N_7224,N_6834,N_6411);
xnor U7225 (N_7225,N_6744,N_6863);
nor U7226 (N_7226,N_6541,N_6455);
or U7227 (N_7227,N_7154,N_6946);
xor U7228 (N_7228,N_7021,N_6985);
and U7229 (N_7229,N_6685,N_6769);
or U7230 (N_7230,N_6443,N_6611);
xnor U7231 (N_7231,N_6811,N_7094);
nor U7232 (N_7232,N_7004,N_7168);
and U7233 (N_7233,N_6560,N_6885);
and U7234 (N_7234,N_6939,N_6518);
and U7235 (N_7235,N_6991,N_7184);
nor U7236 (N_7236,N_6520,N_6798);
and U7237 (N_7237,N_6969,N_6862);
and U7238 (N_7238,N_6514,N_6822);
xnor U7239 (N_7239,N_7091,N_7018);
nor U7240 (N_7240,N_7127,N_6900);
nand U7241 (N_7241,N_6703,N_6406);
or U7242 (N_7242,N_6663,N_6573);
nor U7243 (N_7243,N_6588,N_7017);
xnor U7244 (N_7244,N_6795,N_6548);
or U7245 (N_7245,N_7006,N_6922);
xor U7246 (N_7246,N_6532,N_7079);
xnor U7247 (N_7247,N_6935,N_7022);
or U7248 (N_7248,N_6511,N_7101);
xor U7249 (N_7249,N_6730,N_6925);
xnor U7250 (N_7250,N_6481,N_6478);
or U7251 (N_7251,N_6546,N_6542);
and U7252 (N_7252,N_7077,N_6760);
xnor U7253 (N_7253,N_7063,N_7151);
nor U7254 (N_7254,N_6479,N_6437);
nor U7255 (N_7255,N_6682,N_6642);
nor U7256 (N_7256,N_7157,N_6418);
nor U7257 (N_7257,N_6717,N_6456);
and U7258 (N_7258,N_6934,N_6635);
xnor U7259 (N_7259,N_7137,N_6696);
or U7260 (N_7260,N_6981,N_6659);
nor U7261 (N_7261,N_7034,N_6641);
and U7262 (N_7262,N_7193,N_6712);
xor U7263 (N_7263,N_6757,N_7019);
nand U7264 (N_7264,N_6609,N_7035);
and U7265 (N_7265,N_6817,N_7143);
or U7266 (N_7266,N_7149,N_6743);
and U7267 (N_7267,N_6851,N_6847);
nand U7268 (N_7268,N_6502,N_7047);
xor U7269 (N_7269,N_6876,N_6720);
or U7270 (N_7270,N_6999,N_6438);
nand U7271 (N_7271,N_7083,N_6565);
xnor U7272 (N_7272,N_7032,N_6734);
and U7273 (N_7273,N_6686,N_6937);
nand U7274 (N_7274,N_7142,N_7014);
and U7275 (N_7275,N_6930,N_6854);
nand U7276 (N_7276,N_7183,N_6960);
nand U7277 (N_7277,N_6603,N_6627);
xor U7278 (N_7278,N_7158,N_6904);
and U7279 (N_7279,N_6688,N_6442);
nand U7280 (N_7280,N_6676,N_6736);
and U7281 (N_7281,N_7062,N_6404);
nand U7282 (N_7282,N_6555,N_6445);
nand U7283 (N_7283,N_6733,N_6944);
or U7284 (N_7284,N_6429,N_6462);
nand U7285 (N_7285,N_7080,N_6419);
or U7286 (N_7286,N_6585,N_6756);
nand U7287 (N_7287,N_6907,N_6583);
or U7288 (N_7288,N_6779,N_7177);
and U7289 (N_7289,N_6964,N_6905);
or U7290 (N_7290,N_6766,N_6747);
nand U7291 (N_7291,N_7135,N_6950);
xnor U7292 (N_7292,N_6484,N_6488);
xor U7293 (N_7293,N_7160,N_6807);
xor U7294 (N_7294,N_7164,N_6689);
or U7295 (N_7295,N_7046,N_6668);
xnor U7296 (N_7296,N_6699,N_6533);
xnor U7297 (N_7297,N_6631,N_6804);
or U7298 (N_7298,N_6504,N_6461);
nand U7299 (N_7299,N_6485,N_6874);
xor U7300 (N_7300,N_6896,N_7039);
nand U7301 (N_7301,N_6979,N_6423);
nand U7302 (N_7302,N_6613,N_6503);
xor U7303 (N_7303,N_6649,N_6938);
nor U7304 (N_7304,N_6459,N_6973);
and U7305 (N_7305,N_6739,N_6866);
or U7306 (N_7306,N_6994,N_7003);
xnor U7307 (N_7307,N_7195,N_6868);
nand U7308 (N_7308,N_6653,N_6738);
nor U7309 (N_7309,N_7111,N_6797);
nand U7310 (N_7310,N_6430,N_6634);
nand U7311 (N_7311,N_6489,N_6498);
and U7312 (N_7312,N_7027,N_6951);
nand U7313 (N_7313,N_6775,N_6529);
xnor U7314 (N_7314,N_7144,N_6829);
or U7315 (N_7315,N_6526,N_6652);
and U7316 (N_7316,N_6707,N_6728);
and U7317 (N_7317,N_6710,N_6761);
nand U7318 (N_7318,N_6704,N_6513);
nor U7319 (N_7319,N_6679,N_6838);
nor U7320 (N_7320,N_6616,N_6487);
and U7321 (N_7321,N_6771,N_7178);
nor U7322 (N_7322,N_6790,N_7048);
nand U7323 (N_7323,N_7108,N_7036);
nor U7324 (N_7324,N_7059,N_6803);
nor U7325 (N_7325,N_7124,N_6557);
xor U7326 (N_7326,N_7199,N_6458);
nor U7327 (N_7327,N_7030,N_6449);
and U7328 (N_7328,N_7086,N_7081);
and U7329 (N_7329,N_6493,N_6496);
and U7330 (N_7330,N_6492,N_6844);
nor U7331 (N_7331,N_6692,N_6697);
or U7332 (N_7332,N_6910,N_6523);
and U7333 (N_7333,N_6891,N_6698);
and U7334 (N_7334,N_7029,N_6621);
xnor U7335 (N_7335,N_6898,N_7150);
nor U7336 (N_7336,N_7197,N_6549);
nor U7337 (N_7337,N_6638,N_7185);
or U7338 (N_7338,N_6989,N_6466);
or U7339 (N_7339,N_6660,N_6767);
and U7340 (N_7340,N_7031,N_7087);
or U7341 (N_7341,N_6867,N_6737);
and U7342 (N_7342,N_6924,N_6517);
nand U7343 (N_7343,N_7069,N_6408);
and U7344 (N_7344,N_6619,N_7146);
nor U7345 (N_7345,N_6463,N_6644);
and U7346 (N_7346,N_6879,N_7102);
and U7347 (N_7347,N_6987,N_6793);
xor U7348 (N_7348,N_6967,N_6791);
nand U7349 (N_7349,N_6716,N_6982);
nand U7350 (N_7350,N_6491,N_6632);
nand U7351 (N_7351,N_6672,N_7058);
or U7352 (N_7352,N_6833,N_6869);
xor U7353 (N_7353,N_6467,N_6499);
or U7354 (N_7354,N_6614,N_6519);
nor U7355 (N_7355,N_6836,N_6690);
and U7356 (N_7356,N_6691,N_6949);
or U7357 (N_7357,N_6988,N_6719);
or U7358 (N_7358,N_6932,N_6958);
and U7359 (N_7359,N_6593,N_6572);
or U7360 (N_7360,N_6530,N_7136);
and U7361 (N_7361,N_6886,N_6539);
xnor U7362 (N_7362,N_6482,N_6727);
xor U7363 (N_7363,N_6506,N_6465);
nand U7364 (N_7364,N_6407,N_6528);
and U7365 (N_7365,N_6552,N_6568);
nor U7366 (N_7366,N_6706,N_6911);
and U7367 (N_7367,N_7115,N_6646);
xor U7368 (N_7368,N_6475,N_7033);
and U7369 (N_7369,N_7156,N_6450);
and U7370 (N_7370,N_6596,N_7088);
and U7371 (N_7371,N_6825,N_6505);
and U7372 (N_7372,N_6471,N_6865);
nand U7373 (N_7373,N_6878,N_6516);
and U7374 (N_7374,N_6620,N_6550);
or U7375 (N_7375,N_6674,N_7139);
nand U7376 (N_7376,N_6521,N_7013);
nor U7377 (N_7377,N_6440,N_6801);
xnor U7378 (N_7378,N_7041,N_6909);
and U7379 (N_7379,N_6500,N_7190);
nor U7380 (N_7380,N_7191,N_6575);
nand U7381 (N_7381,N_7009,N_6428);
xnor U7382 (N_7382,N_6476,N_6592);
xor U7383 (N_7383,N_6590,N_6561);
nand U7384 (N_7384,N_6933,N_7052);
and U7385 (N_7385,N_6538,N_7050);
and U7386 (N_7386,N_7140,N_6965);
xor U7387 (N_7387,N_6815,N_6906);
nand U7388 (N_7388,N_6895,N_6840);
nor U7389 (N_7389,N_6759,N_6998);
xnor U7390 (N_7390,N_6892,N_7131);
and U7391 (N_7391,N_6665,N_6402);
nor U7392 (N_7392,N_6883,N_7105);
or U7393 (N_7393,N_6776,N_6884);
nor U7394 (N_7394,N_6955,N_6695);
nand U7395 (N_7395,N_6457,N_7180);
or U7396 (N_7396,N_7075,N_6800);
xor U7397 (N_7397,N_6972,N_6711);
nor U7398 (N_7398,N_7132,N_7056);
nand U7399 (N_7399,N_6623,N_6574);
xnor U7400 (N_7400,N_6810,N_6721);
or U7401 (N_7401,N_6754,N_6952);
or U7402 (N_7402,N_6570,N_7016);
xor U7403 (N_7403,N_6812,N_6400);
and U7404 (N_7404,N_7096,N_6687);
and U7405 (N_7405,N_6431,N_6522);
nand U7406 (N_7406,N_7119,N_6483);
nor U7407 (N_7407,N_6694,N_6954);
or U7408 (N_7408,N_7104,N_6571);
or U7409 (N_7409,N_7020,N_6460);
xnor U7410 (N_7410,N_6882,N_7114);
and U7411 (N_7411,N_6567,N_6433);
xor U7412 (N_7412,N_6486,N_6439);
and U7413 (N_7413,N_7000,N_7130);
nand U7414 (N_7414,N_6681,N_6877);
nor U7415 (N_7415,N_6813,N_6855);
and U7416 (N_7416,N_6763,N_6890);
and U7417 (N_7417,N_6477,N_7179);
nor U7418 (N_7418,N_6628,N_6857);
xor U7419 (N_7419,N_6893,N_6875);
nor U7420 (N_7420,N_7122,N_6831);
and U7421 (N_7421,N_6405,N_7053);
xnor U7422 (N_7422,N_6770,N_6658);
nand U7423 (N_7423,N_6551,N_7188);
nand U7424 (N_7424,N_7161,N_6637);
or U7425 (N_7425,N_6787,N_6984);
and U7426 (N_7426,N_6864,N_7076);
and U7427 (N_7427,N_6780,N_7008);
nand U7428 (N_7428,N_6957,N_7044);
nand U7429 (N_7429,N_6897,N_6669);
nor U7430 (N_7430,N_6713,N_6604);
nand U7431 (N_7431,N_6923,N_7182);
nor U7432 (N_7432,N_7068,N_7074);
and U7433 (N_7433,N_6577,N_6814);
nor U7434 (N_7434,N_7060,N_6683);
nor U7435 (N_7435,N_6888,N_6605);
and U7436 (N_7436,N_7189,N_7107);
and U7437 (N_7437,N_7045,N_6928);
xor U7438 (N_7438,N_6918,N_6781);
nand U7439 (N_7439,N_6902,N_6731);
and U7440 (N_7440,N_6525,N_6701);
nor U7441 (N_7441,N_6643,N_6931);
and U7442 (N_7442,N_6764,N_6835);
or U7443 (N_7443,N_7162,N_6718);
or U7444 (N_7444,N_6678,N_6468);
nor U7445 (N_7445,N_6816,N_6601);
nand U7446 (N_7446,N_7051,N_6448);
or U7447 (N_7447,N_6566,N_7054);
nor U7448 (N_7448,N_6470,N_6941);
or U7449 (N_7449,N_6903,N_6853);
or U7450 (N_7450,N_7196,N_7023);
nor U7451 (N_7451,N_6753,N_6598);
and U7452 (N_7452,N_6639,N_6434);
or U7453 (N_7453,N_6410,N_6921);
xnor U7454 (N_7454,N_6554,N_6626);
xor U7455 (N_7455,N_6742,N_6416);
nand U7456 (N_7456,N_6451,N_6799);
or U7457 (N_7457,N_6708,N_7159);
xor U7458 (N_7458,N_6595,N_7078);
xor U7459 (N_7459,N_6996,N_6427);
nand U7460 (N_7460,N_6661,N_6435);
nand U7461 (N_7461,N_6894,N_7198);
or U7462 (N_7462,N_6714,N_6655);
and U7463 (N_7463,N_6531,N_6610);
nor U7464 (N_7464,N_7026,N_6544);
nand U7465 (N_7465,N_7194,N_7007);
and U7466 (N_7466,N_7172,N_6576);
nand U7467 (N_7467,N_6977,N_6426);
nand U7468 (N_7468,N_7103,N_7070);
nand U7469 (N_7469,N_6929,N_7145);
xor U7470 (N_7470,N_6832,N_6782);
or U7471 (N_7471,N_7098,N_6677);
xor U7472 (N_7472,N_6796,N_6914);
and U7473 (N_7473,N_7002,N_6789);
nand U7474 (N_7474,N_6881,N_6828);
nand U7475 (N_7475,N_6490,N_6830);
nand U7476 (N_7476,N_6846,N_6618);
nand U7477 (N_7477,N_6778,N_7133);
nand U7478 (N_7478,N_6802,N_6412);
nor U7479 (N_7479,N_6995,N_6675);
nor U7480 (N_7480,N_6657,N_6647);
nor U7481 (N_7481,N_7028,N_7134);
nor U7482 (N_7482,N_6786,N_6953);
and U7483 (N_7483,N_7097,N_6648);
and U7484 (N_7484,N_6684,N_6729);
and U7485 (N_7485,N_6421,N_7128);
xor U7486 (N_7486,N_6986,N_7173);
nand U7487 (N_7487,N_6980,N_7055);
nor U7488 (N_7488,N_6794,N_6992);
or U7489 (N_7489,N_7092,N_6725);
nor U7490 (N_7490,N_6494,N_6473);
or U7491 (N_7491,N_6597,N_6602);
or U7492 (N_7492,N_7042,N_6990);
or U7493 (N_7493,N_6956,N_6667);
nand U7494 (N_7494,N_6755,N_6700);
or U7495 (N_7495,N_7084,N_7169);
or U7496 (N_7496,N_6564,N_6553);
nand U7497 (N_7497,N_6976,N_6630);
xor U7498 (N_7498,N_7176,N_6788);
xnor U7499 (N_7499,N_6819,N_7066);
xor U7500 (N_7500,N_6818,N_6765);
nand U7501 (N_7501,N_6722,N_7024);
and U7502 (N_7502,N_6945,N_6664);
nand U7503 (N_7503,N_6959,N_6599);
nor U7504 (N_7504,N_7090,N_6656);
and U7505 (N_7505,N_6413,N_6841);
and U7506 (N_7506,N_6741,N_6971);
nor U7507 (N_7507,N_6792,N_6578);
xnor U7508 (N_7508,N_6705,N_6978);
nand U7509 (N_7509,N_7001,N_6495);
or U7510 (N_7510,N_6420,N_6968);
xor U7511 (N_7511,N_7089,N_7174);
xnor U7512 (N_7512,N_6453,N_6947);
and U7513 (N_7513,N_6591,N_6940);
and U7514 (N_7514,N_6850,N_7167);
or U7515 (N_7515,N_6774,N_6510);
nor U7516 (N_7516,N_7147,N_6962);
xor U7517 (N_7517,N_7166,N_6762);
xnor U7518 (N_7518,N_6750,N_7005);
xnor U7519 (N_7519,N_6915,N_7123);
or U7520 (N_7520,N_6858,N_6908);
nor U7521 (N_7521,N_6856,N_6826);
xor U7522 (N_7522,N_6607,N_6887);
nor U7523 (N_7523,N_7112,N_6414);
and U7524 (N_7524,N_7165,N_6805);
or U7525 (N_7525,N_6622,N_6569);
or U7526 (N_7526,N_6670,N_6422);
and U7527 (N_7527,N_7110,N_6606);
and U7528 (N_7528,N_6446,N_6843);
nor U7529 (N_7529,N_6543,N_6740);
nand U7530 (N_7530,N_6970,N_6654);
and U7531 (N_7531,N_6563,N_7118);
xor U7532 (N_7532,N_6726,N_6600);
nor U7533 (N_7533,N_7057,N_7181);
and U7534 (N_7534,N_7093,N_6645);
xor U7535 (N_7535,N_6993,N_6745);
nor U7536 (N_7536,N_6447,N_6751);
nand U7537 (N_7537,N_6919,N_6842);
xor U7538 (N_7538,N_7043,N_6424);
and U7539 (N_7539,N_6901,N_6415);
nor U7540 (N_7540,N_6650,N_6820);
nand U7541 (N_7541,N_6629,N_6871);
and U7542 (N_7542,N_6587,N_7071);
or U7543 (N_7543,N_7187,N_7175);
xnor U7544 (N_7544,N_6837,N_7186);
nand U7545 (N_7545,N_6732,N_7163);
and U7546 (N_7546,N_6873,N_6748);
and U7547 (N_7547,N_6723,N_6536);
and U7548 (N_7548,N_6527,N_6983);
and U7549 (N_7549,N_6534,N_6640);
nor U7550 (N_7550,N_6912,N_6961);
and U7551 (N_7551,N_6425,N_7085);
or U7552 (N_7552,N_7138,N_7061);
or U7553 (N_7553,N_6783,N_7082);
nor U7554 (N_7554,N_6662,N_6615);
or U7555 (N_7555,N_7025,N_7141);
nand U7556 (N_7556,N_6735,N_6936);
nor U7557 (N_7557,N_6974,N_6889);
or U7558 (N_7558,N_6556,N_6480);
nand U7559 (N_7559,N_6537,N_7012);
xor U7560 (N_7560,N_7192,N_7120);
or U7561 (N_7561,N_6474,N_6617);
or U7562 (N_7562,N_7129,N_6966);
or U7563 (N_7563,N_7121,N_6870);
xor U7564 (N_7564,N_6497,N_6547);
or U7565 (N_7565,N_7072,N_6472);
or U7566 (N_7566,N_6702,N_6927);
or U7567 (N_7567,N_6535,N_6943);
nor U7568 (N_7568,N_6452,N_7109);
xor U7569 (N_7569,N_6899,N_6464);
or U7570 (N_7570,N_6746,N_7049);
xnor U7571 (N_7571,N_6625,N_6589);
or U7572 (N_7572,N_6821,N_6507);
xnor U7573 (N_7573,N_7010,N_6444);
and U7574 (N_7574,N_7067,N_7073);
nand U7575 (N_7575,N_6608,N_7100);
nor U7576 (N_7576,N_6861,N_6824);
or U7577 (N_7577,N_6773,N_6403);
and U7578 (N_7578,N_6749,N_6594);
and U7579 (N_7579,N_6586,N_6680);
or U7580 (N_7580,N_6636,N_7038);
xnor U7581 (N_7581,N_6777,N_6916);
and U7582 (N_7582,N_6823,N_7125);
and U7583 (N_7583,N_6436,N_6963);
nand U7584 (N_7584,N_6512,N_6839);
or U7585 (N_7585,N_7171,N_7015);
nand U7586 (N_7586,N_6508,N_6651);
xor U7587 (N_7587,N_7152,N_7113);
nor U7588 (N_7588,N_6808,N_6441);
xnor U7589 (N_7589,N_6715,N_6913);
xor U7590 (N_7590,N_7065,N_6401);
nor U7591 (N_7591,N_6509,N_6515);
and U7592 (N_7592,N_6942,N_6785);
nand U7593 (N_7593,N_6859,N_7064);
xnor U7594 (N_7594,N_7037,N_6417);
or U7595 (N_7595,N_6752,N_6612);
nand U7596 (N_7596,N_7095,N_6580);
nand U7597 (N_7597,N_6880,N_6666);
nor U7598 (N_7598,N_6582,N_6772);
nor U7599 (N_7599,N_6845,N_6673);
nor U7600 (N_7600,N_6480,N_6804);
xnor U7601 (N_7601,N_6640,N_7005);
or U7602 (N_7602,N_7189,N_6998);
xnor U7603 (N_7603,N_7129,N_6686);
xor U7604 (N_7604,N_6999,N_7048);
nand U7605 (N_7605,N_6992,N_6600);
xnor U7606 (N_7606,N_6920,N_6558);
nor U7607 (N_7607,N_7079,N_7196);
and U7608 (N_7608,N_6652,N_6413);
nor U7609 (N_7609,N_6818,N_6882);
xnor U7610 (N_7610,N_6790,N_6823);
nand U7611 (N_7611,N_6957,N_7157);
nand U7612 (N_7612,N_6502,N_6469);
nand U7613 (N_7613,N_6743,N_7019);
nand U7614 (N_7614,N_6724,N_6761);
nor U7615 (N_7615,N_6683,N_6712);
and U7616 (N_7616,N_6937,N_6903);
and U7617 (N_7617,N_7157,N_6490);
nand U7618 (N_7618,N_6840,N_7015);
or U7619 (N_7619,N_6784,N_7185);
or U7620 (N_7620,N_6753,N_6475);
nor U7621 (N_7621,N_6561,N_6733);
nor U7622 (N_7622,N_6408,N_6603);
nand U7623 (N_7623,N_6787,N_6609);
and U7624 (N_7624,N_7090,N_6778);
nor U7625 (N_7625,N_6998,N_6940);
nor U7626 (N_7626,N_6775,N_6463);
nand U7627 (N_7627,N_6471,N_7084);
xnor U7628 (N_7628,N_7108,N_6599);
or U7629 (N_7629,N_6481,N_6558);
nand U7630 (N_7630,N_7168,N_6973);
nor U7631 (N_7631,N_6863,N_7115);
nand U7632 (N_7632,N_7045,N_6907);
xnor U7633 (N_7633,N_6581,N_6520);
nor U7634 (N_7634,N_6634,N_6560);
xor U7635 (N_7635,N_6910,N_7183);
and U7636 (N_7636,N_6983,N_6714);
nor U7637 (N_7637,N_6596,N_7061);
or U7638 (N_7638,N_6532,N_7035);
xor U7639 (N_7639,N_6962,N_7012);
nand U7640 (N_7640,N_7049,N_7034);
xor U7641 (N_7641,N_6918,N_6788);
nand U7642 (N_7642,N_7124,N_6427);
and U7643 (N_7643,N_6531,N_6991);
or U7644 (N_7644,N_7199,N_6767);
xnor U7645 (N_7645,N_7113,N_6838);
and U7646 (N_7646,N_7101,N_6795);
xnor U7647 (N_7647,N_6832,N_6727);
nand U7648 (N_7648,N_6482,N_7047);
or U7649 (N_7649,N_6643,N_7035);
and U7650 (N_7650,N_7016,N_6767);
nor U7651 (N_7651,N_7123,N_7023);
or U7652 (N_7652,N_6928,N_6483);
and U7653 (N_7653,N_7030,N_6781);
xor U7654 (N_7654,N_6973,N_6692);
nand U7655 (N_7655,N_6725,N_7157);
xor U7656 (N_7656,N_6756,N_7078);
nand U7657 (N_7657,N_6808,N_6525);
and U7658 (N_7658,N_6468,N_7128);
and U7659 (N_7659,N_6668,N_6804);
nor U7660 (N_7660,N_6550,N_6580);
nor U7661 (N_7661,N_6872,N_6914);
nand U7662 (N_7662,N_6761,N_7091);
nor U7663 (N_7663,N_6654,N_6440);
nand U7664 (N_7664,N_7199,N_6555);
nand U7665 (N_7665,N_6750,N_6881);
xnor U7666 (N_7666,N_7127,N_6612);
and U7667 (N_7667,N_7103,N_7025);
nand U7668 (N_7668,N_6750,N_7018);
and U7669 (N_7669,N_6756,N_6939);
and U7670 (N_7670,N_6828,N_6765);
or U7671 (N_7671,N_6575,N_6942);
and U7672 (N_7672,N_6596,N_6820);
nand U7673 (N_7673,N_6869,N_6876);
and U7674 (N_7674,N_6478,N_7024);
or U7675 (N_7675,N_7162,N_7026);
or U7676 (N_7676,N_7045,N_6649);
nor U7677 (N_7677,N_6426,N_7068);
or U7678 (N_7678,N_6800,N_6578);
nor U7679 (N_7679,N_6625,N_6774);
xor U7680 (N_7680,N_7139,N_6624);
or U7681 (N_7681,N_6984,N_6533);
nor U7682 (N_7682,N_7097,N_6460);
xnor U7683 (N_7683,N_7146,N_7143);
nand U7684 (N_7684,N_6846,N_7092);
nor U7685 (N_7685,N_6939,N_7192);
or U7686 (N_7686,N_6651,N_6901);
and U7687 (N_7687,N_7069,N_7107);
nor U7688 (N_7688,N_7061,N_6548);
and U7689 (N_7689,N_6993,N_6553);
or U7690 (N_7690,N_7116,N_6735);
nand U7691 (N_7691,N_6577,N_6678);
or U7692 (N_7692,N_7180,N_6431);
xnor U7693 (N_7693,N_7162,N_6946);
and U7694 (N_7694,N_6986,N_6971);
nand U7695 (N_7695,N_6843,N_6951);
or U7696 (N_7696,N_6874,N_6982);
or U7697 (N_7697,N_7117,N_6593);
nor U7698 (N_7698,N_6821,N_6800);
nor U7699 (N_7699,N_6797,N_6962);
nor U7700 (N_7700,N_6989,N_7094);
nor U7701 (N_7701,N_6596,N_6987);
xor U7702 (N_7702,N_6536,N_7073);
and U7703 (N_7703,N_6553,N_7100);
xor U7704 (N_7704,N_6576,N_6734);
nand U7705 (N_7705,N_6850,N_6872);
xor U7706 (N_7706,N_7166,N_6628);
nand U7707 (N_7707,N_6533,N_6833);
nand U7708 (N_7708,N_6770,N_6682);
nand U7709 (N_7709,N_6467,N_6801);
and U7710 (N_7710,N_6736,N_6578);
xor U7711 (N_7711,N_7185,N_6905);
and U7712 (N_7712,N_6497,N_6579);
nand U7713 (N_7713,N_6981,N_7028);
nor U7714 (N_7714,N_6802,N_6581);
nand U7715 (N_7715,N_6979,N_6882);
nor U7716 (N_7716,N_6597,N_6949);
xnor U7717 (N_7717,N_6462,N_6821);
nor U7718 (N_7718,N_6483,N_6546);
or U7719 (N_7719,N_6959,N_6501);
nand U7720 (N_7720,N_6427,N_7094);
nor U7721 (N_7721,N_6976,N_7195);
nor U7722 (N_7722,N_6742,N_6484);
xnor U7723 (N_7723,N_7132,N_6981);
and U7724 (N_7724,N_6648,N_6737);
nor U7725 (N_7725,N_7085,N_7031);
xor U7726 (N_7726,N_6949,N_6630);
nor U7727 (N_7727,N_7022,N_6995);
nor U7728 (N_7728,N_6918,N_6758);
nand U7729 (N_7729,N_6446,N_6594);
and U7730 (N_7730,N_6438,N_7141);
or U7731 (N_7731,N_6814,N_6816);
nor U7732 (N_7732,N_7070,N_6942);
and U7733 (N_7733,N_6690,N_7061);
nor U7734 (N_7734,N_6420,N_7080);
xor U7735 (N_7735,N_7108,N_6509);
or U7736 (N_7736,N_6474,N_6418);
or U7737 (N_7737,N_7007,N_6851);
nand U7738 (N_7738,N_6652,N_6651);
and U7739 (N_7739,N_7029,N_6807);
xor U7740 (N_7740,N_7002,N_6913);
or U7741 (N_7741,N_6621,N_6847);
xor U7742 (N_7742,N_6947,N_6464);
nor U7743 (N_7743,N_6572,N_7154);
and U7744 (N_7744,N_6898,N_6735);
or U7745 (N_7745,N_6535,N_6550);
nand U7746 (N_7746,N_6472,N_7004);
nand U7747 (N_7747,N_6571,N_6567);
nor U7748 (N_7748,N_6705,N_6424);
xor U7749 (N_7749,N_7068,N_6714);
and U7750 (N_7750,N_7125,N_6518);
nand U7751 (N_7751,N_6611,N_6847);
nor U7752 (N_7752,N_6603,N_6684);
xnor U7753 (N_7753,N_6608,N_6636);
xor U7754 (N_7754,N_6475,N_6975);
xnor U7755 (N_7755,N_6461,N_6683);
nand U7756 (N_7756,N_6992,N_6589);
nor U7757 (N_7757,N_6904,N_6646);
xor U7758 (N_7758,N_6656,N_7140);
xor U7759 (N_7759,N_6487,N_6708);
nand U7760 (N_7760,N_6697,N_6891);
nand U7761 (N_7761,N_6823,N_6630);
or U7762 (N_7762,N_7159,N_6554);
or U7763 (N_7763,N_6505,N_6405);
or U7764 (N_7764,N_7056,N_6503);
and U7765 (N_7765,N_6934,N_6918);
or U7766 (N_7766,N_7076,N_6786);
nand U7767 (N_7767,N_6686,N_6893);
xnor U7768 (N_7768,N_6481,N_7086);
xnor U7769 (N_7769,N_7010,N_6794);
nand U7770 (N_7770,N_6973,N_6775);
xor U7771 (N_7771,N_6568,N_6515);
and U7772 (N_7772,N_6826,N_6818);
and U7773 (N_7773,N_6402,N_6692);
xor U7774 (N_7774,N_6463,N_6755);
nand U7775 (N_7775,N_7199,N_6889);
xnor U7776 (N_7776,N_6705,N_6847);
xor U7777 (N_7777,N_6456,N_6757);
nor U7778 (N_7778,N_6453,N_6486);
or U7779 (N_7779,N_6717,N_6488);
and U7780 (N_7780,N_6474,N_6708);
and U7781 (N_7781,N_6493,N_6902);
or U7782 (N_7782,N_7004,N_6988);
nor U7783 (N_7783,N_6991,N_7190);
xnor U7784 (N_7784,N_6766,N_6869);
or U7785 (N_7785,N_6939,N_6859);
xnor U7786 (N_7786,N_6503,N_6514);
and U7787 (N_7787,N_7100,N_6657);
nor U7788 (N_7788,N_6936,N_6673);
xor U7789 (N_7789,N_6989,N_7132);
xor U7790 (N_7790,N_7168,N_6405);
xor U7791 (N_7791,N_7060,N_7055);
and U7792 (N_7792,N_7167,N_6948);
nor U7793 (N_7793,N_7175,N_7000);
or U7794 (N_7794,N_6825,N_7145);
or U7795 (N_7795,N_6672,N_6431);
nand U7796 (N_7796,N_7058,N_6612);
nand U7797 (N_7797,N_6824,N_6490);
xnor U7798 (N_7798,N_6421,N_6492);
and U7799 (N_7799,N_7188,N_6649);
nand U7800 (N_7800,N_6490,N_6794);
nand U7801 (N_7801,N_6559,N_6779);
nand U7802 (N_7802,N_6502,N_6896);
nor U7803 (N_7803,N_6723,N_6409);
and U7804 (N_7804,N_7016,N_6735);
nor U7805 (N_7805,N_6915,N_6985);
nand U7806 (N_7806,N_6677,N_6645);
xor U7807 (N_7807,N_7089,N_7047);
and U7808 (N_7808,N_7106,N_6524);
and U7809 (N_7809,N_6513,N_6543);
xor U7810 (N_7810,N_6552,N_6737);
xnor U7811 (N_7811,N_6508,N_6978);
or U7812 (N_7812,N_6741,N_6501);
or U7813 (N_7813,N_6942,N_6513);
xnor U7814 (N_7814,N_6625,N_6924);
and U7815 (N_7815,N_6704,N_7199);
nand U7816 (N_7816,N_7173,N_6965);
or U7817 (N_7817,N_6783,N_6877);
xnor U7818 (N_7818,N_6866,N_6558);
or U7819 (N_7819,N_6439,N_7168);
or U7820 (N_7820,N_6936,N_6631);
nand U7821 (N_7821,N_6507,N_7031);
and U7822 (N_7822,N_6684,N_7048);
nand U7823 (N_7823,N_7032,N_6935);
nor U7824 (N_7824,N_7130,N_6619);
or U7825 (N_7825,N_6847,N_6685);
nor U7826 (N_7826,N_6454,N_6479);
or U7827 (N_7827,N_6711,N_6569);
nor U7828 (N_7828,N_7073,N_6522);
and U7829 (N_7829,N_7046,N_7078);
nand U7830 (N_7830,N_6645,N_7025);
nand U7831 (N_7831,N_7067,N_6643);
or U7832 (N_7832,N_6451,N_6561);
or U7833 (N_7833,N_6729,N_6799);
and U7834 (N_7834,N_6419,N_6607);
nor U7835 (N_7835,N_6589,N_6580);
nand U7836 (N_7836,N_6500,N_6768);
xnor U7837 (N_7837,N_6909,N_7002);
nor U7838 (N_7838,N_6777,N_7111);
and U7839 (N_7839,N_6472,N_6450);
or U7840 (N_7840,N_6946,N_6833);
or U7841 (N_7841,N_6602,N_6770);
nor U7842 (N_7842,N_6869,N_6564);
nor U7843 (N_7843,N_6738,N_6434);
nand U7844 (N_7844,N_6681,N_7195);
nor U7845 (N_7845,N_6461,N_6401);
nand U7846 (N_7846,N_6836,N_6986);
nand U7847 (N_7847,N_7126,N_6624);
xnor U7848 (N_7848,N_6615,N_7056);
nand U7849 (N_7849,N_6738,N_6580);
and U7850 (N_7850,N_6798,N_6855);
or U7851 (N_7851,N_6599,N_6595);
and U7852 (N_7852,N_6402,N_6588);
xor U7853 (N_7853,N_7053,N_6536);
xnor U7854 (N_7854,N_6951,N_6936);
xnor U7855 (N_7855,N_6828,N_6976);
nor U7856 (N_7856,N_6881,N_6494);
or U7857 (N_7857,N_6956,N_6516);
nand U7858 (N_7858,N_6956,N_6419);
and U7859 (N_7859,N_7152,N_6478);
or U7860 (N_7860,N_7050,N_6827);
and U7861 (N_7861,N_6939,N_6748);
nor U7862 (N_7862,N_6884,N_6852);
nand U7863 (N_7863,N_6614,N_6960);
nand U7864 (N_7864,N_6764,N_6552);
nor U7865 (N_7865,N_6415,N_6771);
or U7866 (N_7866,N_6710,N_7076);
xor U7867 (N_7867,N_6871,N_6963);
or U7868 (N_7868,N_7127,N_6971);
nand U7869 (N_7869,N_6440,N_6934);
and U7870 (N_7870,N_6642,N_6840);
xor U7871 (N_7871,N_7063,N_7124);
or U7872 (N_7872,N_6625,N_6437);
and U7873 (N_7873,N_6638,N_6409);
and U7874 (N_7874,N_6722,N_6516);
and U7875 (N_7875,N_7076,N_6610);
or U7876 (N_7876,N_6420,N_6829);
and U7877 (N_7877,N_7162,N_7167);
and U7878 (N_7878,N_6902,N_6727);
nor U7879 (N_7879,N_7172,N_6994);
xor U7880 (N_7880,N_6528,N_7060);
nand U7881 (N_7881,N_6424,N_6951);
nor U7882 (N_7882,N_6927,N_6972);
nor U7883 (N_7883,N_7091,N_6921);
nor U7884 (N_7884,N_6494,N_6822);
nor U7885 (N_7885,N_6719,N_6779);
xnor U7886 (N_7886,N_6795,N_6553);
nor U7887 (N_7887,N_7112,N_6683);
xnor U7888 (N_7888,N_6690,N_6937);
or U7889 (N_7889,N_6415,N_7063);
nor U7890 (N_7890,N_6774,N_6986);
nand U7891 (N_7891,N_6907,N_6668);
nand U7892 (N_7892,N_6912,N_7001);
and U7893 (N_7893,N_6893,N_6630);
nand U7894 (N_7894,N_6811,N_6820);
nor U7895 (N_7895,N_6989,N_6429);
and U7896 (N_7896,N_6598,N_6476);
nor U7897 (N_7897,N_6613,N_6787);
or U7898 (N_7898,N_6869,N_6964);
nand U7899 (N_7899,N_6605,N_6598);
and U7900 (N_7900,N_6860,N_6433);
xor U7901 (N_7901,N_6903,N_6884);
and U7902 (N_7902,N_6576,N_6658);
xor U7903 (N_7903,N_7079,N_7165);
or U7904 (N_7904,N_6412,N_7066);
xnor U7905 (N_7905,N_6610,N_6482);
xnor U7906 (N_7906,N_6519,N_6997);
xnor U7907 (N_7907,N_6552,N_6545);
or U7908 (N_7908,N_7016,N_6771);
nand U7909 (N_7909,N_6871,N_6668);
and U7910 (N_7910,N_6910,N_6897);
xor U7911 (N_7911,N_7084,N_6793);
nand U7912 (N_7912,N_7042,N_7121);
nand U7913 (N_7913,N_6489,N_6730);
nand U7914 (N_7914,N_6788,N_6541);
xor U7915 (N_7915,N_6926,N_6488);
nor U7916 (N_7916,N_6813,N_6413);
and U7917 (N_7917,N_6482,N_6868);
and U7918 (N_7918,N_6645,N_7097);
nor U7919 (N_7919,N_6911,N_7184);
xor U7920 (N_7920,N_6850,N_7196);
and U7921 (N_7921,N_6521,N_7017);
nand U7922 (N_7922,N_6487,N_6810);
and U7923 (N_7923,N_7115,N_6866);
xnor U7924 (N_7924,N_6856,N_6914);
and U7925 (N_7925,N_6833,N_6836);
and U7926 (N_7926,N_6892,N_6772);
nor U7927 (N_7927,N_6807,N_6497);
and U7928 (N_7928,N_6883,N_6727);
and U7929 (N_7929,N_6443,N_6735);
or U7930 (N_7930,N_7141,N_6785);
xor U7931 (N_7931,N_6815,N_6597);
and U7932 (N_7932,N_7139,N_6651);
or U7933 (N_7933,N_7050,N_6748);
nand U7934 (N_7934,N_7192,N_6971);
xnor U7935 (N_7935,N_6960,N_6406);
or U7936 (N_7936,N_6416,N_6799);
or U7937 (N_7937,N_7099,N_7123);
and U7938 (N_7938,N_6606,N_7153);
xor U7939 (N_7939,N_6656,N_6640);
xnor U7940 (N_7940,N_6735,N_6521);
nor U7941 (N_7941,N_6702,N_6698);
or U7942 (N_7942,N_7072,N_6646);
nor U7943 (N_7943,N_6581,N_6413);
and U7944 (N_7944,N_7079,N_6421);
and U7945 (N_7945,N_6605,N_6478);
xor U7946 (N_7946,N_7098,N_6642);
and U7947 (N_7947,N_7151,N_7134);
xor U7948 (N_7948,N_6871,N_7133);
xor U7949 (N_7949,N_6791,N_6430);
or U7950 (N_7950,N_7151,N_6556);
and U7951 (N_7951,N_6673,N_6568);
nand U7952 (N_7952,N_6430,N_7175);
xor U7953 (N_7953,N_6631,N_6578);
nand U7954 (N_7954,N_6873,N_6779);
nand U7955 (N_7955,N_7143,N_6739);
xnor U7956 (N_7956,N_7053,N_7185);
or U7957 (N_7957,N_7012,N_6469);
nor U7958 (N_7958,N_6842,N_6497);
nor U7959 (N_7959,N_6441,N_6576);
nand U7960 (N_7960,N_6894,N_6542);
nor U7961 (N_7961,N_6992,N_6863);
or U7962 (N_7962,N_6896,N_7109);
nor U7963 (N_7963,N_6490,N_6947);
nor U7964 (N_7964,N_6722,N_6865);
xor U7965 (N_7965,N_7193,N_6521);
xnor U7966 (N_7966,N_6859,N_6564);
nand U7967 (N_7967,N_6643,N_6664);
xnor U7968 (N_7968,N_6565,N_7022);
and U7969 (N_7969,N_6479,N_6953);
and U7970 (N_7970,N_6646,N_6877);
nor U7971 (N_7971,N_6493,N_7091);
nand U7972 (N_7972,N_6475,N_6485);
nor U7973 (N_7973,N_6877,N_6478);
nor U7974 (N_7974,N_6972,N_7019);
or U7975 (N_7975,N_6746,N_7004);
nand U7976 (N_7976,N_6435,N_6772);
or U7977 (N_7977,N_7077,N_6855);
and U7978 (N_7978,N_7198,N_7179);
xnor U7979 (N_7979,N_7171,N_6450);
nor U7980 (N_7980,N_6659,N_7058);
nand U7981 (N_7981,N_6972,N_6622);
and U7982 (N_7982,N_6948,N_6471);
nand U7983 (N_7983,N_7006,N_6917);
xor U7984 (N_7984,N_7108,N_6801);
nand U7985 (N_7985,N_6743,N_6736);
xnor U7986 (N_7986,N_6780,N_6471);
xor U7987 (N_7987,N_6747,N_7000);
or U7988 (N_7988,N_6450,N_7191);
nor U7989 (N_7989,N_7039,N_6630);
nand U7990 (N_7990,N_6968,N_7096);
nand U7991 (N_7991,N_6986,N_6466);
or U7992 (N_7992,N_6810,N_7074);
or U7993 (N_7993,N_6775,N_6672);
xor U7994 (N_7994,N_7190,N_6730);
nand U7995 (N_7995,N_6694,N_6498);
nand U7996 (N_7996,N_6942,N_6899);
nor U7997 (N_7997,N_6787,N_6907);
or U7998 (N_7998,N_6944,N_6415);
or U7999 (N_7999,N_6595,N_7092);
and U8000 (N_8000,N_7359,N_7540);
and U8001 (N_8001,N_7239,N_7543);
and U8002 (N_8002,N_7646,N_7243);
xor U8003 (N_8003,N_7929,N_7744);
or U8004 (N_8004,N_7278,N_7800);
nand U8005 (N_8005,N_7487,N_7375);
or U8006 (N_8006,N_7514,N_7890);
and U8007 (N_8007,N_7609,N_7286);
nand U8008 (N_8008,N_7712,N_7228);
and U8009 (N_8009,N_7205,N_7805);
nor U8010 (N_8010,N_7496,N_7667);
nand U8011 (N_8011,N_7791,N_7902);
or U8012 (N_8012,N_7383,N_7427);
nand U8013 (N_8013,N_7906,N_7768);
nor U8014 (N_8014,N_7925,N_7743);
nand U8015 (N_8015,N_7645,N_7838);
or U8016 (N_8016,N_7616,N_7698);
or U8017 (N_8017,N_7242,N_7716);
and U8018 (N_8018,N_7985,N_7598);
nand U8019 (N_8019,N_7757,N_7466);
or U8020 (N_8020,N_7888,N_7549);
and U8021 (N_8021,N_7425,N_7649);
and U8022 (N_8022,N_7275,N_7879);
and U8023 (N_8023,N_7300,N_7891);
xnor U8024 (N_8024,N_7745,N_7608);
nand U8025 (N_8025,N_7332,N_7656);
and U8026 (N_8026,N_7264,N_7519);
or U8027 (N_8027,N_7816,N_7672);
nand U8028 (N_8028,N_7450,N_7895);
nand U8029 (N_8029,N_7660,N_7749);
xnor U8030 (N_8030,N_7561,N_7433);
nand U8031 (N_8031,N_7710,N_7727);
and U8032 (N_8032,N_7774,N_7430);
xor U8033 (N_8033,N_7643,N_7234);
or U8034 (N_8034,N_7389,N_7620);
nand U8035 (N_8035,N_7532,N_7265);
nand U8036 (N_8036,N_7545,N_7563);
xnor U8037 (N_8037,N_7361,N_7784);
and U8038 (N_8038,N_7859,N_7615);
xnor U8039 (N_8039,N_7373,N_7814);
and U8040 (N_8040,N_7241,N_7623);
nand U8041 (N_8041,N_7521,N_7453);
nand U8042 (N_8042,N_7410,N_7688);
and U8043 (N_8043,N_7639,N_7328);
and U8044 (N_8044,N_7980,N_7982);
nand U8045 (N_8045,N_7460,N_7594);
or U8046 (N_8046,N_7584,N_7969);
or U8047 (N_8047,N_7517,N_7820);
and U8048 (N_8048,N_7674,N_7246);
nand U8049 (N_8049,N_7964,N_7779);
nand U8050 (N_8050,N_7892,N_7484);
nand U8051 (N_8051,N_7409,N_7834);
xor U8052 (N_8052,N_7229,N_7213);
or U8053 (N_8053,N_7642,N_7404);
nor U8054 (N_8054,N_7270,N_7721);
or U8055 (N_8055,N_7928,N_7970);
nor U8056 (N_8056,N_7381,N_7380);
or U8057 (N_8057,N_7459,N_7288);
nor U8058 (N_8058,N_7932,N_7499);
nor U8059 (N_8059,N_7715,N_7552);
xnor U8060 (N_8060,N_7494,N_7343);
xnor U8061 (N_8061,N_7345,N_7454);
xnor U8062 (N_8062,N_7378,N_7678);
nor U8063 (N_8063,N_7669,N_7537);
or U8064 (N_8064,N_7872,N_7578);
nor U8065 (N_8065,N_7334,N_7962);
or U8066 (N_8066,N_7777,N_7931);
nand U8067 (N_8067,N_7344,N_7438);
nor U8068 (N_8068,N_7350,N_7787);
nor U8069 (N_8069,N_7899,N_7764);
and U8070 (N_8070,N_7445,N_7792);
or U8071 (N_8071,N_7861,N_7534);
nor U8072 (N_8072,N_7556,N_7447);
or U8073 (N_8073,N_7628,N_7668);
nand U8074 (N_8074,N_7780,N_7949);
nor U8075 (N_8075,N_7564,N_7988);
xor U8076 (N_8076,N_7354,N_7823);
nor U8077 (N_8077,N_7612,N_7798);
nand U8078 (N_8078,N_7547,N_7652);
and U8079 (N_8079,N_7386,N_7529);
and U8080 (N_8080,N_7326,N_7480);
and U8081 (N_8081,N_7714,N_7883);
and U8082 (N_8082,N_7392,N_7877);
or U8083 (N_8083,N_7281,N_7737);
nand U8084 (N_8084,N_7390,N_7796);
and U8085 (N_8085,N_7233,N_7840);
and U8086 (N_8086,N_7247,N_7367);
and U8087 (N_8087,N_7588,N_7548);
and U8088 (N_8088,N_7587,N_7349);
nor U8089 (N_8089,N_7299,N_7691);
and U8090 (N_8090,N_7323,N_7795);
xor U8091 (N_8091,N_7808,N_7551);
nor U8092 (N_8092,N_7474,N_7401);
or U8093 (N_8093,N_7277,N_7740);
and U8094 (N_8094,N_7766,N_7842);
xor U8095 (N_8095,N_7283,N_7971);
and U8096 (N_8096,N_7396,N_7684);
nand U8097 (N_8097,N_7218,N_7807);
or U8098 (N_8098,N_7919,N_7975);
or U8099 (N_8099,N_7456,N_7348);
and U8100 (N_8100,N_7833,N_7400);
or U8101 (N_8101,N_7408,N_7618);
nand U8102 (N_8102,N_7759,N_7209);
or U8103 (N_8103,N_7613,N_7599);
and U8104 (N_8104,N_7305,N_7789);
and U8105 (N_8105,N_7702,N_7763);
or U8106 (N_8106,N_7403,N_7388);
nor U8107 (N_8107,N_7933,N_7290);
and U8108 (N_8108,N_7946,N_7307);
or U8109 (N_8109,N_7333,N_7670);
nor U8110 (N_8110,N_7836,N_7516);
nand U8111 (N_8111,N_7295,N_7604);
nor U8112 (N_8112,N_7694,N_7706);
xor U8113 (N_8113,N_7990,N_7738);
or U8114 (N_8114,N_7841,N_7907);
xnor U8115 (N_8115,N_7958,N_7417);
xor U8116 (N_8116,N_7767,N_7268);
nand U8117 (N_8117,N_7202,N_7908);
and U8118 (N_8118,N_7631,N_7995);
or U8119 (N_8119,N_7483,N_7731);
nor U8120 (N_8120,N_7724,N_7274);
nor U8121 (N_8121,N_7812,N_7802);
nand U8122 (N_8122,N_7269,N_7225);
nor U8123 (N_8123,N_7822,N_7314);
or U8124 (N_8124,N_7555,N_7446);
xor U8125 (N_8125,N_7370,N_7530);
and U8126 (N_8126,N_7734,N_7799);
nand U8127 (N_8127,N_7753,N_7916);
xor U8128 (N_8128,N_7340,N_7910);
nor U8129 (N_8129,N_7568,N_7231);
nand U8130 (N_8130,N_7465,N_7352);
xnor U8131 (N_8131,N_7260,N_7904);
or U8132 (N_8132,N_7659,N_7539);
nor U8133 (N_8133,N_7697,N_7546);
nand U8134 (N_8134,N_7923,N_7490);
nand U8135 (N_8135,N_7898,N_7263);
nand U8136 (N_8136,N_7806,N_7809);
or U8137 (N_8137,N_7752,N_7583);
xnor U8138 (N_8138,N_7501,N_7203);
and U8139 (N_8139,N_7909,N_7941);
and U8140 (N_8140,N_7502,N_7482);
and U8141 (N_8141,N_7576,N_7322);
or U8142 (N_8142,N_7874,N_7897);
and U8143 (N_8143,N_7266,N_7586);
xnor U8144 (N_8144,N_7720,N_7204);
and U8145 (N_8145,N_7330,N_7479);
or U8146 (N_8146,N_7863,N_7650);
nand U8147 (N_8147,N_7945,N_7605);
xnor U8148 (N_8148,N_7921,N_7607);
and U8149 (N_8149,N_7419,N_7379);
nor U8150 (N_8150,N_7533,N_7794);
and U8151 (N_8151,N_7978,N_7312);
or U8152 (N_8152,N_7819,N_7986);
and U8153 (N_8153,N_7503,N_7315);
nor U8154 (N_8154,N_7318,N_7216);
nor U8155 (N_8155,N_7913,N_7865);
or U8156 (N_8156,N_7963,N_7735);
or U8157 (N_8157,N_7577,N_7973);
nor U8158 (N_8158,N_7357,N_7316);
nand U8159 (N_8159,N_7633,N_7335);
xnor U8160 (N_8160,N_7857,N_7981);
nand U8161 (N_8161,N_7522,N_7255);
nor U8162 (N_8162,N_7853,N_7625);
xor U8163 (N_8163,N_7513,N_7878);
xor U8164 (N_8164,N_7439,N_7957);
xor U8165 (N_8165,N_7682,N_7291);
and U8166 (N_8166,N_7595,N_7693);
xor U8167 (N_8167,N_7497,N_7428);
xnor U8168 (N_8168,N_7221,N_7271);
or U8169 (N_8169,N_7505,N_7666);
nand U8170 (N_8170,N_7489,N_7920);
or U8171 (N_8171,N_7267,N_7504);
xor U8172 (N_8172,N_7542,N_7602);
or U8173 (N_8173,N_7728,N_7870);
and U8174 (N_8174,N_7309,N_7431);
nor U8175 (N_8175,N_7810,N_7208);
or U8176 (N_8176,N_7847,N_7655);
or U8177 (N_8177,N_7826,N_7952);
and U8178 (N_8178,N_7624,N_7991);
or U8179 (N_8179,N_7416,N_7900);
or U8180 (N_8180,N_7463,N_7717);
and U8181 (N_8181,N_7262,N_7676);
nor U8182 (N_8182,N_7319,N_7593);
or U8183 (N_8183,N_7590,N_7968);
and U8184 (N_8184,N_7560,N_7565);
and U8185 (N_8185,N_7673,N_7236);
xor U8186 (N_8186,N_7253,N_7736);
or U8187 (N_8187,N_7575,N_7654);
and U8188 (N_8188,N_7771,N_7867);
nor U8189 (N_8189,N_7259,N_7881);
xnor U8190 (N_8190,N_7987,N_7455);
nor U8191 (N_8191,N_7781,N_7523);
nor U8192 (N_8192,N_7849,N_7804);
and U8193 (N_8193,N_7954,N_7406);
xnor U8194 (N_8194,N_7821,N_7869);
or U8195 (N_8195,N_7893,N_7418);
or U8196 (N_8196,N_7244,N_7844);
nand U8197 (N_8197,N_7918,N_7875);
nand U8198 (N_8198,N_7770,N_7989);
or U8199 (N_8199,N_7585,N_7882);
and U8200 (N_8200,N_7700,N_7965);
and U8201 (N_8201,N_7797,N_7285);
xor U8202 (N_8202,N_7636,N_7937);
xor U8203 (N_8203,N_7363,N_7562);
and U8204 (N_8204,N_7448,N_7626);
nor U8205 (N_8205,N_7230,N_7825);
xor U8206 (N_8206,N_7432,N_7301);
or U8207 (N_8207,N_7200,N_7531);
nand U8208 (N_8208,N_7365,N_7868);
nor U8209 (N_8209,N_7762,N_7943);
and U8210 (N_8210,N_7374,N_7856);
or U8211 (N_8211,N_7783,N_7589);
nor U8212 (N_8212,N_7393,N_7765);
xnor U8213 (N_8213,N_7828,N_7813);
nor U8214 (N_8214,N_7614,N_7399);
nand U8215 (N_8215,N_7412,N_7782);
nand U8216 (N_8216,N_7414,N_7481);
xnor U8217 (N_8217,N_7689,N_7488);
and U8218 (N_8218,N_7705,N_7364);
nand U8219 (N_8219,N_7424,N_7711);
nand U8220 (N_8220,N_7402,N_7201);
xnor U8221 (N_8221,N_7664,N_7955);
nor U8222 (N_8222,N_7467,N_7475);
nor U8223 (N_8223,N_7596,N_7938);
or U8224 (N_8224,N_7337,N_7681);
or U8225 (N_8225,N_7580,N_7304);
and U8226 (N_8226,N_7491,N_7708);
nor U8227 (N_8227,N_7360,N_7413);
nand U8228 (N_8228,N_7254,N_7866);
nor U8229 (N_8229,N_7747,N_7249);
or U8230 (N_8230,N_7786,N_7211);
xnor U8231 (N_8231,N_7353,N_7788);
xnor U8232 (N_8232,N_7498,N_7544);
nor U8233 (N_8233,N_7742,N_7451);
or U8234 (N_8234,N_7279,N_7889);
or U8235 (N_8235,N_7572,N_7411);
or U8236 (N_8236,N_7368,N_7741);
or U8237 (N_8237,N_7713,N_7331);
and U8238 (N_8238,N_7756,N_7769);
nand U8239 (N_8239,N_7426,N_7997);
or U8240 (N_8240,N_7873,N_7701);
and U8241 (N_8241,N_7336,N_7675);
and U8242 (N_8242,N_7495,N_7457);
nand U8243 (N_8243,N_7718,N_7835);
xor U8244 (N_8244,N_7212,N_7634);
and U8245 (N_8245,N_7739,N_7528);
and U8246 (N_8246,N_7671,N_7458);
or U8247 (N_8247,N_7999,N_7592);
xnor U8248 (N_8248,N_7509,N_7914);
nand U8249 (N_8249,N_7435,N_7934);
nand U8250 (N_8250,N_7321,N_7662);
and U8251 (N_8251,N_7944,N_7905);
or U8252 (N_8252,N_7864,N_7220);
or U8253 (N_8253,N_7648,N_7603);
or U8254 (N_8254,N_7894,N_7293);
xor U8255 (N_8255,N_7478,N_7582);
xnor U8256 (N_8256,N_7967,N_7573);
and U8257 (N_8257,N_7979,N_7935);
nor U8258 (N_8258,N_7984,N_7391);
nor U8259 (N_8259,N_7690,N_7240);
and U8260 (N_8260,N_7831,N_7500);
nand U8261 (N_8261,N_7939,N_7983);
and U8262 (N_8262,N_7930,N_7346);
xor U8263 (N_8263,N_7776,N_7951);
nor U8264 (N_8264,N_7429,N_7617);
and U8265 (N_8265,N_7261,N_7730);
nand U8266 (N_8266,N_7829,N_7518);
and U8267 (N_8267,N_7860,N_7273);
xor U8268 (N_8268,N_7422,N_7630);
or U8269 (N_8269,N_7571,N_7525);
and U8270 (N_8270,N_7839,N_7527);
nor U8271 (N_8271,N_7554,N_7464);
xnor U8272 (N_8272,N_7679,N_7313);
and U8273 (N_8273,N_7287,N_7658);
and U8274 (N_8274,N_7510,N_7297);
and U8275 (N_8275,N_7947,N_7824);
nor U8276 (N_8276,N_7508,N_7966);
or U8277 (N_8277,N_7994,N_7862);
xnor U8278 (N_8278,N_7651,N_7845);
nand U8279 (N_8279,N_7956,N_7760);
or U8280 (N_8280,N_7245,N_7476);
nand U8281 (N_8281,N_7387,N_7257);
nor U8282 (N_8282,N_7683,N_7885);
xor U8283 (N_8283,N_7942,N_7506);
and U8284 (N_8284,N_7423,N_7629);
and U8285 (N_8285,N_7303,N_7507);
nor U8286 (N_8286,N_7663,N_7755);
xnor U8287 (N_8287,N_7773,N_7936);
and U8288 (N_8288,N_7725,N_7310);
nand U8289 (N_8289,N_7512,N_7729);
nand U8290 (N_8290,N_7366,N_7252);
or U8291 (N_8291,N_7559,N_7372);
and U8292 (N_8292,N_7591,N_7473);
nor U8293 (N_8293,N_7515,N_7621);
nor U8294 (N_8294,N_7846,N_7992);
and U8295 (N_8295,N_7719,N_7320);
nand U8296 (N_8296,N_7358,N_7444);
or U8297 (N_8297,N_7723,N_7384);
or U8298 (N_8298,N_7232,N_7884);
xor U8299 (N_8299,N_7886,N_7371);
nor U8300 (N_8300,N_7536,N_7922);
nor U8301 (N_8301,N_7960,N_7680);
nand U8302 (N_8302,N_7722,N_7597);
nand U8303 (N_8303,N_7524,N_7248);
and U8304 (N_8304,N_7790,N_7733);
or U8305 (N_8305,N_7772,N_7217);
and U8306 (N_8306,N_7600,N_7214);
and U8307 (N_8307,N_7726,N_7342);
and U8308 (N_8308,N_7311,N_7355);
nand U8309 (N_8309,N_7852,N_7926);
or U8310 (N_8310,N_7640,N_7855);
and U8311 (N_8311,N_7462,N_7570);
xnor U8312 (N_8312,N_7858,N_7911);
nand U8313 (N_8313,N_7657,N_7811);
or U8314 (N_8314,N_7644,N_7661);
xor U8315 (N_8315,N_7832,N_7704);
or U8316 (N_8316,N_7692,N_7219);
and U8317 (N_8317,N_7526,N_7912);
or U8318 (N_8318,N_7848,N_7574);
nor U8319 (N_8319,N_7850,N_7677);
nor U8320 (N_8320,N_7699,N_7477);
or U8321 (N_8321,N_7296,N_7449);
or U8322 (N_8322,N_7329,N_7953);
nand U8323 (N_8323,N_7761,N_7382);
nor U8324 (N_8324,N_7961,N_7338);
nor U8325 (N_8325,N_7803,N_7437);
nor U8326 (N_8326,N_7915,N_7843);
or U8327 (N_8327,N_7471,N_7685);
nand U8328 (N_8328,N_7638,N_7707);
or U8329 (N_8329,N_7972,N_7421);
and U8330 (N_8330,N_7880,N_7622);
xnor U8331 (N_8331,N_7472,N_7327);
nor U8332 (N_8332,N_7538,N_7732);
xnor U8333 (N_8333,N_7558,N_7601);
or U8334 (N_8334,N_7276,N_7959);
xnor U8335 (N_8335,N_7434,N_7903);
xor U8336 (N_8336,N_7996,N_7420);
and U8337 (N_8337,N_7362,N_7235);
nand U8338 (N_8338,N_7302,N_7407);
nand U8339 (N_8339,N_7837,N_7974);
nor U8340 (N_8340,N_7653,N_7876);
and U8341 (N_8341,N_7492,N_7289);
xnor U8342 (N_8342,N_7703,N_7775);
xnor U8343 (N_8343,N_7535,N_7493);
nand U8344 (N_8344,N_7871,N_7801);
and U8345 (N_8345,N_7976,N_7415);
or U8346 (N_8346,N_7469,N_7940);
xnor U8347 (N_8347,N_7687,N_7611);
or U8348 (N_8348,N_7778,N_7258);
nand U8349 (N_8349,N_7635,N_7632);
xor U8350 (N_8350,N_7394,N_7557);
nand U8351 (N_8351,N_7695,N_7550);
or U8352 (N_8352,N_7222,N_7207);
xor U8353 (N_8353,N_7754,N_7610);
and U8354 (N_8354,N_7292,N_7284);
nor U8355 (N_8355,N_7298,N_7385);
nor U8356 (N_8356,N_7917,N_7553);
nand U8357 (N_8357,N_7793,N_7581);
nor U8358 (N_8358,N_7210,N_7369);
and U8359 (N_8359,N_7441,N_7237);
nand U8360 (N_8360,N_7215,N_7817);
xor U8361 (N_8361,N_7647,N_7377);
nor U8362 (N_8362,N_7461,N_7294);
nand U8363 (N_8363,N_7470,N_7569);
or U8364 (N_8364,N_7686,N_7440);
and U8365 (N_8365,N_7927,N_7567);
or U8366 (N_8366,N_7830,N_7341);
and U8367 (N_8367,N_7339,N_7238);
nor U8368 (N_8368,N_7619,N_7376);
nor U8369 (N_8369,N_7511,N_7827);
or U8370 (N_8370,N_7606,N_7486);
nand U8371 (N_8371,N_7750,N_7785);
or U8372 (N_8372,N_7251,N_7887);
nand U8373 (N_8373,N_7950,N_7452);
nor U8374 (N_8374,N_7665,N_7398);
or U8375 (N_8375,N_7924,N_7854);
nor U8376 (N_8376,N_7579,N_7468);
or U8377 (N_8377,N_7223,N_7436);
and U8378 (N_8378,N_7395,N_7226);
nor U8379 (N_8379,N_7324,N_7351);
nand U8380 (N_8380,N_7206,N_7977);
or U8381 (N_8381,N_7256,N_7901);
nor U8382 (N_8382,N_7758,N_7748);
xnor U8383 (N_8383,N_7851,N_7443);
nor U8384 (N_8384,N_7282,N_7993);
nor U8385 (N_8385,N_7998,N_7405);
xor U8386 (N_8386,N_7541,N_7696);
xor U8387 (N_8387,N_7896,N_7641);
nand U8388 (N_8388,N_7397,N_7224);
nand U8389 (N_8389,N_7709,N_7627);
nand U8390 (N_8390,N_7308,N_7637);
or U8391 (N_8391,N_7818,N_7325);
and U8392 (N_8392,N_7485,N_7566);
nor U8393 (N_8393,N_7442,N_7317);
nor U8394 (N_8394,N_7306,N_7280);
nand U8395 (N_8395,N_7250,N_7356);
or U8396 (N_8396,N_7520,N_7272);
or U8397 (N_8397,N_7227,N_7948);
and U8398 (N_8398,N_7751,N_7347);
and U8399 (N_8399,N_7815,N_7746);
and U8400 (N_8400,N_7301,N_7656);
nand U8401 (N_8401,N_7389,N_7593);
nor U8402 (N_8402,N_7646,N_7860);
and U8403 (N_8403,N_7775,N_7942);
nand U8404 (N_8404,N_7318,N_7316);
or U8405 (N_8405,N_7667,N_7990);
or U8406 (N_8406,N_7751,N_7641);
xnor U8407 (N_8407,N_7819,N_7576);
and U8408 (N_8408,N_7540,N_7442);
and U8409 (N_8409,N_7516,N_7219);
and U8410 (N_8410,N_7246,N_7763);
nor U8411 (N_8411,N_7246,N_7507);
nor U8412 (N_8412,N_7581,N_7338);
xor U8413 (N_8413,N_7774,N_7853);
nor U8414 (N_8414,N_7388,N_7686);
or U8415 (N_8415,N_7384,N_7838);
or U8416 (N_8416,N_7528,N_7524);
and U8417 (N_8417,N_7760,N_7836);
xnor U8418 (N_8418,N_7596,N_7309);
or U8419 (N_8419,N_7816,N_7516);
or U8420 (N_8420,N_7306,N_7403);
and U8421 (N_8421,N_7393,N_7372);
or U8422 (N_8422,N_7363,N_7312);
or U8423 (N_8423,N_7963,N_7230);
or U8424 (N_8424,N_7283,N_7436);
xor U8425 (N_8425,N_7661,N_7830);
and U8426 (N_8426,N_7770,N_7224);
xnor U8427 (N_8427,N_7860,N_7829);
or U8428 (N_8428,N_7884,N_7350);
and U8429 (N_8429,N_7353,N_7511);
nor U8430 (N_8430,N_7979,N_7839);
and U8431 (N_8431,N_7335,N_7474);
nand U8432 (N_8432,N_7577,N_7831);
nand U8433 (N_8433,N_7205,N_7315);
or U8434 (N_8434,N_7364,N_7495);
xnor U8435 (N_8435,N_7552,N_7257);
nor U8436 (N_8436,N_7667,N_7974);
xor U8437 (N_8437,N_7762,N_7343);
or U8438 (N_8438,N_7942,N_7608);
nor U8439 (N_8439,N_7222,N_7612);
and U8440 (N_8440,N_7365,N_7532);
and U8441 (N_8441,N_7452,N_7467);
xnor U8442 (N_8442,N_7609,N_7985);
nand U8443 (N_8443,N_7623,N_7427);
xor U8444 (N_8444,N_7906,N_7808);
or U8445 (N_8445,N_7626,N_7854);
nand U8446 (N_8446,N_7826,N_7970);
nor U8447 (N_8447,N_7415,N_7599);
or U8448 (N_8448,N_7784,N_7732);
and U8449 (N_8449,N_7627,N_7227);
or U8450 (N_8450,N_7550,N_7813);
xnor U8451 (N_8451,N_7834,N_7997);
nand U8452 (N_8452,N_7726,N_7892);
nor U8453 (N_8453,N_7679,N_7714);
xnor U8454 (N_8454,N_7454,N_7902);
nand U8455 (N_8455,N_7915,N_7556);
nand U8456 (N_8456,N_7606,N_7802);
and U8457 (N_8457,N_7402,N_7277);
nand U8458 (N_8458,N_7594,N_7276);
or U8459 (N_8459,N_7418,N_7482);
nor U8460 (N_8460,N_7505,N_7401);
nand U8461 (N_8461,N_7653,N_7500);
and U8462 (N_8462,N_7325,N_7202);
nand U8463 (N_8463,N_7285,N_7578);
and U8464 (N_8464,N_7489,N_7500);
and U8465 (N_8465,N_7549,N_7696);
or U8466 (N_8466,N_7835,N_7876);
or U8467 (N_8467,N_7378,N_7565);
and U8468 (N_8468,N_7254,N_7340);
nand U8469 (N_8469,N_7639,N_7564);
and U8470 (N_8470,N_7973,N_7844);
nand U8471 (N_8471,N_7223,N_7419);
nand U8472 (N_8472,N_7816,N_7576);
or U8473 (N_8473,N_7449,N_7608);
nor U8474 (N_8474,N_7501,N_7957);
or U8475 (N_8475,N_7461,N_7871);
nor U8476 (N_8476,N_7832,N_7403);
nand U8477 (N_8477,N_7586,N_7659);
or U8478 (N_8478,N_7434,N_7698);
nor U8479 (N_8479,N_7829,N_7217);
or U8480 (N_8480,N_7913,N_7764);
nor U8481 (N_8481,N_7810,N_7222);
nand U8482 (N_8482,N_7640,N_7818);
and U8483 (N_8483,N_7343,N_7592);
or U8484 (N_8484,N_7418,N_7911);
xor U8485 (N_8485,N_7902,N_7943);
or U8486 (N_8486,N_7708,N_7315);
nand U8487 (N_8487,N_7497,N_7701);
or U8488 (N_8488,N_7345,N_7284);
nor U8489 (N_8489,N_7740,N_7841);
or U8490 (N_8490,N_7707,N_7286);
xnor U8491 (N_8491,N_7326,N_7336);
nor U8492 (N_8492,N_7674,N_7940);
and U8493 (N_8493,N_7598,N_7271);
nor U8494 (N_8494,N_7518,N_7303);
nor U8495 (N_8495,N_7564,N_7679);
and U8496 (N_8496,N_7879,N_7963);
or U8497 (N_8497,N_7635,N_7824);
xnor U8498 (N_8498,N_7213,N_7711);
or U8499 (N_8499,N_7919,N_7605);
or U8500 (N_8500,N_7286,N_7924);
xor U8501 (N_8501,N_7235,N_7731);
nor U8502 (N_8502,N_7947,N_7932);
xor U8503 (N_8503,N_7637,N_7799);
nor U8504 (N_8504,N_7370,N_7532);
xnor U8505 (N_8505,N_7657,N_7750);
nor U8506 (N_8506,N_7577,N_7274);
nand U8507 (N_8507,N_7908,N_7710);
and U8508 (N_8508,N_7821,N_7956);
xor U8509 (N_8509,N_7327,N_7896);
or U8510 (N_8510,N_7417,N_7850);
and U8511 (N_8511,N_7401,N_7646);
nand U8512 (N_8512,N_7263,N_7405);
or U8513 (N_8513,N_7824,N_7975);
xnor U8514 (N_8514,N_7419,N_7423);
nor U8515 (N_8515,N_7232,N_7498);
and U8516 (N_8516,N_7771,N_7949);
nor U8517 (N_8517,N_7362,N_7701);
xor U8518 (N_8518,N_7459,N_7901);
nor U8519 (N_8519,N_7985,N_7320);
nor U8520 (N_8520,N_7631,N_7340);
nand U8521 (N_8521,N_7581,N_7699);
and U8522 (N_8522,N_7314,N_7864);
nand U8523 (N_8523,N_7787,N_7619);
or U8524 (N_8524,N_7213,N_7271);
and U8525 (N_8525,N_7895,N_7560);
xnor U8526 (N_8526,N_7956,N_7304);
nand U8527 (N_8527,N_7419,N_7488);
xnor U8528 (N_8528,N_7552,N_7698);
and U8529 (N_8529,N_7903,N_7669);
nand U8530 (N_8530,N_7835,N_7600);
xor U8531 (N_8531,N_7732,N_7507);
nand U8532 (N_8532,N_7629,N_7472);
or U8533 (N_8533,N_7873,N_7875);
nand U8534 (N_8534,N_7678,N_7679);
nor U8535 (N_8535,N_7870,N_7704);
nand U8536 (N_8536,N_7212,N_7260);
or U8537 (N_8537,N_7559,N_7770);
and U8538 (N_8538,N_7539,N_7232);
nor U8539 (N_8539,N_7412,N_7729);
or U8540 (N_8540,N_7617,N_7962);
xnor U8541 (N_8541,N_7594,N_7961);
or U8542 (N_8542,N_7698,N_7354);
xnor U8543 (N_8543,N_7959,N_7932);
and U8544 (N_8544,N_7976,N_7776);
or U8545 (N_8545,N_7746,N_7585);
xnor U8546 (N_8546,N_7862,N_7928);
or U8547 (N_8547,N_7653,N_7362);
nor U8548 (N_8548,N_7274,N_7863);
xor U8549 (N_8549,N_7632,N_7779);
nor U8550 (N_8550,N_7629,N_7568);
nand U8551 (N_8551,N_7576,N_7441);
or U8552 (N_8552,N_7257,N_7238);
nor U8553 (N_8553,N_7823,N_7383);
nand U8554 (N_8554,N_7580,N_7998);
xnor U8555 (N_8555,N_7744,N_7687);
and U8556 (N_8556,N_7786,N_7742);
nand U8557 (N_8557,N_7350,N_7771);
and U8558 (N_8558,N_7311,N_7667);
xor U8559 (N_8559,N_7654,N_7480);
nor U8560 (N_8560,N_7347,N_7834);
or U8561 (N_8561,N_7951,N_7582);
and U8562 (N_8562,N_7568,N_7233);
nor U8563 (N_8563,N_7596,N_7703);
and U8564 (N_8564,N_7447,N_7914);
nand U8565 (N_8565,N_7688,N_7322);
or U8566 (N_8566,N_7367,N_7460);
nor U8567 (N_8567,N_7933,N_7575);
and U8568 (N_8568,N_7677,N_7378);
and U8569 (N_8569,N_7313,N_7877);
nand U8570 (N_8570,N_7239,N_7244);
nor U8571 (N_8571,N_7306,N_7455);
and U8572 (N_8572,N_7404,N_7208);
and U8573 (N_8573,N_7677,N_7672);
nand U8574 (N_8574,N_7432,N_7455);
nand U8575 (N_8575,N_7660,N_7457);
xor U8576 (N_8576,N_7417,N_7986);
and U8577 (N_8577,N_7685,N_7782);
xnor U8578 (N_8578,N_7286,N_7819);
or U8579 (N_8579,N_7471,N_7477);
and U8580 (N_8580,N_7657,N_7559);
and U8581 (N_8581,N_7898,N_7312);
nand U8582 (N_8582,N_7978,N_7542);
and U8583 (N_8583,N_7555,N_7627);
and U8584 (N_8584,N_7696,N_7322);
xor U8585 (N_8585,N_7815,N_7429);
nor U8586 (N_8586,N_7345,N_7633);
or U8587 (N_8587,N_7440,N_7629);
nor U8588 (N_8588,N_7313,N_7233);
xnor U8589 (N_8589,N_7501,N_7434);
or U8590 (N_8590,N_7298,N_7836);
nor U8591 (N_8591,N_7577,N_7722);
nor U8592 (N_8592,N_7689,N_7200);
xnor U8593 (N_8593,N_7926,N_7263);
nand U8594 (N_8594,N_7934,N_7480);
or U8595 (N_8595,N_7432,N_7864);
and U8596 (N_8596,N_7990,N_7216);
and U8597 (N_8597,N_7393,N_7946);
xor U8598 (N_8598,N_7318,N_7328);
and U8599 (N_8599,N_7347,N_7831);
xnor U8600 (N_8600,N_7395,N_7389);
and U8601 (N_8601,N_7886,N_7552);
nor U8602 (N_8602,N_7222,N_7329);
or U8603 (N_8603,N_7301,N_7763);
and U8604 (N_8604,N_7486,N_7994);
and U8605 (N_8605,N_7643,N_7663);
nor U8606 (N_8606,N_7462,N_7411);
xnor U8607 (N_8607,N_7934,N_7878);
xnor U8608 (N_8608,N_7837,N_7983);
nand U8609 (N_8609,N_7939,N_7675);
xor U8610 (N_8610,N_7927,N_7626);
xor U8611 (N_8611,N_7652,N_7778);
or U8612 (N_8612,N_7713,N_7563);
nor U8613 (N_8613,N_7406,N_7713);
xnor U8614 (N_8614,N_7244,N_7732);
nand U8615 (N_8615,N_7570,N_7403);
nand U8616 (N_8616,N_7576,N_7842);
xor U8617 (N_8617,N_7326,N_7511);
or U8618 (N_8618,N_7844,N_7267);
nor U8619 (N_8619,N_7611,N_7569);
or U8620 (N_8620,N_7776,N_7893);
nor U8621 (N_8621,N_7270,N_7739);
xor U8622 (N_8622,N_7228,N_7421);
nor U8623 (N_8623,N_7632,N_7247);
nor U8624 (N_8624,N_7827,N_7630);
nor U8625 (N_8625,N_7256,N_7373);
xnor U8626 (N_8626,N_7282,N_7554);
nand U8627 (N_8627,N_7200,N_7807);
nor U8628 (N_8628,N_7642,N_7232);
xnor U8629 (N_8629,N_7448,N_7508);
or U8630 (N_8630,N_7863,N_7876);
nor U8631 (N_8631,N_7827,N_7927);
nor U8632 (N_8632,N_7342,N_7335);
and U8633 (N_8633,N_7733,N_7465);
nand U8634 (N_8634,N_7485,N_7726);
and U8635 (N_8635,N_7992,N_7453);
or U8636 (N_8636,N_7972,N_7293);
nand U8637 (N_8637,N_7927,N_7838);
nand U8638 (N_8638,N_7263,N_7808);
or U8639 (N_8639,N_7465,N_7485);
nand U8640 (N_8640,N_7345,N_7332);
and U8641 (N_8641,N_7591,N_7645);
xnor U8642 (N_8642,N_7612,N_7982);
or U8643 (N_8643,N_7326,N_7293);
nand U8644 (N_8644,N_7708,N_7539);
and U8645 (N_8645,N_7601,N_7602);
nand U8646 (N_8646,N_7960,N_7334);
and U8647 (N_8647,N_7894,N_7654);
and U8648 (N_8648,N_7549,N_7376);
nor U8649 (N_8649,N_7614,N_7293);
nor U8650 (N_8650,N_7938,N_7576);
nor U8651 (N_8651,N_7687,N_7338);
xor U8652 (N_8652,N_7264,N_7504);
and U8653 (N_8653,N_7339,N_7336);
nand U8654 (N_8654,N_7707,N_7391);
nor U8655 (N_8655,N_7669,N_7947);
and U8656 (N_8656,N_7647,N_7778);
and U8657 (N_8657,N_7890,N_7521);
or U8658 (N_8658,N_7596,N_7942);
nand U8659 (N_8659,N_7569,N_7804);
nand U8660 (N_8660,N_7425,N_7365);
and U8661 (N_8661,N_7985,N_7696);
nor U8662 (N_8662,N_7959,N_7969);
xnor U8663 (N_8663,N_7487,N_7610);
or U8664 (N_8664,N_7395,N_7457);
and U8665 (N_8665,N_7768,N_7850);
nand U8666 (N_8666,N_7992,N_7668);
nand U8667 (N_8667,N_7854,N_7921);
xor U8668 (N_8668,N_7572,N_7382);
xor U8669 (N_8669,N_7966,N_7367);
nor U8670 (N_8670,N_7293,N_7884);
nand U8671 (N_8671,N_7394,N_7810);
or U8672 (N_8672,N_7958,N_7639);
nor U8673 (N_8673,N_7951,N_7466);
or U8674 (N_8674,N_7474,N_7900);
nand U8675 (N_8675,N_7880,N_7610);
or U8676 (N_8676,N_7908,N_7211);
xnor U8677 (N_8677,N_7681,N_7264);
xor U8678 (N_8678,N_7382,N_7983);
or U8679 (N_8679,N_7618,N_7347);
and U8680 (N_8680,N_7847,N_7668);
nor U8681 (N_8681,N_7453,N_7804);
and U8682 (N_8682,N_7634,N_7369);
nor U8683 (N_8683,N_7262,N_7699);
and U8684 (N_8684,N_7663,N_7871);
xnor U8685 (N_8685,N_7427,N_7887);
nor U8686 (N_8686,N_7249,N_7885);
nand U8687 (N_8687,N_7935,N_7407);
and U8688 (N_8688,N_7344,N_7529);
nand U8689 (N_8689,N_7788,N_7750);
and U8690 (N_8690,N_7608,N_7245);
nor U8691 (N_8691,N_7686,N_7810);
xnor U8692 (N_8692,N_7456,N_7581);
nand U8693 (N_8693,N_7598,N_7636);
nor U8694 (N_8694,N_7391,N_7814);
nand U8695 (N_8695,N_7348,N_7352);
or U8696 (N_8696,N_7825,N_7545);
and U8697 (N_8697,N_7341,N_7478);
nor U8698 (N_8698,N_7765,N_7712);
nand U8699 (N_8699,N_7278,N_7878);
nor U8700 (N_8700,N_7969,N_7840);
nor U8701 (N_8701,N_7733,N_7989);
xor U8702 (N_8702,N_7444,N_7215);
and U8703 (N_8703,N_7695,N_7579);
and U8704 (N_8704,N_7530,N_7588);
nand U8705 (N_8705,N_7332,N_7265);
or U8706 (N_8706,N_7583,N_7979);
nand U8707 (N_8707,N_7973,N_7823);
nor U8708 (N_8708,N_7958,N_7262);
xor U8709 (N_8709,N_7615,N_7298);
nand U8710 (N_8710,N_7417,N_7646);
nand U8711 (N_8711,N_7792,N_7881);
or U8712 (N_8712,N_7987,N_7639);
or U8713 (N_8713,N_7983,N_7976);
or U8714 (N_8714,N_7550,N_7821);
nand U8715 (N_8715,N_7654,N_7242);
nor U8716 (N_8716,N_7350,N_7679);
nor U8717 (N_8717,N_7921,N_7223);
nand U8718 (N_8718,N_7571,N_7870);
nand U8719 (N_8719,N_7851,N_7592);
nand U8720 (N_8720,N_7449,N_7256);
nand U8721 (N_8721,N_7486,N_7976);
xor U8722 (N_8722,N_7733,N_7344);
xor U8723 (N_8723,N_7805,N_7479);
xor U8724 (N_8724,N_7679,N_7657);
or U8725 (N_8725,N_7591,N_7795);
or U8726 (N_8726,N_7727,N_7663);
and U8727 (N_8727,N_7983,N_7635);
xnor U8728 (N_8728,N_7720,N_7775);
xor U8729 (N_8729,N_7674,N_7517);
nor U8730 (N_8730,N_7527,N_7508);
or U8731 (N_8731,N_7926,N_7344);
or U8732 (N_8732,N_7982,N_7555);
or U8733 (N_8733,N_7817,N_7617);
nor U8734 (N_8734,N_7473,N_7415);
and U8735 (N_8735,N_7652,N_7485);
and U8736 (N_8736,N_7221,N_7211);
nor U8737 (N_8737,N_7943,N_7840);
nor U8738 (N_8738,N_7968,N_7602);
nand U8739 (N_8739,N_7799,N_7281);
and U8740 (N_8740,N_7682,N_7816);
nor U8741 (N_8741,N_7946,N_7622);
nand U8742 (N_8742,N_7653,N_7563);
and U8743 (N_8743,N_7996,N_7693);
nand U8744 (N_8744,N_7870,N_7768);
nand U8745 (N_8745,N_7553,N_7679);
xor U8746 (N_8746,N_7798,N_7575);
nand U8747 (N_8747,N_7281,N_7982);
or U8748 (N_8748,N_7200,N_7206);
nand U8749 (N_8749,N_7647,N_7862);
or U8750 (N_8750,N_7355,N_7643);
nor U8751 (N_8751,N_7603,N_7304);
or U8752 (N_8752,N_7281,N_7888);
nor U8753 (N_8753,N_7919,N_7549);
and U8754 (N_8754,N_7208,N_7313);
or U8755 (N_8755,N_7587,N_7597);
nand U8756 (N_8756,N_7502,N_7371);
nand U8757 (N_8757,N_7885,N_7980);
xnor U8758 (N_8758,N_7756,N_7722);
nor U8759 (N_8759,N_7999,N_7616);
or U8760 (N_8760,N_7260,N_7763);
xor U8761 (N_8761,N_7882,N_7929);
or U8762 (N_8762,N_7500,N_7248);
and U8763 (N_8763,N_7965,N_7842);
nor U8764 (N_8764,N_7718,N_7384);
xor U8765 (N_8765,N_7952,N_7698);
nor U8766 (N_8766,N_7562,N_7942);
xnor U8767 (N_8767,N_7645,N_7452);
xor U8768 (N_8768,N_7214,N_7267);
and U8769 (N_8769,N_7737,N_7641);
nor U8770 (N_8770,N_7609,N_7406);
and U8771 (N_8771,N_7558,N_7562);
or U8772 (N_8772,N_7894,N_7467);
or U8773 (N_8773,N_7238,N_7900);
nand U8774 (N_8774,N_7377,N_7810);
or U8775 (N_8775,N_7349,N_7860);
nor U8776 (N_8776,N_7496,N_7286);
and U8777 (N_8777,N_7253,N_7758);
nand U8778 (N_8778,N_7344,N_7200);
and U8779 (N_8779,N_7802,N_7778);
and U8780 (N_8780,N_7266,N_7414);
and U8781 (N_8781,N_7979,N_7672);
nor U8782 (N_8782,N_7885,N_7244);
xnor U8783 (N_8783,N_7481,N_7614);
nor U8784 (N_8784,N_7391,N_7771);
and U8785 (N_8785,N_7354,N_7258);
nor U8786 (N_8786,N_7471,N_7534);
and U8787 (N_8787,N_7262,N_7983);
nand U8788 (N_8788,N_7267,N_7865);
or U8789 (N_8789,N_7428,N_7723);
or U8790 (N_8790,N_7836,N_7207);
nand U8791 (N_8791,N_7336,N_7886);
xnor U8792 (N_8792,N_7539,N_7619);
or U8793 (N_8793,N_7545,N_7716);
xnor U8794 (N_8794,N_7768,N_7636);
nand U8795 (N_8795,N_7540,N_7966);
nor U8796 (N_8796,N_7837,N_7989);
or U8797 (N_8797,N_7849,N_7603);
nor U8798 (N_8798,N_7868,N_7833);
or U8799 (N_8799,N_7866,N_7948);
nand U8800 (N_8800,N_8188,N_8481);
nand U8801 (N_8801,N_8775,N_8045);
or U8802 (N_8802,N_8435,N_8543);
and U8803 (N_8803,N_8272,N_8461);
nor U8804 (N_8804,N_8055,N_8632);
xor U8805 (N_8805,N_8370,N_8722);
nand U8806 (N_8806,N_8669,N_8639);
or U8807 (N_8807,N_8303,N_8578);
or U8808 (N_8808,N_8372,N_8706);
and U8809 (N_8809,N_8593,N_8193);
nor U8810 (N_8810,N_8128,N_8641);
xnor U8811 (N_8811,N_8287,N_8163);
or U8812 (N_8812,N_8711,N_8605);
or U8813 (N_8813,N_8222,N_8522);
and U8814 (N_8814,N_8262,N_8308);
or U8815 (N_8815,N_8601,N_8337);
xnor U8816 (N_8816,N_8012,N_8375);
nor U8817 (N_8817,N_8268,N_8379);
or U8818 (N_8818,N_8048,N_8073);
or U8819 (N_8819,N_8058,N_8344);
and U8820 (N_8820,N_8071,N_8397);
nor U8821 (N_8821,N_8657,N_8716);
nor U8822 (N_8822,N_8713,N_8220);
and U8823 (N_8823,N_8123,N_8118);
xnor U8824 (N_8824,N_8213,N_8442);
and U8825 (N_8825,N_8021,N_8567);
and U8826 (N_8826,N_8537,N_8033);
nand U8827 (N_8827,N_8340,N_8628);
or U8828 (N_8828,N_8462,N_8078);
or U8829 (N_8829,N_8156,N_8784);
xnor U8830 (N_8830,N_8176,N_8358);
nand U8831 (N_8831,N_8691,N_8398);
xor U8832 (N_8832,N_8394,N_8470);
and U8833 (N_8833,N_8256,N_8650);
nand U8834 (N_8834,N_8257,N_8228);
nor U8835 (N_8835,N_8153,N_8203);
nor U8836 (N_8836,N_8161,N_8009);
nor U8837 (N_8837,N_8672,N_8430);
and U8838 (N_8838,N_8260,N_8539);
nand U8839 (N_8839,N_8062,N_8454);
xnor U8840 (N_8840,N_8647,N_8721);
nand U8841 (N_8841,N_8338,N_8393);
nor U8842 (N_8842,N_8286,N_8141);
or U8843 (N_8843,N_8006,N_8356);
or U8844 (N_8844,N_8757,N_8588);
nor U8845 (N_8845,N_8290,N_8135);
and U8846 (N_8846,N_8793,N_8490);
or U8847 (N_8847,N_8507,N_8771);
nand U8848 (N_8848,N_8486,N_8020);
or U8849 (N_8849,N_8720,N_8703);
nor U8850 (N_8850,N_8634,N_8158);
or U8851 (N_8851,N_8319,N_8038);
xnor U8852 (N_8852,N_8556,N_8190);
and U8853 (N_8853,N_8504,N_8496);
nand U8854 (N_8854,N_8365,N_8354);
and U8855 (N_8855,N_8758,N_8261);
nor U8856 (N_8856,N_8767,N_8705);
nor U8857 (N_8857,N_8041,N_8224);
nand U8858 (N_8858,N_8770,N_8031);
or U8859 (N_8859,N_8205,N_8513);
or U8860 (N_8860,N_8312,N_8534);
or U8861 (N_8861,N_8626,N_8243);
xor U8862 (N_8862,N_8573,N_8113);
nor U8863 (N_8863,N_8212,N_8408);
and U8864 (N_8864,N_8059,N_8659);
or U8865 (N_8865,N_8525,N_8640);
or U8866 (N_8866,N_8446,N_8204);
xor U8867 (N_8867,N_8560,N_8665);
nor U8868 (N_8868,N_8182,N_8562);
and U8869 (N_8869,N_8506,N_8702);
and U8870 (N_8870,N_8414,N_8684);
nor U8871 (N_8871,N_8331,N_8094);
nor U8872 (N_8872,N_8581,N_8503);
xnor U8873 (N_8873,N_8075,N_8599);
xnor U8874 (N_8874,N_8271,N_8277);
and U8875 (N_8875,N_8255,N_8421);
xnor U8876 (N_8876,N_8149,N_8115);
nor U8877 (N_8877,N_8552,N_8388);
or U8878 (N_8878,N_8645,N_8401);
nor U8879 (N_8879,N_8422,N_8744);
or U8880 (N_8880,N_8671,N_8494);
nor U8881 (N_8881,N_8316,N_8072);
or U8882 (N_8882,N_8511,N_8779);
nor U8883 (N_8883,N_8112,N_8416);
xor U8884 (N_8884,N_8371,N_8551);
and U8885 (N_8885,N_8774,N_8472);
or U8886 (N_8886,N_8039,N_8745);
xor U8887 (N_8887,N_8142,N_8281);
xnor U8888 (N_8888,N_8776,N_8196);
or U8889 (N_8889,N_8107,N_8791);
nand U8890 (N_8890,N_8542,N_8291);
nand U8891 (N_8891,N_8509,N_8164);
nor U8892 (N_8892,N_8649,N_8199);
nand U8893 (N_8893,N_8415,N_8780);
xnor U8894 (N_8894,N_8207,N_8748);
xnor U8895 (N_8895,N_8350,N_8307);
nor U8896 (N_8896,N_8417,N_8037);
or U8897 (N_8897,N_8265,N_8455);
or U8898 (N_8898,N_8127,N_8011);
nand U8899 (N_8899,N_8185,N_8318);
nor U8900 (N_8900,N_8610,N_8589);
and U8901 (N_8901,N_8655,N_8437);
xnor U8902 (N_8902,N_8426,N_8413);
nand U8903 (N_8903,N_8679,N_8460);
and U8904 (N_8904,N_8627,N_8574);
xor U8905 (N_8905,N_8476,N_8404);
nor U8906 (N_8906,N_8783,N_8183);
nand U8907 (N_8907,N_8066,N_8051);
nor U8908 (N_8908,N_8150,N_8231);
xor U8909 (N_8909,N_8564,N_8474);
or U8910 (N_8910,N_8607,N_8317);
nand U8911 (N_8911,N_8244,N_8216);
xnor U8912 (N_8912,N_8568,N_8512);
or U8913 (N_8913,N_8355,N_8544);
xor U8914 (N_8914,N_8036,N_8278);
or U8915 (N_8915,N_8615,N_8613);
xor U8916 (N_8916,N_8202,N_8376);
xnor U8917 (N_8917,N_8383,N_8124);
xor U8918 (N_8918,N_8172,N_8138);
nor U8919 (N_8919,N_8391,N_8227);
nand U8920 (N_8920,N_8731,N_8053);
nand U8921 (N_8921,N_8575,N_8042);
nand U8922 (N_8922,N_8034,N_8495);
and U8923 (N_8923,N_8644,N_8248);
nand U8924 (N_8924,N_8425,N_8010);
or U8925 (N_8925,N_8122,N_8154);
nand U8926 (N_8926,N_8366,N_8029);
or U8927 (N_8927,N_8057,N_8368);
xor U8928 (N_8928,N_8184,N_8126);
nor U8929 (N_8929,N_8550,N_8798);
nand U8930 (N_8930,N_8160,N_8019);
nor U8931 (N_8931,N_8483,N_8714);
xnor U8932 (N_8932,N_8710,N_8755);
xnor U8933 (N_8933,N_8590,N_8091);
or U8934 (N_8934,N_8125,N_8535);
nand U8935 (N_8935,N_8345,N_8276);
nand U8936 (N_8936,N_8206,N_8453);
nor U8937 (N_8937,N_8310,N_8274);
nor U8938 (N_8938,N_8546,N_8143);
nor U8939 (N_8939,N_8598,N_8299);
nand U8940 (N_8940,N_8197,N_8616);
nor U8941 (N_8941,N_8173,N_8789);
and U8942 (N_8942,N_8000,N_8389);
or U8943 (N_8943,N_8409,N_8167);
xor U8944 (N_8944,N_8643,N_8467);
xnor U8945 (N_8945,N_8428,N_8768);
or U8946 (N_8946,N_8515,N_8420);
nor U8947 (N_8947,N_8378,N_8517);
nand U8948 (N_8948,N_8580,N_8410);
xnor U8949 (N_8949,N_8781,N_8357);
nor U8950 (N_8950,N_8097,N_8736);
and U8951 (N_8951,N_8148,N_8214);
nand U8952 (N_8952,N_8236,N_8569);
nor U8953 (N_8953,N_8373,N_8471);
nor U8954 (N_8954,N_8166,N_8315);
nor U8955 (N_8955,N_8473,N_8023);
or U8956 (N_8956,N_8364,N_8329);
or U8957 (N_8957,N_8246,N_8549);
or U8958 (N_8958,N_8322,N_8540);
or U8959 (N_8959,N_8129,N_8326);
xor U8960 (N_8960,N_8136,N_8419);
and U8961 (N_8961,N_8050,N_8032);
or U8962 (N_8962,N_8187,N_8336);
and U8963 (N_8963,N_8498,N_8121);
and U8964 (N_8964,N_8445,N_8464);
or U8965 (N_8965,N_8060,N_8024);
nand U8966 (N_8966,N_8772,N_8439);
or U8967 (N_8967,N_8629,N_8762);
and U8968 (N_8968,N_8275,N_8637);
xnor U8969 (N_8969,N_8076,N_8293);
xor U8970 (N_8970,N_8558,N_8225);
or U8971 (N_8971,N_8760,N_8233);
nand U8972 (N_8972,N_8223,N_8014);
and U8973 (N_8973,N_8131,N_8740);
or U8974 (N_8974,N_8186,N_8794);
nand U8975 (N_8975,N_8717,N_8400);
or U8976 (N_8976,N_8480,N_8232);
nand U8977 (N_8977,N_8280,N_8469);
xnor U8978 (N_8978,N_8249,N_8719);
xor U8979 (N_8979,N_8712,N_8374);
or U8980 (N_8980,N_8266,N_8594);
or U8981 (N_8981,N_8418,N_8007);
xnor U8982 (N_8982,N_8104,N_8325);
nor U8983 (N_8983,N_8730,N_8614);
nor U8984 (N_8984,N_8501,N_8254);
xnor U8985 (N_8985,N_8584,N_8510);
and U8986 (N_8986,N_8750,N_8465);
or U8987 (N_8987,N_8282,N_8638);
xnor U8988 (N_8988,N_8683,N_8609);
and U8989 (N_8989,N_8384,N_8521);
xor U8990 (N_8990,N_8001,N_8089);
nand U8991 (N_8991,N_8538,N_8311);
and U8992 (N_8992,N_8458,N_8259);
xor U8993 (N_8993,N_8604,N_8165);
nand U8994 (N_8994,N_8079,N_8238);
and U8995 (N_8995,N_8766,N_8529);
xnor U8996 (N_8996,N_8111,N_8457);
nand U8997 (N_8997,N_8279,N_8102);
xor U8998 (N_8998,N_8074,N_8284);
nand U8999 (N_8999,N_8678,N_8701);
xnor U9000 (N_9000,N_8086,N_8353);
or U9001 (N_9001,N_8219,N_8700);
or U9002 (N_9002,N_8530,N_8668);
xor U9003 (N_9003,N_8352,N_8608);
nor U9004 (N_9004,N_8273,N_8068);
or U9005 (N_9005,N_8570,N_8069);
and U9006 (N_9006,N_8061,N_8606);
or U9007 (N_9007,N_8346,N_8100);
xor U9008 (N_9008,N_8264,N_8734);
or U9009 (N_9009,N_8541,N_8561);
and U9010 (N_9010,N_8170,N_8387);
nand U9011 (N_9011,N_8514,N_8306);
and U9012 (N_9012,N_8497,N_8478);
nor U9013 (N_9013,N_8230,N_8786);
xnor U9014 (N_9014,N_8144,N_8792);
or U9015 (N_9015,N_8587,N_8320);
nand U9016 (N_9016,N_8018,N_8508);
nand U9017 (N_9017,N_8382,N_8399);
xnor U9018 (N_9018,N_8381,N_8162);
nand U9019 (N_9019,N_8585,N_8406);
nor U9020 (N_9020,N_8300,N_8554);
or U9021 (N_9021,N_8013,N_8708);
nand U9022 (N_9022,N_8359,N_8157);
or U9023 (N_9023,N_8052,N_8247);
xnor U9024 (N_9024,N_8433,N_8270);
nor U9025 (N_9025,N_8728,N_8377);
and U9026 (N_9026,N_8690,N_8715);
nor U9027 (N_9027,N_8441,N_8178);
nand U9028 (N_9028,N_8335,N_8309);
nor U9029 (N_9029,N_8002,N_8269);
and U9030 (N_9030,N_8664,N_8524);
and U9031 (N_9031,N_8692,N_8117);
and U9032 (N_9032,N_8682,N_8241);
and U9033 (N_9033,N_8652,N_8630);
nand U9034 (N_9034,N_8595,N_8088);
or U9035 (N_9035,N_8502,N_8674);
or U9036 (N_9036,N_8321,N_8119);
xnor U9037 (N_9037,N_8027,N_8676);
nor U9038 (N_9038,N_8342,N_8092);
or U9039 (N_9039,N_8763,N_8625);
nor U9040 (N_9040,N_8049,N_8407);
or U9041 (N_9041,N_8363,N_8090);
nand U9042 (N_9042,N_8004,N_8545);
or U9043 (N_9043,N_8008,N_8505);
xor U9044 (N_9044,N_8492,N_8695);
xnor U9045 (N_9045,N_8677,N_8648);
nand U9046 (N_9046,N_8210,N_8718);
or U9047 (N_9047,N_8343,N_8171);
or U9048 (N_9048,N_8582,N_8444);
nand U9049 (N_9049,N_8653,N_8084);
and U9050 (N_9050,N_8773,N_8169);
and U9051 (N_9051,N_8189,N_8081);
nor U9052 (N_9052,N_8685,N_8707);
xor U9053 (N_9053,N_8251,N_8137);
and U9054 (N_9054,N_8698,N_8211);
nor U9055 (N_9055,N_8449,N_8566);
or U9056 (N_9056,N_8796,N_8571);
and U9057 (N_9057,N_8016,N_8536);
nand U9058 (N_9058,N_8661,N_8602);
and U9059 (N_9059,N_8603,N_8250);
nor U9060 (N_9060,N_8333,N_8499);
nor U9061 (N_9061,N_8749,N_8330);
and U9062 (N_9062,N_8296,N_8438);
or U9063 (N_9063,N_8611,N_8623);
xor U9064 (N_9064,N_8168,N_8622);
or U9065 (N_9065,N_8459,N_8667);
nor U9066 (N_9066,N_8221,N_8434);
xnor U9067 (N_9067,N_8046,N_8147);
nor U9068 (N_9068,N_8500,N_8636);
nand U9069 (N_9069,N_8132,N_8633);
nand U9070 (N_9070,N_8738,N_8559);
and U9071 (N_9071,N_8283,N_8201);
nor U9072 (N_9072,N_8493,N_8553);
nor U9073 (N_9073,N_8116,N_8047);
and U9074 (N_9074,N_8349,N_8742);
xnor U9075 (N_9075,N_8022,N_8463);
and U9076 (N_9076,N_8479,N_8080);
and U9077 (N_9077,N_8412,N_8452);
or U9078 (N_9078,N_8621,N_8547);
xor U9079 (N_9079,N_8799,N_8294);
nand U9080 (N_9080,N_8596,N_8140);
xnor U9081 (N_9081,N_8101,N_8726);
nand U9082 (N_9082,N_8351,N_8753);
and U9083 (N_9083,N_8735,N_8367);
and U9084 (N_9084,N_8681,N_8323);
nand U9085 (N_9085,N_8488,N_8658);
xor U9086 (N_9086,N_8134,N_8328);
or U9087 (N_9087,N_8332,N_8044);
and U9088 (N_9088,N_8579,N_8788);
nor U9089 (N_9089,N_8313,N_8155);
nor U9090 (N_9090,N_8028,N_8520);
or U9091 (N_9091,N_8724,N_8324);
or U9092 (N_9092,N_8576,N_8181);
or U9093 (N_9093,N_8431,N_8235);
nor U9094 (N_9094,N_8600,N_8258);
or U9095 (N_9095,N_8727,N_8380);
xor U9096 (N_9096,N_8304,N_8477);
nor U9097 (N_9097,N_8531,N_8064);
nand U9098 (N_9098,N_8440,N_8527);
or U9099 (N_9099,N_8747,N_8347);
or U9100 (N_9100,N_8663,N_8240);
nor U9101 (N_9101,N_8145,N_8208);
and U9102 (N_9102,N_8519,N_8234);
nand U9103 (N_9103,N_8109,N_8577);
xnor U9104 (N_9104,N_8572,N_8096);
nor U9105 (N_9105,N_8218,N_8451);
and U9106 (N_9106,N_8723,N_8146);
nor U9107 (N_9107,N_8756,N_8151);
nand U9108 (N_9108,N_8139,N_8586);
nand U9109 (N_9109,N_8015,N_8237);
xnor U9110 (N_9110,N_8289,N_8110);
and U9111 (N_9111,N_8067,N_8253);
xor U9112 (N_9112,N_8194,N_8448);
nor U9113 (N_9113,N_8688,N_8591);
nand U9114 (N_9114,N_8489,N_8790);
xnor U9115 (N_9115,N_8447,N_8764);
and U9116 (N_9116,N_8487,N_8429);
nand U9117 (N_9117,N_8003,N_8026);
nor U9118 (N_9118,N_8741,N_8030);
or U9119 (N_9119,N_8341,N_8005);
and U9120 (N_9120,N_8295,N_8152);
and U9121 (N_9121,N_8689,N_8516);
xor U9122 (N_9122,N_8482,N_8631);
nor U9123 (N_9123,N_8693,N_8436);
xnor U9124 (N_9124,N_8777,N_8518);
and U9125 (N_9125,N_8729,N_8694);
xnor U9126 (N_9126,N_8618,N_8369);
or U9127 (N_9127,N_8746,N_8709);
nor U9128 (N_9128,N_8456,N_8565);
or U9129 (N_9129,N_8159,N_8432);
nor U9130 (N_9130,N_8395,N_8597);
and U9131 (N_9131,N_8769,N_8198);
and U9132 (N_9132,N_8386,N_8646);
xnor U9133 (N_9133,N_8427,N_8195);
nor U9134 (N_9134,N_8635,N_8403);
nor U9135 (N_9135,N_8523,N_8666);
and U9136 (N_9136,N_8675,N_8450);
nand U9137 (N_9137,N_8787,N_8192);
nand U9138 (N_9138,N_8263,N_8177);
and U9139 (N_9139,N_8361,N_8620);
nor U9140 (N_9140,N_8612,N_8095);
or U9141 (N_9141,N_8180,N_8782);
nand U9142 (N_9142,N_8297,N_8670);
xor U9143 (N_9143,N_8179,N_8484);
and U9144 (N_9144,N_8245,N_8298);
nand U9145 (N_9145,N_8108,N_8017);
xor U9146 (N_9146,N_8174,N_8778);
or U9147 (N_9147,N_8348,N_8390);
and U9148 (N_9148,N_8360,N_8392);
or U9149 (N_9149,N_8056,N_8765);
xor U9150 (N_9150,N_8557,N_8120);
nand U9151 (N_9151,N_8642,N_8583);
xor U9152 (N_9152,N_8083,N_8651);
nor U9153 (N_9153,N_8242,N_8733);
xor U9154 (N_9154,N_8686,N_8443);
nand U9155 (N_9155,N_8468,N_8040);
and U9156 (N_9156,N_8114,N_8654);
xnor U9157 (N_9157,N_8035,N_8759);
and U9158 (N_9158,N_8239,N_8305);
nor U9159 (N_9159,N_8085,N_8732);
nor U9160 (N_9160,N_8070,N_8103);
and U9161 (N_9161,N_8215,N_8130);
nor U9162 (N_9162,N_8563,N_8466);
xor U9163 (N_9163,N_8725,N_8334);
xnor U9164 (N_9164,N_8082,N_8697);
nor U9165 (N_9165,N_8217,N_8054);
or U9166 (N_9166,N_8252,N_8405);
xnor U9167 (N_9167,N_8761,N_8025);
nand U9168 (N_9168,N_8362,N_8175);
or U9169 (N_9169,N_8656,N_8209);
and U9170 (N_9170,N_8797,N_8673);
nand U9171 (N_9171,N_8411,N_8475);
nand U9172 (N_9172,N_8065,N_8555);
or U9173 (N_9173,N_8751,N_8226);
or U9174 (N_9174,N_8077,N_8292);
or U9175 (N_9175,N_8285,N_8624);
and U9176 (N_9176,N_8680,N_8485);
and U9177 (N_9177,N_8754,N_8737);
or U9178 (N_9178,N_8785,N_8402);
nand U9179 (N_9179,N_8200,N_8687);
xor U9180 (N_9180,N_8660,N_8043);
xnor U9181 (N_9181,N_8795,N_8696);
or U9182 (N_9182,N_8423,N_8526);
nor U9183 (N_9183,N_8491,N_8619);
or U9184 (N_9184,N_8063,N_8191);
or U9185 (N_9185,N_8532,N_8396);
nand U9186 (N_9186,N_8229,N_8093);
nand U9187 (N_9187,N_8424,N_8267);
nor U9188 (N_9188,N_8301,N_8288);
or U9189 (N_9189,N_8106,N_8662);
nor U9190 (N_9190,N_8133,N_8528);
and U9191 (N_9191,N_8099,N_8385);
nand U9192 (N_9192,N_8087,N_8617);
xnor U9193 (N_9193,N_8592,N_8339);
or U9194 (N_9194,N_8743,N_8704);
or U9195 (N_9195,N_8699,N_8739);
nand U9196 (N_9196,N_8302,N_8752);
xor U9197 (N_9197,N_8533,N_8314);
or U9198 (N_9198,N_8098,N_8548);
nor U9199 (N_9199,N_8105,N_8327);
nand U9200 (N_9200,N_8215,N_8035);
nand U9201 (N_9201,N_8196,N_8568);
nand U9202 (N_9202,N_8093,N_8127);
xor U9203 (N_9203,N_8191,N_8682);
nand U9204 (N_9204,N_8560,N_8081);
nand U9205 (N_9205,N_8529,N_8540);
nand U9206 (N_9206,N_8112,N_8639);
nor U9207 (N_9207,N_8456,N_8743);
or U9208 (N_9208,N_8399,N_8437);
nand U9209 (N_9209,N_8737,N_8411);
xor U9210 (N_9210,N_8339,N_8306);
or U9211 (N_9211,N_8493,N_8432);
or U9212 (N_9212,N_8069,N_8584);
or U9213 (N_9213,N_8351,N_8117);
or U9214 (N_9214,N_8272,N_8370);
or U9215 (N_9215,N_8040,N_8657);
and U9216 (N_9216,N_8279,N_8329);
nor U9217 (N_9217,N_8189,N_8114);
nor U9218 (N_9218,N_8303,N_8443);
or U9219 (N_9219,N_8099,N_8364);
nor U9220 (N_9220,N_8177,N_8535);
nand U9221 (N_9221,N_8003,N_8361);
nor U9222 (N_9222,N_8770,N_8505);
or U9223 (N_9223,N_8581,N_8345);
and U9224 (N_9224,N_8125,N_8245);
or U9225 (N_9225,N_8499,N_8032);
and U9226 (N_9226,N_8075,N_8026);
nor U9227 (N_9227,N_8260,N_8755);
and U9228 (N_9228,N_8658,N_8507);
nand U9229 (N_9229,N_8609,N_8555);
or U9230 (N_9230,N_8741,N_8387);
nand U9231 (N_9231,N_8620,N_8764);
and U9232 (N_9232,N_8557,N_8080);
and U9233 (N_9233,N_8621,N_8020);
or U9234 (N_9234,N_8466,N_8405);
nor U9235 (N_9235,N_8257,N_8408);
and U9236 (N_9236,N_8224,N_8580);
nor U9237 (N_9237,N_8026,N_8636);
or U9238 (N_9238,N_8064,N_8433);
or U9239 (N_9239,N_8046,N_8492);
and U9240 (N_9240,N_8348,N_8263);
or U9241 (N_9241,N_8245,N_8635);
nor U9242 (N_9242,N_8273,N_8384);
xor U9243 (N_9243,N_8253,N_8646);
xor U9244 (N_9244,N_8692,N_8589);
nand U9245 (N_9245,N_8324,N_8691);
and U9246 (N_9246,N_8541,N_8626);
nor U9247 (N_9247,N_8693,N_8555);
nand U9248 (N_9248,N_8557,N_8494);
xnor U9249 (N_9249,N_8614,N_8042);
and U9250 (N_9250,N_8603,N_8346);
or U9251 (N_9251,N_8523,N_8187);
nor U9252 (N_9252,N_8796,N_8191);
xor U9253 (N_9253,N_8278,N_8388);
or U9254 (N_9254,N_8064,N_8749);
nand U9255 (N_9255,N_8035,N_8136);
and U9256 (N_9256,N_8733,N_8750);
or U9257 (N_9257,N_8346,N_8705);
xnor U9258 (N_9258,N_8722,N_8699);
and U9259 (N_9259,N_8751,N_8457);
nor U9260 (N_9260,N_8273,N_8695);
xor U9261 (N_9261,N_8423,N_8686);
and U9262 (N_9262,N_8078,N_8765);
xnor U9263 (N_9263,N_8377,N_8166);
or U9264 (N_9264,N_8195,N_8739);
or U9265 (N_9265,N_8232,N_8120);
xor U9266 (N_9266,N_8483,N_8496);
nor U9267 (N_9267,N_8207,N_8464);
or U9268 (N_9268,N_8311,N_8248);
nor U9269 (N_9269,N_8588,N_8447);
nor U9270 (N_9270,N_8519,N_8719);
and U9271 (N_9271,N_8049,N_8174);
and U9272 (N_9272,N_8077,N_8105);
xor U9273 (N_9273,N_8707,N_8627);
nor U9274 (N_9274,N_8770,N_8111);
and U9275 (N_9275,N_8716,N_8083);
nor U9276 (N_9276,N_8462,N_8603);
xor U9277 (N_9277,N_8345,N_8644);
or U9278 (N_9278,N_8627,N_8697);
xnor U9279 (N_9279,N_8559,N_8156);
or U9280 (N_9280,N_8611,N_8525);
xnor U9281 (N_9281,N_8496,N_8215);
or U9282 (N_9282,N_8330,N_8173);
xor U9283 (N_9283,N_8510,N_8260);
nand U9284 (N_9284,N_8510,N_8180);
nand U9285 (N_9285,N_8729,N_8130);
xnor U9286 (N_9286,N_8540,N_8260);
and U9287 (N_9287,N_8232,N_8417);
and U9288 (N_9288,N_8337,N_8412);
nor U9289 (N_9289,N_8559,N_8741);
nand U9290 (N_9290,N_8130,N_8379);
and U9291 (N_9291,N_8405,N_8506);
and U9292 (N_9292,N_8532,N_8297);
nand U9293 (N_9293,N_8679,N_8006);
nand U9294 (N_9294,N_8247,N_8193);
and U9295 (N_9295,N_8349,N_8123);
and U9296 (N_9296,N_8289,N_8022);
or U9297 (N_9297,N_8116,N_8236);
nand U9298 (N_9298,N_8346,N_8450);
nor U9299 (N_9299,N_8715,N_8584);
nand U9300 (N_9300,N_8766,N_8134);
and U9301 (N_9301,N_8438,N_8390);
nor U9302 (N_9302,N_8114,N_8073);
and U9303 (N_9303,N_8198,N_8095);
or U9304 (N_9304,N_8544,N_8744);
nand U9305 (N_9305,N_8033,N_8150);
nand U9306 (N_9306,N_8438,N_8130);
xor U9307 (N_9307,N_8477,N_8320);
xnor U9308 (N_9308,N_8006,N_8793);
xnor U9309 (N_9309,N_8245,N_8628);
nand U9310 (N_9310,N_8191,N_8495);
xor U9311 (N_9311,N_8588,N_8018);
nand U9312 (N_9312,N_8074,N_8449);
or U9313 (N_9313,N_8509,N_8682);
nor U9314 (N_9314,N_8344,N_8584);
and U9315 (N_9315,N_8238,N_8115);
nand U9316 (N_9316,N_8555,N_8015);
nor U9317 (N_9317,N_8650,N_8430);
or U9318 (N_9318,N_8347,N_8133);
nor U9319 (N_9319,N_8284,N_8476);
xor U9320 (N_9320,N_8103,N_8771);
xnor U9321 (N_9321,N_8651,N_8146);
xnor U9322 (N_9322,N_8201,N_8624);
nor U9323 (N_9323,N_8128,N_8789);
nand U9324 (N_9324,N_8145,N_8780);
or U9325 (N_9325,N_8162,N_8582);
nor U9326 (N_9326,N_8587,N_8173);
nand U9327 (N_9327,N_8604,N_8140);
or U9328 (N_9328,N_8160,N_8539);
and U9329 (N_9329,N_8410,N_8640);
nor U9330 (N_9330,N_8716,N_8093);
nand U9331 (N_9331,N_8446,N_8755);
nand U9332 (N_9332,N_8622,N_8448);
and U9333 (N_9333,N_8589,N_8304);
and U9334 (N_9334,N_8584,N_8370);
or U9335 (N_9335,N_8022,N_8799);
or U9336 (N_9336,N_8322,N_8529);
and U9337 (N_9337,N_8750,N_8177);
or U9338 (N_9338,N_8552,N_8665);
xnor U9339 (N_9339,N_8489,N_8556);
or U9340 (N_9340,N_8686,N_8004);
nand U9341 (N_9341,N_8055,N_8283);
nor U9342 (N_9342,N_8663,N_8010);
and U9343 (N_9343,N_8511,N_8617);
nand U9344 (N_9344,N_8661,N_8709);
nor U9345 (N_9345,N_8304,N_8232);
or U9346 (N_9346,N_8204,N_8072);
or U9347 (N_9347,N_8521,N_8695);
nor U9348 (N_9348,N_8379,N_8275);
nand U9349 (N_9349,N_8588,N_8499);
xnor U9350 (N_9350,N_8278,N_8171);
nor U9351 (N_9351,N_8549,N_8367);
and U9352 (N_9352,N_8512,N_8127);
and U9353 (N_9353,N_8638,N_8385);
and U9354 (N_9354,N_8512,N_8363);
nand U9355 (N_9355,N_8536,N_8124);
nor U9356 (N_9356,N_8010,N_8245);
and U9357 (N_9357,N_8265,N_8070);
xnor U9358 (N_9358,N_8488,N_8219);
nand U9359 (N_9359,N_8745,N_8132);
xor U9360 (N_9360,N_8608,N_8566);
and U9361 (N_9361,N_8670,N_8746);
nand U9362 (N_9362,N_8177,N_8543);
or U9363 (N_9363,N_8476,N_8283);
nand U9364 (N_9364,N_8656,N_8182);
or U9365 (N_9365,N_8304,N_8250);
nand U9366 (N_9366,N_8622,N_8071);
nor U9367 (N_9367,N_8582,N_8670);
or U9368 (N_9368,N_8352,N_8550);
nand U9369 (N_9369,N_8017,N_8547);
nand U9370 (N_9370,N_8467,N_8158);
nand U9371 (N_9371,N_8609,N_8533);
xnor U9372 (N_9372,N_8679,N_8515);
xnor U9373 (N_9373,N_8432,N_8652);
xor U9374 (N_9374,N_8160,N_8380);
nor U9375 (N_9375,N_8030,N_8628);
and U9376 (N_9376,N_8439,N_8586);
nor U9377 (N_9377,N_8665,N_8408);
xor U9378 (N_9378,N_8087,N_8104);
or U9379 (N_9379,N_8483,N_8078);
or U9380 (N_9380,N_8479,N_8560);
nor U9381 (N_9381,N_8219,N_8530);
nand U9382 (N_9382,N_8260,N_8119);
xor U9383 (N_9383,N_8696,N_8361);
and U9384 (N_9384,N_8348,N_8088);
and U9385 (N_9385,N_8047,N_8535);
nand U9386 (N_9386,N_8397,N_8654);
xor U9387 (N_9387,N_8491,N_8627);
xnor U9388 (N_9388,N_8753,N_8187);
and U9389 (N_9389,N_8416,N_8519);
and U9390 (N_9390,N_8333,N_8246);
or U9391 (N_9391,N_8244,N_8631);
xor U9392 (N_9392,N_8389,N_8720);
nand U9393 (N_9393,N_8770,N_8351);
and U9394 (N_9394,N_8619,N_8288);
xor U9395 (N_9395,N_8119,N_8188);
nand U9396 (N_9396,N_8739,N_8728);
nand U9397 (N_9397,N_8433,N_8582);
nor U9398 (N_9398,N_8190,N_8709);
nor U9399 (N_9399,N_8293,N_8170);
xor U9400 (N_9400,N_8139,N_8399);
xor U9401 (N_9401,N_8060,N_8207);
nand U9402 (N_9402,N_8377,N_8152);
nand U9403 (N_9403,N_8427,N_8334);
or U9404 (N_9404,N_8306,N_8296);
or U9405 (N_9405,N_8381,N_8032);
or U9406 (N_9406,N_8791,N_8001);
and U9407 (N_9407,N_8657,N_8112);
nand U9408 (N_9408,N_8784,N_8433);
xnor U9409 (N_9409,N_8359,N_8417);
nand U9410 (N_9410,N_8104,N_8695);
nand U9411 (N_9411,N_8585,N_8730);
nor U9412 (N_9412,N_8414,N_8220);
nand U9413 (N_9413,N_8025,N_8600);
and U9414 (N_9414,N_8081,N_8131);
xor U9415 (N_9415,N_8598,N_8220);
xor U9416 (N_9416,N_8087,N_8253);
xor U9417 (N_9417,N_8384,N_8527);
or U9418 (N_9418,N_8704,N_8269);
nand U9419 (N_9419,N_8413,N_8500);
or U9420 (N_9420,N_8374,N_8025);
nand U9421 (N_9421,N_8679,N_8339);
nor U9422 (N_9422,N_8149,N_8771);
nor U9423 (N_9423,N_8068,N_8595);
or U9424 (N_9424,N_8129,N_8664);
nor U9425 (N_9425,N_8175,N_8476);
and U9426 (N_9426,N_8659,N_8386);
or U9427 (N_9427,N_8538,N_8456);
nor U9428 (N_9428,N_8723,N_8324);
xor U9429 (N_9429,N_8346,N_8696);
or U9430 (N_9430,N_8322,N_8688);
nand U9431 (N_9431,N_8710,N_8727);
nor U9432 (N_9432,N_8036,N_8006);
and U9433 (N_9433,N_8262,N_8770);
and U9434 (N_9434,N_8330,N_8680);
nor U9435 (N_9435,N_8235,N_8522);
or U9436 (N_9436,N_8609,N_8769);
or U9437 (N_9437,N_8452,N_8380);
and U9438 (N_9438,N_8629,N_8667);
nor U9439 (N_9439,N_8186,N_8027);
xnor U9440 (N_9440,N_8443,N_8487);
xnor U9441 (N_9441,N_8754,N_8658);
and U9442 (N_9442,N_8224,N_8025);
nor U9443 (N_9443,N_8041,N_8229);
nor U9444 (N_9444,N_8097,N_8701);
xor U9445 (N_9445,N_8340,N_8305);
or U9446 (N_9446,N_8749,N_8202);
or U9447 (N_9447,N_8233,N_8056);
xnor U9448 (N_9448,N_8720,N_8360);
or U9449 (N_9449,N_8710,N_8389);
and U9450 (N_9450,N_8398,N_8518);
and U9451 (N_9451,N_8336,N_8385);
nor U9452 (N_9452,N_8610,N_8030);
nor U9453 (N_9453,N_8276,N_8705);
nor U9454 (N_9454,N_8288,N_8249);
nor U9455 (N_9455,N_8774,N_8005);
xnor U9456 (N_9456,N_8660,N_8284);
nand U9457 (N_9457,N_8760,N_8665);
xnor U9458 (N_9458,N_8343,N_8498);
nand U9459 (N_9459,N_8310,N_8211);
and U9460 (N_9460,N_8631,N_8562);
and U9461 (N_9461,N_8038,N_8092);
xnor U9462 (N_9462,N_8643,N_8064);
nand U9463 (N_9463,N_8514,N_8782);
nor U9464 (N_9464,N_8003,N_8024);
xor U9465 (N_9465,N_8296,N_8290);
nand U9466 (N_9466,N_8372,N_8782);
or U9467 (N_9467,N_8267,N_8771);
nand U9468 (N_9468,N_8303,N_8257);
and U9469 (N_9469,N_8714,N_8751);
or U9470 (N_9470,N_8610,N_8395);
nand U9471 (N_9471,N_8733,N_8292);
nand U9472 (N_9472,N_8445,N_8323);
and U9473 (N_9473,N_8186,N_8688);
and U9474 (N_9474,N_8733,N_8196);
and U9475 (N_9475,N_8209,N_8470);
nand U9476 (N_9476,N_8498,N_8313);
nand U9477 (N_9477,N_8205,N_8698);
and U9478 (N_9478,N_8538,N_8622);
or U9479 (N_9479,N_8065,N_8507);
nor U9480 (N_9480,N_8789,N_8028);
and U9481 (N_9481,N_8130,N_8577);
or U9482 (N_9482,N_8488,N_8511);
nor U9483 (N_9483,N_8627,N_8308);
nand U9484 (N_9484,N_8626,N_8246);
nand U9485 (N_9485,N_8516,N_8791);
xnor U9486 (N_9486,N_8574,N_8367);
nor U9487 (N_9487,N_8733,N_8780);
and U9488 (N_9488,N_8447,N_8048);
nor U9489 (N_9489,N_8724,N_8154);
xor U9490 (N_9490,N_8074,N_8409);
nor U9491 (N_9491,N_8226,N_8231);
and U9492 (N_9492,N_8578,N_8078);
nand U9493 (N_9493,N_8674,N_8223);
nand U9494 (N_9494,N_8691,N_8353);
xor U9495 (N_9495,N_8792,N_8043);
nand U9496 (N_9496,N_8742,N_8037);
xor U9497 (N_9497,N_8492,N_8266);
nand U9498 (N_9498,N_8244,N_8531);
nand U9499 (N_9499,N_8257,N_8712);
or U9500 (N_9500,N_8281,N_8636);
xnor U9501 (N_9501,N_8140,N_8341);
or U9502 (N_9502,N_8633,N_8642);
xor U9503 (N_9503,N_8311,N_8662);
nor U9504 (N_9504,N_8655,N_8332);
or U9505 (N_9505,N_8320,N_8687);
xnor U9506 (N_9506,N_8465,N_8300);
nand U9507 (N_9507,N_8692,N_8001);
xnor U9508 (N_9508,N_8239,N_8601);
or U9509 (N_9509,N_8125,N_8694);
nand U9510 (N_9510,N_8496,N_8628);
nor U9511 (N_9511,N_8530,N_8595);
or U9512 (N_9512,N_8704,N_8164);
or U9513 (N_9513,N_8782,N_8625);
or U9514 (N_9514,N_8213,N_8526);
nor U9515 (N_9515,N_8704,N_8426);
nor U9516 (N_9516,N_8378,N_8405);
nor U9517 (N_9517,N_8187,N_8255);
nor U9518 (N_9518,N_8638,N_8607);
xor U9519 (N_9519,N_8354,N_8621);
xor U9520 (N_9520,N_8565,N_8745);
nor U9521 (N_9521,N_8082,N_8706);
and U9522 (N_9522,N_8191,N_8565);
and U9523 (N_9523,N_8792,N_8308);
or U9524 (N_9524,N_8495,N_8180);
or U9525 (N_9525,N_8692,N_8198);
nor U9526 (N_9526,N_8077,N_8177);
xor U9527 (N_9527,N_8048,N_8409);
and U9528 (N_9528,N_8029,N_8307);
or U9529 (N_9529,N_8387,N_8092);
and U9530 (N_9530,N_8113,N_8616);
nand U9531 (N_9531,N_8007,N_8270);
nand U9532 (N_9532,N_8456,N_8188);
nand U9533 (N_9533,N_8676,N_8531);
nor U9534 (N_9534,N_8793,N_8141);
nor U9535 (N_9535,N_8672,N_8076);
nand U9536 (N_9536,N_8649,N_8641);
or U9537 (N_9537,N_8583,N_8276);
or U9538 (N_9538,N_8199,N_8255);
nand U9539 (N_9539,N_8498,N_8374);
xnor U9540 (N_9540,N_8456,N_8340);
xnor U9541 (N_9541,N_8084,N_8108);
xor U9542 (N_9542,N_8708,N_8697);
and U9543 (N_9543,N_8373,N_8512);
nand U9544 (N_9544,N_8180,N_8040);
and U9545 (N_9545,N_8783,N_8297);
xnor U9546 (N_9546,N_8587,N_8392);
or U9547 (N_9547,N_8722,N_8451);
xnor U9548 (N_9548,N_8575,N_8419);
nor U9549 (N_9549,N_8708,N_8431);
nor U9550 (N_9550,N_8165,N_8726);
nand U9551 (N_9551,N_8791,N_8773);
xor U9552 (N_9552,N_8075,N_8148);
xor U9553 (N_9553,N_8534,N_8755);
nand U9554 (N_9554,N_8719,N_8155);
nor U9555 (N_9555,N_8029,N_8559);
xor U9556 (N_9556,N_8751,N_8600);
and U9557 (N_9557,N_8543,N_8161);
or U9558 (N_9558,N_8108,N_8501);
and U9559 (N_9559,N_8205,N_8797);
or U9560 (N_9560,N_8420,N_8206);
nor U9561 (N_9561,N_8297,N_8771);
xor U9562 (N_9562,N_8442,N_8641);
nor U9563 (N_9563,N_8483,N_8586);
xnor U9564 (N_9564,N_8465,N_8755);
xnor U9565 (N_9565,N_8073,N_8400);
nand U9566 (N_9566,N_8271,N_8068);
xor U9567 (N_9567,N_8061,N_8490);
nand U9568 (N_9568,N_8593,N_8284);
or U9569 (N_9569,N_8217,N_8009);
xor U9570 (N_9570,N_8425,N_8445);
or U9571 (N_9571,N_8117,N_8216);
xnor U9572 (N_9572,N_8218,N_8399);
and U9573 (N_9573,N_8748,N_8528);
xor U9574 (N_9574,N_8224,N_8661);
nand U9575 (N_9575,N_8198,N_8144);
and U9576 (N_9576,N_8057,N_8625);
nor U9577 (N_9577,N_8180,N_8322);
and U9578 (N_9578,N_8380,N_8487);
nand U9579 (N_9579,N_8258,N_8702);
xnor U9580 (N_9580,N_8793,N_8122);
xor U9581 (N_9581,N_8376,N_8259);
and U9582 (N_9582,N_8019,N_8619);
or U9583 (N_9583,N_8436,N_8110);
nand U9584 (N_9584,N_8032,N_8379);
nand U9585 (N_9585,N_8669,N_8587);
and U9586 (N_9586,N_8177,N_8585);
xnor U9587 (N_9587,N_8360,N_8319);
xor U9588 (N_9588,N_8693,N_8413);
and U9589 (N_9589,N_8790,N_8636);
nor U9590 (N_9590,N_8725,N_8018);
and U9591 (N_9591,N_8686,N_8717);
and U9592 (N_9592,N_8199,N_8261);
nor U9593 (N_9593,N_8579,N_8590);
nand U9594 (N_9594,N_8718,N_8106);
nand U9595 (N_9595,N_8703,N_8132);
or U9596 (N_9596,N_8212,N_8245);
xor U9597 (N_9597,N_8183,N_8776);
or U9598 (N_9598,N_8448,N_8452);
nor U9599 (N_9599,N_8640,N_8066);
xor U9600 (N_9600,N_9020,N_9253);
xnor U9601 (N_9601,N_9372,N_8822);
or U9602 (N_9602,N_8951,N_8808);
or U9603 (N_9603,N_9562,N_9458);
xnor U9604 (N_9604,N_9016,N_9051);
nand U9605 (N_9605,N_9482,N_9468);
or U9606 (N_9606,N_9577,N_9362);
and U9607 (N_9607,N_9420,N_9315);
and U9608 (N_9608,N_9058,N_8872);
nand U9609 (N_9609,N_9258,N_9265);
nor U9610 (N_9610,N_8984,N_8848);
and U9611 (N_9611,N_9392,N_9040);
nand U9612 (N_9612,N_9262,N_9480);
or U9613 (N_9613,N_8871,N_9557);
xnor U9614 (N_9614,N_9101,N_8932);
nand U9615 (N_9615,N_9459,N_8859);
xnor U9616 (N_9616,N_9305,N_9214);
xnor U9617 (N_9617,N_9565,N_9072);
xnor U9618 (N_9618,N_9310,N_9318);
xor U9619 (N_9619,N_9014,N_8837);
and U9620 (N_9620,N_9224,N_9124);
xnor U9621 (N_9621,N_8854,N_9117);
or U9622 (N_9622,N_9580,N_9371);
or U9623 (N_9623,N_9090,N_8802);
and U9624 (N_9624,N_9015,N_8858);
nand U9625 (N_9625,N_9191,N_9381);
nand U9626 (N_9626,N_9170,N_9230);
xnor U9627 (N_9627,N_9326,N_8911);
or U9628 (N_9628,N_8825,N_9240);
or U9629 (N_9629,N_9122,N_9129);
and U9630 (N_9630,N_9142,N_8976);
and U9631 (N_9631,N_8960,N_9281);
or U9632 (N_9632,N_8957,N_9350);
nor U9633 (N_9633,N_9246,N_9188);
nor U9634 (N_9634,N_9138,N_9073);
nand U9635 (N_9635,N_9467,N_9297);
or U9636 (N_9636,N_9210,N_9386);
and U9637 (N_9637,N_8935,N_9450);
and U9638 (N_9638,N_8912,N_9424);
xnor U9639 (N_9639,N_8917,N_9303);
nor U9640 (N_9640,N_9596,N_8986);
xor U9641 (N_9641,N_8941,N_9257);
xor U9642 (N_9642,N_9550,N_9233);
or U9643 (N_9643,N_9013,N_8929);
or U9644 (N_9644,N_8933,N_8982);
nor U9645 (N_9645,N_8916,N_9135);
nand U9646 (N_9646,N_9248,N_8988);
nor U9647 (N_9647,N_9235,N_8809);
nand U9648 (N_9648,N_9416,N_9093);
and U9649 (N_9649,N_9516,N_9493);
nand U9650 (N_9650,N_8923,N_9053);
nand U9651 (N_9651,N_9439,N_9437);
nor U9652 (N_9652,N_9389,N_9156);
and U9653 (N_9653,N_9334,N_9454);
xor U9654 (N_9654,N_8819,N_9376);
and U9655 (N_9655,N_9077,N_8828);
xnor U9656 (N_9656,N_8868,N_9464);
nand U9657 (N_9657,N_9197,N_9509);
nor U9658 (N_9658,N_9027,N_9506);
and U9659 (N_9659,N_9106,N_9299);
or U9660 (N_9660,N_9128,N_8910);
nand U9661 (N_9661,N_9430,N_8826);
and U9662 (N_9662,N_9229,N_9037);
and U9663 (N_9663,N_9290,N_9428);
nor U9664 (N_9664,N_9431,N_9032);
and U9665 (N_9665,N_9126,N_8861);
nor U9666 (N_9666,N_9116,N_9460);
nand U9667 (N_9667,N_9449,N_9242);
or U9668 (N_9668,N_9354,N_9019);
or U9669 (N_9669,N_9064,N_9086);
and U9670 (N_9670,N_8952,N_8849);
and U9671 (N_9671,N_9418,N_9532);
nand U9672 (N_9672,N_8823,N_9484);
and U9673 (N_9673,N_9330,N_9107);
or U9674 (N_9674,N_9538,N_8877);
nand U9675 (N_9675,N_9184,N_9183);
nor U9676 (N_9676,N_9161,N_8840);
xor U9677 (N_9677,N_9042,N_9465);
nand U9678 (N_9678,N_9164,N_9554);
xor U9679 (N_9679,N_9024,N_9226);
xor U9680 (N_9680,N_8895,N_9074);
and U9681 (N_9681,N_9114,N_9581);
and U9682 (N_9682,N_8959,N_9123);
and U9683 (N_9683,N_9515,N_9045);
xor U9684 (N_9684,N_9499,N_9010);
and U9685 (N_9685,N_8817,N_9451);
or U9686 (N_9686,N_8814,N_8853);
xor U9687 (N_9687,N_9218,N_9034);
xor U9688 (N_9688,N_9345,N_9343);
or U9689 (N_9689,N_9154,N_9171);
xnor U9690 (N_9690,N_9455,N_9541);
nand U9691 (N_9691,N_9466,N_9425);
and U9692 (N_9692,N_9213,N_8972);
xnor U9693 (N_9693,N_8964,N_9215);
nor U9694 (N_9694,N_8989,N_9582);
nand U9695 (N_9695,N_9593,N_9001);
or U9696 (N_9696,N_9203,N_9059);
nor U9697 (N_9697,N_9545,N_9169);
or U9698 (N_9698,N_8914,N_9496);
nand U9699 (N_9699,N_9505,N_9176);
nand U9700 (N_9700,N_9308,N_9339);
nand U9701 (N_9701,N_8801,N_8812);
xor U9702 (N_9702,N_9275,N_9195);
or U9703 (N_9703,N_8865,N_8950);
nor U9704 (N_9704,N_8894,N_9384);
or U9705 (N_9705,N_8886,N_9180);
xnor U9706 (N_9706,N_9368,N_9237);
or U9707 (N_9707,N_9473,N_9595);
or U9708 (N_9708,N_9586,N_9205);
xor U9709 (N_9709,N_8897,N_9251);
xnor U9710 (N_9710,N_9139,N_9470);
nand U9711 (N_9711,N_9304,N_8852);
and U9712 (N_9712,N_9151,N_8995);
nand U9713 (N_9713,N_9267,N_9320);
or U9714 (N_9714,N_9574,N_9311);
nor U9715 (N_9715,N_9048,N_9560);
xnor U9716 (N_9716,N_9099,N_9131);
and U9717 (N_9717,N_8906,N_9510);
nand U9718 (N_9718,N_9571,N_9527);
or U9719 (N_9719,N_9052,N_9018);
and U9720 (N_9720,N_9283,N_9471);
nand U9721 (N_9721,N_8813,N_9266);
xor U9722 (N_9722,N_9388,N_8842);
and U9723 (N_9723,N_9137,N_9273);
and U9724 (N_9724,N_8921,N_9274);
xnor U9725 (N_9725,N_9022,N_8881);
and U9726 (N_9726,N_8947,N_8985);
nor U9727 (N_9727,N_8882,N_9033);
nand U9728 (N_9728,N_9462,N_9095);
and U9729 (N_9729,N_9271,N_9380);
nor U9730 (N_9730,N_9427,N_9331);
nand U9731 (N_9731,N_9066,N_9199);
or U9732 (N_9732,N_9278,N_8806);
xor U9733 (N_9733,N_9227,N_9313);
or U9734 (N_9734,N_9092,N_8832);
and U9735 (N_9735,N_9397,N_9316);
nor U9736 (N_9736,N_8829,N_9245);
or U9737 (N_9737,N_9133,N_9168);
and U9738 (N_9738,N_9485,N_9357);
and U9739 (N_9739,N_8997,N_9497);
nor U9740 (N_9740,N_8948,N_8870);
or U9741 (N_9741,N_9435,N_9411);
nor U9742 (N_9742,N_9136,N_8836);
or U9743 (N_9743,N_8949,N_9481);
or U9744 (N_9744,N_9363,N_9157);
nand U9745 (N_9745,N_9494,N_8909);
or U9746 (N_9746,N_9085,N_8994);
nand U9747 (N_9747,N_8876,N_9517);
xnor U9748 (N_9748,N_8908,N_8831);
or U9749 (N_9749,N_9190,N_9108);
and U9750 (N_9750,N_9535,N_8922);
and U9751 (N_9751,N_9125,N_9070);
xor U9752 (N_9752,N_8913,N_8851);
nand U9753 (N_9753,N_9563,N_9280);
or U9754 (N_9754,N_9332,N_9370);
nand U9755 (N_9755,N_8901,N_9444);
xnor U9756 (N_9756,N_9597,N_8804);
nand U9757 (N_9757,N_8953,N_9206);
nand U9758 (N_9758,N_8863,N_9091);
or U9759 (N_9759,N_9236,N_8888);
xnor U9760 (N_9760,N_8937,N_9585);
or U9761 (N_9761,N_9201,N_9118);
xnor U9762 (N_9762,N_8887,N_9256);
and U9763 (N_9763,N_8946,N_9115);
nand U9764 (N_9764,N_9508,N_9094);
xor U9765 (N_9765,N_9490,N_9504);
nand U9766 (N_9766,N_9495,N_9004);
nor U9767 (N_9767,N_9378,N_9202);
nor U9768 (N_9768,N_9222,N_9026);
or U9769 (N_9769,N_8938,N_9269);
nor U9770 (N_9770,N_8838,N_8983);
and U9771 (N_9771,N_9579,N_8968);
xnor U9772 (N_9772,N_9187,N_9573);
nand U9773 (N_9773,N_8915,N_9158);
nor U9774 (N_9774,N_9452,N_9570);
and U9775 (N_9775,N_9009,N_9539);
nand U9776 (N_9776,N_8878,N_9288);
nand U9777 (N_9777,N_9153,N_8925);
xor U9778 (N_9778,N_8843,N_9312);
xor U9779 (N_9779,N_9347,N_9395);
nand U9780 (N_9780,N_8945,N_8818);
nand U9781 (N_9781,N_9342,N_9322);
or U9782 (N_9782,N_9044,N_8860);
and U9783 (N_9783,N_9429,N_9300);
xor U9784 (N_9784,N_9279,N_8991);
nor U9785 (N_9785,N_9383,N_9012);
nand U9786 (N_9786,N_9542,N_8956);
xnor U9787 (N_9787,N_8926,N_8816);
xnor U9788 (N_9788,N_9338,N_8980);
xnor U9789 (N_9789,N_9432,N_9250);
nor U9790 (N_9790,N_9548,N_9518);
nor U9791 (N_9791,N_8979,N_9488);
or U9792 (N_9792,N_9247,N_9522);
nand U9793 (N_9793,N_8967,N_8800);
nor U9794 (N_9794,N_9479,N_8898);
nor U9795 (N_9795,N_9438,N_9160);
and U9796 (N_9796,N_9405,N_9097);
xnor U9797 (N_9797,N_9056,N_9287);
nand U9798 (N_9798,N_9302,N_9145);
nand U9799 (N_9799,N_9592,N_8999);
nand U9800 (N_9800,N_9575,N_9307);
nor U9801 (N_9801,N_9194,N_9196);
nand U9802 (N_9802,N_9149,N_9422);
or U9803 (N_9803,N_9492,N_9078);
nand U9804 (N_9804,N_8805,N_9512);
xor U9805 (N_9805,N_9477,N_8884);
xnor U9806 (N_9806,N_8807,N_9369);
xor U9807 (N_9807,N_9192,N_9546);
or U9808 (N_9808,N_9294,N_9351);
or U9809 (N_9809,N_8830,N_9333);
nand U9810 (N_9810,N_8811,N_9127);
and U9811 (N_9811,N_9584,N_8835);
xor U9812 (N_9812,N_9263,N_9447);
nor U9813 (N_9813,N_9501,N_9232);
nand U9814 (N_9814,N_8875,N_9231);
or U9815 (N_9815,N_8833,N_8918);
or U9816 (N_9816,N_9292,N_9075);
xor U9817 (N_9817,N_9441,N_9039);
nand U9818 (N_9818,N_9513,N_9065);
nand U9819 (N_9819,N_9021,N_9219);
nand U9820 (N_9820,N_8847,N_9293);
nor U9821 (N_9821,N_9005,N_9317);
and U9822 (N_9822,N_9148,N_9319);
or U9823 (N_9823,N_9017,N_9377);
xnor U9824 (N_9824,N_9289,N_9426);
or U9825 (N_9825,N_9068,N_9175);
and U9826 (N_9826,N_9419,N_9352);
nor U9827 (N_9827,N_9109,N_9489);
nand U9828 (N_9828,N_8815,N_9047);
and U9829 (N_9829,N_9212,N_9211);
xnor U9830 (N_9830,N_8857,N_9209);
and U9831 (N_9831,N_9143,N_9483);
xnor U9832 (N_9832,N_8867,N_9547);
nor U9833 (N_9833,N_9113,N_8885);
or U9834 (N_9834,N_8866,N_9448);
or U9835 (N_9835,N_9344,N_9134);
xnor U9836 (N_9836,N_8880,N_9050);
and U9837 (N_9837,N_9152,N_9568);
and U9838 (N_9838,N_8970,N_9514);
xnor U9839 (N_9839,N_8993,N_9216);
or U9840 (N_9840,N_8977,N_9238);
nand U9841 (N_9841,N_9337,N_9401);
and U9842 (N_9842,N_9220,N_9472);
and U9843 (N_9843,N_9088,N_9119);
xnor U9844 (N_9844,N_8850,N_9567);
nand U9845 (N_9845,N_9261,N_8969);
nor U9846 (N_9846,N_8834,N_9404);
or U9847 (N_9847,N_9564,N_9103);
nand U9848 (N_9848,N_9561,N_9069);
or U9849 (N_9849,N_9067,N_9270);
nand U9850 (N_9850,N_9373,N_8966);
and U9851 (N_9851,N_9486,N_9414);
nor U9852 (N_9852,N_9100,N_9081);
nor U9853 (N_9853,N_8905,N_8973);
xnor U9854 (N_9854,N_9355,N_9141);
or U9855 (N_9855,N_8891,N_8862);
nand U9856 (N_9856,N_9207,N_9208);
and U9857 (N_9857,N_9146,N_9559);
and U9858 (N_9858,N_9162,N_9399);
or U9859 (N_9859,N_9589,N_9463);
or U9860 (N_9860,N_9433,N_8869);
nor U9861 (N_9861,N_9023,N_8899);
nor U9862 (N_9862,N_9140,N_9543);
or U9863 (N_9863,N_9277,N_9445);
and U9864 (N_9864,N_8855,N_8824);
nor U9865 (N_9865,N_9374,N_8931);
nor U9866 (N_9866,N_9500,N_9572);
or U9867 (N_9867,N_8902,N_9003);
nor U9868 (N_9868,N_9461,N_9551);
or U9869 (N_9869,N_9007,N_9569);
xnor U9870 (N_9870,N_9361,N_9410);
or U9871 (N_9871,N_9159,N_9181);
nor U9872 (N_9872,N_9254,N_9268);
xnor U9873 (N_9873,N_9442,N_9259);
or U9874 (N_9874,N_9225,N_9144);
and U9875 (N_9875,N_8879,N_9549);
xor U9876 (N_9876,N_9276,N_9112);
xnor U9877 (N_9877,N_8873,N_8920);
and U9878 (N_9878,N_9587,N_9540);
and U9879 (N_9879,N_9029,N_9298);
xor U9880 (N_9880,N_9120,N_9286);
nand U9881 (N_9881,N_9417,N_8971);
or U9882 (N_9882,N_8827,N_8924);
nor U9883 (N_9883,N_9498,N_9002);
nand U9884 (N_9884,N_8845,N_9177);
nor U9885 (N_9885,N_9321,N_8928);
nor U9886 (N_9886,N_9375,N_9163);
or U9887 (N_9887,N_8944,N_9366);
xnor U9888 (N_9888,N_9228,N_9264);
nand U9889 (N_9889,N_9360,N_9193);
xnor U9890 (N_9890,N_9533,N_9475);
nor U9891 (N_9891,N_9525,N_8820);
and U9892 (N_9892,N_9000,N_9174);
nor U9893 (N_9893,N_9327,N_9284);
or U9894 (N_9894,N_8856,N_9111);
nor U9895 (N_9895,N_9036,N_9243);
and U9896 (N_9896,N_9409,N_8987);
or U9897 (N_9897,N_9359,N_9178);
nor U9898 (N_9898,N_8890,N_9110);
nor U9899 (N_9899,N_9349,N_9132);
and U9900 (N_9900,N_9049,N_8936);
nand U9901 (N_9901,N_9030,N_8907);
and U9902 (N_9902,N_9150,N_9011);
and U9903 (N_9903,N_8900,N_8961);
nand U9904 (N_9904,N_9348,N_9387);
and U9905 (N_9905,N_8940,N_9503);
nand U9906 (N_9906,N_9198,N_9167);
nand U9907 (N_9907,N_9221,N_9172);
or U9908 (N_9908,N_9469,N_9061);
and U9909 (N_9909,N_9446,N_9043);
nand U9910 (N_9910,N_8975,N_8963);
and U9911 (N_9911,N_8803,N_9336);
nand U9912 (N_9912,N_9364,N_9255);
and U9913 (N_9913,N_9555,N_9083);
nand U9914 (N_9914,N_9415,N_9412);
and U9915 (N_9915,N_8954,N_9309);
and U9916 (N_9916,N_9189,N_9335);
nor U9917 (N_9917,N_9407,N_9314);
and U9918 (N_9918,N_9536,N_9179);
nor U9919 (N_9919,N_9204,N_9402);
nor U9920 (N_9920,N_9365,N_8839);
and U9921 (N_9921,N_9423,N_9474);
nor U9922 (N_9922,N_9080,N_9063);
or U9923 (N_9923,N_9076,N_9391);
nor U9924 (N_9924,N_9301,N_9394);
and U9925 (N_9925,N_9436,N_9591);
and U9926 (N_9926,N_8996,N_8998);
nand U9927 (N_9927,N_9102,N_9147);
nand U9928 (N_9928,N_9296,N_9006);
nor U9929 (N_9929,N_9367,N_9491);
and U9930 (N_9930,N_9524,N_9537);
xor U9931 (N_9931,N_9443,N_9382);
nor U9932 (N_9932,N_9165,N_9028);
or U9933 (N_9933,N_8958,N_9576);
and U9934 (N_9934,N_9249,N_9223);
nor U9935 (N_9935,N_9379,N_9285);
or U9936 (N_9936,N_9239,N_9252);
or U9937 (N_9937,N_9599,N_8934);
nor U9938 (N_9938,N_9104,N_9185);
and U9939 (N_9939,N_9558,N_9528);
nor U9940 (N_9940,N_9393,N_9583);
or U9941 (N_9941,N_9340,N_9507);
nand U9942 (N_9942,N_9217,N_8974);
and U9943 (N_9943,N_8919,N_9130);
or U9944 (N_9944,N_9588,N_9105);
or U9945 (N_9945,N_9046,N_9556);
nor U9946 (N_9946,N_9598,N_9478);
or U9947 (N_9947,N_9244,N_8889);
xor U9948 (N_9948,N_9329,N_9356);
xor U9949 (N_9949,N_9055,N_9089);
and U9950 (N_9950,N_9084,N_9390);
nor U9951 (N_9951,N_9529,N_9358);
and U9952 (N_9952,N_9173,N_8903);
nand U9953 (N_9953,N_9457,N_9291);
nor U9954 (N_9954,N_8927,N_9421);
nand U9955 (N_9955,N_8978,N_9413);
xnor U9956 (N_9956,N_9054,N_9008);
and U9957 (N_9957,N_9511,N_8990);
and U9958 (N_9958,N_8962,N_8939);
and U9959 (N_9959,N_9062,N_9526);
and U9960 (N_9960,N_9098,N_9323);
xor U9961 (N_9961,N_9594,N_9341);
xor U9962 (N_9962,N_9346,N_8844);
and U9963 (N_9963,N_9031,N_9530);
or U9964 (N_9964,N_9096,N_8893);
nor U9965 (N_9965,N_9400,N_9403);
or U9966 (N_9966,N_9398,N_8955);
nand U9967 (N_9967,N_9234,N_8930);
or U9968 (N_9968,N_9534,N_9523);
or U9969 (N_9969,N_9324,N_9272);
nand U9970 (N_9970,N_9182,N_8864);
or U9971 (N_9971,N_9406,N_9487);
xor U9972 (N_9972,N_9440,N_8943);
and U9973 (N_9973,N_9456,N_9166);
nand U9974 (N_9974,N_9035,N_9295);
xor U9975 (N_9975,N_9434,N_9079);
nor U9976 (N_9976,N_8992,N_9396);
xnor U9977 (N_9977,N_9502,N_9325);
or U9978 (N_9978,N_9578,N_9566);
nor U9979 (N_9979,N_9200,N_8841);
nor U9980 (N_9980,N_9544,N_9041);
nor U9981 (N_9981,N_9328,N_9260);
nor U9982 (N_9982,N_9552,N_8810);
and U9983 (N_9983,N_8965,N_9155);
and U9984 (N_9984,N_9186,N_9385);
or U9985 (N_9985,N_8896,N_9353);
xor U9986 (N_9986,N_9531,N_9071);
nand U9987 (N_9987,N_9121,N_8892);
nor U9988 (N_9988,N_9306,N_8821);
xnor U9989 (N_9989,N_9553,N_8846);
nor U9990 (N_9990,N_8942,N_8981);
nand U9991 (N_9991,N_9060,N_8904);
and U9992 (N_9992,N_9082,N_8874);
nor U9993 (N_9993,N_9282,N_9453);
xnor U9994 (N_9994,N_9590,N_9476);
nor U9995 (N_9995,N_9408,N_9241);
nand U9996 (N_9996,N_9057,N_8883);
xnor U9997 (N_9997,N_9521,N_9520);
and U9998 (N_9998,N_9519,N_9038);
nand U9999 (N_9999,N_9025,N_9087);
xor U10000 (N_10000,N_9078,N_9243);
nand U10001 (N_10001,N_9582,N_8812);
and U10002 (N_10002,N_8958,N_9237);
or U10003 (N_10003,N_9266,N_9294);
nor U10004 (N_10004,N_9224,N_9130);
or U10005 (N_10005,N_8974,N_9477);
and U10006 (N_10006,N_9416,N_9004);
nor U10007 (N_10007,N_9288,N_9223);
or U10008 (N_10008,N_8974,N_9476);
nor U10009 (N_10009,N_9147,N_8881);
nor U10010 (N_10010,N_8825,N_9018);
xnor U10011 (N_10011,N_9095,N_8820);
or U10012 (N_10012,N_9319,N_8948);
xor U10013 (N_10013,N_8969,N_8865);
nor U10014 (N_10014,N_8841,N_9186);
nand U10015 (N_10015,N_8877,N_8889);
xnor U10016 (N_10016,N_8884,N_9432);
nor U10017 (N_10017,N_9115,N_8947);
and U10018 (N_10018,N_9491,N_8913);
xor U10019 (N_10019,N_9446,N_9491);
or U10020 (N_10020,N_9285,N_9212);
and U10021 (N_10021,N_9211,N_9043);
nor U10022 (N_10022,N_9554,N_9550);
nand U10023 (N_10023,N_9532,N_9544);
nor U10024 (N_10024,N_9348,N_9262);
nand U10025 (N_10025,N_9274,N_9173);
or U10026 (N_10026,N_9018,N_9506);
nor U10027 (N_10027,N_9254,N_9178);
nor U10028 (N_10028,N_9547,N_9014);
nor U10029 (N_10029,N_9096,N_9297);
or U10030 (N_10030,N_9394,N_9525);
xnor U10031 (N_10031,N_9007,N_9000);
xor U10032 (N_10032,N_8934,N_8871);
or U10033 (N_10033,N_9376,N_8849);
or U10034 (N_10034,N_9038,N_9530);
and U10035 (N_10035,N_9041,N_9338);
xnor U10036 (N_10036,N_9102,N_9205);
xnor U10037 (N_10037,N_8802,N_9167);
nand U10038 (N_10038,N_9424,N_9144);
or U10039 (N_10039,N_9292,N_8856);
or U10040 (N_10040,N_8969,N_9360);
nand U10041 (N_10041,N_9566,N_8904);
and U10042 (N_10042,N_9448,N_9536);
nand U10043 (N_10043,N_9003,N_9277);
nand U10044 (N_10044,N_9342,N_9591);
or U10045 (N_10045,N_8948,N_9457);
nor U10046 (N_10046,N_9283,N_9159);
nor U10047 (N_10047,N_8890,N_8846);
xnor U10048 (N_10048,N_9334,N_8963);
nand U10049 (N_10049,N_9598,N_9450);
and U10050 (N_10050,N_9255,N_8965);
nand U10051 (N_10051,N_9578,N_9186);
nand U10052 (N_10052,N_8926,N_8869);
or U10053 (N_10053,N_9547,N_9599);
xor U10054 (N_10054,N_9485,N_8957);
xor U10055 (N_10055,N_9484,N_9436);
or U10056 (N_10056,N_8916,N_9327);
nor U10057 (N_10057,N_9532,N_9325);
or U10058 (N_10058,N_9442,N_9358);
or U10059 (N_10059,N_9276,N_8962);
and U10060 (N_10060,N_9577,N_9299);
xor U10061 (N_10061,N_9585,N_9287);
nor U10062 (N_10062,N_9084,N_9224);
xnor U10063 (N_10063,N_9508,N_9068);
nand U10064 (N_10064,N_9279,N_8860);
nand U10065 (N_10065,N_9313,N_9202);
xor U10066 (N_10066,N_9068,N_9201);
nand U10067 (N_10067,N_9355,N_9282);
or U10068 (N_10068,N_9459,N_9000);
nand U10069 (N_10069,N_9528,N_9155);
xnor U10070 (N_10070,N_8992,N_9195);
and U10071 (N_10071,N_9196,N_9432);
or U10072 (N_10072,N_8983,N_9224);
or U10073 (N_10073,N_9333,N_9488);
xnor U10074 (N_10074,N_9099,N_9221);
or U10075 (N_10075,N_9484,N_9055);
or U10076 (N_10076,N_9576,N_9443);
or U10077 (N_10077,N_9371,N_8992);
and U10078 (N_10078,N_9530,N_9356);
nor U10079 (N_10079,N_9272,N_9360);
or U10080 (N_10080,N_9255,N_9587);
and U10081 (N_10081,N_9523,N_9347);
and U10082 (N_10082,N_8817,N_9471);
or U10083 (N_10083,N_8846,N_9140);
and U10084 (N_10084,N_9222,N_9592);
xor U10085 (N_10085,N_9049,N_9548);
and U10086 (N_10086,N_8950,N_9229);
or U10087 (N_10087,N_9456,N_9349);
and U10088 (N_10088,N_8952,N_9017);
and U10089 (N_10089,N_9586,N_9074);
or U10090 (N_10090,N_9576,N_9204);
xor U10091 (N_10091,N_8859,N_9164);
and U10092 (N_10092,N_9094,N_9075);
nor U10093 (N_10093,N_9380,N_8805);
or U10094 (N_10094,N_9321,N_9062);
nand U10095 (N_10095,N_9464,N_9163);
and U10096 (N_10096,N_9163,N_9479);
nand U10097 (N_10097,N_8853,N_9422);
nor U10098 (N_10098,N_9105,N_8961);
xnor U10099 (N_10099,N_9023,N_9210);
nand U10100 (N_10100,N_8952,N_9579);
xor U10101 (N_10101,N_9326,N_8909);
nand U10102 (N_10102,N_9162,N_9228);
nor U10103 (N_10103,N_9358,N_9227);
xor U10104 (N_10104,N_9431,N_8982);
and U10105 (N_10105,N_9029,N_9418);
nor U10106 (N_10106,N_9017,N_9531);
xnor U10107 (N_10107,N_9482,N_9528);
or U10108 (N_10108,N_9579,N_9071);
nand U10109 (N_10109,N_9290,N_9593);
and U10110 (N_10110,N_9381,N_9317);
and U10111 (N_10111,N_9160,N_9096);
or U10112 (N_10112,N_8803,N_9160);
or U10113 (N_10113,N_9148,N_9486);
and U10114 (N_10114,N_9212,N_9401);
nor U10115 (N_10115,N_9228,N_8816);
and U10116 (N_10116,N_8911,N_9236);
or U10117 (N_10117,N_8848,N_8810);
and U10118 (N_10118,N_9255,N_8883);
or U10119 (N_10119,N_9244,N_9570);
xor U10120 (N_10120,N_8978,N_9366);
nand U10121 (N_10121,N_9036,N_8933);
and U10122 (N_10122,N_9042,N_9182);
xnor U10123 (N_10123,N_9575,N_9317);
and U10124 (N_10124,N_9064,N_8905);
nor U10125 (N_10125,N_8876,N_8868);
or U10126 (N_10126,N_9216,N_9338);
xor U10127 (N_10127,N_9251,N_9394);
xnor U10128 (N_10128,N_9226,N_9502);
and U10129 (N_10129,N_9552,N_8897);
or U10130 (N_10130,N_9030,N_9504);
and U10131 (N_10131,N_9103,N_9194);
nand U10132 (N_10132,N_9115,N_9135);
or U10133 (N_10133,N_9040,N_8856);
or U10134 (N_10134,N_9117,N_8849);
or U10135 (N_10135,N_9295,N_8893);
nor U10136 (N_10136,N_8804,N_8948);
nand U10137 (N_10137,N_9124,N_9348);
xor U10138 (N_10138,N_8964,N_9114);
nand U10139 (N_10139,N_9591,N_9510);
and U10140 (N_10140,N_9596,N_9269);
nand U10141 (N_10141,N_9501,N_9390);
nor U10142 (N_10142,N_9288,N_9202);
nand U10143 (N_10143,N_8924,N_8841);
xor U10144 (N_10144,N_8942,N_9136);
xnor U10145 (N_10145,N_9302,N_9032);
xor U10146 (N_10146,N_9161,N_8886);
nor U10147 (N_10147,N_9230,N_9081);
nand U10148 (N_10148,N_9351,N_9048);
and U10149 (N_10149,N_9421,N_9271);
and U10150 (N_10150,N_8963,N_8868);
nor U10151 (N_10151,N_8807,N_9417);
xor U10152 (N_10152,N_9480,N_9127);
or U10153 (N_10153,N_9399,N_9309);
and U10154 (N_10154,N_8958,N_9445);
and U10155 (N_10155,N_8952,N_8963);
or U10156 (N_10156,N_8935,N_9581);
nand U10157 (N_10157,N_9357,N_8859);
and U10158 (N_10158,N_9057,N_9467);
nor U10159 (N_10159,N_8914,N_9162);
nand U10160 (N_10160,N_9309,N_9157);
and U10161 (N_10161,N_9404,N_9300);
xor U10162 (N_10162,N_9294,N_9363);
xor U10163 (N_10163,N_8818,N_9252);
or U10164 (N_10164,N_9542,N_9218);
xnor U10165 (N_10165,N_9162,N_9140);
nor U10166 (N_10166,N_9439,N_8908);
nand U10167 (N_10167,N_9340,N_9127);
or U10168 (N_10168,N_8848,N_9271);
and U10169 (N_10169,N_8843,N_9594);
or U10170 (N_10170,N_8916,N_9448);
nand U10171 (N_10171,N_9104,N_9553);
or U10172 (N_10172,N_8997,N_8940);
xnor U10173 (N_10173,N_9287,N_9455);
nand U10174 (N_10174,N_9373,N_9269);
nand U10175 (N_10175,N_9063,N_9345);
nor U10176 (N_10176,N_8999,N_8804);
nor U10177 (N_10177,N_8983,N_9170);
nor U10178 (N_10178,N_9238,N_8880);
nand U10179 (N_10179,N_9349,N_8845);
xnor U10180 (N_10180,N_9233,N_9404);
or U10181 (N_10181,N_9581,N_9536);
nor U10182 (N_10182,N_8935,N_9103);
or U10183 (N_10183,N_9390,N_9496);
and U10184 (N_10184,N_9363,N_9488);
nor U10185 (N_10185,N_9426,N_9268);
nor U10186 (N_10186,N_8914,N_9574);
nor U10187 (N_10187,N_8816,N_9248);
and U10188 (N_10188,N_8885,N_9183);
nand U10189 (N_10189,N_9043,N_9429);
or U10190 (N_10190,N_9013,N_9462);
nor U10191 (N_10191,N_9204,N_8877);
xor U10192 (N_10192,N_9213,N_8956);
and U10193 (N_10193,N_9330,N_9022);
nand U10194 (N_10194,N_9334,N_8863);
nor U10195 (N_10195,N_9572,N_9040);
nor U10196 (N_10196,N_9117,N_9393);
or U10197 (N_10197,N_9216,N_9365);
nand U10198 (N_10198,N_9374,N_9122);
nor U10199 (N_10199,N_9049,N_9216);
nand U10200 (N_10200,N_9263,N_8937);
or U10201 (N_10201,N_9544,N_9015);
or U10202 (N_10202,N_9557,N_9160);
and U10203 (N_10203,N_9016,N_9581);
xnor U10204 (N_10204,N_8911,N_9433);
xor U10205 (N_10205,N_8935,N_9395);
xor U10206 (N_10206,N_9156,N_9113);
xor U10207 (N_10207,N_9188,N_9100);
xnor U10208 (N_10208,N_9465,N_9411);
nor U10209 (N_10209,N_9454,N_9264);
xnor U10210 (N_10210,N_9393,N_9340);
nor U10211 (N_10211,N_9144,N_9359);
or U10212 (N_10212,N_9278,N_9059);
and U10213 (N_10213,N_9107,N_8988);
xor U10214 (N_10214,N_9131,N_9419);
nor U10215 (N_10215,N_9491,N_9377);
and U10216 (N_10216,N_8803,N_9167);
or U10217 (N_10217,N_8856,N_9587);
and U10218 (N_10218,N_8829,N_9505);
nand U10219 (N_10219,N_9022,N_9318);
or U10220 (N_10220,N_9183,N_9573);
or U10221 (N_10221,N_9406,N_9257);
or U10222 (N_10222,N_9522,N_9419);
and U10223 (N_10223,N_9202,N_9458);
and U10224 (N_10224,N_9567,N_9066);
nand U10225 (N_10225,N_9558,N_9322);
xnor U10226 (N_10226,N_9217,N_8845);
and U10227 (N_10227,N_8992,N_9443);
or U10228 (N_10228,N_9152,N_9369);
nor U10229 (N_10229,N_8861,N_9446);
nand U10230 (N_10230,N_9339,N_9271);
or U10231 (N_10231,N_9132,N_8971);
and U10232 (N_10232,N_9078,N_9583);
or U10233 (N_10233,N_8906,N_9171);
and U10234 (N_10234,N_9470,N_9243);
nand U10235 (N_10235,N_9488,N_9230);
nand U10236 (N_10236,N_8937,N_8883);
and U10237 (N_10237,N_8848,N_9559);
and U10238 (N_10238,N_8866,N_9539);
nor U10239 (N_10239,N_9518,N_9454);
xnor U10240 (N_10240,N_9482,N_9285);
and U10241 (N_10241,N_9579,N_9130);
and U10242 (N_10242,N_9351,N_8860);
nor U10243 (N_10243,N_8992,N_9581);
nor U10244 (N_10244,N_8801,N_9101);
nand U10245 (N_10245,N_9328,N_8930);
xor U10246 (N_10246,N_8984,N_9239);
nand U10247 (N_10247,N_9461,N_9299);
or U10248 (N_10248,N_8901,N_9111);
and U10249 (N_10249,N_9309,N_9368);
and U10250 (N_10250,N_9084,N_9564);
xnor U10251 (N_10251,N_9579,N_9243);
nor U10252 (N_10252,N_9328,N_8853);
or U10253 (N_10253,N_9193,N_8839);
nor U10254 (N_10254,N_8976,N_9375);
and U10255 (N_10255,N_9400,N_8964);
nand U10256 (N_10256,N_9234,N_9361);
nor U10257 (N_10257,N_9509,N_9389);
xor U10258 (N_10258,N_9546,N_9507);
and U10259 (N_10259,N_8816,N_9520);
or U10260 (N_10260,N_9307,N_9319);
and U10261 (N_10261,N_8980,N_9461);
or U10262 (N_10262,N_8829,N_9515);
xnor U10263 (N_10263,N_8978,N_9311);
nand U10264 (N_10264,N_8997,N_9513);
and U10265 (N_10265,N_8816,N_9546);
nor U10266 (N_10266,N_9255,N_9558);
nand U10267 (N_10267,N_8935,N_9482);
nor U10268 (N_10268,N_9106,N_9170);
or U10269 (N_10269,N_9085,N_8846);
and U10270 (N_10270,N_9315,N_9396);
xnor U10271 (N_10271,N_8871,N_9154);
and U10272 (N_10272,N_9324,N_9047);
nand U10273 (N_10273,N_9005,N_9194);
nor U10274 (N_10274,N_9006,N_9464);
nor U10275 (N_10275,N_8812,N_9538);
and U10276 (N_10276,N_9353,N_9226);
nor U10277 (N_10277,N_8836,N_9349);
nor U10278 (N_10278,N_9029,N_8818);
nor U10279 (N_10279,N_9122,N_9501);
nor U10280 (N_10280,N_8845,N_8966);
nand U10281 (N_10281,N_9298,N_8984);
or U10282 (N_10282,N_9586,N_9215);
nor U10283 (N_10283,N_9455,N_8854);
nand U10284 (N_10284,N_9448,N_8903);
and U10285 (N_10285,N_9259,N_8921);
nand U10286 (N_10286,N_9190,N_9432);
nand U10287 (N_10287,N_9234,N_9068);
xnor U10288 (N_10288,N_9322,N_9084);
and U10289 (N_10289,N_8952,N_8921);
nand U10290 (N_10290,N_8963,N_9083);
nor U10291 (N_10291,N_9393,N_9001);
nand U10292 (N_10292,N_9434,N_9354);
or U10293 (N_10293,N_8867,N_8821);
nor U10294 (N_10294,N_9585,N_9039);
nand U10295 (N_10295,N_9433,N_9455);
xor U10296 (N_10296,N_9156,N_9423);
or U10297 (N_10297,N_9487,N_8853);
xnor U10298 (N_10298,N_9522,N_8923);
nand U10299 (N_10299,N_9539,N_9057);
xor U10300 (N_10300,N_9251,N_9071);
or U10301 (N_10301,N_9284,N_9286);
xor U10302 (N_10302,N_9469,N_9182);
and U10303 (N_10303,N_9516,N_9434);
and U10304 (N_10304,N_9591,N_9176);
and U10305 (N_10305,N_9509,N_9391);
and U10306 (N_10306,N_9123,N_9381);
nand U10307 (N_10307,N_8872,N_8881);
nor U10308 (N_10308,N_9224,N_8943);
and U10309 (N_10309,N_9045,N_9588);
or U10310 (N_10310,N_8895,N_9102);
nand U10311 (N_10311,N_9268,N_9418);
and U10312 (N_10312,N_9425,N_8839);
and U10313 (N_10313,N_8886,N_9578);
nor U10314 (N_10314,N_8968,N_9098);
or U10315 (N_10315,N_9199,N_9003);
and U10316 (N_10316,N_9424,N_9094);
nand U10317 (N_10317,N_9072,N_9578);
nor U10318 (N_10318,N_9373,N_9527);
nor U10319 (N_10319,N_9316,N_9248);
and U10320 (N_10320,N_9163,N_9401);
and U10321 (N_10321,N_9098,N_9484);
nand U10322 (N_10322,N_9389,N_9157);
nor U10323 (N_10323,N_8821,N_9376);
or U10324 (N_10324,N_9189,N_8876);
xnor U10325 (N_10325,N_9453,N_8863);
and U10326 (N_10326,N_9589,N_8812);
nand U10327 (N_10327,N_9128,N_9164);
and U10328 (N_10328,N_9588,N_8884);
xor U10329 (N_10329,N_9415,N_9502);
and U10330 (N_10330,N_8934,N_9355);
xnor U10331 (N_10331,N_8986,N_9384);
and U10332 (N_10332,N_9083,N_9484);
xor U10333 (N_10333,N_9248,N_9127);
nand U10334 (N_10334,N_9180,N_9080);
xnor U10335 (N_10335,N_8899,N_9109);
nor U10336 (N_10336,N_9341,N_9392);
or U10337 (N_10337,N_8997,N_9204);
xnor U10338 (N_10338,N_9337,N_8946);
nand U10339 (N_10339,N_9316,N_9575);
and U10340 (N_10340,N_9334,N_9254);
xor U10341 (N_10341,N_9157,N_9278);
and U10342 (N_10342,N_8921,N_8974);
or U10343 (N_10343,N_8806,N_9082);
nand U10344 (N_10344,N_9463,N_9492);
or U10345 (N_10345,N_9233,N_9475);
xor U10346 (N_10346,N_9597,N_9554);
xor U10347 (N_10347,N_8923,N_9428);
xnor U10348 (N_10348,N_9070,N_8851);
and U10349 (N_10349,N_9089,N_9443);
xnor U10350 (N_10350,N_9080,N_9276);
and U10351 (N_10351,N_8825,N_9430);
or U10352 (N_10352,N_9596,N_8928);
nand U10353 (N_10353,N_9083,N_9522);
nand U10354 (N_10354,N_9359,N_9420);
nand U10355 (N_10355,N_9438,N_8934);
nand U10356 (N_10356,N_8878,N_9388);
nand U10357 (N_10357,N_8901,N_9590);
nand U10358 (N_10358,N_9591,N_8915);
nor U10359 (N_10359,N_9300,N_9167);
or U10360 (N_10360,N_9064,N_9338);
and U10361 (N_10361,N_9418,N_9543);
and U10362 (N_10362,N_9397,N_9140);
xor U10363 (N_10363,N_9285,N_9558);
xnor U10364 (N_10364,N_8846,N_9304);
and U10365 (N_10365,N_9523,N_9232);
and U10366 (N_10366,N_8975,N_8910);
xnor U10367 (N_10367,N_9389,N_9079);
xnor U10368 (N_10368,N_9473,N_8959);
nor U10369 (N_10369,N_9349,N_9441);
xnor U10370 (N_10370,N_9120,N_9004);
nor U10371 (N_10371,N_9229,N_8881);
and U10372 (N_10372,N_9487,N_9498);
nor U10373 (N_10373,N_9415,N_9172);
or U10374 (N_10374,N_9192,N_9063);
nor U10375 (N_10375,N_9118,N_9081);
xor U10376 (N_10376,N_9303,N_8834);
xnor U10377 (N_10377,N_9598,N_9152);
nor U10378 (N_10378,N_9034,N_9091);
or U10379 (N_10379,N_9440,N_9354);
or U10380 (N_10380,N_9403,N_9050);
nand U10381 (N_10381,N_9335,N_9275);
nand U10382 (N_10382,N_9413,N_9472);
nor U10383 (N_10383,N_9324,N_8979);
nand U10384 (N_10384,N_8989,N_9077);
and U10385 (N_10385,N_8820,N_9361);
xnor U10386 (N_10386,N_8957,N_9365);
xor U10387 (N_10387,N_9485,N_9323);
or U10388 (N_10388,N_8833,N_9083);
nand U10389 (N_10389,N_9240,N_8859);
nand U10390 (N_10390,N_9152,N_9358);
and U10391 (N_10391,N_9551,N_8821);
nor U10392 (N_10392,N_9442,N_9552);
nor U10393 (N_10393,N_8921,N_9150);
nand U10394 (N_10394,N_9235,N_9015);
and U10395 (N_10395,N_8997,N_8956);
nor U10396 (N_10396,N_9037,N_9456);
and U10397 (N_10397,N_8955,N_9413);
and U10398 (N_10398,N_8843,N_9014);
nand U10399 (N_10399,N_9044,N_9174);
nand U10400 (N_10400,N_9875,N_10168);
nand U10401 (N_10401,N_9664,N_9725);
xor U10402 (N_10402,N_9612,N_10292);
xnor U10403 (N_10403,N_10196,N_10377);
or U10404 (N_10404,N_10156,N_10386);
or U10405 (N_10405,N_10216,N_9615);
nand U10406 (N_10406,N_10353,N_9825);
and U10407 (N_10407,N_9985,N_10065);
nor U10408 (N_10408,N_10212,N_10142);
and U10409 (N_10409,N_9967,N_9915);
nand U10410 (N_10410,N_9837,N_10193);
and U10411 (N_10411,N_10203,N_10385);
nor U10412 (N_10412,N_10122,N_9932);
or U10413 (N_10413,N_10128,N_10069);
and U10414 (N_10414,N_10033,N_9818);
or U10415 (N_10415,N_9833,N_10038);
nand U10416 (N_10416,N_10341,N_9844);
or U10417 (N_10417,N_10008,N_9799);
and U10418 (N_10418,N_9692,N_10324);
xnor U10419 (N_10419,N_10136,N_9756);
xnor U10420 (N_10420,N_9783,N_10003);
xnor U10421 (N_10421,N_9732,N_10223);
and U10422 (N_10422,N_10201,N_9754);
nor U10423 (N_10423,N_9801,N_10296);
nor U10424 (N_10424,N_9919,N_9720);
nand U10425 (N_10425,N_10005,N_9687);
nand U10426 (N_10426,N_9622,N_10100);
xor U10427 (N_10427,N_10250,N_10130);
and U10428 (N_10428,N_10285,N_9872);
or U10429 (N_10429,N_9672,N_10246);
nand U10430 (N_10430,N_9769,N_9751);
nand U10431 (N_10431,N_10176,N_9616);
or U10432 (N_10432,N_10211,N_9807);
or U10433 (N_10433,N_10058,N_10036);
or U10434 (N_10434,N_9847,N_9618);
nand U10435 (N_10435,N_10152,N_9899);
and U10436 (N_10436,N_9701,N_9761);
nor U10437 (N_10437,N_10242,N_10148);
nor U10438 (N_10438,N_9611,N_9924);
and U10439 (N_10439,N_10095,N_10360);
xor U10440 (N_10440,N_9662,N_10145);
xor U10441 (N_10441,N_9954,N_10025);
and U10442 (N_10442,N_9710,N_10253);
xnor U10443 (N_10443,N_10293,N_9930);
xor U10444 (N_10444,N_10303,N_10367);
xnor U10445 (N_10445,N_10396,N_10230);
nand U10446 (N_10446,N_9988,N_10042);
xor U10447 (N_10447,N_10300,N_9714);
nand U10448 (N_10448,N_10037,N_9910);
and U10449 (N_10449,N_10281,N_10147);
xor U10450 (N_10450,N_9690,N_9639);
and U10451 (N_10451,N_10312,N_10260);
or U10452 (N_10452,N_9881,N_10133);
nor U10453 (N_10453,N_10083,N_9738);
and U10454 (N_10454,N_10328,N_9858);
or U10455 (N_10455,N_10101,N_9921);
and U10456 (N_10456,N_10155,N_9685);
nor U10457 (N_10457,N_9834,N_10023);
and U10458 (N_10458,N_10249,N_9607);
nor U10459 (N_10459,N_10080,N_9675);
and U10460 (N_10460,N_9730,N_9992);
or U10461 (N_10461,N_10110,N_9856);
and U10462 (N_10462,N_9909,N_10395);
xnor U10463 (N_10463,N_9700,N_9654);
nand U10464 (N_10464,N_10357,N_9755);
xor U10465 (N_10465,N_10186,N_10141);
xor U10466 (N_10466,N_9901,N_9680);
and U10467 (N_10467,N_9752,N_9952);
or U10468 (N_10468,N_9892,N_10371);
or U10469 (N_10469,N_10368,N_9625);
nand U10470 (N_10470,N_10317,N_10107);
xor U10471 (N_10471,N_9779,N_9614);
nand U10472 (N_10472,N_9841,N_10084);
and U10473 (N_10473,N_9913,N_10335);
and U10474 (N_10474,N_9686,N_9650);
nand U10475 (N_10475,N_9796,N_10092);
and U10476 (N_10476,N_10298,N_10343);
nor U10477 (N_10477,N_10086,N_10344);
nand U10478 (N_10478,N_9931,N_9991);
nand U10479 (N_10479,N_9980,N_10280);
xor U10480 (N_10480,N_9829,N_10184);
and U10481 (N_10481,N_9646,N_9653);
xnor U10482 (N_10482,N_10125,N_10308);
nor U10483 (N_10483,N_9811,N_9998);
and U10484 (N_10484,N_9953,N_10178);
xor U10485 (N_10485,N_9823,N_10181);
or U10486 (N_10486,N_9806,N_10195);
nand U10487 (N_10487,N_10289,N_10007);
nand U10488 (N_10488,N_10073,N_9977);
nand U10489 (N_10489,N_10167,N_9704);
nand U10490 (N_10490,N_10302,N_9603);
or U10491 (N_10491,N_9958,N_9822);
nand U10492 (N_10492,N_10229,N_9842);
and U10493 (N_10493,N_10185,N_10153);
nand U10494 (N_10494,N_9859,N_10102);
and U10495 (N_10495,N_9708,N_9928);
nand U10496 (N_10496,N_9627,N_10235);
or U10497 (N_10497,N_10219,N_10266);
nor U10498 (N_10498,N_9982,N_9969);
nand U10499 (N_10499,N_10275,N_9846);
nand U10500 (N_10500,N_9883,N_10113);
and U10501 (N_10501,N_10217,N_9962);
xnor U10502 (N_10502,N_9869,N_10026);
or U10503 (N_10503,N_9896,N_9864);
and U10504 (N_10504,N_10391,N_10263);
and U10505 (N_10505,N_10162,N_9816);
xnor U10506 (N_10506,N_10019,N_10314);
nand U10507 (N_10507,N_9891,N_9719);
and U10508 (N_10508,N_9854,N_10390);
nand U10509 (N_10509,N_9966,N_9906);
xor U10510 (N_10510,N_9814,N_10127);
nor U10511 (N_10511,N_10261,N_10374);
xnor U10512 (N_10512,N_9666,N_10094);
xor U10513 (N_10513,N_10286,N_10311);
nand U10514 (N_10514,N_10143,N_10331);
and U10515 (N_10515,N_10048,N_9734);
nor U10516 (N_10516,N_9773,N_10067);
nand U10517 (N_10517,N_9792,N_10050);
xnor U10518 (N_10518,N_9624,N_10204);
or U10519 (N_10519,N_9917,N_9623);
xor U10520 (N_10520,N_9983,N_10252);
or U10521 (N_10521,N_10329,N_9688);
nand U10522 (N_10522,N_10149,N_9602);
or U10523 (N_10523,N_9790,N_9750);
and U10524 (N_10524,N_10049,N_10061);
nand U10525 (N_10525,N_9772,N_10154);
nand U10526 (N_10526,N_10109,N_9795);
and U10527 (N_10527,N_9857,N_9873);
xor U10528 (N_10528,N_10233,N_10190);
xnor U10529 (N_10529,N_9741,N_10040);
xnor U10530 (N_10530,N_10258,N_10015);
or U10531 (N_10531,N_10220,N_9999);
nor U10532 (N_10532,N_10332,N_9984);
or U10533 (N_10533,N_10316,N_10089);
xnor U10534 (N_10534,N_10369,N_10081);
xor U10535 (N_10535,N_9762,N_9996);
nand U10536 (N_10536,N_9684,N_10277);
nor U10537 (N_10537,N_9640,N_9956);
nor U10538 (N_10538,N_9871,N_9824);
or U10539 (N_10539,N_9828,N_9944);
and U10540 (N_10540,N_9911,N_9886);
nor U10541 (N_10541,N_9706,N_9948);
or U10542 (N_10542,N_10228,N_10057);
xnor U10543 (N_10543,N_10132,N_9731);
nor U10544 (N_10544,N_9923,N_10175);
or U10545 (N_10545,N_9889,N_9975);
xor U10546 (N_10546,N_9767,N_10001);
xor U10547 (N_10547,N_10160,N_10068);
nand U10548 (N_10548,N_10174,N_10345);
and U10549 (N_10549,N_9939,N_10192);
and U10550 (N_10550,N_10254,N_10375);
nor U10551 (N_10551,N_10268,N_10234);
and U10552 (N_10552,N_10207,N_9938);
xor U10553 (N_10553,N_9691,N_10256);
and U10554 (N_10554,N_9709,N_9771);
or U10555 (N_10555,N_9849,N_10075);
or U10556 (N_10556,N_9964,N_10098);
and U10557 (N_10557,N_10096,N_9884);
and U10558 (N_10558,N_9997,N_10313);
nor U10559 (N_10559,N_10004,N_9723);
nor U10560 (N_10560,N_10010,N_9813);
and U10561 (N_10561,N_10208,N_9876);
xnor U10562 (N_10562,N_10118,N_10151);
or U10563 (N_10563,N_10269,N_9821);
or U10564 (N_10564,N_10271,N_10021);
nor U10565 (N_10565,N_9712,N_9642);
and U10566 (N_10566,N_9718,N_10326);
nor U10567 (N_10567,N_10022,N_10397);
and U10568 (N_10568,N_9788,N_10294);
or U10569 (N_10569,N_9839,N_10224);
xor U10570 (N_10570,N_10044,N_9765);
or U10571 (N_10571,N_9840,N_9610);
nand U10572 (N_10572,N_10123,N_9621);
nand U10573 (N_10573,N_9986,N_10169);
nor U10574 (N_10574,N_9933,N_9798);
xor U10575 (N_10575,N_9781,N_9605);
nor U10576 (N_10576,N_10077,N_9895);
nor U10577 (N_10577,N_10205,N_9743);
nand U10578 (N_10578,N_10350,N_9608);
nand U10579 (N_10579,N_9716,N_10214);
nand U10580 (N_10580,N_10105,N_10020);
xor U10581 (N_10581,N_9914,N_10059);
or U10582 (N_10582,N_10039,N_10334);
nand U10583 (N_10583,N_9705,N_10189);
nor U10584 (N_10584,N_9925,N_10288);
nand U10585 (N_10585,N_9989,N_9733);
or U10586 (N_10586,N_9658,N_9715);
and U10587 (N_10587,N_10278,N_9656);
nor U10588 (N_10588,N_9689,N_10355);
xor U10589 (N_10589,N_10120,N_10180);
and U10590 (N_10590,N_9918,N_9679);
and U10591 (N_10591,N_10115,N_10137);
or U10592 (N_10592,N_9759,N_9673);
nand U10593 (N_10593,N_10315,N_9763);
nor U10594 (N_10594,N_9667,N_10321);
and U10595 (N_10595,N_9641,N_9628);
xor U10596 (N_10596,N_10131,N_10199);
and U10597 (N_10597,N_9668,N_9893);
nor U10598 (N_10598,N_10093,N_9619);
nor U10599 (N_10599,N_10265,N_10140);
nor U10600 (N_10600,N_9870,N_9620);
and U10601 (N_10601,N_9736,N_9676);
nor U10602 (N_10602,N_10247,N_10304);
nand U10603 (N_10603,N_9739,N_10103);
or U10604 (N_10604,N_9636,N_9990);
nand U10605 (N_10605,N_9742,N_10264);
nor U10606 (N_10606,N_10393,N_9946);
and U10607 (N_10607,N_9782,N_10273);
nand U10608 (N_10608,N_10319,N_9951);
xnor U10609 (N_10609,N_10165,N_9696);
nand U10610 (N_10610,N_10309,N_10097);
and U10611 (N_10611,N_10274,N_10215);
or U10612 (N_10612,N_9630,N_9703);
xnor U10613 (N_10613,N_9766,N_9866);
nor U10614 (N_10614,N_10135,N_10342);
nand U10615 (N_10615,N_10177,N_9937);
xor U10616 (N_10616,N_9637,N_9810);
nand U10617 (N_10617,N_9749,N_10138);
xor U10618 (N_10618,N_10336,N_10047);
nand U10619 (N_10619,N_9745,N_9727);
or U10620 (N_10620,N_10222,N_10221);
or U10621 (N_10621,N_9838,N_10259);
or U10622 (N_10622,N_9643,N_9655);
or U10623 (N_10623,N_9764,N_10183);
and U10624 (N_10624,N_10394,N_9970);
nor U10625 (N_10625,N_10164,N_10240);
nand U10626 (N_10626,N_10239,N_9981);
or U10627 (N_10627,N_9916,N_10046);
nand U10628 (N_10628,N_10066,N_10340);
and U10629 (N_10629,N_9827,N_9945);
xnor U10630 (N_10630,N_9855,N_9853);
or U10631 (N_10631,N_9880,N_10284);
and U10632 (N_10632,N_9797,N_9835);
xor U10633 (N_10633,N_10231,N_9809);
nor U10634 (N_10634,N_10041,N_10257);
nor U10635 (N_10635,N_9760,N_9777);
nand U10636 (N_10636,N_9744,N_10173);
or U10637 (N_10637,N_10376,N_9647);
nor U10638 (N_10638,N_9648,N_10055);
and U10639 (N_10639,N_10070,N_10129);
xnor U10640 (N_10640,N_10283,N_9753);
and U10641 (N_10641,N_10099,N_10000);
and U10642 (N_10642,N_10139,N_9860);
nor U10643 (N_10643,N_10063,N_10194);
or U10644 (N_10644,N_10245,N_9845);
xor U10645 (N_10645,N_10398,N_9713);
or U10646 (N_10646,N_9632,N_9697);
nor U10647 (N_10647,N_10232,N_9617);
and U10648 (N_10648,N_10013,N_10327);
nor U10649 (N_10649,N_10226,N_9663);
and U10650 (N_10650,N_10380,N_10062);
or U10651 (N_10651,N_10213,N_10387);
or U10652 (N_10652,N_10060,N_9867);
xnor U10653 (N_10653,N_9757,N_10348);
and U10654 (N_10654,N_10389,N_10337);
xor U10655 (N_10655,N_9631,N_9936);
nand U10656 (N_10656,N_9897,N_10379);
and U10657 (N_10657,N_9638,N_9890);
xor U10658 (N_10658,N_10354,N_9994);
xor U10659 (N_10659,N_9758,N_9670);
nor U10660 (N_10660,N_9768,N_9898);
nand U10661 (N_10661,N_9746,N_9888);
nand U10662 (N_10662,N_10297,N_10209);
nor U10663 (N_10663,N_9702,N_10323);
or U10664 (N_10664,N_10076,N_9874);
nand U10665 (N_10665,N_9695,N_9852);
xor U10666 (N_10666,N_9633,N_10053);
nand U10667 (N_10667,N_9786,N_10157);
nor U10668 (N_10668,N_9912,N_10146);
and U10669 (N_10669,N_9965,N_10104);
and U10670 (N_10670,N_9613,N_9740);
and U10671 (N_10671,N_10363,N_9661);
nor U10672 (N_10672,N_9862,N_10087);
nand U10673 (N_10673,N_9905,N_10392);
nor U10674 (N_10674,N_9800,N_9935);
xnor U10675 (N_10675,N_10006,N_10171);
nor U10676 (N_10676,N_9748,N_10134);
nor U10677 (N_10677,N_10187,N_9717);
nand U10678 (N_10678,N_9728,N_9606);
or U10679 (N_10679,N_9683,N_9882);
nand U10680 (N_10680,N_9803,N_10043);
nor U10681 (N_10681,N_10361,N_9793);
or U10682 (N_10682,N_10002,N_10114);
nor U10683 (N_10683,N_9776,N_10017);
nand U10684 (N_10684,N_9735,N_9922);
nor U10685 (N_10685,N_9600,N_10351);
and U10686 (N_10686,N_9707,N_10279);
xnor U10687 (N_10687,N_9836,N_9729);
xnor U10688 (N_10688,N_10325,N_9963);
xor U10689 (N_10689,N_10035,N_9681);
nand U10690 (N_10690,N_9878,N_10287);
or U10691 (N_10691,N_9787,N_10365);
xor U10692 (N_10692,N_10029,N_9993);
or U10693 (N_10693,N_9894,N_9819);
or U10694 (N_10694,N_10111,N_9861);
and U10695 (N_10695,N_10290,N_9805);
nand U10696 (N_10696,N_9974,N_10248);
nand U10697 (N_10697,N_10262,N_10082);
xor U10698 (N_10698,N_9678,N_9802);
xor U10699 (N_10699,N_10272,N_9942);
nor U10700 (N_10700,N_10014,N_10238);
or U10701 (N_10701,N_10079,N_10306);
and U10702 (N_10702,N_9959,N_10295);
xor U10703 (N_10703,N_9794,N_10191);
or U10704 (N_10704,N_9900,N_9651);
nor U10705 (N_10705,N_9950,N_9721);
and U10706 (N_10706,N_10158,N_10352);
or U10707 (N_10707,N_10072,N_10399);
or U10708 (N_10708,N_9724,N_10244);
nor U10709 (N_10709,N_9961,N_10119);
and U10710 (N_10710,N_9940,N_10056);
and U10711 (N_10711,N_9657,N_10276);
or U10712 (N_10712,N_9789,N_10381);
nor U10713 (N_10713,N_9812,N_9635);
nor U10714 (N_10714,N_10024,N_9671);
nand U10715 (N_10715,N_9955,N_9652);
or U10716 (N_10716,N_9960,N_10200);
xor U10717 (N_10717,N_9629,N_10161);
nand U10718 (N_10718,N_9804,N_10144);
nor U10719 (N_10719,N_10318,N_9868);
nor U10720 (N_10720,N_10267,N_10237);
nand U10721 (N_10721,N_10243,N_9877);
xnor U10722 (N_10722,N_10349,N_9649);
nand U10723 (N_10723,N_10198,N_10126);
nor U10724 (N_10724,N_9775,N_9601);
xnor U10725 (N_10725,N_9885,N_9747);
or U10726 (N_10726,N_10358,N_9850);
nor U10727 (N_10727,N_9820,N_10028);
nand U10728 (N_10728,N_9780,N_9848);
nor U10729 (N_10729,N_9609,N_10030);
or U10730 (N_10730,N_9626,N_9979);
nor U10731 (N_10731,N_9887,N_10378);
xnor U10732 (N_10732,N_10116,N_10346);
nor U10733 (N_10733,N_10112,N_9865);
or U10734 (N_10734,N_9698,N_9815);
or U10735 (N_10735,N_9831,N_10359);
nand U10736 (N_10736,N_10372,N_10291);
and U10737 (N_10737,N_10016,N_10305);
or U10738 (N_10738,N_9903,N_9941);
nand U10739 (N_10739,N_10034,N_10241);
and U10740 (N_10740,N_9902,N_10124);
xnor U10741 (N_10741,N_9947,N_10064);
xnor U10742 (N_10742,N_10188,N_10009);
and U10743 (N_10743,N_9863,N_9711);
or U10744 (N_10744,N_10382,N_9659);
nand U10745 (N_10745,N_10166,N_10051);
and U10746 (N_10746,N_10366,N_9995);
nand U10747 (N_10747,N_10255,N_10085);
nor U10748 (N_10748,N_10011,N_10027);
or U10749 (N_10749,N_9699,N_10074);
xnor U10750 (N_10750,N_10121,N_10388);
nor U10751 (N_10751,N_9785,N_9770);
and U10752 (N_10752,N_9665,N_10054);
nand U10753 (N_10753,N_9604,N_10210);
nand U10754 (N_10754,N_9920,N_10078);
nor U10755 (N_10755,N_10071,N_10117);
xor U10756 (N_10756,N_10383,N_10045);
nand U10757 (N_10757,N_9943,N_9830);
xor U10758 (N_10758,N_10163,N_9826);
nand U10759 (N_10759,N_9674,N_9934);
nand U10760 (N_10760,N_10333,N_9973);
or U10761 (N_10761,N_10362,N_10301);
nor U10762 (N_10762,N_9726,N_10322);
nand U10763 (N_10763,N_10172,N_10251);
nand U10764 (N_10764,N_9645,N_9904);
xor U10765 (N_10765,N_9817,N_10225);
and U10766 (N_10766,N_10307,N_9968);
nor U10767 (N_10767,N_10310,N_10052);
xnor U10768 (N_10768,N_9971,N_10364);
or U10769 (N_10769,N_9949,N_9693);
nor U10770 (N_10770,N_9791,N_10218);
or U10771 (N_10771,N_10170,N_9978);
and U10772 (N_10772,N_9972,N_10236);
nor U10773 (N_10773,N_10202,N_10159);
xor U10774 (N_10774,N_10282,N_10330);
xor U10775 (N_10775,N_10384,N_9851);
nand U10776 (N_10776,N_10031,N_10108);
and U10777 (N_10777,N_10227,N_9644);
nor U10778 (N_10778,N_9634,N_10370);
nand U10779 (N_10779,N_10106,N_9976);
or U10780 (N_10780,N_9774,N_9987);
or U10781 (N_10781,N_10091,N_9660);
nand U10782 (N_10782,N_9879,N_10150);
xor U10783 (N_10783,N_9907,N_9832);
and U10784 (N_10784,N_9957,N_10012);
xnor U10785 (N_10785,N_10320,N_9926);
nand U10786 (N_10786,N_9778,N_9737);
nand U10787 (N_10787,N_9784,N_9694);
nand U10788 (N_10788,N_10270,N_10018);
and U10789 (N_10789,N_9929,N_10197);
nor U10790 (N_10790,N_10299,N_10206);
nor U10791 (N_10791,N_9669,N_10179);
nand U10792 (N_10792,N_10347,N_9808);
xor U10793 (N_10793,N_10032,N_10338);
and U10794 (N_10794,N_9682,N_10373);
xnor U10795 (N_10795,N_9722,N_9908);
nor U10796 (N_10796,N_9927,N_9843);
nor U10797 (N_10797,N_10088,N_10356);
xor U10798 (N_10798,N_10090,N_10182);
xor U10799 (N_10799,N_9677,N_10339);
xnor U10800 (N_10800,N_10392,N_9919);
and U10801 (N_10801,N_9996,N_9779);
nor U10802 (N_10802,N_10087,N_10274);
nor U10803 (N_10803,N_10164,N_10142);
or U10804 (N_10804,N_9705,N_9978);
or U10805 (N_10805,N_10134,N_10267);
nand U10806 (N_10806,N_9848,N_9820);
and U10807 (N_10807,N_10093,N_9651);
xnor U10808 (N_10808,N_9735,N_10068);
or U10809 (N_10809,N_9800,N_10041);
or U10810 (N_10810,N_10096,N_10167);
or U10811 (N_10811,N_10189,N_10011);
and U10812 (N_10812,N_10331,N_9607);
and U10813 (N_10813,N_9758,N_10088);
or U10814 (N_10814,N_9687,N_9740);
xnor U10815 (N_10815,N_9604,N_9805);
nor U10816 (N_10816,N_10266,N_9695);
nand U10817 (N_10817,N_10380,N_10190);
xnor U10818 (N_10818,N_9704,N_10090);
nand U10819 (N_10819,N_9901,N_9758);
nor U10820 (N_10820,N_9989,N_9885);
nor U10821 (N_10821,N_9786,N_10284);
and U10822 (N_10822,N_10238,N_10183);
or U10823 (N_10823,N_9942,N_10034);
nor U10824 (N_10824,N_9824,N_9732);
or U10825 (N_10825,N_10308,N_10200);
and U10826 (N_10826,N_9864,N_9757);
and U10827 (N_10827,N_9694,N_9885);
nand U10828 (N_10828,N_10033,N_10197);
nor U10829 (N_10829,N_10082,N_10196);
and U10830 (N_10830,N_10317,N_9853);
and U10831 (N_10831,N_9844,N_9619);
nand U10832 (N_10832,N_9803,N_10328);
nand U10833 (N_10833,N_10222,N_9704);
xnor U10834 (N_10834,N_9809,N_9890);
nor U10835 (N_10835,N_9727,N_10296);
nand U10836 (N_10836,N_10157,N_10268);
and U10837 (N_10837,N_10069,N_9982);
nand U10838 (N_10838,N_10086,N_9998);
or U10839 (N_10839,N_9803,N_9779);
or U10840 (N_10840,N_9649,N_10399);
nor U10841 (N_10841,N_9922,N_9942);
nand U10842 (N_10842,N_10025,N_9620);
or U10843 (N_10843,N_10344,N_9989);
and U10844 (N_10844,N_9682,N_10092);
nand U10845 (N_10845,N_9885,N_10162);
nor U10846 (N_10846,N_10262,N_10030);
and U10847 (N_10847,N_10235,N_10146);
nand U10848 (N_10848,N_9837,N_9720);
and U10849 (N_10849,N_10024,N_9888);
or U10850 (N_10850,N_10307,N_10301);
or U10851 (N_10851,N_9681,N_10132);
nor U10852 (N_10852,N_10099,N_10320);
xor U10853 (N_10853,N_9700,N_9686);
nor U10854 (N_10854,N_10312,N_9827);
or U10855 (N_10855,N_10133,N_9709);
and U10856 (N_10856,N_9633,N_10292);
or U10857 (N_10857,N_9720,N_9986);
nor U10858 (N_10858,N_9870,N_9600);
nor U10859 (N_10859,N_10357,N_10171);
nand U10860 (N_10860,N_9781,N_9853);
or U10861 (N_10861,N_9942,N_10220);
and U10862 (N_10862,N_10152,N_10289);
and U10863 (N_10863,N_10243,N_9693);
nand U10864 (N_10864,N_9903,N_9878);
nand U10865 (N_10865,N_9753,N_9614);
nand U10866 (N_10866,N_9649,N_9646);
nand U10867 (N_10867,N_10120,N_9810);
nor U10868 (N_10868,N_10247,N_10230);
nand U10869 (N_10869,N_9933,N_9998);
xor U10870 (N_10870,N_10011,N_9890);
xor U10871 (N_10871,N_10011,N_9799);
or U10872 (N_10872,N_10151,N_9808);
nor U10873 (N_10873,N_10378,N_10129);
nor U10874 (N_10874,N_9997,N_10196);
and U10875 (N_10875,N_9773,N_10095);
xor U10876 (N_10876,N_9679,N_10330);
and U10877 (N_10877,N_10136,N_9885);
nor U10878 (N_10878,N_9891,N_10292);
nand U10879 (N_10879,N_10028,N_9609);
nor U10880 (N_10880,N_10349,N_10140);
and U10881 (N_10881,N_10074,N_10047);
and U10882 (N_10882,N_9694,N_9628);
and U10883 (N_10883,N_9883,N_10055);
or U10884 (N_10884,N_9607,N_10230);
nor U10885 (N_10885,N_10010,N_10291);
and U10886 (N_10886,N_9999,N_10341);
nor U10887 (N_10887,N_9651,N_10016);
nand U10888 (N_10888,N_9775,N_9732);
xor U10889 (N_10889,N_10140,N_10058);
nor U10890 (N_10890,N_10247,N_10331);
nand U10891 (N_10891,N_10160,N_9931);
nor U10892 (N_10892,N_9948,N_10396);
xor U10893 (N_10893,N_10380,N_9622);
and U10894 (N_10894,N_10348,N_9735);
xor U10895 (N_10895,N_10369,N_9844);
and U10896 (N_10896,N_10080,N_9759);
or U10897 (N_10897,N_10132,N_10330);
nand U10898 (N_10898,N_9667,N_9872);
xor U10899 (N_10899,N_10065,N_10256);
nor U10900 (N_10900,N_10245,N_10326);
and U10901 (N_10901,N_9656,N_9778);
and U10902 (N_10902,N_9706,N_9910);
and U10903 (N_10903,N_10184,N_9879);
nor U10904 (N_10904,N_9872,N_9977);
nand U10905 (N_10905,N_9626,N_10253);
nand U10906 (N_10906,N_9664,N_9682);
xnor U10907 (N_10907,N_10145,N_10393);
or U10908 (N_10908,N_10261,N_9910);
nand U10909 (N_10909,N_9779,N_9862);
nand U10910 (N_10910,N_9891,N_10230);
nor U10911 (N_10911,N_9786,N_9632);
nor U10912 (N_10912,N_10367,N_9739);
or U10913 (N_10913,N_9774,N_10398);
xor U10914 (N_10914,N_9974,N_10294);
or U10915 (N_10915,N_9773,N_10280);
nand U10916 (N_10916,N_9834,N_10396);
nand U10917 (N_10917,N_9842,N_10086);
and U10918 (N_10918,N_10301,N_9664);
nor U10919 (N_10919,N_10116,N_10033);
and U10920 (N_10920,N_10101,N_10197);
nand U10921 (N_10921,N_10057,N_10069);
or U10922 (N_10922,N_10138,N_10035);
nand U10923 (N_10923,N_9707,N_10249);
xnor U10924 (N_10924,N_10039,N_9934);
xor U10925 (N_10925,N_10287,N_10075);
nor U10926 (N_10926,N_10042,N_9712);
nand U10927 (N_10927,N_9904,N_9737);
nor U10928 (N_10928,N_9869,N_9640);
nor U10929 (N_10929,N_9964,N_10203);
or U10930 (N_10930,N_10031,N_10379);
and U10931 (N_10931,N_9973,N_9705);
and U10932 (N_10932,N_10366,N_10018);
nand U10933 (N_10933,N_9749,N_10262);
xnor U10934 (N_10934,N_9838,N_10298);
and U10935 (N_10935,N_9883,N_9729);
and U10936 (N_10936,N_9722,N_10076);
nand U10937 (N_10937,N_10228,N_10339);
xor U10938 (N_10938,N_10311,N_10260);
or U10939 (N_10939,N_10232,N_9972);
nor U10940 (N_10940,N_10207,N_9930);
nand U10941 (N_10941,N_9800,N_9723);
nand U10942 (N_10942,N_9824,N_9662);
nor U10943 (N_10943,N_10018,N_10344);
xnor U10944 (N_10944,N_10066,N_10356);
xor U10945 (N_10945,N_9788,N_9634);
nor U10946 (N_10946,N_10162,N_10062);
nand U10947 (N_10947,N_10082,N_9840);
or U10948 (N_10948,N_10303,N_9967);
or U10949 (N_10949,N_9779,N_9669);
xor U10950 (N_10950,N_10221,N_10269);
and U10951 (N_10951,N_10389,N_10026);
and U10952 (N_10952,N_10230,N_9799);
or U10953 (N_10953,N_10282,N_9932);
and U10954 (N_10954,N_9722,N_9690);
nand U10955 (N_10955,N_9999,N_9781);
nor U10956 (N_10956,N_10335,N_10186);
nand U10957 (N_10957,N_10046,N_10245);
or U10958 (N_10958,N_9767,N_10078);
or U10959 (N_10959,N_9789,N_10302);
and U10960 (N_10960,N_10115,N_9604);
nand U10961 (N_10961,N_10184,N_10037);
xnor U10962 (N_10962,N_10175,N_10193);
nor U10963 (N_10963,N_10351,N_9647);
xnor U10964 (N_10964,N_9914,N_10009);
and U10965 (N_10965,N_10275,N_10322);
or U10966 (N_10966,N_9668,N_9661);
nand U10967 (N_10967,N_9653,N_9775);
or U10968 (N_10968,N_10087,N_10209);
nand U10969 (N_10969,N_10391,N_9660);
xnor U10970 (N_10970,N_10223,N_9825);
or U10971 (N_10971,N_9878,N_9634);
and U10972 (N_10972,N_10325,N_10278);
nand U10973 (N_10973,N_10293,N_9600);
nand U10974 (N_10974,N_9829,N_10372);
nand U10975 (N_10975,N_10194,N_9784);
nor U10976 (N_10976,N_10092,N_9755);
xor U10977 (N_10977,N_10276,N_10027);
or U10978 (N_10978,N_10010,N_10323);
xnor U10979 (N_10979,N_10044,N_10062);
and U10980 (N_10980,N_10334,N_9785);
or U10981 (N_10981,N_10332,N_10399);
xnor U10982 (N_10982,N_9909,N_9752);
and U10983 (N_10983,N_10331,N_10233);
and U10984 (N_10984,N_10357,N_9911);
and U10985 (N_10985,N_10322,N_9658);
xor U10986 (N_10986,N_9960,N_9935);
or U10987 (N_10987,N_9904,N_10021);
nand U10988 (N_10988,N_9608,N_10163);
nor U10989 (N_10989,N_10076,N_9880);
nand U10990 (N_10990,N_9651,N_10353);
and U10991 (N_10991,N_9760,N_9695);
nand U10992 (N_10992,N_10039,N_10056);
or U10993 (N_10993,N_9895,N_10330);
nand U10994 (N_10994,N_9918,N_9722);
nor U10995 (N_10995,N_9837,N_9849);
and U10996 (N_10996,N_10020,N_9719);
nand U10997 (N_10997,N_10332,N_10092);
xnor U10998 (N_10998,N_10266,N_9920);
xor U10999 (N_10999,N_10087,N_10261);
xnor U11000 (N_11000,N_10196,N_9886);
xnor U11001 (N_11001,N_9803,N_10086);
or U11002 (N_11002,N_10020,N_10350);
xnor U11003 (N_11003,N_9704,N_9660);
nand U11004 (N_11004,N_10211,N_9757);
nand U11005 (N_11005,N_9728,N_10252);
and U11006 (N_11006,N_9909,N_10253);
xnor U11007 (N_11007,N_9678,N_10224);
nor U11008 (N_11008,N_10327,N_9833);
nand U11009 (N_11009,N_9848,N_10001);
nor U11010 (N_11010,N_9615,N_10320);
and U11011 (N_11011,N_10143,N_10199);
and U11012 (N_11012,N_10102,N_9659);
nand U11013 (N_11013,N_10366,N_10079);
nor U11014 (N_11014,N_9793,N_9833);
xnor U11015 (N_11015,N_9757,N_10022);
and U11016 (N_11016,N_9793,N_10034);
xnor U11017 (N_11017,N_10349,N_10134);
xor U11018 (N_11018,N_10181,N_9734);
nand U11019 (N_11019,N_10118,N_9840);
xnor U11020 (N_11020,N_10288,N_9685);
and U11021 (N_11021,N_9678,N_10278);
xnor U11022 (N_11022,N_10148,N_10212);
xnor U11023 (N_11023,N_10260,N_10046);
nand U11024 (N_11024,N_10000,N_10117);
nand U11025 (N_11025,N_9865,N_9935);
or U11026 (N_11026,N_9846,N_9817);
and U11027 (N_11027,N_9676,N_10108);
xor U11028 (N_11028,N_9782,N_9637);
or U11029 (N_11029,N_9951,N_10100);
xor U11030 (N_11030,N_10152,N_10155);
xnor U11031 (N_11031,N_10094,N_9630);
nand U11032 (N_11032,N_9728,N_9683);
or U11033 (N_11033,N_10031,N_9843);
nand U11034 (N_11034,N_10294,N_10219);
nor U11035 (N_11035,N_9613,N_10240);
or U11036 (N_11036,N_10234,N_9888);
and U11037 (N_11037,N_10006,N_10154);
xor U11038 (N_11038,N_9953,N_10367);
nand U11039 (N_11039,N_10081,N_9767);
or U11040 (N_11040,N_10223,N_10278);
and U11041 (N_11041,N_10389,N_10134);
or U11042 (N_11042,N_9750,N_10192);
nor U11043 (N_11043,N_10208,N_10337);
or U11044 (N_11044,N_10148,N_9994);
nand U11045 (N_11045,N_10302,N_9999);
nor U11046 (N_11046,N_9949,N_9701);
nor U11047 (N_11047,N_9811,N_10254);
nor U11048 (N_11048,N_10180,N_10359);
and U11049 (N_11049,N_9897,N_10143);
nor U11050 (N_11050,N_9812,N_9941);
or U11051 (N_11051,N_9758,N_9743);
or U11052 (N_11052,N_9734,N_9945);
nor U11053 (N_11053,N_9969,N_9637);
and U11054 (N_11054,N_10341,N_10022);
nand U11055 (N_11055,N_9783,N_10160);
nor U11056 (N_11056,N_10237,N_9791);
nor U11057 (N_11057,N_9979,N_10206);
and U11058 (N_11058,N_9634,N_10133);
or U11059 (N_11059,N_9691,N_9905);
nor U11060 (N_11060,N_10320,N_10228);
and U11061 (N_11061,N_9713,N_10394);
nand U11062 (N_11062,N_9964,N_9991);
nor U11063 (N_11063,N_9619,N_9780);
or U11064 (N_11064,N_10235,N_10013);
or U11065 (N_11065,N_10203,N_9725);
or U11066 (N_11066,N_9614,N_10003);
xor U11067 (N_11067,N_10122,N_9633);
nand U11068 (N_11068,N_9857,N_10285);
nand U11069 (N_11069,N_10149,N_9653);
and U11070 (N_11070,N_10091,N_10233);
or U11071 (N_11071,N_9795,N_10031);
or U11072 (N_11072,N_10271,N_9661);
or U11073 (N_11073,N_10238,N_9949);
nand U11074 (N_11074,N_9924,N_9672);
nor U11075 (N_11075,N_10000,N_10089);
or U11076 (N_11076,N_9835,N_10085);
and U11077 (N_11077,N_10003,N_10237);
xnor U11078 (N_11078,N_9807,N_10166);
nor U11079 (N_11079,N_10297,N_9738);
nand U11080 (N_11080,N_9855,N_10174);
or U11081 (N_11081,N_10085,N_10348);
nor U11082 (N_11082,N_10135,N_9882);
nand U11083 (N_11083,N_10317,N_10054);
nand U11084 (N_11084,N_9820,N_9776);
and U11085 (N_11085,N_9697,N_10327);
xor U11086 (N_11086,N_9775,N_9995);
xnor U11087 (N_11087,N_9875,N_9869);
and U11088 (N_11088,N_9964,N_10307);
xor U11089 (N_11089,N_9952,N_9810);
nand U11090 (N_11090,N_9981,N_9782);
and U11091 (N_11091,N_10108,N_10238);
and U11092 (N_11092,N_10115,N_10018);
nand U11093 (N_11093,N_9942,N_9648);
and U11094 (N_11094,N_10247,N_10212);
and U11095 (N_11095,N_10392,N_10149);
and U11096 (N_11096,N_9919,N_10321);
and U11097 (N_11097,N_10139,N_9653);
or U11098 (N_11098,N_9913,N_9866);
nand U11099 (N_11099,N_10374,N_10139);
nand U11100 (N_11100,N_9743,N_10334);
and U11101 (N_11101,N_9684,N_9885);
nor U11102 (N_11102,N_9615,N_10322);
and U11103 (N_11103,N_10154,N_10248);
xnor U11104 (N_11104,N_10079,N_9793);
nand U11105 (N_11105,N_10145,N_9909);
nand U11106 (N_11106,N_9759,N_9676);
nand U11107 (N_11107,N_9722,N_9745);
and U11108 (N_11108,N_10017,N_9860);
xnor U11109 (N_11109,N_10376,N_9657);
nand U11110 (N_11110,N_10316,N_9765);
xnor U11111 (N_11111,N_10082,N_9620);
nand U11112 (N_11112,N_10340,N_10358);
and U11113 (N_11113,N_9822,N_9767);
and U11114 (N_11114,N_9814,N_9790);
nor U11115 (N_11115,N_10226,N_10131);
nor U11116 (N_11116,N_10000,N_10036);
or U11117 (N_11117,N_9967,N_10320);
or U11118 (N_11118,N_10225,N_10391);
or U11119 (N_11119,N_9725,N_10093);
nor U11120 (N_11120,N_9885,N_9822);
and U11121 (N_11121,N_10014,N_10167);
xor U11122 (N_11122,N_10150,N_9803);
or U11123 (N_11123,N_10066,N_10206);
xor U11124 (N_11124,N_10387,N_10180);
nand U11125 (N_11125,N_9975,N_9678);
or U11126 (N_11126,N_9635,N_9967);
nor U11127 (N_11127,N_9833,N_10068);
nor U11128 (N_11128,N_9717,N_10340);
and U11129 (N_11129,N_9710,N_10220);
xor U11130 (N_11130,N_10058,N_9840);
or U11131 (N_11131,N_9800,N_9984);
nand U11132 (N_11132,N_10276,N_10109);
xor U11133 (N_11133,N_10059,N_9851);
or U11134 (N_11134,N_9996,N_10066);
nand U11135 (N_11135,N_10272,N_9890);
xnor U11136 (N_11136,N_10221,N_9738);
or U11137 (N_11137,N_9622,N_9605);
nand U11138 (N_11138,N_9828,N_10211);
xnor U11139 (N_11139,N_9846,N_10114);
nand U11140 (N_11140,N_10226,N_9978);
and U11141 (N_11141,N_9647,N_9812);
nor U11142 (N_11142,N_10321,N_10207);
nor U11143 (N_11143,N_10035,N_10327);
or U11144 (N_11144,N_9600,N_9810);
and U11145 (N_11145,N_10370,N_10020);
nor U11146 (N_11146,N_9941,N_10261);
nor U11147 (N_11147,N_9775,N_9766);
xnor U11148 (N_11148,N_10025,N_10204);
and U11149 (N_11149,N_9908,N_10212);
nor U11150 (N_11150,N_10193,N_9998);
nand U11151 (N_11151,N_10394,N_9742);
and U11152 (N_11152,N_10331,N_10323);
or U11153 (N_11153,N_9729,N_10082);
nand U11154 (N_11154,N_10097,N_9805);
xor U11155 (N_11155,N_10241,N_10371);
xor U11156 (N_11156,N_9682,N_10302);
nor U11157 (N_11157,N_10044,N_9963);
nor U11158 (N_11158,N_10346,N_10120);
xnor U11159 (N_11159,N_10148,N_9705);
nand U11160 (N_11160,N_9986,N_9768);
or U11161 (N_11161,N_10043,N_9626);
nand U11162 (N_11162,N_9701,N_10367);
or U11163 (N_11163,N_9827,N_10177);
or U11164 (N_11164,N_9901,N_9883);
and U11165 (N_11165,N_9937,N_9794);
or U11166 (N_11166,N_9757,N_10030);
or U11167 (N_11167,N_10180,N_9653);
nor U11168 (N_11168,N_9805,N_9631);
nand U11169 (N_11169,N_10357,N_10341);
xnor U11170 (N_11170,N_9773,N_10172);
or U11171 (N_11171,N_9856,N_10189);
nor U11172 (N_11172,N_9699,N_9856);
nor U11173 (N_11173,N_10302,N_10016);
nand U11174 (N_11174,N_10268,N_9876);
xor U11175 (N_11175,N_9848,N_9899);
nor U11176 (N_11176,N_9946,N_9745);
xnor U11177 (N_11177,N_10143,N_9959);
nand U11178 (N_11178,N_10046,N_10113);
and U11179 (N_11179,N_9641,N_10285);
nand U11180 (N_11180,N_9995,N_10192);
nor U11181 (N_11181,N_9718,N_9948);
nor U11182 (N_11182,N_10344,N_10105);
xor U11183 (N_11183,N_9874,N_10017);
or U11184 (N_11184,N_10281,N_9789);
and U11185 (N_11185,N_9994,N_9834);
nand U11186 (N_11186,N_10180,N_9720);
or U11187 (N_11187,N_10212,N_9777);
nor U11188 (N_11188,N_10090,N_10322);
or U11189 (N_11189,N_10077,N_10131);
and U11190 (N_11190,N_9848,N_9946);
or U11191 (N_11191,N_10266,N_10058);
or U11192 (N_11192,N_9993,N_10267);
nand U11193 (N_11193,N_9875,N_9938);
nand U11194 (N_11194,N_9735,N_10122);
xnor U11195 (N_11195,N_9914,N_10047);
xor U11196 (N_11196,N_9956,N_10370);
and U11197 (N_11197,N_9847,N_10170);
xor U11198 (N_11198,N_9940,N_10261);
and U11199 (N_11199,N_9921,N_10253);
nor U11200 (N_11200,N_10698,N_10904);
and U11201 (N_11201,N_10605,N_10878);
nor U11202 (N_11202,N_11125,N_11075);
or U11203 (N_11203,N_10990,N_10480);
nand U11204 (N_11204,N_11098,N_10812);
nand U11205 (N_11205,N_10665,N_10838);
or U11206 (N_11206,N_10942,N_11128);
and U11207 (N_11207,N_10500,N_10765);
xnor U11208 (N_11208,N_10711,N_11057);
or U11209 (N_11209,N_10464,N_10481);
or U11210 (N_11210,N_10702,N_11077);
nor U11211 (N_11211,N_10685,N_10503);
and U11212 (N_11212,N_10652,N_10954);
nor U11213 (N_11213,N_10771,N_10463);
or U11214 (N_11214,N_10508,N_10431);
nand U11215 (N_11215,N_10993,N_10417);
or U11216 (N_11216,N_10517,N_10419);
nor U11217 (N_11217,N_11005,N_10400);
and U11218 (N_11218,N_10738,N_10655);
and U11219 (N_11219,N_10582,N_11099);
and U11220 (N_11220,N_10424,N_10509);
xor U11221 (N_11221,N_10718,N_11161);
nor U11222 (N_11222,N_10430,N_10830);
nand U11223 (N_11223,N_11082,N_11089);
nand U11224 (N_11224,N_10604,N_10985);
xnor U11225 (N_11225,N_10953,N_10476);
nand U11226 (N_11226,N_10567,N_11136);
and U11227 (N_11227,N_10518,N_11110);
xnor U11228 (N_11228,N_10930,N_10811);
xor U11229 (N_11229,N_10872,N_11011);
or U11230 (N_11230,N_10641,N_10760);
nor U11231 (N_11231,N_11015,N_10998);
xor U11232 (N_11232,N_11035,N_10465);
and U11233 (N_11233,N_11156,N_10447);
xor U11234 (N_11234,N_10752,N_10704);
nand U11235 (N_11235,N_10853,N_10681);
and U11236 (N_11236,N_11080,N_10809);
and U11237 (N_11237,N_10630,N_10799);
xor U11238 (N_11238,N_10519,N_10826);
nor U11239 (N_11239,N_10624,N_11032);
nor U11240 (N_11240,N_10579,N_11107);
and U11241 (N_11241,N_10468,N_10891);
nand U11242 (N_11242,N_10403,N_10541);
and U11243 (N_11243,N_10761,N_11086);
nand U11244 (N_11244,N_10461,N_11046);
nor U11245 (N_11245,N_10742,N_10848);
xor U11246 (N_11246,N_10627,N_10987);
nor U11247 (N_11247,N_10492,N_10550);
and U11248 (N_11248,N_10635,N_10662);
or U11249 (N_11249,N_11149,N_10610);
nor U11250 (N_11250,N_10535,N_10868);
or U11251 (N_11251,N_10865,N_10515);
nor U11252 (N_11252,N_10608,N_10938);
nand U11253 (N_11253,N_10510,N_11164);
nand U11254 (N_11254,N_10565,N_10625);
or U11255 (N_11255,N_11040,N_11093);
nor U11256 (N_11256,N_10789,N_10974);
nand U11257 (N_11257,N_11143,N_11070);
nand U11258 (N_11258,N_11103,N_11190);
and U11259 (N_11259,N_11023,N_11150);
or U11260 (N_11260,N_10725,N_11183);
and U11261 (N_11261,N_10777,N_10912);
xor U11262 (N_11262,N_11002,N_10745);
nor U11263 (N_11263,N_10860,N_11014);
nand U11264 (N_11264,N_10467,N_11083);
or U11265 (N_11265,N_10970,N_10963);
nand U11266 (N_11266,N_10679,N_10831);
or U11267 (N_11267,N_10670,N_10902);
or U11268 (N_11268,N_10824,N_10941);
and U11269 (N_11269,N_11101,N_10571);
xor U11270 (N_11270,N_10629,N_10678);
xnor U11271 (N_11271,N_10975,N_10653);
xnor U11272 (N_11272,N_11199,N_10421);
or U11273 (N_11273,N_11165,N_11071);
or U11274 (N_11274,N_10986,N_10639);
and U11275 (N_11275,N_10996,N_10566);
and U11276 (N_11276,N_10805,N_10631);
nand U11277 (N_11277,N_11117,N_11142);
or U11278 (N_11278,N_10611,N_11012);
nor U11279 (N_11279,N_10844,N_10818);
nor U11280 (N_11280,N_10731,N_10802);
nor U11281 (N_11281,N_10514,N_10893);
or U11282 (N_11282,N_10800,N_10527);
and U11283 (N_11283,N_10798,N_11187);
and U11284 (N_11284,N_10581,N_10790);
nor U11285 (N_11285,N_10505,N_10645);
nand U11286 (N_11286,N_10699,N_11073);
and U11287 (N_11287,N_10788,N_10660);
or U11288 (N_11288,N_10683,N_10412);
xor U11289 (N_11289,N_11124,N_10956);
nor U11290 (N_11290,N_10516,N_11132);
nor U11291 (N_11291,N_11042,N_10563);
or U11292 (N_11292,N_10433,N_10593);
and U11293 (N_11293,N_10948,N_10422);
nor U11294 (N_11294,N_10825,N_10739);
and U11295 (N_11295,N_10506,N_10766);
and U11296 (N_11296,N_10928,N_10531);
nor U11297 (N_11297,N_10855,N_10889);
xnor U11298 (N_11298,N_10493,N_10892);
xnor U11299 (N_11299,N_10846,N_10915);
xnor U11300 (N_11300,N_11196,N_10806);
xor U11301 (N_11301,N_10816,N_10404);
and U11302 (N_11302,N_11028,N_10471);
or U11303 (N_11303,N_10594,N_11048);
xor U11304 (N_11304,N_11105,N_10602);
or U11305 (N_11305,N_10905,N_11176);
and U11306 (N_11306,N_10744,N_11139);
and U11307 (N_11307,N_11044,N_10874);
nor U11308 (N_11308,N_11109,N_10896);
nand U11309 (N_11309,N_10871,N_10950);
xnor U11310 (N_11310,N_10494,N_10512);
nand U11311 (N_11311,N_10646,N_10551);
xnor U11312 (N_11312,N_11188,N_11100);
nand U11313 (N_11313,N_10663,N_10768);
or U11314 (N_11314,N_10852,N_10589);
and U11315 (N_11315,N_11106,N_11154);
or U11316 (N_11316,N_10944,N_10561);
or U11317 (N_11317,N_10438,N_11181);
xnor U11318 (N_11318,N_10729,N_11084);
nor U11319 (N_11319,N_10960,N_10982);
nand U11320 (N_11320,N_10601,N_10887);
xor U11321 (N_11321,N_10837,N_10600);
and U11322 (N_11322,N_11041,N_11174);
xnor U11323 (N_11323,N_11198,N_10995);
nor U11324 (N_11324,N_10929,N_10451);
and U11325 (N_11325,N_10882,N_10524);
nor U11326 (N_11326,N_10445,N_10910);
nor U11327 (N_11327,N_10885,N_10972);
or U11328 (N_11328,N_10586,N_10857);
xnor U11329 (N_11329,N_11160,N_10688);
or U11330 (N_11330,N_10898,N_10815);
nand U11331 (N_11331,N_10674,N_10906);
xor U11332 (N_11332,N_10499,N_10797);
xor U11333 (N_11333,N_10709,N_10703);
nor U11334 (N_11334,N_10967,N_10978);
or U11335 (N_11335,N_10443,N_10934);
nor U11336 (N_11336,N_11153,N_11001);
xnor U11337 (N_11337,N_11025,N_10714);
xnor U11338 (N_11338,N_10764,N_10979);
nor U11339 (N_11339,N_10875,N_11177);
nor U11340 (N_11340,N_10903,N_11064);
or U11341 (N_11341,N_10574,N_10772);
nor U11342 (N_11342,N_10648,N_10657);
xor U11343 (N_11343,N_11115,N_10854);
nand U11344 (N_11344,N_10521,N_10522);
nor U11345 (N_11345,N_10827,N_11173);
nor U11346 (N_11346,N_10437,N_10769);
and U11347 (N_11347,N_10988,N_10801);
nand U11348 (N_11348,N_10708,N_11022);
or U11349 (N_11349,N_10425,N_11078);
xnor U11350 (N_11350,N_10661,N_10917);
nand U11351 (N_11351,N_11058,N_10459);
or U11352 (N_11352,N_10763,N_11147);
xor U11353 (N_11353,N_10444,N_11144);
nand U11354 (N_11354,N_10585,N_11004);
and U11355 (N_11355,N_10723,N_10472);
nand U11356 (N_11356,N_10836,N_11189);
xor U11357 (N_11357,N_10862,N_10697);
or U11358 (N_11358,N_10534,N_10640);
nor U11359 (N_11359,N_10814,N_10997);
xor U11360 (N_11360,N_10749,N_10864);
nor U11361 (N_11361,N_11138,N_10794);
xnor U11362 (N_11362,N_10823,N_10817);
or U11363 (N_11363,N_10754,N_11079);
nor U11364 (N_11364,N_10787,N_10617);
or U11365 (N_11365,N_10453,N_10529);
xnor U11366 (N_11366,N_10957,N_10520);
or U11367 (N_11367,N_10775,N_10488);
and U11368 (N_11368,N_10402,N_10539);
and U11369 (N_11369,N_10446,N_10575);
xnor U11370 (N_11370,N_10785,N_11137);
and U11371 (N_11371,N_10927,N_10435);
and U11372 (N_11372,N_11087,N_10682);
nor U11373 (N_11373,N_10947,N_10926);
nor U11374 (N_11374,N_11067,N_11059);
and U11375 (N_11375,N_10733,N_11172);
nor U11376 (N_11376,N_10958,N_10606);
xor U11377 (N_11377,N_11088,N_10969);
xor U11378 (N_11378,N_10897,N_10556);
or U11379 (N_11379,N_10717,N_10867);
and U11380 (N_11380,N_10925,N_11027);
and U11381 (N_11381,N_10691,N_11090);
and U11382 (N_11382,N_11121,N_10621);
or U11383 (N_11383,N_11158,N_10884);
and U11384 (N_11384,N_10628,N_11116);
nand U11385 (N_11385,N_10618,N_10548);
or U11386 (N_11386,N_10965,N_10992);
nor U11387 (N_11387,N_10793,N_10828);
and U11388 (N_11388,N_11030,N_10440);
nor U11389 (N_11389,N_10921,N_10686);
or U11390 (N_11390,N_11031,N_10914);
and U11391 (N_11391,N_10866,N_10724);
xnor U11392 (N_11392,N_11013,N_10961);
nor U11393 (N_11393,N_10540,N_10507);
xor U11394 (N_11394,N_10513,N_11074);
or U11395 (N_11395,N_10473,N_10588);
or U11396 (N_11396,N_10533,N_10423);
or U11397 (N_11397,N_11182,N_11047);
or U11398 (N_11398,N_10572,N_11127);
and U11399 (N_11399,N_10498,N_11056);
nor U11400 (N_11400,N_10578,N_10411);
nand U11401 (N_11401,N_10707,N_10780);
and U11402 (N_11402,N_10501,N_10644);
and U11403 (N_11403,N_10804,N_11113);
nor U11404 (N_11404,N_10900,N_10877);
and U11405 (N_11405,N_10543,N_10973);
and U11406 (N_11406,N_10487,N_10647);
nor U11407 (N_11407,N_10770,N_10414);
or U11408 (N_11408,N_11063,N_10450);
nand U11409 (N_11409,N_10418,N_11085);
nor U11410 (N_11410,N_10710,N_10747);
nand U11411 (N_11411,N_10560,N_10803);
and U11412 (N_11412,N_10881,N_10614);
and U11413 (N_11413,N_10615,N_10939);
or U11414 (N_11414,N_10672,N_10455);
or U11415 (N_11415,N_10408,N_10791);
xnor U11416 (N_11416,N_11197,N_10470);
nor U11417 (N_11417,N_10952,N_11191);
nor U11418 (N_11418,N_11166,N_10913);
nand U11419 (N_11419,N_10547,N_10667);
or U11420 (N_11420,N_10656,N_10796);
xor U11421 (N_11421,N_10649,N_10584);
and U11422 (N_11422,N_10466,N_11186);
and U11423 (N_11423,N_10886,N_10994);
xor U11424 (N_11424,N_11060,N_10564);
nor U11425 (N_11425,N_10580,N_10544);
xor U11426 (N_11426,N_10587,N_10951);
xnor U11427 (N_11427,N_10883,N_10715);
xor U11428 (N_11428,N_11021,N_10847);
or U11429 (N_11429,N_10626,N_11016);
xor U11430 (N_11430,N_10721,N_10719);
nand U11431 (N_11431,N_11134,N_11111);
or U11432 (N_11432,N_10504,N_10741);
nand U11433 (N_11433,N_10843,N_10762);
nor U11434 (N_11434,N_11102,N_10612);
xnor U11435 (N_11435,N_10479,N_10429);
nor U11436 (N_11436,N_11194,N_10876);
and U11437 (N_11437,N_10642,N_10964);
xor U11438 (N_11438,N_11066,N_10895);
or U11439 (N_11439,N_11062,N_11108);
nand U11440 (N_11440,N_11045,N_10569);
and U11441 (N_11441,N_11018,N_10695);
or U11442 (N_11442,N_10888,N_10623);
or U11443 (N_11443,N_11178,N_10920);
nand U11444 (N_11444,N_10420,N_10595);
and U11445 (N_11445,N_11119,N_11051);
nand U11446 (N_11446,N_10484,N_10442);
nand U11447 (N_11447,N_11112,N_10583);
or U11448 (N_11448,N_10932,N_10962);
or U11449 (N_11449,N_11065,N_10449);
nor U11450 (N_11450,N_10734,N_11010);
nor U11451 (N_11451,N_10619,N_10406);
nor U11452 (N_11452,N_10636,N_10616);
or U11453 (N_11453,N_10880,N_10555);
or U11454 (N_11454,N_11148,N_11003);
or U11455 (N_11455,N_10658,N_11036);
nor U11456 (N_11456,N_10489,N_10553);
nor U11457 (N_11457,N_11126,N_10822);
nand U11458 (N_11458,N_11133,N_10859);
nor U11459 (N_11459,N_10839,N_11180);
xnor U11460 (N_11460,N_10591,N_10532);
nor U11461 (N_11461,N_10863,N_10728);
nor U11462 (N_11462,N_11168,N_11123);
xor U11463 (N_11463,N_11122,N_10901);
nand U11464 (N_11464,N_10552,N_11146);
nand U11465 (N_11465,N_11081,N_10722);
xor U11466 (N_11466,N_10659,N_11092);
nand U11467 (N_11467,N_10654,N_10576);
or U11468 (N_11468,N_10511,N_11114);
and U11469 (N_11469,N_10736,N_11037);
nor U11470 (N_11470,N_10475,N_10673);
nand U11471 (N_11471,N_10907,N_10792);
or U11472 (N_11472,N_10918,N_10810);
or U11473 (N_11473,N_10720,N_10919);
nor U11474 (N_11474,N_10483,N_11000);
nor U11475 (N_11475,N_10869,N_10474);
xor U11476 (N_11476,N_10746,N_10684);
xnor U11477 (N_11477,N_10620,N_11054);
xnor U11478 (N_11478,N_10959,N_10716);
nand U11479 (N_11479,N_10694,N_10977);
nand U11480 (N_11480,N_10966,N_10946);
or U11481 (N_11481,N_10753,N_10783);
nand U11482 (N_11482,N_10457,N_10922);
xnor U11483 (N_11483,N_10633,N_10677);
nand U11484 (N_11484,N_10955,N_10776);
nor U11485 (N_11485,N_10486,N_10482);
nor U11486 (N_11486,N_10607,N_10712);
xnor U11487 (N_11487,N_10401,N_10478);
or U11488 (N_11488,N_11029,N_10427);
xnor U11489 (N_11489,N_10542,N_10405);
xnor U11490 (N_11490,N_10856,N_10456);
or U11491 (N_11491,N_10598,N_10676);
xnor U11492 (N_11492,N_11052,N_11049);
xnor U11493 (N_11493,N_11076,N_10940);
nand U11494 (N_11494,N_10945,N_10554);
and U11495 (N_11495,N_10671,N_11096);
or U11496 (N_11496,N_10497,N_10454);
nor U11497 (N_11497,N_10758,N_10732);
xor U11498 (N_11498,N_10426,N_10701);
xor U11499 (N_11499,N_10525,N_10832);
and U11500 (N_11500,N_10767,N_10664);
nor U11501 (N_11501,N_10779,N_10562);
and U11502 (N_11502,N_10911,N_10858);
and U11503 (N_11503,N_10687,N_10638);
or U11504 (N_11504,N_10757,N_11020);
nand U11505 (N_11505,N_11167,N_10829);
nor U11506 (N_11506,N_10692,N_10546);
nor U11507 (N_11507,N_10784,N_10807);
nand U11508 (N_11508,N_11159,N_10850);
nand U11509 (N_11509,N_10949,N_10413);
xor U11510 (N_11510,N_10439,N_10407);
nor U11511 (N_11511,N_10786,N_11069);
nand U11512 (N_11512,N_10458,N_11175);
nor U11513 (N_11513,N_10462,N_11050);
nand U11514 (N_11514,N_11072,N_10536);
xnor U11515 (N_11515,N_10637,N_10666);
nand U11516 (N_11516,N_10840,N_11195);
or U11517 (N_11517,N_10751,N_10448);
and U11518 (N_11518,N_11104,N_10819);
nor U11519 (N_11519,N_10841,N_10502);
or U11520 (N_11520,N_10980,N_11185);
or U11521 (N_11521,N_11068,N_11162);
or U11522 (N_11522,N_10696,N_10759);
xor U11523 (N_11523,N_11034,N_10890);
nor U11524 (N_11524,N_11145,N_10740);
xnor U11525 (N_11525,N_10689,N_10923);
or U11526 (N_11526,N_10820,N_11094);
nor U11527 (N_11527,N_11009,N_10968);
or U11528 (N_11528,N_11129,N_10669);
or U11529 (N_11529,N_10545,N_10650);
xor U11530 (N_11530,N_10668,N_10774);
nor U11531 (N_11531,N_10726,N_10894);
nand U11532 (N_11532,N_10452,N_10643);
xor U11533 (N_11533,N_10469,N_10909);
nand U11534 (N_11534,N_10713,N_10599);
xor U11535 (N_11535,N_10495,N_10485);
nand U11536 (N_11536,N_10577,N_10409);
xor U11537 (N_11537,N_10808,N_10813);
or U11538 (N_11538,N_10597,N_11135);
and U11539 (N_11539,N_10557,N_10750);
and U11540 (N_11540,N_10526,N_10795);
and U11541 (N_11541,N_10609,N_11155);
and U11542 (N_11542,N_10899,N_11061);
or U11543 (N_11543,N_10705,N_10937);
xnor U11544 (N_11544,N_10730,N_10690);
nor U11545 (N_11545,N_10834,N_10596);
or U11546 (N_11546,N_10976,N_11017);
and U11547 (N_11547,N_10568,N_11007);
nor U11548 (N_11548,N_10849,N_10706);
and U11549 (N_11549,N_10916,N_10537);
nor U11550 (N_11550,N_10821,N_10835);
nand U11551 (N_11551,N_11055,N_11097);
nand U11552 (N_11552,N_11120,N_11130);
nor U11553 (N_11553,N_11091,N_10999);
or U11554 (N_11554,N_11026,N_10851);
nor U11555 (N_11555,N_11024,N_11192);
nor U11556 (N_11556,N_10981,N_10781);
nand U11557 (N_11557,N_10622,N_10441);
nand U11558 (N_11558,N_11184,N_10870);
or U11559 (N_11559,N_10873,N_11131);
xnor U11560 (N_11560,N_10590,N_10727);
xor U11561 (N_11561,N_10743,N_10991);
nor U11562 (N_11562,N_10632,N_10700);
nand U11563 (N_11563,N_10735,N_10434);
and U11564 (N_11564,N_11008,N_10989);
nand U11565 (N_11565,N_10490,N_10549);
and U11566 (N_11566,N_11095,N_11033);
and U11567 (N_11567,N_10570,N_10778);
nand U11568 (N_11568,N_10936,N_11053);
nor U11569 (N_11569,N_10530,N_10943);
nor U11570 (N_11570,N_11038,N_10496);
and U11571 (N_11571,N_10416,N_11152);
nor U11572 (N_11572,N_10971,N_10491);
or U11573 (N_11573,N_10833,N_10675);
or U11574 (N_11574,N_10756,N_10680);
nand U11575 (N_11575,N_10773,N_10613);
nand U11576 (N_11576,N_10573,N_10931);
and U11577 (N_11577,N_10558,N_10477);
and U11578 (N_11578,N_10528,N_10737);
xnor U11579 (N_11579,N_11170,N_10428);
or U11580 (N_11580,N_10748,N_10924);
and U11581 (N_11581,N_10935,N_11179);
xor U11582 (N_11582,N_10559,N_10693);
nand U11583 (N_11583,N_10436,N_11043);
nand U11584 (N_11584,N_10908,N_11193);
xor U11585 (N_11585,N_11171,N_10755);
xor U11586 (N_11586,N_10523,N_10415);
and U11587 (N_11587,N_10842,N_11019);
and U11588 (N_11588,N_10861,N_10460);
and U11589 (N_11589,N_10592,N_11169);
nand U11590 (N_11590,N_10782,N_10634);
nand U11591 (N_11591,N_11140,N_10984);
and U11592 (N_11592,N_11006,N_10410);
or U11593 (N_11593,N_10933,N_10432);
or U11594 (N_11594,N_10845,N_11141);
and U11595 (N_11595,N_11118,N_11151);
nand U11596 (N_11596,N_11163,N_10603);
nor U11597 (N_11597,N_11157,N_10879);
or U11598 (N_11598,N_11039,N_10983);
nor U11599 (N_11599,N_10538,N_10651);
xnor U11600 (N_11600,N_10826,N_11145);
nor U11601 (N_11601,N_10825,N_10994);
or U11602 (N_11602,N_11019,N_10520);
xor U11603 (N_11603,N_10664,N_10984);
nor U11604 (N_11604,N_10829,N_10961);
nand U11605 (N_11605,N_10879,N_10473);
xnor U11606 (N_11606,N_10534,N_10711);
xor U11607 (N_11607,N_10414,N_10420);
or U11608 (N_11608,N_10760,N_10865);
xor U11609 (N_11609,N_10794,N_10747);
nor U11610 (N_11610,N_11144,N_10982);
nor U11611 (N_11611,N_11155,N_11152);
and U11612 (N_11612,N_10844,N_11073);
nand U11613 (N_11613,N_11169,N_10912);
and U11614 (N_11614,N_10964,N_10472);
and U11615 (N_11615,N_10747,N_10585);
or U11616 (N_11616,N_11067,N_11073);
or U11617 (N_11617,N_10895,N_10720);
nor U11618 (N_11618,N_10501,N_11156);
or U11619 (N_11619,N_10451,N_10845);
nand U11620 (N_11620,N_10442,N_10725);
and U11621 (N_11621,N_10875,N_10690);
or U11622 (N_11622,N_11199,N_10669);
and U11623 (N_11623,N_10504,N_10807);
xnor U11624 (N_11624,N_11152,N_10514);
nand U11625 (N_11625,N_10512,N_10422);
and U11626 (N_11626,N_10546,N_10685);
and U11627 (N_11627,N_10472,N_10525);
nand U11628 (N_11628,N_10925,N_10824);
nand U11629 (N_11629,N_11198,N_10928);
nor U11630 (N_11630,N_10921,N_10730);
xnor U11631 (N_11631,N_10706,N_11179);
xnor U11632 (N_11632,N_10631,N_10585);
xor U11633 (N_11633,N_11069,N_10939);
or U11634 (N_11634,N_10652,N_11195);
and U11635 (N_11635,N_11137,N_10815);
nor U11636 (N_11636,N_10875,N_11110);
or U11637 (N_11637,N_10460,N_10913);
xnor U11638 (N_11638,N_10702,N_10754);
and U11639 (N_11639,N_10965,N_10969);
and U11640 (N_11640,N_10839,N_11058);
and U11641 (N_11641,N_11188,N_10468);
nor U11642 (N_11642,N_10733,N_11102);
nor U11643 (N_11643,N_10774,N_10651);
xor U11644 (N_11644,N_10768,N_10499);
nand U11645 (N_11645,N_10546,N_10637);
or U11646 (N_11646,N_10414,N_10888);
nor U11647 (N_11647,N_10529,N_10640);
nand U11648 (N_11648,N_10738,N_11171);
nand U11649 (N_11649,N_11199,N_11131);
xor U11650 (N_11650,N_10420,N_10685);
and U11651 (N_11651,N_10834,N_10643);
or U11652 (N_11652,N_10595,N_10689);
nand U11653 (N_11653,N_10653,N_10488);
nor U11654 (N_11654,N_11022,N_11107);
xor U11655 (N_11655,N_10503,N_11026);
and U11656 (N_11656,N_10513,N_10427);
or U11657 (N_11657,N_10836,N_10490);
nor U11658 (N_11658,N_10561,N_11128);
or U11659 (N_11659,N_10743,N_11004);
xor U11660 (N_11660,N_10878,N_10990);
nand U11661 (N_11661,N_11006,N_10997);
xor U11662 (N_11662,N_10673,N_10992);
xnor U11663 (N_11663,N_10865,N_11048);
xor U11664 (N_11664,N_10993,N_10728);
xnor U11665 (N_11665,N_10707,N_10651);
or U11666 (N_11666,N_10804,N_10694);
or U11667 (N_11667,N_10709,N_10621);
nor U11668 (N_11668,N_11088,N_10856);
xor U11669 (N_11669,N_10925,N_10561);
xnor U11670 (N_11670,N_10452,N_10647);
nor U11671 (N_11671,N_11054,N_10733);
and U11672 (N_11672,N_10693,N_10731);
nor U11673 (N_11673,N_10564,N_10609);
xor U11674 (N_11674,N_10635,N_10476);
and U11675 (N_11675,N_10855,N_11185);
nor U11676 (N_11676,N_10964,N_10528);
nor U11677 (N_11677,N_10498,N_10816);
and U11678 (N_11678,N_10583,N_11001);
or U11679 (N_11679,N_10573,N_10936);
nand U11680 (N_11680,N_10853,N_10767);
and U11681 (N_11681,N_10835,N_10822);
xor U11682 (N_11682,N_10956,N_11113);
or U11683 (N_11683,N_10678,N_11025);
nand U11684 (N_11684,N_10505,N_10927);
nor U11685 (N_11685,N_10590,N_10556);
or U11686 (N_11686,N_11189,N_11188);
nor U11687 (N_11687,N_10829,N_10644);
xnor U11688 (N_11688,N_10544,N_11182);
or U11689 (N_11689,N_10678,N_11092);
or U11690 (N_11690,N_10866,N_10407);
or U11691 (N_11691,N_10981,N_10710);
and U11692 (N_11692,N_10556,N_10445);
and U11693 (N_11693,N_10474,N_10468);
xnor U11694 (N_11694,N_11153,N_10784);
and U11695 (N_11695,N_10743,N_10771);
nand U11696 (N_11696,N_10540,N_11019);
or U11697 (N_11697,N_10912,N_10943);
or U11698 (N_11698,N_10737,N_11158);
nand U11699 (N_11699,N_10823,N_10634);
and U11700 (N_11700,N_11057,N_11042);
nor U11701 (N_11701,N_10593,N_10768);
or U11702 (N_11702,N_10833,N_11137);
or U11703 (N_11703,N_10854,N_10513);
nand U11704 (N_11704,N_10721,N_10832);
or U11705 (N_11705,N_10846,N_10804);
nor U11706 (N_11706,N_11141,N_11143);
xor U11707 (N_11707,N_10887,N_10787);
nor U11708 (N_11708,N_10524,N_10631);
nor U11709 (N_11709,N_10522,N_10745);
xnor U11710 (N_11710,N_10424,N_10710);
and U11711 (N_11711,N_11018,N_10958);
nand U11712 (N_11712,N_10828,N_11055);
and U11713 (N_11713,N_11191,N_10991);
and U11714 (N_11714,N_10578,N_10750);
and U11715 (N_11715,N_10545,N_11049);
nor U11716 (N_11716,N_10449,N_11033);
xnor U11717 (N_11717,N_11044,N_10723);
nand U11718 (N_11718,N_10667,N_10978);
nor U11719 (N_11719,N_10872,N_10928);
nor U11720 (N_11720,N_10544,N_10432);
nand U11721 (N_11721,N_10864,N_10515);
xnor U11722 (N_11722,N_10836,N_11193);
nor U11723 (N_11723,N_10612,N_10877);
and U11724 (N_11724,N_10982,N_10664);
nor U11725 (N_11725,N_10637,N_10870);
nand U11726 (N_11726,N_10933,N_10725);
xnor U11727 (N_11727,N_10859,N_10796);
nor U11728 (N_11728,N_11083,N_11065);
xor U11729 (N_11729,N_10817,N_10469);
and U11730 (N_11730,N_11106,N_11008);
or U11731 (N_11731,N_10516,N_11108);
nand U11732 (N_11732,N_10989,N_10559);
and U11733 (N_11733,N_10630,N_10976);
xnor U11734 (N_11734,N_10425,N_10685);
and U11735 (N_11735,N_10562,N_10689);
xor U11736 (N_11736,N_11047,N_10490);
or U11737 (N_11737,N_10531,N_10576);
and U11738 (N_11738,N_10983,N_11020);
xnor U11739 (N_11739,N_10905,N_10744);
or U11740 (N_11740,N_10592,N_11114);
nand U11741 (N_11741,N_10602,N_10450);
nor U11742 (N_11742,N_10536,N_11148);
and U11743 (N_11743,N_10835,N_11050);
and U11744 (N_11744,N_10954,N_11033);
nor U11745 (N_11745,N_10706,N_11052);
xnor U11746 (N_11746,N_10636,N_10576);
xor U11747 (N_11747,N_10482,N_10977);
and U11748 (N_11748,N_10956,N_10837);
or U11749 (N_11749,N_10765,N_10585);
nor U11750 (N_11750,N_10589,N_10441);
nor U11751 (N_11751,N_10551,N_11057);
nor U11752 (N_11752,N_10670,N_10441);
xnor U11753 (N_11753,N_10689,N_11088);
or U11754 (N_11754,N_10408,N_10959);
nor U11755 (N_11755,N_10878,N_11000);
or U11756 (N_11756,N_10617,N_10986);
nand U11757 (N_11757,N_10509,N_11144);
xor U11758 (N_11758,N_10541,N_10407);
nor U11759 (N_11759,N_10762,N_10445);
nand U11760 (N_11760,N_10795,N_10409);
or U11761 (N_11761,N_10506,N_10512);
and U11762 (N_11762,N_11017,N_10639);
and U11763 (N_11763,N_10517,N_10621);
xnor U11764 (N_11764,N_10985,N_11082);
xnor U11765 (N_11765,N_11002,N_10746);
nand U11766 (N_11766,N_10619,N_10638);
nand U11767 (N_11767,N_10597,N_11182);
nand U11768 (N_11768,N_11069,N_10707);
or U11769 (N_11769,N_10694,N_11197);
or U11770 (N_11770,N_10656,N_10819);
and U11771 (N_11771,N_10689,N_10859);
and U11772 (N_11772,N_10920,N_10935);
xor U11773 (N_11773,N_11120,N_10958);
nor U11774 (N_11774,N_10469,N_10881);
and U11775 (N_11775,N_10868,N_10757);
nand U11776 (N_11776,N_10617,N_11084);
xor U11777 (N_11777,N_11141,N_10590);
nor U11778 (N_11778,N_11174,N_10746);
and U11779 (N_11779,N_10545,N_10747);
nor U11780 (N_11780,N_10832,N_10802);
nor U11781 (N_11781,N_10853,N_10769);
nand U11782 (N_11782,N_11182,N_11039);
or U11783 (N_11783,N_10768,N_10963);
nand U11784 (N_11784,N_11146,N_10546);
nor U11785 (N_11785,N_10830,N_11124);
and U11786 (N_11786,N_10538,N_10711);
nand U11787 (N_11787,N_10861,N_10948);
nand U11788 (N_11788,N_10853,N_10540);
or U11789 (N_11789,N_10510,N_11191);
nand U11790 (N_11790,N_10993,N_10565);
or U11791 (N_11791,N_11152,N_11020);
or U11792 (N_11792,N_11192,N_10510);
nor U11793 (N_11793,N_10719,N_11002);
xnor U11794 (N_11794,N_11032,N_10679);
or U11795 (N_11795,N_11038,N_11139);
or U11796 (N_11796,N_10660,N_10497);
nor U11797 (N_11797,N_11137,N_10515);
and U11798 (N_11798,N_10982,N_11195);
and U11799 (N_11799,N_11145,N_11106);
or U11800 (N_11800,N_10763,N_11160);
nand U11801 (N_11801,N_10531,N_11193);
and U11802 (N_11802,N_11165,N_10506);
xor U11803 (N_11803,N_10923,N_10511);
nand U11804 (N_11804,N_10898,N_11075);
or U11805 (N_11805,N_10614,N_10414);
xor U11806 (N_11806,N_10719,N_11175);
xor U11807 (N_11807,N_10611,N_11193);
nand U11808 (N_11808,N_10544,N_10780);
xor U11809 (N_11809,N_10899,N_10528);
xnor U11810 (N_11810,N_10485,N_10879);
or U11811 (N_11811,N_10620,N_11008);
xnor U11812 (N_11812,N_10852,N_10502);
xor U11813 (N_11813,N_10423,N_11154);
nor U11814 (N_11814,N_10856,N_10496);
and U11815 (N_11815,N_10506,N_11126);
xnor U11816 (N_11816,N_10483,N_10430);
xor U11817 (N_11817,N_10897,N_11192);
nor U11818 (N_11818,N_10985,N_11101);
or U11819 (N_11819,N_10931,N_11141);
or U11820 (N_11820,N_10953,N_10858);
xnor U11821 (N_11821,N_11023,N_10787);
or U11822 (N_11822,N_10833,N_10858);
and U11823 (N_11823,N_10576,N_11013);
xnor U11824 (N_11824,N_11171,N_10538);
nand U11825 (N_11825,N_11173,N_10965);
nor U11826 (N_11826,N_11077,N_10421);
nor U11827 (N_11827,N_11090,N_11073);
and U11828 (N_11828,N_10557,N_11157);
nand U11829 (N_11829,N_10596,N_10445);
nor U11830 (N_11830,N_10691,N_10495);
or U11831 (N_11831,N_10861,N_11050);
nor U11832 (N_11832,N_10551,N_10632);
nor U11833 (N_11833,N_11057,N_10670);
xor U11834 (N_11834,N_10637,N_11001);
or U11835 (N_11835,N_11030,N_10925);
nor U11836 (N_11836,N_11188,N_10550);
or U11837 (N_11837,N_10454,N_10994);
or U11838 (N_11838,N_11044,N_10815);
nand U11839 (N_11839,N_10549,N_10769);
and U11840 (N_11840,N_11105,N_11046);
nor U11841 (N_11841,N_10990,N_10832);
or U11842 (N_11842,N_10415,N_11084);
nor U11843 (N_11843,N_10969,N_11124);
nor U11844 (N_11844,N_11168,N_11135);
or U11845 (N_11845,N_10467,N_10890);
xnor U11846 (N_11846,N_10615,N_10960);
xnor U11847 (N_11847,N_10617,N_10565);
nand U11848 (N_11848,N_10501,N_10986);
or U11849 (N_11849,N_10615,N_10532);
and U11850 (N_11850,N_10614,N_10706);
nor U11851 (N_11851,N_10737,N_11122);
and U11852 (N_11852,N_10958,N_10853);
and U11853 (N_11853,N_10497,N_11147);
nor U11854 (N_11854,N_10796,N_11063);
or U11855 (N_11855,N_10458,N_11192);
nand U11856 (N_11856,N_10699,N_10605);
and U11857 (N_11857,N_10848,N_11002);
xnor U11858 (N_11858,N_11100,N_10773);
nand U11859 (N_11859,N_10759,N_10496);
nor U11860 (N_11860,N_11193,N_10782);
xor U11861 (N_11861,N_10917,N_11123);
nand U11862 (N_11862,N_10495,N_11064);
and U11863 (N_11863,N_10613,N_10900);
or U11864 (N_11864,N_10519,N_10640);
nor U11865 (N_11865,N_10940,N_10893);
or U11866 (N_11866,N_11021,N_10499);
nand U11867 (N_11867,N_10856,N_10576);
xor U11868 (N_11868,N_10677,N_10868);
or U11869 (N_11869,N_10887,N_10685);
nor U11870 (N_11870,N_10547,N_11083);
nor U11871 (N_11871,N_10785,N_10742);
or U11872 (N_11872,N_10859,N_10984);
and U11873 (N_11873,N_10795,N_11143);
nand U11874 (N_11874,N_10557,N_10477);
and U11875 (N_11875,N_10923,N_11181);
or U11876 (N_11876,N_11010,N_11038);
nor U11877 (N_11877,N_10689,N_11127);
xnor U11878 (N_11878,N_10639,N_10559);
nor U11879 (N_11879,N_10936,N_10483);
or U11880 (N_11880,N_10507,N_10800);
xor U11881 (N_11881,N_10599,N_10994);
xor U11882 (N_11882,N_10753,N_10565);
xor U11883 (N_11883,N_10649,N_10618);
xnor U11884 (N_11884,N_10495,N_11127);
xnor U11885 (N_11885,N_11106,N_11018);
xnor U11886 (N_11886,N_10934,N_11121);
and U11887 (N_11887,N_10950,N_11129);
and U11888 (N_11888,N_10693,N_10415);
nand U11889 (N_11889,N_10414,N_10846);
or U11890 (N_11890,N_10526,N_10995);
nor U11891 (N_11891,N_10840,N_11026);
and U11892 (N_11892,N_11182,N_10623);
xor U11893 (N_11893,N_10450,N_10941);
nor U11894 (N_11894,N_10663,N_10777);
or U11895 (N_11895,N_10503,N_11113);
and U11896 (N_11896,N_11031,N_11174);
nor U11897 (N_11897,N_11057,N_10827);
xnor U11898 (N_11898,N_10573,N_10517);
nor U11899 (N_11899,N_11145,N_11179);
nand U11900 (N_11900,N_11004,N_10779);
nand U11901 (N_11901,N_10556,N_11164);
and U11902 (N_11902,N_10453,N_11036);
nor U11903 (N_11903,N_10727,N_11110);
nand U11904 (N_11904,N_11092,N_10541);
or U11905 (N_11905,N_10840,N_10720);
nand U11906 (N_11906,N_10813,N_10606);
xnor U11907 (N_11907,N_10923,N_10878);
or U11908 (N_11908,N_11138,N_10523);
and U11909 (N_11909,N_10934,N_11093);
xor U11910 (N_11910,N_10458,N_10797);
nor U11911 (N_11911,N_10611,N_10657);
xor U11912 (N_11912,N_10491,N_10747);
and U11913 (N_11913,N_10927,N_10572);
nor U11914 (N_11914,N_10666,N_10578);
xor U11915 (N_11915,N_11197,N_10967);
and U11916 (N_11916,N_10615,N_11048);
or U11917 (N_11917,N_10789,N_10808);
nand U11918 (N_11918,N_10572,N_11104);
and U11919 (N_11919,N_10627,N_10890);
nor U11920 (N_11920,N_10453,N_11075);
and U11921 (N_11921,N_10538,N_10503);
and U11922 (N_11922,N_11085,N_10410);
nor U11923 (N_11923,N_10585,N_11046);
xnor U11924 (N_11924,N_10998,N_10600);
nand U11925 (N_11925,N_10718,N_10410);
xnor U11926 (N_11926,N_10775,N_10474);
xor U11927 (N_11927,N_11042,N_10501);
nand U11928 (N_11928,N_10409,N_10411);
and U11929 (N_11929,N_10593,N_10511);
nand U11930 (N_11930,N_11131,N_11192);
and U11931 (N_11931,N_10704,N_10945);
and U11932 (N_11932,N_10977,N_10753);
or U11933 (N_11933,N_10818,N_11028);
and U11934 (N_11934,N_10725,N_10409);
nand U11935 (N_11935,N_10647,N_10922);
xnor U11936 (N_11936,N_11192,N_10856);
and U11937 (N_11937,N_10595,N_10991);
and U11938 (N_11938,N_11026,N_11159);
xor U11939 (N_11939,N_10549,N_10936);
xor U11940 (N_11940,N_10910,N_10736);
xor U11941 (N_11941,N_10468,N_10545);
and U11942 (N_11942,N_10857,N_11025);
or U11943 (N_11943,N_10819,N_11125);
and U11944 (N_11944,N_10733,N_10837);
nor U11945 (N_11945,N_11152,N_11196);
xnor U11946 (N_11946,N_10700,N_11137);
xnor U11947 (N_11947,N_11174,N_10761);
nor U11948 (N_11948,N_10971,N_10908);
nand U11949 (N_11949,N_10466,N_11002);
nand U11950 (N_11950,N_11114,N_10571);
and U11951 (N_11951,N_11015,N_11013);
and U11952 (N_11952,N_11004,N_11007);
nor U11953 (N_11953,N_10718,N_10751);
nor U11954 (N_11954,N_10447,N_10827);
or U11955 (N_11955,N_10721,N_10992);
nor U11956 (N_11956,N_10404,N_10437);
nand U11957 (N_11957,N_11038,N_11106);
and U11958 (N_11958,N_11016,N_10635);
or U11959 (N_11959,N_10538,N_10661);
or U11960 (N_11960,N_10787,N_10971);
nand U11961 (N_11961,N_10564,N_10665);
nor U11962 (N_11962,N_10446,N_11041);
xnor U11963 (N_11963,N_10741,N_10450);
nor U11964 (N_11964,N_11189,N_10527);
and U11965 (N_11965,N_10804,N_10923);
nor U11966 (N_11966,N_10561,N_10415);
and U11967 (N_11967,N_10573,N_10838);
xnor U11968 (N_11968,N_10425,N_10596);
xnor U11969 (N_11969,N_11107,N_10810);
and U11970 (N_11970,N_10736,N_11172);
nor U11971 (N_11971,N_10528,N_10516);
and U11972 (N_11972,N_11083,N_10573);
nand U11973 (N_11973,N_10740,N_10798);
and U11974 (N_11974,N_11134,N_11135);
nand U11975 (N_11975,N_11051,N_10425);
xor U11976 (N_11976,N_10501,N_10598);
or U11977 (N_11977,N_10923,N_10786);
and U11978 (N_11978,N_10957,N_10418);
or U11979 (N_11979,N_10954,N_11137);
and U11980 (N_11980,N_10448,N_10942);
and U11981 (N_11981,N_11130,N_10678);
and U11982 (N_11982,N_10530,N_10623);
xnor U11983 (N_11983,N_10432,N_10616);
and U11984 (N_11984,N_10985,N_10898);
or U11985 (N_11985,N_10817,N_10419);
and U11986 (N_11986,N_10525,N_11192);
or U11987 (N_11987,N_10525,N_10731);
or U11988 (N_11988,N_10917,N_10502);
and U11989 (N_11989,N_10557,N_10847);
or U11990 (N_11990,N_11058,N_10492);
xor U11991 (N_11991,N_10759,N_10462);
nor U11992 (N_11992,N_10833,N_11076);
nor U11993 (N_11993,N_10775,N_10471);
nor U11994 (N_11994,N_11063,N_10714);
xnor U11995 (N_11995,N_10612,N_10561);
xnor U11996 (N_11996,N_10924,N_10492);
or U11997 (N_11997,N_11184,N_10948);
xor U11998 (N_11998,N_10990,N_10474);
xor U11999 (N_11999,N_11077,N_10453);
nor U12000 (N_12000,N_11755,N_11429);
or U12001 (N_12001,N_11686,N_11524);
or U12002 (N_12002,N_11699,N_11359);
and U12003 (N_12003,N_11488,N_11480);
xor U12004 (N_12004,N_11336,N_11862);
nor U12005 (N_12005,N_11647,N_11337);
or U12006 (N_12006,N_11237,N_11926);
xor U12007 (N_12007,N_11865,N_11709);
nor U12008 (N_12008,N_11323,N_11776);
and U12009 (N_12009,N_11410,N_11291);
or U12010 (N_12010,N_11660,N_11405);
and U12011 (N_12011,N_11556,N_11250);
or U12012 (N_12012,N_11316,N_11550);
and U12013 (N_12013,N_11590,N_11475);
or U12014 (N_12014,N_11907,N_11284);
nand U12015 (N_12015,N_11673,N_11226);
nor U12016 (N_12016,N_11665,N_11852);
or U12017 (N_12017,N_11878,N_11585);
and U12018 (N_12018,N_11838,N_11549);
and U12019 (N_12019,N_11917,N_11333);
nor U12020 (N_12020,N_11381,N_11785);
nor U12021 (N_12021,N_11798,N_11496);
and U12022 (N_12022,N_11218,N_11895);
xor U12023 (N_12023,N_11370,N_11840);
or U12024 (N_12024,N_11882,N_11247);
xor U12025 (N_12025,N_11998,N_11986);
and U12026 (N_12026,N_11815,N_11858);
xnor U12027 (N_12027,N_11697,N_11375);
xnor U12028 (N_12028,N_11501,N_11711);
or U12029 (N_12029,N_11844,N_11757);
xnor U12030 (N_12030,N_11619,N_11351);
or U12031 (N_12031,N_11498,N_11352);
nor U12032 (N_12032,N_11887,N_11422);
or U12033 (N_12033,N_11256,N_11520);
nor U12034 (N_12034,N_11789,N_11521);
xnor U12035 (N_12035,N_11955,N_11557);
and U12036 (N_12036,N_11903,N_11720);
and U12037 (N_12037,N_11530,N_11276);
and U12038 (N_12038,N_11257,N_11857);
or U12039 (N_12039,N_11681,N_11603);
and U12040 (N_12040,N_11418,N_11987);
xor U12041 (N_12041,N_11863,N_11769);
xor U12042 (N_12042,N_11575,N_11210);
nor U12043 (N_12043,N_11649,N_11846);
or U12044 (N_12044,N_11918,N_11784);
nor U12045 (N_12045,N_11794,N_11279);
xor U12046 (N_12046,N_11569,N_11202);
nand U12047 (N_12047,N_11956,N_11529);
xor U12048 (N_12048,N_11365,N_11805);
nand U12049 (N_12049,N_11274,N_11743);
nor U12050 (N_12050,N_11388,N_11357);
xnor U12051 (N_12051,N_11842,N_11935);
xnor U12052 (N_12052,N_11450,N_11985);
or U12053 (N_12053,N_11969,N_11380);
or U12054 (N_12054,N_11654,N_11481);
nand U12055 (N_12055,N_11836,N_11730);
nand U12056 (N_12056,N_11508,N_11942);
nand U12057 (N_12057,N_11558,N_11562);
nand U12058 (N_12058,N_11712,N_11742);
nand U12059 (N_12059,N_11566,N_11261);
xnor U12060 (N_12060,N_11988,N_11632);
xor U12061 (N_12061,N_11317,N_11762);
xnor U12062 (N_12062,N_11203,N_11356);
nor U12063 (N_12063,N_11849,N_11432);
nand U12064 (N_12064,N_11579,N_11652);
nand U12065 (N_12065,N_11555,N_11389);
or U12066 (N_12066,N_11680,N_11507);
nand U12067 (N_12067,N_11298,N_11640);
nand U12068 (N_12068,N_11959,N_11212);
nand U12069 (N_12069,N_11727,N_11461);
nand U12070 (N_12070,N_11814,N_11217);
xnor U12071 (N_12071,N_11833,N_11931);
nor U12072 (N_12072,N_11304,N_11492);
xor U12073 (N_12073,N_11994,N_11295);
xnor U12074 (N_12074,N_11435,N_11296);
and U12075 (N_12075,N_11362,N_11916);
nand U12076 (N_12076,N_11589,N_11433);
nor U12077 (N_12077,N_11717,N_11797);
xnor U12078 (N_12078,N_11385,N_11288);
nand U12079 (N_12079,N_11635,N_11592);
nor U12080 (N_12080,N_11414,N_11285);
and U12081 (N_12081,N_11684,N_11674);
xnor U12082 (N_12082,N_11325,N_11253);
nand U12083 (N_12083,N_11650,N_11315);
nor U12084 (N_12084,N_11387,N_11804);
nor U12085 (N_12085,N_11832,N_11458);
or U12086 (N_12086,N_11509,N_11439);
or U12087 (N_12087,N_11354,N_11309);
and U12088 (N_12088,N_11214,N_11493);
or U12089 (N_12089,N_11913,N_11972);
nor U12090 (N_12090,N_11920,N_11885);
or U12091 (N_12091,N_11305,N_11459);
nand U12092 (N_12092,N_11341,N_11453);
nand U12093 (N_12093,N_11930,N_11672);
xnor U12094 (N_12094,N_11324,N_11514);
xor U12095 (N_12095,N_11273,N_11850);
nor U12096 (N_12096,N_11318,N_11749);
nand U12097 (N_12097,N_11997,N_11421);
nand U12098 (N_12098,N_11747,N_11809);
or U12099 (N_12099,N_11424,N_11978);
and U12100 (N_12100,N_11810,N_11818);
or U12101 (N_12101,N_11426,N_11884);
or U12102 (N_12102,N_11209,N_11806);
or U12103 (N_12103,N_11733,N_11983);
xor U12104 (N_12104,N_11233,N_11827);
nor U12105 (N_12105,N_11398,N_11671);
nand U12106 (N_12106,N_11981,N_11466);
or U12107 (N_12107,N_11397,N_11281);
nor U12108 (N_12108,N_11892,N_11937);
nor U12109 (N_12109,N_11262,N_11413);
nand U12110 (N_12110,N_11801,N_11704);
and U12111 (N_12111,N_11741,N_11889);
and U12112 (N_12112,N_11444,N_11420);
and U12113 (N_12113,N_11392,N_11494);
nand U12114 (N_12114,N_11950,N_11343);
nand U12115 (N_12115,N_11779,N_11744);
xnor U12116 (N_12116,N_11263,N_11229);
nor U12117 (N_12117,N_11581,N_11384);
xnor U12118 (N_12118,N_11452,N_11216);
nand U12119 (N_12119,N_11251,N_11477);
and U12120 (N_12120,N_11476,N_11898);
and U12121 (N_12121,N_11310,N_11313);
nor U12122 (N_12122,N_11912,N_11938);
or U12123 (N_12123,N_11900,N_11236);
or U12124 (N_12124,N_11678,N_11770);
nor U12125 (N_12125,N_11732,N_11676);
nand U12126 (N_12126,N_11729,N_11663);
nor U12127 (N_12127,N_11859,N_11694);
nand U12128 (N_12128,N_11446,N_11928);
nand U12129 (N_12129,N_11613,N_11657);
nor U12130 (N_12130,N_11504,N_11948);
or U12131 (N_12131,N_11778,N_11737);
or U12132 (N_12132,N_11624,N_11200);
xnor U12133 (N_12133,N_11462,N_11754);
xnor U12134 (N_12134,N_11947,N_11706);
nand U12135 (N_12135,N_11817,N_11990);
xnor U12136 (N_12136,N_11723,N_11890);
nor U12137 (N_12137,N_11473,N_11860);
nand U12138 (N_12138,N_11811,N_11830);
and U12139 (N_12139,N_11225,N_11244);
and U12140 (N_12140,N_11946,N_11572);
xnor U12141 (N_12141,N_11787,N_11915);
nand U12142 (N_12142,N_11659,N_11607);
and U12143 (N_12143,N_11490,N_11534);
nand U12144 (N_12144,N_11487,N_11311);
and U12145 (N_12145,N_11303,N_11669);
xor U12146 (N_12146,N_11595,N_11535);
or U12147 (N_12147,N_11834,N_11366);
nor U12148 (N_12148,N_11360,N_11580);
nor U12149 (N_12149,N_11621,N_11875);
or U12150 (N_12150,N_11533,N_11993);
nand U12151 (N_12151,N_11588,N_11503);
or U12152 (N_12152,N_11888,N_11220);
and U12153 (N_12153,N_11249,N_11455);
xnor U12154 (N_12154,N_11552,N_11963);
nand U12155 (N_12155,N_11970,N_11338);
or U12156 (N_12156,N_11896,N_11911);
or U12157 (N_12157,N_11252,N_11953);
and U12158 (N_12158,N_11349,N_11841);
or U12159 (N_12159,N_11611,N_11847);
or U12160 (N_12160,N_11996,N_11745);
nor U12161 (N_12161,N_11499,N_11445);
nand U12162 (N_12162,N_11564,N_11416);
xnor U12163 (N_12163,N_11856,N_11377);
or U12164 (N_12164,N_11799,N_11919);
nand U12165 (N_12165,N_11470,N_11540);
nand U12166 (N_12166,N_11670,N_11726);
and U12167 (N_12167,N_11329,N_11867);
nand U12168 (N_12168,N_11696,N_11264);
nor U12169 (N_12169,N_11792,N_11326);
or U12170 (N_12170,N_11642,N_11240);
and U12171 (N_12171,N_11781,N_11599);
nand U12172 (N_12172,N_11399,N_11353);
or U12173 (N_12173,N_11626,N_11725);
and U12174 (N_12174,N_11334,N_11456);
nor U12175 (N_12175,N_11474,N_11837);
nor U12176 (N_12176,N_11656,N_11764);
or U12177 (N_12177,N_11339,N_11417);
nand U12178 (N_12178,N_11457,N_11979);
nor U12179 (N_12179,N_11927,N_11567);
and U12180 (N_12180,N_11714,N_11440);
nor U12181 (N_12181,N_11835,N_11951);
or U12182 (N_12182,N_11363,N_11666);
nand U12183 (N_12183,N_11322,N_11731);
xor U12184 (N_12184,N_11645,N_11831);
xor U12185 (N_12185,N_11633,N_11977);
nand U12186 (N_12186,N_11629,N_11543);
nor U12187 (N_12187,N_11260,N_11547);
nand U12188 (N_12188,N_11637,N_11302);
nor U12189 (N_12189,N_11695,N_11845);
xnor U12190 (N_12190,N_11812,N_11241);
nor U12191 (N_12191,N_11468,N_11902);
nor U12192 (N_12192,N_11280,N_11355);
nand U12193 (N_12193,N_11961,N_11404);
and U12194 (N_12194,N_11265,N_11495);
or U12195 (N_12195,N_11891,N_11735);
or U12196 (N_12196,N_11932,N_11447);
xor U12197 (N_12197,N_11807,N_11331);
nand U12198 (N_12198,N_11861,N_11658);
or U12199 (N_12199,N_11371,N_11301);
xnor U12200 (N_12200,N_11685,N_11692);
or U12201 (N_12201,N_11786,N_11522);
xor U12202 (N_12202,N_11870,N_11545);
or U12203 (N_12203,N_11312,N_11897);
nor U12204 (N_12204,N_11594,N_11344);
xor U12205 (N_12205,N_11448,N_11713);
or U12206 (N_12206,N_11395,N_11945);
and U12207 (N_12207,N_11653,N_11933);
xnor U12208 (N_12208,N_11268,N_11904);
xnor U12209 (N_12209,N_11269,N_11406);
nand U12210 (N_12210,N_11822,N_11428);
or U12211 (N_12211,N_11204,N_11513);
xor U12212 (N_12212,N_11223,N_11544);
nor U12213 (N_12213,N_11565,N_11957);
or U12214 (N_12214,N_11396,N_11971);
nor U12215 (N_12215,N_11716,N_11430);
and U12216 (N_12216,N_11910,N_11431);
and U12217 (N_12217,N_11819,N_11905);
xor U12218 (N_12218,N_11536,N_11705);
nor U12219 (N_12219,N_11293,N_11703);
xor U12220 (N_12220,N_11824,N_11266);
nor U12221 (N_12221,N_11608,N_11372);
nor U12222 (N_12222,N_11515,N_11449);
and U12223 (N_12223,N_11571,N_11497);
or U12224 (N_12224,N_11369,N_11361);
or U12225 (N_12225,N_11472,N_11719);
or U12226 (N_12226,N_11275,N_11708);
nand U12227 (N_12227,N_11609,N_11829);
xnor U12228 (N_12228,N_11267,N_11936);
nand U12229 (N_12229,N_11750,N_11378);
or U12230 (N_12230,N_11623,N_11965);
and U12231 (N_12231,N_11909,N_11828);
and U12232 (N_12232,N_11782,N_11698);
nor U12233 (N_12233,N_11701,N_11615);
xor U12234 (N_12234,N_11612,N_11636);
nand U12235 (N_12235,N_11736,N_11230);
and U12236 (N_12236,N_11738,N_11728);
nor U12237 (N_12237,N_11601,N_11299);
nand U12238 (N_12238,N_11300,N_11700);
nor U12239 (N_12239,N_11485,N_11502);
or U12240 (N_12240,N_11407,N_11872);
and U12241 (N_12241,N_11553,N_11954);
nor U12242 (N_12242,N_11877,N_11206);
and U12243 (N_12243,N_11873,N_11434);
or U12244 (N_12244,N_11638,N_11437);
nor U12245 (N_12245,N_11221,N_11402);
nor U12246 (N_12246,N_11908,N_11843);
or U12247 (N_12247,N_11707,N_11554);
nor U12248 (N_12248,N_11517,N_11574);
xor U12249 (N_12249,N_11880,N_11826);
nand U12250 (N_12250,N_11816,N_11258);
nand U12251 (N_12251,N_11551,N_11901);
xnor U12252 (N_12252,N_11760,N_11943);
or U12253 (N_12253,N_11941,N_11374);
xnor U12254 (N_12254,N_11655,N_11464);
nand U12255 (N_12255,N_11523,N_11587);
and U12256 (N_12256,N_11821,N_11348);
nand U12257 (N_12257,N_11644,N_11604);
or U12258 (N_12258,N_11791,N_11454);
nand U12259 (N_12259,N_11460,N_11242);
or U12260 (N_12260,N_11583,N_11582);
and U12261 (N_12261,N_11332,N_11982);
or U12262 (N_12262,N_11277,N_11876);
nand U12263 (N_12263,N_11677,N_11777);
and U12264 (N_12264,N_11546,N_11478);
and U12265 (N_12265,N_11286,N_11541);
xor U12266 (N_12266,N_11254,N_11899);
or U12267 (N_12267,N_11393,N_11628);
nor U12268 (N_12268,N_11855,N_11335);
nand U12269 (N_12269,N_11425,N_11625);
nand U12270 (N_12270,N_11602,N_11960);
xnor U12271 (N_12271,N_11330,N_11689);
and U12272 (N_12272,N_11412,N_11914);
xor U12273 (N_12273,N_11929,N_11634);
nor U12274 (N_12274,N_11584,N_11319);
and U12275 (N_12275,N_11668,N_11400);
nor U12276 (N_12276,N_11483,N_11561);
and U12277 (N_12277,N_11871,N_11403);
and U12278 (N_12278,N_11968,N_11246);
nor U12279 (N_12279,N_11622,N_11614);
or U12280 (N_12280,N_11314,N_11925);
or U12281 (N_12281,N_11525,N_11759);
xnor U12282 (N_12282,N_11775,N_11245);
or U12283 (N_12283,N_11702,N_11710);
nor U12284 (N_12284,N_11297,N_11238);
nor U12285 (N_12285,N_11577,N_11271);
nor U12286 (N_12286,N_11228,N_11664);
nor U12287 (N_12287,N_11512,N_11854);
and U12288 (N_12288,N_11989,N_11605);
and U12289 (N_12289,N_11222,N_11610);
xnor U12290 (N_12290,N_11272,N_11679);
xnor U12291 (N_12291,N_11576,N_11617);
xor U12292 (N_12292,N_11227,N_11949);
xor U12293 (N_12293,N_11248,N_11208);
nand U12294 (N_12294,N_11894,N_11598);
xor U12295 (N_12295,N_11687,N_11537);
nand U12296 (N_12296,N_11394,N_11788);
nand U12297 (N_12297,N_11347,N_11758);
or U12298 (N_12298,N_11940,N_11408);
xor U12299 (N_12299,N_11772,N_11766);
nand U12300 (N_12300,N_11964,N_11340);
or U12301 (N_12301,N_11869,N_11234);
nand U12302 (N_12302,N_11548,N_11438);
nand U12303 (N_12303,N_11881,N_11526);
or U12304 (N_12304,N_11294,N_11820);
or U12305 (N_12305,N_11999,N_11489);
and U12306 (N_12306,N_11278,N_11469);
or U12307 (N_12307,N_11427,N_11505);
nand U12308 (N_12308,N_11591,N_11382);
nand U12309 (N_12309,N_11688,N_11825);
nand U12310 (N_12310,N_11390,N_11327);
xnor U12311 (N_12311,N_11290,N_11415);
nand U12312 (N_12312,N_11756,N_11853);
nor U12313 (N_12313,N_11739,N_11506);
nor U12314 (N_12314,N_11205,N_11224);
and U12315 (N_12315,N_11207,N_11538);
nor U12316 (N_12316,N_11491,N_11289);
nor U12317 (N_12317,N_11906,N_11597);
xnor U12318 (N_12318,N_11436,N_11851);
and U12319 (N_12319,N_11573,N_11648);
and U12320 (N_12320,N_11967,N_11767);
and U12321 (N_12321,N_11411,N_11639);
nor U12322 (N_12322,N_11682,N_11691);
or U12323 (N_12323,N_11630,N_11886);
nor U12324 (N_12324,N_11646,N_11974);
or U12325 (N_12325,N_11715,N_11401);
and U12326 (N_12326,N_11321,N_11643);
nand U12327 (N_12327,N_11542,N_11724);
and U12328 (N_12328,N_11528,N_11443);
xnor U12329 (N_12329,N_11868,N_11570);
xor U12330 (N_12330,N_11409,N_11320);
xor U12331 (N_12331,N_11235,N_11255);
xnor U12332 (N_12332,N_11751,N_11376);
nor U12333 (N_12333,N_11934,N_11765);
nor U12334 (N_12334,N_11883,N_11368);
and U12335 (N_12335,N_11373,N_11746);
or U12336 (N_12336,N_11306,N_11282);
or U12337 (N_12337,N_11342,N_11471);
nand U12338 (N_12338,N_11966,N_11667);
nand U12339 (N_12339,N_11568,N_11486);
and U12340 (N_12340,N_11923,N_11451);
nor U12341 (N_12341,N_11662,N_11367);
and U12342 (N_12342,N_11419,N_11813);
and U12343 (N_12343,N_11479,N_11532);
and U12344 (N_12344,N_11596,N_11690);
nand U12345 (N_12345,N_11661,N_11991);
nor U12346 (N_12346,N_11586,N_11527);
nor U12347 (N_12347,N_11802,N_11386);
and U12348 (N_12348,N_11627,N_11718);
xnor U12349 (N_12349,N_11467,N_11922);
xor U12350 (N_12350,N_11292,N_11211);
or U12351 (N_12351,N_11391,N_11465);
or U12352 (N_12352,N_11975,N_11539);
xnor U12353 (N_12353,N_11973,N_11952);
nor U12354 (N_12354,N_11559,N_11740);
nand U12355 (N_12355,N_11995,N_11442);
or U12356 (N_12356,N_11463,N_11823);
and U12357 (N_12357,N_11763,N_11924);
xnor U12358 (N_12358,N_11893,N_11771);
and U12359 (N_12359,N_11848,N_11560);
or U12360 (N_12360,N_11962,N_11358);
and U12361 (N_12361,N_11563,N_11976);
and U12362 (N_12362,N_11423,N_11748);
nor U12363 (N_12363,N_11734,N_11783);
xor U12364 (N_12364,N_11683,N_11808);
nor U12365 (N_12365,N_11379,N_11270);
nand U12366 (N_12366,N_11593,N_11364);
and U12367 (N_12367,N_11879,N_11866);
and U12368 (N_12368,N_11243,N_11921);
nand U12369 (N_12369,N_11308,N_11616);
nand U12370 (N_12370,N_11753,N_11796);
xor U12371 (N_12371,N_11752,N_11773);
xor U12372 (N_12372,N_11231,N_11283);
and U12373 (N_12373,N_11693,N_11780);
nor U12374 (N_12374,N_11958,N_11793);
nor U12375 (N_12375,N_11259,N_11984);
or U12376 (N_12376,N_11350,N_11239);
or U12377 (N_12377,N_11232,N_11774);
or U12378 (N_12378,N_11864,N_11219);
nand U12379 (N_12379,N_11531,N_11795);
and U12380 (N_12380,N_11600,N_11620);
and U12381 (N_12381,N_11874,N_11511);
nand U12382 (N_12382,N_11345,N_11939);
xnor U12383 (N_12383,N_11606,N_11516);
or U12384 (N_12384,N_11839,N_11482);
xor U12385 (N_12385,N_11641,N_11675);
and U12386 (N_12386,N_11992,N_11651);
nor U12387 (N_12387,N_11441,N_11618);
nor U12388 (N_12388,N_11518,N_11944);
and U12389 (N_12389,N_11201,N_11307);
nand U12390 (N_12390,N_11980,N_11346);
nor U12391 (N_12391,N_11383,N_11213);
nor U12392 (N_12392,N_11800,N_11287);
nor U12393 (N_12393,N_11761,N_11721);
xor U12394 (N_12394,N_11768,N_11803);
nand U12395 (N_12395,N_11328,N_11510);
nor U12396 (N_12396,N_11519,N_11578);
or U12397 (N_12397,N_11215,N_11484);
nand U12398 (N_12398,N_11790,N_11500);
nand U12399 (N_12399,N_11722,N_11631);
nand U12400 (N_12400,N_11367,N_11769);
and U12401 (N_12401,N_11688,N_11341);
xor U12402 (N_12402,N_11747,N_11834);
and U12403 (N_12403,N_11529,N_11207);
and U12404 (N_12404,N_11795,N_11357);
and U12405 (N_12405,N_11868,N_11590);
nand U12406 (N_12406,N_11663,N_11938);
nand U12407 (N_12407,N_11700,N_11950);
xor U12408 (N_12408,N_11805,N_11459);
nand U12409 (N_12409,N_11871,N_11501);
and U12410 (N_12410,N_11994,N_11902);
nand U12411 (N_12411,N_11911,N_11941);
xor U12412 (N_12412,N_11505,N_11679);
and U12413 (N_12413,N_11568,N_11287);
or U12414 (N_12414,N_11830,N_11280);
nor U12415 (N_12415,N_11545,N_11695);
and U12416 (N_12416,N_11932,N_11854);
or U12417 (N_12417,N_11366,N_11899);
xnor U12418 (N_12418,N_11602,N_11905);
nand U12419 (N_12419,N_11940,N_11392);
nand U12420 (N_12420,N_11936,N_11810);
nor U12421 (N_12421,N_11929,N_11641);
and U12422 (N_12422,N_11562,N_11421);
and U12423 (N_12423,N_11735,N_11647);
nand U12424 (N_12424,N_11524,N_11373);
nor U12425 (N_12425,N_11402,N_11935);
or U12426 (N_12426,N_11276,N_11237);
xnor U12427 (N_12427,N_11286,N_11894);
nand U12428 (N_12428,N_11499,N_11727);
nor U12429 (N_12429,N_11202,N_11755);
and U12430 (N_12430,N_11986,N_11563);
xnor U12431 (N_12431,N_11292,N_11627);
and U12432 (N_12432,N_11747,N_11837);
xnor U12433 (N_12433,N_11858,N_11255);
xnor U12434 (N_12434,N_11239,N_11445);
nor U12435 (N_12435,N_11719,N_11429);
xor U12436 (N_12436,N_11471,N_11940);
xor U12437 (N_12437,N_11466,N_11563);
nor U12438 (N_12438,N_11850,N_11968);
nand U12439 (N_12439,N_11523,N_11900);
and U12440 (N_12440,N_11265,N_11253);
nand U12441 (N_12441,N_11805,N_11531);
nor U12442 (N_12442,N_11603,N_11739);
xor U12443 (N_12443,N_11337,N_11274);
xnor U12444 (N_12444,N_11749,N_11222);
xor U12445 (N_12445,N_11783,N_11321);
nand U12446 (N_12446,N_11245,N_11806);
nand U12447 (N_12447,N_11559,N_11989);
xor U12448 (N_12448,N_11432,N_11746);
nor U12449 (N_12449,N_11784,N_11593);
and U12450 (N_12450,N_11646,N_11626);
or U12451 (N_12451,N_11950,N_11529);
and U12452 (N_12452,N_11709,N_11891);
nand U12453 (N_12453,N_11321,N_11724);
or U12454 (N_12454,N_11435,N_11352);
nand U12455 (N_12455,N_11234,N_11978);
and U12456 (N_12456,N_11524,N_11965);
nand U12457 (N_12457,N_11440,N_11437);
or U12458 (N_12458,N_11578,N_11620);
xor U12459 (N_12459,N_11229,N_11846);
and U12460 (N_12460,N_11248,N_11329);
xnor U12461 (N_12461,N_11712,N_11861);
xor U12462 (N_12462,N_11386,N_11996);
xor U12463 (N_12463,N_11747,N_11278);
nor U12464 (N_12464,N_11924,N_11494);
nor U12465 (N_12465,N_11289,N_11361);
nor U12466 (N_12466,N_11980,N_11467);
and U12467 (N_12467,N_11749,N_11726);
nand U12468 (N_12468,N_11292,N_11338);
and U12469 (N_12469,N_11391,N_11442);
and U12470 (N_12470,N_11927,N_11376);
xnor U12471 (N_12471,N_11786,N_11898);
nand U12472 (N_12472,N_11972,N_11747);
xnor U12473 (N_12473,N_11984,N_11783);
or U12474 (N_12474,N_11534,N_11293);
nor U12475 (N_12475,N_11314,N_11810);
nand U12476 (N_12476,N_11469,N_11852);
nand U12477 (N_12477,N_11941,N_11820);
and U12478 (N_12478,N_11684,N_11937);
xnor U12479 (N_12479,N_11493,N_11957);
nand U12480 (N_12480,N_11535,N_11385);
nor U12481 (N_12481,N_11794,N_11750);
and U12482 (N_12482,N_11772,N_11869);
xor U12483 (N_12483,N_11628,N_11700);
xor U12484 (N_12484,N_11654,N_11883);
nand U12485 (N_12485,N_11337,N_11526);
xor U12486 (N_12486,N_11219,N_11642);
xor U12487 (N_12487,N_11208,N_11316);
xnor U12488 (N_12488,N_11390,N_11644);
nand U12489 (N_12489,N_11403,N_11301);
nor U12490 (N_12490,N_11443,N_11977);
and U12491 (N_12491,N_11711,N_11993);
nand U12492 (N_12492,N_11402,N_11677);
or U12493 (N_12493,N_11472,N_11422);
nand U12494 (N_12494,N_11561,N_11373);
nand U12495 (N_12495,N_11528,N_11734);
nand U12496 (N_12496,N_11461,N_11406);
or U12497 (N_12497,N_11638,N_11428);
nor U12498 (N_12498,N_11586,N_11294);
xor U12499 (N_12499,N_11616,N_11827);
nor U12500 (N_12500,N_11254,N_11724);
nor U12501 (N_12501,N_11506,N_11939);
nand U12502 (N_12502,N_11373,N_11497);
and U12503 (N_12503,N_11813,N_11304);
nor U12504 (N_12504,N_11359,N_11387);
and U12505 (N_12505,N_11396,N_11513);
xor U12506 (N_12506,N_11382,N_11923);
nor U12507 (N_12507,N_11611,N_11430);
nand U12508 (N_12508,N_11547,N_11501);
nand U12509 (N_12509,N_11758,N_11899);
nor U12510 (N_12510,N_11728,N_11566);
nor U12511 (N_12511,N_11823,N_11250);
xnor U12512 (N_12512,N_11635,N_11844);
or U12513 (N_12513,N_11390,N_11920);
nor U12514 (N_12514,N_11460,N_11259);
and U12515 (N_12515,N_11232,N_11389);
nor U12516 (N_12516,N_11500,N_11651);
xnor U12517 (N_12517,N_11508,N_11979);
nand U12518 (N_12518,N_11719,N_11862);
nor U12519 (N_12519,N_11789,N_11219);
or U12520 (N_12520,N_11784,N_11753);
or U12521 (N_12521,N_11582,N_11960);
nor U12522 (N_12522,N_11237,N_11749);
nor U12523 (N_12523,N_11981,N_11816);
or U12524 (N_12524,N_11869,N_11868);
or U12525 (N_12525,N_11606,N_11846);
and U12526 (N_12526,N_11862,N_11945);
and U12527 (N_12527,N_11881,N_11619);
nand U12528 (N_12528,N_11860,N_11833);
nor U12529 (N_12529,N_11526,N_11313);
nand U12530 (N_12530,N_11445,N_11530);
nand U12531 (N_12531,N_11480,N_11584);
or U12532 (N_12532,N_11843,N_11747);
or U12533 (N_12533,N_11211,N_11322);
or U12534 (N_12534,N_11988,N_11469);
xor U12535 (N_12535,N_11715,N_11755);
nand U12536 (N_12536,N_11752,N_11425);
nand U12537 (N_12537,N_11968,N_11648);
nand U12538 (N_12538,N_11976,N_11411);
and U12539 (N_12539,N_11635,N_11214);
nand U12540 (N_12540,N_11450,N_11599);
and U12541 (N_12541,N_11549,N_11733);
xnor U12542 (N_12542,N_11273,N_11528);
and U12543 (N_12543,N_11935,N_11780);
or U12544 (N_12544,N_11888,N_11219);
nor U12545 (N_12545,N_11950,N_11517);
nor U12546 (N_12546,N_11711,N_11788);
or U12547 (N_12547,N_11237,N_11362);
nand U12548 (N_12548,N_11464,N_11885);
or U12549 (N_12549,N_11446,N_11551);
or U12550 (N_12550,N_11678,N_11894);
xnor U12551 (N_12551,N_11325,N_11473);
or U12552 (N_12552,N_11689,N_11899);
xnor U12553 (N_12553,N_11327,N_11457);
nor U12554 (N_12554,N_11915,N_11490);
and U12555 (N_12555,N_11276,N_11550);
xor U12556 (N_12556,N_11932,N_11218);
nand U12557 (N_12557,N_11266,N_11718);
nor U12558 (N_12558,N_11977,N_11288);
or U12559 (N_12559,N_11386,N_11594);
nand U12560 (N_12560,N_11690,N_11767);
nand U12561 (N_12561,N_11544,N_11681);
nand U12562 (N_12562,N_11790,N_11556);
nand U12563 (N_12563,N_11645,N_11249);
or U12564 (N_12564,N_11749,N_11738);
nor U12565 (N_12565,N_11221,N_11225);
nor U12566 (N_12566,N_11261,N_11224);
or U12567 (N_12567,N_11551,N_11706);
nor U12568 (N_12568,N_11687,N_11226);
nand U12569 (N_12569,N_11649,N_11571);
xnor U12570 (N_12570,N_11288,N_11580);
nor U12571 (N_12571,N_11978,N_11437);
or U12572 (N_12572,N_11411,N_11675);
nor U12573 (N_12573,N_11469,N_11449);
nor U12574 (N_12574,N_11741,N_11718);
nand U12575 (N_12575,N_11630,N_11340);
nor U12576 (N_12576,N_11252,N_11206);
xor U12577 (N_12577,N_11782,N_11618);
xnor U12578 (N_12578,N_11799,N_11774);
nor U12579 (N_12579,N_11932,N_11957);
nand U12580 (N_12580,N_11309,N_11472);
xnor U12581 (N_12581,N_11912,N_11906);
xor U12582 (N_12582,N_11478,N_11579);
xnor U12583 (N_12583,N_11227,N_11916);
and U12584 (N_12584,N_11253,N_11223);
nor U12585 (N_12585,N_11552,N_11298);
xnor U12586 (N_12586,N_11311,N_11710);
nor U12587 (N_12587,N_11554,N_11966);
or U12588 (N_12588,N_11598,N_11656);
nand U12589 (N_12589,N_11281,N_11538);
nor U12590 (N_12590,N_11549,N_11604);
xnor U12591 (N_12591,N_11364,N_11713);
and U12592 (N_12592,N_11777,N_11580);
and U12593 (N_12593,N_11274,N_11226);
or U12594 (N_12594,N_11447,N_11323);
and U12595 (N_12595,N_11827,N_11525);
xor U12596 (N_12596,N_11445,N_11247);
or U12597 (N_12597,N_11492,N_11821);
nor U12598 (N_12598,N_11219,N_11316);
nand U12599 (N_12599,N_11774,N_11723);
or U12600 (N_12600,N_11475,N_11378);
nand U12601 (N_12601,N_11553,N_11546);
nand U12602 (N_12602,N_11324,N_11747);
nand U12603 (N_12603,N_11636,N_11313);
nor U12604 (N_12604,N_11698,N_11563);
nor U12605 (N_12605,N_11228,N_11891);
nor U12606 (N_12606,N_11318,N_11505);
xnor U12607 (N_12607,N_11825,N_11568);
xnor U12608 (N_12608,N_11474,N_11253);
xnor U12609 (N_12609,N_11397,N_11517);
and U12610 (N_12610,N_11514,N_11924);
xnor U12611 (N_12611,N_11599,N_11801);
or U12612 (N_12612,N_11430,N_11438);
nand U12613 (N_12613,N_11735,N_11525);
nor U12614 (N_12614,N_11670,N_11840);
nand U12615 (N_12615,N_11543,N_11404);
xor U12616 (N_12616,N_11401,N_11986);
and U12617 (N_12617,N_11981,N_11941);
or U12618 (N_12618,N_11374,N_11459);
or U12619 (N_12619,N_11977,N_11714);
nand U12620 (N_12620,N_11920,N_11875);
nand U12621 (N_12621,N_11522,N_11652);
xnor U12622 (N_12622,N_11250,N_11537);
nand U12623 (N_12623,N_11878,N_11880);
nor U12624 (N_12624,N_11897,N_11286);
and U12625 (N_12625,N_11788,N_11543);
or U12626 (N_12626,N_11724,N_11271);
or U12627 (N_12627,N_11284,N_11934);
nor U12628 (N_12628,N_11531,N_11895);
xnor U12629 (N_12629,N_11401,N_11396);
xnor U12630 (N_12630,N_11892,N_11953);
and U12631 (N_12631,N_11577,N_11290);
and U12632 (N_12632,N_11915,N_11828);
nor U12633 (N_12633,N_11328,N_11336);
nor U12634 (N_12634,N_11771,N_11348);
or U12635 (N_12635,N_11573,N_11778);
or U12636 (N_12636,N_11863,N_11741);
and U12637 (N_12637,N_11468,N_11688);
and U12638 (N_12638,N_11451,N_11853);
nand U12639 (N_12639,N_11359,N_11755);
nand U12640 (N_12640,N_11867,N_11752);
xor U12641 (N_12641,N_11656,N_11756);
or U12642 (N_12642,N_11313,N_11921);
nor U12643 (N_12643,N_11330,N_11576);
and U12644 (N_12644,N_11918,N_11415);
xnor U12645 (N_12645,N_11276,N_11375);
xor U12646 (N_12646,N_11507,N_11437);
nand U12647 (N_12647,N_11692,N_11965);
nor U12648 (N_12648,N_11782,N_11813);
nand U12649 (N_12649,N_11786,N_11511);
and U12650 (N_12650,N_11801,N_11578);
nand U12651 (N_12651,N_11261,N_11812);
or U12652 (N_12652,N_11507,N_11370);
nand U12653 (N_12653,N_11539,N_11597);
nand U12654 (N_12654,N_11836,N_11799);
nor U12655 (N_12655,N_11845,N_11672);
xor U12656 (N_12656,N_11812,N_11275);
xnor U12657 (N_12657,N_11373,N_11221);
nor U12658 (N_12658,N_11685,N_11884);
nor U12659 (N_12659,N_11938,N_11691);
nand U12660 (N_12660,N_11285,N_11640);
nor U12661 (N_12661,N_11319,N_11494);
and U12662 (N_12662,N_11437,N_11892);
and U12663 (N_12663,N_11324,N_11766);
or U12664 (N_12664,N_11456,N_11917);
xor U12665 (N_12665,N_11305,N_11949);
nor U12666 (N_12666,N_11472,N_11942);
nor U12667 (N_12667,N_11740,N_11581);
nand U12668 (N_12668,N_11641,N_11365);
xnor U12669 (N_12669,N_11927,N_11477);
nand U12670 (N_12670,N_11524,N_11995);
or U12671 (N_12671,N_11612,N_11668);
nor U12672 (N_12672,N_11702,N_11859);
nand U12673 (N_12673,N_11769,N_11727);
xnor U12674 (N_12674,N_11553,N_11880);
and U12675 (N_12675,N_11739,N_11717);
nor U12676 (N_12676,N_11756,N_11700);
or U12677 (N_12677,N_11611,N_11859);
and U12678 (N_12678,N_11652,N_11200);
or U12679 (N_12679,N_11777,N_11318);
or U12680 (N_12680,N_11543,N_11497);
or U12681 (N_12681,N_11845,N_11495);
nor U12682 (N_12682,N_11673,N_11668);
or U12683 (N_12683,N_11496,N_11783);
and U12684 (N_12684,N_11719,N_11723);
nand U12685 (N_12685,N_11317,N_11537);
nor U12686 (N_12686,N_11964,N_11700);
or U12687 (N_12687,N_11594,N_11681);
nand U12688 (N_12688,N_11845,N_11978);
and U12689 (N_12689,N_11511,N_11999);
and U12690 (N_12690,N_11877,N_11596);
nand U12691 (N_12691,N_11514,N_11813);
and U12692 (N_12692,N_11991,N_11396);
nand U12693 (N_12693,N_11698,N_11203);
or U12694 (N_12694,N_11651,N_11738);
or U12695 (N_12695,N_11990,N_11308);
nand U12696 (N_12696,N_11545,N_11957);
nand U12697 (N_12697,N_11957,N_11624);
or U12698 (N_12698,N_11330,N_11651);
xnor U12699 (N_12699,N_11816,N_11368);
and U12700 (N_12700,N_11760,N_11733);
nor U12701 (N_12701,N_11217,N_11637);
xor U12702 (N_12702,N_11233,N_11627);
nor U12703 (N_12703,N_11231,N_11870);
or U12704 (N_12704,N_11541,N_11586);
nand U12705 (N_12705,N_11876,N_11846);
nand U12706 (N_12706,N_11721,N_11506);
xor U12707 (N_12707,N_11934,N_11374);
and U12708 (N_12708,N_11737,N_11565);
or U12709 (N_12709,N_11810,N_11717);
or U12710 (N_12710,N_11708,N_11963);
nor U12711 (N_12711,N_11941,N_11694);
or U12712 (N_12712,N_11214,N_11500);
nand U12713 (N_12713,N_11852,N_11736);
and U12714 (N_12714,N_11911,N_11289);
xnor U12715 (N_12715,N_11547,N_11731);
or U12716 (N_12716,N_11663,N_11284);
nor U12717 (N_12717,N_11896,N_11876);
xor U12718 (N_12718,N_11370,N_11333);
or U12719 (N_12719,N_11479,N_11269);
xor U12720 (N_12720,N_11778,N_11902);
and U12721 (N_12721,N_11701,N_11246);
nor U12722 (N_12722,N_11286,N_11989);
nor U12723 (N_12723,N_11453,N_11429);
or U12724 (N_12724,N_11724,N_11272);
xnor U12725 (N_12725,N_11790,N_11363);
nand U12726 (N_12726,N_11867,N_11326);
or U12727 (N_12727,N_11390,N_11798);
xnor U12728 (N_12728,N_11334,N_11478);
nand U12729 (N_12729,N_11751,N_11448);
and U12730 (N_12730,N_11585,N_11756);
xnor U12731 (N_12731,N_11420,N_11974);
xnor U12732 (N_12732,N_11958,N_11504);
nor U12733 (N_12733,N_11230,N_11914);
nand U12734 (N_12734,N_11466,N_11886);
nand U12735 (N_12735,N_11533,N_11945);
xor U12736 (N_12736,N_11853,N_11629);
and U12737 (N_12737,N_11671,N_11890);
or U12738 (N_12738,N_11569,N_11914);
nor U12739 (N_12739,N_11462,N_11612);
or U12740 (N_12740,N_11552,N_11921);
and U12741 (N_12741,N_11783,N_11646);
and U12742 (N_12742,N_11745,N_11909);
or U12743 (N_12743,N_11689,N_11855);
nor U12744 (N_12744,N_11679,N_11504);
or U12745 (N_12745,N_11615,N_11233);
or U12746 (N_12746,N_11736,N_11759);
and U12747 (N_12747,N_11452,N_11260);
and U12748 (N_12748,N_11587,N_11835);
and U12749 (N_12749,N_11656,N_11205);
or U12750 (N_12750,N_11915,N_11933);
or U12751 (N_12751,N_11339,N_11580);
nand U12752 (N_12752,N_11718,N_11844);
nand U12753 (N_12753,N_11623,N_11985);
or U12754 (N_12754,N_11404,N_11202);
nor U12755 (N_12755,N_11298,N_11754);
and U12756 (N_12756,N_11721,N_11484);
nand U12757 (N_12757,N_11785,N_11314);
xor U12758 (N_12758,N_11941,N_11689);
xor U12759 (N_12759,N_11760,N_11804);
and U12760 (N_12760,N_11484,N_11856);
nand U12761 (N_12761,N_11964,N_11215);
and U12762 (N_12762,N_11646,N_11480);
nand U12763 (N_12763,N_11697,N_11411);
and U12764 (N_12764,N_11268,N_11677);
nor U12765 (N_12765,N_11413,N_11583);
and U12766 (N_12766,N_11787,N_11927);
or U12767 (N_12767,N_11321,N_11635);
or U12768 (N_12768,N_11710,N_11804);
nand U12769 (N_12769,N_11973,N_11400);
or U12770 (N_12770,N_11963,N_11960);
nor U12771 (N_12771,N_11487,N_11518);
nand U12772 (N_12772,N_11577,N_11262);
nand U12773 (N_12773,N_11985,N_11890);
nor U12774 (N_12774,N_11485,N_11895);
or U12775 (N_12775,N_11796,N_11881);
and U12776 (N_12776,N_11904,N_11975);
or U12777 (N_12777,N_11291,N_11872);
nor U12778 (N_12778,N_11693,N_11281);
or U12779 (N_12779,N_11963,N_11485);
and U12780 (N_12780,N_11847,N_11976);
or U12781 (N_12781,N_11365,N_11660);
nor U12782 (N_12782,N_11975,N_11206);
or U12783 (N_12783,N_11322,N_11714);
and U12784 (N_12784,N_11908,N_11853);
and U12785 (N_12785,N_11717,N_11461);
nor U12786 (N_12786,N_11614,N_11976);
nor U12787 (N_12787,N_11948,N_11539);
and U12788 (N_12788,N_11874,N_11560);
xor U12789 (N_12789,N_11309,N_11884);
xor U12790 (N_12790,N_11748,N_11856);
xor U12791 (N_12791,N_11398,N_11514);
nor U12792 (N_12792,N_11775,N_11359);
and U12793 (N_12793,N_11257,N_11416);
nand U12794 (N_12794,N_11285,N_11346);
nor U12795 (N_12795,N_11653,N_11526);
nand U12796 (N_12796,N_11335,N_11252);
xor U12797 (N_12797,N_11212,N_11467);
nand U12798 (N_12798,N_11645,N_11789);
and U12799 (N_12799,N_11514,N_11685);
xnor U12800 (N_12800,N_12007,N_12793);
nand U12801 (N_12801,N_12161,N_12723);
and U12802 (N_12802,N_12246,N_12781);
or U12803 (N_12803,N_12686,N_12774);
xnor U12804 (N_12804,N_12778,N_12738);
or U12805 (N_12805,N_12317,N_12622);
nor U12806 (N_12806,N_12526,N_12340);
nor U12807 (N_12807,N_12357,N_12220);
or U12808 (N_12808,N_12422,N_12114);
and U12809 (N_12809,N_12119,N_12534);
nand U12810 (N_12810,N_12025,N_12201);
xor U12811 (N_12811,N_12057,N_12043);
nand U12812 (N_12812,N_12518,N_12280);
nor U12813 (N_12813,N_12584,N_12790);
and U12814 (N_12814,N_12286,N_12027);
and U12815 (N_12815,N_12536,N_12364);
nand U12816 (N_12816,N_12361,N_12580);
nand U12817 (N_12817,N_12308,N_12578);
nor U12818 (N_12818,N_12756,N_12140);
or U12819 (N_12819,N_12180,N_12232);
and U12820 (N_12820,N_12315,N_12552);
and U12821 (N_12821,N_12276,N_12036);
xnor U12822 (N_12822,N_12309,N_12726);
or U12823 (N_12823,N_12077,N_12743);
and U12824 (N_12824,N_12252,N_12108);
xor U12825 (N_12825,N_12639,N_12399);
nor U12826 (N_12826,N_12478,N_12718);
or U12827 (N_12827,N_12395,N_12771);
and U12828 (N_12828,N_12100,N_12166);
or U12829 (N_12829,N_12666,N_12327);
nor U12830 (N_12830,N_12107,N_12389);
xor U12831 (N_12831,N_12721,N_12342);
nor U12832 (N_12832,N_12241,N_12728);
nand U12833 (N_12833,N_12335,N_12099);
xor U12834 (N_12834,N_12768,N_12056);
nor U12835 (N_12835,N_12504,N_12481);
nand U12836 (N_12836,N_12611,N_12654);
nor U12837 (N_12837,N_12397,N_12544);
nor U12838 (N_12838,N_12625,N_12451);
nor U12839 (N_12839,N_12111,N_12700);
nor U12840 (N_12840,N_12442,N_12343);
nand U12841 (N_12841,N_12329,N_12709);
and U12842 (N_12842,N_12613,N_12633);
nor U12843 (N_12843,N_12486,N_12311);
and U12844 (N_12844,N_12330,N_12670);
or U12845 (N_12845,N_12117,N_12755);
nor U12846 (N_12846,N_12758,N_12199);
and U12847 (N_12847,N_12365,N_12334);
nand U12848 (N_12848,N_12591,N_12603);
nand U12849 (N_12849,N_12352,N_12473);
xor U12850 (N_12850,N_12558,N_12258);
nor U12851 (N_12851,N_12541,N_12200);
nor U12852 (N_12852,N_12013,N_12326);
and U12853 (N_12853,N_12254,N_12414);
nand U12854 (N_12854,N_12185,N_12398);
or U12855 (N_12855,N_12453,N_12701);
or U12856 (N_12856,N_12678,N_12441);
nor U12857 (N_12857,N_12616,N_12685);
nor U12858 (N_12858,N_12174,N_12575);
xor U12859 (N_12859,N_12406,N_12532);
nand U12860 (N_12860,N_12773,N_12015);
nand U12861 (N_12861,N_12448,N_12366);
nand U12862 (N_12862,N_12605,N_12052);
or U12863 (N_12863,N_12629,N_12657);
xnor U12864 (N_12864,N_12150,N_12240);
nand U12865 (N_12865,N_12643,N_12417);
nand U12866 (N_12866,N_12371,N_12144);
and U12867 (N_12867,N_12086,N_12542);
nand U12868 (N_12868,N_12784,N_12332);
and U12869 (N_12869,N_12022,N_12164);
or U12870 (N_12870,N_12391,N_12323);
and U12871 (N_12871,N_12158,N_12551);
nand U12872 (N_12872,N_12206,N_12432);
nor U12873 (N_12873,N_12346,N_12594);
or U12874 (N_12874,N_12725,N_12546);
nor U12875 (N_12875,N_12634,N_12145);
or U12876 (N_12876,N_12418,N_12179);
nand U12877 (N_12877,N_12168,N_12024);
nor U12878 (N_12878,N_12628,N_12533);
or U12879 (N_12879,N_12178,N_12294);
nor U12880 (N_12880,N_12059,N_12132);
xnor U12881 (N_12881,N_12296,N_12596);
or U12882 (N_12882,N_12681,N_12410);
xor U12883 (N_12883,N_12644,N_12285);
nor U12884 (N_12884,N_12118,N_12046);
xor U12885 (N_12885,N_12467,N_12475);
nand U12886 (N_12886,N_12452,N_12275);
or U12887 (N_12887,N_12565,N_12302);
or U12888 (N_12888,N_12236,N_12691);
or U12889 (N_12889,N_12073,N_12494);
and U12890 (N_12890,N_12447,N_12588);
and U12891 (N_12891,N_12281,N_12155);
xor U12892 (N_12892,N_12627,N_12676);
or U12893 (N_12893,N_12677,N_12461);
or U12894 (N_12894,N_12379,N_12067);
nor U12895 (N_12895,N_12690,N_12527);
nand U12896 (N_12896,N_12496,N_12493);
and U12897 (N_12897,N_12297,N_12568);
and U12898 (N_12898,N_12328,N_12171);
or U12899 (N_12899,N_12121,N_12135);
and U12900 (N_12900,N_12706,N_12782);
and U12901 (N_12901,N_12122,N_12050);
nand U12902 (N_12902,N_12030,N_12113);
nor U12903 (N_12903,N_12267,N_12641);
nor U12904 (N_12904,N_12188,N_12714);
or U12905 (N_12905,N_12582,N_12636);
nand U12906 (N_12906,N_12766,N_12028);
xor U12907 (N_12907,N_12060,N_12663);
xnor U12908 (N_12908,N_12423,N_12684);
xnor U12909 (N_12909,N_12257,N_12210);
xnor U12910 (N_12910,N_12384,N_12579);
nor U12911 (N_12911,N_12125,N_12176);
or U12912 (N_12912,N_12522,N_12638);
nor U12913 (N_12913,N_12187,N_12416);
nor U12914 (N_12914,N_12383,N_12464);
nor U12915 (N_12915,N_12078,N_12231);
and U12916 (N_12916,N_12499,N_12312);
nor U12917 (N_12917,N_12704,N_12126);
xnor U12918 (N_12918,N_12157,N_12255);
nor U12919 (N_12919,N_12519,N_12169);
nand U12920 (N_12920,N_12228,N_12087);
and U12921 (N_12921,N_12516,N_12513);
xnor U12922 (N_12922,N_12449,N_12539);
xnor U12923 (N_12923,N_12740,N_12211);
and U12924 (N_12924,N_12731,N_12699);
xnor U12925 (N_12925,N_12459,N_12217);
nand U12926 (N_12926,N_12722,N_12746);
nor U12927 (N_12927,N_12295,N_12660);
or U12928 (N_12928,N_12497,N_12523);
or U12929 (N_12929,N_12750,N_12165);
xor U12930 (N_12930,N_12192,N_12095);
nor U12931 (N_12931,N_12387,N_12433);
nor U12932 (N_12932,N_12313,N_12780);
and U12933 (N_12933,N_12152,N_12783);
or U12934 (N_12934,N_12440,N_12624);
or U12935 (N_12935,N_12018,N_12069);
xnor U12936 (N_12936,N_12711,N_12116);
nor U12937 (N_12937,N_12483,N_12474);
and U12938 (N_12938,N_12599,N_12370);
or U12939 (N_12939,N_12378,N_12377);
nor U12940 (N_12940,N_12054,N_12238);
nand U12941 (N_12941,N_12153,N_12703);
nor U12942 (N_12942,N_12687,N_12322);
and U12943 (N_12943,N_12303,N_12618);
or U12944 (N_12944,N_12053,N_12035);
or U12945 (N_12945,N_12096,N_12549);
xnor U12946 (N_12946,N_12712,N_12112);
or U12947 (N_12947,N_12733,N_12615);
xor U12948 (N_12948,N_12430,N_12251);
nand U12949 (N_12949,N_12610,N_12224);
nand U12950 (N_12950,N_12230,N_12256);
or U12951 (N_12951,N_12041,N_12421);
and U12952 (N_12952,N_12457,N_12487);
xor U12953 (N_12953,N_12265,N_12212);
or U12954 (N_12954,N_12472,N_12601);
and U12955 (N_12955,N_12290,N_12612);
nand U12956 (N_12956,N_12614,N_12012);
nor U12957 (N_12957,N_12291,N_12571);
nand U12958 (N_12958,N_12300,N_12261);
nor U12959 (N_12959,N_12567,N_12697);
nor U12960 (N_12960,N_12495,N_12719);
nor U12961 (N_12961,N_12524,N_12319);
or U12962 (N_12962,N_12626,N_12512);
nor U12963 (N_12963,N_12769,N_12734);
and U12964 (N_12964,N_12465,N_12775);
or U12965 (N_12965,N_12262,N_12359);
nor U12966 (N_12966,N_12072,N_12744);
xor U12967 (N_12967,N_12337,N_12581);
and U12968 (N_12968,N_12356,N_12742);
nor U12969 (N_12969,N_12139,N_12530);
xor U12970 (N_12970,N_12392,N_12149);
xnor U12971 (N_12971,N_12156,N_12445);
or U12972 (N_12972,N_12562,N_12786);
or U12973 (N_12973,N_12219,N_12202);
xor U12974 (N_12974,N_12307,N_12632);
nor U12975 (N_12975,N_12031,N_12754);
xor U12976 (N_12976,N_12282,N_12502);
nor U12977 (N_12977,N_12225,N_12160);
or U12978 (N_12978,N_12757,N_12715);
or U12979 (N_12979,N_12271,N_12767);
or U12980 (N_12980,N_12468,N_12403);
xor U12981 (N_12981,N_12266,N_12141);
xor U12982 (N_12982,N_12463,N_12476);
xor U12983 (N_12983,N_12595,N_12234);
nand U12984 (N_12984,N_12431,N_12602);
nand U12985 (N_12985,N_12159,N_12182);
or U12986 (N_12986,N_12514,N_12216);
and U12987 (N_12987,N_12477,N_12653);
nand U12988 (N_12988,N_12189,N_12272);
or U12989 (N_12989,N_12799,N_12029);
and U12990 (N_12990,N_12696,N_12003);
nand U12991 (N_12991,N_12789,N_12314);
and U12992 (N_12992,N_12586,N_12776);
xor U12993 (N_12993,N_12367,N_12511);
and U12994 (N_12994,N_12093,N_12764);
xor U12995 (N_12995,N_12415,N_12298);
nor U12996 (N_12996,N_12630,N_12386);
and U12997 (N_12997,N_12510,N_12795);
nor U12998 (N_12998,N_12058,N_12409);
nor U12999 (N_12999,N_12123,N_12385);
nor U13000 (N_13000,N_12339,N_12484);
nand U13001 (N_13001,N_12535,N_12606);
and U13002 (N_13002,N_12528,N_12344);
and U13003 (N_13003,N_12205,N_12044);
nand U13004 (N_13004,N_12299,N_12124);
nand U13005 (N_13005,N_12426,N_12587);
and U13006 (N_13006,N_12181,N_12573);
nor U13007 (N_13007,N_12640,N_12318);
nor U13008 (N_13008,N_12515,N_12196);
xor U13009 (N_13009,N_12619,N_12263);
nand U13010 (N_13010,N_12623,N_12097);
or U13011 (N_13011,N_12008,N_12537);
nand U13012 (N_13012,N_12553,N_12195);
nand U13013 (N_13013,N_12175,N_12517);
nor U13014 (N_13014,N_12213,N_12001);
or U13015 (N_13015,N_12358,N_12151);
or U13016 (N_13016,N_12023,N_12090);
and U13017 (N_13017,N_12437,N_12045);
xor U13018 (N_13018,N_12508,N_12429);
nand U13019 (N_13019,N_12407,N_12274);
nor U13020 (N_13020,N_12647,N_12239);
or U13021 (N_13021,N_12362,N_12531);
xor U13022 (N_13022,N_12218,N_12233);
or U13023 (N_13023,N_12436,N_12401);
xnor U13024 (N_13024,N_12146,N_12260);
or U13025 (N_13025,N_12664,N_12085);
nor U13026 (N_13026,N_12642,N_12543);
and U13027 (N_13027,N_12191,N_12170);
nor U13028 (N_13028,N_12652,N_12310);
or U13029 (N_13029,N_12082,N_12101);
xor U13030 (N_13030,N_12450,N_12186);
or U13031 (N_13031,N_12503,N_12102);
xnor U13032 (N_13032,N_12702,N_12270);
nor U13033 (N_13033,N_12011,N_12673);
nor U13034 (N_13034,N_12620,N_12055);
nand U13035 (N_13035,N_12197,N_12739);
nor U13036 (N_13036,N_12745,N_12794);
nor U13037 (N_13037,N_12221,N_12621);
and U13038 (N_13038,N_12498,N_12736);
or U13039 (N_13039,N_12569,N_12645);
or U13040 (N_13040,N_12538,N_12278);
xnor U13041 (N_13041,N_12154,N_12689);
nand U13042 (N_13042,N_12444,N_12462);
and U13043 (N_13043,N_12570,N_12109);
xor U13044 (N_13044,N_12075,N_12287);
xor U13045 (N_13045,N_12729,N_12564);
nand U13046 (N_13046,N_12683,N_12301);
or U13047 (N_13047,N_12033,N_12482);
nand U13048 (N_13048,N_12554,N_12411);
and U13049 (N_13049,N_12325,N_12434);
and U13050 (N_13050,N_12720,N_12713);
or U13051 (N_13051,N_12529,N_12223);
or U13052 (N_13052,N_12348,N_12752);
nor U13053 (N_13053,N_12214,N_12002);
or U13054 (N_13054,N_12460,N_12761);
and U13055 (N_13055,N_12556,N_12269);
xor U13056 (N_13056,N_12490,N_12006);
xor U13057 (N_13057,N_12566,N_12479);
nand U13058 (N_13058,N_12129,N_12042);
nor U13059 (N_13059,N_12545,N_12079);
xnor U13060 (N_13060,N_12204,N_12662);
xnor U13061 (N_13061,N_12115,N_12717);
xnor U13062 (N_13062,N_12369,N_12454);
or U13063 (N_13063,N_12374,N_12143);
and U13064 (N_13064,N_12710,N_12229);
or U13065 (N_13065,N_12000,N_12765);
xnor U13066 (N_13066,N_12649,N_12590);
or U13067 (N_13067,N_12198,N_12128);
nor U13068 (N_13068,N_12138,N_12589);
nor U13069 (N_13069,N_12659,N_12705);
xor U13070 (N_13070,N_12279,N_12304);
nor U13071 (N_13071,N_12521,N_12792);
nor U13072 (N_13072,N_12373,N_12724);
nor U13073 (N_13073,N_12388,N_12617);
and U13074 (N_13074,N_12064,N_12561);
or U13075 (N_13075,N_12062,N_12084);
or U13076 (N_13076,N_12405,N_12080);
xnor U13077 (N_13077,N_12797,N_12787);
xnor U13078 (N_13078,N_12026,N_12458);
xnor U13079 (N_13079,N_12604,N_12247);
and U13080 (N_13080,N_12142,N_12785);
nor U13081 (N_13081,N_12390,N_12469);
nand U13082 (N_13082,N_12708,N_12245);
or U13083 (N_13083,N_12751,N_12034);
nor U13084 (N_13084,N_12572,N_12354);
xnor U13085 (N_13085,N_12032,N_12134);
or U13086 (N_13086,N_12264,N_12509);
or U13087 (N_13087,N_12283,N_12491);
or U13088 (N_13088,N_12694,N_12363);
and U13089 (N_13089,N_12016,N_12404);
or U13090 (N_13090,N_12749,N_12021);
and U13091 (N_13091,N_12777,N_12424);
nor U13092 (N_13092,N_12732,N_12268);
nor U13093 (N_13093,N_12242,N_12350);
and U13094 (N_13094,N_12507,N_12669);
and U13095 (N_13095,N_12695,N_12488);
and U13096 (N_13096,N_12540,N_12737);
or U13097 (N_13097,N_12068,N_12550);
xnor U13098 (N_13098,N_12235,N_12184);
nand U13099 (N_13099,N_12438,N_12548);
xnor U13100 (N_13100,N_12376,N_12762);
nand U13101 (N_13101,N_12063,N_12163);
xnor U13102 (N_13102,N_12408,N_12419);
nor U13103 (N_13103,N_12037,N_12355);
nand U13104 (N_13104,N_12083,N_12248);
nand U13105 (N_13105,N_12576,N_12609);
nand U13106 (N_13106,N_12005,N_12485);
and U13107 (N_13107,N_12456,N_12103);
and U13108 (N_13108,N_12402,N_12305);
nand U13109 (N_13109,N_12104,N_12520);
and U13110 (N_13110,N_12547,N_12577);
nor U13111 (N_13111,N_12071,N_12585);
and U13112 (N_13112,N_12646,N_12796);
or U13113 (N_13113,N_12137,N_12049);
nand U13114 (N_13114,N_12250,N_12321);
nor U13115 (N_13115,N_12707,N_12324);
nor U13116 (N_13116,N_12243,N_12368);
nand U13117 (N_13117,N_12592,N_12375);
nand U13118 (N_13118,N_12688,N_12320);
or U13119 (N_13119,N_12074,N_12209);
and U13120 (N_13120,N_12147,N_12167);
xnor U13121 (N_13121,N_12004,N_12009);
xor U13122 (N_13122,N_12593,N_12396);
or U13123 (N_13123,N_12631,N_12244);
nand U13124 (N_13124,N_12655,N_12088);
or U13125 (N_13125,N_12259,N_12446);
nor U13126 (N_13126,N_12637,N_12559);
nand U13127 (N_13127,N_12607,N_12425);
nor U13128 (N_13128,N_12665,N_12583);
nand U13129 (N_13129,N_12671,N_12289);
nand U13130 (N_13130,N_12455,N_12770);
nor U13131 (N_13131,N_12470,N_12020);
nand U13132 (N_13132,N_12336,N_12306);
xnor U13133 (N_13133,N_12316,N_12039);
xor U13134 (N_13134,N_12380,N_12098);
or U13135 (N_13135,N_12381,N_12560);
and U13136 (N_13136,N_12693,N_12148);
nor U13137 (N_13137,N_12131,N_12372);
nor U13138 (N_13138,N_12500,N_12798);
xor U13139 (N_13139,N_12439,N_12393);
and U13140 (N_13140,N_12412,N_12735);
and U13141 (N_13141,N_12203,N_12555);
xor U13142 (N_13142,N_12038,N_12760);
xor U13143 (N_13143,N_12341,N_12651);
or U13144 (N_13144,N_12215,N_12730);
xnor U13145 (N_13145,N_12656,N_12753);
or U13146 (N_13146,N_12748,N_12505);
xnor U13147 (N_13147,N_12208,N_12333);
or U13148 (N_13148,N_12351,N_12227);
or U13149 (N_13149,N_12061,N_12574);
nand U13150 (N_13150,N_12207,N_12065);
and U13151 (N_13151,N_12506,N_12763);
and U13152 (N_13152,N_12635,N_12608);
or U13153 (N_13153,N_12727,N_12597);
xor U13154 (N_13154,N_12253,N_12716);
or U13155 (N_13155,N_12661,N_12658);
or U13156 (N_13156,N_12136,N_12428);
nor U13157 (N_13157,N_12648,N_12759);
nand U13158 (N_13158,N_12047,N_12489);
nor U13159 (N_13159,N_12127,N_12183);
xnor U13160 (N_13160,N_12177,N_12741);
nor U13161 (N_13161,N_12173,N_12193);
and U13162 (N_13162,N_12674,N_12435);
xnor U13163 (N_13163,N_12443,N_12471);
and U13164 (N_13164,N_12172,N_12277);
nor U13165 (N_13165,N_12682,N_12293);
and U13166 (N_13166,N_12747,N_12480);
nor U13167 (N_13167,N_12598,N_12672);
nand U13168 (N_13168,N_12076,N_12772);
or U13169 (N_13169,N_12133,N_12345);
nand U13170 (N_13170,N_12162,N_12563);
xnor U13171 (N_13171,N_12349,N_12360);
nand U13172 (N_13172,N_12675,N_12413);
xor U13173 (N_13173,N_12237,N_12222);
nor U13174 (N_13174,N_12273,N_12557);
nand U13175 (N_13175,N_12650,N_12019);
or U13176 (N_13176,N_12110,N_12492);
and U13177 (N_13177,N_12089,N_12014);
or U13178 (N_13178,N_12466,N_12680);
nand U13179 (N_13179,N_12070,N_12249);
or U13180 (N_13180,N_12788,N_12382);
or U13181 (N_13181,N_12400,N_12600);
or U13182 (N_13182,N_12668,N_12092);
nand U13183 (N_13183,N_12010,N_12347);
xor U13184 (N_13184,N_12698,N_12190);
nor U13185 (N_13185,N_12120,N_12394);
nor U13186 (N_13186,N_12791,N_12066);
nand U13187 (N_13187,N_12194,N_12288);
nor U13188 (N_13188,N_12105,N_12284);
and U13189 (N_13189,N_12226,N_12292);
and U13190 (N_13190,N_12692,N_12081);
nor U13191 (N_13191,N_12106,N_12331);
nor U13192 (N_13192,N_12051,N_12091);
nor U13193 (N_13193,N_12017,N_12427);
nor U13194 (N_13194,N_12130,N_12420);
nor U13195 (N_13195,N_12679,N_12353);
or U13196 (N_13196,N_12779,N_12501);
nand U13197 (N_13197,N_12667,N_12525);
nand U13198 (N_13198,N_12040,N_12048);
nand U13199 (N_13199,N_12338,N_12094);
xor U13200 (N_13200,N_12072,N_12594);
nand U13201 (N_13201,N_12326,N_12587);
nor U13202 (N_13202,N_12165,N_12722);
nor U13203 (N_13203,N_12103,N_12439);
nor U13204 (N_13204,N_12613,N_12212);
and U13205 (N_13205,N_12100,N_12793);
or U13206 (N_13206,N_12511,N_12461);
or U13207 (N_13207,N_12638,N_12511);
nor U13208 (N_13208,N_12054,N_12100);
or U13209 (N_13209,N_12402,N_12048);
xnor U13210 (N_13210,N_12111,N_12266);
or U13211 (N_13211,N_12153,N_12275);
nand U13212 (N_13212,N_12075,N_12730);
nor U13213 (N_13213,N_12640,N_12726);
nand U13214 (N_13214,N_12189,N_12696);
nand U13215 (N_13215,N_12653,N_12382);
nor U13216 (N_13216,N_12352,N_12243);
and U13217 (N_13217,N_12376,N_12041);
and U13218 (N_13218,N_12125,N_12373);
and U13219 (N_13219,N_12273,N_12151);
or U13220 (N_13220,N_12380,N_12736);
nor U13221 (N_13221,N_12063,N_12548);
or U13222 (N_13222,N_12247,N_12115);
nand U13223 (N_13223,N_12351,N_12406);
nand U13224 (N_13224,N_12538,N_12614);
xor U13225 (N_13225,N_12130,N_12138);
and U13226 (N_13226,N_12748,N_12705);
xnor U13227 (N_13227,N_12696,N_12111);
nor U13228 (N_13228,N_12629,N_12143);
and U13229 (N_13229,N_12542,N_12188);
nor U13230 (N_13230,N_12710,N_12547);
xor U13231 (N_13231,N_12580,N_12053);
nand U13232 (N_13232,N_12097,N_12114);
or U13233 (N_13233,N_12300,N_12591);
and U13234 (N_13234,N_12521,N_12171);
or U13235 (N_13235,N_12248,N_12489);
or U13236 (N_13236,N_12203,N_12617);
nor U13237 (N_13237,N_12086,N_12346);
and U13238 (N_13238,N_12152,N_12196);
or U13239 (N_13239,N_12752,N_12777);
nand U13240 (N_13240,N_12433,N_12538);
nor U13241 (N_13241,N_12000,N_12609);
or U13242 (N_13242,N_12276,N_12100);
nand U13243 (N_13243,N_12435,N_12326);
and U13244 (N_13244,N_12681,N_12066);
xor U13245 (N_13245,N_12730,N_12226);
nor U13246 (N_13246,N_12599,N_12784);
nand U13247 (N_13247,N_12204,N_12537);
nor U13248 (N_13248,N_12271,N_12096);
nand U13249 (N_13249,N_12254,N_12496);
xor U13250 (N_13250,N_12349,N_12249);
xor U13251 (N_13251,N_12212,N_12734);
nand U13252 (N_13252,N_12376,N_12000);
nor U13253 (N_13253,N_12139,N_12268);
or U13254 (N_13254,N_12587,N_12640);
nand U13255 (N_13255,N_12370,N_12411);
and U13256 (N_13256,N_12730,N_12529);
or U13257 (N_13257,N_12121,N_12471);
or U13258 (N_13258,N_12438,N_12484);
xnor U13259 (N_13259,N_12625,N_12387);
nand U13260 (N_13260,N_12526,N_12666);
xor U13261 (N_13261,N_12619,N_12515);
and U13262 (N_13262,N_12277,N_12147);
xor U13263 (N_13263,N_12584,N_12032);
nand U13264 (N_13264,N_12706,N_12730);
xnor U13265 (N_13265,N_12056,N_12253);
xnor U13266 (N_13266,N_12622,N_12247);
or U13267 (N_13267,N_12557,N_12160);
nor U13268 (N_13268,N_12526,N_12252);
or U13269 (N_13269,N_12121,N_12033);
nand U13270 (N_13270,N_12290,N_12261);
nor U13271 (N_13271,N_12396,N_12420);
nor U13272 (N_13272,N_12011,N_12705);
or U13273 (N_13273,N_12374,N_12556);
xnor U13274 (N_13274,N_12051,N_12538);
nor U13275 (N_13275,N_12400,N_12301);
nand U13276 (N_13276,N_12453,N_12116);
xnor U13277 (N_13277,N_12371,N_12573);
xnor U13278 (N_13278,N_12204,N_12095);
nand U13279 (N_13279,N_12513,N_12022);
nand U13280 (N_13280,N_12025,N_12318);
nor U13281 (N_13281,N_12064,N_12321);
or U13282 (N_13282,N_12254,N_12200);
nand U13283 (N_13283,N_12729,N_12459);
nand U13284 (N_13284,N_12677,N_12507);
xor U13285 (N_13285,N_12680,N_12147);
xor U13286 (N_13286,N_12255,N_12623);
xor U13287 (N_13287,N_12151,N_12457);
nor U13288 (N_13288,N_12708,N_12482);
nor U13289 (N_13289,N_12386,N_12352);
and U13290 (N_13290,N_12406,N_12021);
nand U13291 (N_13291,N_12615,N_12793);
nor U13292 (N_13292,N_12485,N_12749);
nand U13293 (N_13293,N_12675,N_12300);
xnor U13294 (N_13294,N_12054,N_12184);
nand U13295 (N_13295,N_12512,N_12256);
nand U13296 (N_13296,N_12678,N_12030);
xor U13297 (N_13297,N_12469,N_12088);
xnor U13298 (N_13298,N_12370,N_12068);
or U13299 (N_13299,N_12649,N_12418);
or U13300 (N_13300,N_12209,N_12028);
or U13301 (N_13301,N_12174,N_12166);
or U13302 (N_13302,N_12367,N_12153);
xnor U13303 (N_13303,N_12210,N_12477);
or U13304 (N_13304,N_12636,N_12409);
and U13305 (N_13305,N_12237,N_12291);
nand U13306 (N_13306,N_12293,N_12186);
nor U13307 (N_13307,N_12163,N_12628);
or U13308 (N_13308,N_12739,N_12760);
nand U13309 (N_13309,N_12113,N_12099);
or U13310 (N_13310,N_12744,N_12708);
nor U13311 (N_13311,N_12639,N_12401);
or U13312 (N_13312,N_12107,N_12355);
nand U13313 (N_13313,N_12387,N_12039);
xnor U13314 (N_13314,N_12742,N_12340);
or U13315 (N_13315,N_12687,N_12796);
nand U13316 (N_13316,N_12425,N_12375);
or U13317 (N_13317,N_12073,N_12040);
xnor U13318 (N_13318,N_12432,N_12450);
nor U13319 (N_13319,N_12049,N_12342);
xor U13320 (N_13320,N_12414,N_12228);
nor U13321 (N_13321,N_12620,N_12011);
nor U13322 (N_13322,N_12465,N_12453);
and U13323 (N_13323,N_12208,N_12293);
or U13324 (N_13324,N_12105,N_12670);
nand U13325 (N_13325,N_12057,N_12222);
and U13326 (N_13326,N_12370,N_12639);
and U13327 (N_13327,N_12582,N_12396);
nand U13328 (N_13328,N_12751,N_12266);
and U13329 (N_13329,N_12752,N_12764);
xnor U13330 (N_13330,N_12260,N_12346);
and U13331 (N_13331,N_12438,N_12255);
and U13332 (N_13332,N_12594,N_12577);
nand U13333 (N_13333,N_12072,N_12313);
xor U13334 (N_13334,N_12409,N_12322);
xor U13335 (N_13335,N_12297,N_12368);
or U13336 (N_13336,N_12444,N_12646);
nand U13337 (N_13337,N_12732,N_12134);
xnor U13338 (N_13338,N_12336,N_12760);
nor U13339 (N_13339,N_12033,N_12431);
nand U13340 (N_13340,N_12081,N_12614);
xor U13341 (N_13341,N_12309,N_12459);
nor U13342 (N_13342,N_12514,N_12542);
or U13343 (N_13343,N_12735,N_12675);
nor U13344 (N_13344,N_12097,N_12474);
nor U13345 (N_13345,N_12732,N_12149);
nor U13346 (N_13346,N_12683,N_12606);
xnor U13347 (N_13347,N_12215,N_12672);
xnor U13348 (N_13348,N_12375,N_12495);
and U13349 (N_13349,N_12738,N_12693);
nand U13350 (N_13350,N_12714,N_12383);
xor U13351 (N_13351,N_12239,N_12250);
or U13352 (N_13352,N_12691,N_12208);
or U13353 (N_13353,N_12229,N_12433);
xor U13354 (N_13354,N_12459,N_12192);
and U13355 (N_13355,N_12751,N_12053);
nand U13356 (N_13356,N_12656,N_12035);
nand U13357 (N_13357,N_12140,N_12546);
nor U13358 (N_13358,N_12626,N_12582);
and U13359 (N_13359,N_12619,N_12722);
nand U13360 (N_13360,N_12472,N_12247);
and U13361 (N_13361,N_12571,N_12583);
xnor U13362 (N_13362,N_12608,N_12300);
nand U13363 (N_13363,N_12782,N_12686);
nor U13364 (N_13364,N_12180,N_12348);
and U13365 (N_13365,N_12027,N_12390);
nand U13366 (N_13366,N_12674,N_12789);
or U13367 (N_13367,N_12076,N_12470);
nand U13368 (N_13368,N_12251,N_12214);
nor U13369 (N_13369,N_12457,N_12299);
and U13370 (N_13370,N_12052,N_12492);
nor U13371 (N_13371,N_12744,N_12673);
nor U13372 (N_13372,N_12181,N_12589);
nand U13373 (N_13373,N_12331,N_12239);
xnor U13374 (N_13374,N_12634,N_12096);
nor U13375 (N_13375,N_12562,N_12547);
nand U13376 (N_13376,N_12631,N_12681);
or U13377 (N_13377,N_12754,N_12712);
or U13378 (N_13378,N_12398,N_12628);
nand U13379 (N_13379,N_12723,N_12308);
xnor U13380 (N_13380,N_12658,N_12531);
or U13381 (N_13381,N_12527,N_12022);
xor U13382 (N_13382,N_12264,N_12222);
nor U13383 (N_13383,N_12481,N_12784);
nor U13384 (N_13384,N_12713,N_12376);
and U13385 (N_13385,N_12349,N_12493);
xor U13386 (N_13386,N_12360,N_12733);
or U13387 (N_13387,N_12154,N_12501);
nor U13388 (N_13388,N_12194,N_12149);
nand U13389 (N_13389,N_12425,N_12514);
xnor U13390 (N_13390,N_12205,N_12325);
nand U13391 (N_13391,N_12425,N_12216);
and U13392 (N_13392,N_12191,N_12339);
nand U13393 (N_13393,N_12002,N_12794);
xnor U13394 (N_13394,N_12162,N_12000);
and U13395 (N_13395,N_12767,N_12182);
or U13396 (N_13396,N_12140,N_12182);
nor U13397 (N_13397,N_12042,N_12429);
or U13398 (N_13398,N_12475,N_12403);
nor U13399 (N_13399,N_12545,N_12051);
nand U13400 (N_13400,N_12553,N_12134);
or U13401 (N_13401,N_12565,N_12556);
and U13402 (N_13402,N_12328,N_12288);
nor U13403 (N_13403,N_12568,N_12592);
xnor U13404 (N_13404,N_12428,N_12157);
or U13405 (N_13405,N_12055,N_12315);
or U13406 (N_13406,N_12737,N_12132);
or U13407 (N_13407,N_12367,N_12378);
nand U13408 (N_13408,N_12567,N_12259);
nand U13409 (N_13409,N_12192,N_12359);
nand U13410 (N_13410,N_12786,N_12081);
or U13411 (N_13411,N_12167,N_12354);
xnor U13412 (N_13412,N_12548,N_12775);
or U13413 (N_13413,N_12279,N_12442);
or U13414 (N_13414,N_12522,N_12382);
or U13415 (N_13415,N_12044,N_12686);
and U13416 (N_13416,N_12664,N_12046);
nand U13417 (N_13417,N_12677,N_12621);
and U13418 (N_13418,N_12006,N_12154);
nor U13419 (N_13419,N_12706,N_12585);
xnor U13420 (N_13420,N_12423,N_12695);
and U13421 (N_13421,N_12716,N_12307);
and U13422 (N_13422,N_12357,N_12482);
xnor U13423 (N_13423,N_12136,N_12184);
nand U13424 (N_13424,N_12046,N_12100);
xor U13425 (N_13425,N_12549,N_12700);
nor U13426 (N_13426,N_12605,N_12748);
or U13427 (N_13427,N_12180,N_12322);
or U13428 (N_13428,N_12188,N_12350);
nor U13429 (N_13429,N_12499,N_12149);
or U13430 (N_13430,N_12012,N_12559);
and U13431 (N_13431,N_12662,N_12592);
and U13432 (N_13432,N_12331,N_12045);
nor U13433 (N_13433,N_12399,N_12373);
nor U13434 (N_13434,N_12768,N_12600);
or U13435 (N_13435,N_12493,N_12578);
nor U13436 (N_13436,N_12454,N_12401);
nand U13437 (N_13437,N_12684,N_12084);
nor U13438 (N_13438,N_12124,N_12644);
nand U13439 (N_13439,N_12299,N_12718);
xor U13440 (N_13440,N_12065,N_12708);
nor U13441 (N_13441,N_12340,N_12792);
or U13442 (N_13442,N_12143,N_12265);
or U13443 (N_13443,N_12233,N_12255);
or U13444 (N_13444,N_12091,N_12062);
or U13445 (N_13445,N_12342,N_12663);
or U13446 (N_13446,N_12761,N_12241);
or U13447 (N_13447,N_12618,N_12527);
nor U13448 (N_13448,N_12720,N_12279);
xor U13449 (N_13449,N_12093,N_12102);
or U13450 (N_13450,N_12403,N_12777);
nand U13451 (N_13451,N_12791,N_12309);
nor U13452 (N_13452,N_12309,N_12201);
xnor U13453 (N_13453,N_12501,N_12054);
and U13454 (N_13454,N_12048,N_12292);
nor U13455 (N_13455,N_12358,N_12226);
and U13456 (N_13456,N_12752,N_12301);
and U13457 (N_13457,N_12344,N_12040);
nor U13458 (N_13458,N_12393,N_12073);
or U13459 (N_13459,N_12379,N_12706);
or U13460 (N_13460,N_12386,N_12721);
nor U13461 (N_13461,N_12138,N_12472);
xnor U13462 (N_13462,N_12214,N_12366);
and U13463 (N_13463,N_12717,N_12267);
nor U13464 (N_13464,N_12102,N_12220);
and U13465 (N_13465,N_12408,N_12566);
nor U13466 (N_13466,N_12189,N_12371);
nor U13467 (N_13467,N_12214,N_12151);
and U13468 (N_13468,N_12657,N_12415);
and U13469 (N_13469,N_12600,N_12166);
nand U13470 (N_13470,N_12693,N_12017);
nor U13471 (N_13471,N_12534,N_12573);
nand U13472 (N_13472,N_12178,N_12787);
xnor U13473 (N_13473,N_12062,N_12584);
or U13474 (N_13474,N_12313,N_12707);
nand U13475 (N_13475,N_12654,N_12233);
nor U13476 (N_13476,N_12296,N_12648);
and U13477 (N_13477,N_12676,N_12052);
and U13478 (N_13478,N_12673,N_12540);
xnor U13479 (N_13479,N_12162,N_12027);
nor U13480 (N_13480,N_12370,N_12469);
nor U13481 (N_13481,N_12402,N_12140);
xnor U13482 (N_13482,N_12612,N_12449);
nor U13483 (N_13483,N_12364,N_12410);
nand U13484 (N_13484,N_12375,N_12075);
xor U13485 (N_13485,N_12793,N_12278);
and U13486 (N_13486,N_12691,N_12263);
nand U13487 (N_13487,N_12122,N_12448);
nand U13488 (N_13488,N_12299,N_12745);
or U13489 (N_13489,N_12108,N_12525);
nand U13490 (N_13490,N_12443,N_12314);
xnor U13491 (N_13491,N_12311,N_12424);
xor U13492 (N_13492,N_12559,N_12292);
and U13493 (N_13493,N_12573,N_12179);
and U13494 (N_13494,N_12608,N_12089);
and U13495 (N_13495,N_12150,N_12483);
xor U13496 (N_13496,N_12796,N_12008);
or U13497 (N_13497,N_12263,N_12286);
or U13498 (N_13498,N_12239,N_12078);
xor U13499 (N_13499,N_12043,N_12512);
xor U13500 (N_13500,N_12317,N_12613);
nor U13501 (N_13501,N_12065,N_12312);
nand U13502 (N_13502,N_12633,N_12328);
and U13503 (N_13503,N_12209,N_12175);
nor U13504 (N_13504,N_12618,N_12519);
and U13505 (N_13505,N_12290,N_12384);
nand U13506 (N_13506,N_12209,N_12013);
or U13507 (N_13507,N_12112,N_12342);
nor U13508 (N_13508,N_12658,N_12107);
nor U13509 (N_13509,N_12172,N_12777);
nand U13510 (N_13510,N_12340,N_12021);
xnor U13511 (N_13511,N_12301,N_12486);
xnor U13512 (N_13512,N_12228,N_12259);
nor U13513 (N_13513,N_12473,N_12271);
xnor U13514 (N_13514,N_12638,N_12309);
and U13515 (N_13515,N_12674,N_12677);
xnor U13516 (N_13516,N_12688,N_12440);
and U13517 (N_13517,N_12389,N_12091);
nor U13518 (N_13518,N_12771,N_12043);
or U13519 (N_13519,N_12675,N_12084);
or U13520 (N_13520,N_12677,N_12350);
nand U13521 (N_13521,N_12545,N_12527);
or U13522 (N_13522,N_12620,N_12180);
nand U13523 (N_13523,N_12554,N_12348);
nand U13524 (N_13524,N_12324,N_12028);
xor U13525 (N_13525,N_12022,N_12064);
nor U13526 (N_13526,N_12118,N_12438);
nand U13527 (N_13527,N_12093,N_12006);
and U13528 (N_13528,N_12621,N_12719);
or U13529 (N_13529,N_12427,N_12381);
nor U13530 (N_13530,N_12381,N_12634);
and U13531 (N_13531,N_12667,N_12132);
or U13532 (N_13532,N_12653,N_12396);
nand U13533 (N_13533,N_12084,N_12239);
nor U13534 (N_13534,N_12259,N_12335);
or U13535 (N_13535,N_12444,N_12736);
and U13536 (N_13536,N_12417,N_12572);
nand U13537 (N_13537,N_12492,N_12422);
nand U13538 (N_13538,N_12434,N_12084);
and U13539 (N_13539,N_12557,N_12118);
nor U13540 (N_13540,N_12737,N_12563);
xor U13541 (N_13541,N_12613,N_12298);
nor U13542 (N_13542,N_12611,N_12523);
nor U13543 (N_13543,N_12321,N_12790);
and U13544 (N_13544,N_12360,N_12378);
nor U13545 (N_13545,N_12496,N_12319);
nor U13546 (N_13546,N_12785,N_12686);
or U13547 (N_13547,N_12170,N_12697);
and U13548 (N_13548,N_12305,N_12507);
or U13549 (N_13549,N_12599,N_12039);
or U13550 (N_13550,N_12044,N_12777);
and U13551 (N_13551,N_12141,N_12676);
or U13552 (N_13552,N_12479,N_12179);
or U13553 (N_13553,N_12663,N_12744);
and U13554 (N_13554,N_12305,N_12152);
and U13555 (N_13555,N_12555,N_12626);
and U13556 (N_13556,N_12312,N_12645);
nor U13557 (N_13557,N_12717,N_12357);
nand U13558 (N_13558,N_12722,N_12549);
and U13559 (N_13559,N_12417,N_12200);
nand U13560 (N_13560,N_12160,N_12427);
nor U13561 (N_13561,N_12578,N_12366);
nor U13562 (N_13562,N_12747,N_12075);
xnor U13563 (N_13563,N_12539,N_12301);
nand U13564 (N_13564,N_12250,N_12287);
and U13565 (N_13565,N_12179,N_12439);
nand U13566 (N_13566,N_12145,N_12671);
nor U13567 (N_13567,N_12167,N_12268);
nor U13568 (N_13568,N_12798,N_12068);
nor U13569 (N_13569,N_12047,N_12722);
and U13570 (N_13570,N_12753,N_12150);
xnor U13571 (N_13571,N_12011,N_12665);
or U13572 (N_13572,N_12562,N_12357);
nor U13573 (N_13573,N_12509,N_12205);
or U13574 (N_13574,N_12700,N_12616);
nand U13575 (N_13575,N_12666,N_12237);
xor U13576 (N_13576,N_12249,N_12293);
xnor U13577 (N_13577,N_12756,N_12350);
nor U13578 (N_13578,N_12523,N_12358);
or U13579 (N_13579,N_12395,N_12613);
xnor U13580 (N_13580,N_12615,N_12745);
xnor U13581 (N_13581,N_12344,N_12127);
or U13582 (N_13582,N_12608,N_12525);
nand U13583 (N_13583,N_12134,N_12091);
or U13584 (N_13584,N_12766,N_12691);
xor U13585 (N_13585,N_12231,N_12531);
xnor U13586 (N_13586,N_12688,N_12752);
nor U13587 (N_13587,N_12535,N_12405);
and U13588 (N_13588,N_12676,N_12704);
nand U13589 (N_13589,N_12189,N_12751);
and U13590 (N_13590,N_12723,N_12007);
or U13591 (N_13591,N_12450,N_12537);
nor U13592 (N_13592,N_12439,N_12526);
nand U13593 (N_13593,N_12793,N_12624);
xor U13594 (N_13594,N_12188,N_12324);
nand U13595 (N_13595,N_12239,N_12560);
or U13596 (N_13596,N_12018,N_12353);
and U13597 (N_13597,N_12454,N_12783);
or U13598 (N_13598,N_12621,N_12293);
nand U13599 (N_13599,N_12707,N_12113);
nand U13600 (N_13600,N_12845,N_13594);
nor U13601 (N_13601,N_13453,N_13539);
nand U13602 (N_13602,N_12912,N_13500);
nand U13603 (N_13603,N_12961,N_13231);
nand U13604 (N_13604,N_13236,N_13335);
nor U13605 (N_13605,N_12995,N_12887);
or U13606 (N_13606,N_13034,N_12896);
xnor U13607 (N_13607,N_13488,N_13502);
or U13608 (N_13608,N_13132,N_13061);
or U13609 (N_13609,N_13441,N_13406);
nor U13610 (N_13610,N_13079,N_13479);
nand U13611 (N_13611,N_13058,N_13420);
nand U13612 (N_13612,N_13591,N_13088);
xnor U13613 (N_13613,N_13509,N_13204);
or U13614 (N_13614,N_12944,N_12948);
nand U13615 (N_13615,N_13511,N_13538);
xor U13616 (N_13616,N_13366,N_12942);
xnor U13617 (N_13617,N_12842,N_13397);
xor U13618 (N_13618,N_13017,N_13575);
and U13619 (N_13619,N_13523,N_13573);
or U13620 (N_13620,N_13277,N_13427);
nand U13621 (N_13621,N_12837,N_12962);
xnor U13622 (N_13622,N_13183,N_13099);
and U13623 (N_13623,N_13542,N_13051);
nor U13624 (N_13624,N_13440,N_13197);
nand U13625 (N_13625,N_13592,N_13216);
nor U13626 (N_13626,N_13283,N_12919);
nand U13627 (N_13627,N_13493,N_13227);
or U13628 (N_13628,N_13124,N_13182);
and U13629 (N_13629,N_13329,N_13060);
nor U13630 (N_13630,N_12821,N_13087);
and U13631 (N_13631,N_13417,N_12983);
nand U13632 (N_13632,N_12931,N_12810);
nor U13633 (N_13633,N_13149,N_12903);
and U13634 (N_13634,N_12872,N_13378);
nand U13635 (N_13635,N_13258,N_13438);
xor U13636 (N_13636,N_13153,N_13497);
nand U13637 (N_13637,N_12823,N_12943);
or U13638 (N_13638,N_13314,N_13385);
or U13639 (N_13639,N_13540,N_12907);
nand U13640 (N_13640,N_12894,N_13095);
nand U13641 (N_13641,N_13167,N_13464);
xnor U13642 (N_13642,N_13190,N_13474);
and U13643 (N_13643,N_13478,N_13568);
nor U13644 (N_13644,N_12926,N_12885);
and U13645 (N_13645,N_13108,N_13173);
xor U13646 (N_13646,N_13485,N_12856);
and U13647 (N_13647,N_13131,N_13262);
or U13648 (N_13648,N_12970,N_13084);
and U13649 (N_13649,N_13271,N_13220);
and U13650 (N_13650,N_13097,N_13172);
and U13651 (N_13651,N_13282,N_13272);
or U13652 (N_13652,N_13424,N_13495);
or U13653 (N_13653,N_13400,N_13285);
xor U13654 (N_13654,N_13484,N_13143);
nor U13655 (N_13655,N_13574,N_13179);
nand U13656 (N_13656,N_13503,N_13462);
xor U13657 (N_13657,N_12922,N_13368);
nand U13658 (N_13658,N_13405,N_13319);
xor U13659 (N_13659,N_13013,N_12947);
and U13660 (N_13660,N_12828,N_12966);
and U13661 (N_13661,N_13007,N_13348);
or U13662 (N_13662,N_13294,N_12928);
and U13663 (N_13663,N_13344,N_13350);
xor U13664 (N_13664,N_13332,N_12997);
or U13665 (N_13665,N_13252,N_12801);
nand U13666 (N_13666,N_13198,N_12937);
nand U13667 (N_13667,N_13546,N_13508);
xnor U13668 (N_13668,N_12863,N_13189);
or U13669 (N_13669,N_13009,N_13414);
xor U13670 (N_13670,N_13171,N_12957);
and U13671 (N_13671,N_12831,N_12851);
and U13672 (N_13672,N_13284,N_12852);
nor U13673 (N_13673,N_12892,N_13138);
xnor U13674 (N_13674,N_12875,N_13073);
or U13675 (N_13675,N_13371,N_13290);
nand U13676 (N_13676,N_13191,N_13422);
xor U13677 (N_13677,N_12990,N_12822);
and U13678 (N_13678,N_12930,N_13547);
or U13679 (N_13679,N_13250,N_13524);
xnor U13680 (N_13680,N_13413,N_13244);
or U13681 (N_13681,N_13388,N_13137);
or U13682 (N_13682,N_13521,N_13567);
nor U13683 (N_13683,N_13025,N_12932);
xnor U13684 (N_13684,N_13450,N_13336);
and U13685 (N_13685,N_13040,N_13577);
and U13686 (N_13686,N_13031,N_13535);
or U13687 (N_13687,N_12844,N_13008);
and U13688 (N_13688,N_13286,N_13045);
nand U13689 (N_13689,N_13295,N_13161);
nand U13690 (N_13690,N_13558,N_13327);
and U13691 (N_13691,N_12946,N_13257);
xnor U13692 (N_13692,N_13349,N_12827);
xor U13693 (N_13693,N_13241,N_12871);
and U13694 (N_13694,N_12954,N_13014);
nor U13695 (N_13695,N_13486,N_13435);
and U13696 (N_13696,N_13576,N_12977);
xor U13697 (N_13697,N_13369,N_13202);
nand U13698 (N_13698,N_13207,N_13387);
and U13699 (N_13699,N_12803,N_13357);
nand U13700 (N_13700,N_13116,N_13548);
xor U13701 (N_13701,N_13482,N_13100);
nand U13702 (N_13702,N_13120,N_13126);
nor U13703 (N_13703,N_13180,N_12992);
xor U13704 (N_13704,N_12911,N_13447);
nand U13705 (N_13705,N_12830,N_13541);
or U13706 (N_13706,N_13028,N_13551);
and U13707 (N_13707,N_12979,N_13103);
and U13708 (N_13708,N_13468,N_13399);
or U13709 (N_13709,N_13062,N_13545);
and U13710 (N_13710,N_12935,N_13069);
xor U13711 (N_13711,N_12988,N_13586);
xor U13712 (N_13712,N_13054,N_13208);
nor U13713 (N_13713,N_13439,N_13597);
and U13714 (N_13714,N_12861,N_13364);
xnor U13715 (N_13715,N_13469,N_12860);
and U13716 (N_13716,N_12952,N_13141);
and U13717 (N_13717,N_13470,N_12834);
or U13718 (N_13718,N_13444,N_12960);
nand U13719 (N_13719,N_13326,N_13145);
nand U13720 (N_13720,N_13050,N_13032);
nor U13721 (N_13721,N_13472,N_13068);
nor U13722 (N_13722,N_12958,N_13359);
nor U13723 (N_13723,N_13264,N_12886);
or U13724 (N_13724,N_12987,N_13537);
nor U13725 (N_13725,N_12832,N_13076);
or U13726 (N_13726,N_13232,N_13446);
and U13727 (N_13727,N_13038,N_12913);
and U13728 (N_13728,N_13052,N_13063);
or U13729 (N_13729,N_13318,N_13499);
nor U13730 (N_13730,N_12806,N_12895);
or U13731 (N_13731,N_13254,N_12900);
or U13732 (N_13732,N_13455,N_13219);
xor U13733 (N_13733,N_13390,N_13561);
nand U13734 (N_13734,N_12804,N_13071);
and U13735 (N_13735,N_13527,N_13037);
nand U13736 (N_13736,N_13233,N_13275);
and U13737 (N_13737,N_13154,N_13181);
and U13738 (N_13738,N_13105,N_13041);
and U13739 (N_13739,N_12956,N_13454);
nor U13740 (N_13740,N_13238,N_13188);
nand U13741 (N_13741,N_13398,N_13312);
nor U13742 (N_13742,N_13057,N_13333);
nand U13743 (N_13743,N_12989,N_13315);
nand U13744 (N_13744,N_13448,N_13102);
nor U13745 (N_13745,N_13334,N_12853);
nand U13746 (N_13746,N_13529,N_13345);
xor U13747 (N_13747,N_13255,N_13512);
or U13748 (N_13748,N_13276,N_13491);
or U13749 (N_13749,N_13156,N_12884);
or U13750 (N_13750,N_12883,N_12864);
or U13751 (N_13751,N_13513,N_13532);
xnor U13752 (N_13752,N_13205,N_13465);
nor U13753 (N_13753,N_12951,N_13245);
and U13754 (N_13754,N_13303,N_13373);
nor U13755 (N_13755,N_13030,N_13270);
nand U13756 (N_13756,N_13432,N_12841);
and U13757 (N_13757,N_13248,N_13101);
nor U13758 (N_13758,N_13544,N_13367);
and U13759 (N_13759,N_13365,N_13408);
and U13760 (N_13760,N_12855,N_12921);
xor U13761 (N_13761,N_13409,N_13118);
and U13762 (N_13762,N_13055,N_13328);
or U13763 (N_13763,N_13112,N_13106);
nand U13764 (N_13764,N_13074,N_12980);
nand U13765 (N_13765,N_13123,N_13256);
xor U13766 (N_13766,N_13260,N_12850);
nand U13767 (N_13767,N_13155,N_13010);
and U13768 (N_13768,N_13184,N_12802);
nor U13769 (N_13769,N_13011,N_12874);
xnor U13770 (N_13770,N_13506,N_13178);
and U13771 (N_13771,N_13048,N_13117);
and U13772 (N_13772,N_13129,N_13237);
and U13773 (N_13773,N_12890,N_13199);
xor U13774 (N_13774,N_13466,N_13451);
nor U13775 (N_13775,N_13431,N_13266);
nand U13776 (N_13776,N_12899,N_12994);
nand U13777 (N_13777,N_13242,N_12865);
or U13778 (N_13778,N_13166,N_13163);
nand U13779 (N_13779,N_13046,N_13514);
nor U13780 (N_13780,N_12901,N_13426);
nand U13781 (N_13781,N_13002,N_13530);
or U13782 (N_13782,N_13082,N_13515);
or U13783 (N_13783,N_13235,N_12972);
xnor U13784 (N_13784,N_13249,N_12807);
nand U13785 (N_13785,N_12839,N_13428);
nor U13786 (N_13786,N_12924,N_12978);
and U13787 (N_13787,N_13125,N_13346);
or U13788 (N_13788,N_13293,N_13559);
nor U13789 (N_13789,N_13376,N_13392);
nor U13790 (N_13790,N_13377,N_12891);
xor U13791 (N_13791,N_13298,N_13351);
and U13792 (N_13792,N_13217,N_13430);
nand U13793 (N_13793,N_12859,N_12933);
nand U13794 (N_13794,N_13504,N_12829);
nand U13795 (N_13795,N_13300,N_12847);
and U13796 (N_13796,N_13218,N_13526);
or U13797 (N_13797,N_12976,N_13419);
nand U13798 (N_13798,N_12925,N_13096);
nand U13799 (N_13799,N_13114,N_12836);
and U13800 (N_13800,N_13104,N_13585);
nor U13801 (N_13801,N_13596,N_13077);
and U13802 (N_13802,N_13598,N_13549);
and U13803 (N_13803,N_13320,N_13085);
and U13804 (N_13804,N_12934,N_13304);
or U13805 (N_13805,N_13020,N_13222);
and U13806 (N_13806,N_13403,N_13589);
nand U13807 (N_13807,N_13361,N_13168);
and U13808 (N_13808,N_13310,N_13228);
nand U13809 (N_13809,N_13210,N_13311);
xnor U13810 (N_13810,N_13433,N_13239);
nand U13811 (N_13811,N_13317,N_13269);
nand U13812 (N_13812,N_12840,N_12953);
or U13813 (N_13813,N_13292,N_13569);
or U13814 (N_13814,N_13230,N_13563);
and U13815 (N_13815,N_13339,N_13572);
xnor U13816 (N_13816,N_13200,N_13380);
nor U13817 (N_13817,N_13595,N_12873);
nand U13818 (N_13818,N_13459,N_12941);
or U13819 (N_13819,N_12862,N_13552);
and U13820 (N_13820,N_13234,N_13225);
or U13821 (N_13821,N_13492,N_13289);
nand U13822 (N_13822,N_12868,N_13193);
nand U13823 (N_13823,N_13386,N_13423);
nand U13824 (N_13824,N_13044,N_13134);
nor U13825 (N_13825,N_13093,N_13185);
nand U13826 (N_13826,N_13473,N_13443);
xor U13827 (N_13827,N_13565,N_13246);
or U13828 (N_13828,N_13587,N_13065);
nand U13829 (N_13829,N_13324,N_13047);
and U13830 (N_13830,N_12969,N_12973);
xnor U13831 (N_13831,N_13562,N_12897);
xor U13832 (N_13832,N_13023,N_13480);
nor U13833 (N_13833,N_12824,N_13240);
nand U13834 (N_13834,N_12893,N_13458);
or U13835 (N_13835,N_13170,N_12870);
or U13836 (N_13836,N_13113,N_13056);
nand U13837 (N_13837,N_13186,N_13412);
and U13838 (N_13838,N_13461,N_13243);
nor U13839 (N_13839,N_13281,N_13554);
xor U13840 (N_13840,N_12917,N_12940);
xor U13841 (N_13841,N_13081,N_13313);
nor U13842 (N_13842,N_12800,N_13338);
xnor U13843 (N_13843,N_13078,N_13229);
or U13844 (N_13844,N_13533,N_13407);
xor U13845 (N_13845,N_13140,N_12880);
or U13846 (N_13846,N_12888,N_13261);
xor U13847 (N_13847,N_13247,N_13042);
and U13848 (N_13848,N_13582,N_13579);
or U13849 (N_13849,N_13507,N_13421);
nand U13850 (N_13850,N_12867,N_12858);
or U13851 (N_13851,N_13599,N_12843);
and U13852 (N_13852,N_13090,N_12878);
xnor U13853 (N_13853,N_13175,N_13353);
xor U13854 (N_13854,N_13445,N_13550);
nor U13855 (N_13855,N_12964,N_13330);
and U13856 (N_13856,N_13518,N_12945);
nand U13857 (N_13857,N_12811,N_13080);
or U13858 (N_13858,N_12986,N_13375);
or U13859 (N_13859,N_13165,N_12902);
and U13860 (N_13860,N_13035,N_13476);
or U13861 (N_13861,N_13018,N_12848);
nand U13862 (N_13862,N_13150,N_13274);
or U13863 (N_13863,N_13543,N_13416);
and U13864 (N_13864,N_12809,N_12805);
xnor U13865 (N_13865,N_12813,N_13026);
and U13866 (N_13866,N_12898,N_13340);
nand U13867 (N_13867,N_13160,N_13389);
nor U13868 (N_13868,N_13401,N_13012);
xnor U13869 (N_13869,N_13302,N_13323);
and U13870 (N_13870,N_13091,N_13158);
nor U13871 (N_13871,N_13590,N_12817);
or U13872 (N_13872,N_13307,N_13280);
or U13873 (N_13873,N_13463,N_13127);
xnor U13874 (N_13874,N_13593,N_13411);
nand U13875 (N_13875,N_13494,N_13206);
nor U13876 (N_13876,N_12906,N_13115);
and U13877 (N_13877,N_13209,N_13094);
nand U13878 (N_13878,N_13162,N_13434);
nand U13879 (N_13879,N_13049,N_13147);
nor U13880 (N_13880,N_13584,N_13251);
or U13881 (N_13881,N_13288,N_13152);
nor U13882 (N_13882,N_13267,N_13517);
nor U13883 (N_13883,N_13211,N_13005);
and U13884 (N_13884,N_13059,N_13296);
and U13885 (N_13885,N_13496,N_12869);
xor U13886 (N_13886,N_13301,N_12999);
and U13887 (N_13887,N_12910,N_13146);
or U13888 (N_13888,N_12905,N_13003);
nand U13889 (N_13889,N_13067,N_13291);
and U13890 (N_13890,N_12939,N_12959);
nor U13891 (N_13891,N_12876,N_12849);
nand U13892 (N_13892,N_13194,N_13107);
or U13893 (N_13893,N_13490,N_13070);
nand U13894 (N_13894,N_13425,N_13321);
and U13895 (N_13895,N_13528,N_13019);
and U13896 (N_13896,N_13477,N_13196);
nor U13897 (N_13897,N_12916,N_13557);
and U13898 (N_13898,N_13024,N_13265);
and U13899 (N_13899,N_13358,N_12838);
nor U13900 (N_13900,N_12981,N_13331);
or U13901 (N_13901,N_13157,N_13525);
nand U13902 (N_13902,N_13053,N_13570);
and U13903 (N_13903,N_13342,N_13043);
xor U13904 (N_13904,N_12820,N_12963);
nand U13905 (N_13905,N_13213,N_13212);
nor U13906 (N_13906,N_12854,N_13571);
xnor U13907 (N_13907,N_12982,N_13456);
nor U13908 (N_13908,N_12814,N_13418);
nand U13909 (N_13909,N_12826,N_12968);
xnor U13910 (N_13910,N_13027,N_12815);
or U13911 (N_13911,N_12998,N_13391);
nor U13912 (N_13912,N_12936,N_12904);
nand U13913 (N_13913,N_12975,N_13516);
xor U13914 (N_13914,N_13064,N_13487);
xnor U13915 (N_13915,N_13534,N_13393);
nor U13916 (N_13916,N_13223,N_13142);
xnor U13917 (N_13917,N_13159,N_13583);
nand U13918 (N_13918,N_13355,N_13483);
nand U13919 (N_13919,N_13467,N_13531);
nor U13920 (N_13920,N_13560,N_13263);
nor U13921 (N_13921,N_12929,N_13356);
nand U13922 (N_13922,N_13588,N_13133);
xor U13923 (N_13923,N_12974,N_13016);
xor U13924 (N_13924,N_13092,N_13384);
xor U13925 (N_13925,N_13164,N_12991);
nand U13926 (N_13926,N_13395,N_13214);
and U13927 (N_13927,N_13436,N_13501);
and U13928 (N_13928,N_12993,N_13151);
and U13929 (N_13929,N_13297,N_13457);
nand U13930 (N_13930,N_13410,N_13452);
and U13931 (N_13931,N_13268,N_13522);
or U13932 (N_13932,N_13475,N_13510);
and U13933 (N_13933,N_13402,N_13226);
or U13934 (N_13934,N_13354,N_13362);
or U13935 (N_13935,N_13083,N_13396);
or U13936 (N_13936,N_13273,N_13505);
nand U13937 (N_13937,N_13404,N_13121);
and U13938 (N_13938,N_13130,N_13253);
nand U13939 (N_13939,N_13429,N_12846);
and U13940 (N_13940,N_13122,N_13379);
xor U13941 (N_13941,N_13174,N_13039);
nand U13942 (N_13942,N_13111,N_13363);
and U13943 (N_13943,N_13308,N_12949);
nor U13944 (N_13944,N_13192,N_13177);
nor U13945 (N_13945,N_13144,N_13381);
and U13946 (N_13946,N_13520,N_13224);
xor U13947 (N_13947,N_13004,N_12927);
and U13948 (N_13948,N_13086,N_13415);
nand U13949 (N_13949,N_13098,N_13022);
or U13950 (N_13950,N_12833,N_13437);
and U13951 (N_13951,N_13578,N_12816);
or U13952 (N_13952,N_12923,N_13519);
nor U13953 (N_13953,N_13442,N_13259);
nor U13954 (N_13954,N_13460,N_13109);
nor U13955 (N_13955,N_12950,N_12818);
xnor U13956 (N_13956,N_12967,N_12889);
xnor U13957 (N_13957,N_13566,N_13119);
nor U13958 (N_13958,N_12857,N_13372);
nand U13959 (N_13959,N_12918,N_13341);
nand U13960 (N_13960,N_13136,N_12984);
nor U13961 (N_13961,N_13148,N_13169);
xnor U13962 (N_13962,N_13135,N_13449);
xor U13963 (N_13963,N_12881,N_13203);
xnor U13964 (N_13964,N_12877,N_13564);
nor U13965 (N_13965,N_12938,N_13343);
and U13966 (N_13966,N_13370,N_13581);
nand U13967 (N_13967,N_13481,N_12808);
nor U13968 (N_13968,N_13221,N_13553);
or U13969 (N_13969,N_13033,N_13382);
and U13970 (N_13970,N_13580,N_13089);
xnor U13971 (N_13971,N_13066,N_13316);
and U13972 (N_13972,N_13306,N_13128);
and U13973 (N_13973,N_12996,N_13021);
xnor U13974 (N_13974,N_13374,N_13278);
xor U13975 (N_13975,N_12909,N_13279);
and U13976 (N_13976,N_13489,N_12985);
nor U13977 (N_13977,N_13394,N_13036);
nor U13978 (N_13978,N_13187,N_13176);
xor U13979 (N_13979,N_12908,N_12920);
xnor U13980 (N_13980,N_13556,N_13555);
nor U13981 (N_13981,N_12879,N_13498);
or U13982 (N_13982,N_13139,N_12835);
xnor U13983 (N_13983,N_13337,N_12965);
xor U13984 (N_13984,N_13325,N_13029);
or U13985 (N_13985,N_13072,N_13215);
xnor U13986 (N_13986,N_12971,N_13322);
xnor U13987 (N_13987,N_13309,N_13536);
nor U13988 (N_13988,N_13001,N_13299);
or U13989 (N_13989,N_12914,N_13201);
xor U13990 (N_13990,N_12955,N_13015);
xnor U13991 (N_13991,N_12915,N_13471);
and U13992 (N_13992,N_12882,N_13383);
nor U13993 (N_13993,N_12819,N_12825);
or U13994 (N_13994,N_13110,N_13075);
nand U13995 (N_13995,N_12866,N_13000);
and U13996 (N_13996,N_12812,N_13352);
nand U13997 (N_13997,N_13347,N_13287);
nor U13998 (N_13998,N_13360,N_13305);
nor U13999 (N_13999,N_13006,N_13195);
and U14000 (N_14000,N_13421,N_13567);
xnor U14001 (N_14001,N_13597,N_13194);
nor U14002 (N_14002,N_13308,N_13232);
nand U14003 (N_14003,N_13062,N_13161);
nand U14004 (N_14004,N_13003,N_12926);
xor U14005 (N_14005,N_12837,N_13257);
nand U14006 (N_14006,N_13490,N_13594);
or U14007 (N_14007,N_13457,N_12918);
or U14008 (N_14008,N_13223,N_13112);
xnor U14009 (N_14009,N_13147,N_13365);
nor U14010 (N_14010,N_13587,N_13005);
xor U14011 (N_14011,N_13409,N_13470);
nor U14012 (N_14012,N_13344,N_13093);
xnor U14013 (N_14013,N_12822,N_13495);
nor U14014 (N_14014,N_13040,N_13154);
xor U14015 (N_14015,N_13013,N_12851);
xor U14016 (N_14016,N_13301,N_13363);
nand U14017 (N_14017,N_13278,N_13024);
and U14018 (N_14018,N_13535,N_13171);
nor U14019 (N_14019,N_13411,N_13497);
nand U14020 (N_14020,N_13155,N_12905);
nor U14021 (N_14021,N_13049,N_13577);
and U14022 (N_14022,N_13288,N_12813);
xor U14023 (N_14023,N_12954,N_12926);
and U14024 (N_14024,N_12904,N_13247);
nand U14025 (N_14025,N_12944,N_13292);
or U14026 (N_14026,N_13184,N_13150);
or U14027 (N_14027,N_13181,N_13454);
xnor U14028 (N_14028,N_13408,N_13286);
or U14029 (N_14029,N_13320,N_13454);
xor U14030 (N_14030,N_12970,N_12937);
or U14031 (N_14031,N_12953,N_13042);
nand U14032 (N_14032,N_13562,N_12866);
xnor U14033 (N_14033,N_13315,N_13327);
xnor U14034 (N_14034,N_13007,N_13403);
nor U14035 (N_14035,N_13173,N_13415);
nor U14036 (N_14036,N_12900,N_12816);
xor U14037 (N_14037,N_13355,N_12886);
and U14038 (N_14038,N_13256,N_13363);
nor U14039 (N_14039,N_13388,N_12928);
nand U14040 (N_14040,N_13100,N_12924);
nor U14041 (N_14041,N_13525,N_13359);
nor U14042 (N_14042,N_12951,N_13065);
nand U14043 (N_14043,N_13185,N_13108);
nor U14044 (N_14044,N_13539,N_13481);
and U14045 (N_14045,N_13435,N_12895);
xor U14046 (N_14046,N_12896,N_12998);
nor U14047 (N_14047,N_13311,N_13199);
nor U14048 (N_14048,N_13453,N_12879);
xnor U14049 (N_14049,N_13362,N_13556);
and U14050 (N_14050,N_13359,N_13317);
xnor U14051 (N_14051,N_13512,N_13338);
or U14052 (N_14052,N_13581,N_13560);
or U14053 (N_14053,N_13380,N_13067);
xor U14054 (N_14054,N_13146,N_13390);
nor U14055 (N_14055,N_12903,N_13233);
nor U14056 (N_14056,N_12888,N_13204);
or U14057 (N_14057,N_13198,N_13495);
nand U14058 (N_14058,N_13383,N_13438);
and U14059 (N_14059,N_12808,N_13418);
nor U14060 (N_14060,N_13086,N_13019);
nand U14061 (N_14061,N_13188,N_13290);
or U14062 (N_14062,N_13339,N_13416);
xnor U14063 (N_14063,N_12816,N_13284);
xor U14064 (N_14064,N_13256,N_13221);
and U14065 (N_14065,N_13050,N_12863);
nand U14066 (N_14066,N_13506,N_13293);
xor U14067 (N_14067,N_13134,N_13226);
nand U14068 (N_14068,N_13331,N_13350);
nand U14069 (N_14069,N_13460,N_13500);
and U14070 (N_14070,N_13546,N_13050);
nand U14071 (N_14071,N_12848,N_13590);
and U14072 (N_14072,N_12820,N_13334);
and U14073 (N_14073,N_13423,N_13095);
and U14074 (N_14074,N_12865,N_13265);
xor U14075 (N_14075,N_13031,N_13274);
nor U14076 (N_14076,N_13363,N_12806);
nand U14077 (N_14077,N_13175,N_13226);
or U14078 (N_14078,N_13265,N_13133);
nand U14079 (N_14079,N_12974,N_13310);
nand U14080 (N_14080,N_13253,N_13386);
xor U14081 (N_14081,N_13318,N_12987);
nand U14082 (N_14082,N_13054,N_13549);
nand U14083 (N_14083,N_13084,N_13019);
xor U14084 (N_14084,N_13594,N_12911);
or U14085 (N_14085,N_13172,N_13037);
and U14086 (N_14086,N_12971,N_13183);
and U14087 (N_14087,N_12989,N_13166);
or U14088 (N_14088,N_12855,N_13463);
xnor U14089 (N_14089,N_13543,N_13209);
and U14090 (N_14090,N_13439,N_13527);
nand U14091 (N_14091,N_13025,N_13101);
and U14092 (N_14092,N_13288,N_13415);
and U14093 (N_14093,N_12852,N_13339);
xor U14094 (N_14094,N_13327,N_12921);
nor U14095 (N_14095,N_12856,N_13527);
xnor U14096 (N_14096,N_13157,N_13127);
or U14097 (N_14097,N_13516,N_13509);
nor U14098 (N_14098,N_13432,N_13439);
and U14099 (N_14099,N_13164,N_13352);
and U14100 (N_14100,N_13346,N_13583);
nor U14101 (N_14101,N_12968,N_12923);
nand U14102 (N_14102,N_13157,N_13485);
nand U14103 (N_14103,N_13507,N_13138);
xnor U14104 (N_14104,N_13521,N_12839);
nand U14105 (N_14105,N_13347,N_13114);
xnor U14106 (N_14106,N_12812,N_13413);
nand U14107 (N_14107,N_13029,N_12914);
nor U14108 (N_14108,N_13452,N_13521);
and U14109 (N_14109,N_13470,N_12813);
or U14110 (N_14110,N_12934,N_12961);
xor U14111 (N_14111,N_13512,N_13389);
xnor U14112 (N_14112,N_13148,N_12870);
nor U14113 (N_14113,N_12817,N_13051);
nor U14114 (N_14114,N_13568,N_13493);
and U14115 (N_14115,N_12909,N_13578);
xnor U14116 (N_14116,N_12957,N_13337);
and U14117 (N_14117,N_13310,N_13235);
or U14118 (N_14118,N_12947,N_12853);
nand U14119 (N_14119,N_13528,N_13178);
nor U14120 (N_14120,N_12879,N_13229);
nand U14121 (N_14121,N_12812,N_13468);
xnor U14122 (N_14122,N_13082,N_13055);
and U14123 (N_14123,N_12927,N_12984);
and U14124 (N_14124,N_13415,N_12988);
nor U14125 (N_14125,N_13165,N_13463);
or U14126 (N_14126,N_13041,N_13508);
nand U14127 (N_14127,N_13025,N_13017);
nor U14128 (N_14128,N_12841,N_12969);
or U14129 (N_14129,N_13041,N_13278);
nand U14130 (N_14130,N_12835,N_12836);
nor U14131 (N_14131,N_13337,N_13373);
and U14132 (N_14132,N_13004,N_13423);
and U14133 (N_14133,N_13240,N_13006);
nand U14134 (N_14134,N_13218,N_13388);
or U14135 (N_14135,N_12964,N_13388);
and U14136 (N_14136,N_13268,N_13388);
nand U14137 (N_14137,N_13135,N_13229);
nand U14138 (N_14138,N_13021,N_13244);
nor U14139 (N_14139,N_13131,N_13488);
xor U14140 (N_14140,N_13176,N_13432);
xnor U14141 (N_14141,N_12957,N_13432);
or U14142 (N_14142,N_13354,N_13522);
and U14143 (N_14143,N_13155,N_12889);
nor U14144 (N_14144,N_12909,N_13408);
nor U14145 (N_14145,N_12959,N_13433);
or U14146 (N_14146,N_13321,N_12883);
or U14147 (N_14147,N_13334,N_13231);
nand U14148 (N_14148,N_12898,N_13104);
xnor U14149 (N_14149,N_12912,N_13434);
nor U14150 (N_14150,N_13276,N_12970);
and U14151 (N_14151,N_13044,N_12982);
nand U14152 (N_14152,N_13386,N_13113);
xor U14153 (N_14153,N_12833,N_12801);
nand U14154 (N_14154,N_13159,N_13274);
nor U14155 (N_14155,N_13071,N_13108);
or U14156 (N_14156,N_12887,N_12845);
nor U14157 (N_14157,N_12818,N_13037);
xnor U14158 (N_14158,N_13183,N_12951);
nor U14159 (N_14159,N_13446,N_13222);
and U14160 (N_14160,N_13566,N_13450);
or U14161 (N_14161,N_13514,N_13047);
or U14162 (N_14162,N_13176,N_13448);
and U14163 (N_14163,N_13405,N_13429);
or U14164 (N_14164,N_13563,N_13212);
or U14165 (N_14165,N_12812,N_12910);
xor U14166 (N_14166,N_13015,N_13218);
or U14167 (N_14167,N_13222,N_13286);
or U14168 (N_14168,N_13537,N_13379);
xnor U14169 (N_14169,N_13038,N_13547);
or U14170 (N_14170,N_13281,N_13585);
or U14171 (N_14171,N_13553,N_13568);
or U14172 (N_14172,N_12954,N_13462);
or U14173 (N_14173,N_13311,N_13271);
nand U14174 (N_14174,N_13342,N_12888);
nand U14175 (N_14175,N_13572,N_13252);
or U14176 (N_14176,N_12841,N_13220);
and U14177 (N_14177,N_13350,N_13473);
and U14178 (N_14178,N_13561,N_13251);
xnor U14179 (N_14179,N_13218,N_13485);
nand U14180 (N_14180,N_13232,N_13314);
or U14181 (N_14181,N_13286,N_13001);
or U14182 (N_14182,N_12886,N_12861);
or U14183 (N_14183,N_13156,N_12905);
or U14184 (N_14184,N_13163,N_13197);
and U14185 (N_14185,N_12943,N_13068);
xnor U14186 (N_14186,N_13202,N_13355);
or U14187 (N_14187,N_13196,N_13059);
and U14188 (N_14188,N_13254,N_12841);
nor U14189 (N_14189,N_13017,N_12878);
or U14190 (N_14190,N_13086,N_12975);
nand U14191 (N_14191,N_13475,N_12987);
nor U14192 (N_14192,N_12945,N_13275);
nor U14193 (N_14193,N_13595,N_13430);
nand U14194 (N_14194,N_13170,N_13024);
and U14195 (N_14195,N_12917,N_12882);
and U14196 (N_14196,N_13202,N_13215);
nor U14197 (N_14197,N_13065,N_12820);
and U14198 (N_14198,N_13557,N_12842);
xor U14199 (N_14199,N_13305,N_13211);
xor U14200 (N_14200,N_12922,N_12839);
xnor U14201 (N_14201,N_12902,N_13447);
nor U14202 (N_14202,N_13451,N_12905);
or U14203 (N_14203,N_13071,N_12958);
nand U14204 (N_14204,N_13194,N_13389);
and U14205 (N_14205,N_12944,N_13520);
nand U14206 (N_14206,N_12817,N_13492);
nand U14207 (N_14207,N_12880,N_12986);
nand U14208 (N_14208,N_12899,N_12803);
xnor U14209 (N_14209,N_13571,N_13223);
xnor U14210 (N_14210,N_13081,N_13495);
xnor U14211 (N_14211,N_13012,N_13389);
nor U14212 (N_14212,N_12934,N_13241);
xor U14213 (N_14213,N_13351,N_13562);
xor U14214 (N_14214,N_13420,N_13205);
nand U14215 (N_14215,N_13555,N_12815);
and U14216 (N_14216,N_12872,N_13567);
nand U14217 (N_14217,N_13142,N_13374);
xnor U14218 (N_14218,N_13248,N_13288);
xnor U14219 (N_14219,N_13459,N_13505);
and U14220 (N_14220,N_12821,N_13568);
nand U14221 (N_14221,N_13051,N_12877);
or U14222 (N_14222,N_12965,N_12803);
or U14223 (N_14223,N_13348,N_12908);
or U14224 (N_14224,N_13016,N_13443);
nand U14225 (N_14225,N_13316,N_12987);
xor U14226 (N_14226,N_13152,N_13467);
nand U14227 (N_14227,N_13197,N_13302);
and U14228 (N_14228,N_13307,N_13105);
xor U14229 (N_14229,N_13499,N_12861);
nand U14230 (N_14230,N_13461,N_13598);
nor U14231 (N_14231,N_12977,N_13488);
nand U14232 (N_14232,N_13455,N_13250);
xnor U14233 (N_14233,N_13304,N_13581);
nor U14234 (N_14234,N_13531,N_13170);
xnor U14235 (N_14235,N_13538,N_13514);
or U14236 (N_14236,N_13313,N_13294);
and U14237 (N_14237,N_13283,N_13100);
nand U14238 (N_14238,N_13482,N_12856);
nand U14239 (N_14239,N_13256,N_12910);
nor U14240 (N_14240,N_12916,N_13370);
nand U14241 (N_14241,N_13520,N_13473);
xnor U14242 (N_14242,N_13131,N_13220);
nor U14243 (N_14243,N_13290,N_13152);
nor U14244 (N_14244,N_13514,N_13511);
xnor U14245 (N_14245,N_13213,N_12912);
or U14246 (N_14246,N_13334,N_13046);
nand U14247 (N_14247,N_13541,N_13143);
nand U14248 (N_14248,N_13498,N_12807);
nor U14249 (N_14249,N_13433,N_12850);
nor U14250 (N_14250,N_13347,N_13498);
nand U14251 (N_14251,N_13260,N_13190);
and U14252 (N_14252,N_13420,N_12893);
nand U14253 (N_14253,N_13023,N_13519);
xor U14254 (N_14254,N_12806,N_13544);
nor U14255 (N_14255,N_12815,N_12933);
or U14256 (N_14256,N_13041,N_12873);
nand U14257 (N_14257,N_13159,N_13181);
nor U14258 (N_14258,N_12972,N_12837);
xnor U14259 (N_14259,N_13454,N_13259);
nor U14260 (N_14260,N_13318,N_13147);
or U14261 (N_14261,N_12970,N_13426);
xnor U14262 (N_14262,N_13432,N_12896);
xor U14263 (N_14263,N_12930,N_13086);
nor U14264 (N_14264,N_12866,N_13324);
and U14265 (N_14265,N_13532,N_13599);
xnor U14266 (N_14266,N_13379,N_12879);
nand U14267 (N_14267,N_13103,N_13186);
nor U14268 (N_14268,N_13356,N_13459);
xnor U14269 (N_14269,N_13557,N_13592);
nand U14270 (N_14270,N_12993,N_13015);
nor U14271 (N_14271,N_12819,N_13217);
and U14272 (N_14272,N_12945,N_13266);
and U14273 (N_14273,N_13081,N_12958);
nand U14274 (N_14274,N_13220,N_13183);
nand U14275 (N_14275,N_13369,N_13374);
or U14276 (N_14276,N_13270,N_12920);
nand U14277 (N_14277,N_13510,N_13181);
nor U14278 (N_14278,N_13091,N_13205);
nand U14279 (N_14279,N_13252,N_13256);
or U14280 (N_14280,N_13221,N_13549);
or U14281 (N_14281,N_13228,N_13283);
and U14282 (N_14282,N_13420,N_13161);
nand U14283 (N_14283,N_13414,N_12873);
nand U14284 (N_14284,N_13504,N_13327);
xnor U14285 (N_14285,N_13334,N_13225);
and U14286 (N_14286,N_13363,N_12975);
nor U14287 (N_14287,N_13420,N_13159);
or U14288 (N_14288,N_13278,N_13502);
and U14289 (N_14289,N_13589,N_12991);
and U14290 (N_14290,N_13109,N_13416);
and U14291 (N_14291,N_13075,N_12837);
nand U14292 (N_14292,N_13067,N_13120);
xnor U14293 (N_14293,N_13347,N_12802);
nor U14294 (N_14294,N_13281,N_13131);
or U14295 (N_14295,N_12811,N_13269);
and U14296 (N_14296,N_13594,N_13241);
nand U14297 (N_14297,N_13298,N_13311);
and U14298 (N_14298,N_13465,N_13509);
and U14299 (N_14299,N_13100,N_12859);
and U14300 (N_14300,N_13153,N_13019);
and U14301 (N_14301,N_13500,N_13525);
nor U14302 (N_14302,N_13571,N_13382);
xnor U14303 (N_14303,N_13443,N_12821);
nor U14304 (N_14304,N_13551,N_13025);
or U14305 (N_14305,N_12958,N_13342);
xor U14306 (N_14306,N_13294,N_13062);
nor U14307 (N_14307,N_12940,N_13028);
and U14308 (N_14308,N_13534,N_13218);
nand U14309 (N_14309,N_13232,N_13352);
nand U14310 (N_14310,N_12921,N_13141);
nand U14311 (N_14311,N_13450,N_12954);
and U14312 (N_14312,N_13415,N_13111);
nand U14313 (N_14313,N_13122,N_13530);
nand U14314 (N_14314,N_13272,N_13138);
nor U14315 (N_14315,N_13194,N_12813);
nor U14316 (N_14316,N_13001,N_12931);
or U14317 (N_14317,N_13337,N_12971);
nor U14318 (N_14318,N_13267,N_13359);
or U14319 (N_14319,N_13400,N_13346);
or U14320 (N_14320,N_12981,N_13360);
nand U14321 (N_14321,N_13393,N_13320);
xnor U14322 (N_14322,N_12818,N_13528);
nor U14323 (N_14323,N_13427,N_12904);
xor U14324 (N_14324,N_13192,N_13103);
or U14325 (N_14325,N_12999,N_13527);
nand U14326 (N_14326,N_13177,N_13255);
nor U14327 (N_14327,N_13500,N_13459);
nand U14328 (N_14328,N_13448,N_13592);
nor U14329 (N_14329,N_12804,N_13310);
and U14330 (N_14330,N_13342,N_13008);
xor U14331 (N_14331,N_13232,N_12979);
nand U14332 (N_14332,N_13248,N_13100);
or U14333 (N_14333,N_13325,N_13267);
nand U14334 (N_14334,N_13151,N_13273);
xor U14335 (N_14335,N_13352,N_12890);
nor U14336 (N_14336,N_13079,N_13335);
and U14337 (N_14337,N_13324,N_13272);
or U14338 (N_14338,N_13133,N_13481);
or U14339 (N_14339,N_13585,N_13319);
nor U14340 (N_14340,N_12934,N_12859);
and U14341 (N_14341,N_13191,N_12814);
and U14342 (N_14342,N_13230,N_13181);
nand U14343 (N_14343,N_13268,N_13022);
and U14344 (N_14344,N_13152,N_13315);
xor U14345 (N_14345,N_12979,N_13049);
xor U14346 (N_14346,N_12976,N_13593);
or U14347 (N_14347,N_13102,N_12841);
nor U14348 (N_14348,N_12828,N_12980);
xor U14349 (N_14349,N_13011,N_13349);
nor U14350 (N_14350,N_12840,N_13065);
and U14351 (N_14351,N_13059,N_13271);
or U14352 (N_14352,N_13589,N_13141);
xor U14353 (N_14353,N_13300,N_13533);
or U14354 (N_14354,N_13367,N_13520);
xor U14355 (N_14355,N_13201,N_12833);
nand U14356 (N_14356,N_13179,N_13513);
nand U14357 (N_14357,N_12969,N_13125);
or U14358 (N_14358,N_12827,N_13428);
or U14359 (N_14359,N_13561,N_12897);
xor U14360 (N_14360,N_13492,N_13419);
nand U14361 (N_14361,N_13524,N_13442);
xnor U14362 (N_14362,N_13347,N_13098);
xnor U14363 (N_14363,N_12813,N_13243);
xnor U14364 (N_14364,N_13344,N_13430);
xnor U14365 (N_14365,N_13242,N_13516);
xnor U14366 (N_14366,N_13075,N_13425);
nor U14367 (N_14367,N_13043,N_12956);
or U14368 (N_14368,N_13440,N_13042);
nor U14369 (N_14369,N_12809,N_13383);
xnor U14370 (N_14370,N_13321,N_13561);
xor U14371 (N_14371,N_13481,N_13112);
or U14372 (N_14372,N_13585,N_13595);
and U14373 (N_14373,N_13373,N_12826);
xor U14374 (N_14374,N_12954,N_13387);
nand U14375 (N_14375,N_13223,N_13091);
and U14376 (N_14376,N_12804,N_13598);
or U14377 (N_14377,N_13364,N_13039);
nand U14378 (N_14378,N_12908,N_13408);
or U14379 (N_14379,N_13558,N_12820);
or U14380 (N_14380,N_13557,N_12957);
or U14381 (N_14381,N_13035,N_13559);
nor U14382 (N_14382,N_13381,N_13187);
nand U14383 (N_14383,N_12942,N_12890);
or U14384 (N_14384,N_13016,N_13284);
nor U14385 (N_14385,N_13416,N_12884);
nor U14386 (N_14386,N_13278,N_13507);
nor U14387 (N_14387,N_13298,N_13201);
xnor U14388 (N_14388,N_13436,N_13155);
nand U14389 (N_14389,N_13150,N_13346);
xnor U14390 (N_14390,N_12911,N_13095);
nand U14391 (N_14391,N_13502,N_13163);
nor U14392 (N_14392,N_13196,N_13527);
xnor U14393 (N_14393,N_13451,N_13569);
and U14394 (N_14394,N_13479,N_13217);
nand U14395 (N_14395,N_13282,N_13095);
nand U14396 (N_14396,N_13066,N_13430);
nor U14397 (N_14397,N_13489,N_13396);
and U14398 (N_14398,N_13238,N_13223);
xor U14399 (N_14399,N_13522,N_13327);
xor U14400 (N_14400,N_14349,N_13959);
and U14401 (N_14401,N_13732,N_14221);
xnor U14402 (N_14402,N_13634,N_13973);
nor U14403 (N_14403,N_13932,N_13798);
xnor U14404 (N_14404,N_14172,N_13906);
nand U14405 (N_14405,N_13686,N_13640);
nor U14406 (N_14406,N_13760,N_13872);
nor U14407 (N_14407,N_13990,N_13968);
nor U14408 (N_14408,N_14034,N_14330);
nand U14409 (N_14409,N_14387,N_14320);
or U14410 (N_14410,N_14323,N_14268);
nor U14411 (N_14411,N_14321,N_14051);
nand U14412 (N_14412,N_14350,N_13832);
or U14413 (N_14413,N_13621,N_13977);
nand U14414 (N_14414,N_13703,N_14252);
or U14415 (N_14415,N_13883,N_13894);
and U14416 (N_14416,N_14041,N_13769);
nand U14417 (N_14417,N_13945,N_13706);
nand U14418 (N_14418,N_14114,N_13645);
and U14419 (N_14419,N_14284,N_13698);
xor U14420 (N_14420,N_13765,N_13991);
nand U14421 (N_14421,N_14100,N_13814);
nand U14422 (N_14422,N_14087,N_13925);
or U14423 (N_14423,N_14331,N_14125);
and U14424 (N_14424,N_14327,N_14032);
nand U14425 (N_14425,N_14245,N_13752);
or U14426 (N_14426,N_13862,N_14399);
nand U14427 (N_14427,N_14202,N_13902);
nor U14428 (N_14428,N_13777,N_13944);
or U14429 (N_14429,N_14184,N_14255);
and U14430 (N_14430,N_14074,N_13723);
nand U14431 (N_14431,N_13705,N_13685);
nor U14432 (N_14432,N_14324,N_14296);
nor U14433 (N_14433,N_14262,N_14118);
xor U14434 (N_14434,N_13728,N_13984);
or U14435 (N_14435,N_13919,N_13650);
nand U14436 (N_14436,N_13840,N_14061);
nor U14437 (N_14437,N_14369,N_14231);
nand U14438 (N_14438,N_14383,N_13873);
and U14439 (N_14439,N_13940,N_13829);
xnor U14440 (N_14440,N_13763,N_13641);
xnor U14441 (N_14441,N_14215,N_13605);
or U14442 (N_14442,N_13976,N_14028);
and U14443 (N_14443,N_13877,N_14169);
nor U14444 (N_14444,N_14097,N_13904);
nor U14445 (N_14445,N_14133,N_13921);
nand U14446 (N_14446,N_13682,N_14137);
xnor U14447 (N_14447,N_14220,N_13871);
xor U14448 (N_14448,N_14025,N_13632);
nor U14449 (N_14449,N_14354,N_14057);
and U14450 (N_14450,N_13701,N_13813);
and U14451 (N_14451,N_13787,N_13941);
or U14452 (N_14452,N_14076,N_14176);
or U14453 (N_14453,N_14195,N_13947);
and U14454 (N_14454,N_14364,N_13891);
or U14455 (N_14455,N_13931,N_13649);
nand U14456 (N_14456,N_13998,N_13954);
and U14457 (N_14457,N_13960,N_13714);
and U14458 (N_14458,N_13850,N_13958);
or U14459 (N_14459,N_13673,N_13799);
nor U14460 (N_14460,N_14388,N_13766);
xor U14461 (N_14461,N_14197,N_14222);
nor U14462 (N_14462,N_13979,N_14166);
and U14463 (N_14463,N_14015,N_13914);
and U14464 (N_14464,N_13704,N_14048);
nor U14465 (N_14465,N_13881,N_14157);
or U14466 (N_14466,N_14343,N_14375);
and U14467 (N_14467,N_14187,N_13803);
xor U14468 (N_14468,N_13992,N_14049);
nor U14469 (N_14469,N_13750,N_14185);
nor U14470 (N_14470,N_14148,N_13729);
nand U14471 (N_14471,N_13933,N_13806);
or U14472 (N_14472,N_14248,N_13671);
or U14473 (N_14473,N_14194,N_13631);
or U14474 (N_14474,N_14386,N_13892);
or U14475 (N_14475,N_13989,N_13694);
nand U14476 (N_14476,N_14122,N_14113);
or U14477 (N_14477,N_13737,N_13863);
and U14478 (N_14478,N_13884,N_13642);
and U14479 (N_14479,N_13983,N_14203);
xnor U14480 (N_14480,N_13784,N_14012);
nand U14481 (N_14481,N_14062,N_14358);
nor U14482 (N_14482,N_14075,N_13950);
or U14483 (N_14483,N_14380,N_14177);
nor U14484 (N_14484,N_14211,N_13845);
xor U14485 (N_14485,N_14193,N_14339);
or U14486 (N_14486,N_14348,N_13629);
nor U14487 (N_14487,N_14163,N_14003);
or U14488 (N_14488,N_14290,N_13609);
nand U14489 (N_14489,N_13851,N_14225);
xnor U14490 (N_14490,N_13779,N_14037);
or U14491 (N_14491,N_13660,N_13889);
xnor U14492 (N_14492,N_14238,N_14355);
nor U14493 (N_14493,N_13712,N_14066);
or U14494 (N_14494,N_13827,N_13690);
nor U14495 (N_14495,N_13697,N_14035);
and U14496 (N_14496,N_13721,N_13710);
or U14497 (N_14497,N_14232,N_13612);
and U14498 (N_14498,N_14138,N_13953);
nor U14499 (N_14499,N_13790,N_14067);
nor U14500 (N_14500,N_13775,N_14344);
and U14501 (N_14501,N_14322,N_14289);
nor U14502 (N_14502,N_13819,N_14024);
nand U14503 (N_14503,N_13951,N_13773);
nand U14504 (N_14504,N_13949,N_13659);
and U14505 (N_14505,N_14340,N_13653);
nand U14506 (N_14506,N_14240,N_14173);
and U14507 (N_14507,N_14207,N_14116);
nor U14508 (N_14508,N_14335,N_13742);
and U14509 (N_14509,N_14283,N_14261);
and U14510 (N_14510,N_14381,N_13600);
or U14511 (N_14511,N_13980,N_14079);
nor U14512 (N_14512,N_14115,N_14027);
nor U14513 (N_14513,N_13797,N_13874);
and U14514 (N_14514,N_13836,N_14101);
and U14515 (N_14515,N_13746,N_13822);
or U14516 (N_14516,N_13607,N_13610);
xor U14517 (N_14517,N_13994,N_13665);
xor U14518 (N_14518,N_13808,N_14056);
nand U14519 (N_14519,N_14300,N_14250);
nand U14520 (N_14520,N_13739,N_13804);
xor U14521 (N_14521,N_13655,N_14174);
or U14522 (N_14522,N_13776,N_13727);
xnor U14523 (N_14523,N_14013,N_14178);
and U14524 (N_14524,N_14314,N_13608);
or U14525 (N_14525,N_14058,N_14069);
nor U14526 (N_14526,N_14368,N_14246);
and U14527 (N_14527,N_14165,N_14191);
or U14528 (N_14528,N_13651,N_14351);
xor U14529 (N_14529,N_14376,N_14162);
and U14530 (N_14530,N_14094,N_13708);
nand U14531 (N_14531,N_13834,N_14171);
and U14532 (N_14532,N_14229,N_14189);
nor U14533 (N_14533,N_13666,N_14153);
or U14534 (N_14534,N_13692,N_14070);
nor U14535 (N_14535,N_14111,N_14291);
or U14536 (N_14536,N_13809,N_13859);
and U14537 (N_14537,N_13759,N_14391);
nand U14538 (N_14538,N_14019,N_13890);
nor U14539 (N_14539,N_14316,N_13611);
nand U14540 (N_14540,N_14333,N_14210);
nor U14541 (N_14541,N_13741,N_14313);
xnor U14542 (N_14542,N_14009,N_13887);
nor U14543 (N_14543,N_14382,N_13757);
nor U14544 (N_14544,N_14083,N_14272);
or U14545 (N_14545,N_14136,N_14361);
nor U14546 (N_14546,N_13747,N_13606);
nand U14547 (N_14547,N_13816,N_13870);
nor U14548 (N_14548,N_14149,N_14288);
and U14549 (N_14549,N_13886,N_14298);
and U14550 (N_14550,N_14275,N_13643);
or U14551 (N_14551,N_13963,N_14164);
nand U14552 (N_14552,N_14346,N_14055);
and U14553 (N_14553,N_13791,N_14328);
nand U14554 (N_14554,N_14278,N_13969);
nor U14555 (N_14555,N_13602,N_14104);
nor U14556 (N_14556,N_13975,N_14373);
nor U14557 (N_14557,N_14224,N_13996);
nand U14558 (N_14558,N_14047,N_13811);
and U14559 (N_14559,N_13821,N_13616);
or U14560 (N_14560,N_13864,N_13943);
nor U14561 (N_14561,N_14198,N_14200);
nand U14562 (N_14562,N_14085,N_13825);
xor U14563 (N_14563,N_13674,N_13652);
or U14564 (N_14564,N_14030,N_14060);
xor U14565 (N_14565,N_14170,N_13658);
or U14566 (N_14566,N_13824,N_14239);
and U14567 (N_14567,N_13619,N_13693);
nand U14568 (N_14568,N_13920,N_14352);
nor U14569 (N_14569,N_13852,N_14129);
nand U14570 (N_14570,N_13835,N_13810);
and U14571 (N_14571,N_14134,N_13638);
nand U14572 (N_14572,N_13930,N_14293);
nand U14573 (N_14573,N_13644,N_14216);
nor U14574 (N_14574,N_14086,N_14160);
xor U14575 (N_14575,N_14254,N_13856);
and U14576 (N_14576,N_13720,N_14117);
or U14577 (N_14577,N_13869,N_14398);
or U14578 (N_14578,N_14108,N_14167);
nor U14579 (N_14579,N_13965,N_13987);
nor U14580 (N_14580,N_13668,N_13722);
xor U14581 (N_14581,N_14265,N_13966);
nand U14582 (N_14582,N_13725,N_13962);
and U14583 (N_14583,N_14384,N_13699);
or U14584 (N_14584,N_13942,N_14217);
nor U14585 (N_14585,N_14237,N_14154);
and U14586 (N_14586,N_14226,N_13795);
xnor U14587 (N_14587,N_13857,N_14110);
nand U14588 (N_14588,N_13833,N_13826);
xor U14589 (N_14589,N_14139,N_13711);
and U14590 (N_14590,N_13922,N_14236);
nor U14591 (N_14591,N_14277,N_13663);
xnor U14592 (N_14592,N_13839,N_14078);
and U14593 (N_14593,N_13885,N_13937);
nor U14594 (N_14594,N_14001,N_13648);
xnor U14595 (N_14595,N_14181,N_14018);
xor U14596 (N_14596,N_14367,N_13923);
or U14597 (N_14597,N_14031,N_13783);
xor U14598 (N_14598,N_14371,N_14159);
and U14599 (N_14599,N_14287,N_14183);
nor U14600 (N_14600,N_13624,N_14093);
and U14601 (N_14601,N_13772,N_14353);
nor U14602 (N_14602,N_13743,N_13604);
xnor U14603 (N_14603,N_14228,N_13781);
and U14604 (N_14604,N_13646,N_13709);
and U14605 (N_14605,N_14276,N_14190);
and U14606 (N_14606,N_14071,N_14064);
or U14607 (N_14607,N_13639,N_14044);
and U14608 (N_14608,N_14068,N_13952);
or U14609 (N_14609,N_13789,N_14090);
xor U14610 (N_14610,N_14038,N_14092);
nand U14611 (N_14611,N_14305,N_14311);
nand U14612 (N_14612,N_13730,N_14251);
nor U14613 (N_14613,N_13867,N_14362);
nor U14614 (N_14614,N_13897,N_14192);
nor U14615 (N_14615,N_14266,N_14196);
and U14616 (N_14616,N_13844,N_14107);
nand U14617 (N_14617,N_13613,N_14043);
or U14618 (N_14618,N_13736,N_14292);
and U14619 (N_14619,N_13936,N_13748);
xor U14620 (N_14620,N_13848,N_14127);
and U14621 (N_14621,N_13918,N_14106);
or U14622 (N_14622,N_14235,N_14036);
xor U14623 (N_14623,N_14046,N_13695);
or U14624 (N_14624,N_13893,N_13909);
xor U14625 (N_14625,N_13929,N_13903);
nand U14626 (N_14626,N_13688,N_14243);
nor U14627 (N_14627,N_14161,N_14084);
xor U14628 (N_14628,N_14285,N_14374);
and U14629 (N_14629,N_14098,N_14033);
nand U14630 (N_14630,N_13786,N_13702);
and U14631 (N_14631,N_13785,N_14007);
or U14632 (N_14632,N_13995,N_14135);
and U14633 (N_14633,N_13882,N_13738);
nor U14634 (N_14634,N_14014,N_14319);
nand U14635 (N_14635,N_13715,N_14312);
xor U14636 (N_14636,N_14155,N_14023);
xnor U14637 (N_14637,N_14310,N_13934);
or U14638 (N_14638,N_14188,N_14103);
nor U14639 (N_14639,N_13675,N_14010);
nand U14640 (N_14640,N_13627,N_14325);
xnor U14641 (N_14641,N_13768,N_13830);
and U14642 (N_14642,N_13788,N_14112);
xor U14643 (N_14643,N_14377,N_13916);
xnor U14644 (N_14644,N_14124,N_14363);
or U14645 (N_14645,N_13978,N_14179);
xor U14646 (N_14646,N_13878,N_13900);
xor U14647 (N_14647,N_13719,N_13672);
and U14648 (N_14648,N_13967,N_13735);
nor U14649 (N_14649,N_14021,N_13875);
and U14650 (N_14650,N_14204,N_13837);
nor U14651 (N_14651,N_13861,N_13865);
and U14652 (N_14652,N_13841,N_14152);
and U14653 (N_14653,N_14294,N_13946);
nor U14654 (N_14654,N_14315,N_13796);
or U14655 (N_14655,N_13948,N_13630);
or U14656 (N_14656,N_14141,N_13774);
and U14657 (N_14657,N_14281,N_13726);
nand U14658 (N_14658,N_13689,N_13667);
xnor U14659 (N_14659,N_13876,N_13761);
or U14660 (N_14660,N_14360,N_14280);
and U14661 (N_14661,N_14218,N_13792);
and U14662 (N_14662,N_13917,N_14230);
or U14663 (N_14663,N_14008,N_14233);
xor U14664 (N_14664,N_14000,N_14273);
nand U14665 (N_14665,N_13749,N_14279);
nand U14666 (N_14666,N_14282,N_13681);
and U14667 (N_14667,N_14227,N_14372);
nor U14668 (N_14668,N_14247,N_14342);
nor U14669 (N_14669,N_14267,N_14143);
nor U14670 (N_14670,N_14081,N_13854);
nor U14671 (N_14671,N_14214,N_13647);
nand U14672 (N_14672,N_14208,N_13764);
xor U14673 (N_14673,N_13683,N_13615);
nor U14674 (N_14674,N_14253,N_13620);
and U14675 (N_14675,N_13676,N_14026);
or U14676 (N_14676,N_13707,N_14004);
or U14677 (N_14677,N_13853,N_13617);
nor U14678 (N_14678,N_13997,N_14053);
and U14679 (N_14679,N_13927,N_14303);
or U14680 (N_14680,N_14379,N_13679);
nand U14681 (N_14681,N_14274,N_14209);
xor U14682 (N_14682,N_14389,N_14102);
xnor U14683 (N_14683,N_13637,N_13982);
xnor U14684 (N_14684,N_14120,N_13911);
or U14685 (N_14685,N_14073,N_14199);
xnor U14686 (N_14686,N_13678,N_13993);
or U14687 (N_14687,N_14270,N_13910);
or U14688 (N_14688,N_14175,N_14308);
and U14689 (N_14689,N_13623,N_13670);
or U14690 (N_14690,N_13912,N_14397);
and U14691 (N_14691,N_14045,N_14182);
nand U14692 (N_14692,N_14006,N_14302);
nor U14693 (N_14693,N_14334,N_13802);
xnor U14694 (N_14694,N_13831,N_14356);
xnor U14695 (N_14695,N_14304,N_14017);
or U14696 (N_14696,N_13661,N_13888);
nor U14697 (N_14697,N_13855,N_13635);
nor U14698 (N_14698,N_14365,N_14260);
or U14699 (N_14699,N_14258,N_13972);
and U14700 (N_14700,N_14307,N_14295);
or U14701 (N_14701,N_13771,N_14123);
nand U14702 (N_14702,N_14130,N_14151);
nor U14703 (N_14703,N_13986,N_13849);
nor U14704 (N_14704,N_14040,N_14180);
nand U14705 (N_14705,N_14002,N_14326);
or U14706 (N_14706,N_14011,N_13842);
xor U14707 (N_14707,N_14234,N_13907);
nor U14708 (N_14708,N_14242,N_14054);
and U14709 (N_14709,N_14206,N_14145);
and U14710 (N_14710,N_13751,N_13731);
xor U14711 (N_14711,N_14140,N_13956);
xor U14712 (N_14712,N_14052,N_13734);
xor U14713 (N_14713,N_13793,N_14016);
or U14714 (N_14714,N_13981,N_13970);
nor U14715 (N_14715,N_14119,N_14212);
nor U14716 (N_14716,N_13618,N_14395);
nand U14717 (N_14717,N_13823,N_13905);
nand U14718 (N_14718,N_13988,N_14394);
and U14719 (N_14719,N_13801,N_13654);
nand U14720 (N_14720,N_13964,N_13664);
xnor U14721 (N_14721,N_13955,N_13669);
or U14722 (N_14722,N_13755,N_13717);
nor U14723 (N_14723,N_14082,N_13908);
nand U14724 (N_14724,N_13778,N_14091);
nand U14725 (N_14725,N_14099,N_13636);
nand U14726 (N_14726,N_13744,N_14357);
xor U14727 (N_14727,N_13691,N_13767);
nand U14728 (N_14728,N_14039,N_13985);
or U14729 (N_14729,N_14338,N_13762);
and U14730 (N_14730,N_13895,N_14020);
nor U14731 (N_14731,N_14144,N_13713);
xor U14732 (N_14732,N_14109,N_14244);
nand U14733 (N_14733,N_14347,N_14150);
nor U14734 (N_14734,N_13622,N_14299);
or U14735 (N_14735,N_14128,N_14105);
nor U14736 (N_14736,N_14345,N_13662);
xor U14737 (N_14737,N_14142,N_13724);
or U14738 (N_14738,N_14050,N_14259);
or U14739 (N_14739,N_13733,N_14146);
nand U14740 (N_14740,N_13858,N_13999);
and U14741 (N_14741,N_13935,N_14089);
and U14742 (N_14742,N_14329,N_14059);
nand U14743 (N_14743,N_13782,N_13847);
xnor U14744 (N_14744,N_14005,N_13939);
nand U14745 (N_14745,N_14223,N_13800);
and U14746 (N_14746,N_14186,N_14359);
or U14747 (N_14747,N_14095,N_13901);
and U14748 (N_14748,N_13812,N_14392);
nand U14749 (N_14749,N_13626,N_13716);
nor U14750 (N_14750,N_14306,N_13913);
nand U14751 (N_14751,N_13625,N_14256);
xnor U14752 (N_14752,N_14131,N_13656);
xor U14753 (N_14753,N_14309,N_14088);
xnor U14754 (N_14754,N_13807,N_14126);
and U14755 (N_14755,N_14201,N_13794);
or U14756 (N_14756,N_14213,N_13770);
xnor U14757 (N_14757,N_14096,N_13601);
or U14758 (N_14758,N_14219,N_14147);
nor U14759 (N_14759,N_14257,N_13879);
nand U14760 (N_14760,N_14378,N_13696);
xor U14761 (N_14761,N_14132,N_13818);
nand U14762 (N_14762,N_13880,N_13718);
nor U14763 (N_14763,N_14332,N_14366);
and U14764 (N_14764,N_13971,N_14249);
and U14765 (N_14765,N_14390,N_14317);
or U14766 (N_14766,N_13846,N_13820);
nor U14767 (N_14767,N_14370,N_14029);
nand U14768 (N_14768,N_14063,N_13633);
nand U14769 (N_14769,N_13899,N_13817);
nand U14770 (N_14770,N_14077,N_13815);
nor U14771 (N_14771,N_14337,N_14121);
nand U14772 (N_14772,N_13700,N_13805);
xnor U14773 (N_14773,N_13680,N_14156);
and U14774 (N_14774,N_13915,N_13928);
nand U14775 (N_14775,N_13974,N_13843);
xor U14776 (N_14776,N_13868,N_13753);
xnor U14777 (N_14777,N_14022,N_13684);
or U14778 (N_14778,N_14271,N_13866);
nand U14779 (N_14779,N_14065,N_13780);
or U14780 (N_14780,N_14269,N_13924);
xor U14781 (N_14781,N_13957,N_13677);
or U14782 (N_14782,N_14042,N_13860);
nor U14783 (N_14783,N_14297,N_14072);
nand U14784 (N_14784,N_13628,N_13828);
and U14785 (N_14785,N_14385,N_14264);
nor U14786 (N_14786,N_14286,N_14168);
or U14787 (N_14787,N_13898,N_14205);
nand U14788 (N_14788,N_13603,N_14318);
nor U14789 (N_14789,N_14396,N_13754);
or U14790 (N_14790,N_14080,N_13756);
and U14791 (N_14791,N_14341,N_14301);
nand U14792 (N_14792,N_14393,N_13938);
nor U14793 (N_14793,N_13657,N_13896);
nor U14794 (N_14794,N_14336,N_14263);
or U14795 (N_14795,N_14241,N_13740);
xnor U14796 (N_14796,N_13838,N_13614);
nor U14797 (N_14797,N_13961,N_13758);
and U14798 (N_14798,N_13687,N_13926);
nand U14799 (N_14799,N_14158,N_13745);
or U14800 (N_14800,N_13672,N_14291);
or U14801 (N_14801,N_13950,N_14067);
nor U14802 (N_14802,N_13976,N_13633);
nand U14803 (N_14803,N_13947,N_14148);
or U14804 (N_14804,N_13797,N_13991);
nand U14805 (N_14805,N_14225,N_13965);
nand U14806 (N_14806,N_13755,N_13870);
xor U14807 (N_14807,N_13942,N_14166);
nor U14808 (N_14808,N_13802,N_13853);
nor U14809 (N_14809,N_14107,N_14162);
nand U14810 (N_14810,N_14250,N_14024);
and U14811 (N_14811,N_14255,N_14348);
nor U14812 (N_14812,N_13891,N_13657);
xor U14813 (N_14813,N_13654,N_14138);
nand U14814 (N_14814,N_13757,N_13984);
or U14815 (N_14815,N_13752,N_13814);
nor U14816 (N_14816,N_14156,N_14203);
nor U14817 (N_14817,N_14027,N_13654);
nor U14818 (N_14818,N_13857,N_14059);
xnor U14819 (N_14819,N_14361,N_14001);
nand U14820 (N_14820,N_13672,N_13753);
xnor U14821 (N_14821,N_14109,N_14359);
nand U14822 (N_14822,N_13840,N_13676);
and U14823 (N_14823,N_13850,N_13983);
and U14824 (N_14824,N_14216,N_14161);
or U14825 (N_14825,N_14397,N_14362);
or U14826 (N_14826,N_13854,N_13691);
nand U14827 (N_14827,N_14348,N_13766);
or U14828 (N_14828,N_14320,N_14013);
nand U14829 (N_14829,N_14206,N_14179);
xor U14830 (N_14830,N_13704,N_14279);
nand U14831 (N_14831,N_14071,N_14062);
nand U14832 (N_14832,N_14179,N_14295);
and U14833 (N_14833,N_13736,N_14047);
nor U14834 (N_14834,N_13766,N_13661);
and U14835 (N_14835,N_14029,N_14049);
xor U14836 (N_14836,N_13856,N_14214);
or U14837 (N_14837,N_13717,N_14123);
nand U14838 (N_14838,N_13816,N_14054);
nand U14839 (N_14839,N_14147,N_14088);
xnor U14840 (N_14840,N_13887,N_13766);
xor U14841 (N_14841,N_13822,N_14196);
nand U14842 (N_14842,N_13678,N_13878);
nand U14843 (N_14843,N_14122,N_14241);
nand U14844 (N_14844,N_13717,N_14008);
nor U14845 (N_14845,N_14057,N_13605);
nor U14846 (N_14846,N_13806,N_14176);
and U14847 (N_14847,N_13659,N_13612);
or U14848 (N_14848,N_14204,N_13775);
nor U14849 (N_14849,N_14388,N_14216);
or U14850 (N_14850,N_13850,N_14028);
or U14851 (N_14851,N_14208,N_14199);
or U14852 (N_14852,N_14136,N_14042);
or U14853 (N_14853,N_14319,N_13922);
nand U14854 (N_14854,N_14067,N_13738);
or U14855 (N_14855,N_14384,N_13631);
or U14856 (N_14856,N_14122,N_14395);
or U14857 (N_14857,N_13763,N_14006);
nand U14858 (N_14858,N_14068,N_13694);
nor U14859 (N_14859,N_14055,N_13809);
xor U14860 (N_14860,N_14234,N_14075);
and U14861 (N_14861,N_13820,N_14365);
and U14862 (N_14862,N_13811,N_13966);
nand U14863 (N_14863,N_13896,N_14279);
nand U14864 (N_14864,N_14226,N_14124);
or U14865 (N_14865,N_14031,N_13955);
or U14866 (N_14866,N_13786,N_14220);
nand U14867 (N_14867,N_14075,N_14052);
xor U14868 (N_14868,N_13745,N_14025);
and U14869 (N_14869,N_13755,N_13820);
xnor U14870 (N_14870,N_14119,N_14095);
and U14871 (N_14871,N_13857,N_13801);
and U14872 (N_14872,N_13990,N_14211);
xor U14873 (N_14873,N_14237,N_14201);
xor U14874 (N_14874,N_13785,N_14255);
xor U14875 (N_14875,N_13985,N_14149);
xor U14876 (N_14876,N_14336,N_13793);
nor U14877 (N_14877,N_14214,N_13701);
or U14878 (N_14878,N_14394,N_14133);
xnor U14879 (N_14879,N_13938,N_13659);
and U14880 (N_14880,N_14079,N_14225);
nand U14881 (N_14881,N_13849,N_14291);
or U14882 (N_14882,N_13842,N_13605);
nand U14883 (N_14883,N_14052,N_13739);
and U14884 (N_14884,N_13824,N_14283);
and U14885 (N_14885,N_13956,N_14281);
nor U14886 (N_14886,N_14305,N_13962);
or U14887 (N_14887,N_13627,N_14285);
or U14888 (N_14888,N_14155,N_13943);
xor U14889 (N_14889,N_13905,N_14352);
nor U14890 (N_14890,N_13944,N_14117);
xor U14891 (N_14891,N_13967,N_13886);
nand U14892 (N_14892,N_14237,N_14368);
nand U14893 (N_14893,N_13861,N_14085);
or U14894 (N_14894,N_14136,N_14399);
nor U14895 (N_14895,N_13774,N_13863);
or U14896 (N_14896,N_13892,N_13641);
nand U14897 (N_14897,N_14161,N_14284);
xnor U14898 (N_14898,N_14361,N_13627);
or U14899 (N_14899,N_13687,N_13872);
xor U14900 (N_14900,N_13762,N_14256);
and U14901 (N_14901,N_14218,N_13889);
nand U14902 (N_14902,N_14026,N_14024);
nand U14903 (N_14903,N_13812,N_13607);
and U14904 (N_14904,N_14091,N_14197);
and U14905 (N_14905,N_13681,N_13631);
or U14906 (N_14906,N_14065,N_14112);
and U14907 (N_14907,N_13730,N_13665);
or U14908 (N_14908,N_13760,N_13664);
xor U14909 (N_14909,N_13887,N_14049);
xor U14910 (N_14910,N_13777,N_14241);
nand U14911 (N_14911,N_14391,N_14032);
xor U14912 (N_14912,N_14336,N_14140);
xnor U14913 (N_14913,N_14259,N_13673);
or U14914 (N_14914,N_14065,N_14052);
or U14915 (N_14915,N_14146,N_13778);
nand U14916 (N_14916,N_13923,N_14262);
or U14917 (N_14917,N_14157,N_13819);
nand U14918 (N_14918,N_13847,N_13711);
or U14919 (N_14919,N_14304,N_13744);
nor U14920 (N_14920,N_13814,N_13675);
nand U14921 (N_14921,N_13958,N_14221);
xor U14922 (N_14922,N_13810,N_13692);
nand U14923 (N_14923,N_14176,N_14314);
nand U14924 (N_14924,N_13782,N_14386);
and U14925 (N_14925,N_14237,N_13784);
xnor U14926 (N_14926,N_14313,N_14181);
and U14927 (N_14927,N_13933,N_14346);
nand U14928 (N_14928,N_13760,N_14186);
nand U14929 (N_14929,N_14173,N_13797);
and U14930 (N_14930,N_13699,N_13957);
nor U14931 (N_14931,N_14336,N_14382);
xnor U14932 (N_14932,N_13880,N_13863);
and U14933 (N_14933,N_13660,N_14382);
nand U14934 (N_14934,N_13820,N_13876);
or U14935 (N_14935,N_13938,N_13668);
xor U14936 (N_14936,N_13781,N_13765);
xor U14937 (N_14937,N_13600,N_14170);
and U14938 (N_14938,N_13704,N_13742);
nor U14939 (N_14939,N_14001,N_13626);
or U14940 (N_14940,N_13846,N_13907);
and U14941 (N_14941,N_13693,N_14293);
xnor U14942 (N_14942,N_14076,N_13718);
nand U14943 (N_14943,N_13772,N_14092);
xor U14944 (N_14944,N_13876,N_13661);
and U14945 (N_14945,N_14348,N_14132);
xor U14946 (N_14946,N_14070,N_13923);
and U14947 (N_14947,N_13905,N_14348);
nor U14948 (N_14948,N_13604,N_14160);
nor U14949 (N_14949,N_14006,N_13734);
or U14950 (N_14950,N_13889,N_14385);
or U14951 (N_14951,N_14024,N_14147);
and U14952 (N_14952,N_14307,N_14096);
and U14953 (N_14953,N_13922,N_13825);
xor U14954 (N_14954,N_13739,N_13835);
nand U14955 (N_14955,N_13794,N_14129);
nor U14956 (N_14956,N_14169,N_14250);
xor U14957 (N_14957,N_14098,N_14326);
and U14958 (N_14958,N_13623,N_13809);
nand U14959 (N_14959,N_13831,N_13747);
nand U14960 (N_14960,N_13953,N_14121);
and U14961 (N_14961,N_13738,N_14091);
and U14962 (N_14962,N_13866,N_13700);
or U14963 (N_14963,N_13791,N_14273);
and U14964 (N_14964,N_13793,N_13651);
or U14965 (N_14965,N_13997,N_14125);
xnor U14966 (N_14966,N_14291,N_14180);
and U14967 (N_14967,N_14027,N_14249);
and U14968 (N_14968,N_13925,N_14075);
or U14969 (N_14969,N_14163,N_14087);
or U14970 (N_14970,N_13744,N_13774);
and U14971 (N_14971,N_13710,N_13995);
xor U14972 (N_14972,N_13616,N_14262);
and U14973 (N_14973,N_13632,N_14208);
and U14974 (N_14974,N_13695,N_13947);
nand U14975 (N_14975,N_14383,N_13604);
nor U14976 (N_14976,N_14307,N_14172);
nor U14977 (N_14977,N_14064,N_13610);
and U14978 (N_14978,N_14347,N_13931);
nor U14979 (N_14979,N_13890,N_14275);
and U14980 (N_14980,N_14231,N_14297);
and U14981 (N_14981,N_14262,N_13749);
and U14982 (N_14982,N_13984,N_13660);
nand U14983 (N_14983,N_14307,N_14252);
or U14984 (N_14984,N_13641,N_13965);
nor U14985 (N_14985,N_14080,N_13920);
nor U14986 (N_14986,N_13861,N_13996);
and U14987 (N_14987,N_14367,N_13681);
nand U14988 (N_14988,N_13701,N_13865);
or U14989 (N_14989,N_14094,N_14053);
xor U14990 (N_14990,N_14337,N_14292);
nand U14991 (N_14991,N_14343,N_13796);
nor U14992 (N_14992,N_13675,N_13621);
and U14993 (N_14993,N_14338,N_13985);
nor U14994 (N_14994,N_13809,N_13982);
and U14995 (N_14995,N_13676,N_13635);
and U14996 (N_14996,N_13809,N_13976);
and U14997 (N_14997,N_14168,N_13854);
and U14998 (N_14998,N_13882,N_14294);
xnor U14999 (N_14999,N_13680,N_13959);
or U15000 (N_15000,N_13703,N_14012);
or U15001 (N_15001,N_13751,N_14071);
xnor U15002 (N_15002,N_14392,N_13666);
nand U15003 (N_15003,N_13844,N_14065);
or U15004 (N_15004,N_14254,N_13892);
xnor U15005 (N_15005,N_13814,N_13689);
xnor U15006 (N_15006,N_13923,N_13953);
nor U15007 (N_15007,N_14052,N_13833);
nand U15008 (N_15008,N_14157,N_13893);
xor U15009 (N_15009,N_14046,N_14277);
and U15010 (N_15010,N_14087,N_13801);
or U15011 (N_15011,N_14067,N_14265);
nor U15012 (N_15012,N_14024,N_14185);
or U15013 (N_15013,N_13915,N_13844);
nor U15014 (N_15014,N_13933,N_14186);
and U15015 (N_15015,N_14398,N_14313);
or U15016 (N_15016,N_14084,N_14260);
nand U15017 (N_15017,N_14219,N_13792);
xor U15018 (N_15018,N_14077,N_13608);
and U15019 (N_15019,N_13978,N_13919);
and U15020 (N_15020,N_14088,N_13653);
and U15021 (N_15021,N_14277,N_14049);
nand U15022 (N_15022,N_13677,N_14392);
nor U15023 (N_15023,N_14258,N_13763);
and U15024 (N_15024,N_13837,N_13870);
and U15025 (N_15025,N_14233,N_13603);
nor U15026 (N_15026,N_14349,N_14196);
and U15027 (N_15027,N_13977,N_14020);
nand U15028 (N_15028,N_13806,N_13872);
nor U15029 (N_15029,N_13929,N_13865);
nand U15030 (N_15030,N_14396,N_14037);
nand U15031 (N_15031,N_14177,N_14368);
xnor U15032 (N_15032,N_14304,N_14390);
xnor U15033 (N_15033,N_13637,N_13880);
nand U15034 (N_15034,N_14085,N_14125);
xnor U15035 (N_15035,N_14083,N_13890);
or U15036 (N_15036,N_13653,N_14010);
or U15037 (N_15037,N_14205,N_13667);
and U15038 (N_15038,N_14216,N_13778);
or U15039 (N_15039,N_14273,N_14303);
nor U15040 (N_15040,N_14160,N_14127);
nand U15041 (N_15041,N_14140,N_13985);
xor U15042 (N_15042,N_14306,N_14297);
nand U15043 (N_15043,N_13834,N_13861);
nor U15044 (N_15044,N_13627,N_14096);
and U15045 (N_15045,N_13659,N_14354);
nor U15046 (N_15046,N_14114,N_14003);
or U15047 (N_15047,N_14176,N_13609);
or U15048 (N_15048,N_13828,N_13709);
and U15049 (N_15049,N_13798,N_13662);
nand U15050 (N_15050,N_14142,N_13926);
or U15051 (N_15051,N_14193,N_14092);
and U15052 (N_15052,N_14343,N_14133);
xnor U15053 (N_15053,N_14008,N_13918);
nor U15054 (N_15054,N_13893,N_13752);
nor U15055 (N_15055,N_14318,N_13800);
nor U15056 (N_15056,N_14221,N_14381);
and U15057 (N_15057,N_14268,N_14315);
and U15058 (N_15058,N_14389,N_14207);
or U15059 (N_15059,N_13915,N_13708);
xnor U15060 (N_15060,N_14023,N_14084);
xor U15061 (N_15061,N_13702,N_14277);
xnor U15062 (N_15062,N_13917,N_14010);
or U15063 (N_15063,N_13829,N_13661);
and U15064 (N_15064,N_14327,N_13772);
or U15065 (N_15065,N_14193,N_13821);
or U15066 (N_15066,N_13841,N_14046);
nand U15067 (N_15067,N_14233,N_14105);
nor U15068 (N_15068,N_14195,N_13984);
nand U15069 (N_15069,N_13821,N_13966);
xor U15070 (N_15070,N_13725,N_13930);
or U15071 (N_15071,N_13829,N_14342);
and U15072 (N_15072,N_14209,N_14395);
xnor U15073 (N_15073,N_13960,N_13842);
and U15074 (N_15074,N_13681,N_13625);
xor U15075 (N_15075,N_14331,N_14277);
or U15076 (N_15076,N_13839,N_14001);
and U15077 (N_15077,N_13849,N_14032);
xnor U15078 (N_15078,N_14096,N_13766);
xnor U15079 (N_15079,N_13697,N_14188);
xnor U15080 (N_15080,N_13664,N_13700);
and U15081 (N_15081,N_14184,N_14105);
or U15082 (N_15082,N_14275,N_14051);
nor U15083 (N_15083,N_13605,N_13768);
or U15084 (N_15084,N_13956,N_13702);
nor U15085 (N_15085,N_14188,N_14398);
or U15086 (N_15086,N_14031,N_14303);
or U15087 (N_15087,N_13666,N_13866);
xnor U15088 (N_15088,N_14168,N_14052);
and U15089 (N_15089,N_13946,N_13713);
and U15090 (N_15090,N_13857,N_13752);
or U15091 (N_15091,N_14159,N_13755);
xnor U15092 (N_15092,N_14275,N_14388);
or U15093 (N_15093,N_13961,N_14135);
and U15094 (N_15094,N_14338,N_14231);
and U15095 (N_15095,N_13950,N_14281);
and U15096 (N_15096,N_13889,N_13954);
nand U15097 (N_15097,N_13686,N_14265);
and U15098 (N_15098,N_13943,N_14000);
xnor U15099 (N_15099,N_14385,N_13894);
xor U15100 (N_15100,N_14396,N_13700);
and U15101 (N_15101,N_14343,N_14241);
xnor U15102 (N_15102,N_14385,N_13718);
and U15103 (N_15103,N_14343,N_14186);
nor U15104 (N_15104,N_13869,N_14171);
nor U15105 (N_15105,N_13951,N_13841);
nand U15106 (N_15106,N_14354,N_14001);
and U15107 (N_15107,N_13932,N_14148);
or U15108 (N_15108,N_14038,N_13614);
nor U15109 (N_15109,N_14240,N_13904);
or U15110 (N_15110,N_14123,N_13809);
and U15111 (N_15111,N_13852,N_13608);
nand U15112 (N_15112,N_14206,N_13716);
nand U15113 (N_15113,N_14347,N_13750);
nor U15114 (N_15114,N_14006,N_14029);
or U15115 (N_15115,N_13704,N_13971);
or U15116 (N_15116,N_13706,N_14257);
or U15117 (N_15117,N_14081,N_13780);
or U15118 (N_15118,N_13846,N_13850);
or U15119 (N_15119,N_13744,N_13990);
nand U15120 (N_15120,N_14203,N_14254);
nand U15121 (N_15121,N_13657,N_14376);
or U15122 (N_15122,N_13822,N_13968);
and U15123 (N_15123,N_13877,N_14134);
or U15124 (N_15124,N_13922,N_13636);
and U15125 (N_15125,N_13940,N_14107);
or U15126 (N_15126,N_13725,N_14032);
nor U15127 (N_15127,N_13987,N_14064);
and U15128 (N_15128,N_13601,N_14212);
nor U15129 (N_15129,N_14342,N_14284);
and U15130 (N_15130,N_14046,N_14302);
nor U15131 (N_15131,N_14289,N_14286);
nor U15132 (N_15132,N_13682,N_14005);
xor U15133 (N_15133,N_13861,N_13833);
nand U15134 (N_15134,N_13683,N_14095);
or U15135 (N_15135,N_14236,N_13729);
and U15136 (N_15136,N_13669,N_13892);
nor U15137 (N_15137,N_14021,N_13855);
and U15138 (N_15138,N_13649,N_13639);
or U15139 (N_15139,N_13685,N_14025);
and U15140 (N_15140,N_14110,N_14341);
or U15141 (N_15141,N_13725,N_14082);
or U15142 (N_15142,N_13766,N_14064);
xnor U15143 (N_15143,N_14367,N_13750);
or U15144 (N_15144,N_13768,N_13779);
and U15145 (N_15145,N_14164,N_14321);
xnor U15146 (N_15146,N_13972,N_14190);
or U15147 (N_15147,N_14339,N_14057);
nor U15148 (N_15148,N_14387,N_13749);
nor U15149 (N_15149,N_14038,N_14337);
and U15150 (N_15150,N_14213,N_13766);
nand U15151 (N_15151,N_14091,N_14176);
nor U15152 (N_15152,N_13878,N_14387);
nand U15153 (N_15153,N_14360,N_13920);
and U15154 (N_15154,N_13750,N_13707);
nor U15155 (N_15155,N_13815,N_13623);
and U15156 (N_15156,N_14122,N_14095);
xnor U15157 (N_15157,N_13631,N_14351);
nor U15158 (N_15158,N_13877,N_13863);
nand U15159 (N_15159,N_13965,N_14229);
xor U15160 (N_15160,N_13981,N_13680);
or U15161 (N_15161,N_14390,N_14359);
nor U15162 (N_15162,N_13977,N_14137);
or U15163 (N_15163,N_13888,N_13643);
and U15164 (N_15164,N_13613,N_13942);
xnor U15165 (N_15165,N_13971,N_14327);
nor U15166 (N_15166,N_14154,N_13841);
and U15167 (N_15167,N_14032,N_13745);
nand U15168 (N_15168,N_14273,N_13827);
nand U15169 (N_15169,N_13705,N_14239);
nor U15170 (N_15170,N_14318,N_13653);
nand U15171 (N_15171,N_13681,N_14145);
and U15172 (N_15172,N_14332,N_14169);
nor U15173 (N_15173,N_13825,N_14073);
xnor U15174 (N_15174,N_13739,N_14026);
and U15175 (N_15175,N_14178,N_13997);
nand U15176 (N_15176,N_14116,N_14037);
or U15177 (N_15177,N_14167,N_13763);
nor U15178 (N_15178,N_13661,N_14316);
nand U15179 (N_15179,N_14133,N_14363);
nand U15180 (N_15180,N_14259,N_13683);
nand U15181 (N_15181,N_14225,N_13804);
and U15182 (N_15182,N_13924,N_13931);
and U15183 (N_15183,N_13932,N_14297);
xor U15184 (N_15184,N_14302,N_14300);
or U15185 (N_15185,N_14147,N_13963);
xor U15186 (N_15186,N_13990,N_14032);
nor U15187 (N_15187,N_13984,N_13732);
xnor U15188 (N_15188,N_13750,N_14318);
nor U15189 (N_15189,N_13867,N_13949);
xor U15190 (N_15190,N_13775,N_13736);
nand U15191 (N_15191,N_13750,N_13886);
nand U15192 (N_15192,N_13794,N_13938);
nand U15193 (N_15193,N_13964,N_14218);
or U15194 (N_15194,N_13994,N_14103);
nand U15195 (N_15195,N_13911,N_14365);
or U15196 (N_15196,N_14280,N_14042);
nor U15197 (N_15197,N_14192,N_13941);
or U15198 (N_15198,N_13919,N_14309);
nor U15199 (N_15199,N_14174,N_14231);
or U15200 (N_15200,N_15074,N_14790);
nor U15201 (N_15201,N_14766,N_15105);
nand U15202 (N_15202,N_14673,N_14944);
nor U15203 (N_15203,N_14430,N_14633);
or U15204 (N_15204,N_15188,N_15155);
xnor U15205 (N_15205,N_15133,N_15176);
nand U15206 (N_15206,N_14784,N_14590);
or U15207 (N_15207,N_14862,N_14823);
xor U15208 (N_15208,N_14435,N_14840);
and U15209 (N_15209,N_14698,N_14973);
xnor U15210 (N_15210,N_14414,N_14429);
and U15211 (N_15211,N_14499,N_14697);
xor U15212 (N_15212,N_14963,N_14609);
nand U15213 (N_15213,N_14871,N_14566);
nor U15214 (N_15214,N_15031,N_14910);
and U15215 (N_15215,N_15180,N_14824);
xor U15216 (N_15216,N_14653,N_15084);
and U15217 (N_15217,N_14972,N_15017);
and U15218 (N_15218,N_14986,N_14737);
xnor U15219 (N_15219,N_14934,N_14561);
nor U15220 (N_15220,N_14714,N_15128);
nand U15221 (N_15221,N_14700,N_14532);
nand U15222 (N_15222,N_15022,N_14756);
or U15223 (N_15223,N_14870,N_15101);
nand U15224 (N_15224,N_15115,N_14449);
xor U15225 (N_15225,N_14912,N_14486);
nand U15226 (N_15226,N_14549,N_14475);
or U15227 (N_15227,N_14624,N_14646);
xnor U15228 (N_15228,N_14488,N_15051);
or U15229 (N_15229,N_14667,N_15187);
or U15230 (N_15230,N_14854,N_14456);
and U15231 (N_15231,N_14782,N_14672);
nor U15232 (N_15232,N_15171,N_14453);
nand U15233 (N_15233,N_14852,N_14664);
nor U15234 (N_15234,N_14471,N_15011);
nor U15235 (N_15235,N_14876,N_14436);
or U15236 (N_15236,N_14647,N_14858);
or U15237 (N_15237,N_15024,N_14713);
nand U15238 (N_15238,N_14631,N_14718);
and U15239 (N_15239,N_14939,N_14805);
nor U15240 (N_15240,N_14778,N_14675);
and U15241 (N_15241,N_14989,N_15106);
nor U15242 (N_15242,N_14514,N_15119);
or U15243 (N_15243,N_14494,N_14534);
nand U15244 (N_15244,N_14531,N_14458);
and U15245 (N_15245,N_14613,N_14855);
xnor U15246 (N_15246,N_15175,N_14620);
nor U15247 (N_15247,N_14418,N_14689);
nand U15248 (N_15248,N_14744,N_14949);
xnor U15249 (N_15249,N_15123,N_14723);
or U15250 (N_15250,N_15195,N_15072);
or U15251 (N_15251,N_14748,N_14819);
xnor U15252 (N_15252,N_15161,N_14965);
or U15253 (N_15253,N_14985,N_15050);
and U15254 (N_15254,N_14717,N_14878);
nor U15255 (N_15255,N_14943,N_14866);
and U15256 (N_15256,N_14961,N_15083);
nand U15257 (N_15257,N_14657,N_14880);
nand U15258 (N_15258,N_14457,N_14841);
xor U15259 (N_15259,N_14892,N_14842);
and U15260 (N_15260,N_14837,N_14911);
nor U15261 (N_15261,N_14898,N_14780);
nor U15262 (N_15262,N_14928,N_14504);
nand U15263 (N_15263,N_14535,N_15117);
nand U15264 (N_15264,N_15097,N_15118);
and U15265 (N_15265,N_14467,N_14420);
or U15266 (N_15266,N_14865,N_15138);
or U15267 (N_15267,N_14632,N_14760);
nor U15268 (N_15268,N_14616,N_14587);
and U15269 (N_15269,N_14922,N_14881);
nand U15270 (N_15270,N_14753,N_14599);
nor U15271 (N_15271,N_14542,N_14650);
xor U15272 (N_15272,N_14726,N_14627);
nand U15273 (N_15273,N_15058,N_14439);
or U15274 (N_15274,N_14563,N_14997);
or U15275 (N_15275,N_14519,N_14891);
or U15276 (N_15276,N_14994,N_14945);
and U15277 (N_15277,N_15141,N_15149);
or U15278 (N_15278,N_14806,N_14802);
nand U15279 (N_15279,N_15007,N_14606);
nand U15280 (N_15280,N_14799,N_14409);
nand U15281 (N_15281,N_14521,N_14530);
nor U15282 (N_15282,N_14797,N_14834);
nand U15283 (N_15283,N_14551,N_14734);
nand U15284 (N_15284,N_14607,N_15116);
nand U15285 (N_15285,N_14591,N_14412);
nand U15286 (N_15286,N_15035,N_15110);
or U15287 (N_15287,N_15094,N_14578);
xor U15288 (N_15288,N_14815,N_14894);
or U15289 (N_15289,N_14422,N_15067);
and U15290 (N_15290,N_15013,N_14827);
or U15291 (N_15291,N_15069,N_14548);
nand U15292 (N_15292,N_15030,N_15156);
xor U15293 (N_15293,N_14592,N_14702);
nor U15294 (N_15294,N_14612,N_14879);
nand U15295 (N_15295,N_15047,N_14450);
xnor U15296 (N_15296,N_14916,N_14847);
nand U15297 (N_15297,N_14820,N_14861);
and U15298 (N_15298,N_14497,N_14953);
and U15299 (N_15299,N_15194,N_15134);
nand U15300 (N_15300,N_14527,N_14400);
or U15301 (N_15301,N_14473,N_14932);
nor U15302 (N_15302,N_15080,N_14401);
and U15303 (N_15303,N_15078,N_14452);
or U15304 (N_15304,N_14623,N_14954);
xor U15305 (N_15305,N_14446,N_14403);
nand U15306 (N_15306,N_14863,N_14528);
nor U15307 (N_15307,N_14860,N_14501);
and U15308 (N_15308,N_14836,N_14728);
nand U15309 (N_15309,N_14517,N_14537);
nor U15310 (N_15310,N_14776,N_14625);
xnor U15311 (N_15311,N_15081,N_15053);
or U15312 (N_15312,N_14921,N_14825);
nand U15313 (N_15313,N_14683,N_14722);
nor U15314 (N_15314,N_14864,N_14908);
and U15315 (N_15315,N_14476,N_15165);
or U15316 (N_15316,N_14597,N_14410);
xor U15317 (N_15317,N_14480,N_14502);
nand U15318 (N_15318,N_14691,N_14424);
xor U15319 (N_15319,N_15198,N_14661);
nor U15320 (N_15320,N_15002,N_14874);
nand U15321 (N_15321,N_14662,N_14843);
nand U15322 (N_15322,N_14937,N_14977);
nand U15323 (N_15323,N_14557,N_14992);
xor U15324 (N_15324,N_15109,N_14987);
and U15325 (N_15325,N_15114,N_14500);
and U15326 (N_15326,N_14765,N_14979);
or U15327 (N_15327,N_14956,N_15189);
xnor U15328 (N_15328,N_15167,N_14838);
xor U15329 (N_15329,N_14955,N_14816);
and U15330 (N_15330,N_15143,N_15100);
nand U15331 (N_15331,N_14626,N_14498);
nor U15332 (N_15332,N_14565,N_14618);
or U15333 (N_15333,N_14506,N_14851);
nand U15334 (N_15334,N_14438,N_15012);
nand U15335 (N_15335,N_14629,N_15038);
nand U15336 (N_15336,N_14853,N_15131);
xnor U15337 (N_15337,N_14707,N_15145);
xnor U15338 (N_15338,N_14421,N_14877);
xnor U15339 (N_15339,N_14508,N_15062);
or U15340 (N_15340,N_14696,N_14669);
nand U15341 (N_15341,N_15193,N_14971);
or U15342 (N_15342,N_15185,N_14919);
nor U15343 (N_15343,N_14596,N_14749);
xnor U15344 (N_15344,N_14895,N_15098);
nand U15345 (N_15345,N_14777,N_14545);
nor U15346 (N_15346,N_14586,N_15163);
xor U15347 (N_15347,N_14523,N_14507);
nand U15348 (N_15348,N_14638,N_14567);
and U15349 (N_15349,N_14513,N_14890);
nor U15350 (N_15350,N_14725,N_14826);
nand U15351 (N_15351,N_14964,N_14583);
and U15352 (N_15352,N_14907,N_15174);
or U15353 (N_15353,N_14594,N_15186);
and U15354 (N_15354,N_15120,N_15019);
xor U15355 (N_15355,N_14572,N_15008);
or U15356 (N_15356,N_14419,N_14693);
xor U15357 (N_15357,N_14741,N_15199);
xor U15358 (N_15358,N_14550,N_14443);
or U15359 (N_15359,N_14644,N_14540);
or U15360 (N_15360,N_14524,N_14670);
nand U15361 (N_15361,N_15124,N_14801);
or U15362 (N_15362,N_15113,N_14974);
or U15363 (N_15363,N_14993,N_14405);
xnor U15364 (N_15364,N_14512,N_14428);
and U15365 (N_15365,N_14788,N_14795);
and U15366 (N_15366,N_14931,N_15173);
nor U15367 (N_15367,N_15041,N_14967);
or U15368 (N_15368,N_14680,N_14995);
nand U15369 (N_15369,N_14455,N_14968);
or U15370 (N_15370,N_14929,N_15040);
nand U15371 (N_15371,N_14743,N_14738);
nor U15372 (N_15372,N_14755,N_14526);
nand U15373 (N_15373,N_15140,N_15162);
xor U15374 (N_15374,N_14639,N_14957);
nor U15375 (N_15375,N_14850,N_14783);
nand U15376 (N_15376,N_14705,N_15056);
or U15377 (N_15377,N_14716,N_15102);
nand U15378 (N_15378,N_14767,N_14999);
nand U15379 (N_15379,N_14990,N_14873);
or U15380 (N_15380,N_15027,N_14712);
nand U15381 (N_15381,N_15028,N_14708);
nand U15382 (N_15382,N_14938,N_14832);
xnor U15383 (N_15383,N_14547,N_14727);
nor U15384 (N_15384,N_14442,N_14630);
or U15385 (N_15385,N_15076,N_14720);
or U15386 (N_15386,N_14897,N_14637);
or U15387 (N_15387,N_15015,N_14759);
nor U15388 (N_15388,N_14692,N_14829);
or U15389 (N_15389,N_14555,N_14688);
xor U15390 (N_15390,N_14773,N_15093);
nor U15391 (N_15391,N_14818,N_14431);
nand U15392 (N_15392,N_14556,N_14411);
nor U15393 (N_15393,N_14466,N_14503);
or U15394 (N_15394,N_14715,N_14694);
or U15395 (N_15395,N_15125,N_14699);
nand U15396 (N_15396,N_14554,N_14918);
xor U15397 (N_15397,N_14984,N_14614);
or U15398 (N_15398,N_15046,N_14786);
and U15399 (N_15399,N_15168,N_14899);
xnor U15400 (N_15400,N_14889,N_14525);
and U15401 (N_15401,N_14859,N_14463);
and U15402 (N_15402,N_14774,N_15079);
xnor U15403 (N_15403,N_14604,N_14615);
nand U15404 (N_15404,N_14883,N_14804);
or U15405 (N_15405,N_15152,N_14413);
and U15406 (N_15406,N_15139,N_14875);
xnor U15407 (N_15407,N_14845,N_14936);
xor U15408 (N_15408,N_14690,N_15026);
and U15409 (N_15409,N_14440,N_14709);
and U15410 (N_15410,N_14792,N_14925);
xor U15411 (N_15411,N_15025,N_14611);
xor U15412 (N_15412,N_14536,N_14747);
or U15413 (N_15413,N_14758,N_14520);
and U15414 (N_15414,N_14654,N_14906);
or U15415 (N_15415,N_14791,N_14679);
and U15416 (N_15416,N_14658,N_14951);
xnor U15417 (N_15417,N_14740,N_14668);
nor U15418 (N_15418,N_14510,N_14573);
or U15419 (N_15419,N_14402,N_14574);
nor U15420 (N_15420,N_14677,N_14745);
nand U15421 (N_15421,N_15068,N_14730);
nor U15422 (N_15422,N_14775,N_14493);
nor U15423 (N_15423,N_15006,N_14509);
and U15424 (N_15424,N_15039,N_14553);
and U15425 (N_15425,N_15052,N_15044);
nor U15426 (N_15426,N_14585,N_14980);
nor U15427 (N_15427,N_15197,N_14946);
xor U15428 (N_15428,N_14433,N_14663);
xnor U15429 (N_15429,N_15042,N_15071);
or U15430 (N_15430,N_14830,N_14762);
nor U15431 (N_15431,N_14605,N_15136);
nor U15432 (N_15432,N_14634,N_14518);
nand U15433 (N_15433,N_15126,N_14404);
and U15434 (N_15434,N_14470,N_14962);
or U15435 (N_15435,N_15048,N_14975);
xor U15436 (N_15436,N_14719,N_15196);
nand U15437 (N_15437,N_14481,N_14900);
xor U15438 (N_15438,N_14541,N_14746);
nor U15439 (N_15439,N_14940,N_14947);
xnor U15440 (N_15440,N_14408,N_15132);
or U15441 (N_15441,N_15032,N_15054);
nand U15442 (N_15442,N_15147,N_14849);
and U15443 (N_15443,N_15169,N_15104);
and U15444 (N_15444,N_15073,N_14868);
xor U15445 (N_15445,N_14909,N_14831);
xor U15446 (N_15446,N_14687,N_14942);
and U15447 (N_15447,N_15066,N_14621);
nor U15448 (N_15448,N_14489,N_14460);
xnor U15449 (N_15449,N_14423,N_14491);
and U15450 (N_15450,N_14477,N_14988);
or U15451 (N_15451,N_14484,N_14655);
nor U15452 (N_15452,N_14576,N_15137);
and U15453 (N_15453,N_15033,N_14562);
and U15454 (N_15454,N_14407,N_15184);
nand U15455 (N_15455,N_14787,N_14848);
nor U15456 (N_15456,N_14811,N_15112);
nand U15457 (N_15457,N_14926,N_14678);
xor U15458 (N_15458,N_14681,N_14495);
nor U15459 (N_15459,N_14462,N_14686);
and U15460 (N_15460,N_14917,N_14872);
or U15461 (N_15461,N_14915,N_14930);
nor U15462 (N_15462,N_14768,N_14807);
xor U15463 (N_15463,N_14996,N_14406);
xnor U15464 (N_15464,N_14803,N_15060);
nand U15465 (N_15465,N_14608,N_14969);
and U15466 (N_15466,N_14483,N_14652);
nor U15467 (N_15467,N_14437,N_14821);
xnor U15468 (N_15468,N_14529,N_15090);
nor U15469 (N_15469,N_14468,N_14432);
xor U15470 (N_15470,N_14622,N_14533);
xnor U15471 (N_15471,N_15000,N_15055);
nand U15472 (N_15472,N_15004,N_14464);
nor U15473 (N_15473,N_15099,N_14735);
or U15474 (N_15474,N_14459,N_14781);
and U15475 (N_15475,N_14703,N_14933);
nand U15476 (N_15476,N_14731,N_15077);
and U15477 (N_15477,N_14581,N_14426);
nor U15478 (N_15478,N_14595,N_14704);
and U15479 (N_15479,N_14732,N_14601);
nand U15480 (N_15480,N_14580,N_14685);
xor U15481 (N_15481,N_14676,N_14885);
or U15482 (N_15482,N_14659,N_15057);
and U15483 (N_15483,N_15121,N_14682);
xor U15484 (N_15484,N_14465,N_14569);
nand U15485 (N_15485,N_14543,N_14461);
nand U15486 (N_15486,N_14635,N_14656);
xnor U15487 (N_15487,N_15144,N_14568);
or U15488 (N_15488,N_14822,N_14695);
xor U15489 (N_15489,N_14779,N_14757);
nand U15490 (N_15490,N_14770,N_14976);
xnor U15491 (N_15491,N_15160,N_14794);
nor U15492 (N_15492,N_15170,N_14813);
and U15493 (N_15493,N_14846,N_14610);
xor U15494 (N_15494,N_14482,N_14427);
or U15495 (N_15495,N_15146,N_14754);
xnor U15496 (N_15496,N_14588,N_15127);
xor U15497 (N_15497,N_14600,N_15037);
nor U15498 (N_15498,N_15034,N_14924);
and U15499 (N_15499,N_14538,N_14516);
xnor U15500 (N_15500,N_14970,N_14771);
nor U15501 (N_15501,N_14844,N_14649);
or U15502 (N_15502,N_14812,N_15122);
and U15503 (N_15503,N_14935,N_15153);
nor U15504 (N_15504,N_14570,N_14867);
or U15505 (N_15505,N_15111,N_15005);
nor U15506 (N_15506,N_14671,N_15045);
nor U15507 (N_15507,N_15183,N_15023);
or U15508 (N_15508,N_14721,N_15089);
and U15509 (N_15509,N_14884,N_15003);
or U15510 (N_15510,N_14701,N_14560);
and U15511 (N_15511,N_14558,N_14736);
or U15512 (N_15512,N_15075,N_14983);
xor U15513 (N_15513,N_14739,N_14642);
nand U15514 (N_15514,N_14978,N_15158);
nor U15515 (N_15515,N_14641,N_15190);
or U15516 (N_15516,N_15029,N_15096);
or U15517 (N_15517,N_14643,N_14950);
or U15518 (N_15518,N_15157,N_14522);
or U15519 (N_15519,N_14598,N_15061);
or U15520 (N_15520,N_14575,N_14835);
nor U15521 (N_15521,N_14948,N_14793);
xor U15522 (N_15522,N_15065,N_14733);
or U15523 (N_15523,N_15063,N_14958);
xnor U15524 (N_15524,N_14941,N_15091);
and U15525 (N_15525,N_15159,N_14544);
xnor U15526 (N_15526,N_14651,N_15172);
or U15527 (N_15527,N_15150,N_15130);
nor U15528 (N_15528,N_14577,N_14991);
and U15529 (N_15529,N_15010,N_14415);
or U15530 (N_15530,N_14952,N_14619);
or U15531 (N_15531,N_15181,N_14905);
and U15532 (N_15532,N_14539,N_14817);
nand U15533 (N_15533,N_15021,N_14810);
xnor U15534 (N_15534,N_15179,N_14579);
nand U15535 (N_15535,N_14665,N_14472);
xor U15536 (N_15536,N_15151,N_14416);
nor U15537 (N_15537,N_14584,N_14490);
and U15538 (N_15538,N_15166,N_14869);
xor U15539 (N_15539,N_14886,N_14814);
and U15540 (N_15540,N_15135,N_15191);
nor U15541 (N_15541,N_14920,N_14496);
or U15542 (N_15542,N_15092,N_14856);
nor U15543 (N_15543,N_14571,N_14769);
or U15544 (N_15544,N_14602,N_14640);
or U15545 (N_15545,N_14434,N_14636);
xnor U15546 (N_15546,N_14603,N_14454);
or U15547 (N_15547,N_14645,N_14750);
nor U15548 (N_15548,N_14448,N_14559);
and U15549 (N_15549,N_15129,N_15095);
and U15550 (N_15550,N_14896,N_14444);
nand U15551 (N_15551,N_14828,N_15177);
and U15552 (N_15552,N_14959,N_14998);
nand U15553 (N_15553,N_15009,N_15178);
nor U15554 (N_15554,N_14789,N_15049);
and U15555 (N_15555,N_14742,N_14711);
nand U15556 (N_15556,N_14882,N_14888);
xor U15557 (N_15557,N_15192,N_15164);
or U15558 (N_15558,N_14960,N_14751);
or U15559 (N_15559,N_14674,N_14887);
nor U15560 (N_15560,N_14469,N_14425);
and U15561 (N_15561,N_15103,N_14684);
xnor U15562 (N_15562,N_15020,N_15088);
or U15563 (N_15563,N_15107,N_14966);
nand U15564 (N_15564,N_14706,N_14893);
nor U15565 (N_15565,N_14752,N_14981);
and U15566 (N_15566,N_15016,N_15085);
nor U15567 (N_15567,N_14511,N_14487);
nor U15568 (N_15568,N_15182,N_14808);
or U15569 (N_15569,N_14515,N_14914);
nor U15570 (N_15570,N_14724,N_14589);
nand U15571 (N_15571,N_14729,N_14796);
nor U15572 (N_15572,N_14648,N_14761);
nor U15573 (N_15573,N_15108,N_15059);
nor U15574 (N_15574,N_14441,N_15014);
and U15575 (N_15575,N_14764,N_15087);
or U15576 (N_15576,N_14903,N_14617);
nand U15577 (N_15577,N_14628,N_14800);
and U15578 (N_15578,N_14902,N_14492);
and U15579 (N_15579,N_14666,N_14546);
and U15580 (N_15580,N_14923,N_14927);
and U15581 (N_15581,N_14478,N_14479);
xnor U15582 (N_15582,N_14593,N_14564);
nor U15583 (N_15583,N_15064,N_14474);
xor U15584 (N_15584,N_14445,N_14857);
and U15585 (N_15585,N_15001,N_14833);
or U15586 (N_15586,N_15142,N_15148);
or U15587 (N_15587,N_15043,N_14710);
nand U15588 (N_15588,N_14913,N_14582);
nand U15589 (N_15589,N_14447,N_15018);
or U15590 (N_15590,N_14798,N_14839);
nor U15591 (N_15591,N_14901,N_15070);
nor U15592 (N_15592,N_14772,N_14809);
xnor U15593 (N_15593,N_14505,N_14660);
and U15594 (N_15594,N_14904,N_14485);
nor U15595 (N_15595,N_15086,N_14785);
and U15596 (N_15596,N_15082,N_14552);
and U15597 (N_15597,N_14982,N_14417);
nand U15598 (N_15598,N_15036,N_15154);
and U15599 (N_15599,N_14451,N_14763);
nor U15600 (N_15600,N_14941,N_14663);
nand U15601 (N_15601,N_14656,N_15003);
or U15602 (N_15602,N_14419,N_14513);
nand U15603 (N_15603,N_14978,N_14785);
nor U15604 (N_15604,N_15057,N_15142);
or U15605 (N_15605,N_14888,N_14581);
nand U15606 (N_15606,N_14937,N_15173);
xor U15607 (N_15607,N_14577,N_14773);
nor U15608 (N_15608,N_15071,N_14994);
nor U15609 (N_15609,N_14401,N_14933);
nand U15610 (N_15610,N_14593,N_14567);
and U15611 (N_15611,N_14667,N_15065);
and U15612 (N_15612,N_14501,N_14761);
and U15613 (N_15613,N_15130,N_15189);
and U15614 (N_15614,N_14605,N_14579);
xnor U15615 (N_15615,N_14968,N_14456);
nand U15616 (N_15616,N_14558,N_15083);
and U15617 (N_15617,N_14964,N_14928);
nor U15618 (N_15618,N_14979,N_14966);
and U15619 (N_15619,N_14934,N_14489);
nand U15620 (N_15620,N_14556,N_14462);
or U15621 (N_15621,N_15040,N_14786);
or U15622 (N_15622,N_14662,N_15182);
nor U15623 (N_15623,N_14601,N_14574);
nor U15624 (N_15624,N_14707,N_14552);
nor U15625 (N_15625,N_14533,N_15149);
or U15626 (N_15626,N_14788,N_14769);
xnor U15627 (N_15627,N_14825,N_14981);
xnor U15628 (N_15628,N_14647,N_14987);
and U15629 (N_15629,N_14845,N_14673);
nor U15630 (N_15630,N_15057,N_14721);
nor U15631 (N_15631,N_14411,N_15136);
xor U15632 (N_15632,N_14554,N_14917);
or U15633 (N_15633,N_15030,N_15037);
and U15634 (N_15634,N_14785,N_14922);
or U15635 (N_15635,N_15091,N_14670);
nor U15636 (N_15636,N_14705,N_14636);
and U15637 (N_15637,N_14558,N_14469);
and U15638 (N_15638,N_14449,N_14739);
or U15639 (N_15639,N_14521,N_15153);
xnor U15640 (N_15640,N_15113,N_15050);
nand U15641 (N_15641,N_14551,N_15174);
nor U15642 (N_15642,N_14480,N_15130);
or U15643 (N_15643,N_15184,N_14528);
or U15644 (N_15644,N_14895,N_14752);
or U15645 (N_15645,N_14779,N_15166);
xor U15646 (N_15646,N_14477,N_15129);
nand U15647 (N_15647,N_14831,N_14870);
xnor U15648 (N_15648,N_14801,N_14802);
nor U15649 (N_15649,N_14694,N_14792);
or U15650 (N_15650,N_15099,N_15032);
and U15651 (N_15651,N_14779,N_14506);
nand U15652 (N_15652,N_14480,N_14694);
nand U15653 (N_15653,N_14585,N_15110);
nand U15654 (N_15654,N_15150,N_14528);
nor U15655 (N_15655,N_15022,N_14532);
nor U15656 (N_15656,N_15085,N_14711);
or U15657 (N_15657,N_15181,N_14919);
nand U15658 (N_15658,N_14870,N_14903);
nor U15659 (N_15659,N_14794,N_14630);
xnor U15660 (N_15660,N_15079,N_14933);
nand U15661 (N_15661,N_14967,N_15049);
xor U15662 (N_15662,N_14715,N_15148);
or U15663 (N_15663,N_14428,N_14835);
nand U15664 (N_15664,N_14549,N_14940);
xor U15665 (N_15665,N_15020,N_14652);
or U15666 (N_15666,N_14845,N_14492);
or U15667 (N_15667,N_14803,N_14958);
or U15668 (N_15668,N_14811,N_14919);
nor U15669 (N_15669,N_14415,N_14875);
and U15670 (N_15670,N_14968,N_14910);
nor U15671 (N_15671,N_14746,N_15034);
nand U15672 (N_15672,N_14691,N_14870);
and U15673 (N_15673,N_14946,N_14741);
nor U15674 (N_15674,N_14819,N_14533);
and U15675 (N_15675,N_14787,N_15034);
or U15676 (N_15676,N_14489,N_14920);
nand U15677 (N_15677,N_15007,N_14642);
nand U15678 (N_15678,N_14708,N_14949);
xor U15679 (N_15679,N_14409,N_14790);
nor U15680 (N_15680,N_15051,N_14655);
and U15681 (N_15681,N_14430,N_14962);
and U15682 (N_15682,N_14793,N_14850);
or U15683 (N_15683,N_14748,N_14635);
nor U15684 (N_15684,N_14859,N_14691);
nand U15685 (N_15685,N_14649,N_14568);
xor U15686 (N_15686,N_15171,N_14524);
nand U15687 (N_15687,N_15102,N_14498);
nand U15688 (N_15688,N_14732,N_15117);
nand U15689 (N_15689,N_14832,N_14663);
nand U15690 (N_15690,N_14774,N_14734);
and U15691 (N_15691,N_14822,N_14923);
xor U15692 (N_15692,N_15192,N_14700);
nor U15693 (N_15693,N_14712,N_14643);
nor U15694 (N_15694,N_15060,N_15005);
nand U15695 (N_15695,N_14702,N_15101);
and U15696 (N_15696,N_15140,N_14609);
and U15697 (N_15697,N_14560,N_14613);
and U15698 (N_15698,N_15170,N_14936);
or U15699 (N_15699,N_14545,N_14679);
and U15700 (N_15700,N_14408,N_14954);
nor U15701 (N_15701,N_15094,N_14483);
or U15702 (N_15702,N_15129,N_14411);
and U15703 (N_15703,N_14973,N_15159);
or U15704 (N_15704,N_14731,N_14953);
and U15705 (N_15705,N_14708,N_14480);
and U15706 (N_15706,N_15158,N_15170);
nand U15707 (N_15707,N_14764,N_14903);
nor U15708 (N_15708,N_14686,N_14443);
nor U15709 (N_15709,N_14452,N_14460);
nor U15710 (N_15710,N_14843,N_14841);
nor U15711 (N_15711,N_14756,N_15184);
xnor U15712 (N_15712,N_14702,N_14729);
xnor U15713 (N_15713,N_14613,N_14726);
xnor U15714 (N_15714,N_14539,N_14730);
nand U15715 (N_15715,N_14825,N_14826);
xnor U15716 (N_15716,N_14401,N_15105);
xnor U15717 (N_15717,N_15007,N_14788);
nor U15718 (N_15718,N_14761,N_14758);
nor U15719 (N_15719,N_14701,N_14946);
xor U15720 (N_15720,N_14548,N_14790);
or U15721 (N_15721,N_14470,N_14404);
nor U15722 (N_15722,N_15134,N_14459);
or U15723 (N_15723,N_14971,N_15035);
or U15724 (N_15724,N_15180,N_14401);
nor U15725 (N_15725,N_14528,N_14799);
and U15726 (N_15726,N_14692,N_14446);
nand U15727 (N_15727,N_14803,N_14480);
nand U15728 (N_15728,N_15170,N_14948);
nor U15729 (N_15729,N_14567,N_14877);
nor U15730 (N_15730,N_14532,N_14983);
xnor U15731 (N_15731,N_14972,N_14933);
xor U15732 (N_15732,N_14642,N_14989);
nor U15733 (N_15733,N_15043,N_14721);
nand U15734 (N_15734,N_14473,N_14712);
and U15735 (N_15735,N_14462,N_14404);
and U15736 (N_15736,N_14829,N_14475);
xor U15737 (N_15737,N_14578,N_15165);
and U15738 (N_15738,N_14575,N_14735);
or U15739 (N_15739,N_15187,N_14594);
nor U15740 (N_15740,N_14620,N_14812);
and U15741 (N_15741,N_15027,N_14717);
nor U15742 (N_15742,N_15195,N_14779);
or U15743 (N_15743,N_14782,N_14560);
xor U15744 (N_15744,N_14612,N_14883);
or U15745 (N_15745,N_14400,N_15015);
nor U15746 (N_15746,N_14404,N_14422);
nor U15747 (N_15747,N_14747,N_15098);
xnor U15748 (N_15748,N_14869,N_14906);
nand U15749 (N_15749,N_14769,N_14831);
nand U15750 (N_15750,N_15000,N_14788);
nand U15751 (N_15751,N_15099,N_14934);
and U15752 (N_15752,N_15032,N_14913);
nor U15753 (N_15753,N_14408,N_14791);
nor U15754 (N_15754,N_14553,N_14668);
and U15755 (N_15755,N_15183,N_15182);
and U15756 (N_15756,N_14577,N_14451);
or U15757 (N_15757,N_14955,N_14562);
nand U15758 (N_15758,N_14516,N_14984);
or U15759 (N_15759,N_15124,N_15008);
nand U15760 (N_15760,N_14586,N_15181);
and U15761 (N_15761,N_14942,N_15055);
nor U15762 (N_15762,N_15012,N_14682);
or U15763 (N_15763,N_14765,N_14892);
xnor U15764 (N_15764,N_14959,N_15056);
nand U15765 (N_15765,N_14909,N_14624);
and U15766 (N_15766,N_15037,N_14899);
or U15767 (N_15767,N_15089,N_14649);
xnor U15768 (N_15768,N_14445,N_14841);
or U15769 (N_15769,N_14739,N_14580);
nand U15770 (N_15770,N_14420,N_14459);
nor U15771 (N_15771,N_14672,N_14705);
and U15772 (N_15772,N_14485,N_14710);
and U15773 (N_15773,N_14850,N_14604);
nor U15774 (N_15774,N_14772,N_14757);
or U15775 (N_15775,N_14784,N_14695);
or U15776 (N_15776,N_14891,N_15100);
nand U15777 (N_15777,N_14604,N_15060);
xor U15778 (N_15778,N_14603,N_14613);
xnor U15779 (N_15779,N_15012,N_15029);
xor U15780 (N_15780,N_14971,N_15144);
and U15781 (N_15781,N_15053,N_15159);
and U15782 (N_15782,N_14673,N_14844);
or U15783 (N_15783,N_14602,N_14966);
or U15784 (N_15784,N_14728,N_14409);
or U15785 (N_15785,N_15038,N_14575);
nand U15786 (N_15786,N_15003,N_14998);
or U15787 (N_15787,N_14755,N_14437);
and U15788 (N_15788,N_14518,N_14652);
nand U15789 (N_15789,N_14654,N_14676);
nor U15790 (N_15790,N_14705,N_14597);
and U15791 (N_15791,N_15080,N_14736);
nand U15792 (N_15792,N_14552,N_15161);
nor U15793 (N_15793,N_14525,N_14821);
and U15794 (N_15794,N_14729,N_14554);
nor U15795 (N_15795,N_14643,N_15083);
nand U15796 (N_15796,N_14519,N_14732);
nand U15797 (N_15797,N_14571,N_14492);
xor U15798 (N_15798,N_14524,N_14617);
and U15799 (N_15799,N_14912,N_14696);
nand U15800 (N_15800,N_15113,N_14988);
xor U15801 (N_15801,N_15162,N_14862);
nand U15802 (N_15802,N_14690,N_14674);
nand U15803 (N_15803,N_14508,N_14428);
nand U15804 (N_15804,N_15049,N_14555);
xnor U15805 (N_15805,N_14673,N_14972);
or U15806 (N_15806,N_15149,N_14929);
nor U15807 (N_15807,N_14530,N_15143);
or U15808 (N_15808,N_14852,N_14597);
and U15809 (N_15809,N_14601,N_14914);
and U15810 (N_15810,N_15037,N_15064);
xnor U15811 (N_15811,N_14626,N_14795);
nor U15812 (N_15812,N_15047,N_14500);
or U15813 (N_15813,N_14517,N_14839);
nor U15814 (N_15814,N_14634,N_14475);
xor U15815 (N_15815,N_15059,N_14605);
or U15816 (N_15816,N_14898,N_14668);
nand U15817 (N_15817,N_15065,N_14885);
nor U15818 (N_15818,N_14876,N_14898);
xnor U15819 (N_15819,N_14681,N_14421);
or U15820 (N_15820,N_14852,N_14776);
or U15821 (N_15821,N_14549,N_14416);
or U15822 (N_15822,N_14443,N_14953);
and U15823 (N_15823,N_15192,N_14564);
and U15824 (N_15824,N_14431,N_15159);
and U15825 (N_15825,N_15057,N_14540);
xnor U15826 (N_15826,N_14441,N_14645);
nor U15827 (N_15827,N_15160,N_15055);
nor U15828 (N_15828,N_14734,N_14548);
nor U15829 (N_15829,N_14979,N_14922);
xnor U15830 (N_15830,N_14809,N_14544);
nor U15831 (N_15831,N_14795,N_15188);
and U15832 (N_15832,N_14928,N_14925);
nand U15833 (N_15833,N_15085,N_15174);
or U15834 (N_15834,N_14843,N_14795);
xor U15835 (N_15835,N_14781,N_14544);
nand U15836 (N_15836,N_15014,N_14648);
nand U15837 (N_15837,N_14534,N_14863);
or U15838 (N_15838,N_14607,N_14799);
or U15839 (N_15839,N_14737,N_14718);
xnor U15840 (N_15840,N_14549,N_14508);
xor U15841 (N_15841,N_15057,N_14819);
nor U15842 (N_15842,N_14815,N_14892);
and U15843 (N_15843,N_14656,N_14564);
nor U15844 (N_15844,N_14627,N_14850);
nand U15845 (N_15845,N_14781,N_15123);
nand U15846 (N_15846,N_14857,N_14513);
or U15847 (N_15847,N_14490,N_15146);
or U15848 (N_15848,N_14492,N_15087);
nor U15849 (N_15849,N_14533,N_14722);
xor U15850 (N_15850,N_15188,N_14854);
nand U15851 (N_15851,N_15114,N_14578);
nor U15852 (N_15852,N_14604,N_14521);
nand U15853 (N_15853,N_14870,N_14702);
xor U15854 (N_15854,N_15121,N_14976);
or U15855 (N_15855,N_14451,N_14503);
nand U15856 (N_15856,N_14730,N_15139);
xor U15857 (N_15857,N_14674,N_14854);
and U15858 (N_15858,N_14905,N_14705);
nand U15859 (N_15859,N_15174,N_15071);
nor U15860 (N_15860,N_15008,N_14809);
xnor U15861 (N_15861,N_14930,N_14693);
nor U15862 (N_15862,N_14993,N_15148);
and U15863 (N_15863,N_14833,N_14650);
nand U15864 (N_15864,N_14616,N_14644);
nand U15865 (N_15865,N_14507,N_14945);
nand U15866 (N_15866,N_14642,N_14552);
and U15867 (N_15867,N_15089,N_14692);
nand U15868 (N_15868,N_15033,N_14962);
and U15869 (N_15869,N_14499,N_14959);
and U15870 (N_15870,N_14732,N_14455);
nand U15871 (N_15871,N_14662,N_14721);
nand U15872 (N_15872,N_14735,N_14876);
xnor U15873 (N_15873,N_14832,N_14599);
xnor U15874 (N_15874,N_14965,N_15121);
and U15875 (N_15875,N_14928,N_15153);
and U15876 (N_15876,N_14462,N_14875);
xor U15877 (N_15877,N_14443,N_14658);
xnor U15878 (N_15878,N_14973,N_14428);
or U15879 (N_15879,N_14687,N_14971);
nand U15880 (N_15880,N_14403,N_14994);
and U15881 (N_15881,N_15068,N_14713);
nor U15882 (N_15882,N_14401,N_15183);
and U15883 (N_15883,N_14492,N_14708);
nor U15884 (N_15884,N_14996,N_14731);
nor U15885 (N_15885,N_15027,N_14674);
and U15886 (N_15886,N_15157,N_14633);
nand U15887 (N_15887,N_14536,N_15062);
nor U15888 (N_15888,N_14729,N_14623);
or U15889 (N_15889,N_14987,N_14531);
or U15890 (N_15890,N_14416,N_14822);
xor U15891 (N_15891,N_15057,N_14989);
or U15892 (N_15892,N_14435,N_14642);
nand U15893 (N_15893,N_14920,N_14873);
nand U15894 (N_15894,N_14488,N_15011);
xnor U15895 (N_15895,N_14949,N_14805);
nand U15896 (N_15896,N_15033,N_14607);
and U15897 (N_15897,N_14669,N_15021);
or U15898 (N_15898,N_14933,N_14874);
nand U15899 (N_15899,N_14884,N_14734);
and U15900 (N_15900,N_14545,N_14561);
nand U15901 (N_15901,N_14921,N_14432);
or U15902 (N_15902,N_14727,N_15043);
or U15903 (N_15903,N_15035,N_14660);
nor U15904 (N_15904,N_14653,N_14579);
nand U15905 (N_15905,N_14488,N_14551);
nand U15906 (N_15906,N_14959,N_14488);
or U15907 (N_15907,N_14790,N_14825);
xor U15908 (N_15908,N_14531,N_14732);
and U15909 (N_15909,N_14513,N_14819);
xnor U15910 (N_15910,N_15005,N_15011);
and U15911 (N_15911,N_14686,N_14403);
nand U15912 (N_15912,N_14993,N_14997);
or U15913 (N_15913,N_14612,N_14437);
and U15914 (N_15914,N_14793,N_14676);
nor U15915 (N_15915,N_14973,N_15177);
nand U15916 (N_15916,N_14582,N_14723);
xnor U15917 (N_15917,N_14730,N_14602);
nand U15918 (N_15918,N_14863,N_15110);
nand U15919 (N_15919,N_14861,N_14842);
nand U15920 (N_15920,N_14599,N_14679);
or U15921 (N_15921,N_14605,N_15171);
and U15922 (N_15922,N_14424,N_15183);
nor U15923 (N_15923,N_14676,N_15004);
or U15924 (N_15924,N_14793,N_14631);
nand U15925 (N_15925,N_15048,N_14955);
nor U15926 (N_15926,N_14871,N_15085);
xor U15927 (N_15927,N_14739,N_15067);
nand U15928 (N_15928,N_14817,N_14965);
nor U15929 (N_15929,N_15097,N_14471);
and U15930 (N_15930,N_14440,N_14509);
or U15931 (N_15931,N_14752,N_15025);
and U15932 (N_15932,N_14838,N_14950);
or U15933 (N_15933,N_15016,N_14872);
xnor U15934 (N_15934,N_15022,N_14869);
xnor U15935 (N_15935,N_14847,N_14739);
xor U15936 (N_15936,N_14712,N_15104);
nor U15937 (N_15937,N_14444,N_14947);
or U15938 (N_15938,N_14584,N_14481);
xor U15939 (N_15939,N_14498,N_14847);
or U15940 (N_15940,N_14475,N_14590);
xor U15941 (N_15941,N_14475,N_15091);
and U15942 (N_15942,N_14807,N_14754);
nor U15943 (N_15943,N_15155,N_14496);
nand U15944 (N_15944,N_14422,N_15001);
or U15945 (N_15945,N_15023,N_15193);
xnor U15946 (N_15946,N_14751,N_14921);
or U15947 (N_15947,N_14620,N_15197);
nand U15948 (N_15948,N_14980,N_14794);
nand U15949 (N_15949,N_14439,N_14837);
xnor U15950 (N_15950,N_14583,N_14977);
xor U15951 (N_15951,N_14849,N_15013);
nor U15952 (N_15952,N_14532,N_14596);
and U15953 (N_15953,N_14831,N_14506);
and U15954 (N_15954,N_14471,N_14627);
or U15955 (N_15955,N_14947,N_14695);
nor U15956 (N_15956,N_14571,N_14703);
xor U15957 (N_15957,N_15067,N_14496);
nor U15958 (N_15958,N_14453,N_15148);
nor U15959 (N_15959,N_14493,N_14733);
or U15960 (N_15960,N_14545,N_14660);
xnor U15961 (N_15961,N_15132,N_15154);
or U15962 (N_15962,N_14922,N_14987);
and U15963 (N_15963,N_14524,N_14407);
or U15964 (N_15964,N_14761,N_14613);
or U15965 (N_15965,N_14979,N_14888);
and U15966 (N_15966,N_14480,N_15085);
nor U15967 (N_15967,N_14944,N_14686);
or U15968 (N_15968,N_14473,N_15125);
nand U15969 (N_15969,N_14770,N_14751);
nor U15970 (N_15970,N_14662,N_15074);
xnor U15971 (N_15971,N_14452,N_14465);
xnor U15972 (N_15972,N_15066,N_14870);
nand U15973 (N_15973,N_14781,N_14416);
or U15974 (N_15974,N_15198,N_14958);
or U15975 (N_15975,N_14727,N_14573);
nor U15976 (N_15976,N_14850,N_14693);
and U15977 (N_15977,N_14575,N_14467);
nor U15978 (N_15978,N_15168,N_14699);
nor U15979 (N_15979,N_14458,N_14497);
and U15980 (N_15980,N_14964,N_14919);
xor U15981 (N_15981,N_14595,N_14938);
xor U15982 (N_15982,N_14532,N_14914);
xor U15983 (N_15983,N_14839,N_14709);
nand U15984 (N_15984,N_14565,N_14843);
and U15985 (N_15985,N_14630,N_15125);
or U15986 (N_15986,N_15167,N_14907);
xnor U15987 (N_15987,N_14981,N_14602);
and U15988 (N_15988,N_15069,N_14495);
nand U15989 (N_15989,N_14514,N_15060);
and U15990 (N_15990,N_14718,N_14698);
nor U15991 (N_15991,N_14771,N_14621);
and U15992 (N_15992,N_14944,N_14736);
and U15993 (N_15993,N_15114,N_14727);
xnor U15994 (N_15994,N_15173,N_14928);
nand U15995 (N_15995,N_15186,N_14769);
nor U15996 (N_15996,N_15121,N_14951);
nand U15997 (N_15997,N_14594,N_14815);
xor U15998 (N_15998,N_14419,N_15146);
xor U15999 (N_15999,N_14792,N_14478);
or U16000 (N_16000,N_15422,N_15453);
xnor U16001 (N_16001,N_15942,N_15745);
nor U16002 (N_16002,N_15738,N_15236);
nor U16003 (N_16003,N_15979,N_15641);
nor U16004 (N_16004,N_15555,N_15892);
nand U16005 (N_16005,N_15430,N_15448);
nand U16006 (N_16006,N_15438,N_15707);
or U16007 (N_16007,N_15984,N_15746);
and U16008 (N_16008,N_15293,N_15951);
xnor U16009 (N_16009,N_15612,N_15418);
or U16010 (N_16010,N_15954,N_15651);
nand U16011 (N_16011,N_15369,N_15306);
xor U16012 (N_16012,N_15724,N_15322);
xnor U16013 (N_16013,N_15292,N_15590);
nand U16014 (N_16014,N_15442,N_15494);
xnor U16015 (N_16015,N_15374,N_15976);
and U16016 (N_16016,N_15224,N_15456);
xnor U16017 (N_16017,N_15841,N_15221);
or U16018 (N_16018,N_15632,N_15474);
and U16019 (N_16019,N_15385,N_15513);
or U16020 (N_16020,N_15330,N_15643);
and U16021 (N_16021,N_15480,N_15327);
or U16022 (N_16022,N_15940,N_15622);
xnor U16023 (N_16023,N_15941,N_15207);
xnor U16024 (N_16024,N_15649,N_15914);
xor U16025 (N_16025,N_15635,N_15929);
or U16026 (N_16026,N_15899,N_15657);
or U16027 (N_16027,N_15329,N_15961);
and U16028 (N_16028,N_15817,N_15286);
nor U16029 (N_16029,N_15432,N_15508);
nor U16030 (N_16030,N_15556,N_15901);
and U16031 (N_16031,N_15604,N_15405);
and U16032 (N_16032,N_15410,N_15301);
nor U16033 (N_16033,N_15821,N_15365);
xor U16034 (N_16034,N_15787,N_15939);
xor U16035 (N_16035,N_15948,N_15227);
nand U16036 (N_16036,N_15989,N_15790);
xor U16037 (N_16037,N_15563,N_15297);
and U16038 (N_16038,N_15888,N_15294);
xor U16039 (N_16039,N_15858,N_15974);
nor U16040 (N_16040,N_15439,N_15501);
and U16041 (N_16041,N_15658,N_15341);
or U16042 (N_16042,N_15462,N_15750);
or U16043 (N_16043,N_15412,N_15211);
nor U16044 (N_16044,N_15402,N_15598);
nor U16045 (N_16045,N_15311,N_15764);
xor U16046 (N_16046,N_15681,N_15434);
and U16047 (N_16047,N_15560,N_15865);
or U16048 (N_16048,N_15775,N_15386);
xor U16049 (N_16049,N_15640,N_15503);
and U16050 (N_16050,N_15584,N_15871);
or U16051 (N_16051,N_15318,N_15844);
nand U16052 (N_16052,N_15723,N_15758);
and U16053 (N_16053,N_15617,N_15532);
xnor U16054 (N_16054,N_15624,N_15677);
xnor U16055 (N_16055,N_15919,N_15546);
xnor U16056 (N_16056,N_15488,N_15392);
xor U16057 (N_16057,N_15482,N_15213);
nand U16058 (N_16058,N_15798,N_15999);
nor U16059 (N_16059,N_15303,N_15446);
and U16060 (N_16060,N_15698,N_15545);
xor U16061 (N_16061,N_15674,N_15689);
xnor U16062 (N_16062,N_15652,N_15934);
and U16063 (N_16063,N_15672,N_15280);
nand U16064 (N_16064,N_15406,N_15815);
xnor U16065 (N_16065,N_15626,N_15421);
nor U16066 (N_16066,N_15611,N_15904);
nand U16067 (N_16067,N_15832,N_15928);
nor U16068 (N_16068,N_15918,N_15490);
or U16069 (N_16069,N_15955,N_15900);
nand U16070 (N_16070,N_15308,N_15427);
xor U16071 (N_16071,N_15634,N_15550);
and U16072 (N_16072,N_15924,N_15248);
nand U16073 (N_16073,N_15466,N_15637);
xnor U16074 (N_16074,N_15302,N_15450);
nor U16075 (N_16075,N_15465,N_15739);
xnor U16076 (N_16076,N_15763,N_15370);
xor U16077 (N_16077,N_15461,N_15295);
or U16078 (N_16078,N_15791,N_15479);
nor U16079 (N_16079,N_15417,N_15389);
nand U16080 (N_16080,N_15331,N_15874);
nor U16081 (N_16081,N_15202,N_15423);
nand U16082 (N_16082,N_15443,N_15922);
nand U16083 (N_16083,N_15522,N_15237);
nor U16084 (N_16084,N_15937,N_15441);
nor U16085 (N_16085,N_15616,N_15769);
nand U16086 (N_16086,N_15338,N_15485);
xor U16087 (N_16087,N_15757,N_15231);
and U16088 (N_16088,N_15251,N_15580);
xnor U16089 (N_16089,N_15978,N_15381);
nor U16090 (N_16090,N_15639,N_15256);
nor U16091 (N_16091,N_15847,N_15263);
and U16092 (N_16092,N_15393,N_15930);
xnor U16093 (N_16093,N_15209,N_15878);
nor U16094 (N_16094,N_15828,N_15887);
nor U16095 (N_16095,N_15952,N_15578);
nor U16096 (N_16096,N_15364,N_15774);
and U16097 (N_16097,N_15458,N_15716);
nor U16098 (N_16098,N_15509,N_15495);
or U16099 (N_16099,N_15933,N_15729);
nor U16100 (N_16100,N_15980,N_15908);
or U16101 (N_16101,N_15850,N_15675);
or U16102 (N_16102,N_15759,N_15523);
xnor U16103 (N_16103,N_15380,N_15367);
and U16104 (N_16104,N_15956,N_15921);
xor U16105 (N_16105,N_15768,N_15464);
nor U16106 (N_16106,N_15968,N_15223);
or U16107 (N_16107,N_15736,N_15923);
and U16108 (N_16108,N_15990,N_15684);
xnor U16109 (N_16109,N_15241,N_15265);
nor U16110 (N_16110,N_15638,N_15820);
nand U16111 (N_16111,N_15363,N_15877);
and U16112 (N_16112,N_15893,N_15205);
xnor U16113 (N_16113,N_15244,N_15264);
nand U16114 (N_16114,N_15694,N_15827);
or U16115 (N_16115,N_15965,N_15797);
xnor U16116 (N_16116,N_15983,N_15521);
and U16117 (N_16117,N_15973,N_15253);
and U16118 (N_16118,N_15667,N_15470);
nand U16119 (N_16119,N_15917,N_15361);
nor U16120 (N_16120,N_15575,N_15299);
nor U16121 (N_16121,N_15399,N_15407);
xor U16122 (N_16122,N_15712,N_15754);
nor U16123 (N_16123,N_15801,N_15778);
or U16124 (N_16124,N_15208,N_15452);
and U16125 (N_16125,N_15972,N_15784);
nor U16126 (N_16126,N_15515,N_15853);
nand U16127 (N_16127,N_15779,N_15574);
nand U16128 (N_16128,N_15680,N_15332);
and U16129 (N_16129,N_15859,N_15950);
or U16130 (N_16130,N_15731,N_15701);
nor U16131 (N_16131,N_15636,N_15749);
nand U16132 (N_16132,N_15375,N_15994);
or U16133 (N_16133,N_15489,N_15535);
and U16134 (N_16134,N_15595,N_15321);
or U16135 (N_16135,N_15996,N_15218);
and U16136 (N_16136,N_15645,N_15862);
nor U16137 (N_16137,N_15666,N_15342);
nand U16138 (N_16138,N_15530,N_15304);
xnor U16139 (N_16139,N_15863,N_15653);
xnor U16140 (N_16140,N_15650,N_15305);
and U16141 (N_16141,N_15291,N_15390);
nor U16142 (N_16142,N_15704,N_15468);
xor U16143 (N_16143,N_15720,N_15500);
and U16144 (N_16144,N_15668,N_15843);
and U16145 (N_16145,N_15685,N_15876);
nor U16146 (N_16146,N_15313,N_15581);
nor U16147 (N_16147,N_15875,N_15662);
and U16148 (N_16148,N_15733,N_15591);
or U16149 (N_16149,N_15340,N_15569);
nand U16150 (N_16150,N_15225,N_15799);
and U16151 (N_16151,N_15814,N_15579);
or U16152 (N_16152,N_15945,N_15492);
or U16153 (N_16153,N_15848,N_15388);
nor U16154 (N_16154,N_15765,N_15686);
or U16155 (N_16155,N_15287,N_15235);
xnor U16156 (N_16156,N_15323,N_15345);
nor U16157 (N_16157,N_15409,N_15457);
and U16158 (N_16158,N_15912,N_15596);
or U16159 (N_16159,N_15573,N_15561);
xnor U16160 (N_16160,N_15629,N_15776);
xor U16161 (N_16161,N_15947,N_15220);
nand U16162 (N_16162,N_15601,N_15346);
xnor U16163 (N_16163,N_15885,N_15800);
xor U16164 (N_16164,N_15661,N_15722);
nand U16165 (N_16165,N_15589,N_15391);
and U16166 (N_16166,N_15376,N_15802);
and U16167 (N_16167,N_15431,N_15206);
nand U16168 (N_16168,N_15665,N_15200);
xnor U16169 (N_16169,N_15794,N_15469);
nor U16170 (N_16170,N_15335,N_15210);
nand U16171 (N_16171,N_15533,N_15927);
nor U16172 (N_16172,N_15891,N_15880);
or U16173 (N_16173,N_15935,N_15803);
nor U16174 (N_16174,N_15384,N_15795);
nor U16175 (N_16175,N_15455,N_15842);
or U16176 (N_16176,N_15460,N_15958);
and U16177 (N_16177,N_15760,N_15325);
nand U16178 (N_16178,N_15873,N_15986);
and U16179 (N_16179,N_15373,N_15627);
and U16180 (N_16180,N_15262,N_15824);
xor U16181 (N_16181,N_15849,N_15328);
xor U16182 (N_16182,N_15362,N_15517);
nor U16183 (N_16183,N_15702,N_15552);
or U16184 (N_16184,N_15770,N_15805);
nand U16185 (N_16185,N_15472,N_15230);
nor U16186 (N_16186,N_15333,N_15710);
or U16187 (N_16187,N_15394,N_15603);
nand U16188 (N_16188,N_15493,N_15426);
or U16189 (N_16189,N_15889,N_15337);
xnor U16190 (N_16190,N_15796,N_15883);
and U16191 (N_16191,N_15679,N_15925);
or U16192 (N_16192,N_15692,N_15851);
xnor U16193 (N_16193,N_15740,N_15314);
nand U16194 (N_16194,N_15215,N_15548);
nor U16195 (N_16195,N_15920,N_15816);
or U16196 (N_16196,N_15440,N_15728);
or U16197 (N_16197,N_15201,N_15551);
xor U16198 (N_16198,N_15780,N_15269);
nor U16199 (N_16199,N_15946,N_15825);
nor U16200 (N_16200,N_15673,N_15261);
and U16201 (N_16201,N_15518,N_15711);
and U16202 (N_16202,N_15631,N_15970);
nand U16203 (N_16203,N_15898,N_15477);
nor U16204 (N_16204,N_15741,N_15504);
nor U16205 (N_16205,N_15926,N_15812);
xnor U16206 (N_16206,N_15382,N_15275);
nand U16207 (N_16207,N_15538,N_15646);
nor U16208 (N_16208,N_15676,N_15993);
nor U16209 (N_16209,N_15300,N_15752);
or U16210 (N_16210,N_15654,N_15756);
nor U16211 (N_16211,N_15602,N_15761);
nand U16212 (N_16212,N_15985,N_15823);
or U16213 (N_16213,N_15613,N_15991);
nand U16214 (N_16214,N_15571,N_15669);
nor U16215 (N_16215,N_15910,N_15204);
nor U16216 (N_16216,N_15310,N_15288);
xor U16217 (N_16217,N_15683,N_15713);
nor U16218 (N_16218,N_15753,N_15378);
nand U16219 (N_16219,N_15238,N_15463);
and U16220 (N_16220,N_15811,N_15356);
nor U16221 (N_16221,N_15837,N_15566);
nor U16222 (N_16222,N_15353,N_15747);
nand U16223 (N_16223,N_15582,N_15425);
and U16224 (N_16224,N_15742,N_15424);
xnor U16225 (N_16225,N_15577,N_15433);
or U16226 (N_16226,N_15343,N_15326);
nor U16227 (N_16227,N_15395,N_15419);
nor U16228 (N_16228,N_15396,N_15840);
xor U16229 (N_16229,N_15895,N_15772);
nand U16230 (N_16230,N_15830,N_15312);
nor U16231 (N_16231,N_15969,N_15719);
nor U16232 (N_16232,N_15852,N_15355);
xnor U16233 (N_16233,N_15870,N_15594);
or U16234 (N_16234,N_15246,N_15833);
nand U16235 (N_16235,N_15705,N_15483);
xor U16236 (N_16236,N_15995,N_15212);
and U16237 (N_16237,N_15902,N_15252);
nand U16238 (N_16238,N_15216,N_15953);
or U16239 (N_16239,N_15558,N_15383);
and U16240 (N_16240,N_15534,N_15525);
nor U16241 (N_16241,N_15415,N_15987);
nand U16242 (N_16242,N_15881,N_15348);
nand U16243 (N_16243,N_15838,N_15943);
or U16244 (N_16244,N_15715,N_15785);
nor U16245 (N_16245,N_15588,N_15621);
or U16246 (N_16246,N_15413,N_15903);
nand U16247 (N_16247,N_15869,N_15240);
nand U16248 (N_16248,N_15687,N_15309);
nand U16249 (N_16249,N_15771,N_15568);
nand U16250 (N_16250,N_15691,N_15408);
and U16251 (N_16251,N_15320,N_15782);
nand U16252 (N_16252,N_15351,N_15975);
or U16253 (N_16253,N_15512,N_15693);
xnor U16254 (N_16254,N_15767,N_15451);
nor U16255 (N_16255,N_15897,N_15911);
or U16256 (N_16256,N_15257,N_15284);
and U16257 (N_16257,N_15285,N_15414);
xnor U16258 (N_16258,N_15514,N_15860);
nor U16259 (N_16259,N_15336,N_15454);
or U16260 (N_16260,N_15502,N_15615);
nand U16261 (N_16261,N_15203,N_15647);
nor U16262 (N_16262,N_15855,N_15334);
or U16263 (N_16263,N_15642,N_15377);
nor U16264 (N_16264,N_15254,N_15670);
or U16265 (N_16265,N_15344,N_15826);
nor U16266 (N_16266,N_15366,N_15938);
nor U16267 (N_16267,N_15296,N_15721);
xnor U16268 (N_16268,N_15316,N_15270);
and U16269 (N_16269,N_15411,N_15909);
nand U16270 (N_16270,N_15717,N_15709);
nor U16271 (N_16271,N_15727,N_15781);
nand U16272 (N_16272,N_15835,N_15549);
xnor U16273 (N_16273,N_15804,N_15743);
xor U16274 (N_16274,N_15540,N_15773);
and U16275 (N_16275,N_15416,N_15398);
xnor U16276 (N_16276,N_15576,N_15690);
and U16277 (N_16277,N_15599,N_15703);
nand U16278 (N_16278,N_15998,N_15682);
nor U16279 (N_16279,N_15671,N_15593);
or U16280 (N_16280,N_15536,N_15981);
xor U16281 (N_16281,N_15586,N_15531);
nor U16282 (N_16282,N_15967,N_15400);
nor U16283 (N_16283,N_15528,N_15699);
nand U16284 (N_16284,N_15663,N_15700);
nor U16285 (N_16285,N_15783,N_15232);
xor U16286 (N_16286,N_15524,N_15890);
and U16287 (N_16287,N_15324,N_15371);
nand U16288 (N_16288,N_15527,N_15319);
xnor U16289 (N_16289,N_15678,N_15537);
nor U16290 (N_16290,N_15447,N_15625);
nand U16291 (N_16291,N_15435,N_15359);
and U16292 (N_16292,N_15648,N_15725);
and U16293 (N_16293,N_15872,N_15744);
and U16294 (N_16294,N_15506,N_15276);
xor U16295 (N_16295,N_15879,N_15478);
nand U16296 (N_16296,N_15813,N_15587);
and U16297 (N_16297,N_15793,N_15818);
nor U16298 (N_16298,N_15553,N_15526);
xnor U16299 (N_16299,N_15884,N_15997);
and U16300 (N_16300,N_15854,N_15255);
and U16301 (N_16301,N_15856,N_15499);
or U16302 (N_16302,N_15266,N_15449);
and U16303 (N_16303,N_15992,N_15623);
or U16304 (N_16304,N_15706,N_15268);
xor U16305 (N_16305,N_15695,N_15708);
or U16306 (N_16306,N_15606,N_15282);
xnor U16307 (N_16307,N_15944,N_15583);
nor U16308 (N_16308,N_15372,N_15916);
and U16309 (N_16309,N_15605,N_15628);
and U16310 (N_16310,N_15307,N_15283);
and U16311 (N_16311,N_15866,N_15554);
xnor U16312 (N_16312,N_15258,N_15429);
xor U16313 (N_16313,N_15792,N_15387);
xnor U16314 (N_16314,N_15279,N_15730);
or U16315 (N_16315,N_15471,N_15913);
nor U16316 (N_16316,N_15260,N_15539);
or U16317 (N_16317,N_15520,N_15529);
xnor U16318 (N_16318,N_15660,N_15547);
xnor U16319 (N_16319,N_15239,N_15473);
nand U16320 (N_16320,N_15559,N_15732);
nand U16321 (N_16321,N_15379,N_15562);
nor U16322 (N_16322,N_15868,N_15397);
and U16323 (N_16323,N_15290,N_15475);
and U16324 (N_16324,N_15789,N_15988);
nor U16325 (N_16325,N_15281,N_15437);
and U16326 (N_16326,N_15608,N_15697);
xor U16327 (N_16327,N_15567,N_15315);
nand U16328 (N_16328,N_15734,N_15233);
xor U16329 (N_16329,N_15222,N_15510);
nor U16330 (N_16330,N_15819,N_15585);
and U16331 (N_16331,N_15592,N_15542);
nand U16332 (N_16332,N_15317,N_15762);
nand U16333 (N_16333,N_15726,N_15352);
nand U16334 (N_16334,N_15420,N_15217);
nand U16335 (N_16335,N_15436,N_15259);
xnor U16336 (N_16336,N_15347,N_15755);
nor U16337 (N_16337,N_15864,N_15907);
xor U16338 (N_16338,N_15949,N_15766);
nor U16339 (N_16339,N_15272,N_15610);
nand U16340 (N_16340,N_15516,N_15278);
nor U16341 (N_16341,N_15339,N_15959);
or U16342 (N_16342,N_15788,N_15619);
nor U16343 (N_16343,N_15932,N_15836);
nand U16344 (N_16344,N_15831,N_15511);
nand U16345 (N_16345,N_15809,N_15894);
nor U16346 (N_16346,N_15688,N_15267);
nor U16347 (N_16347,N_15250,N_15354);
and U16348 (N_16348,N_15403,N_15806);
nor U16349 (N_16349,N_15273,N_15810);
or U16350 (N_16350,N_15476,N_15497);
or U16351 (N_16351,N_15751,N_15620);
and U16352 (N_16352,N_15618,N_15982);
nand U16353 (N_16353,N_15507,N_15839);
nand U16354 (N_16354,N_15845,N_15544);
xnor U16355 (N_16355,N_15861,N_15459);
xor U16356 (N_16356,N_15564,N_15964);
nor U16357 (N_16357,N_15867,N_15971);
and U16358 (N_16358,N_15570,N_15963);
nand U16359 (N_16359,N_15822,N_15936);
nor U16360 (N_16360,N_15368,N_15484);
and U16361 (N_16361,N_15906,N_15630);
and U16362 (N_16362,N_15245,N_15960);
or U16363 (N_16363,N_15214,N_15714);
xor U16364 (N_16364,N_15633,N_15572);
and U16365 (N_16365,N_15243,N_15846);
nor U16366 (N_16366,N_15655,N_15505);
nand U16367 (N_16367,N_15249,N_15644);
nor U16368 (N_16368,N_15808,N_15737);
nand U16369 (N_16369,N_15857,N_15496);
and U16370 (N_16370,N_15519,N_15271);
or U16371 (N_16371,N_15977,N_15428);
xnor U16372 (N_16372,N_15491,N_15234);
nand U16373 (N_16373,N_15748,N_15349);
nor U16374 (N_16374,N_15915,N_15664);
or U16375 (N_16375,N_15543,N_15957);
and U16376 (N_16376,N_15486,N_15886);
or U16377 (N_16377,N_15777,N_15600);
nor U16378 (N_16378,N_15228,N_15607);
nand U16379 (N_16379,N_15467,N_15557);
or U16380 (N_16380,N_15905,N_15289);
and U16381 (N_16381,N_15696,N_15931);
and U16382 (N_16382,N_15656,N_15614);
nand U16383 (N_16383,N_15896,N_15882);
or U16384 (N_16384,N_15219,N_15298);
nand U16385 (N_16385,N_15226,N_15498);
nand U16386 (N_16386,N_15735,N_15445);
xnor U16387 (N_16387,N_15829,N_15481);
and U16388 (N_16388,N_15609,N_15834);
and U16389 (N_16389,N_15401,N_15807);
nand U16390 (N_16390,N_15541,N_15962);
xnor U16391 (N_16391,N_15229,N_15247);
nand U16392 (N_16392,N_15659,N_15565);
or U16393 (N_16393,N_15786,N_15274);
nand U16394 (N_16394,N_15718,N_15358);
nor U16395 (N_16395,N_15350,N_15360);
nor U16396 (N_16396,N_15242,N_15357);
xor U16397 (N_16397,N_15277,N_15966);
xor U16398 (N_16398,N_15404,N_15597);
or U16399 (N_16399,N_15444,N_15487);
nand U16400 (N_16400,N_15415,N_15658);
or U16401 (N_16401,N_15657,N_15699);
xnor U16402 (N_16402,N_15940,N_15749);
and U16403 (N_16403,N_15933,N_15394);
nor U16404 (N_16404,N_15606,N_15454);
xor U16405 (N_16405,N_15682,N_15749);
xor U16406 (N_16406,N_15467,N_15349);
and U16407 (N_16407,N_15755,N_15949);
nand U16408 (N_16408,N_15691,N_15972);
nor U16409 (N_16409,N_15408,N_15378);
xnor U16410 (N_16410,N_15963,N_15314);
or U16411 (N_16411,N_15875,N_15819);
and U16412 (N_16412,N_15360,N_15902);
and U16413 (N_16413,N_15620,N_15983);
or U16414 (N_16414,N_15238,N_15880);
and U16415 (N_16415,N_15437,N_15717);
and U16416 (N_16416,N_15585,N_15385);
or U16417 (N_16417,N_15472,N_15759);
xnor U16418 (N_16418,N_15660,N_15320);
nor U16419 (N_16419,N_15744,N_15961);
xnor U16420 (N_16420,N_15688,N_15532);
nand U16421 (N_16421,N_15763,N_15762);
or U16422 (N_16422,N_15410,N_15848);
or U16423 (N_16423,N_15810,N_15984);
nand U16424 (N_16424,N_15382,N_15977);
nand U16425 (N_16425,N_15671,N_15327);
nand U16426 (N_16426,N_15399,N_15963);
or U16427 (N_16427,N_15500,N_15371);
nand U16428 (N_16428,N_15683,N_15861);
nand U16429 (N_16429,N_15643,N_15273);
xor U16430 (N_16430,N_15259,N_15396);
nor U16431 (N_16431,N_15879,N_15480);
nor U16432 (N_16432,N_15814,N_15823);
xor U16433 (N_16433,N_15463,N_15371);
and U16434 (N_16434,N_15596,N_15297);
nand U16435 (N_16435,N_15857,N_15965);
and U16436 (N_16436,N_15535,N_15670);
nand U16437 (N_16437,N_15989,N_15283);
nand U16438 (N_16438,N_15662,N_15997);
nand U16439 (N_16439,N_15526,N_15799);
xor U16440 (N_16440,N_15564,N_15225);
nor U16441 (N_16441,N_15793,N_15744);
nand U16442 (N_16442,N_15561,N_15697);
nor U16443 (N_16443,N_15941,N_15517);
nand U16444 (N_16444,N_15845,N_15445);
and U16445 (N_16445,N_15322,N_15394);
nand U16446 (N_16446,N_15806,N_15875);
xor U16447 (N_16447,N_15241,N_15773);
and U16448 (N_16448,N_15396,N_15953);
nor U16449 (N_16449,N_15694,N_15685);
nand U16450 (N_16450,N_15909,N_15513);
or U16451 (N_16451,N_15234,N_15812);
or U16452 (N_16452,N_15504,N_15897);
or U16453 (N_16453,N_15897,N_15348);
or U16454 (N_16454,N_15849,N_15370);
or U16455 (N_16455,N_15656,N_15556);
xor U16456 (N_16456,N_15407,N_15496);
xnor U16457 (N_16457,N_15373,N_15212);
xnor U16458 (N_16458,N_15532,N_15430);
and U16459 (N_16459,N_15302,N_15754);
nor U16460 (N_16460,N_15314,N_15651);
nor U16461 (N_16461,N_15461,N_15656);
nor U16462 (N_16462,N_15595,N_15754);
nand U16463 (N_16463,N_15959,N_15691);
nor U16464 (N_16464,N_15913,N_15945);
xor U16465 (N_16465,N_15245,N_15852);
nand U16466 (N_16466,N_15527,N_15386);
nor U16467 (N_16467,N_15300,N_15356);
and U16468 (N_16468,N_15763,N_15391);
or U16469 (N_16469,N_15707,N_15551);
or U16470 (N_16470,N_15405,N_15321);
nor U16471 (N_16471,N_15805,N_15917);
and U16472 (N_16472,N_15369,N_15412);
and U16473 (N_16473,N_15903,N_15989);
nand U16474 (N_16474,N_15438,N_15472);
xor U16475 (N_16475,N_15621,N_15657);
xor U16476 (N_16476,N_15298,N_15366);
or U16477 (N_16477,N_15366,N_15732);
nor U16478 (N_16478,N_15943,N_15885);
or U16479 (N_16479,N_15294,N_15463);
and U16480 (N_16480,N_15349,N_15374);
or U16481 (N_16481,N_15222,N_15626);
and U16482 (N_16482,N_15717,N_15942);
xnor U16483 (N_16483,N_15945,N_15804);
nand U16484 (N_16484,N_15573,N_15470);
and U16485 (N_16485,N_15583,N_15953);
or U16486 (N_16486,N_15983,N_15636);
nor U16487 (N_16487,N_15227,N_15730);
or U16488 (N_16488,N_15554,N_15965);
xor U16489 (N_16489,N_15709,N_15357);
nand U16490 (N_16490,N_15704,N_15391);
nand U16491 (N_16491,N_15314,N_15592);
nand U16492 (N_16492,N_15350,N_15841);
and U16493 (N_16493,N_15607,N_15340);
nor U16494 (N_16494,N_15649,N_15470);
and U16495 (N_16495,N_15953,N_15619);
and U16496 (N_16496,N_15321,N_15594);
xnor U16497 (N_16497,N_15511,N_15730);
nor U16498 (N_16498,N_15793,N_15489);
nor U16499 (N_16499,N_15666,N_15239);
and U16500 (N_16500,N_15344,N_15523);
and U16501 (N_16501,N_15675,N_15376);
xnor U16502 (N_16502,N_15963,N_15307);
nand U16503 (N_16503,N_15896,N_15227);
and U16504 (N_16504,N_15933,N_15338);
nor U16505 (N_16505,N_15821,N_15986);
or U16506 (N_16506,N_15635,N_15471);
nand U16507 (N_16507,N_15530,N_15430);
or U16508 (N_16508,N_15275,N_15535);
and U16509 (N_16509,N_15903,N_15739);
nor U16510 (N_16510,N_15528,N_15567);
xor U16511 (N_16511,N_15860,N_15252);
nor U16512 (N_16512,N_15790,N_15768);
nor U16513 (N_16513,N_15356,N_15810);
xor U16514 (N_16514,N_15367,N_15262);
nand U16515 (N_16515,N_15442,N_15250);
nand U16516 (N_16516,N_15796,N_15248);
or U16517 (N_16517,N_15870,N_15398);
or U16518 (N_16518,N_15678,N_15998);
or U16519 (N_16519,N_15336,N_15576);
xor U16520 (N_16520,N_15742,N_15323);
nand U16521 (N_16521,N_15879,N_15870);
or U16522 (N_16522,N_15398,N_15703);
xnor U16523 (N_16523,N_15696,N_15517);
xnor U16524 (N_16524,N_15623,N_15337);
nand U16525 (N_16525,N_15589,N_15889);
nor U16526 (N_16526,N_15645,N_15209);
nand U16527 (N_16527,N_15358,N_15699);
or U16528 (N_16528,N_15501,N_15245);
nor U16529 (N_16529,N_15877,N_15489);
xnor U16530 (N_16530,N_15433,N_15779);
nand U16531 (N_16531,N_15419,N_15407);
nor U16532 (N_16532,N_15587,N_15427);
or U16533 (N_16533,N_15854,N_15712);
nand U16534 (N_16534,N_15895,N_15396);
nand U16535 (N_16535,N_15984,N_15491);
or U16536 (N_16536,N_15748,N_15545);
nor U16537 (N_16537,N_15849,N_15630);
or U16538 (N_16538,N_15769,N_15356);
nor U16539 (N_16539,N_15543,N_15432);
nand U16540 (N_16540,N_15377,N_15846);
nor U16541 (N_16541,N_15805,N_15371);
and U16542 (N_16542,N_15255,N_15246);
nor U16543 (N_16543,N_15953,N_15644);
nor U16544 (N_16544,N_15788,N_15737);
or U16545 (N_16545,N_15339,N_15496);
nor U16546 (N_16546,N_15399,N_15274);
or U16547 (N_16547,N_15691,N_15679);
nor U16548 (N_16548,N_15686,N_15715);
xor U16549 (N_16549,N_15248,N_15608);
nand U16550 (N_16550,N_15442,N_15220);
nor U16551 (N_16551,N_15747,N_15758);
nor U16552 (N_16552,N_15898,N_15626);
and U16553 (N_16553,N_15383,N_15753);
and U16554 (N_16554,N_15543,N_15783);
nand U16555 (N_16555,N_15936,N_15575);
and U16556 (N_16556,N_15350,N_15278);
and U16557 (N_16557,N_15887,N_15723);
nor U16558 (N_16558,N_15452,N_15424);
xnor U16559 (N_16559,N_15810,N_15858);
xor U16560 (N_16560,N_15770,N_15503);
and U16561 (N_16561,N_15426,N_15293);
nor U16562 (N_16562,N_15949,N_15343);
nor U16563 (N_16563,N_15727,N_15655);
and U16564 (N_16564,N_15435,N_15559);
or U16565 (N_16565,N_15446,N_15717);
or U16566 (N_16566,N_15667,N_15637);
and U16567 (N_16567,N_15579,N_15330);
nand U16568 (N_16568,N_15934,N_15365);
or U16569 (N_16569,N_15558,N_15693);
nor U16570 (N_16570,N_15231,N_15868);
nor U16571 (N_16571,N_15755,N_15701);
nand U16572 (N_16572,N_15715,N_15346);
xnor U16573 (N_16573,N_15655,N_15528);
nand U16574 (N_16574,N_15304,N_15495);
nor U16575 (N_16575,N_15224,N_15672);
nor U16576 (N_16576,N_15992,N_15867);
xor U16577 (N_16577,N_15909,N_15799);
or U16578 (N_16578,N_15913,N_15765);
nor U16579 (N_16579,N_15443,N_15339);
nor U16580 (N_16580,N_15954,N_15960);
or U16581 (N_16581,N_15212,N_15863);
and U16582 (N_16582,N_15458,N_15341);
xor U16583 (N_16583,N_15554,N_15266);
xor U16584 (N_16584,N_15496,N_15777);
or U16585 (N_16585,N_15999,N_15598);
nor U16586 (N_16586,N_15639,N_15903);
xor U16587 (N_16587,N_15524,N_15413);
nand U16588 (N_16588,N_15258,N_15376);
nor U16589 (N_16589,N_15951,N_15994);
and U16590 (N_16590,N_15297,N_15923);
or U16591 (N_16591,N_15332,N_15568);
nor U16592 (N_16592,N_15407,N_15327);
nor U16593 (N_16593,N_15856,N_15231);
xor U16594 (N_16594,N_15941,N_15952);
nand U16595 (N_16595,N_15472,N_15322);
or U16596 (N_16596,N_15578,N_15281);
and U16597 (N_16597,N_15459,N_15487);
or U16598 (N_16598,N_15530,N_15671);
nor U16599 (N_16599,N_15278,N_15698);
nand U16600 (N_16600,N_15573,N_15698);
nor U16601 (N_16601,N_15267,N_15259);
xnor U16602 (N_16602,N_15371,N_15301);
nor U16603 (N_16603,N_15698,N_15476);
and U16604 (N_16604,N_15465,N_15635);
and U16605 (N_16605,N_15791,N_15400);
nor U16606 (N_16606,N_15827,N_15484);
nand U16607 (N_16607,N_15499,N_15554);
nor U16608 (N_16608,N_15476,N_15246);
xnor U16609 (N_16609,N_15802,N_15766);
nand U16610 (N_16610,N_15366,N_15365);
xor U16611 (N_16611,N_15212,N_15631);
or U16612 (N_16612,N_15879,N_15572);
or U16613 (N_16613,N_15555,N_15930);
nand U16614 (N_16614,N_15900,N_15765);
nor U16615 (N_16615,N_15369,N_15948);
xor U16616 (N_16616,N_15533,N_15660);
or U16617 (N_16617,N_15408,N_15786);
and U16618 (N_16618,N_15550,N_15950);
xor U16619 (N_16619,N_15863,N_15889);
nand U16620 (N_16620,N_15409,N_15811);
or U16621 (N_16621,N_15661,N_15289);
or U16622 (N_16622,N_15771,N_15310);
xor U16623 (N_16623,N_15253,N_15348);
xor U16624 (N_16624,N_15771,N_15421);
nor U16625 (N_16625,N_15725,N_15838);
xnor U16626 (N_16626,N_15995,N_15805);
nor U16627 (N_16627,N_15897,N_15960);
and U16628 (N_16628,N_15588,N_15631);
nand U16629 (N_16629,N_15782,N_15674);
and U16630 (N_16630,N_15462,N_15758);
nand U16631 (N_16631,N_15405,N_15267);
nor U16632 (N_16632,N_15968,N_15738);
and U16633 (N_16633,N_15779,N_15421);
or U16634 (N_16634,N_15275,N_15665);
nand U16635 (N_16635,N_15281,N_15833);
nor U16636 (N_16636,N_15697,N_15557);
nor U16637 (N_16637,N_15770,N_15834);
or U16638 (N_16638,N_15215,N_15537);
or U16639 (N_16639,N_15280,N_15579);
nor U16640 (N_16640,N_15456,N_15896);
and U16641 (N_16641,N_15982,N_15687);
nand U16642 (N_16642,N_15349,N_15940);
nor U16643 (N_16643,N_15241,N_15534);
xnor U16644 (N_16644,N_15502,N_15304);
or U16645 (N_16645,N_15700,N_15229);
nor U16646 (N_16646,N_15747,N_15712);
xnor U16647 (N_16647,N_15637,N_15944);
nor U16648 (N_16648,N_15603,N_15417);
and U16649 (N_16649,N_15403,N_15318);
or U16650 (N_16650,N_15329,N_15599);
xnor U16651 (N_16651,N_15367,N_15752);
nand U16652 (N_16652,N_15744,N_15698);
nand U16653 (N_16653,N_15942,N_15496);
nor U16654 (N_16654,N_15637,N_15266);
and U16655 (N_16655,N_15471,N_15914);
nor U16656 (N_16656,N_15664,N_15498);
xnor U16657 (N_16657,N_15952,N_15818);
xor U16658 (N_16658,N_15451,N_15959);
and U16659 (N_16659,N_15222,N_15742);
xor U16660 (N_16660,N_15606,N_15679);
nor U16661 (N_16661,N_15220,N_15624);
nand U16662 (N_16662,N_15640,N_15753);
nand U16663 (N_16663,N_15448,N_15573);
nor U16664 (N_16664,N_15939,N_15337);
and U16665 (N_16665,N_15713,N_15249);
or U16666 (N_16666,N_15212,N_15236);
nor U16667 (N_16667,N_15915,N_15978);
xor U16668 (N_16668,N_15347,N_15766);
nor U16669 (N_16669,N_15422,N_15864);
xnor U16670 (N_16670,N_15844,N_15284);
or U16671 (N_16671,N_15598,N_15678);
xor U16672 (N_16672,N_15305,N_15957);
xnor U16673 (N_16673,N_15427,N_15947);
and U16674 (N_16674,N_15982,N_15609);
xor U16675 (N_16675,N_15343,N_15341);
and U16676 (N_16676,N_15653,N_15982);
xor U16677 (N_16677,N_15568,N_15947);
or U16678 (N_16678,N_15592,N_15676);
xor U16679 (N_16679,N_15200,N_15757);
nor U16680 (N_16680,N_15221,N_15434);
and U16681 (N_16681,N_15865,N_15351);
nor U16682 (N_16682,N_15281,N_15550);
or U16683 (N_16683,N_15505,N_15612);
and U16684 (N_16684,N_15975,N_15451);
xnor U16685 (N_16685,N_15393,N_15254);
nor U16686 (N_16686,N_15800,N_15977);
or U16687 (N_16687,N_15481,N_15659);
or U16688 (N_16688,N_15614,N_15782);
and U16689 (N_16689,N_15710,N_15970);
xor U16690 (N_16690,N_15525,N_15524);
xnor U16691 (N_16691,N_15350,N_15731);
nor U16692 (N_16692,N_15374,N_15239);
or U16693 (N_16693,N_15764,N_15841);
nand U16694 (N_16694,N_15709,N_15404);
xnor U16695 (N_16695,N_15819,N_15787);
nor U16696 (N_16696,N_15674,N_15570);
or U16697 (N_16697,N_15792,N_15949);
nor U16698 (N_16698,N_15524,N_15503);
nand U16699 (N_16699,N_15749,N_15644);
nor U16700 (N_16700,N_15581,N_15945);
nand U16701 (N_16701,N_15595,N_15232);
nand U16702 (N_16702,N_15485,N_15788);
and U16703 (N_16703,N_15714,N_15222);
and U16704 (N_16704,N_15779,N_15509);
xnor U16705 (N_16705,N_15804,N_15234);
nor U16706 (N_16706,N_15222,N_15514);
or U16707 (N_16707,N_15883,N_15888);
and U16708 (N_16708,N_15971,N_15967);
and U16709 (N_16709,N_15407,N_15606);
or U16710 (N_16710,N_15726,N_15662);
xnor U16711 (N_16711,N_15800,N_15861);
or U16712 (N_16712,N_15837,N_15925);
xnor U16713 (N_16713,N_15645,N_15903);
or U16714 (N_16714,N_15516,N_15826);
and U16715 (N_16715,N_15494,N_15350);
xor U16716 (N_16716,N_15568,N_15890);
nor U16717 (N_16717,N_15365,N_15801);
nor U16718 (N_16718,N_15289,N_15389);
or U16719 (N_16719,N_15633,N_15656);
or U16720 (N_16720,N_15245,N_15568);
or U16721 (N_16721,N_15993,N_15768);
nand U16722 (N_16722,N_15835,N_15957);
nand U16723 (N_16723,N_15674,N_15668);
nor U16724 (N_16724,N_15506,N_15264);
xnor U16725 (N_16725,N_15635,N_15384);
and U16726 (N_16726,N_15762,N_15716);
xnor U16727 (N_16727,N_15623,N_15684);
nor U16728 (N_16728,N_15424,N_15621);
or U16729 (N_16729,N_15523,N_15936);
nor U16730 (N_16730,N_15941,N_15813);
nand U16731 (N_16731,N_15687,N_15765);
xnor U16732 (N_16732,N_15844,N_15431);
and U16733 (N_16733,N_15636,N_15885);
xor U16734 (N_16734,N_15964,N_15254);
xnor U16735 (N_16735,N_15302,N_15623);
nor U16736 (N_16736,N_15930,N_15785);
nand U16737 (N_16737,N_15788,N_15298);
or U16738 (N_16738,N_15696,N_15223);
xnor U16739 (N_16739,N_15828,N_15668);
nand U16740 (N_16740,N_15682,N_15971);
nor U16741 (N_16741,N_15240,N_15425);
nand U16742 (N_16742,N_15730,N_15356);
xor U16743 (N_16743,N_15310,N_15355);
xnor U16744 (N_16744,N_15232,N_15617);
xnor U16745 (N_16745,N_15383,N_15905);
xor U16746 (N_16746,N_15836,N_15945);
or U16747 (N_16747,N_15796,N_15928);
nand U16748 (N_16748,N_15530,N_15944);
and U16749 (N_16749,N_15798,N_15466);
xor U16750 (N_16750,N_15311,N_15830);
nor U16751 (N_16751,N_15514,N_15430);
nor U16752 (N_16752,N_15659,N_15393);
and U16753 (N_16753,N_15503,N_15808);
or U16754 (N_16754,N_15969,N_15699);
nand U16755 (N_16755,N_15431,N_15891);
or U16756 (N_16756,N_15632,N_15675);
nand U16757 (N_16757,N_15321,N_15620);
or U16758 (N_16758,N_15211,N_15523);
and U16759 (N_16759,N_15378,N_15203);
nor U16760 (N_16760,N_15282,N_15233);
and U16761 (N_16761,N_15682,N_15353);
nand U16762 (N_16762,N_15834,N_15347);
or U16763 (N_16763,N_15610,N_15516);
and U16764 (N_16764,N_15360,N_15747);
nand U16765 (N_16765,N_15385,N_15396);
or U16766 (N_16766,N_15375,N_15763);
and U16767 (N_16767,N_15285,N_15342);
nand U16768 (N_16768,N_15934,N_15387);
nand U16769 (N_16769,N_15599,N_15951);
or U16770 (N_16770,N_15688,N_15543);
or U16771 (N_16771,N_15697,N_15382);
xor U16772 (N_16772,N_15453,N_15570);
nor U16773 (N_16773,N_15783,N_15238);
nand U16774 (N_16774,N_15729,N_15674);
nand U16775 (N_16775,N_15465,N_15799);
nand U16776 (N_16776,N_15299,N_15419);
nor U16777 (N_16777,N_15289,N_15612);
xnor U16778 (N_16778,N_15512,N_15952);
and U16779 (N_16779,N_15944,N_15782);
nand U16780 (N_16780,N_15817,N_15891);
and U16781 (N_16781,N_15925,N_15236);
nor U16782 (N_16782,N_15578,N_15610);
nand U16783 (N_16783,N_15901,N_15458);
xnor U16784 (N_16784,N_15592,N_15875);
nor U16785 (N_16785,N_15708,N_15731);
or U16786 (N_16786,N_15801,N_15794);
xnor U16787 (N_16787,N_15619,N_15579);
or U16788 (N_16788,N_15742,N_15655);
nand U16789 (N_16789,N_15508,N_15590);
or U16790 (N_16790,N_15503,N_15599);
nand U16791 (N_16791,N_15555,N_15431);
nand U16792 (N_16792,N_15887,N_15524);
nor U16793 (N_16793,N_15980,N_15923);
xor U16794 (N_16794,N_15441,N_15861);
or U16795 (N_16795,N_15522,N_15884);
or U16796 (N_16796,N_15447,N_15418);
nand U16797 (N_16797,N_15675,N_15968);
nor U16798 (N_16798,N_15839,N_15900);
and U16799 (N_16799,N_15725,N_15816);
nand U16800 (N_16800,N_16243,N_16439);
and U16801 (N_16801,N_16650,N_16033);
or U16802 (N_16802,N_16707,N_16431);
and U16803 (N_16803,N_16497,N_16677);
nor U16804 (N_16804,N_16488,N_16610);
xor U16805 (N_16805,N_16603,N_16055);
xnor U16806 (N_16806,N_16391,N_16366);
and U16807 (N_16807,N_16796,N_16302);
or U16808 (N_16808,N_16552,N_16522);
or U16809 (N_16809,N_16674,N_16535);
or U16810 (N_16810,N_16581,N_16763);
nand U16811 (N_16811,N_16339,N_16626);
nand U16812 (N_16812,N_16480,N_16655);
xnor U16813 (N_16813,N_16031,N_16114);
and U16814 (N_16814,N_16649,N_16423);
nor U16815 (N_16815,N_16249,N_16173);
or U16816 (N_16816,N_16560,N_16717);
nor U16817 (N_16817,N_16790,N_16442);
nor U16818 (N_16818,N_16183,N_16182);
nor U16819 (N_16819,N_16609,N_16619);
and U16820 (N_16820,N_16342,N_16333);
xor U16821 (N_16821,N_16065,N_16537);
nor U16822 (N_16822,N_16686,N_16624);
nand U16823 (N_16823,N_16365,N_16135);
and U16824 (N_16824,N_16235,N_16679);
nand U16825 (N_16825,N_16787,N_16505);
xor U16826 (N_16826,N_16292,N_16229);
nor U16827 (N_16827,N_16547,N_16022);
or U16828 (N_16828,N_16580,N_16407);
nor U16829 (N_16829,N_16574,N_16290);
or U16830 (N_16830,N_16553,N_16638);
or U16831 (N_16831,N_16572,N_16565);
nor U16832 (N_16832,N_16490,N_16241);
xor U16833 (N_16833,N_16710,N_16545);
or U16834 (N_16834,N_16095,N_16596);
or U16835 (N_16835,N_16384,N_16299);
nand U16836 (N_16836,N_16563,N_16516);
and U16837 (N_16837,N_16036,N_16695);
xnor U16838 (N_16838,N_16670,N_16434);
and U16839 (N_16839,N_16701,N_16607);
nor U16840 (N_16840,N_16077,N_16589);
and U16841 (N_16841,N_16437,N_16795);
xnor U16842 (N_16842,N_16665,N_16136);
and U16843 (N_16843,N_16378,N_16304);
or U16844 (N_16844,N_16383,N_16094);
nand U16845 (N_16845,N_16016,N_16006);
nor U16846 (N_16846,N_16419,N_16747);
nor U16847 (N_16847,N_16129,N_16486);
or U16848 (N_16848,N_16716,N_16174);
or U16849 (N_16849,N_16557,N_16335);
nor U16850 (N_16850,N_16023,N_16472);
nand U16851 (N_16851,N_16513,N_16770);
or U16852 (N_16852,N_16792,N_16520);
or U16853 (N_16853,N_16237,N_16201);
or U16854 (N_16854,N_16402,N_16024);
nor U16855 (N_16855,N_16138,N_16410);
nor U16856 (N_16856,N_16039,N_16785);
and U16857 (N_16857,N_16131,N_16425);
nor U16858 (N_16858,N_16777,N_16675);
nand U16859 (N_16859,N_16758,N_16618);
or U16860 (N_16860,N_16027,N_16519);
xnor U16861 (N_16861,N_16064,N_16026);
and U16862 (N_16862,N_16773,N_16592);
or U16863 (N_16863,N_16736,N_16528);
nor U16864 (N_16864,N_16145,N_16643);
xnor U16865 (N_16865,N_16030,N_16045);
nand U16866 (N_16866,N_16463,N_16126);
xor U16867 (N_16867,N_16275,N_16521);
nor U16868 (N_16868,N_16307,N_16503);
xor U16869 (N_16869,N_16583,N_16089);
nand U16870 (N_16870,N_16496,N_16133);
or U16871 (N_16871,N_16123,N_16731);
nand U16872 (N_16872,N_16298,N_16197);
and U16873 (N_16873,N_16398,N_16042);
xor U16874 (N_16874,N_16056,N_16086);
and U16875 (N_16875,N_16714,N_16050);
nand U16876 (N_16876,N_16103,N_16169);
xor U16877 (N_16877,N_16191,N_16449);
xor U16878 (N_16878,N_16220,N_16729);
xor U16879 (N_16879,N_16566,N_16376);
xnor U16880 (N_16880,N_16680,N_16272);
xnor U16881 (N_16881,N_16778,N_16389);
or U16882 (N_16882,N_16361,N_16653);
or U16883 (N_16883,N_16689,N_16044);
nand U16884 (N_16884,N_16692,N_16660);
and U16885 (N_16885,N_16484,N_16084);
nand U16886 (N_16886,N_16744,N_16356);
nor U16887 (N_16887,N_16755,N_16189);
and U16888 (N_16888,N_16541,N_16739);
nor U16889 (N_16889,N_16500,N_16244);
nand U16890 (N_16890,N_16119,N_16578);
and U16891 (N_16891,N_16712,N_16097);
and U16892 (N_16892,N_16501,N_16446);
and U16893 (N_16893,N_16113,N_16034);
or U16894 (N_16894,N_16332,N_16186);
nor U16895 (N_16895,N_16313,N_16029);
nand U16896 (N_16896,N_16386,N_16222);
xnor U16897 (N_16897,N_16526,N_16720);
xor U16898 (N_16898,N_16122,N_16794);
xor U16899 (N_16899,N_16028,N_16416);
or U16900 (N_16900,N_16748,N_16047);
and U16901 (N_16901,N_16098,N_16651);
xnor U16902 (N_16902,N_16454,N_16105);
and U16903 (N_16903,N_16198,N_16715);
nor U16904 (N_16904,N_16221,N_16171);
nand U16905 (N_16905,N_16080,N_16424);
or U16906 (N_16906,N_16569,N_16153);
and U16907 (N_16907,N_16190,N_16448);
or U16908 (N_16908,N_16268,N_16057);
nand U16909 (N_16909,N_16540,N_16276);
and U16910 (N_16910,N_16768,N_16432);
xor U16911 (N_16911,N_16600,N_16372);
nor U16912 (N_16912,N_16300,N_16703);
and U16913 (N_16913,N_16798,N_16476);
and U16914 (N_16914,N_16784,N_16512);
nor U16915 (N_16915,N_16783,N_16181);
or U16916 (N_16916,N_16518,N_16387);
and U16917 (N_16917,N_16346,N_16324);
xnor U16918 (N_16918,N_16457,N_16087);
xnor U16919 (N_16919,N_16004,N_16757);
and U16920 (N_16920,N_16724,N_16168);
nand U16921 (N_16921,N_16762,N_16000);
or U16922 (N_16922,N_16265,N_16282);
and U16923 (N_16923,N_16631,N_16752);
nand U16924 (N_16924,N_16465,N_16533);
or U16925 (N_16925,N_16451,N_16749);
xor U16926 (N_16926,N_16306,N_16068);
nor U16927 (N_16927,N_16614,N_16397);
or U16928 (N_16928,N_16212,N_16331);
nor U16929 (N_16929,N_16444,N_16699);
nor U16930 (N_16930,N_16668,N_16115);
nand U16931 (N_16931,N_16112,N_16188);
and U16932 (N_16932,N_16577,N_16037);
or U16933 (N_16933,N_16382,N_16672);
and U16934 (N_16934,N_16256,N_16127);
and U16935 (N_16935,N_16194,N_16110);
and U16936 (N_16936,N_16279,N_16645);
nand U16937 (N_16937,N_16640,N_16470);
nor U16938 (N_16938,N_16775,N_16259);
or U16939 (N_16939,N_16452,N_16664);
xnor U16940 (N_16940,N_16453,N_16481);
or U16941 (N_16941,N_16370,N_16532);
nand U16942 (N_16942,N_16392,N_16791);
nor U16943 (N_16943,N_16013,N_16049);
nor U16944 (N_16944,N_16344,N_16585);
xnor U16945 (N_16945,N_16124,N_16247);
xor U16946 (N_16946,N_16534,N_16628);
nor U16947 (N_16947,N_16662,N_16329);
nor U16948 (N_16948,N_16559,N_16184);
and U16949 (N_16949,N_16269,N_16682);
nand U16950 (N_16950,N_16374,N_16285);
nor U16951 (N_16951,N_16621,N_16311);
and U16952 (N_16952,N_16165,N_16789);
xor U16953 (N_16953,N_16422,N_16576);
xor U16954 (N_16954,N_16380,N_16719);
nand U16955 (N_16955,N_16007,N_16108);
nor U16956 (N_16956,N_16350,N_16334);
and U16957 (N_16957,N_16711,N_16733);
nor U16958 (N_16958,N_16678,N_16730);
xnor U16959 (N_16959,N_16761,N_16627);
or U16960 (N_16960,N_16633,N_16231);
nor U16961 (N_16961,N_16063,N_16353);
nor U16962 (N_16962,N_16141,N_16687);
or U16963 (N_16963,N_16082,N_16012);
or U16964 (N_16964,N_16230,N_16694);
nand U16965 (N_16965,N_16054,N_16504);
xor U16966 (N_16966,N_16517,N_16142);
nor U16967 (N_16967,N_16475,N_16208);
and U16968 (N_16968,N_16240,N_16414);
and U16969 (N_16969,N_16107,N_16009);
nor U16970 (N_16970,N_16742,N_16032);
nand U16971 (N_16971,N_16360,N_16759);
nor U16972 (N_16972,N_16642,N_16588);
nand U16973 (N_16973,N_16284,N_16413);
xor U16974 (N_16974,N_16654,N_16652);
or U16975 (N_16975,N_16223,N_16002);
or U16976 (N_16976,N_16359,N_16255);
nand U16977 (N_16977,N_16530,N_16330);
or U16978 (N_16978,N_16499,N_16176);
nand U16979 (N_16979,N_16134,N_16319);
nor U16980 (N_16980,N_16788,N_16288);
xor U16981 (N_16981,N_16604,N_16215);
nand U16982 (N_16982,N_16315,N_16586);
nor U16983 (N_16983,N_16010,N_16487);
and U16984 (N_16984,N_16700,N_16152);
xor U16985 (N_16985,N_16316,N_16337);
xnor U16986 (N_16986,N_16167,N_16690);
nand U16987 (N_16987,N_16754,N_16573);
and U16988 (N_16988,N_16756,N_16199);
xor U16989 (N_16989,N_16172,N_16558);
nor U16990 (N_16990,N_16226,N_16076);
xnor U16991 (N_16991,N_16646,N_16092);
and U16992 (N_16992,N_16071,N_16379);
or U16993 (N_16993,N_16523,N_16043);
nor U16994 (N_16994,N_16403,N_16154);
nor U16995 (N_16995,N_16549,N_16090);
or U16996 (N_16996,N_16737,N_16641);
nand U16997 (N_16997,N_16697,N_16357);
nor U16998 (N_16998,N_16507,N_16162);
or U16999 (N_16999,N_16294,N_16458);
nor U17000 (N_17000,N_16051,N_16059);
and U17001 (N_17001,N_16343,N_16601);
nor U17002 (N_17002,N_16354,N_16587);
nand U17003 (N_17003,N_16187,N_16326);
or U17004 (N_17004,N_16310,N_16262);
or U17005 (N_17005,N_16018,N_16506);
nand U17006 (N_17006,N_16312,N_16200);
and U17007 (N_17007,N_16671,N_16253);
nand U17008 (N_17008,N_16708,N_16164);
nor U17009 (N_17009,N_16157,N_16260);
nand U17010 (N_17010,N_16227,N_16038);
xnor U17011 (N_17011,N_16494,N_16658);
or U17012 (N_17012,N_16743,N_16732);
or U17013 (N_17013,N_16395,N_16273);
and U17014 (N_17014,N_16769,N_16464);
and U17015 (N_17015,N_16548,N_16192);
xnor U17016 (N_17016,N_16242,N_16706);
or U17017 (N_17017,N_16456,N_16377);
xor U17018 (N_17018,N_16538,N_16467);
xnor U17019 (N_17019,N_16340,N_16156);
xor U17020 (N_17020,N_16204,N_16661);
xnor U17021 (N_17021,N_16726,N_16774);
or U17022 (N_17022,N_16753,N_16786);
nor U17023 (N_17023,N_16020,N_16469);
and U17024 (N_17024,N_16206,N_16417);
or U17025 (N_17025,N_16211,N_16271);
or U17026 (N_17026,N_16623,N_16561);
nor U17027 (N_17027,N_16734,N_16066);
xor U17028 (N_17028,N_16111,N_16551);
nand U17029 (N_17029,N_16236,N_16659);
nand U17030 (N_17030,N_16281,N_16177);
and U17031 (N_17031,N_16676,N_16681);
and U17032 (N_17032,N_16525,N_16369);
nor U17033 (N_17033,N_16477,N_16371);
or U17034 (N_17034,N_16349,N_16263);
or U17035 (N_17035,N_16297,N_16696);
nor U17036 (N_17036,N_16257,N_16225);
nand U17037 (N_17037,N_16612,N_16213);
or U17038 (N_17038,N_16514,N_16025);
nor U17039 (N_17039,N_16772,N_16093);
xnor U17040 (N_17040,N_16629,N_16362);
nor U17041 (N_17041,N_16683,N_16041);
and U17042 (N_17042,N_16104,N_16474);
nand U17043 (N_17043,N_16725,N_16450);
or U17044 (N_17044,N_16375,N_16160);
nand U17045 (N_17045,N_16740,N_16205);
and U17046 (N_17046,N_16195,N_16251);
nor U17047 (N_17047,N_16466,N_16599);
xor U17048 (N_17048,N_16409,N_16562);
or U17049 (N_17049,N_16544,N_16543);
nand U17050 (N_17050,N_16266,N_16613);
or U17051 (N_17051,N_16492,N_16008);
xor U17052 (N_17052,N_16455,N_16611);
or U17053 (N_17053,N_16280,N_16483);
or U17054 (N_17054,N_16401,N_16219);
nor U17055 (N_17055,N_16232,N_16766);
or U17056 (N_17056,N_16224,N_16250);
nor U17057 (N_17057,N_16408,N_16636);
xnor U17058 (N_17058,N_16143,N_16593);
and U17059 (N_17059,N_16555,N_16498);
nand U17060 (N_17060,N_16509,N_16159);
nand U17061 (N_17061,N_16083,N_16396);
xnor U17062 (N_17062,N_16691,N_16515);
nand U17063 (N_17063,N_16254,N_16582);
xor U17064 (N_17064,N_16771,N_16779);
nor U17065 (N_17065,N_16412,N_16399);
or U17066 (N_17066,N_16217,N_16406);
xor U17067 (N_17067,N_16074,N_16308);
or U17068 (N_17068,N_16100,N_16021);
xnor U17069 (N_17069,N_16061,N_16155);
xnor U17070 (N_17070,N_16598,N_16524);
nand U17071 (N_17071,N_16099,N_16267);
and U17072 (N_17072,N_16130,N_16584);
xnor U17073 (N_17073,N_16550,N_16019);
nor U17074 (N_17074,N_16390,N_16358);
or U17075 (N_17075,N_16447,N_16238);
nand U17076 (N_17076,N_16602,N_16673);
nor U17077 (N_17077,N_16776,N_16438);
nand U17078 (N_17078,N_16166,N_16723);
nor U17079 (N_17079,N_16309,N_16075);
nor U17080 (N_17080,N_16301,N_16067);
and U17081 (N_17081,N_16745,N_16291);
and U17082 (N_17082,N_16116,N_16418);
and U17083 (N_17083,N_16283,N_16606);
xor U17084 (N_17084,N_16435,N_16482);
or U17085 (N_17085,N_16289,N_16617);
nor U17086 (N_17086,N_16368,N_16594);
nand U17087 (N_17087,N_16270,N_16616);
nand U17088 (N_17088,N_16210,N_16106);
nand U17089 (N_17089,N_16069,N_16245);
nor U17090 (N_17090,N_16345,N_16214);
nand U17091 (N_17091,N_16072,N_16591);
and U17092 (N_17092,N_16179,N_16035);
nand U17093 (N_17093,N_16385,N_16427);
nor U17094 (N_17094,N_16158,N_16693);
or U17095 (N_17095,N_16539,N_16688);
or U17096 (N_17096,N_16722,N_16073);
nor U17097 (N_17097,N_16702,N_16052);
nor U17098 (N_17098,N_16278,N_16462);
or U17099 (N_17099,N_16128,N_16529);
xor U17100 (N_17100,N_16781,N_16595);
xnor U17101 (N_17101,N_16508,N_16443);
nand U17102 (N_17102,N_16394,N_16568);
xor U17103 (N_17103,N_16328,N_16001);
and U17104 (N_17104,N_16625,N_16070);
nor U17105 (N_17105,N_16293,N_16351);
and U17106 (N_17106,N_16147,N_16760);
nand U17107 (N_17107,N_16175,N_16793);
and U17108 (N_17108,N_16746,N_16139);
xnor U17109 (N_17109,N_16118,N_16295);
and U17110 (N_17110,N_16120,N_16635);
or U17111 (N_17111,N_16764,N_16445);
nor U17112 (N_17112,N_16735,N_16657);
nor U17113 (N_17113,N_16193,N_16323);
nor U17114 (N_17114,N_16388,N_16258);
xor U17115 (N_17115,N_16630,N_16597);
nand U17116 (N_17116,N_16459,N_16048);
nand U17117 (N_17117,N_16228,N_16320);
and U17118 (N_17118,N_16799,N_16202);
or U17119 (N_17119,N_16274,N_16426);
nand U17120 (N_17120,N_16430,N_16149);
and U17121 (N_17121,N_16608,N_16180);
or U17122 (N_17122,N_16140,N_16751);
xnor U17123 (N_17123,N_16489,N_16460);
nand U17124 (N_17124,N_16461,N_16542);
nor U17125 (N_17125,N_16411,N_16579);
xnor U17126 (N_17126,N_16441,N_16570);
nor U17127 (N_17127,N_16421,N_16620);
xor U17128 (N_17128,N_16428,N_16485);
and U17129 (N_17129,N_16101,N_16015);
xnor U17130 (N_17130,N_16348,N_16081);
nand U17131 (N_17131,N_16797,N_16185);
or U17132 (N_17132,N_16338,N_16669);
xor U17133 (N_17133,N_16567,N_16780);
xnor U17134 (N_17134,N_16146,N_16575);
and U17135 (N_17135,N_16656,N_16347);
and U17136 (N_17136,N_16373,N_16234);
or U17137 (N_17137,N_16728,N_16721);
and U17138 (N_17138,N_16058,N_16666);
or U17139 (N_17139,N_16634,N_16364);
xnor U17140 (N_17140,N_16632,N_16121);
nor U17141 (N_17141,N_16161,N_16705);
nor U17142 (N_17142,N_16303,N_16321);
nand U17143 (N_17143,N_16750,N_16404);
xor U17144 (N_17144,N_16554,N_16727);
nor U17145 (N_17145,N_16040,N_16605);
or U17146 (N_17146,N_16252,N_16109);
nand U17147 (N_17147,N_16305,N_16125);
and U17148 (N_17148,N_16325,N_16203);
or U17149 (N_17149,N_16615,N_16698);
xor U17150 (N_17150,N_16314,N_16511);
nand U17151 (N_17151,N_16207,N_16286);
and U17152 (N_17152,N_16556,N_16261);
xnor U17153 (N_17153,N_16479,N_16667);
nand U17154 (N_17154,N_16078,N_16648);
nor U17155 (N_17155,N_16685,N_16393);
or U17156 (N_17156,N_16637,N_16420);
and U17157 (N_17157,N_16493,N_16363);
and U17158 (N_17158,N_16471,N_16546);
nor U17159 (N_17159,N_16218,N_16117);
and U17160 (N_17160,N_16663,N_16248);
and U17161 (N_17161,N_16088,N_16003);
xnor U17162 (N_17162,N_16091,N_16239);
and U17163 (N_17163,N_16322,N_16429);
xnor U17164 (N_17164,N_16132,N_16713);
nor U17165 (N_17165,N_16590,N_16178);
nor U17166 (N_17166,N_16738,N_16096);
and U17167 (N_17167,N_16440,N_16639);
xnor U17168 (N_17168,N_16473,N_16150);
nand U17169 (N_17169,N_16571,N_16709);
xnor U17170 (N_17170,N_16767,N_16287);
or U17171 (N_17171,N_16011,N_16765);
nor U17172 (N_17172,N_16405,N_16531);
nand U17173 (N_17173,N_16148,N_16062);
xor U17174 (N_17174,N_16046,N_16436);
nand U17175 (N_17175,N_16415,N_16478);
nand U17176 (N_17176,N_16233,N_16318);
and U17177 (N_17177,N_16014,N_16622);
and U17178 (N_17178,N_16647,N_16718);
nand U17179 (N_17179,N_16355,N_16527);
xor U17180 (N_17180,N_16510,N_16433);
or U17181 (N_17181,N_16381,N_16196);
and U17182 (N_17182,N_16327,N_16502);
nand U17183 (N_17183,N_16491,N_16367);
and U17184 (N_17184,N_16400,N_16317);
and U17185 (N_17185,N_16216,N_16005);
xor U17186 (N_17186,N_16163,N_16264);
and U17187 (N_17187,N_16495,N_16170);
or U17188 (N_17188,N_16144,N_16277);
nor U17189 (N_17189,N_16246,N_16684);
nand U17190 (N_17190,N_16085,N_16209);
nand U17191 (N_17191,N_16336,N_16468);
nand U17192 (N_17192,N_16053,N_16060);
or U17193 (N_17193,N_16137,N_16564);
and U17194 (N_17194,N_16704,N_16151);
xor U17195 (N_17195,N_16782,N_16644);
and U17196 (N_17196,N_16102,N_16079);
xnor U17197 (N_17197,N_16536,N_16352);
nor U17198 (N_17198,N_16341,N_16741);
nor U17199 (N_17199,N_16017,N_16296);
xor U17200 (N_17200,N_16508,N_16147);
nor U17201 (N_17201,N_16173,N_16445);
xnor U17202 (N_17202,N_16138,N_16002);
xor U17203 (N_17203,N_16600,N_16314);
nor U17204 (N_17204,N_16229,N_16304);
xor U17205 (N_17205,N_16397,N_16410);
and U17206 (N_17206,N_16411,N_16185);
nand U17207 (N_17207,N_16348,N_16675);
nand U17208 (N_17208,N_16048,N_16617);
and U17209 (N_17209,N_16787,N_16380);
and U17210 (N_17210,N_16730,N_16416);
nand U17211 (N_17211,N_16166,N_16208);
and U17212 (N_17212,N_16635,N_16370);
nor U17213 (N_17213,N_16460,N_16677);
or U17214 (N_17214,N_16252,N_16349);
nor U17215 (N_17215,N_16500,N_16056);
and U17216 (N_17216,N_16788,N_16536);
nand U17217 (N_17217,N_16234,N_16301);
xor U17218 (N_17218,N_16106,N_16741);
nand U17219 (N_17219,N_16737,N_16006);
nor U17220 (N_17220,N_16406,N_16707);
nand U17221 (N_17221,N_16564,N_16757);
xnor U17222 (N_17222,N_16521,N_16201);
xor U17223 (N_17223,N_16275,N_16047);
nor U17224 (N_17224,N_16672,N_16484);
nand U17225 (N_17225,N_16272,N_16337);
nand U17226 (N_17226,N_16238,N_16589);
xor U17227 (N_17227,N_16427,N_16215);
nand U17228 (N_17228,N_16220,N_16709);
and U17229 (N_17229,N_16525,N_16290);
or U17230 (N_17230,N_16055,N_16697);
and U17231 (N_17231,N_16628,N_16793);
nand U17232 (N_17232,N_16723,N_16255);
or U17233 (N_17233,N_16197,N_16265);
nand U17234 (N_17234,N_16642,N_16143);
and U17235 (N_17235,N_16317,N_16330);
nand U17236 (N_17236,N_16224,N_16657);
and U17237 (N_17237,N_16619,N_16424);
or U17238 (N_17238,N_16009,N_16504);
xor U17239 (N_17239,N_16289,N_16416);
and U17240 (N_17240,N_16445,N_16681);
nand U17241 (N_17241,N_16741,N_16007);
and U17242 (N_17242,N_16665,N_16401);
nand U17243 (N_17243,N_16541,N_16518);
nor U17244 (N_17244,N_16697,N_16138);
nor U17245 (N_17245,N_16252,N_16455);
or U17246 (N_17246,N_16384,N_16449);
and U17247 (N_17247,N_16482,N_16216);
or U17248 (N_17248,N_16557,N_16153);
and U17249 (N_17249,N_16336,N_16478);
nor U17250 (N_17250,N_16066,N_16546);
or U17251 (N_17251,N_16680,N_16516);
and U17252 (N_17252,N_16410,N_16361);
xor U17253 (N_17253,N_16774,N_16510);
and U17254 (N_17254,N_16575,N_16034);
nor U17255 (N_17255,N_16045,N_16756);
nand U17256 (N_17256,N_16718,N_16799);
nand U17257 (N_17257,N_16112,N_16167);
or U17258 (N_17258,N_16035,N_16055);
and U17259 (N_17259,N_16503,N_16164);
nand U17260 (N_17260,N_16332,N_16365);
or U17261 (N_17261,N_16150,N_16013);
nand U17262 (N_17262,N_16135,N_16174);
and U17263 (N_17263,N_16188,N_16513);
nand U17264 (N_17264,N_16425,N_16397);
xnor U17265 (N_17265,N_16362,N_16373);
and U17266 (N_17266,N_16063,N_16024);
nand U17267 (N_17267,N_16368,N_16058);
or U17268 (N_17268,N_16120,N_16215);
nand U17269 (N_17269,N_16288,N_16025);
nand U17270 (N_17270,N_16493,N_16550);
xnor U17271 (N_17271,N_16272,N_16305);
and U17272 (N_17272,N_16124,N_16649);
or U17273 (N_17273,N_16331,N_16495);
or U17274 (N_17274,N_16027,N_16206);
nor U17275 (N_17275,N_16785,N_16097);
xnor U17276 (N_17276,N_16604,N_16357);
and U17277 (N_17277,N_16558,N_16749);
and U17278 (N_17278,N_16197,N_16565);
xor U17279 (N_17279,N_16414,N_16088);
or U17280 (N_17280,N_16402,N_16583);
and U17281 (N_17281,N_16025,N_16601);
or U17282 (N_17282,N_16365,N_16488);
xnor U17283 (N_17283,N_16337,N_16195);
nor U17284 (N_17284,N_16769,N_16520);
nand U17285 (N_17285,N_16013,N_16529);
and U17286 (N_17286,N_16162,N_16336);
and U17287 (N_17287,N_16546,N_16650);
and U17288 (N_17288,N_16131,N_16572);
or U17289 (N_17289,N_16008,N_16379);
or U17290 (N_17290,N_16634,N_16599);
or U17291 (N_17291,N_16761,N_16762);
xor U17292 (N_17292,N_16407,N_16536);
xnor U17293 (N_17293,N_16443,N_16346);
or U17294 (N_17294,N_16407,N_16726);
nor U17295 (N_17295,N_16186,N_16115);
xor U17296 (N_17296,N_16513,N_16065);
nor U17297 (N_17297,N_16778,N_16403);
nor U17298 (N_17298,N_16473,N_16240);
nor U17299 (N_17299,N_16411,N_16205);
or U17300 (N_17300,N_16166,N_16337);
or U17301 (N_17301,N_16010,N_16146);
nor U17302 (N_17302,N_16799,N_16354);
xor U17303 (N_17303,N_16076,N_16073);
nand U17304 (N_17304,N_16619,N_16615);
and U17305 (N_17305,N_16700,N_16008);
nand U17306 (N_17306,N_16372,N_16018);
xor U17307 (N_17307,N_16401,N_16126);
nand U17308 (N_17308,N_16183,N_16276);
nand U17309 (N_17309,N_16375,N_16303);
and U17310 (N_17310,N_16370,N_16744);
nor U17311 (N_17311,N_16459,N_16303);
or U17312 (N_17312,N_16518,N_16748);
xnor U17313 (N_17313,N_16047,N_16196);
nor U17314 (N_17314,N_16053,N_16609);
xnor U17315 (N_17315,N_16426,N_16661);
or U17316 (N_17316,N_16771,N_16524);
nand U17317 (N_17317,N_16206,N_16677);
or U17318 (N_17318,N_16596,N_16313);
xor U17319 (N_17319,N_16412,N_16034);
nand U17320 (N_17320,N_16483,N_16406);
xor U17321 (N_17321,N_16593,N_16320);
nor U17322 (N_17322,N_16353,N_16597);
xnor U17323 (N_17323,N_16286,N_16188);
and U17324 (N_17324,N_16564,N_16760);
or U17325 (N_17325,N_16402,N_16030);
nand U17326 (N_17326,N_16535,N_16064);
nor U17327 (N_17327,N_16773,N_16244);
or U17328 (N_17328,N_16474,N_16223);
nand U17329 (N_17329,N_16003,N_16441);
and U17330 (N_17330,N_16773,N_16022);
and U17331 (N_17331,N_16051,N_16505);
and U17332 (N_17332,N_16713,N_16304);
nand U17333 (N_17333,N_16719,N_16262);
nand U17334 (N_17334,N_16338,N_16058);
nor U17335 (N_17335,N_16768,N_16533);
or U17336 (N_17336,N_16459,N_16003);
nor U17337 (N_17337,N_16600,N_16755);
nand U17338 (N_17338,N_16024,N_16069);
xnor U17339 (N_17339,N_16186,N_16131);
nand U17340 (N_17340,N_16381,N_16586);
and U17341 (N_17341,N_16151,N_16405);
xor U17342 (N_17342,N_16675,N_16713);
or U17343 (N_17343,N_16742,N_16785);
xor U17344 (N_17344,N_16186,N_16409);
nand U17345 (N_17345,N_16316,N_16032);
xor U17346 (N_17346,N_16502,N_16018);
xnor U17347 (N_17347,N_16079,N_16607);
nand U17348 (N_17348,N_16415,N_16020);
nor U17349 (N_17349,N_16277,N_16426);
nand U17350 (N_17350,N_16686,N_16084);
or U17351 (N_17351,N_16643,N_16500);
xnor U17352 (N_17352,N_16045,N_16090);
xor U17353 (N_17353,N_16155,N_16476);
nor U17354 (N_17354,N_16197,N_16404);
nor U17355 (N_17355,N_16442,N_16757);
nand U17356 (N_17356,N_16443,N_16608);
nor U17357 (N_17357,N_16376,N_16214);
xnor U17358 (N_17358,N_16756,N_16164);
or U17359 (N_17359,N_16696,N_16281);
and U17360 (N_17360,N_16077,N_16763);
xnor U17361 (N_17361,N_16235,N_16373);
xnor U17362 (N_17362,N_16071,N_16446);
or U17363 (N_17363,N_16781,N_16332);
nor U17364 (N_17364,N_16218,N_16061);
nor U17365 (N_17365,N_16289,N_16010);
nor U17366 (N_17366,N_16654,N_16614);
or U17367 (N_17367,N_16404,N_16355);
or U17368 (N_17368,N_16761,N_16292);
or U17369 (N_17369,N_16417,N_16370);
nand U17370 (N_17370,N_16217,N_16070);
and U17371 (N_17371,N_16091,N_16701);
and U17372 (N_17372,N_16717,N_16592);
nor U17373 (N_17373,N_16571,N_16386);
nand U17374 (N_17374,N_16313,N_16022);
xor U17375 (N_17375,N_16356,N_16067);
nand U17376 (N_17376,N_16055,N_16247);
or U17377 (N_17377,N_16135,N_16662);
and U17378 (N_17378,N_16056,N_16685);
xnor U17379 (N_17379,N_16032,N_16772);
or U17380 (N_17380,N_16571,N_16012);
nor U17381 (N_17381,N_16606,N_16591);
and U17382 (N_17382,N_16717,N_16326);
nor U17383 (N_17383,N_16069,N_16708);
nor U17384 (N_17384,N_16485,N_16296);
or U17385 (N_17385,N_16506,N_16588);
nand U17386 (N_17386,N_16732,N_16266);
nor U17387 (N_17387,N_16105,N_16301);
and U17388 (N_17388,N_16503,N_16286);
xnor U17389 (N_17389,N_16532,N_16046);
nor U17390 (N_17390,N_16782,N_16247);
xor U17391 (N_17391,N_16124,N_16161);
nand U17392 (N_17392,N_16482,N_16334);
nor U17393 (N_17393,N_16079,N_16470);
and U17394 (N_17394,N_16759,N_16654);
nand U17395 (N_17395,N_16518,N_16789);
or U17396 (N_17396,N_16698,N_16302);
or U17397 (N_17397,N_16566,N_16568);
or U17398 (N_17398,N_16029,N_16319);
and U17399 (N_17399,N_16657,N_16160);
nand U17400 (N_17400,N_16208,N_16170);
and U17401 (N_17401,N_16319,N_16228);
or U17402 (N_17402,N_16698,N_16183);
nor U17403 (N_17403,N_16513,N_16647);
or U17404 (N_17404,N_16483,N_16645);
nor U17405 (N_17405,N_16651,N_16285);
or U17406 (N_17406,N_16343,N_16365);
nor U17407 (N_17407,N_16680,N_16648);
nor U17408 (N_17408,N_16038,N_16073);
xnor U17409 (N_17409,N_16209,N_16049);
and U17410 (N_17410,N_16787,N_16333);
xor U17411 (N_17411,N_16716,N_16339);
or U17412 (N_17412,N_16731,N_16192);
xnor U17413 (N_17413,N_16273,N_16778);
and U17414 (N_17414,N_16607,N_16100);
nor U17415 (N_17415,N_16361,N_16294);
or U17416 (N_17416,N_16788,N_16527);
nand U17417 (N_17417,N_16470,N_16393);
xor U17418 (N_17418,N_16734,N_16080);
or U17419 (N_17419,N_16728,N_16576);
and U17420 (N_17420,N_16536,N_16730);
nand U17421 (N_17421,N_16352,N_16219);
or U17422 (N_17422,N_16507,N_16240);
or U17423 (N_17423,N_16431,N_16282);
or U17424 (N_17424,N_16742,N_16284);
nor U17425 (N_17425,N_16371,N_16073);
nor U17426 (N_17426,N_16559,N_16242);
nand U17427 (N_17427,N_16588,N_16415);
or U17428 (N_17428,N_16528,N_16534);
xnor U17429 (N_17429,N_16672,N_16322);
nand U17430 (N_17430,N_16050,N_16321);
nor U17431 (N_17431,N_16056,N_16462);
nor U17432 (N_17432,N_16744,N_16671);
nand U17433 (N_17433,N_16395,N_16645);
or U17434 (N_17434,N_16669,N_16180);
nor U17435 (N_17435,N_16442,N_16302);
nor U17436 (N_17436,N_16127,N_16691);
xnor U17437 (N_17437,N_16549,N_16582);
and U17438 (N_17438,N_16775,N_16164);
or U17439 (N_17439,N_16339,N_16080);
nand U17440 (N_17440,N_16786,N_16383);
nor U17441 (N_17441,N_16246,N_16177);
xor U17442 (N_17442,N_16082,N_16253);
and U17443 (N_17443,N_16145,N_16296);
or U17444 (N_17444,N_16506,N_16301);
nand U17445 (N_17445,N_16435,N_16609);
nor U17446 (N_17446,N_16583,N_16447);
nand U17447 (N_17447,N_16591,N_16790);
or U17448 (N_17448,N_16769,N_16693);
xor U17449 (N_17449,N_16112,N_16269);
nand U17450 (N_17450,N_16123,N_16413);
nor U17451 (N_17451,N_16167,N_16625);
xor U17452 (N_17452,N_16479,N_16642);
nor U17453 (N_17453,N_16587,N_16267);
or U17454 (N_17454,N_16790,N_16033);
or U17455 (N_17455,N_16439,N_16173);
or U17456 (N_17456,N_16049,N_16303);
nand U17457 (N_17457,N_16213,N_16264);
or U17458 (N_17458,N_16201,N_16560);
and U17459 (N_17459,N_16261,N_16060);
or U17460 (N_17460,N_16370,N_16630);
nor U17461 (N_17461,N_16019,N_16246);
xor U17462 (N_17462,N_16602,N_16274);
or U17463 (N_17463,N_16345,N_16775);
nor U17464 (N_17464,N_16281,N_16662);
and U17465 (N_17465,N_16432,N_16719);
and U17466 (N_17466,N_16171,N_16479);
or U17467 (N_17467,N_16349,N_16311);
and U17468 (N_17468,N_16046,N_16371);
xnor U17469 (N_17469,N_16782,N_16449);
nand U17470 (N_17470,N_16491,N_16259);
nand U17471 (N_17471,N_16294,N_16031);
nor U17472 (N_17472,N_16200,N_16628);
nand U17473 (N_17473,N_16472,N_16208);
xnor U17474 (N_17474,N_16285,N_16477);
and U17475 (N_17475,N_16206,N_16534);
or U17476 (N_17476,N_16110,N_16653);
xnor U17477 (N_17477,N_16072,N_16701);
nand U17478 (N_17478,N_16264,N_16066);
nand U17479 (N_17479,N_16478,N_16094);
nand U17480 (N_17480,N_16132,N_16454);
nand U17481 (N_17481,N_16026,N_16207);
or U17482 (N_17482,N_16666,N_16501);
nand U17483 (N_17483,N_16206,N_16096);
xor U17484 (N_17484,N_16192,N_16264);
nor U17485 (N_17485,N_16568,N_16037);
nor U17486 (N_17486,N_16227,N_16546);
and U17487 (N_17487,N_16742,N_16563);
nor U17488 (N_17488,N_16607,N_16394);
xnor U17489 (N_17489,N_16579,N_16590);
nand U17490 (N_17490,N_16359,N_16246);
and U17491 (N_17491,N_16173,N_16139);
xor U17492 (N_17492,N_16071,N_16043);
and U17493 (N_17493,N_16638,N_16721);
xnor U17494 (N_17494,N_16264,N_16039);
nand U17495 (N_17495,N_16699,N_16288);
nand U17496 (N_17496,N_16099,N_16191);
nand U17497 (N_17497,N_16017,N_16222);
or U17498 (N_17498,N_16780,N_16758);
nand U17499 (N_17499,N_16127,N_16432);
and U17500 (N_17500,N_16426,N_16015);
and U17501 (N_17501,N_16341,N_16192);
xor U17502 (N_17502,N_16264,N_16286);
nor U17503 (N_17503,N_16264,N_16540);
xor U17504 (N_17504,N_16541,N_16453);
or U17505 (N_17505,N_16665,N_16555);
nand U17506 (N_17506,N_16661,N_16377);
xor U17507 (N_17507,N_16115,N_16497);
xor U17508 (N_17508,N_16783,N_16433);
xnor U17509 (N_17509,N_16574,N_16419);
nor U17510 (N_17510,N_16426,N_16764);
or U17511 (N_17511,N_16553,N_16368);
xor U17512 (N_17512,N_16602,N_16183);
xnor U17513 (N_17513,N_16761,N_16164);
or U17514 (N_17514,N_16631,N_16357);
nor U17515 (N_17515,N_16182,N_16239);
and U17516 (N_17516,N_16518,N_16238);
and U17517 (N_17517,N_16143,N_16146);
and U17518 (N_17518,N_16429,N_16518);
and U17519 (N_17519,N_16011,N_16141);
nor U17520 (N_17520,N_16605,N_16175);
xnor U17521 (N_17521,N_16285,N_16652);
nand U17522 (N_17522,N_16546,N_16004);
nand U17523 (N_17523,N_16382,N_16402);
nor U17524 (N_17524,N_16695,N_16614);
nor U17525 (N_17525,N_16099,N_16159);
nor U17526 (N_17526,N_16228,N_16779);
and U17527 (N_17527,N_16089,N_16161);
and U17528 (N_17528,N_16258,N_16053);
or U17529 (N_17529,N_16182,N_16716);
xnor U17530 (N_17530,N_16187,N_16646);
nor U17531 (N_17531,N_16262,N_16489);
nand U17532 (N_17532,N_16581,N_16268);
or U17533 (N_17533,N_16074,N_16697);
nand U17534 (N_17534,N_16334,N_16232);
nand U17535 (N_17535,N_16395,N_16576);
xnor U17536 (N_17536,N_16192,N_16559);
or U17537 (N_17537,N_16533,N_16753);
nor U17538 (N_17538,N_16581,N_16064);
or U17539 (N_17539,N_16505,N_16172);
and U17540 (N_17540,N_16095,N_16746);
nand U17541 (N_17541,N_16388,N_16453);
or U17542 (N_17542,N_16748,N_16282);
nand U17543 (N_17543,N_16007,N_16720);
nor U17544 (N_17544,N_16746,N_16394);
nand U17545 (N_17545,N_16432,N_16057);
nand U17546 (N_17546,N_16439,N_16518);
or U17547 (N_17547,N_16496,N_16438);
nor U17548 (N_17548,N_16691,N_16251);
xnor U17549 (N_17549,N_16304,N_16249);
or U17550 (N_17550,N_16271,N_16740);
xor U17551 (N_17551,N_16139,N_16213);
nand U17552 (N_17552,N_16716,N_16347);
xor U17553 (N_17553,N_16242,N_16684);
or U17554 (N_17554,N_16057,N_16079);
or U17555 (N_17555,N_16346,N_16630);
nand U17556 (N_17556,N_16459,N_16703);
nand U17557 (N_17557,N_16435,N_16094);
nand U17558 (N_17558,N_16007,N_16452);
and U17559 (N_17559,N_16688,N_16434);
or U17560 (N_17560,N_16120,N_16071);
and U17561 (N_17561,N_16385,N_16744);
and U17562 (N_17562,N_16464,N_16288);
and U17563 (N_17563,N_16732,N_16788);
nand U17564 (N_17564,N_16371,N_16695);
or U17565 (N_17565,N_16001,N_16756);
nor U17566 (N_17566,N_16251,N_16597);
and U17567 (N_17567,N_16166,N_16331);
nand U17568 (N_17568,N_16187,N_16250);
or U17569 (N_17569,N_16199,N_16637);
nand U17570 (N_17570,N_16227,N_16273);
nand U17571 (N_17571,N_16465,N_16144);
nand U17572 (N_17572,N_16705,N_16234);
or U17573 (N_17573,N_16412,N_16014);
nand U17574 (N_17574,N_16258,N_16456);
nor U17575 (N_17575,N_16544,N_16488);
nand U17576 (N_17576,N_16692,N_16297);
xor U17577 (N_17577,N_16762,N_16011);
xor U17578 (N_17578,N_16088,N_16551);
nand U17579 (N_17579,N_16309,N_16462);
and U17580 (N_17580,N_16479,N_16145);
and U17581 (N_17581,N_16107,N_16740);
xor U17582 (N_17582,N_16708,N_16476);
nand U17583 (N_17583,N_16447,N_16349);
xor U17584 (N_17584,N_16630,N_16222);
nand U17585 (N_17585,N_16167,N_16700);
or U17586 (N_17586,N_16439,N_16433);
or U17587 (N_17587,N_16345,N_16425);
and U17588 (N_17588,N_16315,N_16398);
nand U17589 (N_17589,N_16176,N_16359);
xnor U17590 (N_17590,N_16145,N_16511);
and U17591 (N_17591,N_16039,N_16792);
nand U17592 (N_17592,N_16276,N_16265);
nor U17593 (N_17593,N_16793,N_16134);
xor U17594 (N_17594,N_16776,N_16593);
xor U17595 (N_17595,N_16664,N_16387);
nand U17596 (N_17596,N_16076,N_16272);
and U17597 (N_17597,N_16765,N_16120);
nor U17598 (N_17598,N_16565,N_16542);
nand U17599 (N_17599,N_16406,N_16360);
xor U17600 (N_17600,N_17188,N_17005);
nor U17601 (N_17601,N_17305,N_17329);
xor U17602 (N_17602,N_17094,N_16945);
nand U17603 (N_17603,N_17025,N_16916);
or U17604 (N_17604,N_16851,N_17560);
xnor U17605 (N_17605,N_17473,N_16841);
nor U17606 (N_17606,N_17171,N_17032);
and U17607 (N_17607,N_17562,N_16939);
or U17608 (N_17608,N_17599,N_17300);
or U17609 (N_17609,N_17090,N_17549);
and U17610 (N_17610,N_17585,N_17304);
nand U17611 (N_17611,N_17565,N_17347);
nand U17612 (N_17612,N_17014,N_16927);
nor U17613 (N_17613,N_17244,N_17384);
nand U17614 (N_17614,N_17538,N_16863);
nor U17615 (N_17615,N_16985,N_16872);
xnor U17616 (N_17616,N_17264,N_16980);
xor U17617 (N_17617,N_16955,N_17481);
xor U17618 (N_17618,N_17543,N_16970);
nand U17619 (N_17619,N_16990,N_17580);
nor U17620 (N_17620,N_17409,N_17480);
or U17621 (N_17621,N_17333,N_16887);
xnor U17622 (N_17622,N_17542,N_17371);
nor U17623 (N_17623,N_17143,N_17404);
nor U17624 (N_17624,N_17126,N_17127);
and U17625 (N_17625,N_17460,N_17551);
nand U17626 (N_17626,N_16906,N_17085);
or U17627 (N_17627,N_17177,N_17363);
xor U17628 (N_17628,N_17556,N_17167);
and U17629 (N_17629,N_17285,N_17295);
nand U17630 (N_17630,N_17309,N_17525);
and U17631 (N_17631,N_17112,N_16960);
nor U17632 (N_17632,N_17492,N_16921);
nand U17633 (N_17633,N_17572,N_16836);
nor U17634 (N_17634,N_17140,N_16884);
or U17635 (N_17635,N_17507,N_17176);
or U17636 (N_17636,N_17559,N_17401);
nor U17637 (N_17637,N_17458,N_17071);
and U17638 (N_17638,N_17487,N_17399);
xor U17639 (N_17639,N_17569,N_17060);
nand U17640 (N_17640,N_16837,N_17125);
and U17641 (N_17641,N_17446,N_17164);
xor U17642 (N_17642,N_17430,N_17061);
or U17643 (N_17643,N_16840,N_17272);
or U17644 (N_17644,N_16901,N_17489);
or U17645 (N_17645,N_16997,N_17465);
nor U17646 (N_17646,N_16956,N_17021);
and U17647 (N_17647,N_17199,N_17247);
nor U17648 (N_17648,N_17198,N_17332);
nor U17649 (N_17649,N_17224,N_17522);
nor U17650 (N_17650,N_17320,N_16821);
nand U17651 (N_17651,N_17200,N_16994);
and U17652 (N_17652,N_16914,N_16880);
or U17653 (N_17653,N_17083,N_16822);
nand U17654 (N_17654,N_17476,N_17312);
xor U17655 (N_17655,N_16833,N_17318);
and U17656 (N_17656,N_16874,N_17292);
and U17657 (N_17657,N_17521,N_17158);
xnor U17658 (N_17658,N_17201,N_16920);
nor U17659 (N_17659,N_17119,N_17575);
nor U17660 (N_17660,N_16852,N_17087);
or U17661 (N_17661,N_17019,N_17456);
nor U17662 (N_17662,N_17075,N_17053);
nand U17663 (N_17663,N_16926,N_17432);
and U17664 (N_17664,N_17478,N_17524);
nand U17665 (N_17665,N_16907,N_17540);
nand U17666 (N_17666,N_17408,N_17105);
xor U17667 (N_17667,N_17269,N_17110);
or U17668 (N_17668,N_17392,N_16802);
and U17669 (N_17669,N_17003,N_17386);
or U17670 (N_17670,N_17541,N_16832);
and U17671 (N_17671,N_16811,N_16891);
or U17672 (N_17672,N_17115,N_17102);
nand U17673 (N_17673,N_16868,N_17275);
or U17674 (N_17674,N_17331,N_17120);
and U17675 (N_17675,N_16886,N_17076);
xor U17676 (N_17676,N_17360,N_17280);
and U17677 (N_17677,N_17364,N_17470);
nand U17678 (N_17678,N_16904,N_17000);
and U17679 (N_17679,N_17203,N_17302);
nor U17680 (N_17680,N_17374,N_17426);
nand U17681 (N_17681,N_16900,N_16856);
nor U17682 (N_17682,N_17548,N_17172);
nor U17683 (N_17683,N_17040,N_17231);
nand U17684 (N_17684,N_16995,N_16842);
nor U17685 (N_17685,N_17001,N_17131);
xor U17686 (N_17686,N_17425,N_16919);
and U17687 (N_17687,N_17013,N_16831);
xor U17688 (N_17688,N_17051,N_17505);
nor U17689 (N_17689,N_17175,N_17375);
xnor U17690 (N_17690,N_16959,N_16845);
and U17691 (N_17691,N_16964,N_16846);
nor U17692 (N_17692,N_17469,N_17531);
nor U17693 (N_17693,N_17528,N_17322);
or U17694 (N_17694,N_17437,N_17064);
nor U17695 (N_17695,N_17191,N_17070);
and U17696 (N_17696,N_17148,N_17424);
nor U17697 (N_17697,N_17293,N_17045);
xnor U17698 (N_17698,N_16853,N_17555);
nand U17699 (N_17699,N_17475,N_17445);
nor U17700 (N_17700,N_17439,N_17156);
xnor U17701 (N_17701,N_17163,N_17537);
xor U17702 (N_17702,N_17552,N_17587);
and U17703 (N_17703,N_17510,N_17114);
and U17704 (N_17704,N_17296,N_17518);
nor U17705 (N_17705,N_17563,N_17017);
nor U17706 (N_17706,N_17162,N_17454);
nor U17707 (N_17707,N_17576,N_16915);
xor U17708 (N_17708,N_16977,N_17218);
xnor U17709 (N_17709,N_17297,N_17340);
or U17710 (N_17710,N_16930,N_17205);
nand U17711 (N_17711,N_16988,N_17253);
or U17712 (N_17712,N_16950,N_17095);
nor U17713 (N_17713,N_17036,N_16905);
and U17714 (N_17714,N_17078,N_17289);
xor U17715 (N_17715,N_17351,N_16946);
nor U17716 (N_17716,N_17009,N_17453);
and U17717 (N_17717,N_16992,N_16911);
nand U17718 (N_17718,N_17341,N_16944);
xnor U17719 (N_17719,N_17093,N_17417);
or U17720 (N_17720,N_16864,N_17274);
and U17721 (N_17721,N_17512,N_16806);
or U17722 (N_17722,N_17225,N_17260);
nor U17723 (N_17723,N_16897,N_17135);
or U17724 (N_17724,N_17179,N_16825);
and U17725 (N_17725,N_17091,N_17104);
and U17726 (N_17726,N_16932,N_17596);
nor U17727 (N_17727,N_16962,N_17582);
nor U17728 (N_17728,N_16839,N_16935);
xnor U17729 (N_17729,N_16877,N_16876);
or U17730 (N_17730,N_17588,N_17245);
nor U17731 (N_17731,N_17506,N_16892);
nor U17732 (N_17732,N_16871,N_17306);
nor U17733 (N_17733,N_17282,N_17546);
nand U17734 (N_17734,N_17496,N_16898);
xnor U17735 (N_17735,N_17369,N_17405);
nor U17736 (N_17736,N_16986,N_17002);
nor U17737 (N_17737,N_16865,N_17240);
nand U17738 (N_17738,N_17228,N_17047);
and U17739 (N_17739,N_17373,N_16800);
and U17740 (N_17740,N_17035,N_17290);
nor U17741 (N_17741,N_16918,N_17170);
or U17742 (N_17742,N_17130,N_17311);
nand U17743 (N_17743,N_16993,N_17137);
nand U17744 (N_17744,N_17438,N_17041);
and U17745 (N_17745,N_17486,N_17049);
nand U17746 (N_17746,N_16807,N_17361);
and U17747 (N_17747,N_16834,N_17334);
or U17748 (N_17748,N_16828,N_17145);
and U17749 (N_17749,N_16870,N_16931);
or U17750 (N_17750,N_16817,N_17026);
nand U17751 (N_17751,N_16879,N_17080);
nand U17752 (N_17752,N_17046,N_17239);
nand U17753 (N_17753,N_17097,N_17536);
and U17754 (N_17754,N_17284,N_17086);
or U17755 (N_17755,N_16913,N_17263);
or U17756 (N_17756,N_17122,N_16835);
or U17757 (N_17757,N_17431,N_17197);
xor U17758 (N_17758,N_17410,N_17023);
xor U17759 (N_17759,N_16829,N_17419);
xnor U17760 (N_17760,N_17464,N_17220);
xnor U17761 (N_17761,N_16860,N_17301);
or U17762 (N_17762,N_16896,N_17299);
xnor U17763 (N_17763,N_16849,N_17324);
nand U17764 (N_17764,N_17435,N_17307);
xnor U17765 (N_17765,N_17389,N_17367);
or U17766 (N_17766,N_17564,N_16973);
and U17767 (N_17767,N_16801,N_17457);
and U17768 (N_17768,N_17252,N_17530);
and U17769 (N_17769,N_17113,N_17072);
nor U17770 (N_17770,N_17493,N_17268);
or U17771 (N_17771,N_16869,N_17008);
nand U17772 (N_17772,N_17088,N_17511);
and U17773 (N_17773,N_17497,N_17448);
nor U17774 (N_17774,N_17236,N_17461);
and U17775 (N_17775,N_16953,N_17433);
xor U17776 (N_17776,N_17366,N_17149);
or U17777 (N_17777,N_17586,N_17472);
nand U17778 (N_17778,N_17501,N_16978);
nand U17779 (N_17779,N_17362,N_16982);
and U17780 (N_17780,N_17420,N_17593);
nand U17781 (N_17781,N_17339,N_17578);
or U17782 (N_17782,N_17474,N_17273);
xor U17783 (N_17783,N_16971,N_17165);
or U17784 (N_17784,N_17434,N_17037);
and U17785 (N_17785,N_17223,N_17451);
nor U17786 (N_17786,N_17527,N_17050);
and U17787 (N_17787,N_17056,N_17281);
xor U17788 (N_17788,N_17106,N_17155);
xnor U17789 (N_17789,N_17012,N_17081);
nor U17790 (N_17790,N_16951,N_16908);
or U17791 (N_17791,N_17517,N_17313);
xnor U17792 (N_17792,N_17338,N_17452);
nor U17793 (N_17793,N_17421,N_17108);
nor U17794 (N_17794,N_17258,N_17234);
xnor U17795 (N_17795,N_17319,N_16808);
nor U17796 (N_17796,N_16968,N_16844);
xnor U17797 (N_17797,N_17406,N_16889);
nand U17798 (N_17798,N_17230,N_17010);
or U17799 (N_17799,N_17365,N_17411);
and U17800 (N_17800,N_17128,N_16940);
nor U17801 (N_17801,N_17479,N_16882);
or U17802 (N_17802,N_17388,N_17566);
nand U17803 (N_17803,N_17412,N_16983);
xor U17804 (N_17804,N_17346,N_17063);
and U17805 (N_17805,N_17504,N_17467);
or U17806 (N_17806,N_17229,N_17018);
xor U17807 (N_17807,N_17132,N_17092);
xnor U17808 (N_17808,N_16873,N_16899);
or U17809 (N_17809,N_17160,N_17317);
or U17810 (N_17810,N_17577,N_17502);
nand U17811 (N_17811,N_17583,N_16969);
and U17812 (N_17812,N_17161,N_17573);
nand U17813 (N_17813,N_17382,N_17429);
and U17814 (N_17814,N_17571,N_16867);
or U17815 (N_17815,N_16963,N_17394);
nand U17816 (N_17816,N_17196,N_17146);
or U17817 (N_17817,N_17077,N_17490);
and U17818 (N_17818,N_17054,N_17074);
xnor U17819 (N_17819,N_16848,N_17370);
or U17820 (N_17820,N_17241,N_17015);
or U17821 (N_17821,N_17477,N_16937);
and U17822 (N_17822,N_17173,N_16804);
nand U17823 (N_17823,N_17494,N_17116);
or U17824 (N_17824,N_17237,N_17139);
or U17825 (N_17825,N_16974,N_17330);
nor U17826 (N_17826,N_16838,N_17189);
nor U17827 (N_17827,N_17016,N_16989);
nand U17828 (N_17828,N_17589,N_17118);
or U17829 (N_17829,N_16912,N_16809);
and U17830 (N_17830,N_16855,N_17418);
nor U17831 (N_17831,N_16883,N_17416);
nor U17832 (N_17832,N_16890,N_17534);
nor U17833 (N_17833,N_17378,N_17278);
and U17834 (N_17834,N_17251,N_17254);
xor U17835 (N_17835,N_17321,N_17184);
xor U17836 (N_17836,N_16933,N_17027);
nor U17837 (N_17837,N_17463,N_17178);
nor U17838 (N_17838,N_17441,N_17357);
or U17839 (N_17839,N_16861,N_17249);
and U17840 (N_17840,N_16910,N_16981);
and U17841 (N_17841,N_17358,N_17195);
nor U17842 (N_17842,N_17291,N_16996);
xor U17843 (N_17843,N_17535,N_17379);
and U17844 (N_17844,N_17168,N_17561);
xnor U17845 (N_17845,N_17348,N_17383);
xnor U17846 (N_17846,N_17499,N_17436);
xor U17847 (N_17847,N_17052,N_17427);
nand U17848 (N_17848,N_17117,N_17007);
and U17849 (N_17849,N_17235,N_16928);
xnor U17850 (N_17850,N_16943,N_17414);
xnor U17851 (N_17851,N_17208,N_17498);
or U17852 (N_17852,N_17227,N_16965);
or U17853 (N_17853,N_17209,N_17246);
and U17854 (N_17854,N_17422,N_17107);
nand U17855 (N_17855,N_17466,N_17519);
nand U17856 (N_17856,N_16942,N_17157);
or U17857 (N_17857,N_17270,N_17413);
or U17858 (N_17858,N_16922,N_17570);
xor U17859 (N_17859,N_17243,N_17185);
and U17860 (N_17860,N_17030,N_17034);
or U17861 (N_17861,N_17048,N_16888);
nand U17862 (N_17862,N_16826,N_17066);
nor U17863 (N_17863,N_17262,N_17217);
or U17864 (N_17864,N_17271,N_17568);
nor U17865 (N_17865,N_17558,N_17204);
and U17866 (N_17866,N_17028,N_16827);
xor U17867 (N_17867,N_17067,N_17592);
and U17868 (N_17868,N_17385,N_17207);
or U17869 (N_17869,N_17483,N_17508);
nand U17870 (N_17870,N_17387,N_17183);
xor U17871 (N_17871,N_17500,N_17376);
nand U17872 (N_17872,N_16881,N_17442);
nor U17873 (N_17873,N_17238,N_17232);
or U17874 (N_17874,N_17288,N_17211);
and U17875 (N_17875,N_17402,N_17109);
nor U17876 (N_17876,N_17533,N_17287);
xnor U17877 (N_17877,N_17206,N_17342);
or U17878 (N_17878,N_17352,N_16875);
or U17879 (N_17879,N_17257,N_16984);
or U17880 (N_17880,N_17079,N_17256);
nor U17881 (N_17881,N_17327,N_17202);
or U17882 (N_17882,N_17597,N_17396);
nand U17883 (N_17883,N_17044,N_17006);
xnor U17884 (N_17884,N_16895,N_17192);
or U17885 (N_17885,N_16813,N_17462);
or U17886 (N_17886,N_17515,N_17359);
or U17887 (N_17887,N_17350,N_17345);
nand U17888 (N_17888,N_17395,N_17152);
nor U17889 (N_17889,N_17103,N_17447);
nand U17890 (N_17890,N_17190,N_16820);
or U17891 (N_17891,N_16952,N_16812);
xor U17892 (N_17892,N_17099,N_17557);
or U17893 (N_17893,N_17242,N_17354);
and U17894 (N_17894,N_17096,N_17353);
nand U17895 (N_17895,N_16957,N_16936);
and U17896 (N_17896,N_17590,N_17180);
nor U17897 (N_17897,N_17286,N_17503);
nand U17898 (N_17898,N_17062,N_17089);
and U17899 (N_17899,N_17377,N_17101);
nor U17900 (N_17900,N_17356,N_16934);
or U17901 (N_17901,N_16972,N_17403);
or U17902 (N_17902,N_16824,N_17400);
xor U17903 (N_17903,N_17138,N_17193);
xor U17904 (N_17904,N_17574,N_17440);
nor U17905 (N_17905,N_17166,N_17526);
or U17906 (N_17906,N_17449,N_17314);
or U17907 (N_17907,N_16975,N_16961);
or U17908 (N_17908,N_17380,N_17133);
nor U17909 (N_17909,N_17194,N_17491);
or U17910 (N_17910,N_16902,N_16862);
or U17911 (N_17911,N_16949,N_16816);
nand U17912 (N_17912,N_16815,N_16923);
nor U17913 (N_17913,N_17545,N_17134);
xor U17914 (N_17914,N_17181,N_17057);
or U17915 (N_17915,N_17059,N_16850);
or U17916 (N_17916,N_16947,N_16843);
xor U17917 (N_17917,N_17153,N_17174);
xor U17918 (N_17918,N_17276,N_17219);
nor U17919 (N_17919,N_16878,N_17065);
nor U17920 (N_17920,N_16803,N_17186);
nor U17921 (N_17921,N_17415,N_16938);
xor U17922 (N_17922,N_17544,N_17226);
and U17923 (N_17923,N_17516,N_17022);
and U17924 (N_17924,N_16925,N_16810);
xor U17925 (N_17925,N_17266,N_16917);
xor U17926 (N_17926,N_17381,N_17316);
nor U17927 (N_17927,N_17325,N_17221);
nand U17928 (N_17928,N_17423,N_17407);
or U17929 (N_17929,N_17169,N_17267);
xnor U17930 (N_17930,N_17151,N_16893);
or U17931 (N_17931,N_17144,N_17594);
nor U17932 (N_17932,N_17073,N_16818);
and U17933 (N_17933,N_16991,N_17553);
or U17934 (N_17934,N_17315,N_17584);
xor U17935 (N_17935,N_17310,N_17328);
xnor U17936 (N_17936,N_17397,N_17031);
nand U17937 (N_17937,N_17159,N_17233);
or U17938 (N_17938,N_17344,N_17444);
and U17939 (N_17939,N_17450,N_17033);
nor U17940 (N_17940,N_17029,N_17215);
xnor U17941 (N_17941,N_17485,N_17514);
nand U17942 (N_17942,N_17024,N_17368);
nor U17943 (N_17943,N_17595,N_17513);
nand U17944 (N_17944,N_17248,N_17520);
nand U17945 (N_17945,N_17523,N_17279);
and U17946 (N_17946,N_17250,N_17150);
or U17947 (N_17947,N_17482,N_17393);
or U17948 (N_17948,N_16805,N_17277);
or U17949 (N_17949,N_17372,N_16903);
nand U17950 (N_17950,N_16941,N_16854);
or U17951 (N_17951,N_16954,N_17550);
xor U17952 (N_17952,N_16924,N_16858);
nand U17953 (N_17953,N_16894,N_17326);
and U17954 (N_17954,N_17011,N_17154);
and U17955 (N_17955,N_17390,N_17336);
or U17956 (N_17956,N_17141,N_17547);
or U17957 (N_17957,N_17259,N_16929);
or U17958 (N_17958,N_17042,N_17213);
nand U17959 (N_17959,N_16958,N_17038);
nor U17960 (N_17960,N_16814,N_17283);
xor U17961 (N_17961,N_16819,N_17123);
and U17962 (N_17962,N_17084,N_16967);
xor U17963 (N_17963,N_17129,N_17323);
and U17964 (N_17964,N_16909,N_17004);
nor U17965 (N_17965,N_17136,N_17298);
or U17966 (N_17966,N_17391,N_17529);
or U17967 (N_17967,N_17581,N_17222);
xnor U17968 (N_17968,N_16823,N_17182);
nand U17969 (N_17969,N_17398,N_17069);
xnor U17970 (N_17970,N_17082,N_17554);
nand U17971 (N_17971,N_17043,N_17539);
nand U17972 (N_17972,N_17100,N_17455);
xnor U17973 (N_17973,N_17020,N_16885);
nand U17974 (N_17974,N_17355,N_17509);
xor U17975 (N_17975,N_17098,N_17591);
and U17976 (N_17976,N_17294,N_16966);
xor U17977 (N_17977,N_16976,N_16998);
xor U17978 (N_17978,N_16847,N_17471);
nand U17979 (N_17979,N_17261,N_17598);
or U17980 (N_17980,N_17039,N_17142);
or U17981 (N_17981,N_17212,N_17214);
nand U17982 (N_17982,N_17303,N_16857);
nand U17983 (N_17983,N_17579,N_17532);
nand U17984 (N_17984,N_17443,N_17187);
xnor U17985 (N_17985,N_17335,N_17349);
and U17986 (N_17986,N_17058,N_17484);
nor U17987 (N_17987,N_17124,N_17308);
and U17988 (N_17988,N_16948,N_17488);
or U17989 (N_17989,N_17468,N_16830);
nor U17990 (N_17990,N_17567,N_17068);
and U17991 (N_17991,N_16999,N_17343);
xnor U17992 (N_17992,N_17337,N_17428);
or U17993 (N_17993,N_16866,N_17216);
xor U17994 (N_17994,N_17121,N_17055);
nand U17995 (N_17995,N_17255,N_17265);
and U17996 (N_17996,N_17495,N_16987);
xor U17997 (N_17997,N_17210,N_17147);
or U17998 (N_17998,N_16979,N_17459);
nor U17999 (N_17999,N_17111,N_16859);
or U18000 (N_18000,N_17165,N_17598);
nor U18001 (N_18001,N_16828,N_17127);
and U18002 (N_18002,N_16874,N_17537);
xor U18003 (N_18003,N_16991,N_17030);
or U18004 (N_18004,N_17220,N_17454);
nor U18005 (N_18005,N_17527,N_17121);
nor U18006 (N_18006,N_17331,N_16826);
and U18007 (N_18007,N_17445,N_17585);
nand U18008 (N_18008,N_16961,N_17225);
or U18009 (N_18009,N_17372,N_16980);
nor U18010 (N_18010,N_17400,N_17229);
xor U18011 (N_18011,N_16982,N_17241);
nand U18012 (N_18012,N_16926,N_17385);
nor U18013 (N_18013,N_17414,N_17463);
or U18014 (N_18014,N_17473,N_17071);
nor U18015 (N_18015,N_16935,N_16866);
nor U18016 (N_18016,N_17090,N_16848);
xor U18017 (N_18017,N_17434,N_16951);
and U18018 (N_18018,N_16843,N_17150);
nor U18019 (N_18019,N_17573,N_16929);
and U18020 (N_18020,N_17401,N_17066);
nor U18021 (N_18021,N_17365,N_17044);
nand U18022 (N_18022,N_17541,N_16874);
or U18023 (N_18023,N_17526,N_17400);
nor U18024 (N_18024,N_17042,N_17274);
nand U18025 (N_18025,N_17225,N_17532);
nor U18026 (N_18026,N_17203,N_16917);
xnor U18027 (N_18027,N_17234,N_16830);
nor U18028 (N_18028,N_17021,N_17232);
and U18029 (N_18029,N_17115,N_17508);
xor U18030 (N_18030,N_16976,N_17085);
nor U18031 (N_18031,N_17355,N_16872);
and U18032 (N_18032,N_17305,N_16952);
xor U18033 (N_18033,N_16826,N_17214);
and U18034 (N_18034,N_16905,N_17175);
nand U18035 (N_18035,N_17534,N_17026);
xor U18036 (N_18036,N_17544,N_16869);
nor U18037 (N_18037,N_17002,N_17329);
xnor U18038 (N_18038,N_17234,N_17337);
or U18039 (N_18039,N_17417,N_17424);
and U18040 (N_18040,N_17217,N_17452);
xnor U18041 (N_18041,N_17293,N_17296);
or U18042 (N_18042,N_17380,N_17085);
xnor U18043 (N_18043,N_17504,N_17184);
and U18044 (N_18044,N_16904,N_17255);
nor U18045 (N_18045,N_17108,N_17326);
or U18046 (N_18046,N_17154,N_17365);
nor U18047 (N_18047,N_17427,N_17350);
or U18048 (N_18048,N_17274,N_17329);
nand U18049 (N_18049,N_17029,N_16935);
xor U18050 (N_18050,N_16925,N_17086);
and U18051 (N_18051,N_17052,N_17195);
nand U18052 (N_18052,N_16932,N_17236);
nor U18053 (N_18053,N_17303,N_17570);
nor U18054 (N_18054,N_17570,N_16998);
and U18055 (N_18055,N_17254,N_16976);
nor U18056 (N_18056,N_17480,N_17446);
or U18057 (N_18057,N_17357,N_16812);
and U18058 (N_18058,N_16860,N_16847);
xnor U18059 (N_18059,N_17311,N_17197);
and U18060 (N_18060,N_17127,N_17246);
xor U18061 (N_18061,N_16967,N_16994);
and U18062 (N_18062,N_17308,N_17502);
nor U18063 (N_18063,N_17035,N_17286);
nor U18064 (N_18064,N_16988,N_17045);
and U18065 (N_18065,N_17427,N_17289);
nor U18066 (N_18066,N_16947,N_17122);
and U18067 (N_18067,N_17114,N_17207);
nand U18068 (N_18068,N_17149,N_17492);
or U18069 (N_18069,N_17316,N_17505);
nor U18070 (N_18070,N_17230,N_17192);
and U18071 (N_18071,N_17380,N_17564);
nor U18072 (N_18072,N_17464,N_16937);
nand U18073 (N_18073,N_17454,N_17197);
or U18074 (N_18074,N_16987,N_17411);
and U18075 (N_18075,N_17086,N_17319);
and U18076 (N_18076,N_17484,N_17193);
and U18077 (N_18077,N_17041,N_17357);
and U18078 (N_18078,N_16810,N_16935);
and U18079 (N_18079,N_17225,N_17145);
nor U18080 (N_18080,N_17145,N_16948);
and U18081 (N_18081,N_16870,N_17104);
or U18082 (N_18082,N_17472,N_17097);
nor U18083 (N_18083,N_16862,N_17597);
xor U18084 (N_18084,N_17287,N_17210);
or U18085 (N_18085,N_17131,N_16953);
xnor U18086 (N_18086,N_17229,N_17035);
xnor U18087 (N_18087,N_17436,N_16800);
xnor U18088 (N_18088,N_16844,N_16903);
nor U18089 (N_18089,N_17055,N_16949);
nand U18090 (N_18090,N_17585,N_17342);
or U18091 (N_18091,N_17518,N_16893);
or U18092 (N_18092,N_17563,N_17482);
nor U18093 (N_18093,N_17586,N_17133);
nor U18094 (N_18094,N_17558,N_17440);
xor U18095 (N_18095,N_17384,N_17084);
xnor U18096 (N_18096,N_17284,N_16805);
and U18097 (N_18097,N_17101,N_17058);
xor U18098 (N_18098,N_16915,N_17513);
nand U18099 (N_18099,N_17349,N_16882);
or U18100 (N_18100,N_17539,N_16842);
nand U18101 (N_18101,N_17505,N_17537);
or U18102 (N_18102,N_17593,N_17304);
or U18103 (N_18103,N_17526,N_16969);
nand U18104 (N_18104,N_17184,N_17115);
and U18105 (N_18105,N_17480,N_17125);
nand U18106 (N_18106,N_17481,N_17157);
xnor U18107 (N_18107,N_17351,N_17170);
or U18108 (N_18108,N_16911,N_16966);
and U18109 (N_18109,N_16885,N_17226);
xor U18110 (N_18110,N_17092,N_17233);
or U18111 (N_18111,N_17086,N_17269);
and U18112 (N_18112,N_17259,N_17328);
or U18113 (N_18113,N_17180,N_17222);
nor U18114 (N_18114,N_17488,N_17311);
and U18115 (N_18115,N_17219,N_17084);
or U18116 (N_18116,N_17275,N_17506);
xnor U18117 (N_18117,N_17457,N_16906);
and U18118 (N_18118,N_17099,N_17091);
nor U18119 (N_18119,N_16905,N_17329);
nand U18120 (N_18120,N_17342,N_17122);
and U18121 (N_18121,N_17129,N_17311);
xor U18122 (N_18122,N_17455,N_16822);
or U18123 (N_18123,N_17250,N_17103);
and U18124 (N_18124,N_16895,N_17043);
nand U18125 (N_18125,N_17171,N_17018);
nor U18126 (N_18126,N_16902,N_17581);
and U18127 (N_18127,N_16961,N_17297);
xnor U18128 (N_18128,N_16846,N_17461);
nor U18129 (N_18129,N_17148,N_16835);
nor U18130 (N_18130,N_17252,N_16878);
nand U18131 (N_18131,N_16917,N_17259);
or U18132 (N_18132,N_17565,N_17379);
nor U18133 (N_18133,N_17557,N_17271);
nor U18134 (N_18134,N_16821,N_17114);
or U18135 (N_18135,N_17071,N_17591);
or U18136 (N_18136,N_16970,N_17057);
and U18137 (N_18137,N_17297,N_17369);
or U18138 (N_18138,N_17306,N_17379);
nor U18139 (N_18139,N_17097,N_17486);
xnor U18140 (N_18140,N_17288,N_16961);
nor U18141 (N_18141,N_16933,N_17493);
and U18142 (N_18142,N_17495,N_16830);
and U18143 (N_18143,N_17455,N_17196);
or U18144 (N_18144,N_17493,N_16996);
and U18145 (N_18145,N_17097,N_17012);
nand U18146 (N_18146,N_17175,N_17077);
or U18147 (N_18147,N_17580,N_17258);
or U18148 (N_18148,N_17448,N_17107);
nand U18149 (N_18149,N_17443,N_16823);
xor U18150 (N_18150,N_17582,N_17484);
xor U18151 (N_18151,N_16957,N_16954);
nor U18152 (N_18152,N_17439,N_17408);
nor U18153 (N_18153,N_17523,N_17102);
or U18154 (N_18154,N_16887,N_17509);
nor U18155 (N_18155,N_17091,N_17064);
xor U18156 (N_18156,N_17561,N_16921);
or U18157 (N_18157,N_17048,N_17034);
nand U18158 (N_18158,N_17015,N_16919);
nand U18159 (N_18159,N_17092,N_16909);
and U18160 (N_18160,N_17026,N_17097);
xnor U18161 (N_18161,N_17033,N_17414);
xnor U18162 (N_18162,N_17458,N_17218);
nand U18163 (N_18163,N_16877,N_17336);
nand U18164 (N_18164,N_16987,N_17580);
or U18165 (N_18165,N_17061,N_17363);
and U18166 (N_18166,N_16846,N_17150);
nand U18167 (N_18167,N_17076,N_16870);
or U18168 (N_18168,N_17331,N_17573);
and U18169 (N_18169,N_17445,N_17201);
nand U18170 (N_18170,N_16847,N_17149);
nand U18171 (N_18171,N_17165,N_16863);
and U18172 (N_18172,N_17529,N_17141);
nand U18173 (N_18173,N_17149,N_16992);
nor U18174 (N_18174,N_17013,N_17499);
and U18175 (N_18175,N_16867,N_16994);
xor U18176 (N_18176,N_17548,N_17565);
nor U18177 (N_18177,N_17392,N_17425);
nand U18178 (N_18178,N_17392,N_17546);
xor U18179 (N_18179,N_17190,N_17287);
or U18180 (N_18180,N_17264,N_17398);
nor U18181 (N_18181,N_16886,N_17426);
nor U18182 (N_18182,N_17011,N_17157);
or U18183 (N_18183,N_17094,N_17057);
or U18184 (N_18184,N_17589,N_16899);
or U18185 (N_18185,N_16838,N_16834);
nand U18186 (N_18186,N_17240,N_16803);
nand U18187 (N_18187,N_17215,N_17589);
nand U18188 (N_18188,N_17423,N_17194);
or U18189 (N_18189,N_17586,N_17119);
nor U18190 (N_18190,N_17357,N_17279);
nand U18191 (N_18191,N_17472,N_17122);
or U18192 (N_18192,N_17310,N_17112);
xor U18193 (N_18193,N_17407,N_17130);
and U18194 (N_18194,N_17152,N_17587);
and U18195 (N_18195,N_17472,N_17543);
nor U18196 (N_18196,N_17247,N_17311);
xnor U18197 (N_18197,N_16967,N_17472);
nand U18198 (N_18198,N_17227,N_17239);
xnor U18199 (N_18199,N_16952,N_17000);
xnor U18200 (N_18200,N_17442,N_16915);
nor U18201 (N_18201,N_16932,N_17587);
xnor U18202 (N_18202,N_16866,N_16955);
nand U18203 (N_18203,N_17116,N_17422);
xnor U18204 (N_18204,N_17347,N_17409);
and U18205 (N_18205,N_17070,N_17017);
or U18206 (N_18206,N_17381,N_16976);
xnor U18207 (N_18207,N_17312,N_17596);
or U18208 (N_18208,N_17175,N_17517);
nand U18209 (N_18209,N_17550,N_16830);
nand U18210 (N_18210,N_16887,N_17038);
or U18211 (N_18211,N_17082,N_16995);
nand U18212 (N_18212,N_17323,N_16939);
or U18213 (N_18213,N_17526,N_17393);
or U18214 (N_18214,N_16884,N_17316);
nor U18215 (N_18215,N_17214,N_17318);
and U18216 (N_18216,N_17396,N_17529);
nand U18217 (N_18217,N_17102,N_17152);
or U18218 (N_18218,N_16845,N_17168);
nor U18219 (N_18219,N_17320,N_16907);
nor U18220 (N_18220,N_17298,N_17502);
nor U18221 (N_18221,N_17075,N_17123);
nor U18222 (N_18222,N_17494,N_17144);
and U18223 (N_18223,N_17471,N_17306);
nor U18224 (N_18224,N_17278,N_17319);
and U18225 (N_18225,N_17306,N_16923);
nand U18226 (N_18226,N_17474,N_17052);
and U18227 (N_18227,N_17507,N_16848);
xnor U18228 (N_18228,N_16808,N_17297);
and U18229 (N_18229,N_17205,N_17423);
nand U18230 (N_18230,N_17435,N_17405);
nand U18231 (N_18231,N_17159,N_16891);
xnor U18232 (N_18232,N_16935,N_17375);
nand U18233 (N_18233,N_16802,N_17038);
nand U18234 (N_18234,N_16861,N_16810);
nor U18235 (N_18235,N_17554,N_17104);
nor U18236 (N_18236,N_17348,N_17590);
or U18237 (N_18237,N_17386,N_17194);
or U18238 (N_18238,N_16818,N_16965);
xnor U18239 (N_18239,N_16944,N_17131);
nand U18240 (N_18240,N_17075,N_17491);
or U18241 (N_18241,N_17533,N_17204);
nand U18242 (N_18242,N_17486,N_17180);
nand U18243 (N_18243,N_17084,N_17200);
and U18244 (N_18244,N_17588,N_17131);
nand U18245 (N_18245,N_16877,N_16828);
nand U18246 (N_18246,N_17173,N_17509);
or U18247 (N_18247,N_17420,N_17250);
or U18248 (N_18248,N_17466,N_17110);
nor U18249 (N_18249,N_17211,N_16910);
xnor U18250 (N_18250,N_17542,N_17023);
xor U18251 (N_18251,N_17116,N_16948);
and U18252 (N_18252,N_17257,N_17531);
nand U18253 (N_18253,N_17141,N_16913);
nand U18254 (N_18254,N_17599,N_17307);
nand U18255 (N_18255,N_17070,N_17266);
xor U18256 (N_18256,N_17499,N_16932);
xor U18257 (N_18257,N_16845,N_17218);
xnor U18258 (N_18258,N_16865,N_17485);
nand U18259 (N_18259,N_16832,N_17222);
or U18260 (N_18260,N_17541,N_17000);
or U18261 (N_18261,N_16879,N_17561);
or U18262 (N_18262,N_17280,N_17043);
xor U18263 (N_18263,N_17497,N_17235);
and U18264 (N_18264,N_16839,N_16948);
nand U18265 (N_18265,N_17216,N_17572);
or U18266 (N_18266,N_17219,N_17348);
or U18267 (N_18267,N_16897,N_17019);
xor U18268 (N_18268,N_17076,N_16972);
xor U18269 (N_18269,N_16916,N_17220);
xor U18270 (N_18270,N_17310,N_17551);
and U18271 (N_18271,N_17204,N_17205);
xor U18272 (N_18272,N_17278,N_17269);
nor U18273 (N_18273,N_17508,N_17551);
or U18274 (N_18274,N_17213,N_17323);
and U18275 (N_18275,N_17428,N_17334);
or U18276 (N_18276,N_17584,N_16929);
and U18277 (N_18277,N_16971,N_16897);
nand U18278 (N_18278,N_17192,N_17238);
nand U18279 (N_18279,N_17514,N_16885);
nor U18280 (N_18280,N_16956,N_17478);
xnor U18281 (N_18281,N_16960,N_17084);
nand U18282 (N_18282,N_17023,N_17578);
nand U18283 (N_18283,N_17562,N_17319);
or U18284 (N_18284,N_16942,N_17249);
or U18285 (N_18285,N_17448,N_16816);
xor U18286 (N_18286,N_17453,N_17450);
nand U18287 (N_18287,N_17257,N_17194);
or U18288 (N_18288,N_16923,N_16886);
nor U18289 (N_18289,N_17580,N_17077);
nand U18290 (N_18290,N_17128,N_17436);
xnor U18291 (N_18291,N_17448,N_17127);
nor U18292 (N_18292,N_17594,N_17291);
nand U18293 (N_18293,N_17393,N_16913);
and U18294 (N_18294,N_16926,N_16933);
and U18295 (N_18295,N_17537,N_16994);
xor U18296 (N_18296,N_17536,N_17108);
nor U18297 (N_18297,N_17137,N_17235);
or U18298 (N_18298,N_17044,N_16895);
or U18299 (N_18299,N_16910,N_17362);
nor U18300 (N_18300,N_17257,N_17428);
or U18301 (N_18301,N_17524,N_17177);
nand U18302 (N_18302,N_16983,N_17524);
and U18303 (N_18303,N_16887,N_16964);
or U18304 (N_18304,N_17031,N_17516);
xor U18305 (N_18305,N_17581,N_17344);
xnor U18306 (N_18306,N_17292,N_17528);
or U18307 (N_18307,N_17134,N_17004);
nand U18308 (N_18308,N_17168,N_16856);
nor U18309 (N_18309,N_16994,N_17118);
xor U18310 (N_18310,N_17567,N_17343);
and U18311 (N_18311,N_17303,N_16925);
nor U18312 (N_18312,N_17261,N_17541);
and U18313 (N_18313,N_17496,N_16931);
or U18314 (N_18314,N_17056,N_17175);
xor U18315 (N_18315,N_17133,N_16994);
xnor U18316 (N_18316,N_17067,N_17271);
nand U18317 (N_18317,N_16938,N_17089);
nor U18318 (N_18318,N_17368,N_17110);
nand U18319 (N_18319,N_17582,N_16935);
xor U18320 (N_18320,N_17292,N_17439);
or U18321 (N_18321,N_17176,N_17253);
nor U18322 (N_18322,N_17146,N_17241);
or U18323 (N_18323,N_17533,N_16952);
nor U18324 (N_18324,N_16961,N_17255);
nor U18325 (N_18325,N_17308,N_17548);
nor U18326 (N_18326,N_17315,N_17504);
xnor U18327 (N_18327,N_17079,N_17161);
or U18328 (N_18328,N_17072,N_16893);
nor U18329 (N_18329,N_17168,N_16952);
nand U18330 (N_18330,N_17534,N_17418);
nand U18331 (N_18331,N_17526,N_16982);
nand U18332 (N_18332,N_17309,N_17354);
nor U18333 (N_18333,N_17514,N_17232);
nor U18334 (N_18334,N_17325,N_17538);
or U18335 (N_18335,N_16804,N_16973);
xnor U18336 (N_18336,N_17430,N_17277);
and U18337 (N_18337,N_17134,N_17567);
nor U18338 (N_18338,N_17584,N_17086);
or U18339 (N_18339,N_17029,N_16940);
or U18340 (N_18340,N_17170,N_17520);
and U18341 (N_18341,N_17170,N_16999);
or U18342 (N_18342,N_17313,N_17468);
nor U18343 (N_18343,N_17339,N_17343);
nand U18344 (N_18344,N_16998,N_16928);
or U18345 (N_18345,N_16914,N_16837);
nand U18346 (N_18346,N_16985,N_17271);
nor U18347 (N_18347,N_16917,N_17351);
or U18348 (N_18348,N_17119,N_17510);
nand U18349 (N_18349,N_17037,N_17188);
or U18350 (N_18350,N_17461,N_16861);
or U18351 (N_18351,N_16959,N_16889);
and U18352 (N_18352,N_17238,N_17438);
xor U18353 (N_18353,N_16859,N_17188);
nor U18354 (N_18354,N_17484,N_16944);
nand U18355 (N_18355,N_17516,N_16863);
nor U18356 (N_18356,N_17492,N_16912);
xnor U18357 (N_18357,N_17271,N_17327);
nand U18358 (N_18358,N_17582,N_17364);
nor U18359 (N_18359,N_17162,N_17263);
nor U18360 (N_18360,N_17558,N_17417);
or U18361 (N_18361,N_17429,N_16959);
nor U18362 (N_18362,N_16819,N_17364);
nand U18363 (N_18363,N_17543,N_16845);
nor U18364 (N_18364,N_17355,N_16841);
and U18365 (N_18365,N_17274,N_17170);
nor U18366 (N_18366,N_17407,N_16824);
or U18367 (N_18367,N_17525,N_17535);
nand U18368 (N_18368,N_17492,N_16893);
nor U18369 (N_18369,N_17315,N_17558);
nor U18370 (N_18370,N_17420,N_17414);
or U18371 (N_18371,N_17495,N_17539);
nand U18372 (N_18372,N_17303,N_16934);
or U18373 (N_18373,N_16977,N_17171);
or U18374 (N_18374,N_17368,N_17519);
and U18375 (N_18375,N_16994,N_17469);
or U18376 (N_18376,N_17557,N_17576);
nand U18377 (N_18377,N_17397,N_17524);
and U18378 (N_18378,N_17369,N_17309);
nand U18379 (N_18379,N_17038,N_17361);
nand U18380 (N_18380,N_17067,N_17128);
nor U18381 (N_18381,N_17117,N_17579);
and U18382 (N_18382,N_17021,N_17267);
and U18383 (N_18383,N_16937,N_17159);
xnor U18384 (N_18384,N_16816,N_17447);
and U18385 (N_18385,N_17095,N_17556);
xor U18386 (N_18386,N_17245,N_17320);
nor U18387 (N_18387,N_17148,N_17292);
nand U18388 (N_18388,N_17503,N_17593);
nand U18389 (N_18389,N_17169,N_17202);
nand U18390 (N_18390,N_17000,N_16827);
nor U18391 (N_18391,N_17388,N_17039);
or U18392 (N_18392,N_16994,N_17334);
xnor U18393 (N_18393,N_17094,N_17331);
or U18394 (N_18394,N_17038,N_17237);
and U18395 (N_18395,N_17566,N_17544);
and U18396 (N_18396,N_17506,N_17563);
and U18397 (N_18397,N_16889,N_16962);
nand U18398 (N_18398,N_16814,N_17580);
xnor U18399 (N_18399,N_17271,N_17453);
nor U18400 (N_18400,N_17747,N_17997);
nor U18401 (N_18401,N_18110,N_18158);
and U18402 (N_18402,N_18114,N_18310);
nand U18403 (N_18403,N_17638,N_18386);
nor U18404 (N_18404,N_18113,N_17738);
xnor U18405 (N_18405,N_17737,N_18177);
xnor U18406 (N_18406,N_18300,N_17977);
or U18407 (N_18407,N_18013,N_17918);
xor U18408 (N_18408,N_18213,N_17728);
xnor U18409 (N_18409,N_18278,N_17673);
or U18410 (N_18410,N_18341,N_18121);
xor U18411 (N_18411,N_18348,N_17791);
nand U18412 (N_18412,N_17926,N_17627);
nand U18413 (N_18413,N_18159,N_18157);
nand U18414 (N_18414,N_17601,N_18023);
or U18415 (N_18415,N_17809,N_18273);
xor U18416 (N_18416,N_17818,N_17943);
nor U18417 (N_18417,N_17692,N_17713);
xor U18418 (N_18418,N_18365,N_18099);
nor U18419 (N_18419,N_17848,N_17633);
or U18420 (N_18420,N_17605,N_17919);
xor U18421 (N_18421,N_18096,N_18184);
and U18422 (N_18422,N_17635,N_18027);
nand U18423 (N_18423,N_18125,N_18144);
xnor U18424 (N_18424,N_17617,N_17705);
nor U18425 (N_18425,N_17624,N_17701);
xnor U18426 (N_18426,N_18391,N_18396);
nand U18427 (N_18427,N_18281,N_18200);
or U18428 (N_18428,N_18349,N_18091);
and U18429 (N_18429,N_17874,N_18112);
nand U18430 (N_18430,N_17972,N_17929);
nand U18431 (N_18431,N_17801,N_18324);
or U18432 (N_18432,N_18132,N_17654);
or U18433 (N_18433,N_17759,N_18046);
xor U18434 (N_18434,N_18347,N_17726);
or U18435 (N_18435,N_18336,N_17708);
and U18436 (N_18436,N_17651,N_17865);
and U18437 (N_18437,N_18179,N_17664);
or U18438 (N_18438,N_18173,N_18380);
nand U18439 (N_18439,N_18216,N_18176);
nor U18440 (N_18440,N_17625,N_18095);
or U18441 (N_18441,N_17946,N_17922);
or U18442 (N_18442,N_17764,N_17757);
nor U18443 (N_18443,N_17931,N_18215);
and U18444 (N_18444,N_18038,N_17873);
nor U18445 (N_18445,N_17856,N_17942);
or U18446 (N_18446,N_17661,N_17748);
nor U18447 (N_18447,N_17715,N_17973);
or U18448 (N_18448,N_17703,N_17802);
nor U18449 (N_18449,N_17716,N_17915);
nor U18450 (N_18450,N_18131,N_18346);
nand U18451 (N_18451,N_17806,N_17677);
xor U18452 (N_18452,N_18282,N_18171);
or U18453 (N_18453,N_17823,N_18366);
or U18454 (N_18454,N_18235,N_17699);
or U18455 (N_18455,N_17678,N_17666);
and U18456 (N_18456,N_17618,N_17730);
or U18457 (N_18457,N_18207,N_17644);
nand U18458 (N_18458,N_18033,N_17993);
or U18459 (N_18459,N_18355,N_17667);
nand U18460 (N_18460,N_17911,N_17615);
and U18461 (N_18461,N_17777,N_17945);
nand U18462 (N_18462,N_17676,N_18382);
nand U18463 (N_18463,N_17871,N_17976);
and U18464 (N_18464,N_18323,N_17887);
nand U18465 (N_18465,N_18383,N_17690);
nand U18466 (N_18466,N_17729,N_18289);
nor U18467 (N_18467,N_17917,N_18128);
nor U18468 (N_18468,N_18045,N_18206);
or U18469 (N_18469,N_18362,N_18066);
and U18470 (N_18470,N_18149,N_17753);
xnor U18471 (N_18471,N_17832,N_17895);
nor U18472 (N_18472,N_17710,N_18389);
nand U18473 (N_18473,N_18162,N_17826);
xor U18474 (N_18474,N_18118,N_18097);
nand U18475 (N_18475,N_18205,N_18223);
and U18476 (N_18476,N_17657,N_17751);
xnor U18477 (N_18477,N_18369,N_17820);
or U18478 (N_18478,N_17763,N_17797);
xor U18479 (N_18479,N_18250,N_18185);
and U18480 (N_18480,N_17653,N_17902);
or U18481 (N_18481,N_18183,N_17768);
nor U18482 (N_18482,N_18260,N_18228);
xor U18483 (N_18483,N_17960,N_18270);
or U18484 (N_18484,N_18124,N_18364);
and U18485 (N_18485,N_18210,N_18029);
and U18486 (N_18486,N_18318,N_18329);
nand U18487 (N_18487,N_17689,N_17988);
or U18488 (N_18488,N_17670,N_18017);
and U18489 (N_18489,N_17830,N_17967);
nand U18490 (N_18490,N_17884,N_17955);
nor U18491 (N_18491,N_17890,N_17933);
nand U18492 (N_18492,N_18198,N_17805);
xor U18493 (N_18493,N_18202,N_17838);
and U18494 (N_18494,N_17658,N_18302);
or U18495 (N_18495,N_17857,N_17800);
xnor U18496 (N_18496,N_18219,N_18381);
and U18497 (N_18497,N_17813,N_18344);
nor U18498 (N_18498,N_17695,N_17686);
nor U18499 (N_18499,N_18056,N_17810);
and U18500 (N_18500,N_18003,N_17683);
or U18501 (N_18501,N_17603,N_18077);
nor U18502 (N_18502,N_18014,N_17864);
or U18503 (N_18503,N_18280,N_18317);
xor U18504 (N_18504,N_17649,N_17629);
nand U18505 (N_18505,N_18242,N_18005);
or U18506 (N_18506,N_18353,N_18292);
and U18507 (N_18507,N_18330,N_18335);
nand U18508 (N_18508,N_18150,N_17854);
or U18509 (N_18509,N_18286,N_18062);
nor U18510 (N_18510,N_18254,N_18134);
nand U18511 (N_18511,N_18246,N_17652);
nor U18512 (N_18512,N_17900,N_17841);
xor U18513 (N_18513,N_18360,N_18293);
nand U18514 (N_18514,N_18269,N_18039);
or U18515 (N_18515,N_18195,N_17672);
and U18516 (N_18516,N_18049,N_17742);
or U18517 (N_18517,N_17821,N_18079);
and U18518 (N_18518,N_17839,N_18026);
and U18519 (N_18519,N_17965,N_17788);
nand U18520 (N_18520,N_18175,N_17626);
nor U18521 (N_18521,N_18030,N_17935);
xor U18522 (N_18522,N_17698,N_17964);
xor U18523 (N_18523,N_18262,N_18070);
nor U18524 (N_18524,N_18354,N_17790);
and U18525 (N_18525,N_18034,N_18174);
and U18526 (N_18526,N_17991,N_18082);
and U18527 (N_18527,N_17869,N_18322);
nand U18528 (N_18528,N_18040,N_17743);
xnor U18529 (N_18529,N_18052,N_18108);
and U18530 (N_18530,N_18301,N_17794);
xnor U18531 (N_18531,N_18351,N_18140);
or U18532 (N_18532,N_17614,N_18006);
nand U18533 (N_18533,N_18123,N_18116);
and U18534 (N_18534,N_17901,N_17875);
xnor U18535 (N_18535,N_18016,N_18084);
nor U18536 (N_18536,N_17630,N_18387);
or U18537 (N_18537,N_17789,N_17978);
nand U18538 (N_18538,N_18265,N_18368);
xor U18539 (N_18539,N_18352,N_17663);
or U18540 (N_18540,N_17866,N_18000);
and U18541 (N_18541,N_18020,N_18220);
nand U18542 (N_18542,N_18272,N_18343);
nand U18543 (N_18543,N_18284,N_18160);
nor U18544 (N_18544,N_17816,N_18306);
or U18545 (N_18545,N_17799,N_18148);
or U18546 (N_18546,N_17623,N_18231);
nand U18547 (N_18547,N_17606,N_17819);
and U18548 (N_18548,N_17778,N_18204);
or U18549 (N_18549,N_18068,N_17732);
and U18550 (N_18550,N_17659,N_18161);
and U18551 (N_18551,N_17752,N_17923);
nor U18552 (N_18552,N_17662,N_18221);
nand U18553 (N_18553,N_18251,N_17824);
xnor U18554 (N_18554,N_17750,N_17771);
and U18555 (N_18555,N_17693,N_18044);
nand U18556 (N_18556,N_17992,N_17746);
or U18557 (N_18557,N_17712,N_17891);
xor U18558 (N_18558,N_18094,N_17947);
or U18559 (N_18559,N_17928,N_18230);
nand U18560 (N_18560,N_18129,N_18363);
nand U18561 (N_18561,N_17707,N_18305);
nor U18562 (N_18562,N_18345,N_17607);
nor U18563 (N_18563,N_18119,N_18055);
nand U18564 (N_18564,N_17641,N_17787);
xnor U18565 (N_18565,N_17700,N_17880);
or U18566 (N_18566,N_17811,N_17998);
nand U18567 (N_18567,N_18307,N_17984);
or U18568 (N_18568,N_18268,N_18313);
xnor U18569 (N_18569,N_17840,N_17883);
nand U18570 (N_18570,N_17620,N_17671);
xor U18571 (N_18571,N_18007,N_18285);
and U18572 (N_18572,N_17734,N_17969);
xor U18573 (N_18573,N_17674,N_17861);
nand U18574 (N_18574,N_18065,N_18209);
or U18575 (N_18575,N_18130,N_18358);
nor U18576 (N_18576,N_18264,N_17709);
nor U18577 (N_18577,N_17613,N_17688);
xnor U18578 (N_18578,N_18290,N_18390);
xnor U18579 (N_18579,N_17899,N_17814);
and U18580 (N_18580,N_17872,N_17851);
nor U18581 (N_18581,N_18115,N_17879);
nand U18582 (N_18582,N_17975,N_18263);
xnor U18583 (N_18583,N_17985,N_18192);
nor U18584 (N_18584,N_18092,N_17951);
nor U18585 (N_18585,N_17749,N_17995);
and U18586 (N_18586,N_18339,N_17815);
or U18587 (N_18587,N_17980,N_17783);
or U18588 (N_18588,N_18085,N_18241);
nand U18589 (N_18589,N_18249,N_17718);
or U18590 (N_18590,N_17829,N_17648);
and U18591 (N_18591,N_18011,N_18397);
nor U18592 (N_18592,N_17961,N_17665);
nor U18593 (N_18593,N_17850,N_17916);
and U18594 (N_18594,N_18002,N_17956);
or U18595 (N_18595,N_17608,N_18009);
nand U18596 (N_18596,N_18378,N_18088);
nor U18597 (N_18597,N_18021,N_17668);
or U18598 (N_18598,N_18189,N_17912);
or U18599 (N_18599,N_17691,N_18357);
xnor U18600 (N_18600,N_18089,N_18076);
and U18601 (N_18601,N_18093,N_17877);
nand U18602 (N_18602,N_17881,N_17731);
nor U18603 (N_18603,N_18139,N_17650);
nor U18604 (N_18604,N_17979,N_17735);
nand U18605 (N_18605,N_17842,N_18122);
and U18606 (N_18606,N_18145,N_17774);
nor U18607 (N_18607,N_17723,N_18164);
and U18608 (N_18608,N_18187,N_17999);
xnor U18609 (N_18609,N_17619,N_17739);
xnor U18610 (N_18610,N_18277,N_18350);
or U18611 (N_18611,N_18001,N_18111);
or U18612 (N_18612,N_18072,N_18022);
xnor U18613 (N_18613,N_17770,N_17982);
and U18614 (N_18614,N_17682,N_18194);
xor U18615 (N_18615,N_17903,N_17836);
nor U18616 (N_18616,N_18245,N_18047);
or U18617 (N_18617,N_18107,N_18170);
and U18618 (N_18618,N_17745,N_17795);
or U18619 (N_18619,N_18295,N_18253);
or U18620 (N_18620,N_18069,N_18208);
nor U18621 (N_18621,N_18193,N_17934);
nor U18622 (N_18622,N_18057,N_18155);
or U18623 (N_18623,N_18255,N_17876);
nor U18624 (N_18624,N_18308,N_17655);
and U18625 (N_18625,N_17860,N_17906);
nor U18626 (N_18626,N_17827,N_17831);
and U18627 (N_18627,N_17740,N_17858);
nor U18628 (N_18628,N_18053,N_17833);
nor U18629 (N_18629,N_17907,N_18217);
nand U18630 (N_18630,N_18051,N_18063);
and U18631 (N_18631,N_17948,N_18137);
nand U18632 (N_18632,N_18156,N_17642);
or U18633 (N_18633,N_18398,N_17796);
or U18634 (N_18634,N_17958,N_17974);
nand U18635 (N_18635,N_17825,N_17762);
xor U18636 (N_18636,N_17779,N_17904);
nor U18637 (N_18637,N_18303,N_18218);
or U18638 (N_18638,N_17886,N_17761);
xnor U18639 (N_18639,N_18257,N_18178);
and U18640 (N_18640,N_18117,N_18340);
nand U18641 (N_18641,N_17898,N_18147);
nand U18642 (N_18642,N_17636,N_18104);
nor U18643 (N_18643,N_17893,N_17987);
xor U18644 (N_18644,N_18168,N_18247);
xnor U18645 (N_18645,N_17954,N_17639);
xor U18646 (N_18646,N_18212,N_18059);
nor U18647 (N_18647,N_17989,N_18138);
xor U18648 (N_18648,N_18154,N_18276);
nand U18649 (N_18649,N_18239,N_17882);
or U18650 (N_18650,N_18237,N_17938);
or U18651 (N_18651,N_18367,N_18214);
nand U18652 (N_18652,N_17616,N_18298);
and U18653 (N_18653,N_18211,N_17714);
nand U18654 (N_18654,N_17970,N_17910);
and U18655 (N_18655,N_18064,N_17936);
xor U18656 (N_18656,N_17862,N_17957);
nor U18657 (N_18657,N_17610,N_18222);
and U18658 (N_18658,N_18181,N_17645);
nand U18659 (N_18659,N_18165,N_17711);
nor U18660 (N_18660,N_18141,N_17983);
nand U18661 (N_18661,N_17828,N_18120);
nor U18662 (N_18662,N_18325,N_17822);
and U18663 (N_18663,N_17765,N_18126);
or U18664 (N_18664,N_17808,N_17807);
nand U18665 (N_18665,N_18025,N_17843);
nor U18666 (N_18666,N_17849,N_17949);
or U18667 (N_18667,N_18332,N_18287);
xnor U18668 (N_18668,N_17696,N_17798);
or U18669 (N_18669,N_18312,N_17622);
nor U18670 (N_18670,N_17758,N_18394);
or U18671 (N_18671,N_18182,N_18199);
and U18672 (N_18672,N_18060,N_18032);
xor U18673 (N_18673,N_17812,N_17996);
nor U18674 (N_18674,N_18188,N_18041);
or U18675 (N_18675,N_18337,N_17669);
and U18676 (N_18676,N_18248,N_18288);
and U18677 (N_18677,N_17885,N_17769);
nor U18678 (N_18678,N_18393,N_17994);
and U18679 (N_18679,N_18010,N_17859);
nand U18680 (N_18680,N_17835,N_17952);
nor U18681 (N_18681,N_18304,N_17971);
xor U18682 (N_18682,N_18374,N_17932);
nor U18683 (N_18683,N_17896,N_18078);
nand U18684 (N_18684,N_17863,N_18291);
nand U18685 (N_18685,N_18167,N_17717);
nor U18686 (N_18686,N_18196,N_18236);
nand U18687 (N_18687,N_18201,N_18224);
nor U18688 (N_18688,N_17892,N_17817);
or U18689 (N_18689,N_17773,N_18080);
nor U18690 (N_18690,N_18012,N_18048);
or U18691 (N_18691,N_18334,N_18371);
xor U18692 (N_18692,N_18127,N_18018);
xor U18693 (N_18693,N_18042,N_18244);
and U18694 (N_18694,N_17844,N_18311);
or U18695 (N_18695,N_18271,N_18143);
nand U18696 (N_18696,N_18316,N_17981);
xnor U18697 (N_18697,N_18338,N_17782);
nand U18698 (N_18698,N_18163,N_17905);
or U18699 (N_18699,N_17724,N_17611);
or U18700 (N_18700,N_18252,N_17656);
and U18701 (N_18701,N_17754,N_17804);
or U18702 (N_18702,N_17719,N_18342);
nor U18703 (N_18703,N_17602,N_18197);
nor U18704 (N_18704,N_17894,N_17697);
nor U18705 (N_18705,N_18100,N_17744);
nand U18706 (N_18706,N_17687,N_18359);
nor U18707 (N_18707,N_18142,N_18008);
xnor U18708 (N_18708,N_18024,N_17939);
nand U18709 (N_18709,N_18320,N_18399);
nand U18710 (N_18710,N_18388,N_17868);
and U18711 (N_18711,N_17920,N_18135);
nor U18712 (N_18712,N_17959,N_17736);
or U18713 (N_18713,N_17870,N_18151);
or U18714 (N_18714,N_18233,N_18266);
nand U18715 (N_18715,N_18191,N_18275);
or U18716 (N_18716,N_17937,N_17950);
nand U18717 (N_18717,N_17733,N_18385);
nand U18718 (N_18718,N_17781,N_18395);
xor U18719 (N_18719,N_18061,N_18067);
or U18720 (N_18720,N_18296,N_18327);
xor U18721 (N_18721,N_17847,N_17679);
nor U18722 (N_18722,N_18073,N_18172);
or U18723 (N_18723,N_17646,N_17855);
nand U18724 (N_18724,N_18086,N_17852);
and U18725 (N_18725,N_17925,N_17940);
nand U18726 (N_18726,N_18074,N_18050);
nor U18727 (N_18727,N_17741,N_17793);
and U18728 (N_18728,N_18106,N_18136);
xnor U18729 (N_18729,N_18356,N_17704);
and U18730 (N_18730,N_18283,N_17647);
nand U18731 (N_18731,N_17621,N_17681);
and U18732 (N_18732,N_17775,N_18377);
nand U18733 (N_18733,N_17962,N_18294);
and U18734 (N_18734,N_17609,N_18102);
or U18735 (N_18735,N_17776,N_17784);
and U18736 (N_18736,N_18238,N_18180);
and U18737 (N_18737,N_18326,N_17845);
and U18738 (N_18738,N_18152,N_18259);
nand U18739 (N_18739,N_18153,N_18037);
xnor U18740 (N_18740,N_17600,N_17953);
nor U18741 (N_18741,N_18225,N_18054);
xnor U18742 (N_18742,N_18372,N_17846);
nand U18743 (N_18743,N_17722,N_18314);
or U18744 (N_18744,N_18274,N_18169);
nor U18745 (N_18745,N_18258,N_18083);
nor U18746 (N_18746,N_17628,N_17968);
nand U18747 (N_18747,N_18058,N_18019);
nand U18748 (N_18748,N_17640,N_18328);
and U18749 (N_18749,N_17720,N_18321);
xor U18750 (N_18750,N_17721,N_18090);
or U18751 (N_18751,N_17675,N_18015);
or U18752 (N_18752,N_17913,N_17755);
nand U18753 (N_18753,N_18035,N_18146);
nor U18754 (N_18754,N_18256,N_17612);
xnor U18755 (N_18755,N_18309,N_18028);
nand U18756 (N_18756,N_17756,N_17924);
or U18757 (N_18757,N_18279,N_18361);
and U18758 (N_18758,N_17694,N_18319);
and U18759 (N_18759,N_17921,N_18331);
and U18760 (N_18760,N_18379,N_18133);
and U18761 (N_18761,N_17786,N_18376);
or U18762 (N_18762,N_17990,N_18098);
nand U18763 (N_18763,N_17914,N_17727);
xnor U18764 (N_18764,N_18333,N_17643);
or U18765 (N_18765,N_17632,N_18234);
nand U18766 (N_18766,N_18392,N_17680);
or U18767 (N_18767,N_17888,N_17766);
nor U18768 (N_18768,N_17941,N_18243);
nand U18769 (N_18769,N_17637,N_18373);
nor U18770 (N_18770,N_17767,N_17837);
nor U18771 (N_18771,N_17785,N_18232);
or U18772 (N_18772,N_18071,N_17889);
and U18773 (N_18773,N_17878,N_18227);
or U18774 (N_18774,N_17897,N_17772);
nor U18775 (N_18775,N_17834,N_17867);
xnor U18776 (N_18776,N_18043,N_18261);
xnor U18777 (N_18777,N_17685,N_17853);
nor U18778 (N_18778,N_17604,N_17660);
and U18779 (N_18779,N_18240,N_17944);
or U18780 (N_18780,N_17634,N_17908);
nand U18781 (N_18781,N_18375,N_17780);
nand U18782 (N_18782,N_17760,N_18315);
or U18783 (N_18783,N_18105,N_17930);
or U18784 (N_18784,N_17803,N_18203);
nor U18785 (N_18785,N_17706,N_17631);
or U18786 (N_18786,N_18190,N_17927);
nor U18787 (N_18787,N_18101,N_18103);
or U18788 (N_18788,N_18229,N_17725);
xnor U18789 (N_18789,N_18297,N_18109);
nand U18790 (N_18790,N_18081,N_18087);
or U18791 (N_18791,N_18384,N_18075);
or U18792 (N_18792,N_17966,N_18299);
nand U18793 (N_18793,N_17986,N_18370);
nor U18794 (N_18794,N_17684,N_17963);
and U18795 (N_18795,N_18031,N_17909);
nor U18796 (N_18796,N_18166,N_18267);
and U18797 (N_18797,N_18036,N_18186);
xor U18798 (N_18798,N_17792,N_18226);
nor U18799 (N_18799,N_18004,N_17702);
xnor U18800 (N_18800,N_18085,N_17619);
nor U18801 (N_18801,N_18314,N_18074);
or U18802 (N_18802,N_17988,N_17864);
or U18803 (N_18803,N_18196,N_17761);
nand U18804 (N_18804,N_18289,N_18326);
xor U18805 (N_18805,N_17625,N_17772);
or U18806 (N_18806,N_17993,N_17979);
nor U18807 (N_18807,N_17965,N_17636);
and U18808 (N_18808,N_18308,N_17632);
xor U18809 (N_18809,N_17896,N_18094);
nor U18810 (N_18810,N_17824,N_18366);
or U18811 (N_18811,N_18283,N_17848);
or U18812 (N_18812,N_18264,N_17605);
xnor U18813 (N_18813,N_17922,N_17839);
xnor U18814 (N_18814,N_17659,N_17664);
and U18815 (N_18815,N_17824,N_18016);
or U18816 (N_18816,N_17913,N_17885);
nor U18817 (N_18817,N_17935,N_18221);
xnor U18818 (N_18818,N_18147,N_17757);
or U18819 (N_18819,N_18239,N_17737);
nand U18820 (N_18820,N_17647,N_17929);
or U18821 (N_18821,N_18020,N_18301);
and U18822 (N_18822,N_17964,N_18272);
or U18823 (N_18823,N_17930,N_17998);
or U18824 (N_18824,N_18072,N_17647);
and U18825 (N_18825,N_18206,N_17772);
or U18826 (N_18826,N_18149,N_17604);
xor U18827 (N_18827,N_17671,N_18325);
and U18828 (N_18828,N_18344,N_18159);
or U18829 (N_18829,N_18265,N_18186);
nor U18830 (N_18830,N_18059,N_17888);
and U18831 (N_18831,N_17618,N_18325);
nor U18832 (N_18832,N_17756,N_17725);
and U18833 (N_18833,N_18242,N_18013);
nand U18834 (N_18834,N_18068,N_17807);
and U18835 (N_18835,N_18266,N_17645);
or U18836 (N_18836,N_17726,N_18058);
xnor U18837 (N_18837,N_17800,N_18184);
and U18838 (N_18838,N_17853,N_17631);
nor U18839 (N_18839,N_17622,N_17847);
xor U18840 (N_18840,N_18368,N_18013);
nor U18841 (N_18841,N_17732,N_18168);
xnor U18842 (N_18842,N_17813,N_18147);
or U18843 (N_18843,N_17738,N_18280);
nor U18844 (N_18844,N_18039,N_17666);
xor U18845 (N_18845,N_17669,N_17810);
and U18846 (N_18846,N_18150,N_17677);
xor U18847 (N_18847,N_17655,N_18343);
nor U18848 (N_18848,N_18274,N_17609);
and U18849 (N_18849,N_18111,N_18372);
nor U18850 (N_18850,N_17943,N_17767);
nor U18851 (N_18851,N_17640,N_18189);
nand U18852 (N_18852,N_17708,N_17854);
nand U18853 (N_18853,N_17877,N_17667);
nor U18854 (N_18854,N_18058,N_17766);
or U18855 (N_18855,N_18096,N_18040);
nand U18856 (N_18856,N_18198,N_17743);
or U18857 (N_18857,N_18310,N_18193);
nand U18858 (N_18858,N_17703,N_18234);
or U18859 (N_18859,N_17900,N_17885);
or U18860 (N_18860,N_17976,N_17865);
or U18861 (N_18861,N_18091,N_17606);
xor U18862 (N_18862,N_18012,N_17769);
and U18863 (N_18863,N_18313,N_17927);
and U18864 (N_18864,N_17620,N_17988);
nand U18865 (N_18865,N_18230,N_17832);
xor U18866 (N_18866,N_18340,N_18115);
xnor U18867 (N_18867,N_17602,N_18267);
xor U18868 (N_18868,N_17855,N_18378);
nor U18869 (N_18869,N_17765,N_17848);
nand U18870 (N_18870,N_17921,N_18384);
or U18871 (N_18871,N_17802,N_18259);
xor U18872 (N_18872,N_18126,N_17739);
xor U18873 (N_18873,N_18282,N_18194);
nand U18874 (N_18874,N_18247,N_18060);
and U18875 (N_18875,N_18087,N_17988);
nor U18876 (N_18876,N_18333,N_18346);
nand U18877 (N_18877,N_17919,N_18098);
or U18878 (N_18878,N_17844,N_18328);
nor U18879 (N_18879,N_17987,N_18001);
nor U18880 (N_18880,N_17649,N_18060);
and U18881 (N_18881,N_17851,N_18339);
and U18882 (N_18882,N_17916,N_18052);
nor U18883 (N_18883,N_18201,N_18379);
nor U18884 (N_18884,N_18020,N_18208);
nand U18885 (N_18885,N_18026,N_17972);
nand U18886 (N_18886,N_17804,N_18315);
xor U18887 (N_18887,N_17604,N_18293);
nand U18888 (N_18888,N_17937,N_18278);
nor U18889 (N_18889,N_17928,N_18190);
or U18890 (N_18890,N_18308,N_18128);
xnor U18891 (N_18891,N_17732,N_17759);
nand U18892 (N_18892,N_17807,N_17749);
or U18893 (N_18893,N_18023,N_17958);
nor U18894 (N_18894,N_18199,N_17695);
nor U18895 (N_18895,N_17920,N_18243);
or U18896 (N_18896,N_18098,N_17833);
nor U18897 (N_18897,N_17758,N_18321);
nor U18898 (N_18898,N_18309,N_17866);
or U18899 (N_18899,N_17791,N_18002);
nor U18900 (N_18900,N_18138,N_17618);
nand U18901 (N_18901,N_18391,N_17727);
or U18902 (N_18902,N_17806,N_17662);
and U18903 (N_18903,N_17829,N_17900);
xor U18904 (N_18904,N_18279,N_18101);
nor U18905 (N_18905,N_17799,N_17809);
nor U18906 (N_18906,N_17860,N_17947);
nor U18907 (N_18907,N_17938,N_18191);
and U18908 (N_18908,N_17818,N_18206);
and U18909 (N_18909,N_17612,N_18195);
or U18910 (N_18910,N_18240,N_17969);
and U18911 (N_18911,N_18066,N_17736);
nand U18912 (N_18912,N_18095,N_18088);
xnor U18913 (N_18913,N_17777,N_17977);
nand U18914 (N_18914,N_17932,N_18033);
and U18915 (N_18915,N_17731,N_18082);
and U18916 (N_18916,N_17723,N_17969);
nor U18917 (N_18917,N_17704,N_18005);
nand U18918 (N_18918,N_17794,N_18038);
xnor U18919 (N_18919,N_18010,N_17689);
nand U18920 (N_18920,N_18393,N_18356);
xnor U18921 (N_18921,N_18177,N_18164);
or U18922 (N_18922,N_18001,N_17882);
nand U18923 (N_18923,N_17971,N_18098);
nor U18924 (N_18924,N_17717,N_17724);
nand U18925 (N_18925,N_17867,N_18070);
nor U18926 (N_18926,N_18046,N_17865);
and U18927 (N_18927,N_17969,N_17849);
xor U18928 (N_18928,N_18132,N_18236);
xnor U18929 (N_18929,N_17974,N_17690);
nand U18930 (N_18930,N_18087,N_17818);
nand U18931 (N_18931,N_18017,N_17624);
or U18932 (N_18932,N_18046,N_18319);
or U18933 (N_18933,N_18053,N_17993);
xor U18934 (N_18934,N_17732,N_17741);
nor U18935 (N_18935,N_17935,N_17902);
and U18936 (N_18936,N_17685,N_17923);
nand U18937 (N_18937,N_18101,N_18129);
xnor U18938 (N_18938,N_18148,N_17783);
and U18939 (N_18939,N_17644,N_17739);
xnor U18940 (N_18940,N_18314,N_17871);
and U18941 (N_18941,N_18104,N_17677);
and U18942 (N_18942,N_18005,N_18200);
nand U18943 (N_18943,N_18238,N_18192);
or U18944 (N_18944,N_17650,N_17928);
xnor U18945 (N_18945,N_18188,N_17979);
and U18946 (N_18946,N_18267,N_18156);
or U18947 (N_18947,N_18347,N_18294);
and U18948 (N_18948,N_17940,N_18367);
nand U18949 (N_18949,N_18019,N_17984);
or U18950 (N_18950,N_17630,N_17839);
nand U18951 (N_18951,N_18271,N_18107);
nand U18952 (N_18952,N_18331,N_17665);
nor U18953 (N_18953,N_18372,N_17688);
xnor U18954 (N_18954,N_17937,N_18260);
nor U18955 (N_18955,N_18209,N_18082);
nor U18956 (N_18956,N_18119,N_17937);
and U18957 (N_18957,N_18202,N_18179);
nand U18958 (N_18958,N_18220,N_17947);
nand U18959 (N_18959,N_17701,N_18183);
and U18960 (N_18960,N_18027,N_18312);
nand U18961 (N_18961,N_17833,N_17799);
and U18962 (N_18962,N_17701,N_17645);
or U18963 (N_18963,N_17747,N_18267);
nor U18964 (N_18964,N_18146,N_17666);
nand U18965 (N_18965,N_18062,N_17625);
and U18966 (N_18966,N_18385,N_18300);
or U18967 (N_18967,N_18121,N_17876);
xor U18968 (N_18968,N_18151,N_18206);
and U18969 (N_18969,N_17826,N_17738);
nand U18970 (N_18970,N_17771,N_18046);
xor U18971 (N_18971,N_18220,N_18255);
and U18972 (N_18972,N_17874,N_18047);
xor U18973 (N_18973,N_18197,N_18295);
nor U18974 (N_18974,N_17641,N_18247);
and U18975 (N_18975,N_18077,N_17739);
or U18976 (N_18976,N_18155,N_18149);
and U18977 (N_18977,N_18308,N_18282);
nand U18978 (N_18978,N_18136,N_17930);
and U18979 (N_18979,N_18146,N_18055);
or U18980 (N_18980,N_18132,N_17609);
nand U18981 (N_18981,N_17856,N_18376);
nor U18982 (N_18982,N_17650,N_17957);
and U18983 (N_18983,N_18085,N_17861);
or U18984 (N_18984,N_18186,N_17681);
and U18985 (N_18985,N_17923,N_18097);
xnor U18986 (N_18986,N_18323,N_17774);
xnor U18987 (N_18987,N_17910,N_17695);
nor U18988 (N_18988,N_17965,N_17811);
and U18989 (N_18989,N_18307,N_17889);
nor U18990 (N_18990,N_17827,N_18314);
xor U18991 (N_18991,N_17831,N_18010);
nand U18992 (N_18992,N_18113,N_17958);
nor U18993 (N_18993,N_17851,N_17687);
nand U18994 (N_18994,N_17802,N_17650);
and U18995 (N_18995,N_17641,N_17758);
xnor U18996 (N_18996,N_18023,N_18160);
and U18997 (N_18997,N_17758,N_18382);
nand U18998 (N_18998,N_17810,N_17787);
nand U18999 (N_18999,N_18094,N_17854);
nand U19000 (N_19000,N_18259,N_18345);
or U19001 (N_19001,N_18312,N_17870);
xnor U19002 (N_19002,N_17940,N_18275);
nand U19003 (N_19003,N_17687,N_18340);
and U19004 (N_19004,N_18284,N_18060);
xnor U19005 (N_19005,N_17920,N_18157);
nand U19006 (N_19006,N_17924,N_17868);
or U19007 (N_19007,N_18125,N_18120);
xor U19008 (N_19008,N_17849,N_18273);
nand U19009 (N_19009,N_17814,N_18064);
or U19010 (N_19010,N_18363,N_17802);
nand U19011 (N_19011,N_18093,N_18242);
and U19012 (N_19012,N_17886,N_17776);
nor U19013 (N_19013,N_18238,N_18309);
nor U19014 (N_19014,N_17614,N_18354);
nor U19015 (N_19015,N_17992,N_17608);
and U19016 (N_19016,N_18020,N_17770);
nor U19017 (N_19017,N_18193,N_18126);
nor U19018 (N_19018,N_18290,N_18196);
nor U19019 (N_19019,N_18070,N_18126);
xnor U19020 (N_19020,N_17604,N_18036);
and U19021 (N_19021,N_18108,N_18243);
xor U19022 (N_19022,N_17709,N_17760);
or U19023 (N_19023,N_17930,N_17646);
nand U19024 (N_19024,N_18374,N_18171);
nor U19025 (N_19025,N_18264,N_18085);
nand U19026 (N_19026,N_17989,N_18364);
and U19027 (N_19027,N_17766,N_17610);
nand U19028 (N_19028,N_17735,N_17825);
nor U19029 (N_19029,N_18098,N_18257);
nand U19030 (N_19030,N_17689,N_18087);
and U19031 (N_19031,N_17999,N_18219);
xnor U19032 (N_19032,N_18248,N_17853);
and U19033 (N_19033,N_17709,N_18273);
nor U19034 (N_19034,N_17702,N_17740);
xor U19035 (N_19035,N_17876,N_17607);
and U19036 (N_19036,N_17807,N_17639);
or U19037 (N_19037,N_18069,N_18300);
nor U19038 (N_19038,N_18311,N_18048);
nor U19039 (N_19039,N_18248,N_18087);
xor U19040 (N_19040,N_18397,N_17627);
nor U19041 (N_19041,N_17826,N_18153);
nand U19042 (N_19042,N_17620,N_18016);
or U19043 (N_19043,N_18357,N_17930);
and U19044 (N_19044,N_18385,N_18130);
or U19045 (N_19045,N_18208,N_17858);
and U19046 (N_19046,N_18262,N_18368);
xnor U19047 (N_19047,N_17664,N_17953);
or U19048 (N_19048,N_18378,N_17772);
and U19049 (N_19049,N_18002,N_17786);
xnor U19050 (N_19050,N_18332,N_18126);
nand U19051 (N_19051,N_18191,N_18326);
nor U19052 (N_19052,N_18029,N_17917);
nand U19053 (N_19053,N_17798,N_17909);
xnor U19054 (N_19054,N_18240,N_17975);
xor U19055 (N_19055,N_18295,N_18081);
or U19056 (N_19056,N_18171,N_18274);
and U19057 (N_19057,N_17868,N_17938);
nand U19058 (N_19058,N_18006,N_17864);
nor U19059 (N_19059,N_17659,N_18032);
or U19060 (N_19060,N_18061,N_18166);
nand U19061 (N_19061,N_18290,N_18003);
nand U19062 (N_19062,N_17961,N_18255);
xnor U19063 (N_19063,N_18171,N_18087);
nand U19064 (N_19064,N_18243,N_17614);
or U19065 (N_19065,N_17752,N_18302);
or U19066 (N_19066,N_17947,N_17703);
nand U19067 (N_19067,N_18288,N_17683);
or U19068 (N_19068,N_18286,N_17692);
nand U19069 (N_19069,N_18372,N_18200);
nand U19070 (N_19070,N_17944,N_18218);
nor U19071 (N_19071,N_17621,N_17614);
nor U19072 (N_19072,N_18159,N_18102);
and U19073 (N_19073,N_17789,N_17692);
or U19074 (N_19074,N_18193,N_17605);
xnor U19075 (N_19075,N_17860,N_17792);
xnor U19076 (N_19076,N_18058,N_18330);
and U19077 (N_19077,N_18357,N_18037);
nand U19078 (N_19078,N_18070,N_18204);
nand U19079 (N_19079,N_18169,N_17924);
xnor U19080 (N_19080,N_18035,N_18239);
nand U19081 (N_19081,N_18217,N_17809);
xor U19082 (N_19082,N_18150,N_17645);
xor U19083 (N_19083,N_17605,N_17694);
nor U19084 (N_19084,N_18001,N_17707);
nand U19085 (N_19085,N_18304,N_18100);
xor U19086 (N_19086,N_18000,N_18098);
and U19087 (N_19087,N_17848,N_17934);
xor U19088 (N_19088,N_17985,N_18012);
nand U19089 (N_19089,N_17976,N_17841);
and U19090 (N_19090,N_18321,N_18355);
nor U19091 (N_19091,N_18137,N_18300);
xor U19092 (N_19092,N_17904,N_18162);
nor U19093 (N_19093,N_18010,N_17722);
or U19094 (N_19094,N_17657,N_18322);
and U19095 (N_19095,N_18125,N_17695);
or U19096 (N_19096,N_17816,N_17985);
xor U19097 (N_19097,N_17932,N_18294);
nor U19098 (N_19098,N_17839,N_18218);
nand U19099 (N_19099,N_18364,N_17962);
nand U19100 (N_19100,N_18000,N_17953);
nor U19101 (N_19101,N_17735,N_18181);
and U19102 (N_19102,N_18280,N_18016);
and U19103 (N_19103,N_18308,N_18190);
or U19104 (N_19104,N_17620,N_18274);
xnor U19105 (N_19105,N_18274,N_17769);
nor U19106 (N_19106,N_17620,N_17915);
nor U19107 (N_19107,N_18259,N_17986);
or U19108 (N_19108,N_17875,N_18378);
nand U19109 (N_19109,N_17957,N_17836);
or U19110 (N_19110,N_18125,N_17880);
nand U19111 (N_19111,N_17884,N_18339);
xor U19112 (N_19112,N_18382,N_18289);
and U19113 (N_19113,N_17995,N_18057);
nor U19114 (N_19114,N_18125,N_17854);
and U19115 (N_19115,N_17613,N_17965);
nor U19116 (N_19116,N_17617,N_18109);
nor U19117 (N_19117,N_18011,N_18118);
and U19118 (N_19118,N_17826,N_17926);
xnor U19119 (N_19119,N_18358,N_18082);
nand U19120 (N_19120,N_18370,N_17637);
or U19121 (N_19121,N_17831,N_17838);
nand U19122 (N_19122,N_17629,N_18378);
and U19123 (N_19123,N_18117,N_17808);
xor U19124 (N_19124,N_18205,N_18246);
xnor U19125 (N_19125,N_18343,N_18264);
or U19126 (N_19126,N_18133,N_17948);
nor U19127 (N_19127,N_18334,N_18365);
or U19128 (N_19128,N_18291,N_17770);
and U19129 (N_19129,N_18236,N_18067);
nand U19130 (N_19130,N_17902,N_17724);
nor U19131 (N_19131,N_17685,N_18097);
xnor U19132 (N_19132,N_17838,N_18142);
nor U19133 (N_19133,N_18025,N_18169);
nand U19134 (N_19134,N_18098,N_17982);
and U19135 (N_19135,N_17770,N_18362);
or U19136 (N_19136,N_18187,N_18224);
nand U19137 (N_19137,N_17953,N_18018);
nor U19138 (N_19138,N_18357,N_18242);
nor U19139 (N_19139,N_17704,N_18271);
xor U19140 (N_19140,N_18163,N_17989);
or U19141 (N_19141,N_18179,N_17818);
nand U19142 (N_19142,N_17863,N_18207);
or U19143 (N_19143,N_17720,N_18375);
nand U19144 (N_19144,N_18014,N_18310);
and U19145 (N_19145,N_17879,N_17689);
xnor U19146 (N_19146,N_18325,N_18014);
and U19147 (N_19147,N_18099,N_17864);
nand U19148 (N_19148,N_17859,N_18092);
nor U19149 (N_19149,N_18173,N_18293);
or U19150 (N_19150,N_18091,N_18030);
nand U19151 (N_19151,N_18310,N_17618);
nor U19152 (N_19152,N_18199,N_17965);
nor U19153 (N_19153,N_18341,N_18004);
or U19154 (N_19154,N_17703,N_17764);
xnor U19155 (N_19155,N_17867,N_17943);
nand U19156 (N_19156,N_17989,N_17973);
and U19157 (N_19157,N_18189,N_18397);
nor U19158 (N_19158,N_18232,N_17663);
or U19159 (N_19159,N_17649,N_18222);
xnor U19160 (N_19160,N_18214,N_18340);
nand U19161 (N_19161,N_17696,N_17641);
xnor U19162 (N_19162,N_17775,N_17792);
or U19163 (N_19163,N_17853,N_18227);
and U19164 (N_19164,N_18228,N_17678);
or U19165 (N_19165,N_18247,N_18217);
xor U19166 (N_19166,N_17727,N_17792);
xor U19167 (N_19167,N_18361,N_17757);
and U19168 (N_19168,N_17750,N_17772);
or U19169 (N_19169,N_18155,N_18175);
nor U19170 (N_19170,N_18119,N_18296);
nor U19171 (N_19171,N_17859,N_17888);
xor U19172 (N_19172,N_18145,N_18364);
xor U19173 (N_19173,N_18236,N_17874);
or U19174 (N_19174,N_18296,N_18102);
xnor U19175 (N_19175,N_18140,N_17832);
or U19176 (N_19176,N_18262,N_18198);
nor U19177 (N_19177,N_17634,N_17835);
xnor U19178 (N_19178,N_18202,N_17862);
and U19179 (N_19179,N_17745,N_18049);
and U19180 (N_19180,N_17837,N_18270);
nand U19181 (N_19181,N_17787,N_17734);
or U19182 (N_19182,N_17987,N_18325);
nand U19183 (N_19183,N_18228,N_17693);
and U19184 (N_19184,N_17980,N_18060);
nand U19185 (N_19185,N_18316,N_17839);
nor U19186 (N_19186,N_18282,N_17798);
nor U19187 (N_19187,N_18018,N_18364);
and U19188 (N_19188,N_17679,N_18302);
xor U19189 (N_19189,N_17826,N_17965);
and U19190 (N_19190,N_18132,N_18142);
or U19191 (N_19191,N_18078,N_18239);
or U19192 (N_19192,N_18166,N_18213);
xor U19193 (N_19193,N_18019,N_18081);
nand U19194 (N_19194,N_17813,N_18349);
nor U19195 (N_19195,N_17811,N_18199);
nor U19196 (N_19196,N_17639,N_17883);
nand U19197 (N_19197,N_18350,N_17854);
nor U19198 (N_19198,N_18117,N_17840);
or U19199 (N_19199,N_18299,N_18295);
nor U19200 (N_19200,N_18951,N_18822);
and U19201 (N_19201,N_18410,N_18414);
or U19202 (N_19202,N_18767,N_19180);
and U19203 (N_19203,N_18583,N_19034);
or U19204 (N_19204,N_18768,N_18470);
or U19205 (N_19205,N_18983,N_18755);
nor U19206 (N_19206,N_18685,N_19158);
xnor U19207 (N_19207,N_18436,N_18918);
nor U19208 (N_19208,N_18475,N_18692);
and U19209 (N_19209,N_19164,N_18856);
xor U19210 (N_19210,N_19018,N_18878);
xnor U19211 (N_19211,N_18844,N_18502);
xnor U19212 (N_19212,N_18525,N_18834);
nand U19213 (N_19213,N_18461,N_18819);
nand U19214 (N_19214,N_18907,N_19162);
xnor U19215 (N_19215,N_19097,N_18828);
xnor U19216 (N_19216,N_18859,N_19028);
nor U19217 (N_19217,N_18779,N_18508);
xnor U19218 (N_19218,N_19058,N_18809);
or U19219 (N_19219,N_19157,N_18412);
xnor U19220 (N_19220,N_18987,N_18492);
nor U19221 (N_19221,N_18512,N_18625);
nand U19222 (N_19222,N_18615,N_18801);
nor U19223 (N_19223,N_19138,N_19091);
nor U19224 (N_19224,N_18602,N_18686);
and U19225 (N_19225,N_19096,N_18654);
nor U19226 (N_19226,N_19056,N_19196);
nor U19227 (N_19227,N_18810,N_18541);
xnor U19228 (N_19228,N_19137,N_18407);
xor U19229 (N_19229,N_18683,N_18961);
nor U19230 (N_19230,N_18751,N_19008);
or U19231 (N_19231,N_18981,N_19147);
nand U19232 (N_19232,N_19133,N_18415);
xor U19233 (N_19233,N_18714,N_18669);
nor U19234 (N_19234,N_19176,N_18406);
or U19235 (N_19235,N_19057,N_19054);
nor U19236 (N_19236,N_19154,N_18974);
xor U19237 (N_19237,N_18857,N_18617);
xor U19238 (N_19238,N_18902,N_18549);
or U19239 (N_19239,N_18500,N_18531);
nor U19240 (N_19240,N_18404,N_19140);
and U19241 (N_19241,N_18786,N_18627);
and U19242 (N_19242,N_18621,N_18554);
nor U19243 (N_19243,N_18506,N_18573);
nor U19244 (N_19244,N_18558,N_18725);
xnor U19245 (N_19245,N_18874,N_18579);
xor U19246 (N_19246,N_18559,N_18452);
and U19247 (N_19247,N_18928,N_18562);
or U19248 (N_19248,N_18718,N_18776);
nor U19249 (N_19249,N_18504,N_19110);
or U19250 (N_19250,N_18953,N_19111);
and U19251 (N_19251,N_18803,N_19159);
or U19252 (N_19252,N_18816,N_18798);
nand U19253 (N_19253,N_18973,N_18726);
xnor U19254 (N_19254,N_18478,N_18422);
and U19255 (N_19255,N_19193,N_18713);
nor U19256 (N_19256,N_19043,N_18547);
nor U19257 (N_19257,N_18588,N_19168);
or U19258 (N_19258,N_18442,N_18548);
or U19259 (N_19259,N_18870,N_18454);
xnor U19260 (N_19260,N_18693,N_19001);
nand U19261 (N_19261,N_18841,N_18462);
or U19262 (N_19262,N_19003,N_18971);
xnor U19263 (N_19263,N_18451,N_18457);
nand U19264 (N_19264,N_18599,N_18840);
nand U19265 (N_19265,N_19032,N_18425);
nand U19266 (N_19266,N_18688,N_18724);
xor U19267 (N_19267,N_18514,N_19134);
or U19268 (N_19268,N_18813,N_18804);
nand U19269 (N_19269,N_18849,N_18572);
xor U19270 (N_19270,N_18965,N_18649);
nor U19271 (N_19271,N_18523,N_18674);
xnor U19272 (N_19272,N_18889,N_18790);
or U19273 (N_19273,N_18517,N_18424);
xnor U19274 (N_19274,N_18835,N_19095);
nand U19275 (N_19275,N_18642,N_18533);
nand U19276 (N_19276,N_18708,N_18966);
xnor U19277 (N_19277,N_18851,N_18734);
xor U19278 (N_19278,N_18494,N_18991);
and U19279 (N_19279,N_18619,N_18431);
and U19280 (N_19280,N_18493,N_19092);
xnor U19281 (N_19281,N_18648,N_18952);
nor U19282 (N_19282,N_18926,N_18895);
xnor U19283 (N_19283,N_19083,N_18882);
xnor U19284 (N_19284,N_18663,N_19106);
nor U19285 (N_19285,N_19173,N_18439);
or U19286 (N_19286,N_18568,N_18632);
nor U19287 (N_19287,N_19124,N_18984);
or U19288 (N_19288,N_18421,N_18985);
or U19289 (N_19289,N_18400,N_18789);
or U19290 (N_19290,N_18799,N_18885);
and U19291 (N_19291,N_18656,N_19149);
nor U19292 (N_19292,N_18694,N_18887);
nand U19293 (N_19293,N_18581,N_18497);
and U19294 (N_19294,N_19172,N_19100);
nor U19295 (N_19295,N_19181,N_18995);
xnor U19296 (N_19296,N_18879,N_18438);
nand U19297 (N_19297,N_18680,N_18775);
or U19298 (N_19298,N_18975,N_19114);
nor U19299 (N_19299,N_18900,N_18997);
or U19300 (N_19300,N_18495,N_18795);
or U19301 (N_19301,N_18947,N_18608);
nor U19302 (N_19302,N_18867,N_18922);
nor U19303 (N_19303,N_18655,N_18426);
and U19304 (N_19304,N_19152,N_19045);
or U19305 (N_19305,N_18938,N_18658);
nand U19306 (N_19306,N_18488,N_18510);
and U19307 (N_19307,N_18629,N_18905);
xnor U19308 (N_19308,N_18535,N_18700);
nand U19309 (N_19309,N_18865,N_18802);
nor U19310 (N_19310,N_18657,N_19026);
and U19311 (N_19311,N_19109,N_18881);
nand U19312 (N_19312,N_18910,N_18758);
xnor U19313 (N_19313,N_18782,N_18667);
nand U19314 (N_19314,N_18593,N_19025);
and U19315 (N_19315,N_18964,N_18797);
and U19316 (N_19316,N_18747,N_18890);
and U19317 (N_19317,N_18769,N_18532);
xnor U19318 (N_19318,N_18996,N_18827);
nand U19319 (N_19319,N_18456,N_18591);
or U19320 (N_19320,N_18853,N_19126);
nand U19321 (N_19321,N_18862,N_19077);
and U19322 (N_19322,N_19117,N_19103);
nand U19323 (N_19323,N_18759,N_18679);
or U19324 (N_19324,N_19145,N_18706);
and U19325 (N_19325,N_18537,N_18587);
and U19326 (N_19326,N_18603,N_18576);
or U19327 (N_19327,N_19085,N_18528);
xnor U19328 (N_19328,N_18556,N_18899);
nor U19329 (N_19329,N_19087,N_19007);
nand U19330 (N_19330,N_18746,N_18444);
nand U19331 (N_19331,N_18994,N_18678);
and U19332 (N_19332,N_19165,N_19064);
and U19333 (N_19333,N_18972,N_18717);
and U19334 (N_19334,N_18761,N_18875);
xnor U19335 (N_19335,N_18571,N_18771);
nand U19336 (N_19336,N_19023,N_19141);
xnor U19337 (N_19337,N_18474,N_19153);
or U19338 (N_19338,N_18671,N_18607);
and U19339 (N_19339,N_18871,N_19121);
xnor U19340 (N_19340,N_18785,N_18699);
nand U19341 (N_19341,N_18652,N_18850);
or U19342 (N_19342,N_18770,N_18969);
and U19343 (N_19343,N_18565,N_19131);
and U19344 (N_19344,N_18557,N_18943);
or U19345 (N_19345,N_19189,N_18858);
or U19346 (N_19346,N_18598,N_18423);
and U19347 (N_19347,N_18466,N_19136);
nand U19348 (N_19348,N_18638,N_18904);
nor U19349 (N_19349,N_18784,N_18605);
and U19350 (N_19350,N_18703,N_18992);
and U19351 (N_19351,N_18990,N_19199);
or U19352 (N_19352,N_18580,N_18516);
or U19353 (N_19353,N_18518,N_19166);
and U19354 (N_19354,N_18854,N_19127);
and U19355 (N_19355,N_19042,N_18595);
or U19356 (N_19356,N_18738,N_18814);
xor U19357 (N_19357,N_19115,N_18676);
nor U19358 (N_19358,N_19093,N_18846);
and U19359 (N_19359,N_18723,N_19175);
and U19360 (N_19360,N_18869,N_18852);
nand U19361 (N_19361,N_19013,N_18940);
xor U19362 (N_19362,N_19148,N_19021);
nor U19363 (N_19363,N_18949,N_18728);
nand U19364 (N_19364,N_19129,N_18622);
or U19365 (N_19365,N_19050,N_18644);
nor U19366 (N_19366,N_19068,N_19036);
and U19367 (N_19367,N_19030,N_18578);
and U19368 (N_19368,N_18727,N_18513);
xor U19369 (N_19369,N_18886,N_18712);
and U19370 (N_19370,N_19143,N_19182);
nand U19371 (N_19371,N_18760,N_18428);
nor U19372 (N_19372,N_18756,N_19119);
or U19373 (N_19373,N_18752,N_19070);
and U19374 (N_19374,N_18536,N_18732);
nor U19375 (N_19375,N_18818,N_19123);
xor U19376 (N_19376,N_19020,N_18821);
xor U19377 (N_19377,N_18893,N_18610);
xnor U19378 (N_19378,N_18957,N_18464);
xnor U19379 (N_19379,N_18721,N_19192);
or U19380 (N_19380,N_19027,N_18710);
or U19381 (N_19381,N_18577,N_18979);
and U19382 (N_19382,N_18978,N_19055);
nand U19383 (N_19383,N_18792,N_18635);
or U19384 (N_19384,N_19151,N_18939);
and U19385 (N_19385,N_18958,N_18418);
nand U19386 (N_19386,N_18689,N_18673);
and U19387 (N_19387,N_18815,N_19128);
xor U19388 (N_19388,N_19012,N_19075);
and U19389 (N_19389,N_18403,N_18986);
xor U19390 (N_19390,N_18491,N_18794);
nand U19391 (N_19391,N_18805,N_18730);
and U19392 (N_19392,N_18582,N_19051);
or U19393 (N_19393,N_18682,N_18677);
nand U19394 (N_19394,N_18561,N_19074);
xnor U19395 (N_19395,N_18715,N_18914);
nor U19396 (N_19396,N_18783,N_18921);
nand U19397 (N_19397,N_18781,N_18539);
xnor U19398 (N_19398,N_18611,N_18477);
nor U19399 (N_19399,N_18405,N_19048);
or U19400 (N_19400,N_18932,N_18839);
or U19401 (N_19401,N_18778,N_19065);
nor U19402 (N_19402,N_18954,N_18808);
xor U19403 (N_19403,N_18884,N_18735);
and U19404 (N_19404,N_18944,N_18590);
or U19405 (N_19405,N_18567,N_19113);
and U19406 (N_19406,N_19061,N_19073);
or U19407 (N_19407,N_19039,N_19069);
nand U19408 (N_19408,N_18503,N_18913);
or U19409 (N_19409,N_19120,N_18936);
nand U19410 (N_19410,N_19104,N_18534);
and U19411 (N_19411,N_18634,N_19053);
or U19412 (N_19412,N_18524,N_18681);
xor U19413 (N_19413,N_18742,N_18662);
xnor U19414 (N_19414,N_18962,N_18482);
xnor U19415 (N_19415,N_18519,N_18811);
and U19416 (N_19416,N_19002,N_19098);
xnor U19417 (N_19417,N_18739,N_18707);
nor U19418 (N_19418,N_18527,N_18472);
nand U19419 (N_19419,N_19198,N_18897);
nand U19420 (N_19420,N_18485,N_18763);
nand U19421 (N_19421,N_19170,N_18906);
and U19422 (N_19422,N_19040,N_18569);
xnor U19423 (N_19423,N_18695,N_19000);
nor U19424 (N_19424,N_18465,N_18817);
nand U19425 (N_19425,N_18909,N_18765);
and U19426 (N_19426,N_18976,N_18793);
nor U19427 (N_19427,N_18522,N_18823);
nor U19428 (N_19428,N_18645,N_18468);
or U19429 (N_19429,N_18480,N_18570);
or U19430 (N_19430,N_18848,N_19035);
nand U19431 (N_19431,N_18665,N_18753);
nor U19432 (N_19432,N_18633,N_18498);
and U19433 (N_19433,N_18540,N_18545);
nand U19434 (N_19434,N_18427,N_18930);
or U19435 (N_19435,N_18653,N_19178);
nor U19436 (N_19436,N_18743,N_18483);
xnor U19437 (N_19437,N_18993,N_18650);
or U19438 (N_19438,N_19010,N_18529);
xnor U19439 (N_19439,N_18824,N_19094);
nand U19440 (N_19440,N_19011,N_19088);
or U19441 (N_19441,N_18659,N_18505);
nand U19442 (N_19442,N_19169,N_18417);
and U19443 (N_19443,N_18484,N_18443);
or U19444 (N_19444,N_19185,N_19139);
nor U19445 (N_19445,N_18604,N_18898);
nor U19446 (N_19446,N_19122,N_18908);
xor U19447 (N_19447,N_19190,N_18589);
nand U19448 (N_19448,N_18737,N_18521);
nand U19449 (N_19449,N_19132,N_19052);
nor U19450 (N_19450,N_18489,N_18866);
and U19451 (N_19451,N_19084,N_18575);
xor U19452 (N_19452,N_18998,N_18740);
nor U19453 (N_19453,N_18460,N_19031);
nand U19454 (N_19454,N_19197,N_18458);
or U19455 (N_19455,N_18704,N_19105);
and U19456 (N_19456,N_19086,N_19072);
or U19457 (N_19457,N_19099,N_19160);
and U19458 (N_19458,N_18960,N_19016);
nand U19459 (N_19459,N_18845,N_18453);
nand U19460 (N_19460,N_18956,N_18586);
or U19461 (N_19461,N_18630,N_19101);
nand U19462 (N_19462,N_18419,N_18511);
nand U19463 (N_19463,N_18507,N_18892);
or U19464 (N_19464,N_18711,N_19029);
nand U19465 (N_19465,N_19102,N_18748);
xor U19466 (N_19466,N_18744,N_19177);
and U19467 (N_19467,N_18968,N_19179);
xor U19468 (N_19468,N_18433,N_19037);
and U19469 (N_19469,N_18698,N_18788);
xor U19470 (N_19470,N_18796,N_18479);
nor U19471 (N_19471,N_18925,N_18825);
or U19472 (N_19472,N_18432,N_18830);
and U19473 (N_19473,N_18876,N_18600);
xor U19474 (N_19474,N_18820,N_18731);
and U19475 (N_19475,N_18463,N_18501);
or U19476 (N_19476,N_18613,N_18550);
and U19477 (N_19477,N_18745,N_19017);
and U19478 (N_19478,N_18977,N_18896);
nor U19479 (N_19479,N_18441,N_18481);
or U19480 (N_19480,N_18409,N_18620);
or U19481 (N_19481,N_18551,N_18774);
nor U19482 (N_19482,N_19076,N_18408);
xor U19483 (N_19483,N_19135,N_19014);
nand U19484 (N_19484,N_18469,N_18437);
or U19485 (N_19485,N_18413,N_19183);
and U19486 (N_19486,N_18891,N_18563);
or U19487 (N_19487,N_18883,N_18486);
nor U19488 (N_19488,N_18446,N_18915);
or U19489 (N_19489,N_18863,N_18691);
xnor U19490 (N_19490,N_18935,N_18920);
xnor U19491 (N_19491,N_18919,N_18872);
and U19492 (N_19492,N_19082,N_18754);
or U19493 (N_19493,N_19004,N_18912);
nand U19494 (N_19494,N_18709,N_18440);
or U19495 (N_19495,N_18661,N_18459);
nor U19496 (N_19496,N_19015,N_19118);
nand U19497 (N_19497,N_19019,N_18526);
nand U19498 (N_19498,N_18660,N_18624);
or U19499 (N_19499,N_18684,N_18664);
or U19500 (N_19500,N_18670,N_18829);
and U19501 (N_19501,N_18955,N_19184);
nor U19502 (N_19502,N_18473,N_18594);
xor U19503 (N_19503,N_19108,N_18946);
nand U19504 (N_19504,N_19022,N_18948);
nor U19505 (N_19505,N_19063,N_18945);
xnor U19506 (N_19506,N_18628,N_18911);
nor U19507 (N_19507,N_18592,N_18402);
nor U19508 (N_19508,N_18888,N_19080);
and U19509 (N_19509,N_18842,N_18564);
nor U19510 (N_19510,N_18942,N_18530);
and U19511 (N_19511,N_18807,N_18675);
nand U19512 (N_19512,N_18941,N_18980);
xor U19513 (N_19513,N_18959,N_18988);
nor U19514 (N_19514,N_18448,N_18812);
nand U19515 (N_19515,N_18836,N_18429);
nand U19516 (N_19516,N_19062,N_18800);
nand U19517 (N_19517,N_19194,N_19090);
and U19518 (N_19518,N_18719,N_18733);
nand U19519 (N_19519,N_18416,N_18931);
nand U19520 (N_19520,N_19060,N_18705);
xnor U19521 (N_19521,N_18640,N_18467);
or U19522 (N_19522,N_18647,N_19044);
nand U19523 (N_19523,N_18546,N_18773);
nand U19524 (N_19524,N_18687,N_18596);
or U19525 (N_19525,N_18791,N_18455);
xor U19526 (N_19526,N_19038,N_19195);
or U19527 (N_19527,N_19078,N_18741);
nor U19528 (N_19528,N_19188,N_18543);
or U19529 (N_19529,N_19144,N_18832);
nand U19530 (N_19530,N_18449,N_19081);
and U19531 (N_19531,N_18787,N_18766);
and U19532 (N_19532,N_18445,N_18702);
nor U19533 (N_19533,N_18970,N_18873);
nand U19534 (N_19534,N_19047,N_19033);
and U19535 (N_19535,N_18777,N_18762);
and U19536 (N_19536,N_18609,N_18499);
and U19537 (N_19537,N_19156,N_18894);
nor U19538 (N_19538,N_19049,N_18950);
or U19539 (N_19539,N_18967,N_18927);
and U19540 (N_19540,N_18538,N_18636);
nor U19541 (N_19541,N_18933,N_19161);
nor U19542 (N_19542,N_19112,N_19187);
nand U19543 (N_19543,N_18560,N_18544);
or U19544 (N_19544,N_19167,N_18574);
xnor U19545 (N_19545,N_19066,N_19163);
nor U19546 (N_19546,N_18618,N_18716);
or U19547 (N_19547,N_18838,N_18729);
xor U19548 (N_19548,N_18566,N_18606);
xnor U19549 (N_19549,N_19046,N_18903);
nor U19550 (N_19550,N_18916,N_18639);
nor U19551 (N_19551,N_18435,N_18780);
and U19552 (N_19552,N_19009,N_18757);
nor U19553 (N_19553,N_18772,N_19071);
and U19554 (N_19554,N_18847,N_19130);
xor U19555 (N_19555,N_18929,N_18471);
nor U19556 (N_19556,N_18989,N_18999);
nand U19557 (N_19557,N_18401,N_18651);
nor U19558 (N_19558,N_18982,N_19079);
or U19559 (N_19559,N_18934,N_18631);
xnor U19560 (N_19560,N_18963,N_18806);
nand U19561 (N_19561,N_18668,N_19191);
and U19562 (N_19562,N_18696,N_18750);
xor U19563 (N_19563,N_18860,N_18552);
and U19564 (N_19564,N_19146,N_18623);
nor U19565 (N_19565,N_18880,N_19155);
and U19566 (N_19566,N_18720,N_18690);
xor U19567 (N_19567,N_18447,N_18701);
nand U19568 (N_19568,N_18937,N_19041);
nand U19569 (N_19569,N_18601,N_18584);
nor U19570 (N_19570,N_18641,N_18555);
nor U19571 (N_19571,N_18901,N_18612);
nor U19572 (N_19572,N_18450,N_18672);
or U19573 (N_19573,N_18515,N_18487);
or U19574 (N_19574,N_18868,N_18855);
or U19575 (N_19575,N_19171,N_18833);
xnor U19576 (N_19576,N_18585,N_18826);
nor U19577 (N_19577,N_18749,N_18626);
xor U19578 (N_19578,N_18616,N_18434);
and U19579 (N_19579,N_18597,N_18643);
or U19580 (N_19580,N_19005,N_18697);
nor U19581 (N_19581,N_18837,N_18923);
or U19582 (N_19582,N_18831,N_19089);
xnor U19583 (N_19583,N_18861,N_19006);
and U19584 (N_19584,N_19150,N_18614);
or U19585 (N_19585,N_19107,N_18637);
and U19586 (N_19586,N_19059,N_18917);
or U19587 (N_19587,N_18490,N_18666);
nand U19588 (N_19588,N_18764,N_19116);
nor U19589 (N_19589,N_18411,N_19024);
or U19590 (N_19590,N_18646,N_19067);
and U19591 (N_19591,N_18877,N_18843);
and U19592 (N_19592,N_18924,N_18553);
nor U19593 (N_19593,N_19186,N_19125);
or U19594 (N_19594,N_19174,N_18520);
and U19595 (N_19595,N_18509,N_18542);
nor U19596 (N_19596,N_18736,N_19142);
xnor U19597 (N_19597,N_18722,N_18430);
xnor U19598 (N_19598,N_18476,N_18420);
and U19599 (N_19599,N_18864,N_18496);
and U19600 (N_19600,N_18838,N_19184);
nand U19601 (N_19601,N_18646,N_18902);
nor U19602 (N_19602,N_18517,N_18572);
nor U19603 (N_19603,N_18975,N_18655);
nand U19604 (N_19604,N_18566,N_18796);
or U19605 (N_19605,N_18817,N_18998);
or U19606 (N_19606,N_18622,N_18651);
nor U19607 (N_19607,N_18478,N_18923);
and U19608 (N_19608,N_18497,N_18554);
or U19609 (N_19609,N_18619,N_18633);
or U19610 (N_19610,N_18704,N_19196);
and U19611 (N_19611,N_18952,N_19149);
and U19612 (N_19612,N_18891,N_18404);
or U19613 (N_19613,N_18636,N_18537);
and U19614 (N_19614,N_18475,N_19150);
or U19615 (N_19615,N_19168,N_18560);
and U19616 (N_19616,N_19172,N_18510);
nand U19617 (N_19617,N_18486,N_18705);
nor U19618 (N_19618,N_18735,N_19108);
or U19619 (N_19619,N_18765,N_18714);
nand U19620 (N_19620,N_19126,N_19060);
nand U19621 (N_19621,N_18902,N_18664);
and U19622 (N_19622,N_19164,N_18568);
nand U19623 (N_19623,N_18836,N_18944);
or U19624 (N_19624,N_19104,N_18558);
and U19625 (N_19625,N_18779,N_18588);
nand U19626 (N_19626,N_18775,N_18494);
nor U19627 (N_19627,N_18842,N_19196);
or U19628 (N_19628,N_18902,N_18657);
and U19629 (N_19629,N_18567,N_18972);
or U19630 (N_19630,N_18751,N_19132);
or U19631 (N_19631,N_19190,N_19012);
xnor U19632 (N_19632,N_18918,N_19188);
or U19633 (N_19633,N_19121,N_19024);
nor U19634 (N_19634,N_18565,N_18898);
xnor U19635 (N_19635,N_18562,N_18812);
and U19636 (N_19636,N_18484,N_19068);
or U19637 (N_19637,N_19059,N_18520);
nand U19638 (N_19638,N_19037,N_18864);
nor U19639 (N_19639,N_18451,N_18654);
or U19640 (N_19640,N_18527,N_18463);
xnor U19641 (N_19641,N_18476,N_19127);
xnor U19642 (N_19642,N_18600,N_18880);
nand U19643 (N_19643,N_18892,N_19145);
nor U19644 (N_19644,N_18745,N_19029);
nand U19645 (N_19645,N_19185,N_18504);
nor U19646 (N_19646,N_18601,N_18854);
nor U19647 (N_19647,N_18786,N_18953);
xnor U19648 (N_19648,N_18496,N_19103);
nor U19649 (N_19649,N_18825,N_19178);
xor U19650 (N_19650,N_18655,N_18645);
nand U19651 (N_19651,N_18860,N_18965);
xor U19652 (N_19652,N_18505,N_18460);
nor U19653 (N_19653,N_18514,N_18438);
or U19654 (N_19654,N_19171,N_18463);
and U19655 (N_19655,N_18598,N_18461);
xor U19656 (N_19656,N_19055,N_18934);
xor U19657 (N_19657,N_18994,N_18879);
nand U19658 (N_19658,N_18408,N_18538);
xor U19659 (N_19659,N_18759,N_18429);
or U19660 (N_19660,N_18603,N_19169);
nand U19661 (N_19661,N_18805,N_18506);
nand U19662 (N_19662,N_19055,N_18698);
nand U19663 (N_19663,N_18551,N_18634);
or U19664 (N_19664,N_18488,N_18505);
xor U19665 (N_19665,N_18499,N_18850);
xor U19666 (N_19666,N_18643,N_18756);
xnor U19667 (N_19667,N_18955,N_18710);
or U19668 (N_19668,N_18591,N_18563);
or U19669 (N_19669,N_18776,N_18466);
nand U19670 (N_19670,N_18968,N_18916);
and U19671 (N_19671,N_19047,N_19069);
and U19672 (N_19672,N_19083,N_18779);
or U19673 (N_19673,N_19015,N_19132);
nand U19674 (N_19674,N_18519,N_18455);
and U19675 (N_19675,N_18604,N_18537);
nand U19676 (N_19676,N_18841,N_19174);
xnor U19677 (N_19677,N_19188,N_18947);
nand U19678 (N_19678,N_18713,N_18995);
xor U19679 (N_19679,N_18695,N_18687);
and U19680 (N_19680,N_19159,N_19009);
nor U19681 (N_19681,N_19157,N_18407);
nand U19682 (N_19682,N_18901,N_19103);
nand U19683 (N_19683,N_18913,N_19112);
xnor U19684 (N_19684,N_18699,N_18802);
or U19685 (N_19685,N_19023,N_18857);
or U19686 (N_19686,N_18586,N_18831);
and U19687 (N_19687,N_18882,N_18826);
or U19688 (N_19688,N_18559,N_18631);
xor U19689 (N_19689,N_18541,N_18634);
nand U19690 (N_19690,N_18593,N_18872);
or U19691 (N_19691,N_18820,N_18537);
and U19692 (N_19692,N_18584,N_18677);
xor U19693 (N_19693,N_18783,N_18959);
or U19694 (N_19694,N_18417,N_18726);
nand U19695 (N_19695,N_18510,N_18786);
or U19696 (N_19696,N_18940,N_18495);
or U19697 (N_19697,N_18830,N_18747);
or U19698 (N_19698,N_18756,N_18646);
nor U19699 (N_19699,N_18804,N_18552);
nor U19700 (N_19700,N_19140,N_19035);
nor U19701 (N_19701,N_18452,N_18489);
or U19702 (N_19702,N_19184,N_19021);
nor U19703 (N_19703,N_18428,N_19135);
nand U19704 (N_19704,N_18861,N_18463);
nor U19705 (N_19705,N_18696,N_18994);
xor U19706 (N_19706,N_18965,N_18459);
or U19707 (N_19707,N_18767,N_18934);
nor U19708 (N_19708,N_18802,N_18639);
xnor U19709 (N_19709,N_19115,N_18952);
nand U19710 (N_19710,N_19142,N_18983);
nor U19711 (N_19711,N_18743,N_19122);
nor U19712 (N_19712,N_19193,N_18700);
or U19713 (N_19713,N_18679,N_19080);
and U19714 (N_19714,N_18540,N_18562);
or U19715 (N_19715,N_18548,N_18917);
or U19716 (N_19716,N_18506,N_18708);
nor U19717 (N_19717,N_18849,N_18992);
nand U19718 (N_19718,N_18731,N_18607);
nor U19719 (N_19719,N_18562,N_19079);
xor U19720 (N_19720,N_18775,N_18792);
xor U19721 (N_19721,N_19036,N_18987);
and U19722 (N_19722,N_19051,N_18626);
or U19723 (N_19723,N_18575,N_18505);
and U19724 (N_19724,N_18930,N_19148);
nor U19725 (N_19725,N_18835,N_18767);
nor U19726 (N_19726,N_18983,N_18471);
or U19727 (N_19727,N_19043,N_18722);
xor U19728 (N_19728,N_18829,N_18801);
or U19729 (N_19729,N_18417,N_18601);
nor U19730 (N_19730,N_18697,N_19146);
or U19731 (N_19731,N_19156,N_18927);
xnor U19732 (N_19732,N_18480,N_18988);
xor U19733 (N_19733,N_18625,N_19119);
nor U19734 (N_19734,N_18983,N_18443);
nand U19735 (N_19735,N_18411,N_18629);
and U19736 (N_19736,N_19010,N_19190);
or U19737 (N_19737,N_18948,N_19085);
nand U19738 (N_19738,N_18788,N_18529);
xor U19739 (N_19739,N_19047,N_19073);
and U19740 (N_19740,N_18420,N_19104);
xor U19741 (N_19741,N_18586,N_18418);
nor U19742 (N_19742,N_18878,N_18866);
nand U19743 (N_19743,N_18628,N_19040);
nor U19744 (N_19744,N_19038,N_18917);
nor U19745 (N_19745,N_19160,N_19101);
nor U19746 (N_19746,N_18836,N_18677);
nor U19747 (N_19747,N_18872,N_19099);
or U19748 (N_19748,N_18754,N_18404);
xor U19749 (N_19749,N_18442,N_18741);
xnor U19750 (N_19750,N_18806,N_18716);
nor U19751 (N_19751,N_19154,N_19109);
or U19752 (N_19752,N_18953,N_18507);
and U19753 (N_19753,N_19100,N_18930);
nand U19754 (N_19754,N_18749,N_18729);
nor U19755 (N_19755,N_18465,N_19111);
nor U19756 (N_19756,N_19180,N_18545);
or U19757 (N_19757,N_18681,N_19164);
nor U19758 (N_19758,N_18995,N_18980);
or U19759 (N_19759,N_18918,N_18694);
nor U19760 (N_19760,N_19090,N_19010);
xor U19761 (N_19761,N_18973,N_18746);
nand U19762 (N_19762,N_18727,N_19018);
or U19763 (N_19763,N_19031,N_18435);
xnor U19764 (N_19764,N_18459,N_18622);
nor U19765 (N_19765,N_18403,N_19056);
xnor U19766 (N_19766,N_18630,N_19103);
xor U19767 (N_19767,N_18867,N_18625);
xnor U19768 (N_19768,N_18872,N_18541);
xnor U19769 (N_19769,N_18880,N_19014);
nand U19770 (N_19770,N_18882,N_18881);
nand U19771 (N_19771,N_18792,N_18852);
nor U19772 (N_19772,N_18403,N_18683);
or U19773 (N_19773,N_18693,N_18936);
and U19774 (N_19774,N_19149,N_18410);
xor U19775 (N_19775,N_18739,N_18407);
and U19776 (N_19776,N_19069,N_19046);
nand U19777 (N_19777,N_18725,N_18527);
nor U19778 (N_19778,N_19023,N_18880);
nand U19779 (N_19779,N_19087,N_19146);
and U19780 (N_19780,N_18993,N_19028);
nor U19781 (N_19781,N_18900,N_18915);
or U19782 (N_19782,N_18667,N_19125);
xnor U19783 (N_19783,N_18734,N_18488);
nor U19784 (N_19784,N_18658,N_19091);
nand U19785 (N_19785,N_19051,N_19008);
xor U19786 (N_19786,N_18898,N_18682);
nand U19787 (N_19787,N_18855,N_18672);
nor U19788 (N_19788,N_18814,N_18994);
nand U19789 (N_19789,N_19183,N_18833);
xor U19790 (N_19790,N_19178,N_18588);
xnor U19791 (N_19791,N_18785,N_19143);
and U19792 (N_19792,N_18932,N_18781);
or U19793 (N_19793,N_18890,N_18770);
nand U19794 (N_19794,N_18456,N_18604);
xor U19795 (N_19795,N_18723,N_18788);
xor U19796 (N_19796,N_18693,N_18423);
xor U19797 (N_19797,N_18883,N_18944);
and U19798 (N_19798,N_18774,N_19128);
nor U19799 (N_19799,N_18879,N_18903);
and U19800 (N_19800,N_18446,N_18706);
nand U19801 (N_19801,N_18958,N_18980);
xnor U19802 (N_19802,N_19078,N_19092);
or U19803 (N_19803,N_18525,N_19169);
or U19804 (N_19804,N_18656,N_19155);
nand U19805 (N_19805,N_18625,N_18763);
or U19806 (N_19806,N_18788,N_19139);
xnor U19807 (N_19807,N_18836,N_18728);
and U19808 (N_19808,N_18410,N_18947);
nand U19809 (N_19809,N_19069,N_18650);
nand U19810 (N_19810,N_18660,N_18787);
xor U19811 (N_19811,N_18666,N_18411);
xor U19812 (N_19812,N_19028,N_18939);
xnor U19813 (N_19813,N_19087,N_18701);
nor U19814 (N_19814,N_18602,N_19185);
or U19815 (N_19815,N_19089,N_18944);
and U19816 (N_19816,N_18786,N_18519);
or U19817 (N_19817,N_18929,N_18882);
or U19818 (N_19818,N_18825,N_18570);
nor U19819 (N_19819,N_18403,N_18565);
and U19820 (N_19820,N_18792,N_18634);
nand U19821 (N_19821,N_18744,N_18527);
and U19822 (N_19822,N_18477,N_18453);
nand U19823 (N_19823,N_18778,N_19002);
or U19824 (N_19824,N_18971,N_18827);
nand U19825 (N_19825,N_18596,N_18776);
xor U19826 (N_19826,N_19064,N_18497);
and U19827 (N_19827,N_18941,N_18823);
xor U19828 (N_19828,N_19023,N_18748);
nand U19829 (N_19829,N_18856,N_18910);
or U19830 (N_19830,N_18687,N_19039);
or U19831 (N_19831,N_18934,N_18414);
and U19832 (N_19832,N_18733,N_19171);
or U19833 (N_19833,N_18939,N_18585);
or U19834 (N_19834,N_18783,N_18893);
or U19835 (N_19835,N_18931,N_18492);
xnor U19836 (N_19836,N_19094,N_19175);
xnor U19837 (N_19837,N_19118,N_19082);
xnor U19838 (N_19838,N_18547,N_18982);
xor U19839 (N_19839,N_18482,N_18439);
nor U19840 (N_19840,N_18450,N_19125);
nor U19841 (N_19841,N_18558,N_18840);
xnor U19842 (N_19842,N_18701,N_18589);
nor U19843 (N_19843,N_19124,N_18582);
xor U19844 (N_19844,N_18628,N_19146);
and U19845 (N_19845,N_18622,N_19122);
xor U19846 (N_19846,N_19026,N_18862);
and U19847 (N_19847,N_18481,N_18461);
or U19848 (N_19848,N_18655,N_18901);
nor U19849 (N_19849,N_19070,N_19030);
nand U19850 (N_19850,N_18628,N_18439);
xnor U19851 (N_19851,N_19189,N_19096);
nand U19852 (N_19852,N_18810,N_18674);
nand U19853 (N_19853,N_18586,N_19105);
nor U19854 (N_19854,N_19076,N_18699);
nand U19855 (N_19855,N_18520,N_19152);
nor U19856 (N_19856,N_18867,N_18637);
nor U19857 (N_19857,N_18924,N_18747);
nand U19858 (N_19858,N_19052,N_19105);
nor U19859 (N_19859,N_18652,N_18712);
or U19860 (N_19860,N_18852,N_19176);
nor U19861 (N_19861,N_18680,N_18573);
xor U19862 (N_19862,N_19160,N_18507);
or U19863 (N_19863,N_18709,N_19066);
or U19864 (N_19864,N_18485,N_18803);
nor U19865 (N_19865,N_18855,N_18813);
xor U19866 (N_19866,N_19047,N_18915);
and U19867 (N_19867,N_18870,N_18996);
and U19868 (N_19868,N_18523,N_19042);
nand U19869 (N_19869,N_19087,N_19011);
nor U19870 (N_19870,N_18588,N_18932);
nor U19871 (N_19871,N_18894,N_18572);
xor U19872 (N_19872,N_19060,N_18615);
and U19873 (N_19873,N_18778,N_19135);
xor U19874 (N_19874,N_18822,N_18492);
and U19875 (N_19875,N_19078,N_18708);
nand U19876 (N_19876,N_18867,N_19083);
nand U19877 (N_19877,N_18924,N_18579);
nand U19878 (N_19878,N_18456,N_18916);
and U19879 (N_19879,N_18633,N_18968);
nor U19880 (N_19880,N_18755,N_18623);
xor U19881 (N_19881,N_18985,N_18838);
xnor U19882 (N_19882,N_19014,N_18534);
nor U19883 (N_19883,N_18424,N_19195);
or U19884 (N_19884,N_19144,N_18681);
or U19885 (N_19885,N_19119,N_18473);
xnor U19886 (N_19886,N_18445,N_18578);
xor U19887 (N_19887,N_18873,N_18779);
or U19888 (N_19888,N_19180,N_19130);
nor U19889 (N_19889,N_18637,N_18992);
xnor U19890 (N_19890,N_18785,N_18790);
xor U19891 (N_19891,N_18494,N_18489);
nand U19892 (N_19892,N_18485,N_18534);
xnor U19893 (N_19893,N_18507,N_18711);
and U19894 (N_19894,N_18610,N_18892);
nand U19895 (N_19895,N_19046,N_18474);
xnor U19896 (N_19896,N_19151,N_19111);
xor U19897 (N_19897,N_19146,N_18524);
nor U19898 (N_19898,N_18746,N_19169);
and U19899 (N_19899,N_18872,N_18408);
nor U19900 (N_19900,N_18825,N_19138);
nor U19901 (N_19901,N_18627,N_19099);
nor U19902 (N_19902,N_19171,N_18639);
nand U19903 (N_19903,N_18778,N_18516);
nand U19904 (N_19904,N_19076,N_19034);
nand U19905 (N_19905,N_18794,N_18896);
nor U19906 (N_19906,N_19170,N_18654);
or U19907 (N_19907,N_18952,N_18665);
xor U19908 (N_19908,N_18604,N_18805);
or U19909 (N_19909,N_19102,N_18537);
nor U19910 (N_19910,N_18835,N_18690);
nand U19911 (N_19911,N_19098,N_19008);
xor U19912 (N_19912,N_19018,N_19005);
or U19913 (N_19913,N_18917,N_18524);
xnor U19914 (N_19914,N_18705,N_18460);
xor U19915 (N_19915,N_18763,N_18540);
and U19916 (N_19916,N_18875,N_19024);
nor U19917 (N_19917,N_18903,N_18680);
nor U19918 (N_19918,N_18863,N_18948);
or U19919 (N_19919,N_18645,N_18773);
nor U19920 (N_19920,N_18951,N_19131);
or U19921 (N_19921,N_18405,N_19150);
nor U19922 (N_19922,N_18527,N_18605);
or U19923 (N_19923,N_18556,N_18436);
nor U19924 (N_19924,N_18858,N_18404);
and U19925 (N_19925,N_18552,N_18496);
and U19926 (N_19926,N_18576,N_19012);
nand U19927 (N_19927,N_18403,N_19032);
nand U19928 (N_19928,N_19061,N_18949);
xnor U19929 (N_19929,N_18916,N_19174);
or U19930 (N_19930,N_18693,N_18741);
or U19931 (N_19931,N_18495,N_18478);
nand U19932 (N_19932,N_19003,N_18550);
nand U19933 (N_19933,N_18954,N_18668);
or U19934 (N_19934,N_18760,N_18580);
nand U19935 (N_19935,N_19155,N_18629);
nand U19936 (N_19936,N_18484,N_18985);
or U19937 (N_19937,N_19164,N_18918);
xor U19938 (N_19938,N_18556,N_19198);
nand U19939 (N_19939,N_19101,N_19146);
and U19940 (N_19940,N_18422,N_18409);
and U19941 (N_19941,N_19082,N_18541);
nand U19942 (N_19942,N_18527,N_18996);
xor U19943 (N_19943,N_18462,N_18685);
xor U19944 (N_19944,N_19119,N_19105);
nand U19945 (N_19945,N_19191,N_18695);
nor U19946 (N_19946,N_19122,N_18730);
xnor U19947 (N_19947,N_18645,N_19197);
or U19948 (N_19948,N_18598,N_18842);
nand U19949 (N_19949,N_18484,N_18788);
nor U19950 (N_19950,N_18508,N_19109);
nor U19951 (N_19951,N_18432,N_19037);
nor U19952 (N_19952,N_18713,N_18409);
and U19953 (N_19953,N_18496,N_18582);
xor U19954 (N_19954,N_18947,N_18529);
and U19955 (N_19955,N_18553,N_19180);
nor U19956 (N_19956,N_19078,N_18841);
or U19957 (N_19957,N_18686,N_18859);
xor U19958 (N_19958,N_19153,N_18729);
or U19959 (N_19959,N_19103,N_18784);
nand U19960 (N_19960,N_19046,N_18922);
nor U19961 (N_19961,N_18980,N_18687);
nand U19962 (N_19962,N_18483,N_18907);
and U19963 (N_19963,N_18475,N_18433);
and U19964 (N_19964,N_18410,N_18749);
and U19965 (N_19965,N_18712,N_18476);
xor U19966 (N_19966,N_19126,N_18876);
nand U19967 (N_19967,N_19023,N_18555);
or U19968 (N_19968,N_19176,N_18962);
or U19969 (N_19969,N_18588,N_18920);
or U19970 (N_19970,N_18564,N_18519);
and U19971 (N_19971,N_18861,N_19074);
nor U19972 (N_19972,N_19198,N_19119);
nand U19973 (N_19973,N_19192,N_19182);
xnor U19974 (N_19974,N_18821,N_18883);
and U19975 (N_19975,N_18881,N_19050);
nand U19976 (N_19976,N_18508,N_18401);
xnor U19977 (N_19977,N_18903,N_19182);
nand U19978 (N_19978,N_18802,N_18751);
nand U19979 (N_19979,N_18964,N_18440);
nand U19980 (N_19980,N_18999,N_18696);
xor U19981 (N_19981,N_18895,N_18535);
nand U19982 (N_19982,N_18478,N_18461);
nor U19983 (N_19983,N_19084,N_18435);
xnor U19984 (N_19984,N_19093,N_19146);
xnor U19985 (N_19985,N_18823,N_18974);
xnor U19986 (N_19986,N_18935,N_18538);
or U19987 (N_19987,N_18969,N_18496);
or U19988 (N_19988,N_19046,N_18909);
or U19989 (N_19989,N_18916,N_18546);
nor U19990 (N_19990,N_18510,N_18461);
nor U19991 (N_19991,N_19121,N_19140);
and U19992 (N_19992,N_18428,N_19056);
and U19993 (N_19993,N_18658,N_19086);
xor U19994 (N_19994,N_18736,N_18971);
xnor U19995 (N_19995,N_18422,N_18440);
xor U19996 (N_19996,N_18712,N_19109);
and U19997 (N_19997,N_18596,N_18528);
nand U19998 (N_19998,N_18896,N_18892);
and U19999 (N_19999,N_19070,N_18918);
and UO_0 (O_0,N_19753,N_19716);
nand UO_1 (O_1,N_19611,N_19597);
xnor UO_2 (O_2,N_19995,N_19299);
or UO_3 (O_3,N_19605,N_19225);
and UO_4 (O_4,N_19800,N_19454);
nand UO_5 (O_5,N_19896,N_19320);
and UO_6 (O_6,N_19712,N_19651);
or UO_7 (O_7,N_19243,N_19448);
and UO_8 (O_8,N_19237,N_19851);
nor UO_9 (O_9,N_19739,N_19915);
nor UO_10 (O_10,N_19848,N_19941);
or UO_11 (O_11,N_19447,N_19643);
or UO_12 (O_12,N_19734,N_19285);
xnor UO_13 (O_13,N_19562,N_19996);
or UO_14 (O_14,N_19287,N_19613);
nand UO_15 (O_15,N_19376,N_19971);
nor UO_16 (O_16,N_19512,N_19771);
xor UO_17 (O_17,N_19621,N_19819);
xor UO_18 (O_18,N_19560,N_19961);
xor UO_19 (O_19,N_19600,N_19741);
xor UO_20 (O_20,N_19917,N_19650);
xnor UO_21 (O_21,N_19964,N_19524);
or UO_22 (O_22,N_19815,N_19442);
nor UO_23 (O_23,N_19318,N_19238);
xnor UO_24 (O_24,N_19698,N_19968);
nand UO_25 (O_25,N_19797,N_19680);
xor UO_26 (O_26,N_19918,N_19508);
or UO_27 (O_27,N_19947,N_19452);
xor UO_28 (O_28,N_19569,N_19882);
nand UO_29 (O_29,N_19930,N_19521);
or UO_30 (O_30,N_19603,N_19891);
nand UO_31 (O_31,N_19570,N_19488);
or UO_32 (O_32,N_19236,N_19864);
or UO_33 (O_33,N_19558,N_19344);
nand UO_34 (O_34,N_19982,N_19647);
or UO_35 (O_35,N_19247,N_19343);
or UO_36 (O_36,N_19821,N_19765);
xnor UO_37 (O_37,N_19210,N_19718);
and UO_38 (O_38,N_19818,N_19701);
xor UO_39 (O_39,N_19853,N_19214);
xor UO_40 (O_40,N_19474,N_19399);
nand UO_41 (O_41,N_19565,N_19455);
and UO_42 (O_42,N_19519,N_19931);
xnor UO_43 (O_43,N_19586,N_19633);
nand UO_44 (O_44,N_19743,N_19900);
nor UO_45 (O_45,N_19746,N_19531);
nand UO_46 (O_46,N_19298,N_19217);
or UO_47 (O_47,N_19580,N_19678);
and UO_48 (O_48,N_19733,N_19735);
nor UO_49 (O_49,N_19629,N_19654);
or UO_50 (O_50,N_19413,N_19520);
or UO_51 (O_51,N_19387,N_19370);
xnor UO_52 (O_52,N_19581,N_19708);
or UO_53 (O_53,N_19946,N_19942);
and UO_54 (O_54,N_19828,N_19908);
and UO_55 (O_55,N_19468,N_19278);
nand UO_56 (O_56,N_19525,N_19726);
or UO_57 (O_57,N_19705,N_19725);
and UO_58 (O_58,N_19464,N_19628);
and UO_59 (O_59,N_19216,N_19782);
and UO_60 (O_60,N_19596,N_19489);
and UO_61 (O_61,N_19513,N_19740);
and UO_62 (O_62,N_19724,N_19775);
xor UO_63 (O_63,N_19672,N_19847);
and UO_64 (O_64,N_19595,N_19466);
and UO_65 (O_65,N_19538,N_19754);
or UO_66 (O_66,N_19966,N_19663);
or UO_67 (O_67,N_19699,N_19736);
nor UO_68 (O_68,N_19505,N_19655);
xnor UO_69 (O_69,N_19912,N_19806);
and UO_70 (O_70,N_19393,N_19617);
and UO_71 (O_71,N_19213,N_19606);
nand UO_72 (O_72,N_19645,N_19902);
nor UO_73 (O_73,N_19533,N_19446);
or UO_74 (O_74,N_19939,N_19228);
xnor UO_75 (O_75,N_19286,N_19710);
nor UO_76 (O_76,N_19461,N_19737);
xnor UO_77 (O_77,N_19357,N_19421);
nor UO_78 (O_78,N_19316,N_19279);
xor UO_79 (O_79,N_19527,N_19886);
xor UO_80 (O_80,N_19817,N_19414);
xor UO_81 (O_81,N_19683,N_19978);
and UO_82 (O_82,N_19445,N_19437);
and UO_83 (O_83,N_19612,N_19959);
and UO_84 (O_84,N_19630,N_19709);
nand UO_85 (O_85,N_19204,N_19561);
and UO_86 (O_86,N_19635,N_19786);
xnor UO_87 (O_87,N_19410,N_19522);
and UO_88 (O_88,N_19850,N_19954);
nor UO_89 (O_89,N_19273,N_19400);
nor UO_90 (O_90,N_19338,N_19997);
and UO_91 (O_91,N_19591,N_19296);
or UO_92 (O_92,N_19317,N_19755);
nand UO_93 (O_93,N_19773,N_19396);
or UO_94 (O_94,N_19764,N_19648);
nand UO_95 (O_95,N_19785,N_19499);
nor UO_96 (O_96,N_19636,N_19507);
and UO_97 (O_97,N_19252,N_19251);
nand UO_98 (O_98,N_19307,N_19384);
and UO_99 (O_99,N_19266,N_19567);
nor UO_100 (O_100,N_19681,N_19262);
or UO_101 (O_101,N_19496,N_19686);
xnor UO_102 (O_102,N_19665,N_19551);
xor UO_103 (O_103,N_19220,N_19890);
nor UO_104 (O_104,N_19669,N_19319);
nor UO_105 (O_105,N_19267,N_19543);
xnor UO_106 (O_106,N_19984,N_19974);
and UO_107 (O_107,N_19892,N_19436);
xnor UO_108 (O_108,N_19334,N_19844);
or UO_109 (O_109,N_19255,N_19721);
or UO_110 (O_110,N_19294,N_19879);
and UO_111 (O_111,N_19509,N_19469);
and UO_112 (O_112,N_19388,N_19517);
xnor UO_113 (O_113,N_19993,N_19308);
and UO_114 (O_114,N_19728,N_19549);
nor UO_115 (O_115,N_19532,N_19257);
xnor UO_116 (O_116,N_19530,N_19377);
and UO_117 (O_117,N_19662,N_19328);
and UO_118 (O_118,N_19988,N_19829);
nor UO_119 (O_119,N_19932,N_19749);
nor UO_120 (O_120,N_19714,N_19289);
xnor UO_121 (O_121,N_19925,N_19534);
and UO_122 (O_122,N_19443,N_19293);
xnor UO_123 (O_123,N_19608,N_19967);
xor UO_124 (O_124,N_19390,N_19300);
and UO_125 (O_125,N_19420,N_19881);
xnor UO_126 (O_126,N_19638,N_19953);
nand UO_127 (O_127,N_19514,N_19242);
xor UO_128 (O_128,N_19827,N_19837);
xnor UO_129 (O_129,N_19878,N_19835);
nand UO_130 (O_130,N_19667,N_19618);
and UO_131 (O_131,N_19313,N_19899);
and UO_132 (O_132,N_19431,N_19205);
nor UO_133 (O_133,N_19550,N_19620);
and UO_134 (O_134,N_19412,N_19975);
and UO_135 (O_135,N_19843,N_19268);
and UO_136 (O_136,N_19830,N_19417);
and UO_137 (O_137,N_19582,N_19676);
or UO_138 (O_138,N_19234,N_19955);
or UO_139 (O_139,N_19994,N_19703);
or UO_140 (O_140,N_19752,N_19704);
or UO_141 (O_141,N_19398,N_19889);
nor UO_142 (O_142,N_19552,N_19579);
nand UO_143 (O_143,N_19342,N_19641);
or UO_144 (O_144,N_19212,N_19311);
and UO_145 (O_145,N_19240,N_19402);
and UO_146 (O_146,N_19986,N_19875);
nor UO_147 (O_147,N_19463,N_19989);
and UO_148 (O_148,N_19295,N_19555);
xnor UO_149 (O_149,N_19280,N_19483);
and UO_150 (O_150,N_19480,N_19506);
xor UO_151 (O_151,N_19992,N_19671);
xor UO_152 (O_152,N_19987,N_19774);
or UO_153 (O_153,N_19456,N_19924);
or UO_154 (O_154,N_19554,N_19478);
and UO_155 (O_155,N_19487,N_19745);
nor UO_156 (O_156,N_19409,N_19656);
and UO_157 (O_157,N_19965,N_19248);
nand UO_158 (O_158,N_19222,N_19501);
and UO_159 (O_159,N_19223,N_19970);
xor UO_160 (O_160,N_19485,N_19825);
nand UO_161 (O_161,N_19465,N_19516);
nand UO_162 (O_162,N_19305,N_19564);
nor UO_163 (O_163,N_19804,N_19903);
or UO_164 (O_164,N_19623,N_19901);
nor UO_165 (O_165,N_19467,N_19625);
xor UO_166 (O_166,N_19999,N_19691);
nor UO_167 (O_167,N_19253,N_19768);
or UO_168 (O_168,N_19783,N_19833);
nand UO_169 (O_169,N_19679,N_19880);
nor UO_170 (O_170,N_19366,N_19211);
nand UO_171 (O_171,N_19244,N_19491);
nand UO_172 (O_172,N_19365,N_19547);
xnor UO_173 (O_173,N_19484,N_19916);
nand UO_174 (O_174,N_19622,N_19354);
nor UO_175 (O_175,N_19327,N_19218);
and UO_176 (O_176,N_19742,N_19292);
nand UO_177 (O_177,N_19808,N_19738);
xor UO_178 (O_178,N_19258,N_19335);
nor UO_179 (O_179,N_19619,N_19598);
nor UO_180 (O_180,N_19784,N_19867);
xor UO_181 (O_181,N_19938,N_19962);
and UO_182 (O_182,N_19557,N_19624);
and UO_183 (O_183,N_19424,N_19644);
or UO_184 (O_184,N_19688,N_19323);
xor UO_185 (O_185,N_19347,N_19405);
or UO_186 (O_186,N_19788,N_19849);
nand UO_187 (O_187,N_19649,N_19868);
nand UO_188 (O_188,N_19777,N_19927);
nand UO_189 (O_189,N_19846,N_19602);
and UO_190 (O_190,N_19948,N_19919);
nor UO_191 (O_191,N_19814,N_19432);
or UO_192 (O_192,N_19794,N_19492);
xnor UO_193 (O_193,N_19952,N_19796);
xor UO_194 (O_194,N_19497,N_19594);
nand UO_195 (O_195,N_19778,N_19838);
nor UO_196 (O_196,N_19288,N_19711);
nor UO_197 (O_197,N_19274,N_19227);
xor UO_198 (O_198,N_19870,N_19438);
or UO_199 (O_199,N_19760,N_19713);
or UO_200 (O_200,N_19593,N_19763);
xnor UO_201 (O_201,N_19350,N_19254);
nor UO_202 (O_202,N_19553,N_19271);
xor UO_203 (O_203,N_19700,N_19960);
or UO_204 (O_204,N_19291,N_19559);
nand UO_205 (O_205,N_19877,N_19858);
nor UO_206 (O_206,N_19816,N_19799);
xor UO_207 (O_207,N_19418,N_19346);
xnor UO_208 (O_208,N_19857,N_19707);
nand UO_209 (O_209,N_19872,N_19610);
or UO_210 (O_210,N_19859,N_19427);
xnor UO_211 (O_211,N_19284,N_19208);
or UO_212 (O_212,N_19840,N_19360);
nor UO_213 (O_213,N_19841,N_19976);
or UO_214 (O_214,N_19926,N_19661);
and UO_215 (O_215,N_19476,N_19637);
and UO_216 (O_216,N_19601,N_19460);
and UO_217 (O_217,N_19574,N_19382);
and UO_218 (O_218,N_19911,N_19362);
and UO_219 (O_219,N_19950,N_19498);
xnor UO_220 (O_220,N_19407,N_19684);
xnor UO_221 (O_221,N_19440,N_19403);
xor UO_222 (O_222,N_19371,N_19219);
xnor UO_223 (O_223,N_19957,N_19201);
and UO_224 (O_224,N_19395,N_19856);
xnor UO_225 (O_225,N_19949,N_19839);
nand UO_226 (O_226,N_19936,N_19325);
xor UO_227 (O_227,N_19653,N_19331);
or UO_228 (O_228,N_19451,N_19435);
nand UO_229 (O_229,N_19404,N_19290);
and UO_230 (O_230,N_19895,N_19303);
and UO_231 (O_231,N_19425,N_19275);
nor UO_232 (O_232,N_19368,N_19215);
or UO_233 (O_233,N_19545,N_19666);
nand UO_234 (O_234,N_19920,N_19772);
or UO_235 (O_235,N_19529,N_19528);
nand UO_236 (O_236,N_19263,N_19757);
or UO_237 (O_237,N_19202,N_19542);
nor UO_238 (O_238,N_19722,N_19715);
or UO_239 (O_239,N_19477,N_19694);
or UO_240 (O_240,N_19332,N_19646);
or UO_241 (O_241,N_19571,N_19471);
and UO_242 (O_242,N_19401,N_19479);
xnor UO_243 (O_243,N_19614,N_19458);
xnor UO_244 (O_244,N_19495,N_19675);
xor UO_245 (O_245,N_19885,N_19209);
or UO_246 (O_246,N_19909,N_19588);
and UO_247 (O_247,N_19801,N_19758);
nand UO_248 (O_248,N_19563,N_19459);
or UO_249 (O_249,N_19910,N_19259);
and UO_250 (O_250,N_19397,N_19315);
nand UO_251 (O_251,N_19751,N_19807);
and UO_252 (O_252,N_19876,N_19692);
or UO_253 (O_253,N_19793,N_19536);
and UO_254 (O_254,N_19322,N_19353);
or UO_255 (O_255,N_19535,N_19221);
and UO_256 (O_256,N_19824,N_19626);
xnor UO_257 (O_257,N_19803,N_19862);
nand UO_258 (O_258,N_19956,N_19940);
nand UO_259 (O_259,N_19345,N_19207);
nand UO_260 (O_260,N_19659,N_19732);
xor UO_261 (O_261,N_19352,N_19233);
nand UO_262 (O_262,N_19566,N_19750);
xor UO_263 (O_263,N_19983,N_19583);
xor UO_264 (O_264,N_19235,N_19822);
xnor UO_265 (O_265,N_19587,N_19756);
nand UO_266 (O_266,N_19276,N_19355);
nor UO_267 (O_267,N_19852,N_19943);
nand UO_268 (O_268,N_19363,N_19312);
xnor UO_269 (O_269,N_19706,N_19584);
or UO_270 (O_270,N_19423,N_19250);
and UO_271 (O_271,N_19798,N_19906);
nand UO_272 (O_272,N_19609,N_19556);
nor UO_273 (O_273,N_19744,N_19979);
xnor UO_274 (O_274,N_19873,N_19812);
or UO_275 (O_275,N_19282,N_19668);
and UO_276 (O_276,N_19537,N_19504);
xor UO_277 (O_277,N_19523,N_19894);
or UO_278 (O_278,N_19568,N_19702);
nor UO_279 (O_279,N_19866,N_19883);
xor UO_280 (O_280,N_19854,N_19232);
nor UO_281 (O_281,N_19226,N_19391);
and UO_282 (O_282,N_19272,N_19921);
nor UO_283 (O_283,N_19241,N_19802);
or UO_284 (O_284,N_19336,N_19893);
and UO_285 (O_285,N_19406,N_19823);
xnor UO_286 (O_286,N_19657,N_19309);
or UO_287 (O_287,N_19781,N_19748);
and UO_288 (O_288,N_19958,N_19324);
and UO_289 (O_289,N_19206,N_19518);
xnor UO_290 (O_290,N_19935,N_19860);
or UO_291 (O_291,N_19321,N_19639);
or UO_292 (O_292,N_19695,N_19673);
xor UO_293 (O_293,N_19493,N_19791);
or UO_294 (O_294,N_19887,N_19314);
and UO_295 (O_295,N_19720,N_19907);
xnor UO_296 (O_296,N_19502,N_19361);
and UO_297 (O_297,N_19203,N_19717);
and UO_298 (O_298,N_19747,N_19472);
nor UO_299 (O_299,N_19865,N_19426);
or UO_300 (O_300,N_19428,N_19385);
nand UO_301 (O_301,N_19392,N_19977);
nand UO_302 (O_302,N_19905,N_19677);
and UO_303 (O_303,N_19441,N_19546);
or UO_304 (O_304,N_19730,N_19540);
or UO_305 (O_305,N_19230,N_19631);
xnor UO_306 (O_306,N_19769,N_19572);
and UO_307 (O_307,N_19245,N_19340);
xnor UO_308 (O_308,N_19373,N_19378);
and UO_309 (O_309,N_19845,N_19689);
nor UO_310 (O_310,N_19640,N_19836);
and UO_311 (O_311,N_19375,N_19897);
xnor UO_312 (O_312,N_19934,N_19929);
nor UO_313 (O_313,N_19231,N_19482);
and UO_314 (O_314,N_19356,N_19349);
and UO_315 (O_315,N_19246,N_19302);
or UO_316 (O_316,N_19577,N_19810);
nand UO_317 (O_317,N_19515,N_19607);
xor UO_318 (O_318,N_19511,N_19411);
xor UO_319 (O_319,N_19687,N_19674);
or UO_320 (O_320,N_19604,N_19348);
xnor UO_321 (O_321,N_19922,N_19270);
xor UO_322 (O_322,N_19634,N_19381);
and UO_323 (O_323,N_19727,N_19685);
or UO_324 (O_324,N_19383,N_19660);
nand UO_325 (O_325,N_19281,N_19439);
xor UO_326 (O_326,N_19767,N_19380);
nor UO_327 (O_327,N_19337,N_19229);
and UO_328 (O_328,N_19486,N_19690);
xnor UO_329 (O_329,N_19369,N_19449);
xnor UO_330 (O_330,N_19731,N_19855);
or UO_331 (O_331,N_19985,N_19642);
and UO_332 (O_332,N_19913,N_19951);
and UO_333 (O_333,N_19239,N_19386);
and UO_334 (O_334,N_19329,N_19923);
nand UO_335 (O_335,N_19842,N_19379);
nand UO_336 (O_336,N_19945,N_19578);
nand UO_337 (O_337,N_19374,N_19776);
nand UO_338 (O_338,N_19434,N_19470);
xnor UO_339 (O_339,N_19914,N_19548);
and UO_340 (O_340,N_19269,N_19358);
and UO_341 (O_341,N_19541,N_19408);
xnor UO_342 (O_342,N_19792,N_19359);
xor UO_343 (O_343,N_19973,N_19991);
xnor UO_344 (O_344,N_19928,N_19863);
or UO_345 (O_345,N_19503,N_19869);
nand UO_346 (O_346,N_19933,N_19297);
and UO_347 (O_347,N_19200,N_19494);
or UO_348 (O_348,N_19500,N_19585);
nor UO_349 (O_349,N_19790,N_19795);
nor UO_350 (O_350,N_19589,N_19990);
and UO_351 (O_351,N_19590,N_19310);
and UO_352 (O_352,N_19576,N_19980);
nand UO_353 (O_353,N_19341,N_19770);
nand UO_354 (O_354,N_19433,N_19389);
and UO_355 (O_355,N_19416,N_19615);
xnor UO_356 (O_356,N_19696,N_19969);
nor UO_357 (O_357,N_19333,N_19723);
nor UO_358 (O_358,N_19539,N_19450);
nor UO_359 (O_359,N_19481,N_19719);
nand UO_360 (O_360,N_19670,N_19544);
nand UO_361 (O_361,N_19789,N_19820);
nand UO_362 (O_362,N_19430,N_19861);
and UO_363 (O_363,N_19762,N_19224);
xor UO_364 (O_364,N_19616,N_19832);
and UO_365 (O_365,N_19277,N_19510);
or UO_366 (O_366,N_19658,N_19573);
nor UO_367 (O_367,N_19805,N_19265);
xnor UO_368 (O_368,N_19998,N_19599);
xnor UO_369 (O_369,N_19473,N_19415);
and UO_370 (O_370,N_19834,N_19972);
or UO_371 (O_371,N_19575,N_19627);
or UO_372 (O_372,N_19787,N_19394);
and UO_373 (O_373,N_19888,N_19632);
or UO_374 (O_374,N_19697,N_19831);
nor UO_375 (O_375,N_19283,N_19761);
nor UO_376 (O_376,N_19826,N_19429);
nand UO_377 (O_377,N_19729,N_19264);
xor UO_378 (O_378,N_19811,N_19944);
or UO_379 (O_379,N_19871,N_19367);
nor UO_380 (O_380,N_19526,N_19664);
nand UO_381 (O_381,N_19937,N_19981);
xnor UO_382 (O_382,N_19304,N_19904);
or UO_383 (O_383,N_19372,N_19963);
nand UO_384 (O_384,N_19592,N_19780);
and UO_385 (O_385,N_19682,N_19766);
and UO_386 (O_386,N_19874,N_19306);
and UO_387 (O_387,N_19249,N_19260);
or UO_388 (O_388,N_19339,N_19475);
or UO_389 (O_389,N_19444,N_19261);
or UO_390 (O_390,N_19351,N_19453);
xor UO_391 (O_391,N_19364,N_19462);
and UO_392 (O_392,N_19759,N_19457);
nand UO_393 (O_393,N_19301,N_19652);
xor UO_394 (O_394,N_19809,N_19884);
and UO_395 (O_395,N_19898,N_19490);
or UO_396 (O_396,N_19330,N_19813);
xor UO_397 (O_397,N_19326,N_19779);
xnor UO_398 (O_398,N_19693,N_19422);
or UO_399 (O_399,N_19419,N_19256);
or UO_400 (O_400,N_19330,N_19682);
or UO_401 (O_401,N_19659,N_19926);
nand UO_402 (O_402,N_19472,N_19574);
xor UO_403 (O_403,N_19895,N_19334);
or UO_404 (O_404,N_19391,N_19289);
and UO_405 (O_405,N_19296,N_19806);
nand UO_406 (O_406,N_19740,N_19921);
nand UO_407 (O_407,N_19631,N_19345);
and UO_408 (O_408,N_19331,N_19378);
nand UO_409 (O_409,N_19204,N_19536);
or UO_410 (O_410,N_19467,N_19501);
xor UO_411 (O_411,N_19653,N_19679);
or UO_412 (O_412,N_19966,N_19823);
xor UO_413 (O_413,N_19231,N_19852);
or UO_414 (O_414,N_19382,N_19315);
nand UO_415 (O_415,N_19939,N_19595);
and UO_416 (O_416,N_19796,N_19841);
xnor UO_417 (O_417,N_19871,N_19489);
nand UO_418 (O_418,N_19645,N_19609);
nand UO_419 (O_419,N_19307,N_19646);
xor UO_420 (O_420,N_19571,N_19261);
xor UO_421 (O_421,N_19269,N_19255);
xor UO_422 (O_422,N_19564,N_19467);
or UO_423 (O_423,N_19375,N_19958);
nor UO_424 (O_424,N_19209,N_19386);
nand UO_425 (O_425,N_19344,N_19549);
nand UO_426 (O_426,N_19671,N_19814);
nand UO_427 (O_427,N_19611,N_19513);
or UO_428 (O_428,N_19620,N_19825);
and UO_429 (O_429,N_19405,N_19355);
nand UO_430 (O_430,N_19634,N_19734);
nand UO_431 (O_431,N_19847,N_19717);
xor UO_432 (O_432,N_19544,N_19401);
or UO_433 (O_433,N_19721,N_19923);
or UO_434 (O_434,N_19540,N_19575);
and UO_435 (O_435,N_19879,N_19428);
xor UO_436 (O_436,N_19964,N_19316);
nand UO_437 (O_437,N_19205,N_19784);
and UO_438 (O_438,N_19922,N_19275);
nand UO_439 (O_439,N_19267,N_19406);
and UO_440 (O_440,N_19895,N_19472);
xor UO_441 (O_441,N_19808,N_19522);
xnor UO_442 (O_442,N_19336,N_19537);
nand UO_443 (O_443,N_19724,N_19707);
or UO_444 (O_444,N_19214,N_19276);
nor UO_445 (O_445,N_19253,N_19762);
nor UO_446 (O_446,N_19286,N_19484);
nand UO_447 (O_447,N_19459,N_19493);
and UO_448 (O_448,N_19486,N_19532);
nand UO_449 (O_449,N_19360,N_19533);
or UO_450 (O_450,N_19733,N_19655);
nand UO_451 (O_451,N_19517,N_19311);
nand UO_452 (O_452,N_19802,N_19243);
or UO_453 (O_453,N_19435,N_19975);
and UO_454 (O_454,N_19284,N_19447);
or UO_455 (O_455,N_19816,N_19865);
or UO_456 (O_456,N_19894,N_19469);
xnor UO_457 (O_457,N_19406,N_19328);
xor UO_458 (O_458,N_19679,N_19700);
and UO_459 (O_459,N_19346,N_19537);
nand UO_460 (O_460,N_19541,N_19524);
nor UO_461 (O_461,N_19460,N_19589);
nand UO_462 (O_462,N_19288,N_19528);
nand UO_463 (O_463,N_19719,N_19883);
and UO_464 (O_464,N_19757,N_19381);
xnor UO_465 (O_465,N_19388,N_19890);
or UO_466 (O_466,N_19471,N_19854);
or UO_467 (O_467,N_19739,N_19533);
and UO_468 (O_468,N_19221,N_19457);
or UO_469 (O_469,N_19228,N_19785);
or UO_470 (O_470,N_19969,N_19397);
xor UO_471 (O_471,N_19941,N_19785);
nor UO_472 (O_472,N_19324,N_19392);
nor UO_473 (O_473,N_19271,N_19344);
nand UO_474 (O_474,N_19325,N_19436);
nand UO_475 (O_475,N_19450,N_19927);
and UO_476 (O_476,N_19502,N_19623);
and UO_477 (O_477,N_19755,N_19607);
or UO_478 (O_478,N_19676,N_19358);
or UO_479 (O_479,N_19979,N_19738);
nand UO_480 (O_480,N_19359,N_19206);
or UO_481 (O_481,N_19799,N_19741);
and UO_482 (O_482,N_19204,N_19433);
xnor UO_483 (O_483,N_19226,N_19984);
or UO_484 (O_484,N_19555,N_19831);
nor UO_485 (O_485,N_19597,N_19272);
and UO_486 (O_486,N_19538,N_19321);
nand UO_487 (O_487,N_19503,N_19510);
or UO_488 (O_488,N_19207,N_19969);
nand UO_489 (O_489,N_19538,N_19618);
and UO_490 (O_490,N_19809,N_19692);
or UO_491 (O_491,N_19289,N_19992);
nand UO_492 (O_492,N_19267,N_19562);
xor UO_493 (O_493,N_19828,N_19296);
xor UO_494 (O_494,N_19809,N_19584);
nor UO_495 (O_495,N_19535,N_19324);
xor UO_496 (O_496,N_19894,N_19778);
nand UO_497 (O_497,N_19588,N_19547);
xor UO_498 (O_498,N_19930,N_19544);
nand UO_499 (O_499,N_19891,N_19226);
nor UO_500 (O_500,N_19605,N_19254);
nand UO_501 (O_501,N_19818,N_19610);
nand UO_502 (O_502,N_19790,N_19263);
or UO_503 (O_503,N_19862,N_19929);
nor UO_504 (O_504,N_19445,N_19217);
nor UO_505 (O_505,N_19554,N_19298);
and UO_506 (O_506,N_19331,N_19389);
and UO_507 (O_507,N_19386,N_19516);
and UO_508 (O_508,N_19685,N_19608);
nand UO_509 (O_509,N_19739,N_19308);
and UO_510 (O_510,N_19486,N_19833);
xor UO_511 (O_511,N_19993,N_19851);
nand UO_512 (O_512,N_19858,N_19487);
nand UO_513 (O_513,N_19350,N_19909);
and UO_514 (O_514,N_19967,N_19613);
and UO_515 (O_515,N_19466,N_19266);
and UO_516 (O_516,N_19671,N_19659);
and UO_517 (O_517,N_19781,N_19347);
nor UO_518 (O_518,N_19792,N_19436);
or UO_519 (O_519,N_19912,N_19693);
nand UO_520 (O_520,N_19250,N_19860);
nand UO_521 (O_521,N_19232,N_19832);
and UO_522 (O_522,N_19484,N_19344);
nor UO_523 (O_523,N_19518,N_19419);
nor UO_524 (O_524,N_19262,N_19808);
nand UO_525 (O_525,N_19694,N_19776);
and UO_526 (O_526,N_19570,N_19485);
and UO_527 (O_527,N_19593,N_19531);
and UO_528 (O_528,N_19261,N_19511);
nand UO_529 (O_529,N_19297,N_19694);
nand UO_530 (O_530,N_19713,N_19949);
nand UO_531 (O_531,N_19334,N_19689);
nand UO_532 (O_532,N_19670,N_19491);
or UO_533 (O_533,N_19614,N_19771);
or UO_534 (O_534,N_19842,N_19695);
xnor UO_535 (O_535,N_19644,N_19917);
or UO_536 (O_536,N_19586,N_19784);
nand UO_537 (O_537,N_19576,N_19676);
nor UO_538 (O_538,N_19686,N_19321);
nand UO_539 (O_539,N_19702,N_19435);
or UO_540 (O_540,N_19784,N_19820);
nand UO_541 (O_541,N_19948,N_19698);
nand UO_542 (O_542,N_19883,N_19860);
or UO_543 (O_543,N_19582,N_19706);
xnor UO_544 (O_544,N_19677,N_19290);
nand UO_545 (O_545,N_19268,N_19255);
or UO_546 (O_546,N_19437,N_19356);
nor UO_547 (O_547,N_19917,N_19580);
xor UO_548 (O_548,N_19256,N_19737);
nand UO_549 (O_549,N_19353,N_19612);
or UO_550 (O_550,N_19312,N_19667);
nand UO_551 (O_551,N_19273,N_19239);
nand UO_552 (O_552,N_19607,N_19324);
nor UO_553 (O_553,N_19844,N_19662);
and UO_554 (O_554,N_19446,N_19629);
or UO_555 (O_555,N_19206,N_19329);
or UO_556 (O_556,N_19278,N_19317);
nor UO_557 (O_557,N_19725,N_19992);
nand UO_558 (O_558,N_19847,N_19589);
and UO_559 (O_559,N_19327,N_19489);
nor UO_560 (O_560,N_19533,N_19606);
or UO_561 (O_561,N_19704,N_19623);
nand UO_562 (O_562,N_19976,N_19474);
and UO_563 (O_563,N_19760,N_19892);
xor UO_564 (O_564,N_19291,N_19539);
and UO_565 (O_565,N_19876,N_19381);
nor UO_566 (O_566,N_19655,N_19516);
xor UO_567 (O_567,N_19211,N_19998);
nor UO_568 (O_568,N_19471,N_19849);
and UO_569 (O_569,N_19836,N_19818);
or UO_570 (O_570,N_19204,N_19318);
nor UO_571 (O_571,N_19222,N_19252);
and UO_572 (O_572,N_19761,N_19937);
and UO_573 (O_573,N_19479,N_19342);
and UO_574 (O_574,N_19528,N_19560);
nand UO_575 (O_575,N_19332,N_19839);
nor UO_576 (O_576,N_19516,N_19923);
and UO_577 (O_577,N_19959,N_19722);
nor UO_578 (O_578,N_19548,N_19570);
and UO_579 (O_579,N_19696,N_19718);
or UO_580 (O_580,N_19650,N_19549);
or UO_581 (O_581,N_19260,N_19660);
or UO_582 (O_582,N_19745,N_19952);
nor UO_583 (O_583,N_19561,N_19784);
or UO_584 (O_584,N_19799,N_19895);
and UO_585 (O_585,N_19726,N_19515);
xnor UO_586 (O_586,N_19923,N_19728);
and UO_587 (O_587,N_19913,N_19392);
and UO_588 (O_588,N_19445,N_19520);
and UO_589 (O_589,N_19371,N_19517);
xnor UO_590 (O_590,N_19532,N_19305);
and UO_591 (O_591,N_19372,N_19853);
and UO_592 (O_592,N_19861,N_19947);
xor UO_593 (O_593,N_19697,N_19227);
xnor UO_594 (O_594,N_19731,N_19217);
nor UO_595 (O_595,N_19635,N_19944);
and UO_596 (O_596,N_19351,N_19488);
nor UO_597 (O_597,N_19952,N_19299);
xor UO_598 (O_598,N_19354,N_19588);
nand UO_599 (O_599,N_19217,N_19437);
or UO_600 (O_600,N_19640,N_19448);
nor UO_601 (O_601,N_19552,N_19559);
nor UO_602 (O_602,N_19771,N_19370);
nand UO_603 (O_603,N_19426,N_19560);
nor UO_604 (O_604,N_19567,N_19539);
nor UO_605 (O_605,N_19971,N_19500);
xnor UO_606 (O_606,N_19498,N_19804);
or UO_607 (O_607,N_19801,N_19482);
nor UO_608 (O_608,N_19784,N_19922);
nor UO_609 (O_609,N_19487,N_19352);
and UO_610 (O_610,N_19680,N_19393);
and UO_611 (O_611,N_19269,N_19747);
and UO_612 (O_612,N_19535,N_19313);
and UO_613 (O_613,N_19974,N_19387);
or UO_614 (O_614,N_19490,N_19597);
or UO_615 (O_615,N_19777,N_19818);
nor UO_616 (O_616,N_19803,N_19447);
or UO_617 (O_617,N_19489,N_19449);
nand UO_618 (O_618,N_19866,N_19766);
and UO_619 (O_619,N_19685,N_19474);
or UO_620 (O_620,N_19840,N_19239);
nand UO_621 (O_621,N_19791,N_19899);
xnor UO_622 (O_622,N_19378,N_19636);
nor UO_623 (O_623,N_19559,N_19647);
xnor UO_624 (O_624,N_19817,N_19982);
and UO_625 (O_625,N_19350,N_19278);
or UO_626 (O_626,N_19373,N_19283);
nand UO_627 (O_627,N_19403,N_19625);
xor UO_628 (O_628,N_19609,N_19803);
or UO_629 (O_629,N_19507,N_19780);
nor UO_630 (O_630,N_19402,N_19709);
nor UO_631 (O_631,N_19657,N_19498);
or UO_632 (O_632,N_19514,N_19250);
and UO_633 (O_633,N_19230,N_19904);
nand UO_634 (O_634,N_19584,N_19640);
nor UO_635 (O_635,N_19921,N_19658);
xor UO_636 (O_636,N_19902,N_19722);
or UO_637 (O_637,N_19714,N_19695);
xor UO_638 (O_638,N_19572,N_19780);
nor UO_639 (O_639,N_19406,N_19262);
xnor UO_640 (O_640,N_19905,N_19783);
xnor UO_641 (O_641,N_19410,N_19944);
and UO_642 (O_642,N_19810,N_19646);
xnor UO_643 (O_643,N_19248,N_19396);
nor UO_644 (O_644,N_19717,N_19236);
nor UO_645 (O_645,N_19946,N_19736);
and UO_646 (O_646,N_19799,N_19617);
nand UO_647 (O_647,N_19320,N_19711);
nand UO_648 (O_648,N_19546,N_19450);
and UO_649 (O_649,N_19875,N_19535);
xnor UO_650 (O_650,N_19252,N_19301);
nor UO_651 (O_651,N_19362,N_19612);
nand UO_652 (O_652,N_19578,N_19417);
nor UO_653 (O_653,N_19526,N_19706);
nor UO_654 (O_654,N_19361,N_19397);
or UO_655 (O_655,N_19458,N_19203);
xor UO_656 (O_656,N_19534,N_19372);
and UO_657 (O_657,N_19539,N_19234);
and UO_658 (O_658,N_19345,N_19517);
or UO_659 (O_659,N_19201,N_19826);
or UO_660 (O_660,N_19761,N_19805);
and UO_661 (O_661,N_19929,N_19296);
xor UO_662 (O_662,N_19756,N_19860);
or UO_663 (O_663,N_19342,N_19968);
and UO_664 (O_664,N_19934,N_19428);
xor UO_665 (O_665,N_19542,N_19894);
and UO_666 (O_666,N_19223,N_19904);
and UO_667 (O_667,N_19387,N_19858);
or UO_668 (O_668,N_19236,N_19967);
xnor UO_669 (O_669,N_19203,N_19601);
nor UO_670 (O_670,N_19228,N_19896);
nor UO_671 (O_671,N_19796,N_19913);
or UO_672 (O_672,N_19955,N_19474);
nand UO_673 (O_673,N_19611,N_19703);
nand UO_674 (O_674,N_19209,N_19315);
nand UO_675 (O_675,N_19853,N_19762);
xor UO_676 (O_676,N_19489,N_19688);
nand UO_677 (O_677,N_19397,N_19810);
and UO_678 (O_678,N_19534,N_19279);
and UO_679 (O_679,N_19519,N_19596);
or UO_680 (O_680,N_19494,N_19836);
nand UO_681 (O_681,N_19924,N_19758);
or UO_682 (O_682,N_19993,N_19801);
nor UO_683 (O_683,N_19238,N_19552);
or UO_684 (O_684,N_19800,N_19772);
nand UO_685 (O_685,N_19293,N_19322);
and UO_686 (O_686,N_19516,N_19750);
nand UO_687 (O_687,N_19309,N_19300);
and UO_688 (O_688,N_19331,N_19589);
and UO_689 (O_689,N_19889,N_19804);
xnor UO_690 (O_690,N_19736,N_19956);
nor UO_691 (O_691,N_19623,N_19445);
and UO_692 (O_692,N_19626,N_19864);
or UO_693 (O_693,N_19900,N_19424);
xor UO_694 (O_694,N_19420,N_19602);
or UO_695 (O_695,N_19220,N_19452);
xor UO_696 (O_696,N_19693,N_19465);
and UO_697 (O_697,N_19262,N_19431);
nand UO_698 (O_698,N_19575,N_19829);
and UO_699 (O_699,N_19536,N_19380);
nand UO_700 (O_700,N_19408,N_19444);
and UO_701 (O_701,N_19897,N_19651);
xnor UO_702 (O_702,N_19293,N_19983);
nand UO_703 (O_703,N_19278,N_19776);
nor UO_704 (O_704,N_19507,N_19839);
nand UO_705 (O_705,N_19941,N_19229);
nand UO_706 (O_706,N_19674,N_19602);
nor UO_707 (O_707,N_19358,N_19631);
xnor UO_708 (O_708,N_19329,N_19650);
xnor UO_709 (O_709,N_19804,N_19639);
xor UO_710 (O_710,N_19960,N_19915);
xnor UO_711 (O_711,N_19205,N_19780);
and UO_712 (O_712,N_19758,N_19614);
xnor UO_713 (O_713,N_19513,N_19255);
nand UO_714 (O_714,N_19249,N_19229);
and UO_715 (O_715,N_19432,N_19333);
nand UO_716 (O_716,N_19925,N_19393);
or UO_717 (O_717,N_19645,N_19737);
nand UO_718 (O_718,N_19430,N_19844);
or UO_719 (O_719,N_19668,N_19910);
and UO_720 (O_720,N_19860,N_19419);
nand UO_721 (O_721,N_19407,N_19291);
or UO_722 (O_722,N_19485,N_19833);
or UO_723 (O_723,N_19691,N_19471);
and UO_724 (O_724,N_19655,N_19393);
or UO_725 (O_725,N_19846,N_19496);
and UO_726 (O_726,N_19617,N_19700);
or UO_727 (O_727,N_19995,N_19342);
xor UO_728 (O_728,N_19379,N_19678);
or UO_729 (O_729,N_19844,N_19221);
nor UO_730 (O_730,N_19846,N_19714);
nand UO_731 (O_731,N_19860,N_19343);
nand UO_732 (O_732,N_19749,N_19397);
xnor UO_733 (O_733,N_19510,N_19845);
nor UO_734 (O_734,N_19861,N_19748);
nor UO_735 (O_735,N_19611,N_19873);
nand UO_736 (O_736,N_19733,N_19695);
nor UO_737 (O_737,N_19731,N_19494);
nor UO_738 (O_738,N_19319,N_19922);
xor UO_739 (O_739,N_19293,N_19269);
nor UO_740 (O_740,N_19744,N_19222);
nand UO_741 (O_741,N_19240,N_19924);
nor UO_742 (O_742,N_19547,N_19868);
nor UO_743 (O_743,N_19368,N_19946);
nor UO_744 (O_744,N_19666,N_19274);
and UO_745 (O_745,N_19612,N_19536);
nand UO_746 (O_746,N_19821,N_19899);
nand UO_747 (O_747,N_19754,N_19697);
nor UO_748 (O_748,N_19349,N_19853);
xnor UO_749 (O_749,N_19520,N_19645);
or UO_750 (O_750,N_19593,N_19711);
or UO_751 (O_751,N_19955,N_19693);
xnor UO_752 (O_752,N_19899,N_19579);
and UO_753 (O_753,N_19944,N_19222);
nand UO_754 (O_754,N_19214,N_19442);
or UO_755 (O_755,N_19692,N_19361);
xnor UO_756 (O_756,N_19587,N_19783);
and UO_757 (O_757,N_19496,N_19524);
or UO_758 (O_758,N_19926,N_19913);
nand UO_759 (O_759,N_19927,N_19650);
xnor UO_760 (O_760,N_19665,N_19254);
or UO_761 (O_761,N_19548,N_19577);
xor UO_762 (O_762,N_19423,N_19913);
nor UO_763 (O_763,N_19849,N_19916);
nor UO_764 (O_764,N_19953,N_19755);
and UO_765 (O_765,N_19738,N_19617);
nor UO_766 (O_766,N_19854,N_19719);
or UO_767 (O_767,N_19378,N_19696);
nand UO_768 (O_768,N_19321,N_19645);
nor UO_769 (O_769,N_19565,N_19862);
or UO_770 (O_770,N_19561,N_19231);
and UO_771 (O_771,N_19356,N_19970);
nor UO_772 (O_772,N_19901,N_19566);
nor UO_773 (O_773,N_19809,N_19230);
xor UO_774 (O_774,N_19590,N_19815);
or UO_775 (O_775,N_19787,N_19801);
nand UO_776 (O_776,N_19948,N_19525);
nor UO_777 (O_777,N_19882,N_19314);
nor UO_778 (O_778,N_19454,N_19265);
and UO_779 (O_779,N_19782,N_19543);
nand UO_780 (O_780,N_19377,N_19825);
nor UO_781 (O_781,N_19830,N_19224);
xnor UO_782 (O_782,N_19815,N_19953);
nand UO_783 (O_783,N_19376,N_19405);
xor UO_784 (O_784,N_19916,N_19271);
and UO_785 (O_785,N_19846,N_19512);
xor UO_786 (O_786,N_19713,N_19457);
and UO_787 (O_787,N_19691,N_19347);
nand UO_788 (O_788,N_19885,N_19337);
nand UO_789 (O_789,N_19990,N_19967);
and UO_790 (O_790,N_19352,N_19920);
xnor UO_791 (O_791,N_19806,N_19734);
nor UO_792 (O_792,N_19718,N_19835);
and UO_793 (O_793,N_19310,N_19960);
nor UO_794 (O_794,N_19456,N_19959);
or UO_795 (O_795,N_19689,N_19915);
and UO_796 (O_796,N_19469,N_19675);
and UO_797 (O_797,N_19348,N_19803);
and UO_798 (O_798,N_19783,N_19939);
or UO_799 (O_799,N_19926,N_19786);
and UO_800 (O_800,N_19807,N_19761);
and UO_801 (O_801,N_19648,N_19763);
nand UO_802 (O_802,N_19715,N_19674);
and UO_803 (O_803,N_19629,N_19874);
nor UO_804 (O_804,N_19322,N_19722);
nor UO_805 (O_805,N_19855,N_19213);
and UO_806 (O_806,N_19249,N_19364);
nor UO_807 (O_807,N_19558,N_19618);
nand UO_808 (O_808,N_19484,N_19547);
nor UO_809 (O_809,N_19769,N_19467);
nor UO_810 (O_810,N_19879,N_19908);
or UO_811 (O_811,N_19526,N_19255);
nand UO_812 (O_812,N_19607,N_19948);
and UO_813 (O_813,N_19312,N_19651);
xnor UO_814 (O_814,N_19654,N_19450);
nor UO_815 (O_815,N_19987,N_19585);
xnor UO_816 (O_816,N_19229,N_19572);
nor UO_817 (O_817,N_19955,N_19450);
and UO_818 (O_818,N_19220,N_19563);
and UO_819 (O_819,N_19501,N_19809);
nand UO_820 (O_820,N_19207,N_19372);
nand UO_821 (O_821,N_19292,N_19966);
or UO_822 (O_822,N_19217,N_19825);
xnor UO_823 (O_823,N_19406,N_19438);
nand UO_824 (O_824,N_19256,N_19624);
or UO_825 (O_825,N_19594,N_19753);
nand UO_826 (O_826,N_19223,N_19839);
nand UO_827 (O_827,N_19619,N_19486);
nor UO_828 (O_828,N_19270,N_19439);
or UO_829 (O_829,N_19258,N_19726);
or UO_830 (O_830,N_19746,N_19892);
xnor UO_831 (O_831,N_19437,N_19424);
nand UO_832 (O_832,N_19671,N_19862);
xor UO_833 (O_833,N_19396,N_19330);
and UO_834 (O_834,N_19655,N_19701);
nor UO_835 (O_835,N_19888,N_19687);
nor UO_836 (O_836,N_19249,N_19493);
and UO_837 (O_837,N_19255,N_19974);
nand UO_838 (O_838,N_19316,N_19272);
nor UO_839 (O_839,N_19439,N_19592);
nor UO_840 (O_840,N_19837,N_19202);
xnor UO_841 (O_841,N_19469,N_19545);
and UO_842 (O_842,N_19404,N_19723);
nand UO_843 (O_843,N_19777,N_19664);
or UO_844 (O_844,N_19659,N_19583);
and UO_845 (O_845,N_19455,N_19998);
xnor UO_846 (O_846,N_19204,N_19614);
and UO_847 (O_847,N_19977,N_19782);
and UO_848 (O_848,N_19769,N_19884);
nor UO_849 (O_849,N_19237,N_19329);
and UO_850 (O_850,N_19386,N_19528);
xnor UO_851 (O_851,N_19243,N_19220);
or UO_852 (O_852,N_19998,N_19468);
nor UO_853 (O_853,N_19824,N_19364);
and UO_854 (O_854,N_19337,N_19387);
xnor UO_855 (O_855,N_19205,N_19519);
nand UO_856 (O_856,N_19608,N_19678);
xor UO_857 (O_857,N_19663,N_19358);
nand UO_858 (O_858,N_19753,N_19806);
xor UO_859 (O_859,N_19883,N_19835);
xor UO_860 (O_860,N_19653,N_19644);
or UO_861 (O_861,N_19923,N_19732);
or UO_862 (O_862,N_19537,N_19842);
and UO_863 (O_863,N_19811,N_19926);
nand UO_864 (O_864,N_19746,N_19995);
nand UO_865 (O_865,N_19831,N_19974);
xnor UO_866 (O_866,N_19200,N_19556);
nand UO_867 (O_867,N_19713,N_19979);
or UO_868 (O_868,N_19857,N_19548);
xnor UO_869 (O_869,N_19503,N_19861);
nand UO_870 (O_870,N_19801,N_19435);
nand UO_871 (O_871,N_19967,N_19371);
and UO_872 (O_872,N_19386,N_19344);
xnor UO_873 (O_873,N_19648,N_19784);
nand UO_874 (O_874,N_19727,N_19614);
xor UO_875 (O_875,N_19442,N_19945);
nor UO_876 (O_876,N_19637,N_19463);
nand UO_877 (O_877,N_19660,N_19521);
xnor UO_878 (O_878,N_19487,N_19547);
nor UO_879 (O_879,N_19942,N_19332);
xor UO_880 (O_880,N_19602,N_19368);
xnor UO_881 (O_881,N_19644,N_19410);
or UO_882 (O_882,N_19633,N_19606);
xor UO_883 (O_883,N_19452,N_19829);
nor UO_884 (O_884,N_19220,N_19493);
nand UO_885 (O_885,N_19513,N_19843);
xor UO_886 (O_886,N_19538,N_19376);
and UO_887 (O_887,N_19277,N_19473);
xor UO_888 (O_888,N_19852,N_19933);
or UO_889 (O_889,N_19907,N_19321);
or UO_890 (O_890,N_19523,N_19584);
nand UO_891 (O_891,N_19353,N_19287);
and UO_892 (O_892,N_19202,N_19419);
nand UO_893 (O_893,N_19705,N_19624);
and UO_894 (O_894,N_19971,N_19817);
nor UO_895 (O_895,N_19866,N_19318);
or UO_896 (O_896,N_19983,N_19572);
xor UO_897 (O_897,N_19898,N_19747);
and UO_898 (O_898,N_19801,N_19311);
and UO_899 (O_899,N_19256,N_19978);
or UO_900 (O_900,N_19291,N_19827);
or UO_901 (O_901,N_19870,N_19978);
nor UO_902 (O_902,N_19374,N_19994);
xor UO_903 (O_903,N_19285,N_19221);
nand UO_904 (O_904,N_19692,N_19654);
nor UO_905 (O_905,N_19960,N_19552);
and UO_906 (O_906,N_19263,N_19797);
nor UO_907 (O_907,N_19650,N_19987);
nor UO_908 (O_908,N_19687,N_19400);
nand UO_909 (O_909,N_19383,N_19201);
or UO_910 (O_910,N_19273,N_19947);
and UO_911 (O_911,N_19686,N_19566);
xnor UO_912 (O_912,N_19845,N_19580);
nor UO_913 (O_913,N_19407,N_19397);
nand UO_914 (O_914,N_19286,N_19249);
xnor UO_915 (O_915,N_19723,N_19705);
nand UO_916 (O_916,N_19557,N_19273);
nand UO_917 (O_917,N_19204,N_19863);
nand UO_918 (O_918,N_19438,N_19658);
nor UO_919 (O_919,N_19917,N_19307);
nor UO_920 (O_920,N_19568,N_19559);
or UO_921 (O_921,N_19809,N_19319);
nor UO_922 (O_922,N_19845,N_19619);
nand UO_923 (O_923,N_19202,N_19296);
xor UO_924 (O_924,N_19815,N_19319);
xnor UO_925 (O_925,N_19890,N_19860);
nor UO_926 (O_926,N_19265,N_19674);
nor UO_927 (O_927,N_19776,N_19681);
or UO_928 (O_928,N_19456,N_19699);
or UO_929 (O_929,N_19309,N_19649);
and UO_930 (O_930,N_19423,N_19765);
xnor UO_931 (O_931,N_19452,N_19739);
or UO_932 (O_932,N_19573,N_19778);
nand UO_933 (O_933,N_19375,N_19857);
nor UO_934 (O_934,N_19215,N_19830);
nand UO_935 (O_935,N_19346,N_19926);
xor UO_936 (O_936,N_19382,N_19599);
xnor UO_937 (O_937,N_19230,N_19978);
nor UO_938 (O_938,N_19791,N_19641);
or UO_939 (O_939,N_19418,N_19905);
nor UO_940 (O_940,N_19307,N_19246);
or UO_941 (O_941,N_19355,N_19391);
xnor UO_942 (O_942,N_19478,N_19967);
or UO_943 (O_943,N_19731,N_19339);
nand UO_944 (O_944,N_19856,N_19642);
nor UO_945 (O_945,N_19864,N_19314);
nor UO_946 (O_946,N_19398,N_19535);
and UO_947 (O_947,N_19692,N_19384);
xor UO_948 (O_948,N_19550,N_19761);
nor UO_949 (O_949,N_19905,N_19578);
nor UO_950 (O_950,N_19976,N_19415);
xor UO_951 (O_951,N_19534,N_19422);
xnor UO_952 (O_952,N_19860,N_19868);
nand UO_953 (O_953,N_19499,N_19626);
xnor UO_954 (O_954,N_19899,N_19722);
and UO_955 (O_955,N_19459,N_19665);
nand UO_956 (O_956,N_19367,N_19544);
and UO_957 (O_957,N_19519,N_19420);
and UO_958 (O_958,N_19740,N_19562);
and UO_959 (O_959,N_19999,N_19430);
nand UO_960 (O_960,N_19473,N_19635);
and UO_961 (O_961,N_19370,N_19888);
nand UO_962 (O_962,N_19624,N_19323);
nand UO_963 (O_963,N_19849,N_19918);
or UO_964 (O_964,N_19476,N_19966);
nor UO_965 (O_965,N_19238,N_19263);
nor UO_966 (O_966,N_19430,N_19332);
nand UO_967 (O_967,N_19336,N_19361);
or UO_968 (O_968,N_19923,N_19543);
or UO_969 (O_969,N_19266,N_19298);
nor UO_970 (O_970,N_19690,N_19348);
or UO_971 (O_971,N_19940,N_19501);
and UO_972 (O_972,N_19384,N_19643);
xor UO_973 (O_973,N_19859,N_19204);
and UO_974 (O_974,N_19427,N_19521);
xor UO_975 (O_975,N_19466,N_19829);
nor UO_976 (O_976,N_19848,N_19761);
nor UO_977 (O_977,N_19818,N_19956);
and UO_978 (O_978,N_19902,N_19567);
nor UO_979 (O_979,N_19474,N_19776);
xnor UO_980 (O_980,N_19647,N_19471);
and UO_981 (O_981,N_19897,N_19889);
and UO_982 (O_982,N_19602,N_19256);
xor UO_983 (O_983,N_19908,N_19575);
and UO_984 (O_984,N_19350,N_19705);
nand UO_985 (O_985,N_19952,N_19571);
xor UO_986 (O_986,N_19849,N_19922);
and UO_987 (O_987,N_19477,N_19455);
or UO_988 (O_988,N_19782,N_19892);
and UO_989 (O_989,N_19646,N_19385);
nor UO_990 (O_990,N_19434,N_19746);
nor UO_991 (O_991,N_19898,N_19930);
xor UO_992 (O_992,N_19493,N_19953);
or UO_993 (O_993,N_19849,N_19931);
nand UO_994 (O_994,N_19890,N_19422);
nor UO_995 (O_995,N_19838,N_19318);
nor UO_996 (O_996,N_19996,N_19910);
or UO_997 (O_997,N_19465,N_19832);
nand UO_998 (O_998,N_19364,N_19929);
nor UO_999 (O_999,N_19571,N_19547);
nor UO_1000 (O_1000,N_19849,N_19251);
xnor UO_1001 (O_1001,N_19301,N_19457);
and UO_1002 (O_1002,N_19318,N_19660);
nand UO_1003 (O_1003,N_19206,N_19866);
xnor UO_1004 (O_1004,N_19689,N_19546);
or UO_1005 (O_1005,N_19326,N_19994);
nor UO_1006 (O_1006,N_19531,N_19556);
or UO_1007 (O_1007,N_19562,N_19885);
xnor UO_1008 (O_1008,N_19624,N_19969);
nor UO_1009 (O_1009,N_19755,N_19238);
and UO_1010 (O_1010,N_19945,N_19872);
nand UO_1011 (O_1011,N_19912,N_19434);
or UO_1012 (O_1012,N_19928,N_19947);
and UO_1013 (O_1013,N_19687,N_19397);
and UO_1014 (O_1014,N_19342,N_19966);
or UO_1015 (O_1015,N_19814,N_19906);
nor UO_1016 (O_1016,N_19555,N_19416);
xor UO_1017 (O_1017,N_19761,N_19711);
and UO_1018 (O_1018,N_19621,N_19977);
nand UO_1019 (O_1019,N_19496,N_19322);
and UO_1020 (O_1020,N_19795,N_19221);
xor UO_1021 (O_1021,N_19793,N_19971);
nor UO_1022 (O_1022,N_19366,N_19581);
and UO_1023 (O_1023,N_19223,N_19389);
nor UO_1024 (O_1024,N_19536,N_19238);
and UO_1025 (O_1025,N_19771,N_19986);
nand UO_1026 (O_1026,N_19211,N_19639);
nor UO_1027 (O_1027,N_19621,N_19949);
nor UO_1028 (O_1028,N_19663,N_19811);
nor UO_1029 (O_1029,N_19963,N_19967);
xor UO_1030 (O_1030,N_19866,N_19386);
nand UO_1031 (O_1031,N_19377,N_19849);
or UO_1032 (O_1032,N_19699,N_19806);
or UO_1033 (O_1033,N_19516,N_19701);
nor UO_1034 (O_1034,N_19653,N_19343);
or UO_1035 (O_1035,N_19934,N_19206);
nor UO_1036 (O_1036,N_19925,N_19816);
and UO_1037 (O_1037,N_19458,N_19808);
and UO_1038 (O_1038,N_19341,N_19296);
nand UO_1039 (O_1039,N_19872,N_19759);
or UO_1040 (O_1040,N_19958,N_19950);
nor UO_1041 (O_1041,N_19739,N_19539);
and UO_1042 (O_1042,N_19215,N_19474);
and UO_1043 (O_1043,N_19343,N_19986);
nand UO_1044 (O_1044,N_19409,N_19276);
or UO_1045 (O_1045,N_19854,N_19727);
or UO_1046 (O_1046,N_19372,N_19558);
or UO_1047 (O_1047,N_19310,N_19753);
xnor UO_1048 (O_1048,N_19890,N_19596);
xor UO_1049 (O_1049,N_19480,N_19748);
nor UO_1050 (O_1050,N_19617,N_19820);
nor UO_1051 (O_1051,N_19969,N_19220);
and UO_1052 (O_1052,N_19602,N_19923);
xnor UO_1053 (O_1053,N_19656,N_19828);
xnor UO_1054 (O_1054,N_19573,N_19633);
xnor UO_1055 (O_1055,N_19445,N_19253);
and UO_1056 (O_1056,N_19910,N_19419);
or UO_1057 (O_1057,N_19313,N_19743);
nand UO_1058 (O_1058,N_19785,N_19704);
nand UO_1059 (O_1059,N_19456,N_19267);
xnor UO_1060 (O_1060,N_19336,N_19323);
or UO_1061 (O_1061,N_19940,N_19224);
xor UO_1062 (O_1062,N_19289,N_19462);
and UO_1063 (O_1063,N_19671,N_19910);
or UO_1064 (O_1064,N_19762,N_19468);
nand UO_1065 (O_1065,N_19275,N_19396);
or UO_1066 (O_1066,N_19962,N_19997);
and UO_1067 (O_1067,N_19493,N_19410);
xnor UO_1068 (O_1068,N_19352,N_19309);
or UO_1069 (O_1069,N_19260,N_19524);
and UO_1070 (O_1070,N_19447,N_19578);
xor UO_1071 (O_1071,N_19283,N_19383);
nand UO_1072 (O_1072,N_19955,N_19377);
nor UO_1073 (O_1073,N_19818,N_19462);
xnor UO_1074 (O_1074,N_19769,N_19423);
or UO_1075 (O_1075,N_19929,N_19355);
or UO_1076 (O_1076,N_19645,N_19412);
or UO_1077 (O_1077,N_19798,N_19353);
nand UO_1078 (O_1078,N_19620,N_19875);
and UO_1079 (O_1079,N_19226,N_19890);
or UO_1080 (O_1080,N_19791,N_19767);
nand UO_1081 (O_1081,N_19458,N_19213);
or UO_1082 (O_1082,N_19721,N_19816);
nor UO_1083 (O_1083,N_19259,N_19996);
and UO_1084 (O_1084,N_19381,N_19295);
nor UO_1085 (O_1085,N_19778,N_19900);
xor UO_1086 (O_1086,N_19667,N_19844);
nor UO_1087 (O_1087,N_19486,N_19946);
or UO_1088 (O_1088,N_19866,N_19265);
nand UO_1089 (O_1089,N_19273,N_19634);
xnor UO_1090 (O_1090,N_19632,N_19246);
nand UO_1091 (O_1091,N_19205,N_19245);
xor UO_1092 (O_1092,N_19988,N_19862);
nor UO_1093 (O_1093,N_19920,N_19878);
or UO_1094 (O_1094,N_19606,N_19346);
and UO_1095 (O_1095,N_19940,N_19255);
xnor UO_1096 (O_1096,N_19865,N_19872);
and UO_1097 (O_1097,N_19872,N_19819);
nand UO_1098 (O_1098,N_19914,N_19282);
nand UO_1099 (O_1099,N_19670,N_19938);
or UO_1100 (O_1100,N_19851,N_19908);
and UO_1101 (O_1101,N_19419,N_19765);
and UO_1102 (O_1102,N_19887,N_19354);
nand UO_1103 (O_1103,N_19642,N_19730);
or UO_1104 (O_1104,N_19358,N_19846);
and UO_1105 (O_1105,N_19736,N_19201);
nand UO_1106 (O_1106,N_19807,N_19780);
and UO_1107 (O_1107,N_19912,N_19598);
nor UO_1108 (O_1108,N_19971,N_19430);
xnor UO_1109 (O_1109,N_19808,N_19962);
xnor UO_1110 (O_1110,N_19954,N_19288);
nor UO_1111 (O_1111,N_19453,N_19259);
nor UO_1112 (O_1112,N_19790,N_19636);
and UO_1113 (O_1113,N_19291,N_19965);
nand UO_1114 (O_1114,N_19469,N_19763);
xnor UO_1115 (O_1115,N_19364,N_19829);
nor UO_1116 (O_1116,N_19464,N_19347);
or UO_1117 (O_1117,N_19693,N_19768);
nor UO_1118 (O_1118,N_19494,N_19510);
nand UO_1119 (O_1119,N_19329,N_19400);
xor UO_1120 (O_1120,N_19650,N_19315);
or UO_1121 (O_1121,N_19987,N_19633);
or UO_1122 (O_1122,N_19571,N_19401);
and UO_1123 (O_1123,N_19731,N_19513);
and UO_1124 (O_1124,N_19983,N_19564);
nor UO_1125 (O_1125,N_19225,N_19272);
nor UO_1126 (O_1126,N_19310,N_19912);
xnor UO_1127 (O_1127,N_19771,N_19376);
nand UO_1128 (O_1128,N_19280,N_19745);
nor UO_1129 (O_1129,N_19745,N_19898);
nor UO_1130 (O_1130,N_19280,N_19651);
and UO_1131 (O_1131,N_19618,N_19727);
and UO_1132 (O_1132,N_19213,N_19931);
nand UO_1133 (O_1133,N_19353,N_19463);
nor UO_1134 (O_1134,N_19330,N_19569);
xnor UO_1135 (O_1135,N_19228,N_19486);
and UO_1136 (O_1136,N_19367,N_19769);
and UO_1137 (O_1137,N_19862,N_19481);
nand UO_1138 (O_1138,N_19983,N_19609);
and UO_1139 (O_1139,N_19919,N_19914);
nand UO_1140 (O_1140,N_19676,N_19991);
and UO_1141 (O_1141,N_19514,N_19660);
or UO_1142 (O_1142,N_19231,N_19859);
and UO_1143 (O_1143,N_19628,N_19704);
or UO_1144 (O_1144,N_19486,N_19852);
nand UO_1145 (O_1145,N_19844,N_19764);
xor UO_1146 (O_1146,N_19299,N_19637);
nor UO_1147 (O_1147,N_19943,N_19913);
nand UO_1148 (O_1148,N_19959,N_19746);
and UO_1149 (O_1149,N_19670,N_19992);
xnor UO_1150 (O_1150,N_19502,N_19537);
xor UO_1151 (O_1151,N_19910,N_19657);
or UO_1152 (O_1152,N_19891,N_19839);
nand UO_1153 (O_1153,N_19519,N_19961);
or UO_1154 (O_1154,N_19796,N_19792);
xor UO_1155 (O_1155,N_19920,N_19699);
xnor UO_1156 (O_1156,N_19637,N_19623);
nand UO_1157 (O_1157,N_19658,N_19640);
and UO_1158 (O_1158,N_19441,N_19683);
or UO_1159 (O_1159,N_19710,N_19589);
xnor UO_1160 (O_1160,N_19526,N_19733);
xor UO_1161 (O_1161,N_19692,N_19676);
or UO_1162 (O_1162,N_19621,N_19515);
or UO_1163 (O_1163,N_19274,N_19992);
xor UO_1164 (O_1164,N_19541,N_19961);
nand UO_1165 (O_1165,N_19330,N_19944);
or UO_1166 (O_1166,N_19555,N_19809);
xor UO_1167 (O_1167,N_19293,N_19523);
xor UO_1168 (O_1168,N_19575,N_19301);
nand UO_1169 (O_1169,N_19400,N_19541);
nor UO_1170 (O_1170,N_19859,N_19533);
or UO_1171 (O_1171,N_19864,N_19679);
nand UO_1172 (O_1172,N_19404,N_19958);
nor UO_1173 (O_1173,N_19964,N_19924);
xnor UO_1174 (O_1174,N_19276,N_19990);
nand UO_1175 (O_1175,N_19720,N_19315);
xor UO_1176 (O_1176,N_19499,N_19261);
nor UO_1177 (O_1177,N_19727,N_19203);
nor UO_1178 (O_1178,N_19976,N_19523);
nor UO_1179 (O_1179,N_19337,N_19973);
or UO_1180 (O_1180,N_19513,N_19973);
xnor UO_1181 (O_1181,N_19566,N_19436);
and UO_1182 (O_1182,N_19706,N_19812);
or UO_1183 (O_1183,N_19791,N_19881);
xor UO_1184 (O_1184,N_19275,N_19608);
or UO_1185 (O_1185,N_19935,N_19245);
nor UO_1186 (O_1186,N_19716,N_19996);
nand UO_1187 (O_1187,N_19870,N_19678);
or UO_1188 (O_1188,N_19743,N_19401);
nand UO_1189 (O_1189,N_19455,N_19703);
nor UO_1190 (O_1190,N_19572,N_19885);
and UO_1191 (O_1191,N_19996,N_19991);
xnor UO_1192 (O_1192,N_19275,N_19638);
nand UO_1193 (O_1193,N_19201,N_19849);
or UO_1194 (O_1194,N_19310,N_19961);
xnor UO_1195 (O_1195,N_19927,N_19681);
nand UO_1196 (O_1196,N_19887,N_19368);
xnor UO_1197 (O_1197,N_19395,N_19671);
xor UO_1198 (O_1198,N_19300,N_19360);
xor UO_1199 (O_1199,N_19999,N_19289);
and UO_1200 (O_1200,N_19753,N_19514);
and UO_1201 (O_1201,N_19942,N_19226);
and UO_1202 (O_1202,N_19223,N_19556);
nor UO_1203 (O_1203,N_19651,N_19244);
or UO_1204 (O_1204,N_19562,N_19631);
xnor UO_1205 (O_1205,N_19730,N_19976);
nor UO_1206 (O_1206,N_19620,N_19943);
xor UO_1207 (O_1207,N_19946,N_19624);
nand UO_1208 (O_1208,N_19999,N_19262);
and UO_1209 (O_1209,N_19223,N_19384);
nor UO_1210 (O_1210,N_19886,N_19871);
nor UO_1211 (O_1211,N_19269,N_19619);
nand UO_1212 (O_1212,N_19822,N_19541);
xnor UO_1213 (O_1213,N_19433,N_19962);
nor UO_1214 (O_1214,N_19640,N_19555);
xor UO_1215 (O_1215,N_19869,N_19320);
nand UO_1216 (O_1216,N_19350,N_19987);
xor UO_1217 (O_1217,N_19919,N_19478);
xnor UO_1218 (O_1218,N_19368,N_19337);
or UO_1219 (O_1219,N_19920,N_19876);
or UO_1220 (O_1220,N_19707,N_19207);
or UO_1221 (O_1221,N_19270,N_19262);
and UO_1222 (O_1222,N_19277,N_19354);
nor UO_1223 (O_1223,N_19620,N_19643);
and UO_1224 (O_1224,N_19879,N_19901);
and UO_1225 (O_1225,N_19278,N_19268);
or UO_1226 (O_1226,N_19601,N_19779);
xor UO_1227 (O_1227,N_19426,N_19443);
nor UO_1228 (O_1228,N_19218,N_19236);
xor UO_1229 (O_1229,N_19284,N_19769);
nor UO_1230 (O_1230,N_19506,N_19620);
xor UO_1231 (O_1231,N_19815,N_19702);
nand UO_1232 (O_1232,N_19775,N_19808);
or UO_1233 (O_1233,N_19621,N_19366);
nand UO_1234 (O_1234,N_19707,N_19581);
xnor UO_1235 (O_1235,N_19866,N_19788);
and UO_1236 (O_1236,N_19642,N_19607);
xnor UO_1237 (O_1237,N_19307,N_19346);
xor UO_1238 (O_1238,N_19594,N_19516);
or UO_1239 (O_1239,N_19414,N_19975);
and UO_1240 (O_1240,N_19620,N_19663);
or UO_1241 (O_1241,N_19427,N_19308);
nor UO_1242 (O_1242,N_19604,N_19517);
or UO_1243 (O_1243,N_19833,N_19274);
and UO_1244 (O_1244,N_19966,N_19872);
xor UO_1245 (O_1245,N_19699,N_19762);
xor UO_1246 (O_1246,N_19647,N_19253);
and UO_1247 (O_1247,N_19729,N_19843);
or UO_1248 (O_1248,N_19588,N_19784);
nor UO_1249 (O_1249,N_19747,N_19761);
nand UO_1250 (O_1250,N_19337,N_19444);
nor UO_1251 (O_1251,N_19546,N_19971);
nor UO_1252 (O_1252,N_19704,N_19827);
nand UO_1253 (O_1253,N_19488,N_19802);
or UO_1254 (O_1254,N_19618,N_19435);
nor UO_1255 (O_1255,N_19779,N_19862);
and UO_1256 (O_1256,N_19854,N_19502);
and UO_1257 (O_1257,N_19223,N_19440);
nand UO_1258 (O_1258,N_19323,N_19375);
or UO_1259 (O_1259,N_19986,N_19412);
or UO_1260 (O_1260,N_19259,N_19436);
or UO_1261 (O_1261,N_19856,N_19346);
xnor UO_1262 (O_1262,N_19583,N_19710);
nand UO_1263 (O_1263,N_19963,N_19316);
and UO_1264 (O_1264,N_19348,N_19424);
xnor UO_1265 (O_1265,N_19946,N_19349);
or UO_1266 (O_1266,N_19795,N_19309);
xor UO_1267 (O_1267,N_19484,N_19569);
or UO_1268 (O_1268,N_19357,N_19310);
nor UO_1269 (O_1269,N_19548,N_19677);
or UO_1270 (O_1270,N_19626,N_19834);
xor UO_1271 (O_1271,N_19399,N_19361);
nor UO_1272 (O_1272,N_19387,N_19470);
and UO_1273 (O_1273,N_19767,N_19276);
or UO_1274 (O_1274,N_19229,N_19802);
xnor UO_1275 (O_1275,N_19366,N_19384);
and UO_1276 (O_1276,N_19443,N_19357);
or UO_1277 (O_1277,N_19717,N_19241);
nand UO_1278 (O_1278,N_19979,N_19553);
nand UO_1279 (O_1279,N_19726,N_19757);
nand UO_1280 (O_1280,N_19932,N_19959);
xnor UO_1281 (O_1281,N_19910,N_19284);
xnor UO_1282 (O_1282,N_19315,N_19928);
nor UO_1283 (O_1283,N_19225,N_19887);
or UO_1284 (O_1284,N_19329,N_19854);
nand UO_1285 (O_1285,N_19770,N_19543);
or UO_1286 (O_1286,N_19253,N_19985);
nor UO_1287 (O_1287,N_19209,N_19376);
nor UO_1288 (O_1288,N_19587,N_19232);
and UO_1289 (O_1289,N_19398,N_19486);
nand UO_1290 (O_1290,N_19270,N_19426);
nand UO_1291 (O_1291,N_19791,N_19866);
nand UO_1292 (O_1292,N_19940,N_19251);
nand UO_1293 (O_1293,N_19271,N_19909);
nand UO_1294 (O_1294,N_19977,N_19673);
and UO_1295 (O_1295,N_19872,N_19616);
or UO_1296 (O_1296,N_19416,N_19998);
nand UO_1297 (O_1297,N_19884,N_19604);
nor UO_1298 (O_1298,N_19821,N_19919);
or UO_1299 (O_1299,N_19219,N_19267);
xor UO_1300 (O_1300,N_19417,N_19932);
or UO_1301 (O_1301,N_19726,N_19931);
nor UO_1302 (O_1302,N_19720,N_19577);
and UO_1303 (O_1303,N_19752,N_19647);
xor UO_1304 (O_1304,N_19654,N_19815);
nor UO_1305 (O_1305,N_19797,N_19336);
and UO_1306 (O_1306,N_19860,N_19686);
and UO_1307 (O_1307,N_19820,N_19897);
nor UO_1308 (O_1308,N_19404,N_19542);
or UO_1309 (O_1309,N_19986,N_19563);
nor UO_1310 (O_1310,N_19821,N_19401);
or UO_1311 (O_1311,N_19821,N_19888);
nand UO_1312 (O_1312,N_19803,N_19735);
xnor UO_1313 (O_1313,N_19996,N_19862);
and UO_1314 (O_1314,N_19537,N_19458);
and UO_1315 (O_1315,N_19582,N_19221);
nor UO_1316 (O_1316,N_19977,N_19825);
xnor UO_1317 (O_1317,N_19717,N_19675);
or UO_1318 (O_1318,N_19954,N_19857);
or UO_1319 (O_1319,N_19413,N_19310);
and UO_1320 (O_1320,N_19596,N_19701);
nand UO_1321 (O_1321,N_19530,N_19427);
or UO_1322 (O_1322,N_19375,N_19599);
xnor UO_1323 (O_1323,N_19581,N_19565);
and UO_1324 (O_1324,N_19666,N_19951);
and UO_1325 (O_1325,N_19561,N_19315);
xnor UO_1326 (O_1326,N_19241,N_19894);
and UO_1327 (O_1327,N_19338,N_19871);
nor UO_1328 (O_1328,N_19704,N_19626);
nand UO_1329 (O_1329,N_19657,N_19224);
nand UO_1330 (O_1330,N_19428,N_19249);
and UO_1331 (O_1331,N_19392,N_19763);
xor UO_1332 (O_1332,N_19870,N_19324);
xor UO_1333 (O_1333,N_19448,N_19705);
nor UO_1334 (O_1334,N_19639,N_19461);
nor UO_1335 (O_1335,N_19210,N_19927);
nand UO_1336 (O_1336,N_19210,N_19297);
and UO_1337 (O_1337,N_19432,N_19886);
nor UO_1338 (O_1338,N_19245,N_19417);
and UO_1339 (O_1339,N_19731,N_19905);
and UO_1340 (O_1340,N_19957,N_19873);
xor UO_1341 (O_1341,N_19784,N_19615);
nor UO_1342 (O_1342,N_19744,N_19711);
nor UO_1343 (O_1343,N_19685,N_19265);
nor UO_1344 (O_1344,N_19818,N_19640);
and UO_1345 (O_1345,N_19678,N_19778);
nor UO_1346 (O_1346,N_19959,N_19254);
nor UO_1347 (O_1347,N_19455,N_19672);
nand UO_1348 (O_1348,N_19564,N_19664);
nand UO_1349 (O_1349,N_19506,N_19681);
xnor UO_1350 (O_1350,N_19817,N_19413);
nor UO_1351 (O_1351,N_19489,N_19234);
nor UO_1352 (O_1352,N_19658,N_19986);
and UO_1353 (O_1353,N_19371,N_19790);
nand UO_1354 (O_1354,N_19269,N_19297);
and UO_1355 (O_1355,N_19242,N_19932);
or UO_1356 (O_1356,N_19560,N_19824);
nand UO_1357 (O_1357,N_19507,N_19460);
or UO_1358 (O_1358,N_19207,N_19630);
xnor UO_1359 (O_1359,N_19731,N_19664);
xor UO_1360 (O_1360,N_19602,N_19924);
and UO_1361 (O_1361,N_19247,N_19589);
or UO_1362 (O_1362,N_19407,N_19238);
nand UO_1363 (O_1363,N_19203,N_19652);
nand UO_1364 (O_1364,N_19601,N_19565);
or UO_1365 (O_1365,N_19416,N_19649);
nor UO_1366 (O_1366,N_19631,N_19910);
nand UO_1367 (O_1367,N_19736,N_19951);
or UO_1368 (O_1368,N_19257,N_19355);
xor UO_1369 (O_1369,N_19666,N_19311);
or UO_1370 (O_1370,N_19570,N_19633);
and UO_1371 (O_1371,N_19268,N_19679);
nand UO_1372 (O_1372,N_19362,N_19808);
nand UO_1373 (O_1373,N_19482,N_19438);
xor UO_1374 (O_1374,N_19629,N_19859);
and UO_1375 (O_1375,N_19667,N_19895);
and UO_1376 (O_1376,N_19631,N_19859);
xnor UO_1377 (O_1377,N_19895,N_19440);
or UO_1378 (O_1378,N_19916,N_19436);
nand UO_1379 (O_1379,N_19681,N_19989);
or UO_1380 (O_1380,N_19372,N_19324);
and UO_1381 (O_1381,N_19682,N_19302);
nor UO_1382 (O_1382,N_19495,N_19245);
or UO_1383 (O_1383,N_19612,N_19222);
and UO_1384 (O_1384,N_19673,N_19503);
nor UO_1385 (O_1385,N_19975,N_19796);
nor UO_1386 (O_1386,N_19640,N_19998);
xnor UO_1387 (O_1387,N_19819,N_19885);
nor UO_1388 (O_1388,N_19686,N_19791);
or UO_1389 (O_1389,N_19498,N_19436);
nor UO_1390 (O_1390,N_19271,N_19929);
and UO_1391 (O_1391,N_19967,N_19756);
or UO_1392 (O_1392,N_19858,N_19333);
nor UO_1393 (O_1393,N_19848,N_19389);
nand UO_1394 (O_1394,N_19508,N_19521);
xor UO_1395 (O_1395,N_19404,N_19649);
nand UO_1396 (O_1396,N_19525,N_19752);
xor UO_1397 (O_1397,N_19581,N_19747);
or UO_1398 (O_1398,N_19823,N_19806);
and UO_1399 (O_1399,N_19651,N_19228);
nand UO_1400 (O_1400,N_19610,N_19803);
or UO_1401 (O_1401,N_19722,N_19602);
nor UO_1402 (O_1402,N_19601,N_19281);
or UO_1403 (O_1403,N_19415,N_19524);
or UO_1404 (O_1404,N_19697,N_19966);
and UO_1405 (O_1405,N_19549,N_19456);
nor UO_1406 (O_1406,N_19237,N_19717);
xor UO_1407 (O_1407,N_19857,N_19560);
or UO_1408 (O_1408,N_19921,N_19909);
xor UO_1409 (O_1409,N_19946,N_19958);
nor UO_1410 (O_1410,N_19884,N_19550);
or UO_1411 (O_1411,N_19707,N_19476);
xor UO_1412 (O_1412,N_19509,N_19336);
nor UO_1413 (O_1413,N_19686,N_19958);
xnor UO_1414 (O_1414,N_19693,N_19852);
xnor UO_1415 (O_1415,N_19621,N_19557);
or UO_1416 (O_1416,N_19792,N_19429);
xnor UO_1417 (O_1417,N_19512,N_19401);
or UO_1418 (O_1418,N_19239,N_19600);
or UO_1419 (O_1419,N_19235,N_19878);
xnor UO_1420 (O_1420,N_19469,N_19230);
and UO_1421 (O_1421,N_19612,N_19655);
nor UO_1422 (O_1422,N_19767,N_19673);
nor UO_1423 (O_1423,N_19922,N_19643);
nor UO_1424 (O_1424,N_19873,N_19679);
nor UO_1425 (O_1425,N_19420,N_19607);
xor UO_1426 (O_1426,N_19385,N_19363);
or UO_1427 (O_1427,N_19968,N_19598);
nor UO_1428 (O_1428,N_19492,N_19612);
and UO_1429 (O_1429,N_19529,N_19892);
nand UO_1430 (O_1430,N_19830,N_19234);
nand UO_1431 (O_1431,N_19312,N_19974);
and UO_1432 (O_1432,N_19974,N_19663);
or UO_1433 (O_1433,N_19905,N_19463);
nand UO_1434 (O_1434,N_19268,N_19242);
and UO_1435 (O_1435,N_19665,N_19253);
xnor UO_1436 (O_1436,N_19518,N_19889);
xor UO_1437 (O_1437,N_19835,N_19480);
and UO_1438 (O_1438,N_19363,N_19957);
and UO_1439 (O_1439,N_19368,N_19495);
or UO_1440 (O_1440,N_19516,N_19908);
xnor UO_1441 (O_1441,N_19779,N_19994);
or UO_1442 (O_1442,N_19935,N_19240);
xnor UO_1443 (O_1443,N_19443,N_19586);
or UO_1444 (O_1444,N_19448,N_19434);
or UO_1445 (O_1445,N_19220,N_19277);
and UO_1446 (O_1446,N_19661,N_19826);
or UO_1447 (O_1447,N_19937,N_19614);
nand UO_1448 (O_1448,N_19836,N_19734);
nor UO_1449 (O_1449,N_19270,N_19226);
xnor UO_1450 (O_1450,N_19602,N_19684);
nand UO_1451 (O_1451,N_19723,N_19375);
and UO_1452 (O_1452,N_19505,N_19933);
and UO_1453 (O_1453,N_19973,N_19425);
and UO_1454 (O_1454,N_19526,N_19524);
nand UO_1455 (O_1455,N_19208,N_19596);
nor UO_1456 (O_1456,N_19688,N_19254);
nor UO_1457 (O_1457,N_19794,N_19748);
nor UO_1458 (O_1458,N_19303,N_19776);
nand UO_1459 (O_1459,N_19495,N_19566);
xnor UO_1460 (O_1460,N_19336,N_19753);
xor UO_1461 (O_1461,N_19324,N_19976);
nor UO_1462 (O_1462,N_19982,N_19325);
and UO_1463 (O_1463,N_19262,N_19708);
nor UO_1464 (O_1464,N_19662,N_19278);
xor UO_1465 (O_1465,N_19801,N_19356);
xor UO_1466 (O_1466,N_19789,N_19967);
xnor UO_1467 (O_1467,N_19738,N_19360);
or UO_1468 (O_1468,N_19508,N_19445);
and UO_1469 (O_1469,N_19846,N_19807);
and UO_1470 (O_1470,N_19442,N_19569);
and UO_1471 (O_1471,N_19317,N_19930);
nor UO_1472 (O_1472,N_19861,N_19597);
nor UO_1473 (O_1473,N_19508,N_19805);
xnor UO_1474 (O_1474,N_19712,N_19232);
nor UO_1475 (O_1475,N_19585,N_19562);
xor UO_1476 (O_1476,N_19989,N_19598);
and UO_1477 (O_1477,N_19743,N_19920);
nor UO_1478 (O_1478,N_19460,N_19585);
nor UO_1479 (O_1479,N_19899,N_19383);
nor UO_1480 (O_1480,N_19943,N_19589);
nor UO_1481 (O_1481,N_19516,N_19432);
or UO_1482 (O_1482,N_19279,N_19404);
or UO_1483 (O_1483,N_19556,N_19312);
and UO_1484 (O_1484,N_19559,N_19487);
and UO_1485 (O_1485,N_19540,N_19310);
nand UO_1486 (O_1486,N_19604,N_19721);
or UO_1487 (O_1487,N_19513,N_19482);
or UO_1488 (O_1488,N_19322,N_19483);
nor UO_1489 (O_1489,N_19232,N_19653);
and UO_1490 (O_1490,N_19699,N_19818);
and UO_1491 (O_1491,N_19219,N_19226);
nand UO_1492 (O_1492,N_19741,N_19826);
xor UO_1493 (O_1493,N_19586,N_19449);
nor UO_1494 (O_1494,N_19380,N_19724);
xor UO_1495 (O_1495,N_19758,N_19832);
or UO_1496 (O_1496,N_19507,N_19804);
nand UO_1497 (O_1497,N_19812,N_19690);
nand UO_1498 (O_1498,N_19672,N_19391);
xor UO_1499 (O_1499,N_19563,N_19704);
nand UO_1500 (O_1500,N_19562,N_19319);
nand UO_1501 (O_1501,N_19643,N_19496);
nor UO_1502 (O_1502,N_19908,N_19824);
xor UO_1503 (O_1503,N_19347,N_19994);
and UO_1504 (O_1504,N_19858,N_19819);
nor UO_1505 (O_1505,N_19751,N_19909);
nor UO_1506 (O_1506,N_19748,N_19414);
and UO_1507 (O_1507,N_19229,N_19732);
or UO_1508 (O_1508,N_19310,N_19484);
nand UO_1509 (O_1509,N_19441,N_19316);
xor UO_1510 (O_1510,N_19255,N_19626);
nand UO_1511 (O_1511,N_19653,N_19848);
nor UO_1512 (O_1512,N_19352,N_19256);
xnor UO_1513 (O_1513,N_19768,N_19579);
nor UO_1514 (O_1514,N_19499,N_19320);
nand UO_1515 (O_1515,N_19376,N_19521);
and UO_1516 (O_1516,N_19546,N_19746);
and UO_1517 (O_1517,N_19350,N_19529);
and UO_1518 (O_1518,N_19844,N_19587);
or UO_1519 (O_1519,N_19269,N_19278);
or UO_1520 (O_1520,N_19362,N_19503);
nor UO_1521 (O_1521,N_19873,N_19507);
and UO_1522 (O_1522,N_19426,N_19967);
nor UO_1523 (O_1523,N_19495,N_19772);
or UO_1524 (O_1524,N_19407,N_19577);
nand UO_1525 (O_1525,N_19441,N_19344);
nand UO_1526 (O_1526,N_19927,N_19497);
nand UO_1527 (O_1527,N_19520,N_19996);
nand UO_1528 (O_1528,N_19809,N_19412);
xnor UO_1529 (O_1529,N_19556,N_19982);
xor UO_1530 (O_1530,N_19417,N_19688);
xnor UO_1531 (O_1531,N_19341,N_19241);
xor UO_1532 (O_1532,N_19459,N_19760);
and UO_1533 (O_1533,N_19957,N_19712);
nor UO_1534 (O_1534,N_19624,N_19385);
xnor UO_1535 (O_1535,N_19482,N_19882);
nand UO_1536 (O_1536,N_19986,N_19273);
nor UO_1537 (O_1537,N_19986,N_19285);
nand UO_1538 (O_1538,N_19271,N_19842);
and UO_1539 (O_1539,N_19585,N_19715);
or UO_1540 (O_1540,N_19234,N_19426);
nor UO_1541 (O_1541,N_19871,N_19544);
nand UO_1542 (O_1542,N_19494,N_19788);
nor UO_1543 (O_1543,N_19980,N_19953);
nand UO_1544 (O_1544,N_19963,N_19545);
or UO_1545 (O_1545,N_19215,N_19523);
or UO_1546 (O_1546,N_19900,N_19473);
or UO_1547 (O_1547,N_19381,N_19747);
or UO_1548 (O_1548,N_19455,N_19799);
or UO_1549 (O_1549,N_19222,N_19503);
nand UO_1550 (O_1550,N_19402,N_19202);
and UO_1551 (O_1551,N_19889,N_19477);
nor UO_1552 (O_1552,N_19654,N_19813);
or UO_1553 (O_1553,N_19213,N_19254);
nand UO_1554 (O_1554,N_19683,N_19713);
xor UO_1555 (O_1555,N_19379,N_19573);
or UO_1556 (O_1556,N_19314,N_19839);
nor UO_1557 (O_1557,N_19999,N_19457);
nand UO_1558 (O_1558,N_19476,N_19508);
nand UO_1559 (O_1559,N_19280,N_19614);
xnor UO_1560 (O_1560,N_19426,N_19943);
nand UO_1561 (O_1561,N_19564,N_19934);
or UO_1562 (O_1562,N_19879,N_19552);
and UO_1563 (O_1563,N_19612,N_19823);
or UO_1564 (O_1564,N_19767,N_19712);
nor UO_1565 (O_1565,N_19917,N_19628);
xor UO_1566 (O_1566,N_19251,N_19659);
and UO_1567 (O_1567,N_19752,N_19405);
or UO_1568 (O_1568,N_19477,N_19693);
and UO_1569 (O_1569,N_19861,N_19581);
and UO_1570 (O_1570,N_19377,N_19481);
or UO_1571 (O_1571,N_19730,N_19748);
or UO_1572 (O_1572,N_19987,N_19449);
and UO_1573 (O_1573,N_19480,N_19826);
and UO_1574 (O_1574,N_19592,N_19878);
xor UO_1575 (O_1575,N_19829,N_19662);
xor UO_1576 (O_1576,N_19693,N_19247);
and UO_1577 (O_1577,N_19407,N_19706);
xor UO_1578 (O_1578,N_19521,N_19641);
and UO_1579 (O_1579,N_19450,N_19585);
nand UO_1580 (O_1580,N_19492,N_19913);
or UO_1581 (O_1581,N_19693,N_19834);
and UO_1582 (O_1582,N_19312,N_19477);
or UO_1583 (O_1583,N_19705,N_19628);
or UO_1584 (O_1584,N_19248,N_19765);
nor UO_1585 (O_1585,N_19276,N_19667);
nor UO_1586 (O_1586,N_19817,N_19988);
nand UO_1587 (O_1587,N_19788,N_19458);
nand UO_1588 (O_1588,N_19546,N_19933);
xnor UO_1589 (O_1589,N_19749,N_19443);
nor UO_1590 (O_1590,N_19435,N_19966);
and UO_1591 (O_1591,N_19780,N_19269);
or UO_1592 (O_1592,N_19775,N_19357);
nor UO_1593 (O_1593,N_19771,N_19937);
nand UO_1594 (O_1594,N_19258,N_19333);
nand UO_1595 (O_1595,N_19307,N_19577);
nor UO_1596 (O_1596,N_19448,N_19645);
xor UO_1597 (O_1597,N_19902,N_19270);
or UO_1598 (O_1598,N_19226,N_19941);
nor UO_1599 (O_1599,N_19246,N_19635);
xor UO_1600 (O_1600,N_19271,N_19360);
xnor UO_1601 (O_1601,N_19710,N_19381);
nor UO_1602 (O_1602,N_19560,N_19753);
nor UO_1603 (O_1603,N_19679,N_19738);
or UO_1604 (O_1604,N_19989,N_19591);
nand UO_1605 (O_1605,N_19856,N_19287);
nand UO_1606 (O_1606,N_19827,N_19372);
or UO_1607 (O_1607,N_19576,N_19244);
nor UO_1608 (O_1608,N_19389,N_19707);
xor UO_1609 (O_1609,N_19855,N_19251);
and UO_1610 (O_1610,N_19301,N_19491);
nor UO_1611 (O_1611,N_19625,N_19782);
nand UO_1612 (O_1612,N_19686,N_19363);
and UO_1613 (O_1613,N_19348,N_19563);
and UO_1614 (O_1614,N_19464,N_19618);
xnor UO_1615 (O_1615,N_19995,N_19638);
xnor UO_1616 (O_1616,N_19891,N_19208);
and UO_1617 (O_1617,N_19707,N_19267);
nand UO_1618 (O_1618,N_19239,N_19577);
xnor UO_1619 (O_1619,N_19695,N_19381);
or UO_1620 (O_1620,N_19266,N_19503);
xnor UO_1621 (O_1621,N_19646,N_19834);
nor UO_1622 (O_1622,N_19421,N_19646);
and UO_1623 (O_1623,N_19459,N_19615);
nand UO_1624 (O_1624,N_19876,N_19566);
or UO_1625 (O_1625,N_19351,N_19929);
xnor UO_1626 (O_1626,N_19413,N_19270);
and UO_1627 (O_1627,N_19876,N_19399);
or UO_1628 (O_1628,N_19971,N_19726);
nand UO_1629 (O_1629,N_19525,N_19324);
or UO_1630 (O_1630,N_19211,N_19304);
xnor UO_1631 (O_1631,N_19962,N_19495);
or UO_1632 (O_1632,N_19620,N_19952);
nor UO_1633 (O_1633,N_19808,N_19507);
nor UO_1634 (O_1634,N_19278,N_19446);
or UO_1635 (O_1635,N_19374,N_19610);
nand UO_1636 (O_1636,N_19275,N_19816);
or UO_1637 (O_1637,N_19427,N_19356);
xnor UO_1638 (O_1638,N_19373,N_19673);
nand UO_1639 (O_1639,N_19287,N_19245);
nor UO_1640 (O_1640,N_19848,N_19608);
nor UO_1641 (O_1641,N_19805,N_19818);
xnor UO_1642 (O_1642,N_19250,N_19719);
nor UO_1643 (O_1643,N_19465,N_19291);
nor UO_1644 (O_1644,N_19282,N_19272);
nand UO_1645 (O_1645,N_19236,N_19924);
nand UO_1646 (O_1646,N_19584,N_19434);
and UO_1647 (O_1647,N_19908,N_19595);
nor UO_1648 (O_1648,N_19906,N_19853);
or UO_1649 (O_1649,N_19821,N_19981);
nand UO_1650 (O_1650,N_19920,N_19435);
nor UO_1651 (O_1651,N_19674,N_19629);
and UO_1652 (O_1652,N_19252,N_19663);
nor UO_1653 (O_1653,N_19738,N_19660);
nand UO_1654 (O_1654,N_19647,N_19211);
nor UO_1655 (O_1655,N_19672,N_19980);
nand UO_1656 (O_1656,N_19277,N_19716);
xnor UO_1657 (O_1657,N_19428,N_19637);
or UO_1658 (O_1658,N_19272,N_19307);
nor UO_1659 (O_1659,N_19952,N_19514);
nor UO_1660 (O_1660,N_19795,N_19907);
xnor UO_1661 (O_1661,N_19429,N_19861);
nand UO_1662 (O_1662,N_19633,N_19512);
nor UO_1663 (O_1663,N_19544,N_19299);
or UO_1664 (O_1664,N_19691,N_19975);
or UO_1665 (O_1665,N_19580,N_19961);
and UO_1666 (O_1666,N_19898,N_19923);
xor UO_1667 (O_1667,N_19591,N_19557);
nor UO_1668 (O_1668,N_19269,N_19927);
and UO_1669 (O_1669,N_19647,N_19670);
xnor UO_1670 (O_1670,N_19393,N_19765);
xnor UO_1671 (O_1671,N_19990,N_19908);
and UO_1672 (O_1672,N_19363,N_19922);
or UO_1673 (O_1673,N_19941,N_19977);
xnor UO_1674 (O_1674,N_19213,N_19800);
nor UO_1675 (O_1675,N_19310,N_19457);
nand UO_1676 (O_1676,N_19705,N_19551);
or UO_1677 (O_1677,N_19433,N_19359);
or UO_1678 (O_1678,N_19210,N_19457);
or UO_1679 (O_1679,N_19711,N_19559);
xnor UO_1680 (O_1680,N_19276,N_19799);
and UO_1681 (O_1681,N_19859,N_19831);
or UO_1682 (O_1682,N_19583,N_19812);
and UO_1683 (O_1683,N_19418,N_19787);
and UO_1684 (O_1684,N_19588,N_19924);
nand UO_1685 (O_1685,N_19371,N_19754);
or UO_1686 (O_1686,N_19742,N_19220);
xor UO_1687 (O_1687,N_19995,N_19651);
nor UO_1688 (O_1688,N_19312,N_19913);
nor UO_1689 (O_1689,N_19596,N_19366);
nor UO_1690 (O_1690,N_19579,N_19922);
or UO_1691 (O_1691,N_19711,N_19224);
nand UO_1692 (O_1692,N_19721,N_19242);
and UO_1693 (O_1693,N_19533,N_19724);
or UO_1694 (O_1694,N_19258,N_19987);
nor UO_1695 (O_1695,N_19677,N_19288);
nor UO_1696 (O_1696,N_19214,N_19635);
or UO_1697 (O_1697,N_19426,N_19995);
or UO_1698 (O_1698,N_19580,N_19535);
xnor UO_1699 (O_1699,N_19858,N_19645);
nand UO_1700 (O_1700,N_19662,N_19882);
and UO_1701 (O_1701,N_19904,N_19558);
and UO_1702 (O_1702,N_19768,N_19557);
or UO_1703 (O_1703,N_19558,N_19633);
or UO_1704 (O_1704,N_19659,N_19971);
xnor UO_1705 (O_1705,N_19373,N_19588);
or UO_1706 (O_1706,N_19250,N_19667);
nand UO_1707 (O_1707,N_19764,N_19933);
xnor UO_1708 (O_1708,N_19616,N_19511);
or UO_1709 (O_1709,N_19914,N_19740);
xnor UO_1710 (O_1710,N_19285,N_19240);
and UO_1711 (O_1711,N_19871,N_19854);
nand UO_1712 (O_1712,N_19325,N_19767);
nand UO_1713 (O_1713,N_19222,N_19935);
nor UO_1714 (O_1714,N_19894,N_19363);
nand UO_1715 (O_1715,N_19447,N_19432);
and UO_1716 (O_1716,N_19865,N_19252);
and UO_1717 (O_1717,N_19237,N_19932);
nor UO_1718 (O_1718,N_19617,N_19352);
nand UO_1719 (O_1719,N_19561,N_19463);
or UO_1720 (O_1720,N_19262,N_19363);
nand UO_1721 (O_1721,N_19310,N_19348);
nor UO_1722 (O_1722,N_19895,N_19818);
xnor UO_1723 (O_1723,N_19942,N_19398);
xnor UO_1724 (O_1724,N_19768,N_19915);
and UO_1725 (O_1725,N_19526,N_19896);
nor UO_1726 (O_1726,N_19315,N_19990);
and UO_1727 (O_1727,N_19809,N_19556);
and UO_1728 (O_1728,N_19416,N_19866);
and UO_1729 (O_1729,N_19563,N_19536);
nand UO_1730 (O_1730,N_19576,N_19989);
nor UO_1731 (O_1731,N_19716,N_19431);
nand UO_1732 (O_1732,N_19580,N_19331);
nand UO_1733 (O_1733,N_19643,N_19269);
or UO_1734 (O_1734,N_19405,N_19976);
or UO_1735 (O_1735,N_19673,N_19932);
and UO_1736 (O_1736,N_19826,N_19604);
xnor UO_1737 (O_1737,N_19333,N_19753);
nand UO_1738 (O_1738,N_19768,N_19778);
nor UO_1739 (O_1739,N_19409,N_19690);
nor UO_1740 (O_1740,N_19809,N_19408);
xor UO_1741 (O_1741,N_19416,N_19785);
and UO_1742 (O_1742,N_19838,N_19925);
xnor UO_1743 (O_1743,N_19989,N_19293);
xnor UO_1744 (O_1744,N_19733,N_19539);
xnor UO_1745 (O_1745,N_19600,N_19608);
or UO_1746 (O_1746,N_19799,N_19541);
or UO_1747 (O_1747,N_19546,N_19462);
and UO_1748 (O_1748,N_19443,N_19953);
xnor UO_1749 (O_1749,N_19242,N_19753);
and UO_1750 (O_1750,N_19281,N_19284);
nor UO_1751 (O_1751,N_19850,N_19449);
nor UO_1752 (O_1752,N_19362,N_19532);
or UO_1753 (O_1753,N_19901,N_19812);
nand UO_1754 (O_1754,N_19931,N_19465);
or UO_1755 (O_1755,N_19456,N_19440);
nor UO_1756 (O_1756,N_19610,N_19508);
and UO_1757 (O_1757,N_19408,N_19606);
nor UO_1758 (O_1758,N_19301,N_19584);
and UO_1759 (O_1759,N_19525,N_19787);
and UO_1760 (O_1760,N_19236,N_19249);
or UO_1761 (O_1761,N_19940,N_19972);
or UO_1762 (O_1762,N_19641,N_19971);
nor UO_1763 (O_1763,N_19218,N_19566);
nor UO_1764 (O_1764,N_19245,N_19506);
nand UO_1765 (O_1765,N_19264,N_19341);
or UO_1766 (O_1766,N_19737,N_19553);
nand UO_1767 (O_1767,N_19376,N_19316);
nor UO_1768 (O_1768,N_19467,N_19544);
and UO_1769 (O_1769,N_19206,N_19550);
and UO_1770 (O_1770,N_19663,N_19750);
or UO_1771 (O_1771,N_19578,N_19454);
xnor UO_1772 (O_1772,N_19742,N_19616);
nor UO_1773 (O_1773,N_19524,N_19779);
or UO_1774 (O_1774,N_19647,N_19896);
nand UO_1775 (O_1775,N_19401,N_19866);
or UO_1776 (O_1776,N_19289,N_19771);
nor UO_1777 (O_1777,N_19997,N_19865);
xor UO_1778 (O_1778,N_19225,N_19525);
xor UO_1779 (O_1779,N_19524,N_19623);
nor UO_1780 (O_1780,N_19441,N_19892);
xor UO_1781 (O_1781,N_19561,N_19764);
nand UO_1782 (O_1782,N_19974,N_19839);
xor UO_1783 (O_1783,N_19635,N_19317);
and UO_1784 (O_1784,N_19654,N_19357);
nor UO_1785 (O_1785,N_19242,N_19301);
and UO_1786 (O_1786,N_19540,N_19896);
nand UO_1787 (O_1787,N_19997,N_19384);
or UO_1788 (O_1788,N_19661,N_19642);
nand UO_1789 (O_1789,N_19549,N_19669);
and UO_1790 (O_1790,N_19809,N_19860);
and UO_1791 (O_1791,N_19469,N_19760);
nor UO_1792 (O_1792,N_19287,N_19590);
nor UO_1793 (O_1793,N_19581,N_19443);
nand UO_1794 (O_1794,N_19432,N_19592);
and UO_1795 (O_1795,N_19987,N_19389);
and UO_1796 (O_1796,N_19603,N_19846);
or UO_1797 (O_1797,N_19612,N_19995);
xnor UO_1798 (O_1798,N_19386,N_19583);
or UO_1799 (O_1799,N_19514,N_19390);
xnor UO_1800 (O_1800,N_19944,N_19637);
or UO_1801 (O_1801,N_19925,N_19870);
nor UO_1802 (O_1802,N_19223,N_19270);
or UO_1803 (O_1803,N_19377,N_19790);
and UO_1804 (O_1804,N_19237,N_19514);
and UO_1805 (O_1805,N_19939,N_19951);
nor UO_1806 (O_1806,N_19808,N_19628);
and UO_1807 (O_1807,N_19489,N_19392);
or UO_1808 (O_1808,N_19557,N_19357);
xor UO_1809 (O_1809,N_19523,N_19423);
nand UO_1810 (O_1810,N_19519,N_19864);
and UO_1811 (O_1811,N_19684,N_19296);
or UO_1812 (O_1812,N_19897,N_19417);
nand UO_1813 (O_1813,N_19604,N_19421);
or UO_1814 (O_1814,N_19333,N_19262);
nor UO_1815 (O_1815,N_19218,N_19443);
nand UO_1816 (O_1816,N_19538,N_19817);
nand UO_1817 (O_1817,N_19727,N_19376);
xnor UO_1818 (O_1818,N_19866,N_19969);
xnor UO_1819 (O_1819,N_19681,N_19490);
nand UO_1820 (O_1820,N_19647,N_19875);
and UO_1821 (O_1821,N_19682,N_19617);
nand UO_1822 (O_1822,N_19590,N_19464);
and UO_1823 (O_1823,N_19499,N_19433);
nand UO_1824 (O_1824,N_19740,N_19263);
and UO_1825 (O_1825,N_19936,N_19809);
nand UO_1826 (O_1826,N_19230,N_19651);
nor UO_1827 (O_1827,N_19927,N_19482);
nor UO_1828 (O_1828,N_19950,N_19476);
nor UO_1829 (O_1829,N_19797,N_19720);
nand UO_1830 (O_1830,N_19725,N_19542);
or UO_1831 (O_1831,N_19433,N_19906);
nor UO_1832 (O_1832,N_19668,N_19767);
nor UO_1833 (O_1833,N_19520,N_19220);
nand UO_1834 (O_1834,N_19417,N_19665);
xor UO_1835 (O_1835,N_19494,N_19578);
or UO_1836 (O_1836,N_19822,N_19696);
nand UO_1837 (O_1837,N_19366,N_19691);
and UO_1838 (O_1838,N_19665,N_19651);
nor UO_1839 (O_1839,N_19366,N_19551);
xor UO_1840 (O_1840,N_19964,N_19637);
or UO_1841 (O_1841,N_19647,N_19439);
or UO_1842 (O_1842,N_19650,N_19216);
and UO_1843 (O_1843,N_19450,N_19579);
nor UO_1844 (O_1844,N_19911,N_19387);
or UO_1845 (O_1845,N_19774,N_19829);
nand UO_1846 (O_1846,N_19478,N_19205);
and UO_1847 (O_1847,N_19500,N_19684);
nand UO_1848 (O_1848,N_19619,N_19777);
xnor UO_1849 (O_1849,N_19667,N_19943);
nor UO_1850 (O_1850,N_19329,N_19699);
xor UO_1851 (O_1851,N_19426,N_19665);
nand UO_1852 (O_1852,N_19384,N_19949);
nor UO_1853 (O_1853,N_19598,N_19783);
or UO_1854 (O_1854,N_19946,N_19208);
xor UO_1855 (O_1855,N_19381,N_19285);
nand UO_1856 (O_1856,N_19215,N_19529);
or UO_1857 (O_1857,N_19513,N_19578);
and UO_1858 (O_1858,N_19886,N_19660);
or UO_1859 (O_1859,N_19273,N_19941);
xnor UO_1860 (O_1860,N_19214,N_19412);
xnor UO_1861 (O_1861,N_19596,N_19723);
or UO_1862 (O_1862,N_19533,N_19604);
or UO_1863 (O_1863,N_19870,N_19310);
nand UO_1864 (O_1864,N_19749,N_19933);
nor UO_1865 (O_1865,N_19909,N_19495);
or UO_1866 (O_1866,N_19235,N_19305);
or UO_1867 (O_1867,N_19717,N_19741);
nand UO_1868 (O_1868,N_19540,N_19521);
nand UO_1869 (O_1869,N_19940,N_19220);
or UO_1870 (O_1870,N_19794,N_19272);
or UO_1871 (O_1871,N_19454,N_19975);
xnor UO_1872 (O_1872,N_19262,N_19235);
nor UO_1873 (O_1873,N_19452,N_19219);
or UO_1874 (O_1874,N_19295,N_19610);
nand UO_1875 (O_1875,N_19316,N_19604);
nor UO_1876 (O_1876,N_19283,N_19965);
or UO_1877 (O_1877,N_19633,N_19344);
nor UO_1878 (O_1878,N_19922,N_19608);
nand UO_1879 (O_1879,N_19356,N_19256);
or UO_1880 (O_1880,N_19864,N_19585);
or UO_1881 (O_1881,N_19792,N_19595);
nor UO_1882 (O_1882,N_19955,N_19507);
nor UO_1883 (O_1883,N_19995,N_19334);
and UO_1884 (O_1884,N_19611,N_19648);
nor UO_1885 (O_1885,N_19599,N_19656);
nand UO_1886 (O_1886,N_19828,N_19416);
and UO_1887 (O_1887,N_19700,N_19531);
nor UO_1888 (O_1888,N_19437,N_19414);
or UO_1889 (O_1889,N_19684,N_19983);
and UO_1890 (O_1890,N_19329,N_19350);
and UO_1891 (O_1891,N_19267,N_19788);
nor UO_1892 (O_1892,N_19724,N_19867);
nor UO_1893 (O_1893,N_19697,N_19583);
xor UO_1894 (O_1894,N_19859,N_19939);
or UO_1895 (O_1895,N_19312,N_19401);
and UO_1896 (O_1896,N_19524,N_19770);
or UO_1897 (O_1897,N_19255,N_19731);
and UO_1898 (O_1898,N_19635,N_19380);
nand UO_1899 (O_1899,N_19741,N_19349);
nor UO_1900 (O_1900,N_19760,N_19960);
or UO_1901 (O_1901,N_19849,N_19299);
and UO_1902 (O_1902,N_19699,N_19624);
nand UO_1903 (O_1903,N_19494,N_19617);
xnor UO_1904 (O_1904,N_19690,N_19563);
or UO_1905 (O_1905,N_19519,N_19856);
and UO_1906 (O_1906,N_19231,N_19272);
or UO_1907 (O_1907,N_19746,N_19308);
and UO_1908 (O_1908,N_19459,N_19517);
xnor UO_1909 (O_1909,N_19332,N_19581);
or UO_1910 (O_1910,N_19576,N_19278);
nand UO_1911 (O_1911,N_19963,N_19765);
nor UO_1912 (O_1912,N_19896,N_19382);
xor UO_1913 (O_1913,N_19611,N_19415);
xor UO_1914 (O_1914,N_19629,N_19313);
nand UO_1915 (O_1915,N_19556,N_19820);
or UO_1916 (O_1916,N_19538,N_19484);
nand UO_1917 (O_1917,N_19391,N_19556);
nor UO_1918 (O_1918,N_19788,N_19980);
xor UO_1919 (O_1919,N_19865,N_19359);
or UO_1920 (O_1920,N_19867,N_19420);
and UO_1921 (O_1921,N_19667,N_19355);
and UO_1922 (O_1922,N_19864,N_19532);
and UO_1923 (O_1923,N_19648,N_19689);
or UO_1924 (O_1924,N_19716,N_19992);
and UO_1925 (O_1925,N_19270,N_19705);
or UO_1926 (O_1926,N_19328,N_19628);
nand UO_1927 (O_1927,N_19944,N_19943);
nor UO_1928 (O_1928,N_19869,N_19419);
and UO_1929 (O_1929,N_19227,N_19983);
xor UO_1930 (O_1930,N_19597,N_19806);
xnor UO_1931 (O_1931,N_19595,N_19699);
or UO_1932 (O_1932,N_19932,N_19616);
or UO_1933 (O_1933,N_19400,N_19845);
and UO_1934 (O_1934,N_19242,N_19656);
xor UO_1935 (O_1935,N_19477,N_19921);
and UO_1936 (O_1936,N_19822,N_19247);
nand UO_1937 (O_1937,N_19471,N_19335);
and UO_1938 (O_1938,N_19640,N_19368);
xnor UO_1939 (O_1939,N_19980,N_19504);
and UO_1940 (O_1940,N_19855,N_19452);
or UO_1941 (O_1941,N_19472,N_19374);
nand UO_1942 (O_1942,N_19923,N_19454);
xor UO_1943 (O_1943,N_19462,N_19788);
nand UO_1944 (O_1944,N_19290,N_19787);
or UO_1945 (O_1945,N_19698,N_19376);
or UO_1946 (O_1946,N_19901,N_19474);
nand UO_1947 (O_1947,N_19940,N_19486);
nor UO_1948 (O_1948,N_19260,N_19504);
xor UO_1949 (O_1949,N_19490,N_19403);
nand UO_1950 (O_1950,N_19345,N_19774);
or UO_1951 (O_1951,N_19895,N_19862);
or UO_1952 (O_1952,N_19928,N_19814);
nand UO_1953 (O_1953,N_19573,N_19447);
nand UO_1954 (O_1954,N_19921,N_19838);
and UO_1955 (O_1955,N_19534,N_19600);
xor UO_1956 (O_1956,N_19527,N_19245);
xor UO_1957 (O_1957,N_19512,N_19714);
or UO_1958 (O_1958,N_19932,N_19820);
nor UO_1959 (O_1959,N_19570,N_19881);
or UO_1960 (O_1960,N_19804,N_19446);
nand UO_1961 (O_1961,N_19439,N_19664);
and UO_1962 (O_1962,N_19519,N_19343);
nand UO_1963 (O_1963,N_19871,N_19528);
nor UO_1964 (O_1964,N_19224,N_19422);
nand UO_1965 (O_1965,N_19825,N_19591);
or UO_1966 (O_1966,N_19616,N_19519);
or UO_1967 (O_1967,N_19730,N_19704);
nand UO_1968 (O_1968,N_19621,N_19993);
nand UO_1969 (O_1969,N_19237,N_19654);
or UO_1970 (O_1970,N_19910,N_19946);
nand UO_1971 (O_1971,N_19675,N_19673);
or UO_1972 (O_1972,N_19890,N_19713);
nand UO_1973 (O_1973,N_19619,N_19865);
and UO_1974 (O_1974,N_19774,N_19513);
nand UO_1975 (O_1975,N_19201,N_19423);
or UO_1976 (O_1976,N_19606,N_19714);
or UO_1977 (O_1977,N_19623,N_19635);
nor UO_1978 (O_1978,N_19322,N_19972);
nand UO_1979 (O_1979,N_19944,N_19605);
nand UO_1980 (O_1980,N_19953,N_19568);
nor UO_1981 (O_1981,N_19635,N_19220);
nor UO_1982 (O_1982,N_19353,N_19229);
xnor UO_1983 (O_1983,N_19919,N_19266);
or UO_1984 (O_1984,N_19364,N_19576);
and UO_1985 (O_1985,N_19389,N_19913);
nand UO_1986 (O_1986,N_19791,N_19444);
and UO_1987 (O_1987,N_19543,N_19727);
nor UO_1988 (O_1988,N_19933,N_19232);
xor UO_1989 (O_1989,N_19301,N_19732);
and UO_1990 (O_1990,N_19851,N_19455);
nor UO_1991 (O_1991,N_19713,N_19416);
nor UO_1992 (O_1992,N_19405,N_19845);
nand UO_1993 (O_1993,N_19982,N_19993);
nand UO_1994 (O_1994,N_19796,N_19290);
nand UO_1995 (O_1995,N_19922,N_19900);
nand UO_1996 (O_1996,N_19237,N_19454);
nor UO_1997 (O_1997,N_19566,N_19311);
xor UO_1998 (O_1998,N_19906,N_19747);
nor UO_1999 (O_1999,N_19751,N_19589);
nor UO_2000 (O_2000,N_19293,N_19798);
nor UO_2001 (O_2001,N_19741,N_19303);
xor UO_2002 (O_2002,N_19219,N_19875);
xor UO_2003 (O_2003,N_19874,N_19562);
or UO_2004 (O_2004,N_19450,N_19767);
nand UO_2005 (O_2005,N_19506,N_19477);
and UO_2006 (O_2006,N_19624,N_19594);
xnor UO_2007 (O_2007,N_19492,N_19560);
xor UO_2008 (O_2008,N_19339,N_19724);
or UO_2009 (O_2009,N_19473,N_19921);
nor UO_2010 (O_2010,N_19490,N_19301);
xor UO_2011 (O_2011,N_19814,N_19716);
xnor UO_2012 (O_2012,N_19511,N_19969);
nand UO_2013 (O_2013,N_19248,N_19646);
nor UO_2014 (O_2014,N_19202,N_19227);
nor UO_2015 (O_2015,N_19661,N_19253);
nand UO_2016 (O_2016,N_19326,N_19636);
and UO_2017 (O_2017,N_19909,N_19499);
xor UO_2018 (O_2018,N_19248,N_19598);
nand UO_2019 (O_2019,N_19791,N_19648);
or UO_2020 (O_2020,N_19386,N_19718);
and UO_2021 (O_2021,N_19621,N_19231);
and UO_2022 (O_2022,N_19855,N_19960);
or UO_2023 (O_2023,N_19470,N_19698);
nand UO_2024 (O_2024,N_19848,N_19800);
and UO_2025 (O_2025,N_19892,N_19920);
or UO_2026 (O_2026,N_19614,N_19826);
nor UO_2027 (O_2027,N_19909,N_19597);
nand UO_2028 (O_2028,N_19869,N_19308);
xor UO_2029 (O_2029,N_19579,N_19305);
or UO_2030 (O_2030,N_19285,N_19786);
nor UO_2031 (O_2031,N_19926,N_19567);
xor UO_2032 (O_2032,N_19371,N_19808);
nand UO_2033 (O_2033,N_19741,N_19801);
xor UO_2034 (O_2034,N_19684,N_19497);
nand UO_2035 (O_2035,N_19286,N_19434);
and UO_2036 (O_2036,N_19239,N_19512);
xnor UO_2037 (O_2037,N_19368,N_19467);
nand UO_2038 (O_2038,N_19611,N_19974);
nor UO_2039 (O_2039,N_19929,N_19879);
nand UO_2040 (O_2040,N_19557,N_19648);
nand UO_2041 (O_2041,N_19398,N_19342);
nand UO_2042 (O_2042,N_19498,N_19751);
nor UO_2043 (O_2043,N_19656,N_19884);
nor UO_2044 (O_2044,N_19499,N_19649);
or UO_2045 (O_2045,N_19266,N_19244);
nor UO_2046 (O_2046,N_19201,N_19407);
nand UO_2047 (O_2047,N_19337,N_19285);
or UO_2048 (O_2048,N_19466,N_19454);
xor UO_2049 (O_2049,N_19762,N_19489);
and UO_2050 (O_2050,N_19412,N_19309);
and UO_2051 (O_2051,N_19733,N_19446);
nor UO_2052 (O_2052,N_19421,N_19996);
xnor UO_2053 (O_2053,N_19632,N_19977);
xnor UO_2054 (O_2054,N_19938,N_19701);
xnor UO_2055 (O_2055,N_19560,N_19640);
nor UO_2056 (O_2056,N_19611,N_19929);
and UO_2057 (O_2057,N_19361,N_19337);
nor UO_2058 (O_2058,N_19637,N_19440);
xnor UO_2059 (O_2059,N_19640,N_19225);
xnor UO_2060 (O_2060,N_19773,N_19829);
and UO_2061 (O_2061,N_19453,N_19833);
or UO_2062 (O_2062,N_19871,N_19881);
and UO_2063 (O_2063,N_19298,N_19872);
and UO_2064 (O_2064,N_19791,N_19279);
and UO_2065 (O_2065,N_19417,N_19721);
xor UO_2066 (O_2066,N_19731,N_19493);
and UO_2067 (O_2067,N_19450,N_19583);
nand UO_2068 (O_2068,N_19724,N_19204);
and UO_2069 (O_2069,N_19392,N_19669);
xor UO_2070 (O_2070,N_19410,N_19927);
or UO_2071 (O_2071,N_19322,N_19220);
nand UO_2072 (O_2072,N_19396,N_19853);
xnor UO_2073 (O_2073,N_19530,N_19644);
or UO_2074 (O_2074,N_19957,N_19646);
nand UO_2075 (O_2075,N_19360,N_19950);
nor UO_2076 (O_2076,N_19959,N_19987);
nand UO_2077 (O_2077,N_19850,N_19260);
nor UO_2078 (O_2078,N_19567,N_19554);
nand UO_2079 (O_2079,N_19672,N_19882);
xnor UO_2080 (O_2080,N_19337,N_19624);
or UO_2081 (O_2081,N_19919,N_19915);
xor UO_2082 (O_2082,N_19697,N_19647);
or UO_2083 (O_2083,N_19999,N_19920);
xor UO_2084 (O_2084,N_19317,N_19264);
and UO_2085 (O_2085,N_19338,N_19208);
and UO_2086 (O_2086,N_19404,N_19333);
or UO_2087 (O_2087,N_19999,N_19740);
nand UO_2088 (O_2088,N_19980,N_19577);
and UO_2089 (O_2089,N_19887,N_19841);
or UO_2090 (O_2090,N_19958,N_19526);
xnor UO_2091 (O_2091,N_19860,N_19222);
and UO_2092 (O_2092,N_19748,N_19888);
or UO_2093 (O_2093,N_19972,N_19489);
or UO_2094 (O_2094,N_19501,N_19667);
or UO_2095 (O_2095,N_19542,N_19251);
nor UO_2096 (O_2096,N_19518,N_19720);
xnor UO_2097 (O_2097,N_19910,N_19380);
xnor UO_2098 (O_2098,N_19352,N_19335);
and UO_2099 (O_2099,N_19456,N_19874);
nor UO_2100 (O_2100,N_19463,N_19768);
nand UO_2101 (O_2101,N_19816,N_19598);
nor UO_2102 (O_2102,N_19475,N_19307);
or UO_2103 (O_2103,N_19309,N_19418);
and UO_2104 (O_2104,N_19382,N_19629);
nor UO_2105 (O_2105,N_19751,N_19601);
nor UO_2106 (O_2106,N_19931,N_19816);
or UO_2107 (O_2107,N_19836,N_19464);
or UO_2108 (O_2108,N_19469,N_19241);
nor UO_2109 (O_2109,N_19579,N_19671);
xor UO_2110 (O_2110,N_19543,N_19628);
nor UO_2111 (O_2111,N_19701,N_19950);
nand UO_2112 (O_2112,N_19710,N_19736);
and UO_2113 (O_2113,N_19752,N_19795);
and UO_2114 (O_2114,N_19359,N_19565);
or UO_2115 (O_2115,N_19938,N_19706);
nand UO_2116 (O_2116,N_19888,N_19971);
xnor UO_2117 (O_2117,N_19970,N_19580);
nor UO_2118 (O_2118,N_19662,N_19519);
xor UO_2119 (O_2119,N_19645,N_19761);
xor UO_2120 (O_2120,N_19897,N_19869);
nor UO_2121 (O_2121,N_19950,N_19263);
nor UO_2122 (O_2122,N_19200,N_19829);
nand UO_2123 (O_2123,N_19452,N_19682);
nand UO_2124 (O_2124,N_19904,N_19614);
nand UO_2125 (O_2125,N_19339,N_19707);
nor UO_2126 (O_2126,N_19457,N_19227);
nand UO_2127 (O_2127,N_19696,N_19724);
nor UO_2128 (O_2128,N_19562,N_19200);
and UO_2129 (O_2129,N_19614,N_19605);
and UO_2130 (O_2130,N_19345,N_19887);
nand UO_2131 (O_2131,N_19240,N_19542);
nor UO_2132 (O_2132,N_19202,N_19368);
or UO_2133 (O_2133,N_19967,N_19202);
and UO_2134 (O_2134,N_19829,N_19270);
or UO_2135 (O_2135,N_19969,N_19661);
nand UO_2136 (O_2136,N_19795,N_19586);
and UO_2137 (O_2137,N_19670,N_19958);
nor UO_2138 (O_2138,N_19876,N_19353);
xnor UO_2139 (O_2139,N_19641,N_19790);
or UO_2140 (O_2140,N_19828,N_19533);
nand UO_2141 (O_2141,N_19718,N_19442);
and UO_2142 (O_2142,N_19739,N_19207);
or UO_2143 (O_2143,N_19923,N_19794);
nor UO_2144 (O_2144,N_19246,N_19236);
nand UO_2145 (O_2145,N_19793,N_19290);
nand UO_2146 (O_2146,N_19556,N_19368);
nand UO_2147 (O_2147,N_19543,N_19401);
nand UO_2148 (O_2148,N_19814,N_19498);
xor UO_2149 (O_2149,N_19679,N_19427);
or UO_2150 (O_2150,N_19906,N_19472);
nand UO_2151 (O_2151,N_19489,N_19786);
or UO_2152 (O_2152,N_19424,N_19987);
or UO_2153 (O_2153,N_19758,N_19630);
nor UO_2154 (O_2154,N_19887,N_19535);
and UO_2155 (O_2155,N_19812,N_19965);
nand UO_2156 (O_2156,N_19662,N_19638);
and UO_2157 (O_2157,N_19405,N_19858);
nand UO_2158 (O_2158,N_19711,N_19296);
nor UO_2159 (O_2159,N_19768,N_19305);
or UO_2160 (O_2160,N_19899,N_19836);
and UO_2161 (O_2161,N_19478,N_19879);
nand UO_2162 (O_2162,N_19915,N_19882);
or UO_2163 (O_2163,N_19335,N_19887);
nand UO_2164 (O_2164,N_19545,N_19447);
xnor UO_2165 (O_2165,N_19333,N_19870);
and UO_2166 (O_2166,N_19530,N_19710);
or UO_2167 (O_2167,N_19430,N_19476);
and UO_2168 (O_2168,N_19551,N_19613);
nand UO_2169 (O_2169,N_19500,N_19486);
and UO_2170 (O_2170,N_19373,N_19681);
xor UO_2171 (O_2171,N_19368,N_19522);
or UO_2172 (O_2172,N_19733,N_19916);
nand UO_2173 (O_2173,N_19371,N_19881);
xor UO_2174 (O_2174,N_19769,N_19556);
and UO_2175 (O_2175,N_19894,N_19507);
xnor UO_2176 (O_2176,N_19501,N_19511);
xnor UO_2177 (O_2177,N_19362,N_19297);
or UO_2178 (O_2178,N_19804,N_19738);
nand UO_2179 (O_2179,N_19410,N_19645);
nor UO_2180 (O_2180,N_19258,N_19368);
or UO_2181 (O_2181,N_19285,N_19375);
and UO_2182 (O_2182,N_19658,N_19204);
nand UO_2183 (O_2183,N_19764,N_19205);
xor UO_2184 (O_2184,N_19719,N_19860);
xor UO_2185 (O_2185,N_19308,N_19443);
xnor UO_2186 (O_2186,N_19471,N_19886);
xor UO_2187 (O_2187,N_19309,N_19221);
or UO_2188 (O_2188,N_19281,N_19815);
xor UO_2189 (O_2189,N_19548,N_19803);
nor UO_2190 (O_2190,N_19329,N_19603);
or UO_2191 (O_2191,N_19693,N_19917);
and UO_2192 (O_2192,N_19811,N_19808);
nand UO_2193 (O_2193,N_19524,N_19391);
or UO_2194 (O_2194,N_19848,N_19473);
and UO_2195 (O_2195,N_19809,N_19485);
nor UO_2196 (O_2196,N_19262,N_19652);
or UO_2197 (O_2197,N_19255,N_19888);
and UO_2198 (O_2198,N_19802,N_19921);
nor UO_2199 (O_2199,N_19322,N_19926);
and UO_2200 (O_2200,N_19998,N_19252);
nand UO_2201 (O_2201,N_19561,N_19547);
nor UO_2202 (O_2202,N_19552,N_19428);
xnor UO_2203 (O_2203,N_19544,N_19268);
nand UO_2204 (O_2204,N_19230,N_19267);
and UO_2205 (O_2205,N_19603,N_19746);
nor UO_2206 (O_2206,N_19821,N_19595);
xnor UO_2207 (O_2207,N_19599,N_19861);
and UO_2208 (O_2208,N_19212,N_19312);
xnor UO_2209 (O_2209,N_19858,N_19431);
and UO_2210 (O_2210,N_19370,N_19602);
nand UO_2211 (O_2211,N_19562,N_19503);
nand UO_2212 (O_2212,N_19766,N_19537);
nor UO_2213 (O_2213,N_19911,N_19834);
nand UO_2214 (O_2214,N_19453,N_19982);
nor UO_2215 (O_2215,N_19868,N_19918);
nor UO_2216 (O_2216,N_19806,N_19536);
or UO_2217 (O_2217,N_19416,N_19915);
nand UO_2218 (O_2218,N_19331,N_19946);
and UO_2219 (O_2219,N_19218,N_19722);
nor UO_2220 (O_2220,N_19680,N_19890);
or UO_2221 (O_2221,N_19617,N_19392);
nor UO_2222 (O_2222,N_19634,N_19245);
and UO_2223 (O_2223,N_19458,N_19577);
nand UO_2224 (O_2224,N_19215,N_19203);
nor UO_2225 (O_2225,N_19901,N_19744);
nand UO_2226 (O_2226,N_19228,N_19492);
xor UO_2227 (O_2227,N_19745,N_19963);
or UO_2228 (O_2228,N_19673,N_19374);
nand UO_2229 (O_2229,N_19510,N_19696);
or UO_2230 (O_2230,N_19364,N_19727);
xor UO_2231 (O_2231,N_19303,N_19876);
nor UO_2232 (O_2232,N_19457,N_19506);
nand UO_2233 (O_2233,N_19696,N_19434);
nand UO_2234 (O_2234,N_19382,N_19409);
nor UO_2235 (O_2235,N_19698,N_19626);
nand UO_2236 (O_2236,N_19637,N_19914);
nand UO_2237 (O_2237,N_19820,N_19422);
nor UO_2238 (O_2238,N_19443,N_19522);
xor UO_2239 (O_2239,N_19906,N_19903);
or UO_2240 (O_2240,N_19614,N_19310);
or UO_2241 (O_2241,N_19388,N_19929);
and UO_2242 (O_2242,N_19252,N_19513);
xnor UO_2243 (O_2243,N_19702,N_19834);
xor UO_2244 (O_2244,N_19383,N_19680);
xor UO_2245 (O_2245,N_19887,N_19799);
and UO_2246 (O_2246,N_19270,N_19484);
nand UO_2247 (O_2247,N_19371,N_19406);
nand UO_2248 (O_2248,N_19742,N_19970);
nor UO_2249 (O_2249,N_19597,N_19300);
nand UO_2250 (O_2250,N_19961,N_19858);
or UO_2251 (O_2251,N_19841,N_19550);
and UO_2252 (O_2252,N_19633,N_19951);
xnor UO_2253 (O_2253,N_19803,N_19439);
or UO_2254 (O_2254,N_19527,N_19619);
nor UO_2255 (O_2255,N_19229,N_19744);
xor UO_2256 (O_2256,N_19553,N_19600);
nand UO_2257 (O_2257,N_19894,N_19791);
and UO_2258 (O_2258,N_19972,N_19530);
xnor UO_2259 (O_2259,N_19764,N_19209);
and UO_2260 (O_2260,N_19347,N_19345);
nor UO_2261 (O_2261,N_19454,N_19919);
xor UO_2262 (O_2262,N_19237,N_19644);
or UO_2263 (O_2263,N_19477,N_19791);
nor UO_2264 (O_2264,N_19497,N_19819);
nand UO_2265 (O_2265,N_19205,N_19876);
nand UO_2266 (O_2266,N_19953,N_19562);
xnor UO_2267 (O_2267,N_19881,N_19663);
or UO_2268 (O_2268,N_19259,N_19356);
nor UO_2269 (O_2269,N_19443,N_19878);
nor UO_2270 (O_2270,N_19783,N_19908);
nand UO_2271 (O_2271,N_19303,N_19547);
and UO_2272 (O_2272,N_19789,N_19417);
xnor UO_2273 (O_2273,N_19244,N_19984);
and UO_2274 (O_2274,N_19321,N_19298);
or UO_2275 (O_2275,N_19821,N_19707);
nand UO_2276 (O_2276,N_19963,N_19308);
or UO_2277 (O_2277,N_19662,N_19221);
or UO_2278 (O_2278,N_19812,N_19333);
and UO_2279 (O_2279,N_19404,N_19993);
nand UO_2280 (O_2280,N_19965,N_19930);
or UO_2281 (O_2281,N_19629,N_19520);
nand UO_2282 (O_2282,N_19362,N_19335);
nor UO_2283 (O_2283,N_19946,N_19769);
or UO_2284 (O_2284,N_19573,N_19606);
and UO_2285 (O_2285,N_19202,N_19312);
xnor UO_2286 (O_2286,N_19562,N_19642);
or UO_2287 (O_2287,N_19386,N_19947);
nor UO_2288 (O_2288,N_19576,N_19714);
nor UO_2289 (O_2289,N_19780,N_19492);
nor UO_2290 (O_2290,N_19667,N_19702);
xnor UO_2291 (O_2291,N_19579,N_19709);
and UO_2292 (O_2292,N_19734,N_19360);
xnor UO_2293 (O_2293,N_19540,N_19650);
xnor UO_2294 (O_2294,N_19577,N_19388);
or UO_2295 (O_2295,N_19296,N_19419);
and UO_2296 (O_2296,N_19346,N_19848);
xor UO_2297 (O_2297,N_19860,N_19241);
xor UO_2298 (O_2298,N_19927,N_19576);
xor UO_2299 (O_2299,N_19640,N_19782);
and UO_2300 (O_2300,N_19547,N_19436);
xnor UO_2301 (O_2301,N_19654,N_19983);
xnor UO_2302 (O_2302,N_19536,N_19878);
xor UO_2303 (O_2303,N_19501,N_19368);
nand UO_2304 (O_2304,N_19228,N_19764);
or UO_2305 (O_2305,N_19249,N_19948);
or UO_2306 (O_2306,N_19250,N_19978);
or UO_2307 (O_2307,N_19859,N_19245);
xor UO_2308 (O_2308,N_19931,N_19634);
or UO_2309 (O_2309,N_19729,N_19323);
and UO_2310 (O_2310,N_19624,N_19672);
or UO_2311 (O_2311,N_19351,N_19355);
nor UO_2312 (O_2312,N_19288,N_19443);
nand UO_2313 (O_2313,N_19558,N_19743);
nand UO_2314 (O_2314,N_19867,N_19399);
nand UO_2315 (O_2315,N_19868,N_19433);
nor UO_2316 (O_2316,N_19603,N_19617);
nand UO_2317 (O_2317,N_19621,N_19399);
or UO_2318 (O_2318,N_19639,N_19875);
nand UO_2319 (O_2319,N_19359,N_19897);
and UO_2320 (O_2320,N_19208,N_19949);
or UO_2321 (O_2321,N_19924,N_19928);
xnor UO_2322 (O_2322,N_19645,N_19205);
or UO_2323 (O_2323,N_19475,N_19444);
xnor UO_2324 (O_2324,N_19362,N_19957);
and UO_2325 (O_2325,N_19296,N_19612);
or UO_2326 (O_2326,N_19890,N_19434);
xnor UO_2327 (O_2327,N_19449,N_19778);
and UO_2328 (O_2328,N_19513,N_19203);
nand UO_2329 (O_2329,N_19760,N_19797);
nor UO_2330 (O_2330,N_19525,N_19434);
or UO_2331 (O_2331,N_19384,N_19239);
xor UO_2332 (O_2332,N_19524,N_19826);
and UO_2333 (O_2333,N_19764,N_19667);
nor UO_2334 (O_2334,N_19369,N_19249);
and UO_2335 (O_2335,N_19438,N_19397);
nand UO_2336 (O_2336,N_19684,N_19858);
or UO_2337 (O_2337,N_19272,N_19698);
and UO_2338 (O_2338,N_19368,N_19886);
nand UO_2339 (O_2339,N_19975,N_19400);
xnor UO_2340 (O_2340,N_19213,N_19323);
nand UO_2341 (O_2341,N_19834,N_19743);
and UO_2342 (O_2342,N_19472,N_19599);
or UO_2343 (O_2343,N_19371,N_19689);
or UO_2344 (O_2344,N_19684,N_19391);
or UO_2345 (O_2345,N_19519,N_19349);
or UO_2346 (O_2346,N_19293,N_19760);
xnor UO_2347 (O_2347,N_19840,N_19431);
and UO_2348 (O_2348,N_19851,N_19572);
xor UO_2349 (O_2349,N_19704,N_19507);
xnor UO_2350 (O_2350,N_19727,N_19666);
and UO_2351 (O_2351,N_19669,N_19672);
nand UO_2352 (O_2352,N_19280,N_19284);
nor UO_2353 (O_2353,N_19577,N_19297);
xnor UO_2354 (O_2354,N_19738,N_19856);
xnor UO_2355 (O_2355,N_19309,N_19289);
and UO_2356 (O_2356,N_19622,N_19285);
xor UO_2357 (O_2357,N_19888,N_19229);
and UO_2358 (O_2358,N_19468,N_19599);
and UO_2359 (O_2359,N_19636,N_19797);
xor UO_2360 (O_2360,N_19207,N_19606);
and UO_2361 (O_2361,N_19804,N_19562);
and UO_2362 (O_2362,N_19470,N_19286);
and UO_2363 (O_2363,N_19592,N_19735);
and UO_2364 (O_2364,N_19458,N_19661);
and UO_2365 (O_2365,N_19961,N_19296);
xnor UO_2366 (O_2366,N_19621,N_19344);
or UO_2367 (O_2367,N_19756,N_19503);
nor UO_2368 (O_2368,N_19917,N_19459);
nand UO_2369 (O_2369,N_19435,N_19653);
nor UO_2370 (O_2370,N_19324,N_19385);
nor UO_2371 (O_2371,N_19671,N_19894);
nand UO_2372 (O_2372,N_19858,N_19519);
nor UO_2373 (O_2373,N_19618,N_19926);
and UO_2374 (O_2374,N_19427,N_19353);
nor UO_2375 (O_2375,N_19687,N_19995);
and UO_2376 (O_2376,N_19276,N_19244);
nand UO_2377 (O_2377,N_19561,N_19217);
nand UO_2378 (O_2378,N_19728,N_19968);
nor UO_2379 (O_2379,N_19844,N_19307);
nand UO_2380 (O_2380,N_19932,N_19857);
nor UO_2381 (O_2381,N_19418,N_19584);
xnor UO_2382 (O_2382,N_19790,N_19438);
and UO_2383 (O_2383,N_19660,N_19524);
or UO_2384 (O_2384,N_19432,N_19847);
or UO_2385 (O_2385,N_19439,N_19683);
nor UO_2386 (O_2386,N_19721,N_19270);
xnor UO_2387 (O_2387,N_19611,N_19856);
nor UO_2388 (O_2388,N_19618,N_19772);
nor UO_2389 (O_2389,N_19850,N_19675);
and UO_2390 (O_2390,N_19723,N_19996);
and UO_2391 (O_2391,N_19814,N_19211);
nand UO_2392 (O_2392,N_19669,N_19905);
or UO_2393 (O_2393,N_19782,N_19219);
xnor UO_2394 (O_2394,N_19446,N_19300);
and UO_2395 (O_2395,N_19774,N_19882);
and UO_2396 (O_2396,N_19326,N_19387);
or UO_2397 (O_2397,N_19519,N_19439);
xor UO_2398 (O_2398,N_19754,N_19297);
nand UO_2399 (O_2399,N_19471,N_19912);
and UO_2400 (O_2400,N_19839,N_19278);
nor UO_2401 (O_2401,N_19272,N_19507);
xor UO_2402 (O_2402,N_19436,N_19560);
nor UO_2403 (O_2403,N_19895,N_19606);
or UO_2404 (O_2404,N_19730,N_19861);
xnor UO_2405 (O_2405,N_19748,N_19565);
xor UO_2406 (O_2406,N_19470,N_19229);
xor UO_2407 (O_2407,N_19317,N_19852);
or UO_2408 (O_2408,N_19730,N_19298);
nand UO_2409 (O_2409,N_19962,N_19892);
and UO_2410 (O_2410,N_19781,N_19234);
and UO_2411 (O_2411,N_19473,N_19242);
nand UO_2412 (O_2412,N_19604,N_19953);
xnor UO_2413 (O_2413,N_19443,N_19805);
xor UO_2414 (O_2414,N_19519,N_19632);
xor UO_2415 (O_2415,N_19394,N_19870);
nor UO_2416 (O_2416,N_19668,N_19644);
and UO_2417 (O_2417,N_19876,N_19609);
and UO_2418 (O_2418,N_19973,N_19781);
or UO_2419 (O_2419,N_19933,N_19981);
and UO_2420 (O_2420,N_19206,N_19267);
or UO_2421 (O_2421,N_19578,N_19366);
nor UO_2422 (O_2422,N_19747,N_19517);
and UO_2423 (O_2423,N_19242,N_19444);
nand UO_2424 (O_2424,N_19912,N_19217);
or UO_2425 (O_2425,N_19766,N_19667);
or UO_2426 (O_2426,N_19880,N_19931);
nor UO_2427 (O_2427,N_19953,N_19795);
or UO_2428 (O_2428,N_19693,N_19655);
nor UO_2429 (O_2429,N_19254,N_19370);
xor UO_2430 (O_2430,N_19880,N_19481);
and UO_2431 (O_2431,N_19655,N_19543);
xnor UO_2432 (O_2432,N_19775,N_19915);
xor UO_2433 (O_2433,N_19664,N_19239);
xor UO_2434 (O_2434,N_19422,N_19557);
or UO_2435 (O_2435,N_19505,N_19437);
and UO_2436 (O_2436,N_19453,N_19317);
nor UO_2437 (O_2437,N_19648,N_19543);
xor UO_2438 (O_2438,N_19958,N_19748);
xor UO_2439 (O_2439,N_19204,N_19441);
xnor UO_2440 (O_2440,N_19356,N_19930);
and UO_2441 (O_2441,N_19782,N_19906);
nand UO_2442 (O_2442,N_19896,N_19632);
or UO_2443 (O_2443,N_19854,N_19867);
and UO_2444 (O_2444,N_19364,N_19631);
xnor UO_2445 (O_2445,N_19515,N_19526);
xnor UO_2446 (O_2446,N_19464,N_19334);
and UO_2447 (O_2447,N_19760,N_19668);
nor UO_2448 (O_2448,N_19901,N_19792);
xor UO_2449 (O_2449,N_19279,N_19851);
nand UO_2450 (O_2450,N_19962,N_19425);
and UO_2451 (O_2451,N_19839,N_19760);
or UO_2452 (O_2452,N_19954,N_19555);
xnor UO_2453 (O_2453,N_19475,N_19580);
xnor UO_2454 (O_2454,N_19961,N_19795);
xor UO_2455 (O_2455,N_19776,N_19224);
and UO_2456 (O_2456,N_19870,N_19966);
and UO_2457 (O_2457,N_19421,N_19874);
nor UO_2458 (O_2458,N_19788,N_19400);
or UO_2459 (O_2459,N_19379,N_19744);
and UO_2460 (O_2460,N_19832,N_19318);
and UO_2461 (O_2461,N_19386,N_19326);
or UO_2462 (O_2462,N_19553,N_19202);
or UO_2463 (O_2463,N_19263,N_19468);
nand UO_2464 (O_2464,N_19950,N_19739);
xor UO_2465 (O_2465,N_19629,N_19356);
nor UO_2466 (O_2466,N_19394,N_19596);
nand UO_2467 (O_2467,N_19619,N_19456);
or UO_2468 (O_2468,N_19556,N_19746);
nand UO_2469 (O_2469,N_19556,N_19380);
and UO_2470 (O_2470,N_19796,N_19380);
nor UO_2471 (O_2471,N_19292,N_19800);
xnor UO_2472 (O_2472,N_19775,N_19360);
nor UO_2473 (O_2473,N_19896,N_19640);
and UO_2474 (O_2474,N_19754,N_19953);
nand UO_2475 (O_2475,N_19547,N_19664);
or UO_2476 (O_2476,N_19805,N_19976);
nand UO_2477 (O_2477,N_19670,N_19271);
and UO_2478 (O_2478,N_19772,N_19371);
xor UO_2479 (O_2479,N_19526,N_19674);
or UO_2480 (O_2480,N_19715,N_19393);
nand UO_2481 (O_2481,N_19607,N_19512);
and UO_2482 (O_2482,N_19299,N_19220);
nor UO_2483 (O_2483,N_19667,N_19512);
nor UO_2484 (O_2484,N_19479,N_19857);
nor UO_2485 (O_2485,N_19682,N_19881);
nand UO_2486 (O_2486,N_19947,N_19326);
xnor UO_2487 (O_2487,N_19697,N_19855);
xor UO_2488 (O_2488,N_19835,N_19354);
nand UO_2489 (O_2489,N_19275,N_19540);
xor UO_2490 (O_2490,N_19230,N_19806);
nand UO_2491 (O_2491,N_19703,N_19848);
nand UO_2492 (O_2492,N_19766,N_19566);
xor UO_2493 (O_2493,N_19927,N_19827);
xnor UO_2494 (O_2494,N_19646,N_19722);
xor UO_2495 (O_2495,N_19826,N_19809);
xnor UO_2496 (O_2496,N_19564,N_19264);
xnor UO_2497 (O_2497,N_19710,N_19566);
nor UO_2498 (O_2498,N_19206,N_19256);
or UO_2499 (O_2499,N_19917,N_19414);
endmodule