module basic_1500_15000_2000_3_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10002,N_10003,N_10004,N_10005,N_10007,N_10008,N_10009,N_10010,N_10011,N_10014,N_10015,N_10016,N_10018,N_10019,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10048,N_10050,N_10051,N_10052,N_10053,N_10054,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10068,N_10069,N_10070,N_10071,N_10072,N_10075,N_10076,N_10077,N_10078,N_10080,N_10082,N_10084,N_10085,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10100,N_10101,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10118,N_10119,N_10121,N_10122,N_10123,N_10125,N_10126,N_10128,N_10129,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10145,N_10146,N_10147,N_10148,N_10150,N_10151,N_10154,N_10155,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10179,N_10181,N_10182,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10194,N_10195,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10235,N_10236,N_10240,N_10242,N_10243,N_10244,N_10245,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10257,N_10258,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10305,N_10307,N_10308,N_10309,N_10310,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10323,N_10324,N_10325,N_10326,N_10327,N_10330,N_10331,N_10333,N_10334,N_10335,N_10336,N_10338,N_10339,N_10340,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10358,N_10359,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10370,N_10371,N_10373,N_10374,N_10375,N_10377,N_10379,N_10382,N_10383,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10399,N_10400,N_10401,N_10402,N_10403,N_10405,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10425,N_10427,N_10428,N_10429,N_10430,N_10431,N_10433,N_10434,N_10436,N_10437,N_10438,N_10439,N_10441,N_10442,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10454,N_10456,N_10457,N_10458,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10474,N_10475,N_10476,N_10477,N_10478,N_10480,N_10481,N_10482,N_10485,N_10486,N_10487,N_10491,N_10493,N_10494,N_10495,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10517,N_10519,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10529,N_10531,N_10532,N_10533,N_10534,N_10535,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10547,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10558,N_10561,N_10562,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10611,N_10613,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10622,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10675,N_10677,N_10678,N_10680,N_10681,N_10682,N_10683,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10709,N_10710,N_10711,N_10712,N_10714,N_10715,N_10717,N_10718,N_10721,N_10722,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10757,N_10758,N_10762,N_10763,N_10765,N_10766,N_10767,N_10768,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10796,N_10798,N_10799,N_10800,N_10802,N_10803,N_10804,N_10805,N_10806,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10820,N_10821,N_10822,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10831,N_10832,N_10833,N_10834,N_10836,N_10838,N_10839,N_10840,N_10841,N_10843,N_10845,N_10846,N_10847,N_10848,N_10849,N_10851,N_10852,N_10854,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10875,N_10878,N_10879,N_10881,N_10882,N_10884,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10897,N_10898,N_10899,N_10900,N_10901,N_10904,N_10905,N_10906,N_10907,N_10909,N_10910,N_10911,N_10912,N_10914,N_10918,N_10919,N_10920,N_10921,N_10922,N_10925,N_10926,N_10927,N_10928,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10937,N_10939,N_10940,N_10941,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10966,N_10967,N_10969,N_10970,N_10974,N_10976,N_10978,N_10979,N_10980,N_10981,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10995,N_10996,N_10997,N_10998,N_11000,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11047,N_11048,N_11049,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11065,N_11066,N_11067,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11096,N_11097,N_11098,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11114,N_11115,N_11116,N_11117,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11130,N_11133,N_11135,N_11136,N_11137,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11146,N_11148,N_11149,N_11150,N_11151,N_11153,N_11154,N_11156,N_11157,N_11159,N_11160,N_11161,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11196,N_11197,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11209,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11227,N_11228,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11245,N_11247,N_11249,N_11250,N_11251,N_11252,N_11253,N_11255,N_11256,N_11258,N_11259,N_11260,N_11262,N_11263,N_11264,N_11266,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11288,N_11289,N_11290,N_11292,N_11293,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11304,N_11305,N_11306,N_11307,N_11308,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11335,N_11336,N_11338,N_11339,N_11341,N_11342,N_11345,N_11346,N_11347,N_11348,N_11350,N_11351,N_11352,N_11355,N_11356,N_11357,N_11359,N_11360,N_11361,N_11363,N_11364,N_11365,N_11367,N_11368,N_11369,N_11371,N_11373,N_11374,N_11375,N_11378,N_11379,N_11380,N_11381,N_11382,N_11384,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11406,N_11407,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11436,N_11438,N_11441,N_11442,N_11443,N_11445,N_11446,N_11447,N_11450,N_11452,N_11454,N_11455,N_11457,N_11458,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11501,N_11502,N_11503,N_11504,N_11507,N_11509,N_11510,N_11511,N_11512,N_11513,N_11515,N_11516,N_11517,N_11518,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11529,N_11530,N_11531,N_11532,N_11534,N_11535,N_11536,N_11537,N_11538,N_11541,N_11542,N_11544,N_11545,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11555,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11580,N_11582,N_11583,N_11584,N_11586,N_11588,N_11589,N_11590,N_11592,N_11593,N_11594,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11613,N_11615,N_11616,N_11617,N_11618,N_11619,N_11621,N_11622,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11643,N_11644,N_11645,N_11647,N_11649,N_11650,N_11651,N_11652,N_11654,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11665,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11688,N_11689,N_11691,N_11693,N_11694,N_11695,N_11696,N_11697,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11716,N_11717,N_11719,N_11721,N_11723,N_11724,N_11725,N_11726,N_11727,N_11729,N_11730,N_11731,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11748,N_11749,N_11750,N_11751,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11767,N_11768,N_11769,N_11770,N_11772,N_11773,N_11774,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11799,N_11801,N_11802,N_11803,N_11804,N_11805,N_11807,N_11809,N_11810,N_11811,N_11812,N_11813,N_11817,N_11818,N_11820,N_11821,N_11822,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11835,N_11836,N_11837,N_11839,N_11840,N_11841,N_11845,N_11846,N_11848,N_11849,N_11850,N_11851,N_11852,N_11854,N_11855,N_11858,N_11859,N_11860,N_11862,N_11863,N_11864,N_11865,N_11866,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11875,N_11876,N_11877,N_11880,N_11881,N_11886,N_11887,N_11889,N_11891,N_11892,N_11895,N_11896,N_11897,N_11898,N_11899,N_11901,N_11902,N_11903,N_11904,N_11906,N_11908,N_11909,N_11912,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11922,N_11923,N_11924,N_11926,N_11927,N_11929,N_11932,N_11933,N_11935,N_11936,N_11937,N_11940,N_11941,N_11943,N_11944,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11981,N_11982,N_11983,N_11984,N_11986,N_11987,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12017,N_12018,N_12020,N_12021,N_12022,N_12024,N_12025,N_12026,N_12027,N_12031,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12063,N_12064,N_12067,N_12069,N_12070,N_12071,N_12072,N_12074,N_12075,N_12076,N_12077,N_12079,N_12080,N_12081,N_12082,N_12083,N_12085,N_12086,N_12087,N_12089,N_12090,N_12091,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12107,N_12109,N_12110,N_12112,N_12113,N_12114,N_12116,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12127,N_12128,N_12130,N_12132,N_12133,N_12134,N_12135,N_12137,N_12138,N_12139,N_12141,N_12142,N_12143,N_12144,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12193,N_12194,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12210,N_12211,N_12212,N_12214,N_12215,N_12216,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12236,N_12237,N_12238,N_12239,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12254,N_12255,N_12256,N_12257,N_12259,N_12260,N_12261,N_12263,N_12265,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12281,N_12282,N_12283,N_12286,N_12288,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12297,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12319,N_12321,N_12322,N_12323,N_12324,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12336,N_12337,N_12338,N_12339,N_12342,N_12343,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12368,N_12369,N_12370,N_12372,N_12373,N_12374,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12407,N_12411,N_12413,N_12414,N_12416,N_12417,N_12418,N_12419,N_12421,N_12422,N_12424,N_12425,N_12427,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12444,N_12445,N_12448,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12458,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12469,N_12470,N_12472,N_12473,N_12474,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12485,N_12486,N_12487,N_12488,N_12491,N_12493,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12520,N_12521,N_12522,N_12523,N_12524,N_12528,N_12531,N_12532,N_12534,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12561,N_12563,N_12564,N_12565,N_12566,N_12567,N_12570,N_12572,N_12573,N_12574,N_12575,N_12577,N_12578,N_12579,N_12580,N_12583,N_12584,N_12585,N_12586,N_12587,N_12589,N_12590,N_12592,N_12593,N_12595,N_12596,N_12598,N_12599,N_12601,N_12603,N_12604,N_12605,N_12608,N_12609,N_12610,N_12613,N_12614,N_12615,N_12616,N_12617,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12641,N_12642,N_12643,N_12645,N_12647,N_12648,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12661,N_12662,N_12664,N_12665,N_12666,N_12667,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12679,N_12680,N_12681,N_12682,N_12683,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12696,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12723,N_12725,N_12726,N_12727,N_12729,N_12730,N_12731,N_12732,N_12733,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12750,N_12751,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12773,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12799,N_12800,N_12801,N_12802,N_12804,N_12805,N_12806,N_12807,N_12809,N_12810,N_12811,N_12812,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12822,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12835,N_12836,N_12838,N_12840,N_12841,N_12842,N_12843,N_12844,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12864,N_12865,N_12866,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12878,N_12879,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12896,N_12897,N_12901,N_12902,N_12904,N_12905,N_12906,N_12907,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12928,N_12929,N_12930,N_12933,N_12934,N_12935,N_12936,N_12938,N_12939,N_12941,N_12943,N_12944,N_12945,N_12947,N_12949,N_12950,N_12951,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12983,N_12984,N_12985,N_12988,N_12989,N_12990,N_12991,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13007,N_13008,N_13011,N_13012,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13023,N_13024,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13033,N_13034,N_13035,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13046,N_13048,N_13049,N_13052,N_13054,N_13055,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13065,N_13066,N_13067,N_13068,N_13070,N_13073,N_13075,N_13078,N_13079,N_13080,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13089,N_13090,N_13091,N_13092,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13108,N_13109,N_13110,N_13111,N_13113,N_13115,N_13117,N_13119,N_13120,N_13121,N_13122,N_13123,N_13125,N_13126,N_13127,N_13129,N_13131,N_13133,N_13135,N_13136,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13146,N_13147,N_13148,N_13150,N_13151,N_13152,N_13154,N_13155,N_13157,N_13158,N_13159,N_13160,N_13162,N_13163,N_13165,N_13166,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13218,N_13219,N_13220,N_13221,N_13223,N_13224,N_13225,N_13226,N_13228,N_13229,N_13230,N_13231,N_13232,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13242,N_13244,N_13245,N_13246,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13281,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13293,N_13294,N_13295,N_13297,N_13298,N_13300,N_13302,N_13303,N_13304,N_13306,N_13307,N_13308,N_13309,N_13310,N_13312,N_13313,N_13314,N_13315,N_13316,N_13319,N_13320,N_13322,N_13325,N_13327,N_13328,N_13329,N_13331,N_13332,N_13333,N_13334,N_13337,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13349,N_13350,N_13351,N_13352,N_13355,N_13356,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13383,N_13384,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13417,N_13418,N_13419,N_13420,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13430,N_13433,N_13434,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13485,N_13486,N_13487,N_13488,N_13489,N_13491,N_13492,N_13493,N_13495,N_13497,N_13498,N_13499,N_13500,N_13503,N_13504,N_13505,N_13506,N_13507,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13534,N_13535,N_13536,N_13537,N_13538,N_13540,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13549,N_13550,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13584,N_13585,N_13586,N_13587,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13618,N_13619,N_13620,N_13621,N_13623,N_13624,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13650,N_13651,N_13652,N_13655,N_13656,N_13657,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13675,N_13676,N_13677,N_13679,N_13680,N_13681,N_13682,N_13684,N_13686,N_13687,N_13688,N_13689,N_13690,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13702,N_13704,N_13705,N_13708,N_13709,N_13710,N_13711,N_13712,N_13714,N_13716,N_13717,N_13718,N_13720,N_13721,N_13722,N_13723,N_13724,N_13726,N_13728,N_13730,N_13731,N_13733,N_13735,N_13736,N_13737,N_13739,N_13740,N_13742,N_13743,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13755,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13807,N_13808,N_13809,N_13811,N_13812,N_13813,N_13814,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13839,N_13840,N_13842,N_13843,N_13844,N_13846,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13858,N_13859,N_13860,N_13862,N_13863,N_13864,N_13865,N_13866,N_13868,N_13869,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13878,N_13879,N_13880,N_13881,N_13883,N_13884,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13904,N_13907,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13919,N_13920,N_13921,N_13922,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13940,N_13941,N_13942,N_13943,N_13945,N_13946,N_13947,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13962,N_13963,N_13964,N_13965,N_13966,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13979,N_13980,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13996,N_13998,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14021,N_14023,N_14024,N_14025,N_14026,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14055,N_14056,N_14057,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14068,N_14069,N_14070,N_14071,N_14072,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14081,N_14082,N_14084,N_14085,N_14086,N_14087,N_14089,N_14090,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14100,N_14101,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14113,N_14115,N_14116,N_14117,N_14120,N_14122,N_14124,N_14125,N_14126,N_14127,N_14129,N_14130,N_14131,N_14133,N_14134,N_14135,N_14137,N_14138,N_14139,N_14140,N_14143,N_14144,N_14146,N_14147,N_14148,N_14150,N_14152,N_14153,N_14154,N_14156,N_14157,N_14158,N_14159,N_14162,N_14163,N_14165,N_14166,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14186,N_14187,N_14188,N_14189,N_14191,N_14193,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14237,N_14238,N_14239,N_14240,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14251,N_14252,N_14253,N_14254,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14265,N_14266,N_14267,N_14268,N_14271,N_14272,N_14273,N_14275,N_14277,N_14278,N_14279,N_14280,N_14281,N_14283,N_14284,N_14285,N_14287,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14300,N_14301,N_14303,N_14304,N_14305,N_14306,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14349,N_14350,N_14351,N_14353,N_14355,N_14356,N_14358,N_14359,N_14360,N_14361,N_14362,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14374,N_14375,N_14376,N_14377,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14409,N_14411,N_14414,N_14415,N_14416,N_14417,N_14419,N_14420,N_14422,N_14428,N_14429,N_14432,N_14433,N_14436,N_14437,N_14438,N_14439,N_14441,N_14442,N_14444,N_14445,N_14446,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14466,N_14467,N_14468,N_14469,N_14471,N_14472,N_14473,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14498,N_14499,N_14500,N_14501,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14513,N_14514,N_14515,N_14517,N_14518,N_14519,N_14520,N_14521,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14549,N_14551,N_14552,N_14553,N_14554,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14563,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14575,N_14576,N_14577,N_14578,N_14579,N_14581,N_14582,N_14583,N_14584,N_14585,N_14587,N_14588,N_14589,N_14590,N_14592,N_14593,N_14594,N_14595,N_14597,N_14599,N_14601,N_14602,N_14603,N_14605,N_14606,N_14607,N_14608,N_14610,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14634,N_14635,N_14636,N_14637,N_14639,N_14641,N_14642,N_14643,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14657,N_14658,N_14659,N_14660,N_14662,N_14663,N_14664,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14674,N_14675,N_14676,N_14677,N_14678,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14699,N_14700,N_14702,N_14703,N_14704,N_14705,N_14706,N_14708,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14738,N_14740,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14762,N_14763,N_14764,N_14765,N_14767,N_14768,N_14769,N_14770,N_14772,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14785,N_14786,N_14787,N_14789,N_14791,N_14792,N_14793,N_14794,N_14795,N_14798,N_14801,N_14804,N_14808,N_14809,N_14810,N_14811,N_14812,N_14814,N_14815,N_14816,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14826,N_14827,N_14828,N_14831,N_14832,N_14833,N_14834,N_14836,N_14837,N_14838,N_14839,N_14841,N_14843,N_14844,N_14845,N_14846,N_14848,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14876,N_14877,N_14878,N_14882,N_14886,N_14887,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14898,N_14899,N_14900,N_14901,N_14903,N_14905,N_14907,N_14909,N_14910,N_14912,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14940,N_14941,N_14942,N_14943,N_14945,N_14946,N_14947,N_14948,N_14949,N_14952,N_14953,N_14955,N_14956,N_14959,N_14960,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14969,N_14972,N_14973,N_14974,N_14975,N_14976,N_14978,N_14979,N_14980,N_14982,N_14984,N_14985,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_566,In_1096);
xor U1 (N_1,In_1107,In_17);
or U2 (N_2,In_1086,In_1487);
nor U3 (N_3,In_28,In_706);
or U4 (N_4,In_1159,In_72);
or U5 (N_5,In_1099,In_798);
and U6 (N_6,In_1040,In_108);
and U7 (N_7,In_784,In_818);
and U8 (N_8,In_1121,In_302);
xnor U9 (N_9,In_387,In_982);
xor U10 (N_10,In_53,In_1043);
nor U11 (N_11,In_13,In_648);
nand U12 (N_12,In_456,In_173);
or U13 (N_13,In_696,In_1452);
nand U14 (N_14,In_628,In_59);
and U15 (N_15,In_1006,In_662);
xnor U16 (N_16,In_211,In_86);
nand U17 (N_17,In_1387,In_144);
xnor U18 (N_18,In_555,In_699);
xor U19 (N_19,In_1325,In_783);
or U20 (N_20,In_484,In_560);
xor U21 (N_21,In_862,In_1402);
and U22 (N_22,In_1477,In_272);
xnor U23 (N_23,In_407,In_329);
xor U24 (N_24,In_604,In_1418);
nand U25 (N_25,In_74,In_1163);
xor U26 (N_26,In_301,In_1364);
nor U27 (N_27,In_1062,In_40);
xor U28 (N_28,In_508,In_1181);
xnor U29 (N_29,In_256,In_1247);
or U30 (N_30,In_747,In_148);
nand U31 (N_31,In_386,In_803);
or U32 (N_32,In_469,In_477);
and U33 (N_33,In_1157,In_522);
xor U34 (N_34,In_889,In_1237);
or U35 (N_35,In_1041,In_1015);
nand U36 (N_36,In_663,In_1125);
nor U37 (N_37,In_182,In_1478);
xor U38 (N_38,In_621,In_330);
nor U39 (N_39,In_1182,In_741);
xnor U40 (N_40,In_828,In_1025);
nor U41 (N_41,In_379,In_1180);
and U42 (N_42,In_929,In_43);
or U43 (N_43,In_757,In_539);
or U44 (N_44,In_760,In_106);
nand U45 (N_45,In_1432,In_1276);
xnor U46 (N_46,In_516,In_579);
or U47 (N_47,In_1369,In_599);
nand U48 (N_48,In_898,In_1162);
and U49 (N_49,In_179,In_135);
nor U50 (N_50,In_138,In_934);
and U51 (N_51,In_219,In_961);
or U52 (N_52,In_25,In_1484);
and U53 (N_53,In_670,In_808);
nor U54 (N_54,In_1372,In_232);
nor U55 (N_55,In_1283,In_492);
xnor U56 (N_56,In_56,In_843);
nand U57 (N_57,In_820,In_1155);
xor U58 (N_58,In_61,In_856);
xor U59 (N_59,In_1227,In_475);
or U60 (N_60,In_117,In_901);
nor U61 (N_61,In_583,In_42);
xor U62 (N_62,In_928,In_447);
nor U63 (N_63,In_1454,In_18);
and U64 (N_64,In_1053,In_78);
and U65 (N_65,In_1021,In_1463);
or U66 (N_66,In_432,In_422);
nand U67 (N_67,In_542,In_831);
nand U68 (N_68,In_515,In_355);
nand U69 (N_69,In_323,In_707);
nor U70 (N_70,In_1442,In_943);
and U71 (N_71,In_999,In_1330);
xor U72 (N_72,In_1289,In_596);
xor U73 (N_73,In_781,In_526);
nor U74 (N_74,In_1279,In_1148);
nor U75 (N_75,In_444,In_580);
or U76 (N_76,In_766,In_708);
or U77 (N_77,In_631,In_639);
or U78 (N_78,In_1116,In_949);
nand U79 (N_79,In_738,In_813);
and U80 (N_80,In_1327,In_45);
or U81 (N_81,In_1368,In_1355);
or U82 (N_82,In_792,In_1490);
xor U83 (N_83,In_367,In_1035);
or U84 (N_84,In_390,In_60);
and U85 (N_85,In_260,In_569);
nor U86 (N_86,In_932,In_1225);
nor U87 (N_87,In_391,In_224);
nand U88 (N_88,In_350,In_689);
nor U89 (N_89,In_673,In_240);
xnor U90 (N_90,In_395,In_1022);
or U91 (N_91,In_38,In_963);
and U92 (N_92,In_491,In_234);
and U93 (N_93,In_1337,In_421);
nand U94 (N_94,In_361,In_554);
nand U95 (N_95,In_1329,In_630);
xnor U96 (N_96,In_47,In_1293);
xnor U97 (N_97,In_352,In_1004);
or U98 (N_98,In_922,In_1098);
or U99 (N_99,In_880,In_279);
and U100 (N_100,In_415,In_490);
nor U101 (N_101,In_75,In_220);
or U102 (N_102,In_80,In_658);
nor U103 (N_103,In_1232,In_1271);
nand U104 (N_104,In_496,In_991);
nand U105 (N_105,In_1353,In_568);
or U106 (N_106,In_607,In_810);
or U107 (N_107,In_561,In_67);
or U108 (N_108,In_845,In_433);
or U109 (N_109,In_890,In_1229);
xor U110 (N_110,In_1095,In_971);
xor U111 (N_111,In_837,In_94);
nor U112 (N_112,In_50,In_557);
and U113 (N_113,In_482,In_692);
nand U114 (N_114,In_251,In_1331);
nor U115 (N_115,In_701,In_328);
or U116 (N_116,In_528,In_112);
xnor U117 (N_117,In_1497,In_1333);
and U118 (N_118,In_170,In_1030);
and U119 (N_119,In_382,In_672);
nor U120 (N_120,In_1071,In_1158);
or U121 (N_121,In_57,In_981);
xor U122 (N_122,In_95,In_1453);
or U123 (N_123,In_996,In_548);
or U124 (N_124,In_129,In_1370);
and U125 (N_125,In_551,In_1458);
nor U126 (N_126,In_521,In_109);
or U127 (N_127,In_1093,In_643);
xnor U128 (N_128,In_545,In_1115);
nor U129 (N_129,In_1019,In_867);
or U130 (N_130,In_461,In_640);
nor U131 (N_131,In_200,In_398);
and U132 (N_132,In_1152,In_720);
or U133 (N_133,In_247,In_917);
or U134 (N_134,In_851,In_869);
nor U135 (N_135,In_962,In_71);
nand U136 (N_136,In_776,In_1020);
nand U137 (N_137,In_1440,In_1304);
nand U138 (N_138,In_1416,In_137);
nand U139 (N_139,In_894,In_1054);
nand U140 (N_140,In_1287,In_1083);
nand U141 (N_141,In_502,In_27);
xor U142 (N_142,In_416,In_574);
and U143 (N_143,In_498,In_474);
and U144 (N_144,In_1184,In_1087);
nand U145 (N_145,In_334,In_752);
or U146 (N_146,In_771,In_925);
or U147 (N_147,In_998,In_1113);
nand U148 (N_148,In_36,In_363);
or U149 (N_149,In_313,In_839);
nand U150 (N_150,In_1036,In_1139);
nor U151 (N_151,In_1081,In_19);
xnor U152 (N_152,In_503,In_1244);
or U153 (N_153,In_1424,In_172);
nor U154 (N_154,In_29,In_543);
nor U155 (N_155,In_846,In_1485);
nand U156 (N_156,In_231,In_742);
xor U157 (N_157,In_429,In_393);
nand U158 (N_158,In_1014,In_1217);
nand U159 (N_159,In_1383,In_202);
nor U160 (N_160,In_91,In_1420);
or U161 (N_161,In_177,In_481);
nor U162 (N_162,In_76,In_312);
and U163 (N_163,In_737,In_331);
or U164 (N_164,In_1316,In_879);
nor U165 (N_165,In_1334,In_1417);
nor U166 (N_166,In_1366,In_1348);
nand U167 (N_167,In_1027,In_1309);
and U168 (N_168,In_800,In_436);
nor U169 (N_169,In_300,In_956);
nor U170 (N_170,In_616,In_921);
or U171 (N_171,In_276,In_980);
or U172 (N_172,In_1307,In_1342);
xor U173 (N_173,In_435,In_473);
and U174 (N_174,In_93,In_1167);
xor U175 (N_175,In_595,In_1018);
xor U176 (N_176,In_605,In_1318);
nor U177 (N_177,In_450,In_1361);
nand U178 (N_178,In_1322,In_400);
nand U179 (N_179,In_228,In_1352);
xor U180 (N_180,In_396,In_1412);
and U181 (N_181,In_212,In_1308);
and U182 (N_182,In_243,In_1142);
nand U183 (N_183,In_1349,In_501);
and U184 (N_184,In_322,In_852);
and U185 (N_185,In_1396,In_1140);
nor U186 (N_186,In_1356,In_622);
xnor U187 (N_187,In_30,In_812);
and U188 (N_188,In_1373,In_48);
and U189 (N_189,In_1038,In_190);
or U190 (N_190,In_479,In_126);
nor U191 (N_191,In_1468,In_855);
or U192 (N_192,In_1431,In_1386);
and U193 (N_193,In_591,In_610);
or U194 (N_194,In_578,In_602);
and U195 (N_195,In_357,In_537);
or U196 (N_196,In_532,In_278);
nor U197 (N_197,In_1210,In_1270);
xnor U198 (N_198,In_446,In_115);
nor U199 (N_199,In_1393,In_1314);
and U200 (N_200,In_295,In_1483);
nand U201 (N_201,In_601,In_1186);
nand U202 (N_202,In_863,In_695);
xnor U203 (N_203,In_1437,In_406);
and U204 (N_204,In_341,In_983);
xnor U205 (N_205,In_1141,In_1010);
or U206 (N_206,In_62,In_634);
nor U207 (N_207,In_385,In_751);
or U208 (N_208,In_1489,In_168);
nand U209 (N_209,In_635,In_1259);
nor U210 (N_210,In_365,In_154);
or U211 (N_211,In_1470,In_1258);
or U212 (N_212,In_266,In_558);
nor U213 (N_213,In_68,In_169);
or U214 (N_214,In_426,In_32);
and U215 (N_215,In_957,In_891);
and U216 (N_216,In_1112,In_665);
xnor U217 (N_217,In_966,In_158);
xor U218 (N_218,In_1436,In_1100);
and U219 (N_219,In_793,In_586);
and U220 (N_220,In_589,In_656);
or U221 (N_221,In_320,In_1132);
xnor U222 (N_222,In_1428,In_726);
xnor U223 (N_223,In_1242,In_1301);
nor U224 (N_224,In_1223,In_754);
xnor U225 (N_225,In_1438,In_1255);
xnor U226 (N_226,In_11,In_703);
or U227 (N_227,In_1039,In_759);
xnor U228 (N_228,In_134,In_209);
nor U229 (N_229,In_33,In_788);
or U230 (N_230,In_1400,In_609);
or U231 (N_231,In_1060,In_324);
and U232 (N_232,In_1187,In_413);
or U233 (N_233,In_1399,In_253);
xor U234 (N_234,In_505,In_124);
or U235 (N_235,In_442,In_1291);
xnor U236 (N_236,In_12,In_414);
nor U237 (N_237,In_1084,In_1492);
xor U238 (N_238,In_215,In_1042);
and U239 (N_239,In_1066,In_920);
nor U240 (N_240,In_684,In_1074);
nor U241 (N_241,In_1249,In_1268);
and U242 (N_242,In_318,In_1192);
nand U243 (N_243,In_1389,In_1392);
nor U244 (N_244,In_1034,In_1195);
or U245 (N_245,In_466,In_1029);
nor U246 (N_246,In_517,In_440);
and U247 (N_247,In_778,In_1257);
and U248 (N_248,In_919,In_1310);
nand U249 (N_249,In_372,In_1008);
and U250 (N_250,In_1124,In_121);
nand U251 (N_251,In_1292,In_66);
or U252 (N_252,In_1415,In_875);
nor U253 (N_253,In_1009,In_1168);
xnor U254 (N_254,In_1441,In_651);
nor U255 (N_255,In_822,In_55);
or U256 (N_256,In_139,In_369);
nand U257 (N_257,In_308,In_499);
or U258 (N_258,In_368,In_1344);
and U259 (N_259,In_785,In_773);
or U260 (N_260,In_418,In_685);
nand U261 (N_261,In_805,In_175);
nor U262 (N_262,In_735,In_1434);
nand U263 (N_263,In_676,In_1089);
and U264 (N_264,In_1256,In_404);
nand U265 (N_265,In_235,In_1120);
nor U266 (N_266,In_834,In_1494);
nand U267 (N_267,In_1376,In_277);
or U268 (N_268,In_1446,In_697);
nand U269 (N_269,In_1456,In_723);
nor U270 (N_270,In_326,In_1179);
nor U271 (N_271,In_0,In_1090);
or U272 (N_272,In_509,In_188);
nand U273 (N_273,In_252,In_988);
nand U274 (N_274,In_1126,In_96);
and U275 (N_275,In_840,In_314);
nand U276 (N_276,In_1164,In_575);
nand U277 (N_277,In_455,In_1384);
nor U278 (N_278,In_1243,In_582);
nand U279 (N_279,In_1178,In_304);
nand U280 (N_280,In_1103,In_958);
nand U281 (N_281,In_487,In_1153);
nand U282 (N_282,In_1226,In_1101);
xor U283 (N_283,In_608,In_281);
nor U284 (N_284,In_930,In_1231);
and U285 (N_285,In_947,In_675);
nand U286 (N_286,In_270,In_791);
or U287 (N_287,In_530,In_222);
xor U288 (N_288,In_842,In_687);
nand U289 (N_289,In_512,In_571);
nand U290 (N_290,In_23,In_122);
and U291 (N_291,In_1207,In_241);
and U292 (N_292,In_397,In_1350);
and U293 (N_293,In_1003,In_1050);
nand U294 (N_294,In_293,In_133);
or U295 (N_295,In_772,In_1273);
nor U296 (N_296,In_223,In_176);
nor U297 (N_297,In_1080,In_375);
or U298 (N_298,In_916,In_1251);
nor U299 (N_299,In_208,In_192);
nand U300 (N_300,In_289,In_1254);
or U301 (N_301,In_632,In_495);
xor U302 (N_302,In_1149,In_832);
xor U303 (N_303,In_739,In_162);
and U304 (N_304,In_908,In_1421);
nand U305 (N_305,In_335,In_1471);
nor U306 (N_306,In_815,In_373);
or U307 (N_307,In_716,In_1013);
nor U308 (N_308,In_242,In_437);
nor U309 (N_309,In_199,In_360);
or U310 (N_310,In_448,In_948);
or U311 (N_311,In_1445,In_1144);
nor U312 (N_312,In_1374,In_1351);
nor U313 (N_313,In_915,In_953);
and U314 (N_314,In_912,In_693);
nor U315 (N_315,In_633,In_721);
xor U316 (N_316,In_1375,In_160);
or U317 (N_317,In_860,In_1209);
or U318 (N_318,In_668,In_1215);
and U319 (N_319,In_306,In_857);
nor U320 (N_320,In_615,In_213);
xnor U321 (N_321,In_873,In_258);
and U322 (N_322,In_841,In_1151);
nand U323 (N_323,In_7,In_1323);
and U324 (N_324,In_906,In_58);
xor U325 (N_325,In_394,In_893);
or U326 (N_326,In_205,In_248);
nor U327 (N_327,In_618,In_489);
xnor U328 (N_328,In_1092,In_853);
or U329 (N_329,In_140,In_1341);
xor U330 (N_330,In_1185,In_885);
nor U331 (N_331,In_65,In_339);
nor U332 (N_332,In_606,In_1447);
nand U333 (N_333,In_698,In_1338);
xnor U334 (N_334,In_644,In_180);
xnor U335 (N_335,In_1295,In_700);
or U336 (N_336,In_844,In_283);
xnor U337 (N_337,In_1306,In_682);
nor U338 (N_338,In_494,In_54);
nor U339 (N_339,In_995,In_585);
nor U340 (N_340,In_340,In_567);
xnor U341 (N_341,In_1024,In_49);
nor U342 (N_342,In_287,In_770);
nand U343 (N_343,In_1413,In_854);
xnor U344 (N_344,In_736,In_904);
and U345 (N_345,In_214,In_730);
nand U346 (N_346,In_233,In_364);
nor U347 (N_347,In_826,In_1057);
nor U348 (N_348,In_165,In_657);
and U349 (N_349,In_1114,In_167);
or U350 (N_350,In_729,In_1065);
nand U351 (N_351,In_523,In_303);
xor U352 (N_352,In_954,In_577);
xnor U353 (N_353,In_1193,In_125);
nand U354 (N_354,In_1346,In_10);
or U355 (N_355,In_1406,In_46);
nor U356 (N_356,In_924,In_1319);
xnor U357 (N_357,In_811,In_1320);
nand U358 (N_358,In_681,In_311);
nor U359 (N_359,In_1390,In_1200);
nand U360 (N_360,In_753,In_882);
nand U361 (N_361,In_927,In_659);
xor U362 (N_362,In_614,In_598);
nor U363 (N_363,In_319,In_1281);
and U364 (N_364,In_733,In_679);
nand U365 (N_365,In_1462,In_1052);
and U366 (N_366,In_102,In_305);
xnor U367 (N_367,In_110,In_892);
and U368 (N_368,In_556,In_409);
nor U369 (N_369,In_524,In_250);
nand U370 (N_370,In_835,In_774);
nor U371 (N_371,In_143,In_1260);
nand U372 (N_372,In_178,In_207);
nor U373 (N_373,In_381,In_1457);
nand U374 (N_374,In_849,In_288);
and U375 (N_375,In_768,In_1422);
xnor U376 (N_376,In_1482,In_359);
xor U377 (N_377,In_913,In_861);
nor U378 (N_378,In_203,In_206);
nor U379 (N_379,In_732,In_1377);
xnor U380 (N_380,In_443,In_244);
xnor U381 (N_381,In_1105,In_236);
and U382 (N_382,In_1357,In_787);
xnor U383 (N_383,In_85,In_819);
nor U384 (N_384,In_864,In_338);
xor U385 (N_385,In_533,In_171);
or U386 (N_386,In_21,In_1297);
nand U387 (N_387,In_540,In_1343);
xnor U388 (N_388,In_358,In_597);
nor U389 (N_389,In_1480,In_717);
or U390 (N_390,In_1068,In_297);
xnor U391 (N_391,In_119,In_186);
and U392 (N_392,In_83,In_677);
or U393 (N_393,In_789,In_467);
or U394 (N_394,In_384,In_713);
and U395 (N_395,In_550,In_1439);
and U396 (N_396,In_902,In_1206);
xnor U397 (N_397,In_325,In_346);
and U398 (N_398,In_1423,In_198);
nor U399 (N_399,In_950,In_128);
nand U400 (N_400,In_127,In_638);
xor U401 (N_401,In_1133,In_1430);
xor U402 (N_402,In_189,In_830);
and U403 (N_403,In_1028,In_1302);
or U404 (N_404,In_588,In_594);
and U405 (N_405,In_118,In_749);
xnor U406 (N_406,In_529,In_249);
or U407 (N_407,In_430,In_113);
nand U408 (N_408,In_645,In_777);
nand U409 (N_409,In_976,In_955);
nor U410 (N_410,In_419,In_427);
and U411 (N_411,In_1267,In_1411);
xnor U412 (N_412,In_184,In_1380);
and U413 (N_413,In_485,In_1236);
nor U414 (N_414,In_1177,In_1194);
nand U415 (N_415,In_868,In_725);
xor U416 (N_416,In_1241,In_1363);
or U417 (N_417,In_1174,In_52);
nand U418 (N_418,In_1203,In_458);
and U419 (N_419,In_411,In_1212);
nand U420 (N_420,In_1044,In_507);
and U421 (N_421,In_967,In_896);
or U422 (N_422,In_1051,In_518);
xor U423 (N_423,In_1001,In_1026);
nor U424 (N_424,In_333,In_513);
and U425 (N_425,In_973,In_1138);
or U426 (N_426,In_1303,In_1197);
nand U427 (N_427,In_472,In_895);
nand U428 (N_428,In_470,In_153);
or U429 (N_429,In_187,In_653);
nand U430 (N_430,In_370,In_1444);
nor U431 (N_431,In_1311,In_309);
or U432 (N_432,In_587,In_945);
or U433 (N_433,In_878,In_756);
and U434 (N_434,In_1261,In_100);
nor U435 (N_435,In_691,In_1127);
nand U436 (N_436,In_1294,In_226);
nor U437 (N_437,In_420,In_41);
nand U438 (N_438,In_259,In_275);
nand U439 (N_439,In_116,In_745);
nor U440 (N_440,In_87,In_412);
or U441 (N_441,In_463,In_592);
or U442 (N_442,In_960,In_459);
xor U443 (N_443,In_709,In_183);
xnor U444 (N_444,In_977,In_923);
or U445 (N_445,In_1448,In_541);
nor U446 (N_446,In_918,In_762);
nand U447 (N_447,In_796,In_1239);
xor U448 (N_448,In_342,In_221);
or U449 (N_449,In_559,In_194);
xor U450 (N_450,In_870,In_16);
nor U451 (N_451,In_402,In_850);
xnor U452 (N_452,In_2,In_1064);
xor U453 (N_453,In_683,In_1296);
xor U454 (N_454,In_1136,In_625);
or U455 (N_455,In_1154,In_1262);
and U456 (N_456,In_666,In_1213);
nor U457 (N_457,In_1037,In_510);
nand U458 (N_458,In_974,In_1070);
or U459 (N_459,In_1016,In_1102);
nor U460 (N_460,In_264,In_356);
or U461 (N_461,In_377,In_984);
or U462 (N_462,In_911,In_197);
nand U463 (N_463,In_1464,In_994);
or U464 (N_464,In_1228,In_1085);
and U465 (N_465,In_859,In_1216);
and U466 (N_466,In_823,In_1449);
or U467 (N_467,In_702,In_1118);
or U468 (N_468,In_1094,In_1312);
and U469 (N_469,In_99,In_553);
xnor U470 (N_470,In_201,In_268);
nor U471 (N_471,In_1011,In_824);
nor U472 (N_472,In_1298,In_239);
xor U473 (N_473,In_63,In_858);
nand U474 (N_474,In_727,In_722);
xnor U475 (N_475,In_669,In_1173);
nand U476 (N_476,In_590,In_979);
or U477 (N_477,In_185,In_1046);
or U478 (N_478,In_1201,In_89);
xor U479 (N_479,In_344,In_978);
and U480 (N_480,In_989,In_262);
nand U481 (N_481,In_1069,In_576);
nand U482 (N_482,In_619,In_1275);
or U483 (N_483,In_655,In_1474);
and U484 (N_484,In_1278,In_196);
xor U485 (N_485,In_1450,In_1077);
nor U486 (N_486,In_14,In_775);
or U487 (N_487,In_1465,In_937);
and U488 (N_488,In_649,In_88);
or U489 (N_489,In_1313,In_1233);
xor U490 (N_490,In_686,In_990);
and U491 (N_491,In_82,In_1479);
xnor U492 (N_492,In_159,In_620);
nand U493 (N_493,In_1460,In_968);
nand U494 (N_494,In_98,In_806);
and U495 (N_495,In_1335,In_438);
and U496 (N_496,In_1495,In_876);
xor U497 (N_497,In_718,In_969);
and U498 (N_498,In_972,In_941);
xnor U499 (N_499,In_802,In_1245);
nand U500 (N_500,In_804,In_1385);
and U501 (N_501,In_1111,In_1145);
and U502 (N_502,In_1317,In_514);
or U503 (N_503,In_1122,In_424);
and U504 (N_504,In_809,In_265);
and U505 (N_505,In_299,In_688);
and U506 (N_506,In_1345,In_1476);
nand U507 (N_507,In_678,In_97);
and U508 (N_508,In_807,In_44);
xnor U509 (N_509,In_821,In_1147);
nand U510 (N_510,In_1461,In_204);
or U511 (N_511,In_714,In_546);
and U512 (N_512,In_1403,In_603);
or U513 (N_513,In_343,In_39);
nand U514 (N_514,In_1191,In_650);
and U515 (N_515,In_69,In_1367);
and U516 (N_516,In_1117,In_1328);
and U517 (N_517,In_1156,In_536);
or U518 (N_518,In_291,In_1204);
nand U519 (N_519,In_1360,In_1425);
or U520 (N_520,In_1097,In_157);
xnor U521 (N_521,In_769,In_1176);
xnor U522 (N_522,In_786,In_1214);
nand U523 (N_523,In_146,In_131);
nand U524 (N_524,In_337,In_354);
or U525 (N_525,In_403,In_1202);
nor U526 (N_526,In_105,In_938);
and U527 (N_527,In_1410,In_156);
and U528 (N_528,In_626,In_81);
or U529 (N_529,In_1175,In_1002);
or U530 (N_530,In_900,In_1059);
nand U531 (N_531,In_1129,In_1196);
nor U532 (N_532,In_531,In_1288);
nor U533 (N_533,In_1171,In_674);
xor U534 (N_534,In_195,In_1012);
or U535 (N_535,In_975,In_103);
or U536 (N_536,In_1079,In_431);
or U537 (N_537,In_600,In_660);
and U538 (N_538,In_405,In_827);
nor U539 (N_539,In_1221,In_1272);
nand U540 (N_540,In_881,In_51);
and U541 (N_541,In_1473,In_1378);
nor U542 (N_542,In_1250,In_84);
nand U543 (N_543,In_452,In_926);
and U544 (N_544,In_336,In_952);
or U545 (N_545,In_497,In_1045);
and U546 (N_546,In_959,In_1286);
xnor U547 (N_547,In_3,In_993);
nand U548 (N_548,In_480,In_936);
xor U549 (N_549,In_935,In_210);
and U550 (N_550,In_1189,In_163);
nand U551 (N_551,In_883,In_573);
or U552 (N_552,In_246,In_145);
xnor U553 (N_553,In_903,In_1198);
and U554 (N_554,In_286,In_794);
and U555 (N_555,In_641,In_1326);
and U556 (N_556,In_149,In_1466);
and U557 (N_557,In_1072,In_1280);
nand U558 (N_558,In_1467,In_761);
nand U559 (N_559,In_1486,In_24);
nand U560 (N_560,In_1211,In_1205);
nor U561 (N_561,In_150,In_970);
xor U562 (N_562,In_801,In_1091);
or U563 (N_563,In_942,In_1419);
xor U564 (N_564,In_401,In_392);
or U565 (N_565,In_1119,In_1208);
nand U566 (N_566,In_345,In_562);
and U567 (N_567,In_410,In_1190);
xor U568 (N_568,In_445,In_1253);
xnor U569 (N_569,In_255,In_4);
nor U570 (N_570,In_1248,In_940);
or U571 (N_571,In_1224,In_1031);
nor U572 (N_572,In_230,In_1381);
or U573 (N_573,In_374,In_848);
nor U574 (N_574,In_1498,In_267);
xor U575 (N_575,In_817,In_570);
xor U576 (N_576,In_292,In_296);
nand U577 (N_577,In_453,In_1265);
nand U578 (N_578,In_77,In_130);
xnor U579 (N_579,In_728,In_1023);
nor U580 (N_580,In_1235,In_504);
nor U581 (N_581,In_572,In_1274);
and U582 (N_582,In_767,In_191);
nor U583 (N_583,In_611,In_1398);
nor U584 (N_584,In_642,In_1332);
xor U585 (N_585,In_327,In_1073);
and U586 (N_586,In_64,In_1240);
nor U587 (N_587,In_1063,In_298);
nor U588 (N_588,In_174,In_886);
nand U589 (N_589,In_1188,In_871);
nor U590 (N_590,In_1161,In_1305);
nand U591 (N_591,In_376,In_1088);
nand U592 (N_592,In_1000,In_120);
xor U593 (N_593,In_525,In_471);
or U594 (N_594,In_1362,In_1131);
xnor U595 (N_595,In_238,In_617);
nand U596 (N_596,In_269,In_1282);
and U597 (N_597,In_1277,In_1172);
and U598 (N_598,In_910,In_389);
or U599 (N_599,In_9,In_613);
nor U600 (N_600,In_181,In_1427);
xnor U601 (N_601,In_1339,In_464);
nor U602 (N_602,In_944,In_1455);
or U603 (N_603,In_1222,In_1382);
and U604 (N_604,In_887,In_70);
or U605 (N_605,In_1252,In_321);
nor U606 (N_606,In_765,In_26);
xnor U607 (N_607,In_245,In_740);
and U608 (N_608,In_476,In_1108);
nand U609 (N_609,In_667,In_1166);
nand U610 (N_610,In_434,In_671);
nor U611 (N_611,In_520,In_166);
nand U612 (N_612,In_1238,In_782);
or U613 (N_613,In_141,In_15);
nand U614 (N_614,In_425,In_865);
and U615 (N_615,In_1299,In_985);
nand U616 (N_616,In_274,In_1005);
nand U617 (N_617,In_31,In_1146);
xor U618 (N_618,In_284,In_1429);
nand U619 (N_619,In_1391,In_997);
and U620 (N_620,In_680,In_462);
nor U621 (N_621,In_227,In_22);
nand U622 (N_622,In_280,In_899);
nand U623 (N_623,In_564,In_294);
xnor U624 (N_624,In_1049,In_866);
and U625 (N_625,In_914,In_1408);
xnor U626 (N_626,In_290,In_1426);
and U627 (N_627,In_1358,In_347);
and U628 (N_628,In_1143,In_388);
and U629 (N_629,In_282,In_884);
nand U630 (N_630,In_511,In_1414);
xor U631 (N_631,In_483,In_1150);
or U632 (N_632,In_353,In_833);
and U633 (N_633,In_399,In_317);
nand U634 (N_634,In_1365,In_654);
xnor U635 (N_635,In_519,In_34);
and U636 (N_636,In_1032,In_457);
nand U637 (N_637,In_451,In_549);
or U638 (N_638,In_1379,In_711);
or U639 (N_639,In_612,In_1493);
or U640 (N_640,In_1324,In_1048);
xor U641 (N_641,In_1169,In_563);
or U642 (N_642,In_101,In_694);
nor U643 (N_643,In_1459,In_731);
nor U644 (N_644,In_652,In_1472);
nor U645 (N_645,In_1128,In_1104);
or U646 (N_646,In_744,In_271);
nand U647 (N_647,In_261,In_1218);
nand U648 (N_648,In_986,In_623);
nor U649 (N_649,In_423,In_1404);
or U650 (N_650,In_951,In_763);
xor U651 (N_651,In_946,In_1170);
nand U652 (N_652,In_362,In_629);
or U653 (N_653,In_1481,In_1183);
xor U654 (N_654,In_829,In_132);
and U655 (N_655,In_565,In_547);
or U656 (N_656,In_1082,In_161);
or U657 (N_657,In_454,In_1220);
or U658 (N_658,In_1246,In_1266);
or U659 (N_659,In_1135,In_1263);
or U660 (N_660,In_366,In_965);
nor U661 (N_661,In_104,In_1130);
nand U662 (N_662,In_351,In_1300);
or U663 (N_663,In_1433,In_734);
nor U664 (N_664,In_1137,In_705);
nand U665 (N_665,In_217,In_90);
or U666 (N_666,In_332,In_1078);
nand U667 (N_667,In_748,In_1475);
nor U668 (N_668,In_229,In_593);
and U669 (N_669,In_1285,In_710);
nand U670 (N_670,In_316,In_1491);
and U671 (N_671,In_838,In_193);
nand U672 (N_672,In_1076,In_897);
xor U673 (N_673,In_719,In_378);
nand U674 (N_674,In_535,In_380);
nor U675 (N_675,In_500,In_1397);
nor U676 (N_676,In_114,In_872);
nor U677 (N_677,In_816,In_1388);
nand U678 (N_678,In_661,In_825);
and U679 (N_679,In_704,In_1075);
nand U680 (N_680,In_493,In_1340);
xnor U681 (N_681,In_646,In_307);
or U682 (N_682,In_1496,In_743);
and U683 (N_683,In_35,In_315);
nand U684 (N_684,In_1315,In_147);
or U685 (N_685,In_449,In_814);
or U686 (N_686,In_1401,In_584);
xor U687 (N_687,In_724,In_371);
and U688 (N_688,In_136,In_428);
nand U689 (N_689,In_764,In_1134);
xnor U690 (N_690,In_285,In_1269);
xor U691 (N_691,In_383,In_715);
nand U692 (N_692,In_1007,In_439);
xor U693 (N_693,In_1047,In_664);
or U694 (N_694,In_488,In_874);
nand U695 (N_695,In_152,In_797);
nand U696 (N_696,In_690,In_37);
nor U697 (N_697,In_1110,In_799);
xnor U698 (N_698,In_417,In_758);
or U699 (N_699,In_1058,In_478);
nand U700 (N_700,In_527,In_225);
xor U701 (N_701,In_506,In_581);
nand U702 (N_702,In_1109,In_1321);
and U703 (N_703,In_1199,In_1354);
and U704 (N_704,In_987,In_1469);
nand U705 (N_705,In_1290,In_647);
and U706 (N_706,In_712,In_1234);
xnor U707 (N_707,In_6,In_847);
xor U708 (N_708,In_273,In_1);
or U709 (N_709,In_750,In_1394);
nand U710 (N_710,In_155,In_218);
or U711 (N_711,In_1435,In_534);
xor U712 (N_712,In_636,In_1488);
nand U713 (N_713,In_1056,In_907);
and U714 (N_714,In_111,In_780);
nand U715 (N_715,In_142,In_909);
and U716 (N_716,In_755,In_552);
and U717 (N_717,In_1061,In_888);
xnor U718 (N_718,In_1106,In_1451);
xnor U719 (N_719,In_1395,In_465);
xnor U720 (N_720,In_92,In_5);
or U721 (N_721,In_263,In_964);
nor U722 (N_722,In_746,In_790);
or U723 (N_723,In_257,In_1165);
nor U724 (N_724,In_933,In_931);
xnor U725 (N_725,In_1160,In_349);
xor U726 (N_726,In_310,In_151);
nand U727 (N_727,In_1264,In_1017);
xor U728 (N_728,In_441,In_486);
nor U729 (N_729,In_795,In_1123);
nor U730 (N_730,In_538,In_836);
nand U731 (N_731,In_79,In_1347);
nor U732 (N_732,In_877,In_1055);
and U733 (N_733,In_1067,In_992);
nor U734 (N_734,In_779,In_1230);
and U735 (N_735,In_939,In_1033);
or U736 (N_736,In_73,In_123);
nor U737 (N_737,In_905,In_1219);
and U738 (N_738,In_1336,In_1359);
xnor U739 (N_739,In_624,In_460);
or U740 (N_740,In_216,In_20);
or U741 (N_741,In_107,In_1405);
or U742 (N_742,In_627,In_1407);
xor U743 (N_743,In_237,In_254);
xnor U744 (N_744,In_1499,In_468);
nand U745 (N_745,In_1371,In_348);
and U746 (N_746,In_1443,In_637);
and U747 (N_747,In_1409,In_544);
nand U748 (N_748,In_164,In_8);
and U749 (N_749,In_408,In_1284);
and U750 (N_750,In_835,In_532);
xnor U751 (N_751,In_1146,In_1304);
nor U752 (N_752,In_215,In_1211);
nand U753 (N_753,In_1392,In_604);
xnor U754 (N_754,In_239,In_144);
or U755 (N_755,In_148,In_175);
nor U756 (N_756,In_1468,In_410);
nor U757 (N_757,In_349,In_1092);
nor U758 (N_758,In_1330,In_777);
nand U759 (N_759,In_193,In_1463);
and U760 (N_760,In_1198,In_1361);
and U761 (N_761,In_613,In_1331);
nand U762 (N_762,In_801,In_1497);
nor U763 (N_763,In_1261,In_477);
and U764 (N_764,In_527,In_721);
xor U765 (N_765,In_336,In_791);
nand U766 (N_766,In_244,In_64);
and U767 (N_767,In_1302,In_437);
nand U768 (N_768,In_1090,In_1231);
nor U769 (N_769,In_104,In_945);
xnor U770 (N_770,In_443,In_485);
nand U771 (N_771,In_382,In_114);
and U772 (N_772,In_978,In_318);
xnor U773 (N_773,In_1180,In_213);
xnor U774 (N_774,In_1193,In_1286);
nor U775 (N_775,In_1176,In_938);
or U776 (N_776,In_1082,In_9);
and U777 (N_777,In_171,In_375);
xor U778 (N_778,In_247,In_1008);
or U779 (N_779,In_990,In_484);
xnor U780 (N_780,In_1489,In_25);
and U781 (N_781,In_1153,In_336);
nand U782 (N_782,In_455,In_1163);
or U783 (N_783,In_198,In_622);
and U784 (N_784,In_1221,In_1181);
xnor U785 (N_785,In_291,In_1183);
and U786 (N_786,In_1494,In_1314);
nand U787 (N_787,In_312,In_1019);
xor U788 (N_788,In_390,In_428);
nand U789 (N_789,In_404,In_934);
xnor U790 (N_790,In_591,In_1459);
or U791 (N_791,In_623,In_1318);
nand U792 (N_792,In_1265,In_210);
xnor U793 (N_793,In_161,In_1219);
nor U794 (N_794,In_701,In_1286);
nand U795 (N_795,In_199,In_1227);
nor U796 (N_796,In_581,In_779);
and U797 (N_797,In_767,In_810);
or U798 (N_798,In_868,In_1265);
xnor U799 (N_799,In_9,In_422);
and U800 (N_800,In_1347,In_74);
nand U801 (N_801,In_801,In_286);
and U802 (N_802,In_1399,In_911);
xnor U803 (N_803,In_809,In_1056);
or U804 (N_804,In_169,In_613);
and U805 (N_805,In_1415,In_275);
and U806 (N_806,In_860,In_170);
nand U807 (N_807,In_672,In_598);
nand U808 (N_808,In_948,In_612);
xnor U809 (N_809,In_829,In_1454);
xor U810 (N_810,In_819,In_321);
xnor U811 (N_811,In_260,In_1476);
nor U812 (N_812,In_17,In_1246);
nor U813 (N_813,In_336,In_1175);
and U814 (N_814,In_434,In_128);
xnor U815 (N_815,In_499,In_171);
nand U816 (N_816,In_427,In_95);
nor U817 (N_817,In_1367,In_1456);
and U818 (N_818,In_1480,In_442);
nand U819 (N_819,In_442,In_834);
or U820 (N_820,In_633,In_227);
nor U821 (N_821,In_580,In_1284);
or U822 (N_822,In_1485,In_1477);
nand U823 (N_823,In_36,In_871);
nor U824 (N_824,In_431,In_1296);
nand U825 (N_825,In_485,In_496);
or U826 (N_826,In_1277,In_932);
and U827 (N_827,In_1130,In_1120);
nand U828 (N_828,In_451,In_789);
nand U829 (N_829,In_995,In_1473);
or U830 (N_830,In_852,In_834);
or U831 (N_831,In_1259,In_1199);
nor U832 (N_832,In_887,In_1018);
and U833 (N_833,In_18,In_588);
and U834 (N_834,In_726,In_172);
nand U835 (N_835,In_201,In_126);
xnor U836 (N_836,In_1396,In_74);
nand U837 (N_837,In_702,In_709);
nand U838 (N_838,In_993,In_748);
nor U839 (N_839,In_56,In_739);
nor U840 (N_840,In_331,In_1214);
nand U841 (N_841,In_769,In_991);
and U842 (N_842,In_1252,In_552);
or U843 (N_843,In_1442,In_144);
and U844 (N_844,In_711,In_908);
xor U845 (N_845,In_1478,In_1462);
and U846 (N_846,In_1486,In_1266);
xnor U847 (N_847,In_34,In_652);
nor U848 (N_848,In_332,In_271);
and U849 (N_849,In_263,In_1485);
or U850 (N_850,In_1465,In_1454);
and U851 (N_851,In_8,In_1286);
nand U852 (N_852,In_1281,In_721);
nand U853 (N_853,In_865,In_257);
or U854 (N_854,In_1054,In_605);
or U855 (N_855,In_1392,In_60);
and U856 (N_856,In_751,In_1202);
xnor U857 (N_857,In_779,In_230);
xnor U858 (N_858,In_765,In_629);
and U859 (N_859,In_465,In_1228);
and U860 (N_860,In_124,In_585);
xor U861 (N_861,In_776,In_1281);
or U862 (N_862,In_1418,In_671);
or U863 (N_863,In_246,In_186);
nor U864 (N_864,In_822,In_91);
nand U865 (N_865,In_1481,In_96);
nand U866 (N_866,In_533,In_557);
nor U867 (N_867,In_372,In_715);
nand U868 (N_868,In_324,In_1042);
or U869 (N_869,In_482,In_1376);
nand U870 (N_870,In_833,In_430);
xnor U871 (N_871,In_60,In_630);
xnor U872 (N_872,In_407,In_595);
and U873 (N_873,In_81,In_211);
nand U874 (N_874,In_257,In_157);
xor U875 (N_875,In_1454,In_295);
nor U876 (N_876,In_516,In_830);
nor U877 (N_877,In_601,In_266);
nor U878 (N_878,In_1260,In_1186);
nand U879 (N_879,In_838,In_1157);
nand U880 (N_880,In_1095,In_305);
nor U881 (N_881,In_845,In_1244);
xor U882 (N_882,In_1282,In_1490);
nand U883 (N_883,In_486,In_412);
nand U884 (N_884,In_1406,In_240);
or U885 (N_885,In_1189,In_1461);
nand U886 (N_886,In_146,In_1022);
nand U887 (N_887,In_1332,In_1328);
and U888 (N_888,In_1184,In_974);
xnor U889 (N_889,In_560,In_1279);
xnor U890 (N_890,In_150,In_935);
nand U891 (N_891,In_258,In_1129);
xor U892 (N_892,In_427,In_114);
or U893 (N_893,In_1422,In_1212);
or U894 (N_894,In_1006,In_754);
or U895 (N_895,In_961,In_375);
xor U896 (N_896,In_351,In_1446);
or U897 (N_897,In_73,In_226);
and U898 (N_898,In_674,In_811);
or U899 (N_899,In_311,In_154);
nand U900 (N_900,In_216,In_808);
nor U901 (N_901,In_949,In_215);
or U902 (N_902,In_757,In_301);
or U903 (N_903,In_909,In_758);
and U904 (N_904,In_837,In_1369);
xnor U905 (N_905,In_858,In_1478);
nor U906 (N_906,In_504,In_1490);
xor U907 (N_907,In_309,In_557);
xor U908 (N_908,In_1247,In_814);
xor U909 (N_909,In_510,In_430);
xnor U910 (N_910,In_994,In_877);
and U911 (N_911,In_629,In_750);
or U912 (N_912,In_1467,In_266);
and U913 (N_913,In_275,In_833);
and U914 (N_914,In_1447,In_120);
nor U915 (N_915,In_4,In_724);
nor U916 (N_916,In_649,In_943);
nor U917 (N_917,In_1126,In_944);
nand U918 (N_918,In_1189,In_1111);
nor U919 (N_919,In_18,In_386);
xor U920 (N_920,In_429,In_952);
and U921 (N_921,In_788,In_864);
xor U922 (N_922,In_163,In_1390);
or U923 (N_923,In_1474,In_645);
xor U924 (N_924,In_1434,In_897);
xor U925 (N_925,In_1009,In_506);
and U926 (N_926,In_1025,In_421);
or U927 (N_927,In_129,In_95);
or U928 (N_928,In_1163,In_1242);
nor U929 (N_929,In_695,In_389);
nand U930 (N_930,In_1138,In_476);
xor U931 (N_931,In_1212,In_157);
or U932 (N_932,In_1003,In_733);
xnor U933 (N_933,In_729,In_924);
nor U934 (N_934,In_404,In_1168);
or U935 (N_935,In_321,In_953);
nand U936 (N_936,In_751,In_202);
nor U937 (N_937,In_1416,In_1100);
xnor U938 (N_938,In_358,In_255);
and U939 (N_939,In_345,In_323);
xnor U940 (N_940,In_1423,In_639);
and U941 (N_941,In_445,In_1451);
xor U942 (N_942,In_627,In_156);
or U943 (N_943,In_447,In_1289);
nand U944 (N_944,In_679,In_524);
or U945 (N_945,In_1221,In_1230);
nand U946 (N_946,In_900,In_775);
and U947 (N_947,In_103,In_87);
xnor U948 (N_948,In_522,In_820);
nor U949 (N_949,In_399,In_876);
nor U950 (N_950,In_1143,In_1240);
xnor U951 (N_951,In_284,In_500);
xor U952 (N_952,In_356,In_1451);
nor U953 (N_953,In_79,In_1479);
and U954 (N_954,In_172,In_184);
nand U955 (N_955,In_857,In_1478);
nor U956 (N_956,In_523,In_125);
nor U957 (N_957,In_1309,In_8);
nand U958 (N_958,In_1400,In_1195);
or U959 (N_959,In_234,In_979);
nand U960 (N_960,In_1000,In_334);
and U961 (N_961,In_702,In_1078);
nand U962 (N_962,In_1415,In_415);
nor U963 (N_963,In_487,In_590);
and U964 (N_964,In_30,In_135);
nand U965 (N_965,In_1155,In_1085);
or U966 (N_966,In_656,In_720);
xnor U967 (N_967,In_1230,In_1047);
and U968 (N_968,In_1346,In_261);
and U969 (N_969,In_1111,In_232);
or U970 (N_970,In_545,In_502);
xnor U971 (N_971,In_490,In_380);
xnor U972 (N_972,In_705,In_1302);
nor U973 (N_973,In_944,In_560);
or U974 (N_974,In_298,In_754);
nor U975 (N_975,In_869,In_835);
xor U976 (N_976,In_538,In_1099);
nor U977 (N_977,In_279,In_87);
and U978 (N_978,In_465,In_928);
xor U979 (N_979,In_249,In_1190);
and U980 (N_980,In_656,In_133);
nor U981 (N_981,In_498,In_866);
xor U982 (N_982,In_654,In_1451);
nand U983 (N_983,In_415,In_406);
nand U984 (N_984,In_617,In_854);
xor U985 (N_985,In_338,In_306);
or U986 (N_986,In_641,In_76);
xnor U987 (N_987,In_1207,In_748);
and U988 (N_988,In_686,In_218);
nor U989 (N_989,In_194,In_456);
or U990 (N_990,In_226,In_63);
and U991 (N_991,In_816,In_567);
xor U992 (N_992,In_684,In_1422);
or U993 (N_993,In_245,In_774);
and U994 (N_994,In_1118,In_1491);
and U995 (N_995,In_357,In_665);
and U996 (N_996,In_405,In_585);
nor U997 (N_997,In_715,In_520);
xor U998 (N_998,In_572,In_1407);
or U999 (N_999,In_1306,In_603);
nor U1000 (N_1000,In_359,In_890);
nand U1001 (N_1001,In_940,In_183);
nor U1002 (N_1002,In_590,In_1411);
xnor U1003 (N_1003,In_1247,In_1227);
or U1004 (N_1004,In_897,In_309);
nor U1005 (N_1005,In_314,In_1445);
and U1006 (N_1006,In_1043,In_417);
or U1007 (N_1007,In_869,In_930);
or U1008 (N_1008,In_172,In_670);
nor U1009 (N_1009,In_680,In_373);
nand U1010 (N_1010,In_1392,In_855);
xnor U1011 (N_1011,In_1245,In_475);
nor U1012 (N_1012,In_961,In_381);
or U1013 (N_1013,In_1303,In_1232);
nor U1014 (N_1014,In_1478,In_693);
and U1015 (N_1015,In_1085,In_682);
or U1016 (N_1016,In_1395,In_989);
and U1017 (N_1017,In_1386,In_623);
or U1018 (N_1018,In_1175,In_256);
xor U1019 (N_1019,In_649,In_1282);
nand U1020 (N_1020,In_399,In_746);
nand U1021 (N_1021,In_448,In_1332);
or U1022 (N_1022,In_1486,In_644);
or U1023 (N_1023,In_649,In_187);
or U1024 (N_1024,In_453,In_593);
nor U1025 (N_1025,In_924,In_188);
xnor U1026 (N_1026,In_517,In_1467);
nand U1027 (N_1027,In_1122,In_519);
xor U1028 (N_1028,In_68,In_456);
and U1029 (N_1029,In_283,In_629);
xor U1030 (N_1030,In_355,In_28);
or U1031 (N_1031,In_1405,In_1337);
or U1032 (N_1032,In_1157,In_922);
nor U1033 (N_1033,In_320,In_1046);
nor U1034 (N_1034,In_412,In_67);
and U1035 (N_1035,In_94,In_340);
nor U1036 (N_1036,In_906,In_168);
nand U1037 (N_1037,In_765,In_30);
nor U1038 (N_1038,In_519,In_1333);
or U1039 (N_1039,In_1315,In_112);
nor U1040 (N_1040,In_87,In_59);
nand U1041 (N_1041,In_908,In_703);
or U1042 (N_1042,In_721,In_863);
nor U1043 (N_1043,In_1385,In_326);
nor U1044 (N_1044,In_1428,In_1008);
nor U1045 (N_1045,In_82,In_1455);
or U1046 (N_1046,In_1241,In_937);
xnor U1047 (N_1047,In_1378,In_413);
nand U1048 (N_1048,In_501,In_1380);
nor U1049 (N_1049,In_1252,In_1064);
nand U1050 (N_1050,In_32,In_1207);
nand U1051 (N_1051,In_505,In_1489);
nor U1052 (N_1052,In_1156,In_545);
nor U1053 (N_1053,In_371,In_142);
xor U1054 (N_1054,In_448,In_820);
and U1055 (N_1055,In_595,In_1263);
nand U1056 (N_1056,In_774,In_376);
xor U1057 (N_1057,In_214,In_1148);
nand U1058 (N_1058,In_1103,In_1166);
and U1059 (N_1059,In_171,In_598);
or U1060 (N_1060,In_62,In_1109);
nor U1061 (N_1061,In_583,In_1375);
and U1062 (N_1062,In_1249,In_1288);
nor U1063 (N_1063,In_916,In_840);
and U1064 (N_1064,In_1493,In_1209);
nand U1065 (N_1065,In_774,In_1136);
nor U1066 (N_1066,In_1332,In_770);
or U1067 (N_1067,In_308,In_950);
nand U1068 (N_1068,In_739,In_1478);
and U1069 (N_1069,In_613,In_452);
and U1070 (N_1070,In_624,In_64);
and U1071 (N_1071,In_484,In_690);
nor U1072 (N_1072,In_28,In_935);
nor U1073 (N_1073,In_356,In_475);
nand U1074 (N_1074,In_307,In_103);
xnor U1075 (N_1075,In_941,In_119);
and U1076 (N_1076,In_642,In_1030);
nor U1077 (N_1077,In_444,In_434);
xnor U1078 (N_1078,In_7,In_349);
nor U1079 (N_1079,In_741,In_1059);
or U1080 (N_1080,In_413,In_474);
xor U1081 (N_1081,In_144,In_1358);
or U1082 (N_1082,In_1461,In_1370);
nand U1083 (N_1083,In_799,In_443);
xnor U1084 (N_1084,In_428,In_647);
nor U1085 (N_1085,In_346,In_856);
and U1086 (N_1086,In_996,In_921);
or U1087 (N_1087,In_938,In_567);
and U1088 (N_1088,In_1361,In_509);
or U1089 (N_1089,In_1140,In_804);
or U1090 (N_1090,In_665,In_1233);
xor U1091 (N_1091,In_107,In_401);
and U1092 (N_1092,In_1377,In_817);
and U1093 (N_1093,In_137,In_1111);
and U1094 (N_1094,In_740,In_1179);
and U1095 (N_1095,In_436,In_201);
xnor U1096 (N_1096,In_1080,In_474);
nor U1097 (N_1097,In_770,In_180);
and U1098 (N_1098,In_1464,In_60);
or U1099 (N_1099,In_27,In_1122);
xor U1100 (N_1100,In_939,In_715);
nor U1101 (N_1101,In_794,In_834);
and U1102 (N_1102,In_994,In_33);
nand U1103 (N_1103,In_1014,In_1097);
nand U1104 (N_1104,In_811,In_272);
nor U1105 (N_1105,In_517,In_479);
nand U1106 (N_1106,In_590,In_771);
or U1107 (N_1107,In_928,In_140);
xnor U1108 (N_1108,In_929,In_22);
xor U1109 (N_1109,In_967,In_1391);
xor U1110 (N_1110,In_1031,In_172);
nand U1111 (N_1111,In_638,In_1176);
nor U1112 (N_1112,In_435,In_653);
nor U1113 (N_1113,In_189,In_1357);
and U1114 (N_1114,In_946,In_1270);
xor U1115 (N_1115,In_1342,In_1282);
xnor U1116 (N_1116,In_573,In_1148);
nand U1117 (N_1117,In_49,In_228);
and U1118 (N_1118,In_1337,In_1386);
nor U1119 (N_1119,In_893,In_1451);
xor U1120 (N_1120,In_208,In_366);
xor U1121 (N_1121,In_931,In_1107);
and U1122 (N_1122,In_1096,In_487);
nor U1123 (N_1123,In_889,In_867);
nand U1124 (N_1124,In_778,In_428);
xor U1125 (N_1125,In_412,In_1082);
nor U1126 (N_1126,In_1046,In_912);
and U1127 (N_1127,In_64,In_385);
nor U1128 (N_1128,In_1171,In_1201);
nor U1129 (N_1129,In_468,In_712);
nor U1130 (N_1130,In_395,In_844);
and U1131 (N_1131,In_1384,In_913);
xnor U1132 (N_1132,In_735,In_1394);
xor U1133 (N_1133,In_145,In_1249);
xor U1134 (N_1134,In_1140,In_55);
or U1135 (N_1135,In_142,In_660);
nor U1136 (N_1136,In_210,In_653);
xor U1137 (N_1137,In_1389,In_1066);
or U1138 (N_1138,In_991,In_251);
nor U1139 (N_1139,In_1453,In_434);
or U1140 (N_1140,In_1325,In_1217);
and U1141 (N_1141,In_689,In_1200);
or U1142 (N_1142,In_185,In_319);
xnor U1143 (N_1143,In_751,In_275);
xor U1144 (N_1144,In_179,In_1424);
and U1145 (N_1145,In_1067,In_620);
or U1146 (N_1146,In_892,In_776);
nor U1147 (N_1147,In_1091,In_478);
or U1148 (N_1148,In_564,In_62);
nor U1149 (N_1149,In_1254,In_1013);
and U1150 (N_1150,In_1256,In_1204);
nand U1151 (N_1151,In_419,In_811);
or U1152 (N_1152,In_116,In_764);
nor U1153 (N_1153,In_188,In_1082);
nor U1154 (N_1154,In_1467,In_1439);
nor U1155 (N_1155,In_877,In_417);
nand U1156 (N_1156,In_505,In_497);
and U1157 (N_1157,In_536,In_1170);
nor U1158 (N_1158,In_1037,In_1246);
or U1159 (N_1159,In_139,In_525);
nor U1160 (N_1160,In_827,In_760);
xor U1161 (N_1161,In_1369,In_153);
and U1162 (N_1162,In_526,In_1433);
and U1163 (N_1163,In_1173,In_1099);
or U1164 (N_1164,In_959,In_664);
or U1165 (N_1165,In_444,In_355);
nand U1166 (N_1166,In_827,In_625);
or U1167 (N_1167,In_1017,In_1372);
or U1168 (N_1168,In_401,In_748);
or U1169 (N_1169,In_961,In_253);
or U1170 (N_1170,In_579,In_1011);
or U1171 (N_1171,In_127,In_380);
xnor U1172 (N_1172,In_1408,In_822);
and U1173 (N_1173,In_583,In_1263);
nor U1174 (N_1174,In_928,In_1011);
nand U1175 (N_1175,In_548,In_863);
or U1176 (N_1176,In_801,In_1299);
xnor U1177 (N_1177,In_161,In_846);
and U1178 (N_1178,In_600,In_799);
xnor U1179 (N_1179,In_1311,In_1419);
xnor U1180 (N_1180,In_389,In_991);
or U1181 (N_1181,In_462,In_756);
xor U1182 (N_1182,In_58,In_829);
nor U1183 (N_1183,In_1133,In_296);
and U1184 (N_1184,In_296,In_728);
and U1185 (N_1185,In_919,In_396);
nor U1186 (N_1186,In_1216,In_1011);
xor U1187 (N_1187,In_947,In_162);
xnor U1188 (N_1188,In_1084,In_432);
or U1189 (N_1189,In_514,In_830);
nor U1190 (N_1190,In_403,In_661);
nor U1191 (N_1191,In_1436,In_1019);
or U1192 (N_1192,In_739,In_476);
and U1193 (N_1193,In_1450,In_103);
nand U1194 (N_1194,In_369,In_225);
xnor U1195 (N_1195,In_403,In_79);
nor U1196 (N_1196,In_868,In_431);
nor U1197 (N_1197,In_492,In_467);
xor U1198 (N_1198,In_218,In_300);
nand U1199 (N_1199,In_315,In_1236);
nand U1200 (N_1200,In_625,In_269);
and U1201 (N_1201,In_1370,In_40);
nand U1202 (N_1202,In_688,In_1276);
and U1203 (N_1203,In_1421,In_805);
and U1204 (N_1204,In_1106,In_1473);
or U1205 (N_1205,In_848,In_228);
xor U1206 (N_1206,In_914,In_81);
nand U1207 (N_1207,In_10,In_381);
nor U1208 (N_1208,In_640,In_1486);
and U1209 (N_1209,In_625,In_718);
nor U1210 (N_1210,In_1348,In_522);
or U1211 (N_1211,In_118,In_1090);
nor U1212 (N_1212,In_812,In_813);
nor U1213 (N_1213,In_1265,In_248);
and U1214 (N_1214,In_397,In_0);
or U1215 (N_1215,In_906,In_814);
or U1216 (N_1216,In_230,In_746);
or U1217 (N_1217,In_1245,In_1425);
xnor U1218 (N_1218,In_1035,In_782);
and U1219 (N_1219,In_306,In_66);
xor U1220 (N_1220,In_1228,In_546);
nand U1221 (N_1221,In_336,In_1472);
xor U1222 (N_1222,In_1004,In_966);
or U1223 (N_1223,In_1069,In_799);
xnor U1224 (N_1224,In_471,In_360);
or U1225 (N_1225,In_14,In_598);
nor U1226 (N_1226,In_408,In_114);
nand U1227 (N_1227,In_1261,In_868);
xnor U1228 (N_1228,In_90,In_876);
and U1229 (N_1229,In_467,In_1301);
nand U1230 (N_1230,In_32,In_66);
nor U1231 (N_1231,In_751,In_852);
xnor U1232 (N_1232,In_1166,In_339);
nand U1233 (N_1233,In_562,In_473);
xnor U1234 (N_1234,In_1246,In_598);
and U1235 (N_1235,In_354,In_1355);
nor U1236 (N_1236,In_1094,In_404);
xor U1237 (N_1237,In_1388,In_1235);
nand U1238 (N_1238,In_1118,In_1369);
nand U1239 (N_1239,In_1136,In_1191);
or U1240 (N_1240,In_110,In_354);
and U1241 (N_1241,In_406,In_419);
or U1242 (N_1242,In_734,In_858);
nor U1243 (N_1243,In_118,In_464);
and U1244 (N_1244,In_719,In_1121);
nor U1245 (N_1245,In_937,In_1403);
nand U1246 (N_1246,In_843,In_1457);
nor U1247 (N_1247,In_54,In_253);
nor U1248 (N_1248,In_959,In_105);
xnor U1249 (N_1249,In_319,In_400);
xor U1250 (N_1250,In_680,In_898);
nor U1251 (N_1251,In_854,In_630);
nand U1252 (N_1252,In_461,In_883);
and U1253 (N_1253,In_568,In_1266);
nor U1254 (N_1254,In_609,In_188);
and U1255 (N_1255,In_926,In_1249);
nand U1256 (N_1256,In_286,In_585);
and U1257 (N_1257,In_949,In_966);
xor U1258 (N_1258,In_429,In_16);
and U1259 (N_1259,In_44,In_511);
nand U1260 (N_1260,In_202,In_823);
nand U1261 (N_1261,In_984,In_1288);
xor U1262 (N_1262,In_1361,In_1129);
nor U1263 (N_1263,In_1425,In_679);
and U1264 (N_1264,In_147,In_474);
and U1265 (N_1265,In_993,In_1310);
nand U1266 (N_1266,In_776,In_819);
xnor U1267 (N_1267,In_539,In_1008);
nand U1268 (N_1268,In_1319,In_462);
nor U1269 (N_1269,In_825,In_869);
nand U1270 (N_1270,In_496,In_719);
nand U1271 (N_1271,In_912,In_207);
nor U1272 (N_1272,In_1109,In_666);
nor U1273 (N_1273,In_1204,In_1460);
or U1274 (N_1274,In_607,In_239);
nand U1275 (N_1275,In_646,In_130);
nor U1276 (N_1276,In_761,In_218);
or U1277 (N_1277,In_111,In_932);
nor U1278 (N_1278,In_862,In_158);
xor U1279 (N_1279,In_304,In_1313);
nor U1280 (N_1280,In_1015,In_307);
or U1281 (N_1281,In_519,In_1377);
or U1282 (N_1282,In_619,In_1459);
nand U1283 (N_1283,In_690,In_182);
xor U1284 (N_1284,In_1469,In_814);
or U1285 (N_1285,In_13,In_133);
and U1286 (N_1286,In_813,In_973);
and U1287 (N_1287,In_976,In_1480);
and U1288 (N_1288,In_438,In_187);
or U1289 (N_1289,In_1496,In_73);
xnor U1290 (N_1290,In_479,In_791);
nand U1291 (N_1291,In_787,In_1482);
nor U1292 (N_1292,In_195,In_371);
or U1293 (N_1293,In_718,In_347);
or U1294 (N_1294,In_1163,In_1362);
nor U1295 (N_1295,In_269,In_475);
nor U1296 (N_1296,In_1027,In_705);
or U1297 (N_1297,In_785,In_63);
and U1298 (N_1298,In_793,In_1146);
and U1299 (N_1299,In_1281,In_1014);
and U1300 (N_1300,In_650,In_456);
nor U1301 (N_1301,In_1347,In_1075);
or U1302 (N_1302,In_375,In_1339);
nand U1303 (N_1303,In_872,In_821);
xnor U1304 (N_1304,In_1399,In_1172);
xor U1305 (N_1305,In_926,In_1322);
nor U1306 (N_1306,In_198,In_923);
nor U1307 (N_1307,In_494,In_1495);
nor U1308 (N_1308,In_599,In_1105);
nor U1309 (N_1309,In_1159,In_245);
xor U1310 (N_1310,In_1156,In_1153);
and U1311 (N_1311,In_788,In_362);
xnor U1312 (N_1312,In_1341,In_1388);
xnor U1313 (N_1313,In_1494,In_104);
nand U1314 (N_1314,In_1402,In_261);
nor U1315 (N_1315,In_611,In_1316);
or U1316 (N_1316,In_631,In_720);
xnor U1317 (N_1317,In_905,In_673);
and U1318 (N_1318,In_389,In_1241);
or U1319 (N_1319,In_329,In_629);
or U1320 (N_1320,In_581,In_574);
or U1321 (N_1321,In_595,In_373);
or U1322 (N_1322,In_1340,In_768);
xnor U1323 (N_1323,In_1310,In_124);
nand U1324 (N_1324,In_107,In_797);
or U1325 (N_1325,In_697,In_1257);
or U1326 (N_1326,In_1249,In_172);
xnor U1327 (N_1327,In_940,In_74);
or U1328 (N_1328,In_19,In_898);
or U1329 (N_1329,In_693,In_965);
nand U1330 (N_1330,In_256,In_297);
xor U1331 (N_1331,In_989,In_241);
or U1332 (N_1332,In_1392,In_432);
or U1333 (N_1333,In_306,In_206);
or U1334 (N_1334,In_1019,In_1359);
nor U1335 (N_1335,In_776,In_15);
nor U1336 (N_1336,In_1478,In_730);
xor U1337 (N_1337,In_1441,In_569);
xor U1338 (N_1338,In_629,In_124);
xor U1339 (N_1339,In_1349,In_1095);
or U1340 (N_1340,In_1474,In_269);
nand U1341 (N_1341,In_589,In_953);
nand U1342 (N_1342,In_1403,In_1368);
nor U1343 (N_1343,In_833,In_1488);
xnor U1344 (N_1344,In_873,In_1203);
nor U1345 (N_1345,In_1393,In_1291);
xnor U1346 (N_1346,In_1255,In_1289);
and U1347 (N_1347,In_137,In_1055);
or U1348 (N_1348,In_261,In_1333);
nor U1349 (N_1349,In_1226,In_409);
xor U1350 (N_1350,In_485,In_312);
nor U1351 (N_1351,In_1290,In_562);
nand U1352 (N_1352,In_272,In_1330);
nor U1353 (N_1353,In_311,In_1498);
or U1354 (N_1354,In_1428,In_516);
and U1355 (N_1355,In_310,In_870);
and U1356 (N_1356,In_719,In_181);
or U1357 (N_1357,In_451,In_453);
nand U1358 (N_1358,In_264,In_1154);
nor U1359 (N_1359,In_933,In_1202);
xnor U1360 (N_1360,In_675,In_714);
or U1361 (N_1361,In_354,In_531);
and U1362 (N_1362,In_1286,In_310);
or U1363 (N_1363,In_517,In_1156);
and U1364 (N_1364,In_661,In_685);
nand U1365 (N_1365,In_166,In_1119);
xnor U1366 (N_1366,In_1470,In_485);
or U1367 (N_1367,In_1198,In_514);
nor U1368 (N_1368,In_1162,In_368);
nor U1369 (N_1369,In_1145,In_1306);
nand U1370 (N_1370,In_970,In_1190);
xor U1371 (N_1371,In_100,In_921);
nor U1372 (N_1372,In_164,In_604);
or U1373 (N_1373,In_943,In_470);
and U1374 (N_1374,In_1499,In_252);
nor U1375 (N_1375,In_833,In_1461);
nor U1376 (N_1376,In_1378,In_661);
xnor U1377 (N_1377,In_17,In_284);
nand U1378 (N_1378,In_453,In_1315);
nand U1379 (N_1379,In_129,In_832);
and U1380 (N_1380,In_449,In_1496);
and U1381 (N_1381,In_1393,In_916);
and U1382 (N_1382,In_633,In_178);
or U1383 (N_1383,In_816,In_1483);
or U1384 (N_1384,In_1164,In_14);
nor U1385 (N_1385,In_312,In_1068);
and U1386 (N_1386,In_1108,In_392);
xor U1387 (N_1387,In_505,In_930);
nor U1388 (N_1388,In_630,In_1422);
or U1389 (N_1389,In_134,In_1003);
nand U1390 (N_1390,In_125,In_144);
or U1391 (N_1391,In_35,In_1124);
or U1392 (N_1392,In_139,In_947);
nand U1393 (N_1393,In_786,In_371);
and U1394 (N_1394,In_467,In_1465);
and U1395 (N_1395,In_1348,In_962);
xnor U1396 (N_1396,In_115,In_47);
and U1397 (N_1397,In_616,In_965);
and U1398 (N_1398,In_758,In_981);
nand U1399 (N_1399,In_1310,In_142);
nand U1400 (N_1400,In_445,In_326);
and U1401 (N_1401,In_695,In_478);
nand U1402 (N_1402,In_250,In_1493);
nor U1403 (N_1403,In_1168,In_650);
nor U1404 (N_1404,In_976,In_1017);
and U1405 (N_1405,In_934,In_788);
xnor U1406 (N_1406,In_323,In_1382);
nand U1407 (N_1407,In_184,In_24);
xnor U1408 (N_1408,In_696,In_1355);
nor U1409 (N_1409,In_96,In_1334);
nor U1410 (N_1410,In_1152,In_1134);
xor U1411 (N_1411,In_478,In_5);
or U1412 (N_1412,In_640,In_418);
nor U1413 (N_1413,In_229,In_1186);
xnor U1414 (N_1414,In_937,In_404);
nor U1415 (N_1415,In_703,In_538);
and U1416 (N_1416,In_1046,In_526);
or U1417 (N_1417,In_140,In_271);
xnor U1418 (N_1418,In_1494,In_1022);
xor U1419 (N_1419,In_858,In_770);
and U1420 (N_1420,In_911,In_1037);
xnor U1421 (N_1421,In_605,In_601);
and U1422 (N_1422,In_628,In_1021);
or U1423 (N_1423,In_1064,In_249);
and U1424 (N_1424,In_703,In_965);
nor U1425 (N_1425,In_463,In_1317);
and U1426 (N_1426,In_1353,In_511);
or U1427 (N_1427,In_1096,In_1482);
nand U1428 (N_1428,In_875,In_1490);
xor U1429 (N_1429,In_794,In_486);
xnor U1430 (N_1430,In_288,In_681);
xnor U1431 (N_1431,In_443,In_150);
and U1432 (N_1432,In_246,In_35);
xor U1433 (N_1433,In_1186,In_604);
and U1434 (N_1434,In_1489,In_1023);
nand U1435 (N_1435,In_792,In_1266);
nand U1436 (N_1436,In_808,In_1090);
or U1437 (N_1437,In_121,In_1105);
nand U1438 (N_1438,In_1315,In_619);
and U1439 (N_1439,In_776,In_674);
xor U1440 (N_1440,In_1283,In_1032);
nand U1441 (N_1441,In_1497,In_1152);
nor U1442 (N_1442,In_458,In_40);
nand U1443 (N_1443,In_1267,In_613);
or U1444 (N_1444,In_1073,In_722);
nand U1445 (N_1445,In_841,In_834);
or U1446 (N_1446,In_1335,In_1385);
nand U1447 (N_1447,In_968,In_975);
or U1448 (N_1448,In_605,In_1290);
nor U1449 (N_1449,In_745,In_726);
nor U1450 (N_1450,In_916,In_992);
nor U1451 (N_1451,In_972,In_208);
xnor U1452 (N_1452,In_668,In_340);
nor U1453 (N_1453,In_258,In_837);
and U1454 (N_1454,In_144,In_1101);
and U1455 (N_1455,In_774,In_384);
xor U1456 (N_1456,In_974,In_156);
and U1457 (N_1457,In_1233,In_882);
and U1458 (N_1458,In_120,In_1298);
and U1459 (N_1459,In_956,In_437);
xnor U1460 (N_1460,In_108,In_699);
xnor U1461 (N_1461,In_839,In_1475);
xnor U1462 (N_1462,In_1296,In_724);
xnor U1463 (N_1463,In_1312,In_925);
and U1464 (N_1464,In_632,In_996);
nor U1465 (N_1465,In_880,In_130);
nor U1466 (N_1466,In_1354,In_380);
xor U1467 (N_1467,In_39,In_571);
xor U1468 (N_1468,In_547,In_427);
and U1469 (N_1469,In_252,In_968);
and U1470 (N_1470,In_497,In_609);
nor U1471 (N_1471,In_1163,In_1196);
or U1472 (N_1472,In_771,In_18);
xor U1473 (N_1473,In_251,In_708);
nand U1474 (N_1474,In_329,In_1305);
and U1475 (N_1475,In_232,In_124);
nor U1476 (N_1476,In_989,In_839);
nor U1477 (N_1477,In_21,In_569);
nor U1478 (N_1478,In_925,In_1045);
nand U1479 (N_1479,In_1022,In_1340);
xor U1480 (N_1480,In_1062,In_1092);
or U1481 (N_1481,In_374,In_1339);
xor U1482 (N_1482,In_1080,In_1115);
xnor U1483 (N_1483,In_63,In_9);
xnor U1484 (N_1484,In_528,In_134);
and U1485 (N_1485,In_581,In_1156);
or U1486 (N_1486,In_557,In_568);
nor U1487 (N_1487,In_895,In_1426);
or U1488 (N_1488,In_1382,In_207);
nor U1489 (N_1489,In_61,In_129);
or U1490 (N_1490,In_32,In_228);
or U1491 (N_1491,In_1142,In_1484);
and U1492 (N_1492,In_250,In_1266);
or U1493 (N_1493,In_837,In_1045);
xor U1494 (N_1494,In_812,In_47);
and U1495 (N_1495,In_761,In_253);
and U1496 (N_1496,In_766,In_1473);
and U1497 (N_1497,In_362,In_459);
nand U1498 (N_1498,In_561,In_811);
or U1499 (N_1499,In_935,In_1487);
nor U1500 (N_1500,In_442,In_1130);
nand U1501 (N_1501,In_1180,In_1013);
nor U1502 (N_1502,In_375,In_227);
xnor U1503 (N_1503,In_735,In_621);
and U1504 (N_1504,In_1338,In_458);
and U1505 (N_1505,In_1099,In_1111);
or U1506 (N_1506,In_313,In_847);
xnor U1507 (N_1507,In_42,In_464);
xor U1508 (N_1508,In_88,In_774);
nand U1509 (N_1509,In_135,In_1447);
or U1510 (N_1510,In_1416,In_199);
nor U1511 (N_1511,In_1477,In_966);
nor U1512 (N_1512,In_1181,In_40);
nand U1513 (N_1513,In_614,In_900);
nand U1514 (N_1514,In_87,In_107);
nand U1515 (N_1515,In_320,In_1437);
and U1516 (N_1516,In_1226,In_423);
or U1517 (N_1517,In_1174,In_543);
nor U1518 (N_1518,In_1065,In_7);
nand U1519 (N_1519,In_960,In_300);
xor U1520 (N_1520,In_579,In_955);
or U1521 (N_1521,In_1026,In_271);
nor U1522 (N_1522,In_1358,In_145);
nand U1523 (N_1523,In_1102,In_1086);
nand U1524 (N_1524,In_1268,In_1385);
nand U1525 (N_1525,In_1328,In_1239);
and U1526 (N_1526,In_52,In_259);
xor U1527 (N_1527,In_1367,In_1250);
xnor U1528 (N_1528,In_1317,In_77);
and U1529 (N_1529,In_546,In_853);
nand U1530 (N_1530,In_1236,In_1033);
nand U1531 (N_1531,In_192,In_985);
nand U1532 (N_1532,In_622,In_647);
xor U1533 (N_1533,In_737,In_910);
nor U1534 (N_1534,In_985,In_515);
nor U1535 (N_1535,In_987,In_1042);
nor U1536 (N_1536,In_845,In_678);
nand U1537 (N_1537,In_432,In_203);
nor U1538 (N_1538,In_653,In_1027);
nor U1539 (N_1539,In_1371,In_1399);
nand U1540 (N_1540,In_923,In_250);
and U1541 (N_1541,In_963,In_1313);
xor U1542 (N_1542,In_78,In_138);
xnor U1543 (N_1543,In_928,In_1492);
nor U1544 (N_1544,In_467,In_1277);
nor U1545 (N_1545,In_944,In_1094);
and U1546 (N_1546,In_379,In_524);
and U1547 (N_1547,In_838,In_1160);
or U1548 (N_1548,In_1141,In_854);
or U1549 (N_1549,In_832,In_535);
and U1550 (N_1550,In_1477,In_450);
and U1551 (N_1551,In_341,In_1186);
nand U1552 (N_1552,In_23,In_1388);
nand U1553 (N_1553,In_125,In_525);
xnor U1554 (N_1554,In_116,In_379);
xor U1555 (N_1555,In_491,In_487);
nand U1556 (N_1556,In_462,In_353);
or U1557 (N_1557,In_1328,In_215);
nor U1558 (N_1558,In_146,In_1336);
or U1559 (N_1559,In_1273,In_501);
or U1560 (N_1560,In_254,In_266);
and U1561 (N_1561,In_275,In_1329);
and U1562 (N_1562,In_1309,In_548);
nor U1563 (N_1563,In_1489,In_843);
nand U1564 (N_1564,In_1257,In_89);
or U1565 (N_1565,In_594,In_943);
and U1566 (N_1566,In_1412,In_412);
and U1567 (N_1567,In_1055,In_431);
nand U1568 (N_1568,In_527,In_1305);
nor U1569 (N_1569,In_94,In_1222);
nor U1570 (N_1570,In_953,In_322);
or U1571 (N_1571,In_1270,In_952);
and U1572 (N_1572,In_1476,In_1428);
xnor U1573 (N_1573,In_465,In_1129);
or U1574 (N_1574,In_1286,In_1045);
xor U1575 (N_1575,In_1387,In_293);
xor U1576 (N_1576,In_652,In_1294);
xor U1577 (N_1577,In_328,In_142);
nand U1578 (N_1578,In_1226,In_235);
xnor U1579 (N_1579,In_617,In_655);
nand U1580 (N_1580,In_554,In_613);
and U1581 (N_1581,In_952,In_948);
and U1582 (N_1582,In_1242,In_1364);
or U1583 (N_1583,In_329,In_909);
or U1584 (N_1584,In_414,In_1067);
nand U1585 (N_1585,In_1466,In_1413);
nand U1586 (N_1586,In_72,In_1093);
or U1587 (N_1587,In_1285,In_924);
nor U1588 (N_1588,In_571,In_394);
nand U1589 (N_1589,In_1132,In_69);
and U1590 (N_1590,In_663,In_32);
xnor U1591 (N_1591,In_230,In_365);
nand U1592 (N_1592,In_1270,In_227);
nor U1593 (N_1593,In_1030,In_484);
xor U1594 (N_1594,In_419,In_1292);
nand U1595 (N_1595,In_913,In_1495);
and U1596 (N_1596,In_1071,In_1456);
or U1597 (N_1597,In_1269,In_1435);
xor U1598 (N_1598,In_760,In_1482);
nor U1599 (N_1599,In_450,In_254);
xnor U1600 (N_1600,In_1488,In_1392);
xor U1601 (N_1601,In_84,In_1467);
xnor U1602 (N_1602,In_890,In_640);
nor U1603 (N_1603,In_616,In_1486);
or U1604 (N_1604,In_789,In_1207);
nor U1605 (N_1605,In_1106,In_495);
nor U1606 (N_1606,In_372,In_1122);
and U1607 (N_1607,In_484,In_194);
or U1608 (N_1608,In_1203,In_1445);
xor U1609 (N_1609,In_808,In_1246);
or U1610 (N_1610,In_217,In_307);
xnor U1611 (N_1611,In_136,In_62);
nand U1612 (N_1612,In_529,In_545);
or U1613 (N_1613,In_584,In_789);
and U1614 (N_1614,In_86,In_1282);
nor U1615 (N_1615,In_87,In_193);
and U1616 (N_1616,In_221,In_934);
and U1617 (N_1617,In_1468,In_65);
nor U1618 (N_1618,In_210,In_1203);
and U1619 (N_1619,In_31,In_71);
nand U1620 (N_1620,In_1439,In_1383);
nand U1621 (N_1621,In_1201,In_189);
and U1622 (N_1622,In_563,In_997);
or U1623 (N_1623,In_165,In_1371);
nor U1624 (N_1624,In_111,In_1346);
nand U1625 (N_1625,In_155,In_312);
nand U1626 (N_1626,In_581,In_336);
or U1627 (N_1627,In_1032,In_43);
or U1628 (N_1628,In_1067,In_587);
xor U1629 (N_1629,In_75,In_1307);
nand U1630 (N_1630,In_99,In_989);
nor U1631 (N_1631,In_493,In_1382);
nand U1632 (N_1632,In_413,In_351);
or U1633 (N_1633,In_237,In_1356);
xor U1634 (N_1634,In_174,In_503);
nand U1635 (N_1635,In_844,In_710);
xor U1636 (N_1636,In_817,In_1015);
nand U1637 (N_1637,In_1208,In_288);
xnor U1638 (N_1638,In_190,In_209);
nor U1639 (N_1639,In_699,In_1012);
xnor U1640 (N_1640,In_441,In_1141);
nand U1641 (N_1641,In_1419,In_524);
nand U1642 (N_1642,In_679,In_1472);
xor U1643 (N_1643,In_241,In_1437);
nand U1644 (N_1644,In_251,In_1014);
xor U1645 (N_1645,In_140,In_317);
nand U1646 (N_1646,In_1460,In_356);
or U1647 (N_1647,In_1389,In_390);
nand U1648 (N_1648,In_1395,In_353);
nor U1649 (N_1649,In_815,In_399);
and U1650 (N_1650,In_721,In_1403);
nand U1651 (N_1651,In_852,In_1210);
and U1652 (N_1652,In_318,In_819);
nor U1653 (N_1653,In_91,In_730);
and U1654 (N_1654,In_399,In_968);
or U1655 (N_1655,In_1351,In_1202);
or U1656 (N_1656,In_1128,In_124);
and U1657 (N_1657,In_381,In_77);
nand U1658 (N_1658,In_275,In_1379);
or U1659 (N_1659,In_110,In_1441);
or U1660 (N_1660,In_942,In_343);
and U1661 (N_1661,In_562,In_715);
or U1662 (N_1662,In_245,In_394);
and U1663 (N_1663,In_526,In_84);
xor U1664 (N_1664,In_78,In_524);
nand U1665 (N_1665,In_321,In_1149);
nand U1666 (N_1666,In_355,In_609);
or U1667 (N_1667,In_90,In_865);
or U1668 (N_1668,In_1427,In_1311);
xnor U1669 (N_1669,In_1193,In_1098);
and U1670 (N_1670,In_1288,In_936);
or U1671 (N_1671,In_854,In_1432);
nand U1672 (N_1672,In_666,In_507);
nand U1673 (N_1673,In_215,In_465);
nand U1674 (N_1674,In_210,In_682);
and U1675 (N_1675,In_471,In_591);
nand U1676 (N_1676,In_245,In_1129);
xor U1677 (N_1677,In_1322,In_629);
nand U1678 (N_1678,In_1419,In_1021);
nand U1679 (N_1679,In_120,In_293);
nor U1680 (N_1680,In_1339,In_897);
or U1681 (N_1681,In_363,In_1059);
and U1682 (N_1682,In_152,In_939);
nor U1683 (N_1683,In_511,In_1189);
and U1684 (N_1684,In_261,In_425);
nand U1685 (N_1685,In_1125,In_473);
nor U1686 (N_1686,In_939,In_1223);
xnor U1687 (N_1687,In_350,In_139);
nand U1688 (N_1688,In_635,In_334);
or U1689 (N_1689,In_1416,In_66);
nor U1690 (N_1690,In_1329,In_797);
nor U1691 (N_1691,In_263,In_124);
and U1692 (N_1692,In_797,In_865);
and U1693 (N_1693,In_414,In_874);
nand U1694 (N_1694,In_83,In_1382);
nor U1695 (N_1695,In_1130,In_463);
or U1696 (N_1696,In_209,In_1401);
nor U1697 (N_1697,In_1356,In_683);
or U1698 (N_1698,In_1415,In_1217);
or U1699 (N_1699,In_62,In_297);
and U1700 (N_1700,In_1351,In_978);
nor U1701 (N_1701,In_1299,In_371);
xor U1702 (N_1702,In_663,In_1463);
or U1703 (N_1703,In_1466,In_972);
nor U1704 (N_1704,In_594,In_1302);
nor U1705 (N_1705,In_38,In_823);
nor U1706 (N_1706,In_1273,In_1163);
nand U1707 (N_1707,In_1004,In_1049);
nand U1708 (N_1708,In_728,In_994);
and U1709 (N_1709,In_1257,In_33);
xnor U1710 (N_1710,In_1386,In_1429);
nor U1711 (N_1711,In_288,In_147);
xor U1712 (N_1712,In_714,In_73);
and U1713 (N_1713,In_1281,In_246);
nand U1714 (N_1714,In_1073,In_585);
nor U1715 (N_1715,In_1074,In_401);
nand U1716 (N_1716,In_982,In_1139);
nand U1717 (N_1717,In_951,In_1457);
nor U1718 (N_1718,In_1239,In_1479);
or U1719 (N_1719,In_1351,In_977);
nand U1720 (N_1720,In_1466,In_1196);
nor U1721 (N_1721,In_857,In_620);
and U1722 (N_1722,In_60,In_849);
and U1723 (N_1723,In_1437,In_896);
nor U1724 (N_1724,In_800,In_551);
or U1725 (N_1725,In_322,In_283);
nand U1726 (N_1726,In_992,In_125);
nand U1727 (N_1727,In_807,In_937);
nand U1728 (N_1728,In_251,In_144);
and U1729 (N_1729,In_777,In_362);
nand U1730 (N_1730,In_180,In_1013);
xor U1731 (N_1731,In_172,In_545);
xnor U1732 (N_1732,In_179,In_621);
and U1733 (N_1733,In_516,In_1357);
nor U1734 (N_1734,In_1290,In_570);
xnor U1735 (N_1735,In_1317,In_473);
nor U1736 (N_1736,In_475,In_350);
or U1737 (N_1737,In_691,In_961);
nor U1738 (N_1738,In_1251,In_733);
nor U1739 (N_1739,In_403,In_1391);
and U1740 (N_1740,In_790,In_1346);
and U1741 (N_1741,In_951,In_1107);
xor U1742 (N_1742,In_216,In_853);
nand U1743 (N_1743,In_1278,In_798);
or U1744 (N_1744,In_361,In_559);
and U1745 (N_1745,In_1056,In_949);
or U1746 (N_1746,In_993,In_211);
nor U1747 (N_1747,In_421,In_555);
xnor U1748 (N_1748,In_988,In_468);
or U1749 (N_1749,In_1166,In_390);
or U1750 (N_1750,In_769,In_1351);
and U1751 (N_1751,In_590,In_356);
nor U1752 (N_1752,In_308,In_1167);
or U1753 (N_1753,In_164,In_314);
or U1754 (N_1754,In_1227,In_856);
or U1755 (N_1755,In_405,In_264);
or U1756 (N_1756,In_441,In_495);
or U1757 (N_1757,In_194,In_1358);
and U1758 (N_1758,In_591,In_1038);
and U1759 (N_1759,In_1190,In_1308);
and U1760 (N_1760,In_662,In_593);
nand U1761 (N_1761,In_1064,In_460);
nor U1762 (N_1762,In_583,In_718);
or U1763 (N_1763,In_467,In_1116);
nor U1764 (N_1764,In_934,In_986);
nor U1765 (N_1765,In_559,In_360);
nand U1766 (N_1766,In_42,In_155);
xnor U1767 (N_1767,In_689,In_1294);
xnor U1768 (N_1768,In_762,In_203);
and U1769 (N_1769,In_57,In_714);
xnor U1770 (N_1770,In_1304,In_140);
or U1771 (N_1771,In_815,In_28);
nand U1772 (N_1772,In_1333,In_491);
or U1773 (N_1773,In_1273,In_942);
or U1774 (N_1774,In_1300,In_508);
xnor U1775 (N_1775,In_1361,In_156);
nand U1776 (N_1776,In_1450,In_113);
or U1777 (N_1777,In_1479,In_699);
nor U1778 (N_1778,In_833,In_267);
nor U1779 (N_1779,In_512,In_509);
nor U1780 (N_1780,In_788,In_277);
xnor U1781 (N_1781,In_1043,In_349);
nor U1782 (N_1782,In_842,In_415);
nand U1783 (N_1783,In_1058,In_1431);
nor U1784 (N_1784,In_272,In_1173);
xor U1785 (N_1785,In_916,In_1259);
xor U1786 (N_1786,In_423,In_574);
nor U1787 (N_1787,In_1254,In_1175);
and U1788 (N_1788,In_726,In_331);
and U1789 (N_1789,In_73,In_1277);
nand U1790 (N_1790,In_102,In_321);
xor U1791 (N_1791,In_1239,In_437);
or U1792 (N_1792,In_918,In_496);
and U1793 (N_1793,In_1345,In_324);
and U1794 (N_1794,In_762,In_1393);
xnor U1795 (N_1795,In_759,In_279);
and U1796 (N_1796,In_964,In_53);
and U1797 (N_1797,In_956,In_1408);
xnor U1798 (N_1798,In_1449,In_1095);
and U1799 (N_1799,In_835,In_53);
nand U1800 (N_1800,In_306,In_98);
nor U1801 (N_1801,In_363,In_757);
and U1802 (N_1802,In_1491,In_924);
and U1803 (N_1803,In_908,In_409);
nand U1804 (N_1804,In_1204,In_930);
xnor U1805 (N_1805,In_1358,In_1413);
nand U1806 (N_1806,In_617,In_315);
or U1807 (N_1807,In_756,In_218);
or U1808 (N_1808,In_939,In_411);
and U1809 (N_1809,In_1205,In_295);
xor U1810 (N_1810,In_978,In_1229);
nand U1811 (N_1811,In_33,In_1015);
xor U1812 (N_1812,In_1234,In_1473);
nand U1813 (N_1813,In_882,In_69);
and U1814 (N_1814,In_521,In_186);
and U1815 (N_1815,In_1012,In_176);
and U1816 (N_1816,In_170,In_1464);
or U1817 (N_1817,In_973,In_814);
xnor U1818 (N_1818,In_862,In_1334);
nand U1819 (N_1819,In_110,In_1317);
or U1820 (N_1820,In_515,In_519);
and U1821 (N_1821,In_1161,In_1202);
nand U1822 (N_1822,In_22,In_859);
nor U1823 (N_1823,In_1421,In_234);
xor U1824 (N_1824,In_770,In_343);
xnor U1825 (N_1825,In_518,In_33);
nor U1826 (N_1826,In_1126,In_1211);
and U1827 (N_1827,In_701,In_617);
and U1828 (N_1828,In_247,In_935);
nand U1829 (N_1829,In_609,In_425);
nand U1830 (N_1830,In_1275,In_856);
nor U1831 (N_1831,In_1173,In_1431);
or U1832 (N_1832,In_1314,In_1235);
or U1833 (N_1833,In_269,In_387);
and U1834 (N_1834,In_114,In_1025);
and U1835 (N_1835,In_356,In_1219);
and U1836 (N_1836,In_794,In_1176);
nand U1837 (N_1837,In_235,In_281);
nor U1838 (N_1838,In_1071,In_1272);
or U1839 (N_1839,In_1077,In_1148);
xnor U1840 (N_1840,In_1327,In_1447);
xor U1841 (N_1841,In_1169,In_58);
nor U1842 (N_1842,In_1476,In_507);
xor U1843 (N_1843,In_1184,In_727);
xor U1844 (N_1844,In_157,In_1484);
xnor U1845 (N_1845,In_218,In_1039);
nand U1846 (N_1846,In_37,In_172);
or U1847 (N_1847,In_1468,In_1289);
xor U1848 (N_1848,In_1489,In_507);
nand U1849 (N_1849,In_715,In_137);
xnor U1850 (N_1850,In_1075,In_284);
nor U1851 (N_1851,In_433,In_588);
nor U1852 (N_1852,In_15,In_1021);
nand U1853 (N_1853,In_192,In_1491);
nor U1854 (N_1854,In_708,In_1230);
and U1855 (N_1855,In_1112,In_922);
xor U1856 (N_1856,In_640,In_1181);
xnor U1857 (N_1857,In_301,In_1499);
xnor U1858 (N_1858,In_1134,In_1014);
nor U1859 (N_1859,In_820,In_752);
nor U1860 (N_1860,In_1291,In_694);
nor U1861 (N_1861,In_1317,In_1103);
nor U1862 (N_1862,In_410,In_414);
or U1863 (N_1863,In_133,In_650);
or U1864 (N_1864,In_619,In_1418);
or U1865 (N_1865,In_723,In_681);
nor U1866 (N_1866,In_642,In_1401);
and U1867 (N_1867,In_65,In_1493);
or U1868 (N_1868,In_229,In_357);
xor U1869 (N_1869,In_1215,In_439);
and U1870 (N_1870,In_293,In_804);
xor U1871 (N_1871,In_667,In_1117);
nand U1872 (N_1872,In_189,In_673);
nand U1873 (N_1873,In_660,In_262);
nor U1874 (N_1874,In_599,In_537);
xor U1875 (N_1875,In_1064,In_1066);
nor U1876 (N_1876,In_535,In_1355);
nor U1877 (N_1877,In_1361,In_862);
xor U1878 (N_1878,In_1121,In_1158);
nand U1879 (N_1879,In_212,In_701);
nor U1880 (N_1880,In_903,In_1161);
xnor U1881 (N_1881,In_322,In_612);
nor U1882 (N_1882,In_71,In_1407);
xnor U1883 (N_1883,In_1201,In_623);
nor U1884 (N_1884,In_941,In_959);
xnor U1885 (N_1885,In_341,In_42);
xnor U1886 (N_1886,In_1385,In_1017);
xnor U1887 (N_1887,In_1193,In_420);
or U1888 (N_1888,In_448,In_475);
xor U1889 (N_1889,In_92,In_151);
nor U1890 (N_1890,In_680,In_304);
nand U1891 (N_1891,In_292,In_61);
xor U1892 (N_1892,In_1355,In_1383);
or U1893 (N_1893,In_1489,In_36);
xnor U1894 (N_1894,In_961,In_59);
nor U1895 (N_1895,In_546,In_375);
nand U1896 (N_1896,In_379,In_390);
nor U1897 (N_1897,In_1089,In_160);
xor U1898 (N_1898,In_136,In_1036);
xnor U1899 (N_1899,In_1206,In_1024);
and U1900 (N_1900,In_55,In_719);
xor U1901 (N_1901,In_37,In_1326);
or U1902 (N_1902,In_1168,In_377);
and U1903 (N_1903,In_1444,In_1327);
or U1904 (N_1904,In_109,In_504);
nand U1905 (N_1905,In_31,In_149);
nand U1906 (N_1906,In_696,In_824);
xor U1907 (N_1907,In_145,In_1010);
nor U1908 (N_1908,In_72,In_1371);
nand U1909 (N_1909,In_1306,In_245);
nand U1910 (N_1910,In_1356,In_698);
nor U1911 (N_1911,In_1298,In_974);
xor U1912 (N_1912,In_670,In_703);
nand U1913 (N_1913,In_503,In_604);
nor U1914 (N_1914,In_1144,In_1057);
or U1915 (N_1915,In_41,In_1398);
nand U1916 (N_1916,In_195,In_931);
xor U1917 (N_1917,In_819,In_316);
nor U1918 (N_1918,In_11,In_1212);
nor U1919 (N_1919,In_1309,In_479);
and U1920 (N_1920,In_108,In_1156);
xnor U1921 (N_1921,In_142,In_835);
nor U1922 (N_1922,In_280,In_181);
nor U1923 (N_1923,In_555,In_132);
or U1924 (N_1924,In_2,In_1245);
nor U1925 (N_1925,In_562,In_1164);
nor U1926 (N_1926,In_1020,In_783);
xnor U1927 (N_1927,In_1488,In_1321);
nor U1928 (N_1928,In_1278,In_767);
nor U1929 (N_1929,In_1416,In_834);
or U1930 (N_1930,In_1123,In_1495);
and U1931 (N_1931,In_1220,In_808);
nand U1932 (N_1932,In_241,In_1227);
and U1933 (N_1933,In_1085,In_122);
nand U1934 (N_1934,In_445,In_1350);
and U1935 (N_1935,In_998,In_19);
and U1936 (N_1936,In_984,In_1075);
xor U1937 (N_1937,In_432,In_1250);
nand U1938 (N_1938,In_1249,In_1179);
nor U1939 (N_1939,In_1296,In_494);
and U1940 (N_1940,In_1486,In_993);
nand U1941 (N_1941,In_954,In_261);
nand U1942 (N_1942,In_1066,In_657);
and U1943 (N_1943,In_244,In_980);
nand U1944 (N_1944,In_578,In_125);
and U1945 (N_1945,In_123,In_1263);
or U1946 (N_1946,In_1408,In_381);
and U1947 (N_1947,In_1420,In_335);
or U1948 (N_1948,In_616,In_111);
nor U1949 (N_1949,In_1009,In_1184);
nand U1950 (N_1950,In_681,In_1356);
nor U1951 (N_1951,In_1255,In_126);
xnor U1952 (N_1952,In_1317,In_1426);
nand U1953 (N_1953,In_1236,In_973);
xor U1954 (N_1954,In_583,In_683);
and U1955 (N_1955,In_1435,In_269);
nand U1956 (N_1956,In_1491,In_776);
and U1957 (N_1957,In_932,In_1359);
and U1958 (N_1958,In_690,In_184);
nor U1959 (N_1959,In_1125,In_810);
xnor U1960 (N_1960,In_135,In_39);
nor U1961 (N_1961,In_1,In_1470);
nor U1962 (N_1962,In_46,In_706);
or U1963 (N_1963,In_334,In_1427);
xor U1964 (N_1964,In_400,In_611);
xor U1965 (N_1965,In_997,In_976);
nor U1966 (N_1966,In_1017,In_553);
and U1967 (N_1967,In_632,In_1077);
or U1968 (N_1968,In_843,In_131);
or U1969 (N_1969,In_312,In_1072);
and U1970 (N_1970,In_502,In_1466);
or U1971 (N_1971,In_986,In_741);
or U1972 (N_1972,In_1155,In_276);
nor U1973 (N_1973,In_912,In_1180);
and U1974 (N_1974,In_1221,In_185);
or U1975 (N_1975,In_1388,In_708);
nor U1976 (N_1976,In_955,In_704);
nand U1977 (N_1977,In_1186,In_739);
xor U1978 (N_1978,In_369,In_635);
xnor U1979 (N_1979,In_1314,In_1334);
nand U1980 (N_1980,In_1317,In_105);
nand U1981 (N_1981,In_27,In_1019);
and U1982 (N_1982,In_1443,In_1444);
nand U1983 (N_1983,In_3,In_240);
nand U1984 (N_1984,In_597,In_776);
xnor U1985 (N_1985,In_344,In_672);
xnor U1986 (N_1986,In_1095,In_844);
or U1987 (N_1987,In_1273,In_988);
nand U1988 (N_1988,In_643,In_883);
or U1989 (N_1989,In_548,In_76);
nor U1990 (N_1990,In_94,In_247);
or U1991 (N_1991,In_780,In_585);
nor U1992 (N_1992,In_638,In_300);
nand U1993 (N_1993,In_274,In_525);
xnor U1994 (N_1994,In_122,In_822);
or U1995 (N_1995,In_540,In_826);
nor U1996 (N_1996,In_507,In_1340);
nand U1997 (N_1997,In_1230,In_886);
nor U1998 (N_1998,In_388,In_1324);
and U1999 (N_1999,In_155,In_720);
xor U2000 (N_2000,In_513,In_811);
nand U2001 (N_2001,In_765,In_986);
or U2002 (N_2002,In_1472,In_1352);
xnor U2003 (N_2003,In_1053,In_389);
and U2004 (N_2004,In_33,In_202);
and U2005 (N_2005,In_750,In_438);
xor U2006 (N_2006,In_715,In_178);
and U2007 (N_2007,In_1345,In_647);
and U2008 (N_2008,In_721,In_932);
or U2009 (N_2009,In_699,In_1060);
nand U2010 (N_2010,In_1316,In_507);
nand U2011 (N_2011,In_957,In_461);
nor U2012 (N_2012,In_102,In_482);
nor U2013 (N_2013,In_107,In_530);
xor U2014 (N_2014,In_1141,In_1169);
nor U2015 (N_2015,In_904,In_754);
nor U2016 (N_2016,In_551,In_594);
nor U2017 (N_2017,In_819,In_186);
xnor U2018 (N_2018,In_1432,In_683);
xor U2019 (N_2019,In_254,In_1251);
xor U2020 (N_2020,In_1257,In_135);
and U2021 (N_2021,In_1372,In_1429);
and U2022 (N_2022,In_1159,In_1311);
nor U2023 (N_2023,In_1332,In_401);
xor U2024 (N_2024,In_1262,In_716);
or U2025 (N_2025,In_1463,In_1282);
nand U2026 (N_2026,In_307,In_696);
xnor U2027 (N_2027,In_727,In_186);
nand U2028 (N_2028,In_534,In_1381);
or U2029 (N_2029,In_963,In_1005);
xnor U2030 (N_2030,In_1075,In_455);
or U2031 (N_2031,In_1183,In_97);
or U2032 (N_2032,In_104,In_863);
nor U2033 (N_2033,In_1316,In_888);
nor U2034 (N_2034,In_379,In_529);
or U2035 (N_2035,In_1018,In_1262);
or U2036 (N_2036,In_492,In_1322);
nand U2037 (N_2037,In_712,In_905);
nor U2038 (N_2038,In_1221,In_928);
and U2039 (N_2039,In_1169,In_1330);
or U2040 (N_2040,In_156,In_169);
xnor U2041 (N_2041,In_1453,In_1001);
nor U2042 (N_2042,In_1374,In_145);
nand U2043 (N_2043,In_30,In_147);
or U2044 (N_2044,In_93,In_1226);
nand U2045 (N_2045,In_38,In_808);
or U2046 (N_2046,In_769,In_42);
nor U2047 (N_2047,In_54,In_1164);
xor U2048 (N_2048,In_374,In_487);
xor U2049 (N_2049,In_1054,In_344);
nor U2050 (N_2050,In_1494,In_1223);
nand U2051 (N_2051,In_1036,In_1440);
nor U2052 (N_2052,In_19,In_152);
nand U2053 (N_2053,In_1170,In_507);
xor U2054 (N_2054,In_1116,In_1220);
nor U2055 (N_2055,In_780,In_320);
nor U2056 (N_2056,In_1430,In_721);
nor U2057 (N_2057,In_1167,In_454);
and U2058 (N_2058,In_626,In_714);
xor U2059 (N_2059,In_138,In_385);
xnor U2060 (N_2060,In_289,In_22);
and U2061 (N_2061,In_1404,In_398);
nand U2062 (N_2062,In_1355,In_1366);
nand U2063 (N_2063,In_114,In_21);
or U2064 (N_2064,In_719,In_880);
nand U2065 (N_2065,In_1111,In_965);
and U2066 (N_2066,In_900,In_1467);
nand U2067 (N_2067,In_56,In_169);
xnor U2068 (N_2068,In_1494,In_854);
or U2069 (N_2069,In_57,In_554);
and U2070 (N_2070,In_1431,In_364);
nand U2071 (N_2071,In_1214,In_627);
xnor U2072 (N_2072,In_1069,In_483);
xnor U2073 (N_2073,In_1327,In_1483);
nor U2074 (N_2074,In_208,In_918);
and U2075 (N_2075,In_1084,In_1414);
nand U2076 (N_2076,In_740,In_302);
or U2077 (N_2077,In_1038,In_276);
or U2078 (N_2078,In_1383,In_1478);
nor U2079 (N_2079,In_655,In_753);
and U2080 (N_2080,In_1325,In_785);
nor U2081 (N_2081,In_609,In_316);
nand U2082 (N_2082,In_621,In_317);
nor U2083 (N_2083,In_131,In_425);
nand U2084 (N_2084,In_436,In_1019);
or U2085 (N_2085,In_1129,In_1005);
xor U2086 (N_2086,In_832,In_1421);
nand U2087 (N_2087,In_800,In_600);
nor U2088 (N_2088,In_909,In_1338);
nor U2089 (N_2089,In_1264,In_1350);
nor U2090 (N_2090,In_1399,In_101);
xnor U2091 (N_2091,In_820,In_414);
and U2092 (N_2092,In_445,In_890);
xor U2093 (N_2093,In_1264,In_944);
or U2094 (N_2094,In_437,In_601);
xnor U2095 (N_2095,In_1390,In_590);
nor U2096 (N_2096,In_988,In_36);
and U2097 (N_2097,In_786,In_1049);
and U2098 (N_2098,In_1104,In_1398);
or U2099 (N_2099,In_530,In_210);
or U2100 (N_2100,In_477,In_1297);
nor U2101 (N_2101,In_1302,In_910);
nor U2102 (N_2102,In_741,In_688);
nand U2103 (N_2103,In_749,In_20);
nand U2104 (N_2104,In_1284,In_1147);
and U2105 (N_2105,In_588,In_311);
xor U2106 (N_2106,In_923,In_1062);
nand U2107 (N_2107,In_34,In_1281);
nand U2108 (N_2108,In_716,In_121);
and U2109 (N_2109,In_1306,In_747);
or U2110 (N_2110,In_831,In_310);
nor U2111 (N_2111,In_872,In_47);
or U2112 (N_2112,In_766,In_1236);
nand U2113 (N_2113,In_1126,In_561);
or U2114 (N_2114,In_1213,In_184);
or U2115 (N_2115,In_249,In_515);
or U2116 (N_2116,In_418,In_1322);
xnor U2117 (N_2117,In_264,In_1331);
and U2118 (N_2118,In_412,In_723);
or U2119 (N_2119,In_443,In_1099);
nand U2120 (N_2120,In_1079,In_264);
or U2121 (N_2121,In_516,In_590);
nor U2122 (N_2122,In_404,In_1404);
nand U2123 (N_2123,In_797,In_362);
and U2124 (N_2124,In_1421,In_713);
nor U2125 (N_2125,In_166,In_102);
or U2126 (N_2126,In_1331,In_638);
or U2127 (N_2127,In_879,In_1135);
xnor U2128 (N_2128,In_1348,In_1415);
or U2129 (N_2129,In_1384,In_1304);
xor U2130 (N_2130,In_1446,In_1363);
xor U2131 (N_2131,In_1400,In_726);
or U2132 (N_2132,In_631,In_784);
nand U2133 (N_2133,In_757,In_1382);
nand U2134 (N_2134,In_391,In_1286);
and U2135 (N_2135,In_440,In_949);
and U2136 (N_2136,In_291,In_369);
xor U2137 (N_2137,In_1341,In_178);
nand U2138 (N_2138,In_325,In_1270);
nor U2139 (N_2139,In_526,In_157);
xor U2140 (N_2140,In_1045,In_343);
nand U2141 (N_2141,In_242,In_1033);
nand U2142 (N_2142,In_1122,In_891);
or U2143 (N_2143,In_267,In_496);
and U2144 (N_2144,In_1001,In_362);
and U2145 (N_2145,In_668,In_1194);
or U2146 (N_2146,In_78,In_803);
nand U2147 (N_2147,In_581,In_1223);
xor U2148 (N_2148,In_743,In_993);
or U2149 (N_2149,In_229,In_375);
nand U2150 (N_2150,In_297,In_1146);
xnor U2151 (N_2151,In_1135,In_874);
and U2152 (N_2152,In_951,In_870);
nand U2153 (N_2153,In_1329,In_1155);
nand U2154 (N_2154,In_658,In_813);
or U2155 (N_2155,In_367,In_600);
nor U2156 (N_2156,In_854,In_739);
nand U2157 (N_2157,In_252,In_934);
or U2158 (N_2158,In_112,In_167);
xor U2159 (N_2159,In_277,In_489);
nand U2160 (N_2160,In_1118,In_485);
and U2161 (N_2161,In_1042,In_116);
or U2162 (N_2162,In_393,In_659);
nor U2163 (N_2163,In_316,In_1485);
nor U2164 (N_2164,In_1095,In_1480);
and U2165 (N_2165,In_1442,In_1208);
xnor U2166 (N_2166,In_52,In_590);
or U2167 (N_2167,In_1049,In_417);
nand U2168 (N_2168,In_445,In_976);
or U2169 (N_2169,In_606,In_63);
and U2170 (N_2170,In_1005,In_13);
or U2171 (N_2171,In_632,In_1108);
nor U2172 (N_2172,In_975,In_696);
nor U2173 (N_2173,In_1495,In_329);
and U2174 (N_2174,In_1012,In_407);
or U2175 (N_2175,In_838,In_596);
nand U2176 (N_2176,In_795,In_1383);
and U2177 (N_2177,In_433,In_323);
nor U2178 (N_2178,In_477,In_1404);
nor U2179 (N_2179,In_1130,In_501);
nand U2180 (N_2180,In_925,In_725);
nor U2181 (N_2181,In_1411,In_900);
or U2182 (N_2182,In_105,In_174);
xor U2183 (N_2183,In_664,In_137);
and U2184 (N_2184,In_710,In_1376);
xor U2185 (N_2185,In_200,In_735);
nor U2186 (N_2186,In_277,In_328);
nor U2187 (N_2187,In_94,In_933);
nor U2188 (N_2188,In_1273,In_175);
and U2189 (N_2189,In_556,In_1130);
nand U2190 (N_2190,In_1085,In_807);
nand U2191 (N_2191,In_1240,In_654);
xor U2192 (N_2192,In_340,In_34);
and U2193 (N_2193,In_1447,In_534);
nor U2194 (N_2194,In_471,In_1087);
or U2195 (N_2195,In_971,In_1081);
xnor U2196 (N_2196,In_1156,In_729);
nor U2197 (N_2197,In_802,In_17);
and U2198 (N_2198,In_491,In_1115);
xnor U2199 (N_2199,In_761,In_561);
or U2200 (N_2200,In_949,In_970);
and U2201 (N_2201,In_790,In_347);
or U2202 (N_2202,In_349,In_568);
xor U2203 (N_2203,In_425,In_1215);
nor U2204 (N_2204,In_275,In_822);
xnor U2205 (N_2205,In_40,In_474);
xor U2206 (N_2206,In_703,In_117);
nor U2207 (N_2207,In_1205,In_1473);
or U2208 (N_2208,In_785,In_694);
and U2209 (N_2209,In_1010,In_47);
and U2210 (N_2210,In_971,In_201);
and U2211 (N_2211,In_0,In_1259);
xnor U2212 (N_2212,In_484,In_522);
or U2213 (N_2213,In_1150,In_726);
nor U2214 (N_2214,In_1496,In_332);
nand U2215 (N_2215,In_996,In_242);
or U2216 (N_2216,In_255,In_790);
and U2217 (N_2217,In_608,In_358);
nand U2218 (N_2218,In_346,In_208);
nand U2219 (N_2219,In_10,In_153);
and U2220 (N_2220,In_495,In_811);
nor U2221 (N_2221,In_1382,In_1495);
and U2222 (N_2222,In_1137,In_880);
and U2223 (N_2223,In_29,In_337);
nor U2224 (N_2224,In_548,In_1087);
or U2225 (N_2225,In_183,In_929);
or U2226 (N_2226,In_204,In_979);
nand U2227 (N_2227,In_413,In_1163);
nand U2228 (N_2228,In_357,In_1396);
nand U2229 (N_2229,In_299,In_1467);
xor U2230 (N_2230,In_1237,In_593);
nand U2231 (N_2231,In_1085,In_1405);
nor U2232 (N_2232,In_482,In_582);
nand U2233 (N_2233,In_574,In_1489);
or U2234 (N_2234,In_1254,In_578);
nand U2235 (N_2235,In_136,In_1301);
and U2236 (N_2236,In_693,In_89);
nand U2237 (N_2237,In_208,In_99);
nor U2238 (N_2238,In_481,In_140);
or U2239 (N_2239,In_246,In_979);
nor U2240 (N_2240,In_399,In_1017);
or U2241 (N_2241,In_1446,In_34);
xor U2242 (N_2242,In_331,In_1023);
or U2243 (N_2243,In_140,In_467);
and U2244 (N_2244,In_266,In_341);
nor U2245 (N_2245,In_577,In_236);
nand U2246 (N_2246,In_37,In_923);
xnor U2247 (N_2247,In_1259,In_456);
and U2248 (N_2248,In_1173,In_989);
and U2249 (N_2249,In_1412,In_572);
nand U2250 (N_2250,In_965,In_540);
nand U2251 (N_2251,In_900,In_746);
or U2252 (N_2252,In_1044,In_475);
xor U2253 (N_2253,In_1141,In_652);
xnor U2254 (N_2254,In_312,In_713);
or U2255 (N_2255,In_525,In_1262);
nand U2256 (N_2256,In_1420,In_146);
and U2257 (N_2257,In_765,In_461);
and U2258 (N_2258,In_242,In_667);
nor U2259 (N_2259,In_660,In_646);
xor U2260 (N_2260,In_1306,In_107);
xor U2261 (N_2261,In_1318,In_327);
nor U2262 (N_2262,In_1354,In_1324);
nor U2263 (N_2263,In_254,In_535);
or U2264 (N_2264,In_455,In_203);
xnor U2265 (N_2265,In_1276,In_610);
xor U2266 (N_2266,In_1282,In_574);
and U2267 (N_2267,In_1330,In_564);
or U2268 (N_2268,In_437,In_356);
and U2269 (N_2269,In_967,In_185);
xnor U2270 (N_2270,In_434,In_571);
and U2271 (N_2271,In_884,In_1255);
nand U2272 (N_2272,In_1099,In_1183);
or U2273 (N_2273,In_252,In_961);
and U2274 (N_2274,In_775,In_674);
or U2275 (N_2275,In_1443,In_1170);
and U2276 (N_2276,In_37,In_545);
xnor U2277 (N_2277,In_381,In_494);
nor U2278 (N_2278,In_372,In_1058);
or U2279 (N_2279,In_197,In_313);
nand U2280 (N_2280,In_860,In_618);
nor U2281 (N_2281,In_1245,In_516);
nand U2282 (N_2282,In_1038,In_333);
or U2283 (N_2283,In_1155,In_1460);
nor U2284 (N_2284,In_1273,In_285);
xnor U2285 (N_2285,In_302,In_444);
xor U2286 (N_2286,In_888,In_483);
nor U2287 (N_2287,In_695,In_1031);
nand U2288 (N_2288,In_758,In_1157);
nand U2289 (N_2289,In_119,In_47);
and U2290 (N_2290,In_694,In_179);
nor U2291 (N_2291,In_1434,In_580);
or U2292 (N_2292,In_838,In_218);
nand U2293 (N_2293,In_718,In_439);
nor U2294 (N_2294,In_1076,In_467);
and U2295 (N_2295,In_1290,In_1013);
nor U2296 (N_2296,In_1431,In_1156);
or U2297 (N_2297,In_1302,In_365);
nand U2298 (N_2298,In_572,In_1103);
and U2299 (N_2299,In_169,In_1260);
and U2300 (N_2300,In_1310,In_348);
nor U2301 (N_2301,In_120,In_582);
or U2302 (N_2302,In_1041,In_224);
nor U2303 (N_2303,In_1029,In_694);
and U2304 (N_2304,In_537,In_1372);
or U2305 (N_2305,In_1229,In_288);
and U2306 (N_2306,In_277,In_547);
nor U2307 (N_2307,In_848,In_530);
nand U2308 (N_2308,In_18,In_1430);
or U2309 (N_2309,In_413,In_1395);
or U2310 (N_2310,In_1258,In_1156);
nand U2311 (N_2311,In_860,In_219);
xor U2312 (N_2312,In_1300,In_931);
nor U2313 (N_2313,In_548,In_649);
nand U2314 (N_2314,In_93,In_804);
nand U2315 (N_2315,In_1009,In_257);
nand U2316 (N_2316,In_473,In_1269);
xnor U2317 (N_2317,In_1474,In_489);
and U2318 (N_2318,In_1473,In_855);
and U2319 (N_2319,In_513,In_118);
nand U2320 (N_2320,In_358,In_1437);
xnor U2321 (N_2321,In_1461,In_978);
and U2322 (N_2322,In_171,In_183);
nand U2323 (N_2323,In_536,In_165);
nand U2324 (N_2324,In_1420,In_1305);
or U2325 (N_2325,In_1273,In_884);
xnor U2326 (N_2326,In_554,In_735);
or U2327 (N_2327,In_85,In_1151);
or U2328 (N_2328,In_1127,In_119);
and U2329 (N_2329,In_1275,In_1117);
or U2330 (N_2330,In_842,In_852);
or U2331 (N_2331,In_106,In_442);
xor U2332 (N_2332,In_866,In_620);
nand U2333 (N_2333,In_38,In_579);
and U2334 (N_2334,In_475,In_893);
nor U2335 (N_2335,In_1454,In_914);
or U2336 (N_2336,In_554,In_358);
nor U2337 (N_2337,In_683,In_1188);
and U2338 (N_2338,In_1385,In_502);
nand U2339 (N_2339,In_952,In_283);
and U2340 (N_2340,In_1445,In_793);
nor U2341 (N_2341,In_294,In_600);
xnor U2342 (N_2342,In_1011,In_268);
nand U2343 (N_2343,In_920,In_583);
or U2344 (N_2344,In_1003,In_1);
xnor U2345 (N_2345,In_570,In_936);
nand U2346 (N_2346,In_689,In_383);
and U2347 (N_2347,In_192,In_437);
and U2348 (N_2348,In_1054,In_7);
nand U2349 (N_2349,In_1156,In_73);
xor U2350 (N_2350,In_1086,In_303);
and U2351 (N_2351,In_84,In_1482);
xnor U2352 (N_2352,In_547,In_1088);
nor U2353 (N_2353,In_642,In_326);
xor U2354 (N_2354,In_1412,In_50);
nand U2355 (N_2355,In_969,In_638);
and U2356 (N_2356,In_876,In_1035);
nor U2357 (N_2357,In_1112,In_1003);
nand U2358 (N_2358,In_1137,In_698);
and U2359 (N_2359,In_1390,In_259);
and U2360 (N_2360,In_1404,In_802);
xnor U2361 (N_2361,In_1326,In_307);
xnor U2362 (N_2362,In_1203,In_580);
nor U2363 (N_2363,In_788,In_1182);
and U2364 (N_2364,In_36,In_867);
or U2365 (N_2365,In_1003,In_580);
or U2366 (N_2366,In_1125,In_1406);
nor U2367 (N_2367,In_847,In_572);
nand U2368 (N_2368,In_1091,In_576);
nor U2369 (N_2369,In_867,In_357);
or U2370 (N_2370,In_415,In_1386);
nand U2371 (N_2371,In_1189,In_1039);
xnor U2372 (N_2372,In_599,In_251);
or U2373 (N_2373,In_970,In_1020);
nor U2374 (N_2374,In_1130,In_1420);
or U2375 (N_2375,In_1055,In_780);
or U2376 (N_2376,In_841,In_6);
nand U2377 (N_2377,In_1391,In_582);
nand U2378 (N_2378,In_28,In_445);
nand U2379 (N_2379,In_10,In_47);
and U2380 (N_2380,In_1074,In_595);
and U2381 (N_2381,In_935,In_833);
nor U2382 (N_2382,In_1459,In_673);
nand U2383 (N_2383,In_991,In_617);
xnor U2384 (N_2384,In_947,In_217);
nand U2385 (N_2385,In_290,In_46);
and U2386 (N_2386,In_431,In_129);
xor U2387 (N_2387,In_994,In_119);
nand U2388 (N_2388,In_703,In_907);
nand U2389 (N_2389,In_365,In_809);
xor U2390 (N_2390,In_323,In_452);
nand U2391 (N_2391,In_1335,In_808);
and U2392 (N_2392,In_1037,In_1468);
xnor U2393 (N_2393,In_596,In_1122);
xnor U2394 (N_2394,In_1250,In_1214);
xor U2395 (N_2395,In_191,In_971);
and U2396 (N_2396,In_1400,In_651);
or U2397 (N_2397,In_1455,In_374);
nor U2398 (N_2398,In_803,In_1449);
or U2399 (N_2399,In_53,In_260);
xor U2400 (N_2400,In_1043,In_846);
and U2401 (N_2401,In_986,In_1320);
nand U2402 (N_2402,In_1334,In_1454);
nand U2403 (N_2403,In_1193,In_1495);
xor U2404 (N_2404,In_1191,In_1485);
and U2405 (N_2405,In_467,In_1046);
and U2406 (N_2406,In_739,In_202);
or U2407 (N_2407,In_1466,In_82);
nand U2408 (N_2408,In_662,In_58);
xnor U2409 (N_2409,In_35,In_531);
nand U2410 (N_2410,In_267,In_590);
xnor U2411 (N_2411,In_350,In_968);
xor U2412 (N_2412,In_60,In_55);
nand U2413 (N_2413,In_547,In_1182);
nor U2414 (N_2414,In_1448,In_870);
or U2415 (N_2415,In_1116,In_808);
xor U2416 (N_2416,In_942,In_1086);
xor U2417 (N_2417,In_920,In_1176);
nor U2418 (N_2418,In_201,In_1488);
or U2419 (N_2419,In_514,In_813);
or U2420 (N_2420,In_324,In_964);
nand U2421 (N_2421,In_682,In_749);
and U2422 (N_2422,In_741,In_127);
nor U2423 (N_2423,In_1389,In_846);
and U2424 (N_2424,In_541,In_127);
nor U2425 (N_2425,In_942,In_540);
xor U2426 (N_2426,In_359,In_1351);
nand U2427 (N_2427,In_863,In_1201);
xor U2428 (N_2428,In_1077,In_789);
nor U2429 (N_2429,In_383,In_194);
nand U2430 (N_2430,In_1383,In_4);
or U2431 (N_2431,In_368,In_601);
and U2432 (N_2432,In_930,In_1482);
nand U2433 (N_2433,In_1114,In_371);
or U2434 (N_2434,In_528,In_173);
nor U2435 (N_2435,In_420,In_78);
or U2436 (N_2436,In_992,In_257);
or U2437 (N_2437,In_935,In_1155);
and U2438 (N_2438,In_139,In_764);
and U2439 (N_2439,In_1412,In_436);
xor U2440 (N_2440,In_1412,In_1048);
nor U2441 (N_2441,In_8,In_90);
nor U2442 (N_2442,In_193,In_821);
and U2443 (N_2443,In_1228,In_1129);
nand U2444 (N_2444,In_575,In_44);
and U2445 (N_2445,In_617,In_549);
and U2446 (N_2446,In_922,In_1221);
and U2447 (N_2447,In_972,In_1306);
xor U2448 (N_2448,In_486,In_973);
nor U2449 (N_2449,In_1090,In_926);
xor U2450 (N_2450,In_1103,In_1075);
and U2451 (N_2451,In_1342,In_649);
or U2452 (N_2452,In_458,In_444);
nor U2453 (N_2453,In_802,In_1140);
nand U2454 (N_2454,In_160,In_571);
nand U2455 (N_2455,In_1154,In_905);
nand U2456 (N_2456,In_384,In_77);
nand U2457 (N_2457,In_1482,In_1420);
xnor U2458 (N_2458,In_926,In_1068);
and U2459 (N_2459,In_707,In_1164);
and U2460 (N_2460,In_488,In_875);
nand U2461 (N_2461,In_1076,In_1166);
and U2462 (N_2462,In_311,In_293);
nand U2463 (N_2463,In_1227,In_1487);
nand U2464 (N_2464,In_568,In_1468);
nand U2465 (N_2465,In_794,In_1043);
or U2466 (N_2466,In_202,In_640);
nand U2467 (N_2467,In_954,In_898);
or U2468 (N_2468,In_1084,In_878);
xnor U2469 (N_2469,In_672,In_624);
xnor U2470 (N_2470,In_23,In_752);
and U2471 (N_2471,In_1256,In_1477);
or U2472 (N_2472,In_1339,In_667);
xnor U2473 (N_2473,In_1347,In_1329);
nor U2474 (N_2474,In_428,In_816);
nor U2475 (N_2475,In_650,In_1291);
and U2476 (N_2476,In_1011,In_1242);
nor U2477 (N_2477,In_1183,In_537);
nor U2478 (N_2478,In_495,In_1337);
or U2479 (N_2479,In_1355,In_1357);
nand U2480 (N_2480,In_545,In_1384);
and U2481 (N_2481,In_1302,In_209);
nand U2482 (N_2482,In_1036,In_1034);
nor U2483 (N_2483,In_1333,In_1359);
or U2484 (N_2484,In_1314,In_571);
nand U2485 (N_2485,In_1486,In_234);
and U2486 (N_2486,In_96,In_1403);
or U2487 (N_2487,In_1475,In_1456);
nor U2488 (N_2488,In_1025,In_753);
or U2489 (N_2489,In_1312,In_834);
nor U2490 (N_2490,In_1047,In_723);
xnor U2491 (N_2491,In_1430,In_735);
nand U2492 (N_2492,In_210,In_1067);
or U2493 (N_2493,In_1429,In_1393);
nand U2494 (N_2494,In_1081,In_428);
and U2495 (N_2495,In_457,In_1407);
xor U2496 (N_2496,In_1153,In_1226);
nand U2497 (N_2497,In_723,In_372);
or U2498 (N_2498,In_892,In_512);
xnor U2499 (N_2499,In_887,In_26);
xor U2500 (N_2500,In_1001,In_1010);
nand U2501 (N_2501,In_170,In_1460);
or U2502 (N_2502,In_45,In_153);
nand U2503 (N_2503,In_279,In_407);
and U2504 (N_2504,In_482,In_607);
nand U2505 (N_2505,In_965,In_1450);
or U2506 (N_2506,In_656,In_1085);
nor U2507 (N_2507,In_884,In_1259);
and U2508 (N_2508,In_902,In_954);
or U2509 (N_2509,In_336,In_1380);
or U2510 (N_2510,In_162,In_290);
and U2511 (N_2511,In_1292,In_120);
nor U2512 (N_2512,In_261,In_970);
xnor U2513 (N_2513,In_585,In_607);
nor U2514 (N_2514,In_152,In_532);
and U2515 (N_2515,In_883,In_1384);
or U2516 (N_2516,In_173,In_558);
and U2517 (N_2517,In_327,In_422);
or U2518 (N_2518,In_1011,In_1278);
or U2519 (N_2519,In_265,In_1408);
or U2520 (N_2520,In_1027,In_1351);
and U2521 (N_2521,In_125,In_435);
and U2522 (N_2522,In_296,In_828);
and U2523 (N_2523,In_1263,In_355);
or U2524 (N_2524,In_793,In_1042);
and U2525 (N_2525,In_1353,In_1405);
xnor U2526 (N_2526,In_1170,In_909);
and U2527 (N_2527,In_489,In_1453);
nor U2528 (N_2528,In_1279,In_190);
nor U2529 (N_2529,In_997,In_1074);
xnor U2530 (N_2530,In_1128,In_357);
xnor U2531 (N_2531,In_631,In_787);
nor U2532 (N_2532,In_1223,In_1197);
nand U2533 (N_2533,In_268,In_570);
and U2534 (N_2534,In_179,In_1444);
xnor U2535 (N_2535,In_1344,In_970);
or U2536 (N_2536,In_64,In_393);
or U2537 (N_2537,In_639,In_1461);
nor U2538 (N_2538,In_1102,In_104);
nor U2539 (N_2539,In_1408,In_1121);
or U2540 (N_2540,In_233,In_254);
or U2541 (N_2541,In_793,In_790);
nor U2542 (N_2542,In_846,In_1180);
nand U2543 (N_2543,In_1056,In_1402);
or U2544 (N_2544,In_449,In_104);
nor U2545 (N_2545,In_1212,In_940);
or U2546 (N_2546,In_1243,In_1260);
and U2547 (N_2547,In_812,In_1205);
and U2548 (N_2548,In_1424,In_1426);
or U2549 (N_2549,In_1239,In_852);
xnor U2550 (N_2550,In_929,In_868);
or U2551 (N_2551,In_1305,In_1266);
nor U2552 (N_2552,In_162,In_812);
xor U2553 (N_2553,In_1195,In_606);
nor U2554 (N_2554,In_443,In_719);
nor U2555 (N_2555,In_305,In_211);
nand U2556 (N_2556,In_265,In_755);
and U2557 (N_2557,In_950,In_1287);
or U2558 (N_2558,In_1251,In_280);
nor U2559 (N_2559,In_434,In_1242);
and U2560 (N_2560,In_107,In_140);
xor U2561 (N_2561,In_1467,In_1309);
and U2562 (N_2562,In_1303,In_245);
nor U2563 (N_2563,In_755,In_1496);
xnor U2564 (N_2564,In_122,In_998);
and U2565 (N_2565,In_1304,In_1217);
nand U2566 (N_2566,In_1416,In_574);
nand U2567 (N_2567,In_884,In_631);
or U2568 (N_2568,In_648,In_379);
or U2569 (N_2569,In_743,In_165);
xor U2570 (N_2570,In_1218,In_1288);
nor U2571 (N_2571,In_559,In_417);
or U2572 (N_2572,In_835,In_540);
xor U2573 (N_2573,In_1211,In_8);
nand U2574 (N_2574,In_643,In_1209);
nor U2575 (N_2575,In_113,In_155);
nand U2576 (N_2576,In_1339,In_198);
or U2577 (N_2577,In_1007,In_1279);
or U2578 (N_2578,In_1218,In_145);
nand U2579 (N_2579,In_1263,In_1271);
nor U2580 (N_2580,In_423,In_615);
nand U2581 (N_2581,In_333,In_795);
xor U2582 (N_2582,In_413,In_922);
and U2583 (N_2583,In_1138,In_556);
nand U2584 (N_2584,In_460,In_1334);
nor U2585 (N_2585,In_889,In_1159);
and U2586 (N_2586,In_640,In_638);
nor U2587 (N_2587,In_1238,In_1076);
and U2588 (N_2588,In_810,In_1385);
and U2589 (N_2589,In_208,In_1393);
xor U2590 (N_2590,In_801,In_1173);
or U2591 (N_2591,In_1465,In_136);
nor U2592 (N_2592,In_1237,In_25);
xnor U2593 (N_2593,In_831,In_878);
and U2594 (N_2594,In_808,In_1397);
or U2595 (N_2595,In_1133,In_754);
nand U2596 (N_2596,In_624,In_823);
or U2597 (N_2597,In_1410,In_793);
nor U2598 (N_2598,In_1072,In_1358);
and U2599 (N_2599,In_1332,In_568);
nor U2600 (N_2600,In_491,In_247);
or U2601 (N_2601,In_731,In_995);
nor U2602 (N_2602,In_1272,In_391);
and U2603 (N_2603,In_714,In_1339);
and U2604 (N_2604,In_950,In_53);
xnor U2605 (N_2605,In_593,In_1418);
xnor U2606 (N_2606,In_525,In_54);
xor U2607 (N_2607,In_1305,In_1402);
xor U2608 (N_2608,In_788,In_467);
nor U2609 (N_2609,In_654,In_1088);
nor U2610 (N_2610,In_862,In_638);
nor U2611 (N_2611,In_603,In_890);
nor U2612 (N_2612,In_371,In_1431);
nand U2613 (N_2613,In_1357,In_966);
or U2614 (N_2614,In_360,In_1255);
and U2615 (N_2615,In_984,In_1156);
nand U2616 (N_2616,In_852,In_77);
xnor U2617 (N_2617,In_1178,In_866);
or U2618 (N_2618,In_993,In_1311);
xnor U2619 (N_2619,In_1211,In_1295);
nand U2620 (N_2620,In_225,In_1373);
xnor U2621 (N_2621,In_479,In_430);
nand U2622 (N_2622,In_880,In_1330);
or U2623 (N_2623,In_1051,In_312);
nor U2624 (N_2624,In_8,In_1007);
and U2625 (N_2625,In_483,In_629);
xnor U2626 (N_2626,In_175,In_881);
or U2627 (N_2627,In_520,In_655);
and U2628 (N_2628,In_581,In_165);
or U2629 (N_2629,In_322,In_217);
xnor U2630 (N_2630,In_1195,In_660);
nand U2631 (N_2631,In_606,In_88);
and U2632 (N_2632,In_799,In_912);
and U2633 (N_2633,In_354,In_520);
xnor U2634 (N_2634,In_692,In_346);
or U2635 (N_2635,In_1400,In_679);
and U2636 (N_2636,In_171,In_258);
or U2637 (N_2637,In_777,In_74);
and U2638 (N_2638,In_397,In_66);
nor U2639 (N_2639,In_1242,In_1378);
and U2640 (N_2640,In_596,In_356);
and U2641 (N_2641,In_610,In_1270);
or U2642 (N_2642,In_623,In_830);
nor U2643 (N_2643,In_855,In_1423);
and U2644 (N_2644,In_94,In_1227);
and U2645 (N_2645,In_901,In_1104);
nand U2646 (N_2646,In_439,In_606);
nand U2647 (N_2647,In_1079,In_452);
and U2648 (N_2648,In_431,In_1021);
xor U2649 (N_2649,In_1336,In_1405);
nand U2650 (N_2650,In_57,In_424);
nor U2651 (N_2651,In_1184,In_64);
nand U2652 (N_2652,In_1311,In_444);
and U2653 (N_2653,In_431,In_172);
nor U2654 (N_2654,In_385,In_37);
nand U2655 (N_2655,In_413,In_269);
xor U2656 (N_2656,In_235,In_90);
nor U2657 (N_2657,In_135,In_482);
xor U2658 (N_2658,In_106,In_829);
nand U2659 (N_2659,In_496,In_1261);
nand U2660 (N_2660,In_588,In_322);
xor U2661 (N_2661,In_107,In_245);
nand U2662 (N_2662,In_2,In_1364);
nor U2663 (N_2663,In_75,In_213);
and U2664 (N_2664,In_880,In_250);
or U2665 (N_2665,In_354,In_864);
xor U2666 (N_2666,In_816,In_1160);
nand U2667 (N_2667,In_1269,In_1129);
and U2668 (N_2668,In_598,In_1286);
and U2669 (N_2669,In_1295,In_11);
nand U2670 (N_2670,In_1029,In_622);
or U2671 (N_2671,In_879,In_827);
nand U2672 (N_2672,In_943,In_170);
nand U2673 (N_2673,In_1206,In_1028);
xor U2674 (N_2674,In_686,In_605);
or U2675 (N_2675,In_874,In_240);
or U2676 (N_2676,In_632,In_864);
nand U2677 (N_2677,In_38,In_553);
nor U2678 (N_2678,In_751,In_141);
nand U2679 (N_2679,In_910,In_1473);
and U2680 (N_2680,In_441,In_505);
nor U2681 (N_2681,In_1469,In_1264);
nor U2682 (N_2682,In_266,In_98);
and U2683 (N_2683,In_181,In_496);
nor U2684 (N_2684,In_544,In_1029);
nor U2685 (N_2685,In_1168,In_1075);
or U2686 (N_2686,In_319,In_1426);
nand U2687 (N_2687,In_792,In_218);
and U2688 (N_2688,In_1311,In_288);
xor U2689 (N_2689,In_605,In_630);
xnor U2690 (N_2690,In_1479,In_42);
or U2691 (N_2691,In_233,In_862);
and U2692 (N_2692,In_1054,In_0);
or U2693 (N_2693,In_1312,In_1478);
and U2694 (N_2694,In_263,In_1156);
and U2695 (N_2695,In_1027,In_840);
xor U2696 (N_2696,In_1169,In_910);
and U2697 (N_2697,In_1199,In_386);
xor U2698 (N_2698,In_1400,In_853);
or U2699 (N_2699,In_1373,In_461);
nor U2700 (N_2700,In_1429,In_1059);
and U2701 (N_2701,In_129,In_546);
xnor U2702 (N_2702,In_1146,In_1182);
nand U2703 (N_2703,In_762,In_864);
nor U2704 (N_2704,In_1000,In_44);
nor U2705 (N_2705,In_1487,In_76);
or U2706 (N_2706,In_1138,In_420);
or U2707 (N_2707,In_967,In_910);
xnor U2708 (N_2708,In_819,In_669);
and U2709 (N_2709,In_266,In_1412);
nand U2710 (N_2710,In_133,In_313);
xnor U2711 (N_2711,In_925,In_179);
nor U2712 (N_2712,In_1042,In_1054);
or U2713 (N_2713,In_0,In_1224);
and U2714 (N_2714,In_1051,In_580);
and U2715 (N_2715,In_1139,In_855);
or U2716 (N_2716,In_351,In_1321);
xor U2717 (N_2717,In_675,In_1268);
or U2718 (N_2718,In_295,In_1342);
and U2719 (N_2719,In_963,In_948);
xnor U2720 (N_2720,In_1008,In_808);
nand U2721 (N_2721,In_486,In_7);
nand U2722 (N_2722,In_412,In_766);
and U2723 (N_2723,In_573,In_385);
or U2724 (N_2724,In_1076,In_435);
nor U2725 (N_2725,In_779,In_1264);
and U2726 (N_2726,In_135,In_218);
nand U2727 (N_2727,In_281,In_1138);
nand U2728 (N_2728,In_95,In_9);
nand U2729 (N_2729,In_519,In_986);
and U2730 (N_2730,In_23,In_770);
nand U2731 (N_2731,In_897,In_153);
and U2732 (N_2732,In_745,In_712);
nand U2733 (N_2733,In_27,In_1066);
or U2734 (N_2734,In_10,In_208);
xnor U2735 (N_2735,In_857,In_707);
nor U2736 (N_2736,In_425,In_240);
nor U2737 (N_2737,In_892,In_777);
nand U2738 (N_2738,In_481,In_1452);
nand U2739 (N_2739,In_1153,In_964);
or U2740 (N_2740,In_544,In_1234);
or U2741 (N_2741,In_821,In_803);
nand U2742 (N_2742,In_1004,In_407);
xnor U2743 (N_2743,In_1414,In_540);
or U2744 (N_2744,In_415,In_906);
nor U2745 (N_2745,In_245,In_1111);
and U2746 (N_2746,In_601,In_688);
xnor U2747 (N_2747,In_191,In_221);
xor U2748 (N_2748,In_881,In_1427);
xnor U2749 (N_2749,In_681,In_199);
or U2750 (N_2750,In_723,In_1139);
or U2751 (N_2751,In_305,In_746);
xnor U2752 (N_2752,In_967,In_1138);
nand U2753 (N_2753,In_621,In_1386);
nor U2754 (N_2754,In_1361,In_244);
nand U2755 (N_2755,In_849,In_1123);
or U2756 (N_2756,In_698,In_349);
and U2757 (N_2757,In_332,In_1107);
xnor U2758 (N_2758,In_584,In_212);
xnor U2759 (N_2759,In_949,In_16);
nor U2760 (N_2760,In_1448,In_16);
and U2761 (N_2761,In_202,In_989);
xnor U2762 (N_2762,In_1378,In_834);
nor U2763 (N_2763,In_1086,In_1368);
nor U2764 (N_2764,In_325,In_1204);
nor U2765 (N_2765,In_833,In_1341);
and U2766 (N_2766,In_1264,In_682);
nand U2767 (N_2767,In_1146,In_782);
xnor U2768 (N_2768,In_1326,In_1452);
and U2769 (N_2769,In_1362,In_336);
and U2770 (N_2770,In_534,In_955);
or U2771 (N_2771,In_793,In_1061);
nor U2772 (N_2772,In_744,In_1368);
xor U2773 (N_2773,In_446,In_1000);
nand U2774 (N_2774,In_106,In_9);
nor U2775 (N_2775,In_1073,In_1360);
xor U2776 (N_2776,In_585,In_1131);
xor U2777 (N_2777,In_54,In_261);
and U2778 (N_2778,In_1039,In_1102);
nor U2779 (N_2779,In_1336,In_244);
or U2780 (N_2780,In_1372,In_1495);
or U2781 (N_2781,In_670,In_915);
nand U2782 (N_2782,In_711,In_668);
or U2783 (N_2783,In_660,In_209);
and U2784 (N_2784,In_194,In_450);
nand U2785 (N_2785,In_557,In_132);
or U2786 (N_2786,In_1150,In_797);
or U2787 (N_2787,In_882,In_434);
xor U2788 (N_2788,In_918,In_120);
or U2789 (N_2789,In_695,In_645);
and U2790 (N_2790,In_778,In_549);
nand U2791 (N_2791,In_151,In_875);
or U2792 (N_2792,In_954,In_882);
xor U2793 (N_2793,In_724,In_1052);
and U2794 (N_2794,In_820,In_824);
nand U2795 (N_2795,In_504,In_777);
nand U2796 (N_2796,In_1352,In_152);
or U2797 (N_2797,In_1020,In_130);
or U2798 (N_2798,In_716,In_1353);
nor U2799 (N_2799,In_916,In_1382);
nor U2800 (N_2800,In_360,In_1125);
and U2801 (N_2801,In_1101,In_1353);
and U2802 (N_2802,In_868,In_190);
nand U2803 (N_2803,In_69,In_1373);
and U2804 (N_2804,In_1366,In_1259);
nor U2805 (N_2805,In_1183,In_336);
nand U2806 (N_2806,In_578,In_907);
xor U2807 (N_2807,In_115,In_1391);
xor U2808 (N_2808,In_1130,In_1452);
nand U2809 (N_2809,In_1406,In_374);
and U2810 (N_2810,In_348,In_785);
or U2811 (N_2811,In_1176,In_469);
and U2812 (N_2812,In_289,In_1297);
or U2813 (N_2813,In_661,In_1205);
nor U2814 (N_2814,In_846,In_892);
nand U2815 (N_2815,In_406,In_60);
and U2816 (N_2816,In_446,In_176);
nand U2817 (N_2817,In_543,In_782);
nand U2818 (N_2818,In_1418,In_863);
or U2819 (N_2819,In_1399,In_1024);
or U2820 (N_2820,In_268,In_1094);
nand U2821 (N_2821,In_1427,In_297);
nor U2822 (N_2822,In_729,In_765);
xor U2823 (N_2823,In_532,In_173);
nand U2824 (N_2824,In_275,In_857);
or U2825 (N_2825,In_238,In_661);
and U2826 (N_2826,In_468,In_965);
xor U2827 (N_2827,In_66,In_1150);
nor U2828 (N_2828,In_987,In_109);
xnor U2829 (N_2829,In_439,In_493);
or U2830 (N_2830,In_1024,In_139);
and U2831 (N_2831,In_578,In_488);
or U2832 (N_2832,In_257,In_763);
xnor U2833 (N_2833,In_232,In_777);
nor U2834 (N_2834,In_89,In_474);
xor U2835 (N_2835,In_1009,In_888);
nand U2836 (N_2836,In_655,In_640);
nor U2837 (N_2837,In_340,In_1361);
nor U2838 (N_2838,In_1013,In_795);
and U2839 (N_2839,In_1362,In_1271);
or U2840 (N_2840,In_1401,In_964);
nand U2841 (N_2841,In_1363,In_992);
and U2842 (N_2842,In_409,In_1087);
nand U2843 (N_2843,In_80,In_813);
nand U2844 (N_2844,In_1250,In_303);
nor U2845 (N_2845,In_292,In_623);
xnor U2846 (N_2846,In_193,In_496);
or U2847 (N_2847,In_1231,In_1433);
and U2848 (N_2848,In_335,In_809);
nand U2849 (N_2849,In_1168,In_1126);
xnor U2850 (N_2850,In_1365,In_799);
xor U2851 (N_2851,In_19,In_1470);
nand U2852 (N_2852,In_77,In_269);
or U2853 (N_2853,In_143,In_734);
nor U2854 (N_2854,In_471,In_1359);
xor U2855 (N_2855,In_1112,In_325);
nor U2856 (N_2856,In_1068,In_1194);
xnor U2857 (N_2857,In_1034,In_34);
nor U2858 (N_2858,In_713,In_1387);
xnor U2859 (N_2859,In_1098,In_41);
xnor U2860 (N_2860,In_643,In_1387);
xnor U2861 (N_2861,In_566,In_1359);
xor U2862 (N_2862,In_1147,In_845);
xnor U2863 (N_2863,In_608,In_854);
or U2864 (N_2864,In_672,In_484);
nand U2865 (N_2865,In_847,In_301);
nand U2866 (N_2866,In_1299,In_989);
or U2867 (N_2867,In_222,In_1340);
or U2868 (N_2868,In_1214,In_1206);
and U2869 (N_2869,In_3,In_541);
xor U2870 (N_2870,In_1340,In_1132);
nand U2871 (N_2871,In_840,In_278);
nor U2872 (N_2872,In_1427,In_1298);
nor U2873 (N_2873,In_417,In_966);
nand U2874 (N_2874,In_1438,In_220);
or U2875 (N_2875,In_883,In_1348);
nand U2876 (N_2876,In_1066,In_1232);
nor U2877 (N_2877,In_1252,In_33);
and U2878 (N_2878,In_913,In_201);
nand U2879 (N_2879,In_312,In_637);
or U2880 (N_2880,In_1443,In_452);
nand U2881 (N_2881,In_86,In_827);
nand U2882 (N_2882,In_1427,In_820);
and U2883 (N_2883,In_1116,In_572);
nand U2884 (N_2884,In_581,In_1427);
nand U2885 (N_2885,In_1287,In_576);
nand U2886 (N_2886,In_458,In_968);
or U2887 (N_2887,In_42,In_1264);
and U2888 (N_2888,In_1313,In_348);
nor U2889 (N_2889,In_566,In_337);
and U2890 (N_2890,In_156,In_536);
xnor U2891 (N_2891,In_256,In_1065);
and U2892 (N_2892,In_1478,In_72);
nor U2893 (N_2893,In_669,In_592);
nor U2894 (N_2894,In_1111,In_1456);
or U2895 (N_2895,In_1307,In_676);
nor U2896 (N_2896,In_1057,In_80);
nand U2897 (N_2897,In_109,In_1226);
nor U2898 (N_2898,In_1477,In_811);
nor U2899 (N_2899,In_1173,In_25);
and U2900 (N_2900,In_1436,In_504);
or U2901 (N_2901,In_905,In_753);
nor U2902 (N_2902,In_801,In_279);
nand U2903 (N_2903,In_229,In_919);
or U2904 (N_2904,In_607,In_216);
and U2905 (N_2905,In_985,In_920);
xnor U2906 (N_2906,In_816,In_74);
nand U2907 (N_2907,In_700,In_1337);
xnor U2908 (N_2908,In_49,In_244);
or U2909 (N_2909,In_870,In_1128);
and U2910 (N_2910,In_637,In_73);
or U2911 (N_2911,In_600,In_146);
xnor U2912 (N_2912,In_1110,In_818);
or U2913 (N_2913,In_205,In_115);
nand U2914 (N_2914,In_0,In_785);
nor U2915 (N_2915,In_1460,In_1308);
nor U2916 (N_2916,In_1495,In_541);
nand U2917 (N_2917,In_1491,In_1192);
or U2918 (N_2918,In_518,In_1147);
xor U2919 (N_2919,In_191,In_108);
or U2920 (N_2920,In_750,In_986);
nand U2921 (N_2921,In_1391,In_1316);
xnor U2922 (N_2922,In_139,In_84);
nor U2923 (N_2923,In_837,In_1094);
and U2924 (N_2924,In_777,In_1481);
xor U2925 (N_2925,In_392,In_558);
or U2926 (N_2926,In_325,In_204);
or U2927 (N_2927,In_1241,In_462);
xnor U2928 (N_2928,In_365,In_313);
nand U2929 (N_2929,In_1204,In_1054);
nor U2930 (N_2930,In_973,In_884);
and U2931 (N_2931,In_361,In_1317);
nand U2932 (N_2932,In_753,In_342);
nor U2933 (N_2933,In_1426,In_1430);
or U2934 (N_2934,In_661,In_66);
nand U2935 (N_2935,In_776,In_736);
nor U2936 (N_2936,In_443,In_888);
nor U2937 (N_2937,In_66,In_1147);
or U2938 (N_2938,In_598,In_925);
and U2939 (N_2939,In_69,In_233);
nand U2940 (N_2940,In_1279,In_148);
and U2941 (N_2941,In_1316,In_442);
and U2942 (N_2942,In_810,In_42);
nand U2943 (N_2943,In_1395,In_893);
nand U2944 (N_2944,In_1422,In_242);
xor U2945 (N_2945,In_1313,In_1226);
nor U2946 (N_2946,In_1497,In_1049);
xnor U2947 (N_2947,In_1478,In_1484);
xnor U2948 (N_2948,In_688,In_410);
or U2949 (N_2949,In_136,In_694);
or U2950 (N_2950,In_97,In_1391);
and U2951 (N_2951,In_708,In_843);
nor U2952 (N_2952,In_413,In_425);
or U2953 (N_2953,In_1003,In_1479);
and U2954 (N_2954,In_55,In_64);
nor U2955 (N_2955,In_1067,In_207);
or U2956 (N_2956,In_939,In_761);
nor U2957 (N_2957,In_635,In_1315);
or U2958 (N_2958,In_494,In_114);
xor U2959 (N_2959,In_680,In_676);
or U2960 (N_2960,In_872,In_917);
nor U2961 (N_2961,In_608,In_832);
and U2962 (N_2962,In_586,In_1086);
nor U2963 (N_2963,In_1111,In_807);
or U2964 (N_2964,In_594,In_287);
nand U2965 (N_2965,In_1066,In_305);
and U2966 (N_2966,In_866,In_36);
nand U2967 (N_2967,In_264,In_1448);
nor U2968 (N_2968,In_241,In_528);
and U2969 (N_2969,In_149,In_1276);
nor U2970 (N_2970,In_1208,In_263);
xor U2971 (N_2971,In_1346,In_492);
nor U2972 (N_2972,In_1065,In_512);
xnor U2973 (N_2973,In_938,In_1164);
and U2974 (N_2974,In_632,In_1392);
or U2975 (N_2975,In_438,In_480);
and U2976 (N_2976,In_708,In_1034);
xor U2977 (N_2977,In_352,In_1469);
or U2978 (N_2978,In_954,In_1219);
xnor U2979 (N_2979,In_1414,In_62);
xnor U2980 (N_2980,In_1206,In_389);
or U2981 (N_2981,In_593,In_1254);
xor U2982 (N_2982,In_1263,In_850);
or U2983 (N_2983,In_1311,In_551);
xnor U2984 (N_2984,In_33,In_1416);
and U2985 (N_2985,In_1381,In_1487);
nand U2986 (N_2986,In_1320,In_18);
nand U2987 (N_2987,In_959,In_904);
nand U2988 (N_2988,In_81,In_1482);
xnor U2989 (N_2989,In_1062,In_1414);
nand U2990 (N_2990,In_957,In_245);
and U2991 (N_2991,In_491,In_404);
nor U2992 (N_2992,In_1144,In_297);
xnor U2993 (N_2993,In_617,In_742);
or U2994 (N_2994,In_1371,In_358);
nand U2995 (N_2995,In_404,In_1478);
nor U2996 (N_2996,In_610,In_579);
or U2997 (N_2997,In_1016,In_546);
nor U2998 (N_2998,In_1023,In_1002);
nand U2999 (N_2999,In_537,In_1159);
and U3000 (N_3000,In_1177,In_40);
and U3001 (N_3001,In_714,In_1188);
nor U3002 (N_3002,In_922,In_300);
or U3003 (N_3003,In_889,In_906);
xor U3004 (N_3004,In_1194,In_1439);
or U3005 (N_3005,In_178,In_799);
xnor U3006 (N_3006,In_142,In_267);
or U3007 (N_3007,In_907,In_653);
nor U3008 (N_3008,In_1215,In_831);
and U3009 (N_3009,In_825,In_752);
nand U3010 (N_3010,In_1027,In_148);
xor U3011 (N_3011,In_942,In_730);
and U3012 (N_3012,In_1265,In_1230);
and U3013 (N_3013,In_1073,In_454);
nor U3014 (N_3014,In_1036,In_260);
xnor U3015 (N_3015,In_386,In_990);
xnor U3016 (N_3016,In_955,In_593);
nand U3017 (N_3017,In_931,In_845);
or U3018 (N_3018,In_1410,In_174);
or U3019 (N_3019,In_640,In_1479);
or U3020 (N_3020,In_549,In_1289);
xnor U3021 (N_3021,In_1492,In_1204);
xnor U3022 (N_3022,In_1289,In_996);
and U3023 (N_3023,In_1216,In_556);
and U3024 (N_3024,In_13,In_1182);
xor U3025 (N_3025,In_345,In_1370);
and U3026 (N_3026,In_762,In_226);
or U3027 (N_3027,In_190,In_684);
or U3028 (N_3028,In_979,In_677);
and U3029 (N_3029,In_1184,In_465);
or U3030 (N_3030,In_1412,In_201);
nor U3031 (N_3031,In_501,In_877);
xor U3032 (N_3032,In_943,In_1469);
nand U3033 (N_3033,In_772,In_393);
xor U3034 (N_3034,In_63,In_1245);
xnor U3035 (N_3035,In_352,In_1218);
nor U3036 (N_3036,In_751,In_75);
nor U3037 (N_3037,In_1252,In_1128);
xnor U3038 (N_3038,In_1117,In_1474);
and U3039 (N_3039,In_1224,In_427);
nand U3040 (N_3040,In_801,In_1044);
xor U3041 (N_3041,In_1414,In_806);
xor U3042 (N_3042,In_439,In_1013);
nor U3043 (N_3043,In_269,In_704);
or U3044 (N_3044,In_434,In_215);
xor U3045 (N_3045,In_943,In_831);
and U3046 (N_3046,In_453,In_485);
and U3047 (N_3047,In_1407,In_1009);
nand U3048 (N_3048,In_265,In_816);
or U3049 (N_3049,In_344,In_220);
nor U3050 (N_3050,In_1296,In_312);
and U3051 (N_3051,In_728,In_1260);
nor U3052 (N_3052,In_1383,In_387);
or U3053 (N_3053,In_1088,In_1165);
or U3054 (N_3054,In_784,In_977);
or U3055 (N_3055,In_804,In_371);
and U3056 (N_3056,In_1482,In_1383);
nand U3057 (N_3057,In_1429,In_1334);
or U3058 (N_3058,In_1214,In_45);
nor U3059 (N_3059,In_239,In_822);
nor U3060 (N_3060,In_33,In_309);
nor U3061 (N_3061,In_1184,In_1294);
nor U3062 (N_3062,In_1437,In_87);
nand U3063 (N_3063,In_1447,In_1435);
and U3064 (N_3064,In_1433,In_765);
xor U3065 (N_3065,In_706,In_1389);
nand U3066 (N_3066,In_560,In_1171);
nor U3067 (N_3067,In_1350,In_978);
or U3068 (N_3068,In_974,In_746);
or U3069 (N_3069,In_1323,In_706);
xnor U3070 (N_3070,In_1005,In_1120);
or U3071 (N_3071,In_1414,In_1094);
nand U3072 (N_3072,In_1236,In_624);
nand U3073 (N_3073,In_1412,In_680);
and U3074 (N_3074,In_903,In_75);
xnor U3075 (N_3075,In_1058,In_660);
and U3076 (N_3076,In_802,In_1223);
xor U3077 (N_3077,In_1443,In_797);
nor U3078 (N_3078,In_671,In_623);
nor U3079 (N_3079,In_524,In_1457);
xnor U3080 (N_3080,In_1412,In_484);
nor U3081 (N_3081,In_1332,In_606);
or U3082 (N_3082,In_713,In_245);
xnor U3083 (N_3083,In_1450,In_637);
or U3084 (N_3084,In_487,In_34);
or U3085 (N_3085,In_591,In_473);
nand U3086 (N_3086,In_636,In_590);
nand U3087 (N_3087,In_1417,In_1347);
or U3088 (N_3088,In_447,In_595);
nand U3089 (N_3089,In_137,In_755);
or U3090 (N_3090,In_5,In_414);
xnor U3091 (N_3091,In_640,In_1017);
xor U3092 (N_3092,In_645,In_654);
nand U3093 (N_3093,In_1143,In_428);
xor U3094 (N_3094,In_211,In_152);
and U3095 (N_3095,In_479,In_1374);
xnor U3096 (N_3096,In_178,In_895);
xor U3097 (N_3097,In_391,In_992);
nand U3098 (N_3098,In_942,In_419);
nand U3099 (N_3099,In_214,In_680);
nand U3100 (N_3100,In_500,In_1168);
xor U3101 (N_3101,In_717,In_221);
nand U3102 (N_3102,In_251,In_1419);
nand U3103 (N_3103,In_1068,In_929);
nor U3104 (N_3104,In_1106,In_304);
nor U3105 (N_3105,In_1196,In_826);
nand U3106 (N_3106,In_1195,In_1030);
nand U3107 (N_3107,In_416,In_471);
nand U3108 (N_3108,In_24,In_204);
nor U3109 (N_3109,In_262,In_1262);
nor U3110 (N_3110,In_1487,In_745);
or U3111 (N_3111,In_187,In_731);
nor U3112 (N_3112,In_767,In_898);
or U3113 (N_3113,In_432,In_609);
xnor U3114 (N_3114,In_1259,In_197);
nand U3115 (N_3115,In_1008,In_342);
nor U3116 (N_3116,In_298,In_325);
or U3117 (N_3117,In_1494,In_1174);
nand U3118 (N_3118,In_37,In_541);
nor U3119 (N_3119,In_869,In_740);
and U3120 (N_3120,In_1323,In_388);
nand U3121 (N_3121,In_893,In_748);
or U3122 (N_3122,In_1071,In_478);
or U3123 (N_3123,In_905,In_14);
or U3124 (N_3124,In_932,In_688);
or U3125 (N_3125,In_161,In_1045);
nor U3126 (N_3126,In_334,In_578);
and U3127 (N_3127,In_882,In_309);
and U3128 (N_3128,In_1369,In_1437);
and U3129 (N_3129,In_566,In_1211);
xnor U3130 (N_3130,In_143,In_659);
nand U3131 (N_3131,In_233,In_1164);
nand U3132 (N_3132,In_1450,In_283);
xor U3133 (N_3133,In_1181,In_528);
and U3134 (N_3134,In_1242,In_176);
nor U3135 (N_3135,In_399,In_456);
nor U3136 (N_3136,In_1153,In_956);
xor U3137 (N_3137,In_1292,In_835);
and U3138 (N_3138,In_434,In_1239);
or U3139 (N_3139,In_30,In_1148);
or U3140 (N_3140,In_888,In_1136);
xnor U3141 (N_3141,In_537,In_225);
and U3142 (N_3142,In_1359,In_454);
or U3143 (N_3143,In_1086,In_224);
nor U3144 (N_3144,In_559,In_84);
nand U3145 (N_3145,In_364,In_433);
nand U3146 (N_3146,In_1175,In_80);
nand U3147 (N_3147,In_46,In_677);
nor U3148 (N_3148,In_1094,In_696);
xnor U3149 (N_3149,In_922,In_670);
xnor U3150 (N_3150,In_1324,In_1430);
nor U3151 (N_3151,In_1267,In_359);
nor U3152 (N_3152,In_1491,In_44);
or U3153 (N_3153,In_479,In_529);
and U3154 (N_3154,In_427,In_1112);
and U3155 (N_3155,In_460,In_5);
and U3156 (N_3156,In_1197,In_622);
and U3157 (N_3157,In_713,In_487);
or U3158 (N_3158,In_1097,In_84);
or U3159 (N_3159,In_699,In_429);
nor U3160 (N_3160,In_697,In_1283);
and U3161 (N_3161,In_933,In_302);
and U3162 (N_3162,In_161,In_924);
nor U3163 (N_3163,In_407,In_1399);
xnor U3164 (N_3164,In_892,In_803);
xor U3165 (N_3165,In_267,In_270);
xnor U3166 (N_3166,In_1252,In_756);
xor U3167 (N_3167,In_107,In_523);
nand U3168 (N_3168,In_400,In_997);
nand U3169 (N_3169,In_949,In_448);
nor U3170 (N_3170,In_438,In_181);
or U3171 (N_3171,In_1166,In_1256);
or U3172 (N_3172,In_964,In_860);
xor U3173 (N_3173,In_1303,In_1208);
xnor U3174 (N_3174,In_537,In_991);
and U3175 (N_3175,In_1202,In_979);
or U3176 (N_3176,In_1465,In_231);
and U3177 (N_3177,In_896,In_677);
xnor U3178 (N_3178,In_15,In_153);
nand U3179 (N_3179,In_590,In_1283);
xnor U3180 (N_3180,In_21,In_224);
xnor U3181 (N_3181,In_18,In_966);
or U3182 (N_3182,In_1377,In_302);
nand U3183 (N_3183,In_572,In_1361);
and U3184 (N_3184,In_1084,In_73);
xnor U3185 (N_3185,In_619,In_341);
or U3186 (N_3186,In_123,In_191);
xor U3187 (N_3187,In_742,In_958);
nand U3188 (N_3188,In_1181,In_306);
xor U3189 (N_3189,In_785,In_1204);
and U3190 (N_3190,In_245,In_800);
xor U3191 (N_3191,In_787,In_366);
or U3192 (N_3192,In_318,In_472);
xnor U3193 (N_3193,In_1147,In_1050);
xnor U3194 (N_3194,In_583,In_930);
nor U3195 (N_3195,In_267,In_1020);
xor U3196 (N_3196,In_1235,In_135);
xor U3197 (N_3197,In_281,In_155);
xor U3198 (N_3198,In_501,In_1069);
nand U3199 (N_3199,In_913,In_333);
or U3200 (N_3200,In_175,In_883);
and U3201 (N_3201,In_725,In_168);
nor U3202 (N_3202,In_217,In_1304);
nor U3203 (N_3203,In_763,In_46);
nor U3204 (N_3204,In_884,In_1358);
nor U3205 (N_3205,In_1360,In_1267);
and U3206 (N_3206,In_1201,In_287);
xnor U3207 (N_3207,In_1480,In_792);
nand U3208 (N_3208,In_811,In_441);
xor U3209 (N_3209,In_1217,In_190);
xnor U3210 (N_3210,In_100,In_443);
xnor U3211 (N_3211,In_874,In_680);
nor U3212 (N_3212,In_1420,In_197);
xnor U3213 (N_3213,In_223,In_1033);
and U3214 (N_3214,In_1343,In_367);
nand U3215 (N_3215,In_677,In_479);
and U3216 (N_3216,In_837,In_870);
xnor U3217 (N_3217,In_597,In_1426);
nand U3218 (N_3218,In_739,In_890);
or U3219 (N_3219,In_1056,In_865);
xor U3220 (N_3220,In_310,In_75);
nand U3221 (N_3221,In_715,In_882);
and U3222 (N_3222,In_160,In_546);
nand U3223 (N_3223,In_184,In_138);
nor U3224 (N_3224,In_1486,In_287);
nand U3225 (N_3225,In_1074,In_10);
nand U3226 (N_3226,In_1346,In_137);
nor U3227 (N_3227,In_108,In_1468);
xor U3228 (N_3228,In_1076,In_968);
or U3229 (N_3229,In_315,In_518);
nand U3230 (N_3230,In_1461,In_83);
and U3231 (N_3231,In_1318,In_63);
nand U3232 (N_3232,In_1320,In_417);
xnor U3233 (N_3233,In_703,In_235);
and U3234 (N_3234,In_1041,In_1214);
or U3235 (N_3235,In_801,In_1192);
and U3236 (N_3236,In_52,In_1232);
nor U3237 (N_3237,In_506,In_650);
nor U3238 (N_3238,In_411,In_894);
nor U3239 (N_3239,In_1454,In_672);
nor U3240 (N_3240,In_651,In_937);
nand U3241 (N_3241,In_642,In_862);
nor U3242 (N_3242,In_124,In_1484);
or U3243 (N_3243,In_943,In_142);
nand U3244 (N_3244,In_386,In_810);
nor U3245 (N_3245,In_376,In_1029);
xnor U3246 (N_3246,In_102,In_362);
or U3247 (N_3247,In_1338,In_77);
nor U3248 (N_3248,In_642,In_1212);
nand U3249 (N_3249,In_1332,In_759);
nor U3250 (N_3250,In_770,In_339);
nand U3251 (N_3251,In_543,In_200);
xnor U3252 (N_3252,In_654,In_1318);
and U3253 (N_3253,In_340,In_454);
or U3254 (N_3254,In_1041,In_257);
nor U3255 (N_3255,In_18,In_719);
xor U3256 (N_3256,In_633,In_395);
nor U3257 (N_3257,In_846,In_1207);
or U3258 (N_3258,In_593,In_1295);
or U3259 (N_3259,In_413,In_1022);
or U3260 (N_3260,In_862,In_1417);
nand U3261 (N_3261,In_897,In_608);
xor U3262 (N_3262,In_625,In_1364);
or U3263 (N_3263,In_872,In_123);
xnor U3264 (N_3264,In_144,In_52);
or U3265 (N_3265,In_826,In_1408);
or U3266 (N_3266,In_769,In_215);
nor U3267 (N_3267,In_549,In_720);
nand U3268 (N_3268,In_213,In_698);
nor U3269 (N_3269,In_209,In_511);
nor U3270 (N_3270,In_63,In_486);
nor U3271 (N_3271,In_1405,In_1241);
nand U3272 (N_3272,In_950,In_884);
nor U3273 (N_3273,In_898,In_754);
nand U3274 (N_3274,In_681,In_1450);
and U3275 (N_3275,In_152,In_554);
and U3276 (N_3276,In_519,In_514);
and U3277 (N_3277,In_430,In_632);
and U3278 (N_3278,In_770,In_248);
nor U3279 (N_3279,In_182,In_52);
nor U3280 (N_3280,In_864,In_1089);
nand U3281 (N_3281,In_967,In_1479);
or U3282 (N_3282,In_1148,In_853);
xnor U3283 (N_3283,In_177,In_321);
nand U3284 (N_3284,In_1174,In_876);
or U3285 (N_3285,In_875,In_861);
nor U3286 (N_3286,In_176,In_621);
nor U3287 (N_3287,In_979,In_300);
nor U3288 (N_3288,In_1417,In_160);
nand U3289 (N_3289,In_351,In_627);
or U3290 (N_3290,In_1096,In_112);
nor U3291 (N_3291,In_1399,In_1042);
nand U3292 (N_3292,In_884,In_1186);
nor U3293 (N_3293,In_940,In_835);
nor U3294 (N_3294,In_1481,In_110);
or U3295 (N_3295,In_1268,In_707);
and U3296 (N_3296,In_132,In_406);
nor U3297 (N_3297,In_419,In_1145);
nor U3298 (N_3298,In_101,In_887);
or U3299 (N_3299,In_1263,In_107);
or U3300 (N_3300,In_667,In_1162);
xnor U3301 (N_3301,In_1063,In_641);
and U3302 (N_3302,In_438,In_1079);
nand U3303 (N_3303,In_570,In_988);
nor U3304 (N_3304,In_798,In_942);
and U3305 (N_3305,In_1208,In_1277);
nor U3306 (N_3306,In_1358,In_751);
nand U3307 (N_3307,In_951,In_205);
nand U3308 (N_3308,In_1319,In_1492);
xnor U3309 (N_3309,In_1314,In_375);
or U3310 (N_3310,In_44,In_806);
nand U3311 (N_3311,In_285,In_1427);
nand U3312 (N_3312,In_18,In_284);
xnor U3313 (N_3313,In_989,In_1154);
nand U3314 (N_3314,In_118,In_1262);
or U3315 (N_3315,In_1024,In_1478);
nand U3316 (N_3316,In_1168,In_1390);
xor U3317 (N_3317,In_1354,In_482);
nor U3318 (N_3318,In_8,In_454);
nand U3319 (N_3319,In_1023,In_60);
or U3320 (N_3320,In_861,In_229);
or U3321 (N_3321,In_1350,In_1025);
or U3322 (N_3322,In_1441,In_1390);
xor U3323 (N_3323,In_1108,In_714);
xor U3324 (N_3324,In_919,In_355);
nand U3325 (N_3325,In_682,In_1136);
nand U3326 (N_3326,In_107,In_358);
and U3327 (N_3327,In_87,In_558);
nor U3328 (N_3328,In_673,In_339);
or U3329 (N_3329,In_734,In_36);
xor U3330 (N_3330,In_499,In_1018);
nor U3331 (N_3331,In_675,In_1101);
and U3332 (N_3332,In_102,In_246);
nor U3333 (N_3333,In_878,In_548);
or U3334 (N_3334,In_494,In_409);
or U3335 (N_3335,In_236,In_1346);
and U3336 (N_3336,In_1368,In_1451);
nand U3337 (N_3337,In_1371,In_260);
nand U3338 (N_3338,In_71,In_1496);
xnor U3339 (N_3339,In_406,In_1278);
nand U3340 (N_3340,In_611,In_396);
xor U3341 (N_3341,In_465,In_1137);
nand U3342 (N_3342,In_912,In_875);
nand U3343 (N_3343,In_1137,In_428);
xnor U3344 (N_3344,In_884,In_1396);
nand U3345 (N_3345,In_60,In_129);
or U3346 (N_3346,In_693,In_1299);
nor U3347 (N_3347,In_893,In_114);
xor U3348 (N_3348,In_1161,In_782);
or U3349 (N_3349,In_1310,In_1232);
nor U3350 (N_3350,In_123,In_1015);
xor U3351 (N_3351,In_92,In_1298);
nor U3352 (N_3352,In_129,In_168);
and U3353 (N_3353,In_117,In_1218);
nand U3354 (N_3354,In_1182,In_853);
and U3355 (N_3355,In_39,In_188);
xnor U3356 (N_3356,In_1446,In_165);
nor U3357 (N_3357,In_15,In_905);
or U3358 (N_3358,In_765,In_1077);
or U3359 (N_3359,In_1278,In_974);
nand U3360 (N_3360,In_650,In_665);
or U3361 (N_3361,In_258,In_401);
nand U3362 (N_3362,In_697,In_559);
xor U3363 (N_3363,In_616,In_1397);
xnor U3364 (N_3364,In_587,In_999);
xor U3365 (N_3365,In_964,In_44);
nor U3366 (N_3366,In_51,In_701);
and U3367 (N_3367,In_604,In_192);
or U3368 (N_3368,In_1356,In_1150);
and U3369 (N_3369,In_981,In_792);
or U3370 (N_3370,In_100,In_591);
or U3371 (N_3371,In_916,In_525);
xor U3372 (N_3372,In_1265,In_1477);
and U3373 (N_3373,In_333,In_927);
xor U3374 (N_3374,In_456,In_264);
xnor U3375 (N_3375,In_557,In_1271);
xor U3376 (N_3376,In_1454,In_69);
and U3377 (N_3377,In_330,In_1314);
and U3378 (N_3378,In_959,In_1308);
xnor U3379 (N_3379,In_1442,In_273);
or U3380 (N_3380,In_1240,In_550);
and U3381 (N_3381,In_167,In_774);
and U3382 (N_3382,In_1120,In_1233);
xor U3383 (N_3383,In_90,In_744);
xor U3384 (N_3384,In_60,In_358);
or U3385 (N_3385,In_261,In_1071);
xnor U3386 (N_3386,In_1006,In_1486);
xnor U3387 (N_3387,In_859,In_725);
nand U3388 (N_3388,In_1198,In_126);
nor U3389 (N_3389,In_938,In_1135);
nor U3390 (N_3390,In_907,In_1323);
xor U3391 (N_3391,In_746,In_1021);
nand U3392 (N_3392,In_768,In_175);
nand U3393 (N_3393,In_1085,In_575);
nor U3394 (N_3394,In_738,In_164);
and U3395 (N_3395,In_140,In_1386);
and U3396 (N_3396,In_930,In_628);
xnor U3397 (N_3397,In_718,In_1100);
nand U3398 (N_3398,In_1482,In_1286);
and U3399 (N_3399,In_368,In_207);
xor U3400 (N_3400,In_259,In_686);
xor U3401 (N_3401,In_508,In_539);
xor U3402 (N_3402,In_567,In_625);
xor U3403 (N_3403,In_888,In_1038);
nand U3404 (N_3404,In_1077,In_35);
nor U3405 (N_3405,In_1185,In_1044);
and U3406 (N_3406,In_39,In_92);
or U3407 (N_3407,In_851,In_1173);
nand U3408 (N_3408,In_995,In_1112);
and U3409 (N_3409,In_1376,In_521);
and U3410 (N_3410,In_1046,In_496);
or U3411 (N_3411,In_88,In_984);
nor U3412 (N_3412,In_559,In_1432);
or U3413 (N_3413,In_568,In_949);
or U3414 (N_3414,In_1091,In_1062);
nand U3415 (N_3415,In_109,In_1269);
or U3416 (N_3416,In_289,In_1434);
nor U3417 (N_3417,In_313,In_647);
and U3418 (N_3418,In_1392,In_375);
or U3419 (N_3419,In_1315,In_1345);
or U3420 (N_3420,In_337,In_564);
nand U3421 (N_3421,In_454,In_83);
nand U3422 (N_3422,In_209,In_198);
xor U3423 (N_3423,In_1074,In_1217);
and U3424 (N_3424,In_568,In_473);
xor U3425 (N_3425,In_428,In_1092);
nand U3426 (N_3426,In_572,In_407);
nor U3427 (N_3427,In_756,In_27);
or U3428 (N_3428,In_959,In_107);
xor U3429 (N_3429,In_1057,In_1370);
xnor U3430 (N_3430,In_983,In_675);
nand U3431 (N_3431,In_696,In_320);
or U3432 (N_3432,In_124,In_42);
or U3433 (N_3433,In_1407,In_1135);
xor U3434 (N_3434,In_86,In_371);
xor U3435 (N_3435,In_1371,In_1184);
and U3436 (N_3436,In_776,In_1456);
and U3437 (N_3437,In_869,In_606);
and U3438 (N_3438,In_1394,In_733);
nand U3439 (N_3439,In_638,In_755);
xnor U3440 (N_3440,In_362,In_313);
nor U3441 (N_3441,In_796,In_1472);
and U3442 (N_3442,In_5,In_27);
or U3443 (N_3443,In_678,In_1275);
nor U3444 (N_3444,In_159,In_1486);
or U3445 (N_3445,In_555,In_591);
or U3446 (N_3446,In_500,In_372);
nor U3447 (N_3447,In_306,In_380);
xor U3448 (N_3448,In_1047,In_863);
or U3449 (N_3449,In_771,In_1487);
nand U3450 (N_3450,In_1394,In_403);
and U3451 (N_3451,In_1449,In_1145);
xnor U3452 (N_3452,In_204,In_1424);
xor U3453 (N_3453,In_1362,In_925);
and U3454 (N_3454,In_682,In_801);
and U3455 (N_3455,In_121,In_66);
nor U3456 (N_3456,In_929,In_432);
nor U3457 (N_3457,In_1053,In_1268);
or U3458 (N_3458,In_281,In_1235);
and U3459 (N_3459,In_493,In_1394);
xnor U3460 (N_3460,In_1331,In_508);
nor U3461 (N_3461,In_419,In_492);
and U3462 (N_3462,In_723,In_408);
nor U3463 (N_3463,In_1204,In_249);
or U3464 (N_3464,In_600,In_1053);
xnor U3465 (N_3465,In_1131,In_732);
nand U3466 (N_3466,In_398,In_1162);
and U3467 (N_3467,In_491,In_393);
and U3468 (N_3468,In_1264,In_1371);
nand U3469 (N_3469,In_1375,In_1249);
or U3470 (N_3470,In_682,In_436);
nor U3471 (N_3471,In_1165,In_1487);
nand U3472 (N_3472,In_578,In_1310);
nor U3473 (N_3473,In_318,In_1405);
or U3474 (N_3474,In_1239,In_430);
nor U3475 (N_3475,In_604,In_717);
xnor U3476 (N_3476,In_354,In_226);
or U3477 (N_3477,In_1492,In_738);
nand U3478 (N_3478,In_1203,In_430);
nand U3479 (N_3479,In_668,In_954);
nor U3480 (N_3480,In_934,In_311);
and U3481 (N_3481,In_1278,In_838);
nand U3482 (N_3482,In_754,In_1448);
and U3483 (N_3483,In_130,In_1422);
xnor U3484 (N_3484,In_1019,In_1465);
and U3485 (N_3485,In_1434,In_360);
nor U3486 (N_3486,In_207,In_130);
nand U3487 (N_3487,In_709,In_336);
nor U3488 (N_3488,In_948,In_263);
xor U3489 (N_3489,In_764,In_452);
nor U3490 (N_3490,In_546,In_490);
or U3491 (N_3491,In_1429,In_994);
and U3492 (N_3492,In_559,In_1112);
or U3493 (N_3493,In_796,In_317);
and U3494 (N_3494,In_1266,In_790);
and U3495 (N_3495,In_742,In_618);
and U3496 (N_3496,In_1105,In_339);
or U3497 (N_3497,In_159,In_950);
xnor U3498 (N_3498,In_236,In_1183);
xnor U3499 (N_3499,In_1278,In_877);
and U3500 (N_3500,In_1127,In_358);
xor U3501 (N_3501,In_1202,In_383);
xor U3502 (N_3502,In_243,In_1279);
or U3503 (N_3503,In_1393,In_59);
xnor U3504 (N_3504,In_334,In_466);
and U3505 (N_3505,In_1212,In_1452);
or U3506 (N_3506,In_1240,In_1204);
or U3507 (N_3507,In_593,In_1472);
and U3508 (N_3508,In_471,In_4);
nand U3509 (N_3509,In_554,In_511);
and U3510 (N_3510,In_421,In_132);
or U3511 (N_3511,In_947,In_632);
nand U3512 (N_3512,In_290,In_1087);
and U3513 (N_3513,In_547,In_221);
and U3514 (N_3514,In_83,In_939);
nand U3515 (N_3515,In_1274,In_1156);
or U3516 (N_3516,In_855,In_762);
xor U3517 (N_3517,In_625,In_1013);
and U3518 (N_3518,In_969,In_844);
or U3519 (N_3519,In_680,In_587);
xor U3520 (N_3520,In_1357,In_955);
nand U3521 (N_3521,In_139,In_272);
or U3522 (N_3522,In_450,In_1279);
nand U3523 (N_3523,In_1407,In_1335);
xor U3524 (N_3524,In_1380,In_1127);
xnor U3525 (N_3525,In_497,In_841);
and U3526 (N_3526,In_1286,In_581);
or U3527 (N_3527,In_435,In_162);
nand U3528 (N_3528,In_1467,In_454);
and U3529 (N_3529,In_1490,In_1452);
nor U3530 (N_3530,In_855,In_1179);
nand U3531 (N_3531,In_1170,In_752);
and U3532 (N_3532,In_1013,In_243);
or U3533 (N_3533,In_515,In_610);
xnor U3534 (N_3534,In_1073,In_691);
xnor U3535 (N_3535,In_439,In_9);
xnor U3536 (N_3536,In_836,In_1086);
nor U3537 (N_3537,In_772,In_224);
or U3538 (N_3538,In_981,In_11);
xor U3539 (N_3539,In_1260,In_1293);
nor U3540 (N_3540,In_1230,In_357);
nor U3541 (N_3541,In_264,In_1070);
nor U3542 (N_3542,In_79,In_229);
or U3543 (N_3543,In_1463,In_97);
or U3544 (N_3544,In_696,In_703);
nand U3545 (N_3545,In_472,In_713);
or U3546 (N_3546,In_1450,In_1069);
nor U3547 (N_3547,In_641,In_1245);
and U3548 (N_3548,In_115,In_1194);
or U3549 (N_3549,In_397,In_1195);
nor U3550 (N_3550,In_540,In_69);
or U3551 (N_3551,In_960,In_693);
nor U3552 (N_3552,In_1154,In_1099);
xor U3553 (N_3553,In_92,In_456);
or U3554 (N_3554,In_925,In_1156);
xor U3555 (N_3555,In_1295,In_57);
nor U3556 (N_3556,In_467,In_774);
or U3557 (N_3557,In_875,In_1050);
nor U3558 (N_3558,In_395,In_128);
and U3559 (N_3559,In_1433,In_750);
nor U3560 (N_3560,In_1328,In_1068);
or U3561 (N_3561,In_696,In_1231);
or U3562 (N_3562,In_992,In_1481);
or U3563 (N_3563,In_1468,In_83);
and U3564 (N_3564,In_119,In_70);
nor U3565 (N_3565,In_29,In_293);
and U3566 (N_3566,In_489,In_1266);
nand U3567 (N_3567,In_1434,In_1025);
and U3568 (N_3568,In_545,In_785);
xnor U3569 (N_3569,In_427,In_1035);
nand U3570 (N_3570,In_414,In_910);
or U3571 (N_3571,In_248,In_352);
or U3572 (N_3572,In_261,In_1279);
xnor U3573 (N_3573,In_1409,In_831);
nor U3574 (N_3574,In_481,In_80);
and U3575 (N_3575,In_1426,In_974);
and U3576 (N_3576,In_505,In_967);
xor U3577 (N_3577,In_65,In_1158);
and U3578 (N_3578,In_1347,In_620);
nor U3579 (N_3579,In_1054,In_467);
nand U3580 (N_3580,In_1019,In_854);
nand U3581 (N_3581,In_1270,In_39);
or U3582 (N_3582,In_49,In_983);
or U3583 (N_3583,In_751,In_338);
nor U3584 (N_3584,In_276,In_46);
and U3585 (N_3585,In_1127,In_1166);
nor U3586 (N_3586,In_282,In_1014);
and U3587 (N_3587,In_882,In_1385);
nor U3588 (N_3588,In_285,In_72);
and U3589 (N_3589,In_398,In_152);
or U3590 (N_3590,In_506,In_1013);
xor U3591 (N_3591,In_113,In_678);
and U3592 (N_3592,In_965,In_653);
nand U3593 (N_3593,In_1247,In_1459);
nand U3594 (N_3594,In_585,In_682);
nor U3595 (N_3595,In_57,In_870);
or U3596 (N_3596,In_608,In_276);
and U3597 (N_3597,In_262,In_530);
and U3598 (N_3598,In_694,In_1322);
or U3599 (N_3599,In_1187,In_1100);
nand U3600 (N_3600,In_1474,In_633);
nand U3601 (N_3601,In_72,In_777);
or U3602 (N_3602,In_855,In_1074);
nor U3603 (N_3603,In_703,In_143);
nor U3604 (N_3604,In_748,In_615);
nand U3605 (N_3605,In_959,In_1342);
nand U3606 (N_3606,In_1346,In_83);
and U3607 (N_3607,In_1340,In_1443);
nand U3608 (N_3608,In_1423,In_709);
nand U3609 (N_3609,In_465,In_623);
xnor U3610 (N_3610,In_378,In_1332);
nor U3611 (N_3611,In_367,In_512);
xor U3612 (N_3612,In_483,In_79);
or U3613 (N_3613,In_336,In_170);
nand U3614 (N_3614,In_346,In_358);
nand U3615 (N_3615,In_720,In_299);
and U3616 (N_3616,In_1499,In_423);
or U3617 (N_3617,In_96,In_1314);
xor U3618 (N_3618,In_911,In_488);
nand U3619 (N_3619,In_777,In_85);
or U3620 (N_3620,In_180,In_346);
nand U3621 (N_3621,In_974,In_1270);
or U3622 (N_3622,In_1158,In_1481);
or U3623 (N_3623,In_623,In_724);
xor U3624 (N_3624,In_1339,In_84);
nand U3625 (N_3625,In_1105,In_67);
and U3626 (N_3626,In_1355,In_1301);
xnor U3627 (N_3627,In_916,In_1083);
or U3628 (N_3628,In_1274,In_1299);
nor U3629 (N_3629,In_923,In_1369);
or U3630 (N_3630,In_439,In_494);
or U3631 (N_3631,In_1002,In_415);
nor U3632 (N_3632,In_1368,In_582);
xor U3633 (N_3633,In_924,In_1420);
nand U3634 (N_3634,In_197,In_304);
xor U3635 (N_3635,In_1076,In_887);
nor U3636 (N_3636,In_1316,In_259);
nor U3637 (N_3637,In_709,In_1441);
xor U3638 (N_3638,In_578,In_994);
and U3639 (N_3639,In_59,In_278);
and U3640 (N_3640,In_1424,In_641);
nand U3641 (N_3641,In_1264,In_210);
xor U3642 (N_3642,In_310,In_1491);
and U3643 (N_3643,In_300,In_1351);
nor U3644 (N_3644,In_1231,In_925);
or U3645 (N_3645,In_883,In_422);
nor U3646 (N_3646,In_40,In_1063);
nor U3647 (N_3647,In_1275,In_514);
nor U3648 (N_3648,In_142,In_1313);
and U3649 (N_3649,In_353,In_1230);
nor U3650 (N_3650,In_1127,In_636);
xor U3651 (N_3651,In_114,In_1195);
xnor U3652 (N_3652,In_612,In_460);
and U3653 (N_3653,In_414,In_1071);
or U3654 (N_3654,In_44,In_1479);
nor U3655 (N_3655,In_594,In_507);
and U3656 (N_3656,In_707,In_193);
xor U3657 (N_3657,In_990,In_1482);
or U3658 (N_3658,In_1466,In_81);
nor U3659 (N_3659,In_640,In_943);
or U3660 (N_3660,In_513,In_1010);
xnor U3661 (N_3661,In_1445,In_1016);
xor U3662 (N_3662,In_120,In_197);
nor U3663 (N_3663,In_614,In_780);
or U3664 (N_3664,In_1020,In_969);
and U3665 (N_3665,In_80,In_1439);
nor U3666 (N_3666,In_1250,In_892);
nor U3667 (N_3667,In_643,In_904);
and U3668 (N_3668,In_488,In_306);
or U3669 (N_3669,In_1141,In_1059);
and U3670 (N_3670,In_1496,In_435);
or U3671 (N_3671,In_385,In_408);
nand U3672 (N_3672,In_293,In_1142);
nand U3673 (N_3673,In_292,In_816);
and U3674 (N_3674,In_1271,In_553);
or U3675 (N_3675,In_1213,In_862);
xor U3676 (N_3676,In_1140,In_996);
and U3677 (N_3677,In_595,In_631);
xor U3678 (N_3678,In_802,In_750);
nand U3679 (N_3679,In_22,In_862);
nand U3680 (N_3680,In_988,In_487);
or U3681 (N_3681,In_296,In_427);
and U3682 (N_3682,In_292,In_1230);
nor U3683 (N_3683,In_1183,In_1064);
or U3684 (N_3684,In_124,In_203);
and U3685 (N_3685,In_22,In_1086);
xor U3686 (N_3686,In_279,In_1);
nand U3687 (N_3687,In_556,In_1433);
nand U3688 (N_3688,In_633,In_864);
xnor U3689 (N_3689,In_795,In_1079);
xnor U3690 (N_3690,In_1055,In_1085);
nand U3691 (N_3691,In_942,In_836);
or U3692 (N_3692,In_871,In_362);
xnor U3693 (N_3693,In_265,In_514);
nor U3694 (N_3694,In_1251,In_858);
nand U3695 (N_3695,In_22,In_721);
and U3696 (N_3696,In_93,In_119);
or U3697 (N_3697,In_607,In_958);
xor U3698 (N_3698,In_194,In_471);
and U3699 (N_3699,In_295,In_1401);
and U3700 (N_3700,In_1113,In_945);
nand U3701 (N_3701,In_442,In_1116);
nand U3702 (N_3702,In_312,In_827);
and U3703 (N_3703,In_16,In_1159);
nand U3704 (N_3704,In_757,In_845);
nor U3705 (N_3705,In_717,In_314);
and U3706 (N_3706,In_743,In_246);
xnor U3707 (N_3707,In_690,In_294);
and U3708 (N_3708,In_709,In_974);
xnor U3709 (N_3709,In_555,In_379);
or U3710 (N_3710,In_18,In_746);
nand U3711 (N_3711,In_792,In_280);
and U3712 (N_3712,In_689,In_1337);
xnor U3713 (N_3713,In_467,In_1372);
nand U3714 (N_3714,In_553,In_29);
nand U3715 (N_3715,In_683,In_444);
and U3716 (N_3716,In_674,In_1102);
nor U3717 (N_3717,In_879,In_721);
nand U3718 (N_3718,In_658,In_850);
xnor U3719 (N_3719,In_344,In_882);
xor U3720 (N_3720,In_951,In_1384);
nand U3721 (N_3721,In_357,In_1247);
nand U3722 (N_3722,In_1348,In_98);
nor U3723 (N_3723,In_945,In_1472);
xnor U3724 (N_3724,In_951,In_744);
and U3725 (N_3725,In_338,In_1466);
nand U3726 (N_3726,In_606,In_275);
or U3727 (N_3727,In_1137,In_711);
nand U3728 (N_3728,In_238,In_857);
nand U3729 (N_3729,In_424,In_1142);
and U3730 (N_3730,In_557,In_718);
nor U3731 (N_3731,In_138,In_121);
and U3732 (N_3732,In_946,In_496);
or U3733 (N_3733,In_236,In_1132);
or U3734 (N_3734,In_241,In_1139);
nor U3735 (N_3735,In_1411,In_1175);
nor U3736 (N_3736,In_1414,In_169);
and U3737 (N_3737,In_757,In_198);
nor U3738 (N_3738,In_254,In_1375);
or U3739 (N_3739,In_323,In_1018);
nor U3740 (N_3740,In_462,In_1389);
nor U3741 (N_3741,In_486,In_1230);
nor U3742 (N_3742,In_935,In_1197);
nand U3743 (N_3743,In_409,In_1050);
and U3744 (N_3744,In_979,In_314);
nand U3745 (N_3745,In_997,In_842);
nor U3746 (N_3746,In_1344,In_1469);
or U3747 (N_3747,In_931,In_707);
nand U3748 (N_3748,In_1047,In_361);
or U3749 (N_3749,In_1431,In_145);
or U3750 (N_3750,In_1109,In_1438);
nand U3751 (N_3751,In_164,In_1251);
nand U3752 (N_3752,In_296,In_1158);
xnor U3753 (N_3753,In_185,In_117);
nor U3754 (N_3754,In_795,In_715);
xnor U3755 (N_3755,In_3,In_1428);
or U3756 (N_3756,In_2,In_865);
nand U3757 (N_3757,In_88,In_677);
xor U3758 (N_3758,In_539,In_1334);
nand U3759 (N_3759,In_1489,In_1291);
and U3760 (N_3760,In_1422,In_188);
and U3761 (N_3761,In_391,In_421);
and U3762 (N_3762,In_478,In_1412);
and U3763 (N_3763,In_834,In_203);
nand U3764 (N_3764,In_443,In_1144);
nand U3765 (N_3765,In_845,In_340);
nor U3766 (N_3766,In_599,In_1166);
and U3767 (N_3767,In_426,In_946);
xor U3768 (N_3768,In_1309,In_1318);
nor U3769 (N_3769,In_538,In_203);
and U3770 (N_3770,In_780,In_67);
xor U3771 (N_3771,In_159,In_1145);
nand U3772 (N_3772,In_580,In_1254);
and U3773 (N_3773,In_442,In_280);
nand U3774 (N_3774,In_534,In_1328);
xor U3775 (N_3775,In_1303,In_290);
or U3776 (N_3776,In_10,In_392);
nor U3777 (N_3777,In_183,In_753);
or U3778 (N_3778,In_436,In_1435);
or U3779 (N_3779,In_1200,In_1208);
nor U3780 (N_3780,In_1255,In_235);
or U3781 (N_3781,In_340,In_1192);
or U3782 (N_3782,In_1001,In_1287);
nor U3783 (N_3783,In_1265,In_1458);
and U3784 (N_3784,In_836,In_445);
or U3785 (N_3785,In_128,In_1040);
xnor U3786 (N_3786,In_1130,In_692);
nor U3787 (N_3787,In_26,In_289);
and U3788 (N_3788,In_115,In_151);
nor U3789 (N_3789,In_873,In_92);
and U3790 (N_3790,In_1209,In_692);
xor U3791 (N_3791,In_913,In_135);
or U3792 (N_3792,In_85,In_1330);
xor U3793 (N_3793,In_318,In_95);
or U3794 (N_3794,In_1361,In_710);
nand U3795 (N_3795,In_376,In_57);
nand U3796 (N_3796,In_5,In_544);
and U3797 (N_3797,In_1068,In_1462);
nor U3798 (N_3798,In_260,In_991);
xnor U3799 (N_3799,In_252,In_81);
nor U3800 (N_3800,In_1451,In_791);
xnor U3801 (N_3801,In_1180,In_706);
nand U3802 (N_3802,In_149,In_380);
nor U3803 (N_3803,In_166,In_666);
xnor U3804 (N_3804,In_1205,In_14);
nand U3805 (N_3805,In_105,In_538);
nor U3806 (N_3806,In_926,In_141);
and U3807 (N_3807,In_1371,In_893);
xor U3808 (N_3808,In_1140,In_649);
xnor U3809 (N_3809,In_113,In_381);
and U3810 (N_3810,In_1386,In_1258);
and U3811 (N_3811,In_1135,In_1056);
or U3812 (N_3812,In_1269,In_394);
xor U3813 (N_3813,In_1304,In_985);
xor U3814 (N_3814,In_990,In_1393);
nor U3815 (N_3815,In_123,In_337);
xor U3816 (N_3816,In_970,In_967);
and U3817 (N_3817,In_795,In_928);
nand U3818 (N_3818,In_1029,In_1355);
nor U3819 (N_3819,In_648,In_328);
and U3820 (N_3820,In_531,In_125);
or U3821 (N_3821,In_139,In_1300);
or U3822 (N_3822,In_6,In_733);
nor U3823 (N_3823,In_1346,In_370);
xor U3824 (N_3824,In_173,In_1287);
nand U3825 (N_3825,In_1365,In_855);
nor U3826 (N_3826,In_925,In_454);
or U3827 (N_3827,In_1234,In_1196);
and U3828 (N_3828,In_312,In_285);
and U3829 (N_3829,In_1224,In_422);
or U3830 (N_3830,In_213,In_1031);
or U3831 (N_3831,In_1119,In_632);
nor U3832 (N_3832,In_1210,In_857);
nor U3833 (N_3833,In_119,In_1397);
and U3834 (N_3834,In_1300,In_1351);
or U3835 (N_3835,In_1428,In_918);
and U3836 (N_3836,In_693,In_1194);
and U3837 (N_3837,In_955,In_746);
nand U3838 (N_3838,In_287,In_1044);
xnor U3839 (N_3839,In_141,In_766);
xnor U3840 (N_3840,In_3,In_916);
nand U3841 (N_3841,In_61,In_876);
or U3842 (N_3842,In_858,In_236);
or U3843 (N_3843,In_106,In_626);
nand U3844 (N_3844,In_702,In_293);
or U3845 (N_3845,In_1013,In_1009);
nor U3846 (N_3846,In_569,In_733);
nor U3847 (N_3847,In_1193,In_298);
nor U3848 (N_3848,In_374,In_99);
or U3849 (N_3849,In_1022,In_715);
nor U3850 (N_3850,In_512,In_918);
or U3851 (N_3851,In_1072,In_164);
nand U3852 (N_3852,In_146,In_1238);
nand U3853 (N_3853,In_102,In_211);
and U3854 (N_3854,In_16,In_1325);
nand U3855 (N_3855,In_356,In_327);
nor U3856 (N_3856,In_1272,In_1065);
and U3857 (N_3857,In_875,In_119);
xnor U3858 (N_3858,In_646,In_1025);
nor U3859 (N_3859,In_428,In_396);
xor U3860 (N_3860,In_310,In_758);
nand U3861 (N_3861,In_350,In_90);
nand U3862 (N_3862,In_595,In_909);
nand U3863 (N_3863,In_260,In_1153);
xnor U3864 (N_3864,In_1008,In_631);
nand U3865 (N_3865,In_1452,In_1174);
nor U3866 (N_3866,In_945,In_295);
nand U3867 (N_3867,In_731,In_424);
xnor U3868 (N_3868,In_1405,In_812);
nand U3869 (N_3869,In_147,In_206);
xnor U3870 (N_3870,In_1402,In_559);
xnor U3871 (N_3871,In_1488,In_965);
or U3872 (N_3872,In_1473,In_59);
nand U3873 (N_3873,In_955,In_17);
or U3874 (N_3874,In_1058,In_60);
nor U3875 (N_3875,In_1076,In_688);
xor U3876 (N_3876,In_709,In_1139);
xor U3877 (N_3877,In_1479,In_1431);
xor U3878 (N_3878,In_514,In_81);
xor U3879 (N_3879,In_1428,In_1258);
nand U3880 (N_3880,In_1127,In_397);
and U3881 (N_3881,In_1179,In_1397);
and U3882 (N_3882,In_550,In_1472);
nor U3883 (N_3883,In_1441,In_1391);
nor U3884 (N_3884,In_1283,In_423);
or U3885 (N_3885,In_586,In_489);
xor U3886 (N_3886,In_867,In_944);
and U3887 (N_3887,In_358,In_1093);
or U3888 (N_3888,In_926,In_847);
xnor U3889 (N_3889,In_724,In_594);
nor U3890 (N_3890,In_833,In_952);
or U3891 (N_3891,In_121,In_267);
and U3892 (N_3892,In_680,In_798);
nand U3893 (N_3893,In_1255,In_5);
xor U3894 (N_3894,In_568,In_609);
nor U3895 (N_3895,In_1379,In_137);
and U3896 (N_3896,In_1374,In_262);
nor U3897 (N_3897,In_375,In_1207);
xor U3898 (N_3898,In_74,In_1422);
or U3899 (N_3899,In_1123,In_860);
or U3900 (N_3900,In_708,In_924);
nor U3901 (N_3901,In_657,In_1380);
nand U3902 (N_3902,In_1029,In_1303);
nor U3903 (N_3903,In_1136,In_491);
nand U3904 (N_3904,In_1069,In_379);
nor U3905 (N_3905,In_73,In_1175);
and U3906 (N_3906,In_602,In_909);
or U3907 (N_3907,In_243,In_1411);
and U3908 (N_3908,In_368,In_224);
or U3909 (N_3909,In_768,In_1289);
nor U3910 (N_3910,In_1466,In_671);
and U3911 (N_3911,In_455,In_267);
nand U3912 (N_3912,In_1230,In_647);
and U3913 (N_3913,In_971,In_1196);
or U3914 (N_3914,In_144,In_949);
or U3915 (N_3915,In_714,In_1201);
nand U3916 (N_3916,In_293,In_1153);
nor U3917 (N_3917,In_1305,In_1079);
or U3918 (N_3918,In_156,In_12);
nand U3919 (N_3919,In_1140,In_88);
and U3920 (N_3920,In_362,In_751);
nand U3921 (N_3921,In_73,In_538);
or U3922 (N_3922,In_612,In_112);
nor U3923 (N_3923,In_1071,In_847);
xor U3924 (N_3924,In_207,In_1414);
nor U3925 (N_3925,In_1439,In_494);
or U3926 (N_3926,In_655,In_1483);
and U3927 (N_3927,In_781,In_417);
and U3928 (N_3928,In_1365,In_53);
xnor U3929 (N_3929,In_1460,In_764);
nor U3930 (N_3930,In_346,In_496);
nand U3931 (N_3931,In_334,In_1225);
or U3932 (N_3932,In_163,In_543);
or U3933 (N_3933,In_655,In_213);
nor U3934 (N_3934,In_1183,In_978);
nor U3935 (N_3935,In_1057,In_1467);
nand U3936 (N_3936,In_858,In_21);
and U3937 (N_3937,In_101,In_161);
nand U3938 (N_3938,In_797,In_1159);
nor U3939 (N_3939,In_852,In_56);
nand U3940 (N_3940,In_785,In_1388);
nor U3941 (N_3941,In_326,In_587);
nand U3942 (N_3942,In_439,In_1105);
or U3943 (N_3943,In_834,In_1167);
and U3944 (N_3944,In_408,In_1227);
and U3945 (N_3945,In_1020,In_1250);
nand U3946 (N_3946,In_491,In_735);
or U3947 (N_3947,In_163,In_762);
or U3948 (N_3948,In_1426,In_745);
nor U3949 (N_3949,In_468,In_925);
nor U3950 (N_3950,In_25,In_667);
and U3951 (N_3951,In_1013,In_719);
xnor U3952 (N_3952,In_1176,In_151);
nand U3953 (N_3953,In_473,In_492);
nand U3954 (N_3954,In_976,In_893);
or U3955 (N_3955,In_153,In_1276);
xnor U3956 (N_3956,In_393,In_1214);
nand U3957 (N_3957,In_253,In_172);
and U3958 (N_3958,In_234,In_48);
nand U3959 (N_3959,In_1473,In_204);
nand U3960 (N_3960,In_740,In_504);
xnor U3961 (N_3961,In_1479,In_500);
nand U3962 (N_3962,In_958,In_3);
nand U3963 (N_3963,In_150,In_200);
or U3964 (N_3964,In_95,In_102);
nand U3965 (N_3965,In_705,In_543);
nand U3966 (N_3966,In_27,In_672);
nor U3967 (N_3967,In_1373,In_237);
and U3968 (N_3968,In_677,In_1218);
nand U3969 (N_3969,In_1105,In_666);
xnor U3970 (N_3970,In_185,In_342);
and U3971 (N_3971,In_1225,In_787);
nand U3972 (N_3972,In_539,In_126);
xnor U3973 (N_3973,In_968,In_992);
nand U3974 (N_3974,In_765,In_915);
nor U3975 (N_3975,In_806,In_514);
and U3976 (N_3976,In_434,In_1054);
nand U3977 (N_3977,In_706,In_1235);
and U3978 (N_3978,In_1064,In_1135);
nor U3979 (N_3979,In_849,In_222);
xor U3980 (N_3980,In_386,In_737);
or U3981 (N_3981,In_432,In_261);
nand U3982 (N_3982,In_72,In_1082);
nor U3983 (N_3983,In_400,In_117);
and U3984 (N_3984,In_540,In_804);
and U3985 (N_3985,In_75,In_384);
and U3986 (N_3986,In_179,In_273);
xnor U3987 (N_3987,In_73,In_412);
nand U3988 (N_3988,In_635,In_1024);
or U3989 (N_3989,In_1166,In_1367);
nor U3990 (N_3990,In_743,In_162);
or U3991 (N_3991,In_1101,In_1069);
xnor U3992 (N_3992,In_609,In_917);
nand U3993 (N_3993,In_641,In_487);
nand U3994 (N_3994,In_1092,In_672);
nor U3995 (N_3995,In_767,In_303);
xnor U3996 (N_3996,In_10,In_1077);
nor U3997 (N_3997,In_635,In_922);
nor U3998 (N_3998,In_539,In_299);
nand U3999 (N_3999,In_496,In_870);
xnor U4000 (N_4000,In_1237,In_1275);
nor U4001 (N_4001,In_989,In_959);
xnor U4002 (N_4002,In_1110,In_1006);
and U4003 (N_4003,In_115,In_1085);
nand U4004 (N_4004,In_1385,In_922);
or U4005 (N_4005,In_1089,In_1284);
nand U4006 (N_4006,In_1133,In_418);
xnor U4007 (N_4007,In_267,In_855);
and U4008 (N_4008,In_42,In_142);
nor U4009 (N_4009,In_581,In_1098);
or U4010 (N_4010,In_708,In_785);
or U4011 (N_4011,In_203,In_1481);
nand U4012 (N_4012,In_526,In_532);
or U4013 (N_4013,In_485,In_708);
nand U4014 (N_4014,In_702,In_491);
xor U4015 (N_4015,In_343,In_1487);
nor U4016 (N_4016,In_687,In_1382);
and U4017 (N_4017,In_761,In_821);
nor U4018 (N_4018,In_423,In_776);
nor U4019 (N_4019,In_1168,In_1232);
nand U4020 (N_4020,In_972,In_200);
nor U4021 (N_4021,In_601,In_533);
or U4022 (N_4022,In_1048,In_418);
xnor U4023 (N_4023,In_942,In_174);
and U4024 (N_4024,In_358,In_542);
and U4025 (N_4025,In_825,In_1151);
xor U4026 (N_4026,In_921,In_1407);
or U4027 (N_4027,In_765,In_714);
xnor U4028 (N_4028,In_1340,In_658);
xor U4029 (N_4029,In_1059,In_1120);
nor U4030 (N_4030,In_402,In_1294);
and U4031 (N_4031,In_1483,In_596);
xor U4032 (N_4032,In_203,In_828);
nand U4033 (N_4033,In_876,In_972);
nor U4034 (N_4034,In_131,In_919);
and U4035 (N_4035,In_1246,In_122);
xor U4036 (N_4036,In_68,In_1111);
xor U4037 (N_4037,In_307,In_1044);
and U4038 (N_4038,In_1247,In_365);
and U4039 (N_4039,In_1091,In_1152);
nor U4040 (N_4040,In_243,In_1260);
xor U4041 (N_4041,In_839,In_437);
nor U4042 (N_4042,In_435,In_1275);
or U4043 (N_4043,In_390,In_1108);
or U4044 (N_4044,In_1448,In_160);
or U4045 (N_4045,In_1336,In_61);
or U4046 (N_4046,In_1190,In_1230);
xnor U4047 (N_4047,In_1462,In_625);
or U4048 (N_4048,In_1354,In_416);
and U4049 (N_4049,In_768,In_688);
nor U4050 (N_4050,In_1098,In_1093);
or U4051 (N_4051,In_340,In_496);
nor U4052 (N_4052,In_48,In_1197);
xnor U4053 (N_4053,In_63,In_138);
xor U4054 (N_4054,In_679,In_637);
xor U4055 (N_4055,In_604,In_190);
or U4056 (N_4056,In_531,In_281);
nand U4057 (N_4057,In_508,In_1437);
nor U4058 (N_4058,In_471,In_860);
or U4059 (N_4059,In_243,In_1176);
nor U4060 (N_4060,In_307,In_1095);
or U4061 (N_4061,In_240,In_813);
nor U4062 (N_4062,In_508,In_258);
nor U4063 (N_4063,In_438,In_1462);
nor U4064 (N_4064,In_1326,In_1468);
xor U4065 (N_4065,In_1212,In_911);
or U4066 (N_4066,In_607,In_1245);
nor U4067 (N_4067,In_1277,In_1263);
and U4068 (N_4068,In_609,In_848);
nand U4069 (N_4069,In_1089,In_278);
nand U4070 (N_4070,In_1143,In_878);
nand U4071 (N_4071,In_1327,In_137);
or U4072 (N_4072,In_1007,In_141);
or U4073 (N_4073,In_1047,In_138);
nand U4074 (N_4074,In_1207,In_749);
and U4075 (N_4075,In_256,In_1135);
xnor U4076 (N_4076,In_413,In_242);
xor U4077 (N_4077,In_429,In_177);
nand U4078 (N_4078,In_586,In_1203);
and U4079 (N_4079,In_201,In_840);
and U4080 (N_4080,In_1314,In_48);
or U4081 (N_4081,In_826,In_177);
and U4082 (N_4082,In_883,In_1421);
nand U4083 (N_4083,In_193,In_589);
nand U4084 (N_4084,In_13,In_1225);
nand U4085 (N_4085,In_424,In_1380);
nand U4086 (N_4086,In_34,In_105);
nor U4087 (N_4087,In_401,In_194);
nand U4088 (N_4088,In_1017,In_1379);
nor U4089 (N_4089,In_967,In_720);
xor U4090 (N_4090,In_1402,In_1311);
nand U4091 (N_4091,In_14,In_745);
or U4092 (N_4092,In_41,In_320);
nor U4093 (N_4093,In_759,In_360);
xor U4094 (N_4094,In_830,In_806);
and U4095 (N_4095,In_353,In_336);
xnor U4096 (N_4096,In_74,In_883);
nand U4097 (N_4097,In_171,In_930);
nor U4098 (N_4098,In_253,In_1428);
nand U4099 (N_4099,In_553,In_662);
nand U4100 (N_4100,In_1189,In_202);
nor U4101 (N_4101,In_232,In_1261);
nand U4102 (N_4102,In_901,In_145);
nand U4103 (N_4103,In_107,In_370);
and U4104 (N_4104,In_1074,In_115);
xor U4105 (N_4105,In_1462,In_409);
xor U4106 (N_4106,In_988,In_174);
or U4107 (N_4107,In_1005,In_870);
nand U4108 (N_4108,In_1003,In_1352);
xnor U4109 (N_4109,In_273,In_357);
nor U4110 (N_4110,In_200,In_306);
or U4111 (N_4111,In_391,In_521);
nor U4112 (N_4112,In_1124,In_317);
nor U4113 (N_4113,In_1351,In_1055);
xnor U4114 (N_4114,In_1057,In_433);
nor U4115 (N_4115,In_121,In_881);
xnor U4116 (N_4116,In_1319,In_452);
and U4117 (N_4117,In_1373,In_64);
and U4118 (N_4118,In_612,In_1057);
nor U4119 (N_4119,In_591,In_363);
xor U4120 (N_4120,In_446,In_630);
nand U4121 (N_4121,In_670,In_837);
and U4122 (N_4122,In_18,In_252);
nand U4123 (N_4123,In_1331,In_429);
nor U4124 (N_4124,In_432,In_1353);
nand U4125 (N_4125,In_451,In_174);
or U4126 (N_4126,In_213,In_525);
nand U4127 (N_4127,In_1176,In_1362);
and U4128 (N_4128,In_417,In_809);
nor U4129 (N_4129,In_452,In_230);
nor U4130 (N_4130,In_1173,In_119);
xor U4131 (N_4131,In_264,In_1315);
and U4132 (N_4132,In_99,In_1081);
xnor U4133 (N_4133,In_976,In_1099);
nor U4134 (N_4134,In_869,In_457);
or U4135 (N_4135,In_757,In_181);
nand U4136 (N_4136,In_883,In_704);
xor U4137 (N_4137,In_438,In_394);
nand U4138 (N_4138,In_187,In_840);
and U4139 (N_4139,In_512,In_510);
and U4140 (N_4140,In_1171,In_352);
or U4141 (N_4141,In_307,In_1212);
or U4142 (N_4142,In_67,In_900);
nor U4143 (N_4143,In_707,In_352);
and U4144 (N_4144,In_1459,In_578);
xor U4145 (N_4145,In_367,In_1434);
nand U4146 (N_4146,In_324,In_413);
nand U4147 (N_4147,In_333,In_1278);
xor U4148 (N_4148,In_408,In_126);
nand U4149 (N_4149,In_752,In_415);
or U4150 (N_4150,In_212,In_570);
and U4151 (N_4151,In_409,In_807);
or U4152 (N_4152,In_134,In_1180);
xor U4153 (N_4153,In_241,In_1205);
xor U4154 (N_4154,In_635,In_851);
or U4155 (N_4155,In_1345,In_687);
nor U4156 (N_4156,In_123,In_124);
or U4157 (N_4157,In_450,In_769);
xnor U4158 (N_4158,In_861,In_1256);
and U4159 (N_4159,In_1423,In_296);
and U4160 (N_4160,In_1105,In_1489);
nor U4161 (N_4161,In_670,In_487);
or U4162 (N_4162,In_1121,In_601);
xor U4163 (N_4163,In_746,In_714);
nand U4164 (N_4164,In_243,In_71);
xor U4165 (N_4165,In_1219,In_1070);
nor U4166 (N_4166,In_676,In_35);
and U4167 (N_4167,In_332,In_444);
nor U4168 (N_4168,In_211,In_865);
and U4169 (N_4169,In_1124,In_249);
and U4170 (N_4170,In_1404,In_203);
and U4171 (N_4171,In_1127,In_1294);
and U4172 (N_4172,In_315,In_546);
or U4173 (N_4173,In_905,In_408);
or U4174 (N_4174,In_170,In_570);
nor U4175 (N_4175,In_1057,In_24);
nand U4176 (N_4176,In_1499,In_318);
nor U4177 (N_4177,In_1059,In_1051);
and U4178 (N_4178,In_1150,In_395);
nor U4179 (N_4179,In_510,In_81);
or U4180 (N_4180,In_905,In_470);
xor U4181 (N_4181,In_1071,In_483);
nor U4182 (N_4182,In_164,In_201);
or U4183 (N_4183,In_910,In_1151);
and U4184 (N_4184,In_390,In_934);
xor U4185 (N_4185,In_41,In_1115);
nor U4186 (N_4186,In_529,In_380);
or U4187 (N_4187,In_150,In_1198);
xnor U4188 (N_4188,In_503,In_960);
nand U4189 (N_4189,In_1174,In_1110);
xnor U4190 (N_4190,In_553,In_162);
or U4191 (N_4191,In_501,In_1170);
or U4192 (N_4192,In_1123,In_628);
and U4193 (N_4193,In_559,In_1236);
nor U4194 (N_4194,In_400,In_1063);
nand U4195 (N_4195,In_997,In_1035);
or U4196 (N_4196,In_1446,In_939);
xor U4197 (N_4197,In_1249,In_689);
and U4198 (N_4198,In_1389,In_358);
nand U4199 (N_4199,In_390,In_1103);
and U4200 (N_4200,In_154,In_1123);
nand U4201 (N_4201,In_1167,In_1057);
nor U4202 (N_4202,In_463,In_10);
or U4203 (N_4203,In_23,In_73);
or U4204 (N_4204,In_408,In_557);
nor U4205 (N_4205,In_801,In_419);
nor U4206 (N_4206,In_1116,In_904);
nor U4207 (N_4207,In_1259,In_1306);
xor U4208 (N_4208,In_377,In_716);
nand U4209 (N_4209,In_1107,In_517);
nor U4210 (N_4210,In_1456,In_1059);
or U4211 (N_4211,In_205,In_717);
or U4212 (N_4212,In_1439,In_584);
xor U4213 (N_4213,In_803,In_281);
nand U4214 (N_4214,In_382,In_251);
or U4215 (N_4215,In_1468,In_1257);
or U4216 (N_4216,In_1484,In_1227);
xor U4217 (N_4217,In_340,In_1331);
and U4218 (N_4218,In_314,In_70);
nor U4219 (N_4219,In_1352,In_1385);
or U4220 (N_4220,In_1244,In_1375);
xnor U4221 (N_4221,In_1046,In_470);
or U4222 (N_4222,In_1374,In_1426);
or U4223 (N_4223,In_139,In_429);
nand U4224 (N_4224,In_732,In_795);
and U4225 (N_4225,In_921,In_435);
nor U4226 (N_4226,In_1197,In_956);
and U4227 (N_4227,In_823,In_1288);
xor U4228 (N_4228,In_984,In_904);
nor U4229 (N_4229,In_671,In_908);
nor U4230 (N_4230,In_1239,In_19);
nand U4231 (N_4231,In_25,In_341);
xor U4232 (N_4232,In_949,In_179);
and U4233 (N_4233,In_602,In_644);
or U4234 (N_4234,In_131,In_1310);
nor U4235 (N_4235,In_789,In_917);
nor U4236 (N_4236,In_688,In_254);
nand U4237 (N_4237,In_390,In_34);
and U4238 (N_4238,In_1471,In_1009);
nand U4239 (N_4239,In_1078,In_524);
xnor U4240 (N_4240,In_279,In_988);
nand U4241 (N_4241,In_1241,In_1120);
xor U4242 (N_4242,In_590,In_840);
and U4243 (N_4243,In_1067,In_408);
or U4244 (N_4244,In_376,In_712);
nand U4245 (N_4245,In_640,In_776);
nor U4246 (N_4246,In_232,In_1394);
xor U4247 (N_4247,In_445,In_1088);
xor U4248 (N_4248,In_1149,In_134);
xor U4249 (N_4249,In_1099,In_548);
nor U4250 (N_4250,In_93,In_1285);
xnor U4251 (N_4251,In_221,In_591);
or U4252 (N_4252,In_619,In_703);
nor U4253 (N_4253,In_577,In_549);
nor U4254 (N_4254,In_84,In_1171);
nand U4255 (N_4255,In_799,In_888);
and U4256 (N_4256,In_257,In_380);
xor U4257 (N_4257,In_1044,In_148);
or U4258 (N_4258,In_1202,In_1257);
nor U4259 (N_4259,In_815,In_1480);
and U4260 (N_4260,In_1439,In_627);
xnor U4261 (N_4261,In_643,In_126);
nor U4262 (N_4262,In_1041,In_932);
or U4263 (N_4263,In_1324,In_311);
or U4264 (N_4264,In_249,In_1141);
xnor U4265 (N_4265,In_21,In_1181);
nand U4266 (N_4266,In_107,In_393);
or U4267 (N_4267,In_613,In_160);
xor U4268 (N_4268,In_755,In_676);
nand U4269 (N_4269,In_560,In_451);
xor U4270 (N_4270,In_554,In_1031);
xor U4271 (N_4271,In_1083,In_983);
and U4272 (N_4272,In_542,In_725);
xnor U4273 (N_4273,In_1049,In_434);
nor U4274 (N_4274,In_569,In_476);
xnor U4275 (N_4275,In_573,In_1269);
and U4276 (N_4276,In_1128,In_1257);
or U4277 (N_4277,In_1287,In_1260);
or U4278 (N_4278,In_280,In_586);
and U4279 (N_4279,In_1275,In_625);
nor U4280 (N_4280,In_1186,In_1334);
and U4281 (N_4281,In_991,In_874);
xor U4282 (N_4282,In_175,In_230);
nor U4283 (N_4283,In_47,In_1444);
or U4284 (N_4284,In_671,In_827);
nor U4285 (N_4285,In_1409,In_1115);
nand U4286 (N_4286,In_1001,In_1115);
nor U4287 (N_4287,In_1322,In_356);
or U4288 (N_4288,In_282,In_212);
nor U4289 (N_4289,In_1192,In_920);
and U4290 (N_4290,In_1350,In_59);
and U4291 (N_4291,In_21,In_3);
nor U4292 (N_4292,In_516,In_414);
nand U4293 (N_4293,In_1435,In_1338);
and U4294 (N_4294,In_1034,In_808);
nor U4295 (N_4295,In_134,In_780);
xnor U4296 (N_4296,In_663,In_542);
nor U4297 (N_4297,In_1204,In_1324);
and U4298 (N_4298,In_209,In_725);
nand U4299 (N_4299,In_193,In_1022);
and U4300 (N_4300,In_475,In_1162);
or U4301 (N_4301,In_1342,In_607);
and U4302 (N_4302,In_1079,In_374);
and U4303 (N_4303,In_375,In_167);
nor U4304 (N_4304,In_422,In_235);
nor U4305 (N_4305,In_1473,In_1236);
xor U4306 (N_4306,In_1305,In_1426);
and U4307 (N_4307,In_764,In_1056);
nor U4308 (N_4308,In_415,In_30);
and U4309 (N_4309,In_1461,In_380);
and U4310 (N_4310,In_992,In_1401);
nand U4311 (N_4311,In_215,In_1093);
or U4312 (N_4312,In_857,In_756);
nand U4313 (N_4313,In_1195,In_975);
xor U4314 (N_4314,In_102,In_66);
or U4315 (N_4315,In_1310,In_1131);
nor U4316 (N_4316,In_717,In_1346);
and U4317 (N_4317,In_574,In_920);
or U4318 (N_4318,In_449,In_5);
nand U4319 (N_4319,In_1000,In_675);
nand U4320 (N_4320,In_82,In_929);
and U4321 (N_4321,In_966,In_195);
and U4322 (N_4322,In_1160,In_583);
or U4323 (N_4323,In_382,In_106);
nand U4324 (N_4324,In_1448,In_1422);
nand U4325 (N_4325,In_112,In_402);
and U4326 (N_4326,In_1290,In_195);
or U4327 (N_4327,In_147,In_1296);
nand U4328 (N_4328,In_963,In_1254);
nand U4329 (N_4329,In_1484,In_973);
nand U4330 (N_4330,In_1267,In_950);
or U4331 (N_4331,In_922,In_195);
xnor U4332 (N_4332,In_1046,In_951);
xor U4333 (N_4333,In_929,In_1081);
nand U4334 (N_4334,In_63,In_651);
nor U4335 (N_4335,In_415,In_1040);
or U4336 (N_4336,In_626,In_885);
nor U4337 (N_4337,In_1093,In_1392);
xor U4338 (N_4338,In_1206,In_1257);
nor U4339 (N_4339,In_414,In_300);
and U4340 (N_4340,In_35,In_41);
nand U4341 (N_4341,In_123,In_613);
xor U4342 (N_4342,In_1105,In_282);
or U4343 (N_4343,In_270,In_1336);
nor U4344 (N_4344,In_312,In_341);
nor U4345 (N_4345,In_357,In_1433);
xnor U4346 (N_4346,In_1429,In_865);
nor U4347 (N_4347,In_848,In_404);
and U4348 (N_4348,In_56,In_851);
nand U4349 (N_4349,In_1218,In_566);
and U4350 (N_4350,In_865,In_416);
or U4351 (N_4351,In_641,In_994);
xor U4352 (N_4352,In_1454,In_913);
nor U4353 (N_4353,In_874,In_1300);
nor U4354 (N_4354,In_465,In_442);
nand U4355 (N_4355,In_38,In_348);
nand U4356 (N_4356,In_801,In_249);
nor U4357 (N_4357,In_860,In_703);
or U4358 (N_4358,In_393,In_120);
or U4359 (N_4359,In_1114,In_1266);
xnor U4360 (N_4360,In_1344,In_536);
xnor U4361 (N_4361,In_136,In_1322);
xor U4362 (N_4362,In_151,In_1293);
nor U4363 (N_4363,In_349,In_503);
and U4364 (N_4364,In_995,In_912);
or U4365 (N_4365,In_720,In_928);
xnor U4366 (N_4366,In_1335,In_787);
nand U4367 (N_4367,In_1333,In_1015);
and U4368 (N_4368,In_713,In_1303);
xnor U4369 (N_4369,In_928,In_1209);
nand U4370 (N_4370,In_426,In_1139);
xnor U4371 (N_4371,In_448,In_406);
nand U4372 (N_4372,In_1452,In_1191);
nor U4373 (N_4373,In_1239,In_1156);
nor U4374 (N_4374,In_756,In_70);
nor U4375 (N_4375,In_1106,In_690);
nand U4376 (N_4376,In_223,In_1035);
nand U4377 (N_4377,In_464,In_1142);
xor U4378 (N_4378,In_260,In_343);
nor U4379 (N_4379,In_830,In_1212);
nand U4380 (N_4380,In_623,In_575);
and U4381 (N_4381,In_875,In_652);
xor U4382 (N_4382,In_598,In_988);
nor U4383 (N_4383,In_124,In_1466);
xnor U4384 (N_4384,In_1284,In_1132);
or U4385 (N_4385,In_1361,In_916);
or U4386 (N_4386,In_1233,In_852);
xor U4387 (N_4387,In_697,In_67);
nor U4388 (N_4388,In_1096,In_470);
and U4389 (N_4389,In_1119,In_635);
or U4390 (N_4390,In_203,In_613);
xnor U4391 (N_4391,In_555,In_999);
nor U4392 (N_4392,In_1323,In_142);
nor U4393 (N_4393,In_1496,In_313);
or U4394 (N_4394,In_144,In_1232);
or U4395 (N_4395,In_198,In_224);
xnor U4396 (N_4396,In_1373,In_215);
or U4397 (N_4397,In_97,In_113);
and U4398 (N_4398,In_110,In_864);
or U4399 (N_4399,In_983,In_169);
nand U4400 (N_4400,In_489,In_620);
and U4401 (N_4401,In_718,In_1293);
nor U4402 (N_4402,In_1149,In_1427);
nand U4403 (N_4403,In_481,In_1445);
and U4404 (N_4404,In_81,In_1354);
xnor U4405 (N_4405,In_853,In_867);
nand U4406 (N_4406,In_705,In_185);
and U4407 (N_4407,In_1245,In_552);
and U4408 (N_4408,In_478,In_776);
nand U4409 (N_4409,In_316,In_306);
or U4410 (N_4410,In_811,In_1451);
nor U4411 (N_4411,In_1380,In_792);
nor U4412 (N_4412,In_1363,In_199);
and U4413 (N_4413,In_868,In_1311);
nand U4414 (N_4414,In_1246,In_1015);
xor U4415 (N_4415,In_190,In_336);
nand U4416 (N_4416,In_1473,In_461);
nor U4417 (N_4417,In_1180,In_315);
nand U4418 (N_4418,In_101,In_988);
xor U4419 (N_4419,In_92,In_536);
nand U4420 (N_4420,In_879,In_650);
or U4421 (N_4421,In_675,In_1059);
and U4422 (N_4422,In_41,In_901);
and U4423 (N_4423,In_161,In_16);
xnor U4424 (N_4424,In_818,In_626);
and U4425 (N_4425,In_1478,In_539);
xor U4426 (N_4426,In_518,In_1477);
xor U4427 (N_4427,In_1132,In_1474);
and U4428 (N_4428,In_433,In_1007);
and U4429 (N_4429,In_359,In_204);
nor U4430 (N_4430,In_101,In_923);
nor U4431 (N_4431,In_1371,In_701);
xor U4432 (N_4432,In_1498,In_293);
xnor U4433 (N_4433,In_1070,In_60);
and U4434 (N_4434,In_514,In_21);
nor U4435 (N_4435,In_222,In_1073);
or U4436 (N_4436,In_1211,In_1297);
xor U4437 (N_4437,In_914,In_419);
nor U4438 (N_4438,In_1233,In_1005);
or U4439 (N_4439,In_317,In_206);
nand U4440 (N_4440,In_158,In_881);
nand U4441 (N_4441,In_226,In_702);
xor U4442 (N_4442,In_988,In_462);
nor U4443 (N_4443,In_584,In_794);
nor U4444 (N_4444,In_475,In_1384);
xnor U4445 (N_4445,In_914,In_136);
and U4446 (N_4446,In_389,In_255);
nor U4447 (N_4447,In_719,In_1455);
xor U4448 (N_4448,In_279,In_158);
and U4449 (N_4449,In_462,In_197);
nand U4450 (N_4450,In_897,In_1086);
or U4451 (N_4451,In_1051,In_390);
or U4452 (N_4452,In_135,In_625);
and U4453 (N_4453,In_941,In_853);
nand U4454 (N_4454,In_241,In_797);
xnor U4455 (N_4455,In_1002,In_1152);
xor U4456 (N_4456,In_954,In_205);
xor U4457 (N_4457,In_599,In_51);
xor U4458 (N_4458,In_1416,In_448);
or U4459 (N_4459,In_1201,In_1236);
or U4460 (N_4460,In_1404,In_76);
and U4461 (N_4461,In_981,In_1344);
xor U4462 (N_4462,In_110,In_139);
and U4463 (N_4463,In_917,In_1185);
or U4464 (N_4464,In_454,In_1238);
xnor U4465 (N_4465,In_500,In_523);
nand U4466 (N_4466,In_1410,In_1254);
nor U4467 (N_4467,In_1375,In_1167);
nand U4468 (N_4468,In_347,In_1266);
and U4469 (N_4469,In_409,In_1318);
and U4470 (N_4470,In_1148,In_83);
nor U4471 (N_4471,In_482,In_155);
xnor U4472 (N_4472,In_281,In_1030);
nand U4473 (N_4473,In_836,In_312);
or U4474 (N_4474,In_1128,In_701);
nand U4475 (N_4475,In_657,In_1383);
nand U4476 (N_4476,In_118,In_179);
nor U4477 (N_4477,In_1351,In_1430);
and U4478 (N_4478,In_223,In_1188);
and U4479 (N_4479,In_148,In_416);
nand U4480 (N_4480,In_126,In_1020);
and U4481 (N_4481,In_252,In_1175);
nor U4482 (N_4482,In_589,In_1059);
and U4483 (N_4483,In_769,In_678);
nand U4484 (N_4484,In_1413,In_204);
and U4485 (N_4485,In_408,In_450);
and U4486 (N_4486,In_1492,In_660);
and U4487 (N_4487,In_1208,In_519);
xor U4488 (N_4488,In_1493,In_374);
or U4489 (N_4489,In_1030,In_453);
nand U4490 (N_4490,In_1012,In_380);
and U4491 (N_4491,In_176,In_611);
nor U4492 (N_4492,In_661,In_627);
nand U4493 (N_4493,In_148,In_536);
nor U4494 (N_4494,In_322,In_362);
or U4495 (N_4495,In_271,In_126);
and U4496 (N_4496,In_622,In_882);
or U4497 (N_4497,In_582,In_996);
or U4498 (N_4498,In_1261,In_812);
nor U4499 (N_4499,In_824,In_805);
or U4500 (N_4500,In_786,In_1066);
and U4501 (N_4501,In_632,In_80);
and U4502 (N_4502,In_467,In_677);
nand U4503 (N_4503,In_593,In_87);
nor U4504 (N_4504,In_1459,In_219);
and U4505 (N_4505,In_568,In_219);
and U4506 (N_4506,In_610,In_90);
nand U4507 (N_4507,In_822,In_466);
nand U4508 (N_4508,In_92,In_994);
or U4509 (N_4509,In_308,In_322);
or U4510 (N_4510,In_1042,In_693);
nand U4511 (N_4511,In_1441,In_25);
nor U4512 (N_4512,In_123,In_242);
nand U4513 (N_4513,In_626,In_634);
or U4514 (N_4514,In_1435,In_563);
nor U4515 (N_4515,In_67,In_917);
nor U4516 (N_4516,In_1376,In_522);
and U4517 (N_4517,In_821,In_407);
xnor U4518 (N_4518,In_238,In_811);
xor U4519 (N_4519,In_101,In_320);
nand U4520 (N_4520,In_986,In_1249);
nor U4521 (N_4521,In_609,In_1081);
xor U4522 (N_4522,In_153,In_442);
nor U4523 (N_4523,In_1120,In_756);
nand U4524 (N_4524,In_317,In_554);
nor U4525 (N_4525,In_383,In_326);
nor U4526 (N_4526,In_188,In_638);
and U4527 (N_4527,In_1190,In_51);
or U4528 (N_4528,In_856,In_1333);
xnor U4529 (N_4529,In_939,In_588);
nor U4530 (N_4530,In_48,In_859);
or U4531 (N_4531,In_1243,In_1425);
and U4532 (N_4532,In_534,In_265);
nand U4533 (N_4533,In_399,In_595);
xor U4534 (N_4534,In_1473,In_575);
nand U4535 (N_4535,In_816,In_209);
and U4536 (N_4536,In_314,In_779);
or U4537 (N_4537,In_814,In_103);
and U4538 (N_4538,In_101,In_225);
xor U4539 (N_4539,In_530,In_172);
or U4540 (N_4540,In_1021,In_731);
and U4541 (N_4541,In_1225,In_531);
nor U4542 (N_4542,In_650,In_1177);
and U4543 (N_4543,In_490,In_436);
xor U4544 (N_4544,In_1488,In_1020);
or U4545 (N_4545,In_235,In_603);
and U4546 (N_4546,In_983,In_442);
nand U4547 (N_4547,In_799,In_701);
xnor U4548 (N_4548,In_4,In_146);
nor U4549 (N_4549,In_320,In_711);
and U4550 (N_4550,In_998,In_452);
xnor U4551 (N_4551,In_931,In_1260);
nor U4552 (N_4552,In_1314,In_1476);
and U4553 (N_4553,In_294,In_1209);
nand U4554 (N_4554,In_1084,In_26);
nor U4555 (N_4555,In_574,In_1467);
xnor U4556 (N_4556,In_1300,In_632);
nor U4557 (N_4557,In_752,In_1391);
or U4558 (N_4558,In_356,In_126);
or U4559 (N_4559,In_38,In_1091);
xnor U4560 (N_4560,In_1440,In_1057);
and U4561 (N_4561,In_798,In_1282);
xor U4562 (N_4562,In_612,In_998);
or U4563 (N_4563,In_546,In_1397);
xor U4564 (N_4564,In_871,In_82);
nor U4565 (N_4565,In_1040,In_386);
and U4566 (N_4566,In_1477,In_1416);
xor U4567 (N_4567,In_238,In_1045);
or U4568 (N_4568,In_371,In_390);
and U4569 (N_4569,In_294,In_1254);
xnor U4570 (N_4570,In_77,In_480);
or U4571 (N_4571,In_1413,In_827);
xnor U4572 (N_4572,In_42,In_532);
nand U4573 (N_4573,In_931,In_12);
and U4574 (N_4574,In_1066,In_1080);
or U4575 (N_4575,In_378,In_1129);
xnor U4576 (N_4576,In_684,In_1030);
and U4577 (N_4577,In_1491,In_1002);
nor U4578 (N_4578,In_1298,In_1267);
nor U4579 (N_4579,In_1154,In_811);
xnor U4580 (N_4580,In_862,In_328);
nor U4581 (N_4581,In_324,In_119);
nor U4582 (N_4582,In_1440,In_1381);
nand U4583 (N_4583,In_817,In_834);
xnor U4584 (N_4584,In_842,In_1281);
and U4585 (N_4585,In_941,In_760);
xor U4586 (N_4586,In_963,In_1312);
or U4587 (N_4587,In_1357,In_1490);
or U4588 (N_4588,In_513,In_1223);
and U4589 (N_4589,In_214,In_44);
nor U4590 (N_4590,In_890,In_185);
or U4591 (N_4591,In_556,In_1491);
nand U4592 (N_4592,In_553,In_172);
and U4593 (N_4593,In_56,In_967);
nor U4594 (N_4594,In_121,In_1019);
nor U4595 (N_4595,In_1192,In_817);
nand U4596 (N_4596,In_437,In_898);
and U4597 (N_4597,In_1154,In_988);
or U4598 (N_4598,In_1436,In_659);
nor U4599 (N_4599,In_888,In_606);
nand U4600 (N_4600,In_196,In_937);
xnor U4601 (N_4601,In_319,In_250);
nand U4602 (N_4602,In_825,In_1421);
nand U4603 (N_4603,In_379,In_505);
nor U4604 (N_4604,In_1322,In_643);
and U4605 (N_4605,In_1132,In_1497);
nor U4606 (N_4606,In_1361,In_484);
xnor U4607 (N_4607,In_673,In_727);
or U4608 (N_4608,In_635,In_424);
nand U4609 (N_4609,In_920,In_18);
or U4610 (N_4610,In_1052,In_431);
and U4611 (N_4611,In_1466,In_781);
nand U4612 (N_4612,In_106,In_595);
or U4613 (N_4613,In_1122,In_517);
nor U4614 (N_4614,In_553,In_1006);
or U4615 (N_4615,In_248,In_1182);
and U4616 (N_4616,In_174,In_227);
or U4617 (N_4617,In_1332,In_1040);
or U4618 (N_4618,In_1193,In_867);
nand U4619 (N_4619,In_291,In_25);
or U4620 (N_4620,In_398,In_465);
xnor U4621 (N_4621,In_498,In_1318);
xnor U4622 (N_4622,In_258,In_621);
xor U4623 (N_4623,In_1446,In_574);
and U4624 (N_4624,In_774,In_640);
and U4625 (N_4625,In_1111,In_1299);
or U4626 (N_4626,In_584,In_606);
nor U4627 (N_4627,In_1235,In_431);
nor U4628 (N_4628,In_772,In_748);
nand U4629 (N_4629,In_173,In_885);
xnor U4630 (N_4630,In_752,In_1444);
xor U4631 (N_4631,In_431,In_819);
and U4632 (N_4632,In_223,In_235);
nand U4633 (N_4633,In_895,In_216);
xor U4634 (N_4634,In_223,In_1481);
nand U4635 (N_4635,In_759,In_726);
and U4636 (N_4636,In_964,In_762);
nor U4637 (N_4637,In_1068,In_651);
or U4638 (N_4638,In_998,In_299);
or U4639 (N_4639,In_691,In_1094);
xnor U4640 (N_4640,In_1021,In_1059);
and U4641 (N_4641,In_205,In_1412);
nor U4642 (N_4642,In_1148,In_823);
and U4643 (N_4643,In_572,In_1356);
nor U4644 (N_4644,In_1424,In_740);
xor U4645 (N_4645,In_563,In_1446);
and U4646 (N_4646,In_1381,In_1353);
nor U4647 (N_4647,In_749,In_631);
or U4648 (N_4648,In_500,In_549);
and U4649 (N_4649,In_1183,In_233);
xnor U4650 (N_4650,In_169,In_180);
xor U4651 (N_4651,In_210,In_312);
and U4652 (N_4652,In_640,In_331);
or U4653 (N_4653,In_352,In_431);
nor U4654 (N_4654,In_1414,In_38);
xnor U4655 (N_4655,In_863,In_29);
or U4656 (N_4656,In_411,In_773);
nand U4657 (N_4657,In_1361,In_707);
nor U4658 (N_4658,In_384,In_78);
nor U4659 (N_4659,In_178,In_300);
nor U4660 (N_4660,In_479,In_880);
or U4661 (N_4661,In_1470,In_39);
xnor U4662 (N_4662,In_127,In_1458);
nand U4663 (N_4663,In_860,In_1134);
nor U4664 (N_4664,In_983,In_247);
nand U4665 (N_4665,In_306,In_1496);
nor U4666 (N_4666,In_365,In_39);
or U4667 (N_4667,In_456,In_28);
nor U4668 (N_4668,In_599,In_561);
nor U4669 (N_4669,In_33,In_673);
and U4670 (N_4670,In_8,In_727);
nand U4671 (N_4671,In_1029,In_1375);
xnor U4672 (N_4672,In_740,In_856);
xnor U4673 (N_4673,In_206,In_561);
nand U4674 (N_4674,In_242,In_537);
or U4675 (N_4675,In_733,In_594);
nand U4676 (N_4676,In_1142,In_90);
nand U4677 (N_4677,In_598,In_278);
xnor U4678 (N_4678,In_1378,In_358);
xor U4679 (N_4679,In_88,In_751);
nor U4680 (N_4680,In_1272,In_1189);
xor U4681 (N_4681,In_307,In_433);
xor U4682 (N_4682,In_676,In_764);
and U4683 (N_4683,In_751,In_764);
nand U4684 (N_4684,In_318,In_81);
nor U4685 (N_4685,In_1250,In_570);
and U4686 (N_4686,In_250,In_1034);
and U4687 (N_4687,In_605,In_748);
or U4688 (N_4688,In_1410,In_889);
and U4689 (N_4689,In_1090,In_183);
or U4690 (N_4690,In_137,In_485);
nand U4691 (N_4691,In_1309,In_262);
nand U4692 (N_4692,In_770,In_667);
or U4693 (N_4693,In_918,In_519);
and U4694 (N_4694,In_209,In_170);
and U4695 (N_4695,In_1126,In_414);
xnor U4696 (N_4696,In_357,In_713);
and U4697 (N_4697,In_102,In_1332);
nor U4698 (N_4698,In_173,In_1145);
xnor U4699 (N_4699,In_201,In_1392);
or U4700 (N_4700,In_1090,In_1194);
xor U4701 (N_4701,In_364,In_1092);
or U4702 (N_4702,In_1341,In_687);
or U4703 (N_4703,In_1015,In_1179);
nand U4704 (N_4704,In_82,In_608);
xor U4705 (N_4705,In_1112,In_878);
nand U4706 (N_4706,In_1079,In_1482);
xnor U4707 (N_4707,In_7,In_1275);
and U4708 (N_4708,In_158,In_98);
or U4709 (N_4709,In_481,In_134);
nand U4710 (N_4710,In_804,In_1243);
and U4711 (N_4711,In_997,In_351);
nand U4712 (N_4712,In_396,In_1147);
or U4713 (N_4713,In_938,In_1430);
nand U4714 (N_4714,In_1057,In_425);
and U4715 (N_4715,In_498,In_151);
or U4716 (N_4716,In_1349,In_961);
nor U4717 (N_4717,In_1227,In_283);
nand U4718 (N_4718,In_531,In_475);
nor U4719 (N_4719,In_216,In_1074);
nor U4720 (N_4720,In_851,In_1402);
xor U4721 (N_4721,In_799,In_161);
xor U4722 (N_4722,In_730,In_442);
nand U4723 (N_4723,In_1450,In_32);
xor U4724 (N_4724,In_1160,In_88);
xnor U4725 (N_4725,In_1041,In_966);
nor U4726 (N_4726,In_93,In_450);
nand U4727 (N_4727,In_111,In_504);
xnor U4728 (N_4728,In_767,In_136);
nor U4729 (N_4729,In_1256,In_384);
nor U4730 (N_4730,In_47,In_713);
and U4731 (N_4731,In_1156,In_453);
nand U4732 (N_4732,In_815,In_678);
xnor U4733 (N_4733,In_634,In_897);
nor U4734 (N_4734,In_720,In_10);
xnor U4735 (N_4735,In_400,In_829);
and U4736 (N_4736,In_848,In_646);
xnor U4737 (N_4737,In_398,In_25);
nand U4738 (N_4738,In_1475,In_473);
or U4739 (N_4739,In_293,In_96);
nor U4740 (N_4740,In_50,In_176);
xor U4741 (N_4741,In_1011,In_854);
or U4742 (N_4742,In_887,In_1230);
xnor U4743 (N_4743,In_1349,In_1106);
xnor U4744 (N_4744,In_365,In_990);
nand U4745 (N_4745,In_342,In_496);
or U4746 (N_4746,In_9,In_290);
nor U4747 (N_4747,In_316,In_989);
nand U4748 (N_4748,In_656,In_250);
or U4749 (N_4749,In_1271,In_1475);
xnor U4750 (N_4750,In_40,In_177);
and U4751 (N_4751,In_1152,In_932);
xor U4752 (N_4752,In_869,In_1071);
xor U4753 (N_4753,In_624,In_575);
or U4754 (N_4754,In_300,In_521);
nand U4755 (N_4755,In_1388,In_1296);
nor U4756 (N_4756,In_1407,In_1254);
nor U4757 (N_4757,In_1262,In_558);
or U4758 (N_4758,In_99,In_1350);
nor U4759 (N_4759,In_817,In_11);
or U4760 (N_4760,In_873,In_671);
and U4761 (N_4761,In_511,In_345);
nor U4762 (N_4762,In_5,In_827);
and U4763 (N_4763,In_17,In_781);
and U4764 (N_4764,In_1052,In_942);
or U4765 (N_4765,In_9,In_1377);
nor U4766 (N_4766,In_1085,In_1326);
nor U4767 (N_4767,In_1099,In_255);
nor U4768 (N_4768,In_601,In_836);
nor U4769 (N_4769,In_549,In_880);
nand U4770 (N_4770,In_81,In_673);
nand U4771 (N_4771,In_460,In_1129);
xnor U4772 (N_4772,In_572,In_530);
and U4773 (N_4773,In_124,In_945);
nand U4774 (N_4774,In_1418,In_1379);
or U4775 (N_4775,In_809,In_240);
or U4776 (N_4776,In_617,In_184);
or U4777 (N_4777,In_232,In_351);
or U4778 (N_4778,In_1154,In_1480);
nand U4779 (N_4779,In_1076,In_1311);
xnor U4780 (N_4780,In_731,In_95);
and U4781 (N_4781,In_971,In_1010);
or U4782 (N_4782,In_138,In_793);
nand U4783 (N_4783,In_603,In_428);
or U4784 (N_4784,In_992,In_778);
nor U4785 (N_4785,In_1046,In_76);
or U4786 (N_4786,In_1189,In_416);
xor U4787 (N_4787,In_304,In_512);
nand U4788 (N_4788,In_535,In_405);
nand U4789 (N_4789,In_1335,In_1274);
nor U4790 (N_4790,In_1411,In_578);
xor U4791 (N_4791,In_675,In_849);
nor U4792 (N_4792,In_590,In_649);
or U4793 (N_4793,In_547,In_434);
or U4794 (N_4794,In_491,In_1300);
xnor U4795 (N_4795,In_1051,In_735);
nor U4796 (N_4796,In_271,In_964);
nor U4797 (N_4797,In_615,In_1150);
xnor U4798 (N_4798,In_675,In_258);
xnor U4799 (N_4799,In_63,In_812);
nand U4800 (N_4800,In_50,In_119);
nand U4801 (N_4801,In_1467,In_240);
xor U4802 (N_4802,In_73,In_640);
and U4803 (N_4803,In_166,In_125);
or U4804 (N_4804,In_500,In_816);
nor U4805 (N_4805,In_1158,In_1002);
nand U4806 (N_4806,In_1147,In_32);
nor U4807 (N_4807,In_226,In_1350);
nand U4808 (N_4808,In_518,In_1446);
xor U4809 (N_4809,In_292,In_1499);
nand U4810 (N_4810,In_850,In_1060);
nor U4811 (N_4811,In_507,In_519);
or U4812 (N_4812,In_363,In_1337);
or U4813 (N_4813,In_354,In_1401);
nand U4814 (N_4814,In_1485,In_249);
or U4815 (N_4815,In_1043,In_1361);
or U4816 (N_4816,In_493,In_386);
or U4817 (N_4817,In_1321,In_9);
xor U4818 (N_4818,In_556,In_1016);
nor U4819 (N_4819,In_1327,In_784);
nand U4820 (N_4820,In_438,In_550);
and U4821 (N_4821,In_80,In_1040);
or U4822 (N_4822,In_362,In_532);
or U4823 (N_4823,In_958,In_726);
nand U4824 (N_4824,In_889,In_339);
nor U4825 (N_4825,In_1321,In_1105);
and U4826 (N_4826,In_571,In_627);
xnor U4827 (N_4827,In_590,In_960);
xor U4828 (N_4828,In_144,In_1095);
nor U4829 (N_4829,In_391,In_212);
and U4830 (N_4830,In_595,In_253);
or U4831 (N_4831,In_1262,In_726);
and U4832 (N_4832,In_320,In_69);
nand U4833 (N_4833,In_5,In_945);
nor U4834 (N_4834,In_645,In_996);
or U4835 (N_4835,In_882,In_1106);
nor U4836 (N_4836,In_1069,In_807);
nand U4837 (N_4837,In_562,In_229);
xor U4838 (N_4838,In_840,In_446);
nand U4839 (N_4839,In_1309,In_504);
nand U4840 (N_4840,In_1070,In_1159);
xor U4841 (N_4841,In_309,In_817);
nor U4842 (N_4842,In_1409,In_619);
xnor U4843 (N_4843,In_1157,In_1153);
and U4844 (N_4844,In_1306,In_1207);
nor U4845 (N_4845,In_1417,In_1182);
xnor U4846 (N_4846,In_496,In_22);
and U4847 (N_4847,In_903,In_667);
nand U4848 (N_4848,In_1390,In_1269);
or U4849 (N_4849,In_882,In_1057);
and U4850 (N_4850,In_495,In_66);
and U4851 (N_4851,In_696,In_1349);
nand U4852 (N_4852,In_921,In_1309);
nand U4853 (N_4853,In_1306,In_1180);
xnor U4854 (N_4854,In_153,In_21);
nand U4855 (N_4855,In_396,In_594);
or U4856 (N_4856,In_1348,In_459);
xor U4857 (N_4857,In_1140,In_447);
xnor U4858 (N_4858,In_1209,In_247);
xor U4859 (N_4859,In_1239,In_1493);
nor U4860 (N_4860,In_1323,In_385);
xnor U4861 (N_4861,In_356,In_120);
nor U4862 (N_4862,In_389,In_103);
nand U4863 (N_4863,In_1260,In_1345);
nor U4864 (N_4864,In_665,In_483);
xnor U4865 (N_4865,In_1020,In_1235);
or U4866 (N_4866,In_746,In_1277);
and U4867 (N_4867,In_600,In_347);
xnor U4868 (N_4868,In_884,In_1204);
or U4869 (N_4869,In_896,In_835);
nor U4870 (N_4870,In_48,In_194);
nand U4871 (N_4871,In_386,In_1222);
nor U4872 (N_4872,In_364,In_795);
nand U4873 (N_4873,In_692,In_1195);
xnor U4874 (N_4874,In_1096,In_1219);
nand U4875 (N_4875,In_835,In_1165);
nor U4876 (N_4876,In_1185,In_737);
and U4877 (N_4877,In_1111,In_999);
xnor U4878 (N_4878,In_1085,In_483);
nor U4879 (N_4879,In_1400,In_1272);
nor U4880 (N_4880,In_485,In_170);
nor U4881 (N_4881,In_1077,In_889);
or U4882 (N_4882,In_1182,In_505);
or U4883 (N_4883,In_1360,In_945);
or U4884 (N_4884,In_284,In_926);
nor U4885 (N_4885,In_915,In_1467);
nand U4886 (N_4886,In_1226,In_953);
nor U4887 (N_4887,In_1265,In_429);
nand U4888 (N_4888,In_857,In_635);
or U4889 (N_4889,In_1335,In_1413);
nand U4890 (N_4890,In_954,In_597);
nor U4891 (N_4891,In_12,In_1266);
xor U4892 (N_4892,In_314,In_597);
or U4893 (N_4893,In_720,In_387);
xor U4894 (N_4894,In_286,In_607);
nand U4895 (N_4895,In_865,In_202);
xnor U4896 (N_4896,In_438,In_1129);
or U4897 (N_4897,In_330,In_46);
or U4898 (N_4898,In_1045,In_1278);
and U4899 (N_4899,In_1058,In_189);
xnor U4900 (N_4900,In_20,In_311);
nand U4901 (N_4901,In_733,In_959);
or U4902 (N_4902,In_736,In_1285);
nand U4903 (N_4903,In_181,In_1433);
and U4904 (N_4904,In_643,In_139);
xor U4905 (N_4905,In_1437,In_771);
nand U4906 (N_4906,In_516,In_63);
nor U4907 (N_4907,In_288,In_1158);
nand U4908 (N_4908,In_408,In_239);
nand U4909 (N_4909,In_1337,In_731);
or U4910 (N_4910,In_1452,In_1128);
nand U4911 (N_4911,In_1112,In_593);
and U4912 (N_4912,In_255,In_1073);
xnor U4913 (N_4913,In_1149,In_201);
nand U4914 (N_4914,In_914,In_712);
or U4915 (N_4915,In_1102,In_1228);
and U4916 (N_4916,In_1065,In_950);
xor U4917 (N_4917,In_623,In_923);
nor U4918 (N_4918,In_1320,In_400);
nand U4919 (N_4919,In_300,In_98);
nand U4920 (N_4920,In_1215,In_942);
nand U4921 (N_4921,In_549,In_1304);
or U4922 (N_4922,In_407,In_508);
or U4923 (N_4923,In_1235,In_1408);
xnor U4924 (N_4924,In_655,In_913);
xor U4925 (N_4925,In_1342,In_1469);
nand U4926 (N_4926,In_873,In_115);
and U4927 (N_4927,In_716,In_685);
and U4928 (N_4928,In_306,In_82);
or U4929 (N_4929,In_986,In_674);
nor U4930 (N_4930,In_969,In_519);
nand U4931 (N_4931,In_758,In_124);
and U4932 (N_4932,In_1389,In_1231);
nand U4933 (N_4933,In_283,In_1458);
nor U4934 (N_4934,In_265,In_363);
and U4935 (N_4935,In_1227,In_1215);
nor U4936 (N_4936,In_1224,In_1078);
and U4937 (N_4937,In_1303,In_1247);
nand U4938 (N_4938,In_724,In_763);
xnor U4939 (N_4939,In_1462,In_103);
or U4940 (N_4940,In_543,In_360);
and U4941 (N_4941,In_1080,In_422);
nor U4942 (N_4942,In_34,In_214);
or U4943 (N_4943,In_1490,In_1333);
nor U4944 (N_4944,In_1267,In_433);
xor U4945 (N_4945,In_20,In_416);
xnor U4946 (N_4946,In_767,In_68);
or U4947 (N_4947,In_954,In_75);
nand U4948 (N_4948,In_511,In_159);
and U4949 (N_4949,In_1239,In_64);
nand U4950 (N_4950,In_548,In_867);
and U4951 (N_4951,In_467,In_1207);
nand U4952 (N_4952,In_771,In_580);
nand U4953 (N_4953,In_20,In_1322);
and U4954 (N_4954,In_911,In_1077);
nand U4955 (N_4955,In_1149,In_1414);
xnor U4956 (N_4956,In_497,In_865);
nand U4957 (N_4957,In_1317,In_1406);
xor U4958 (N_4958,In_1201,In_857);
and U4959 (N_4959,In_197,In_165);
and U4960 (N_4960,In_1438,In_867);
or U4961 (N_4961,In_507,In_186);
nor U4962 (N_4962,In_1466,In_1095);
and U4963 (N_4963,In_33,In_1490);
xnor U4964 (N_4964,In_541,In_271);
xnor U4965 (N_4965,In_1203,In_74);
nor U4966 (N_4966,In_1000,In_546);
xnor U4967 (N_4967,In_20,In_762);
nor U4968 (N_4968,In_1103,In_613);
xnor U4969 (N_4969,In_1452,In_264);
nand U4970 (N_4970,In_1368,In_736);
and U4971 (N_4971,In_140,In_1377);
nand U4972 (N_4972,In_86,In_590);
and U4973 (N_4973,In_517,In_556);
xnor U4974 (N_4974,In_863,In_1087);
nand U4975 (N_4975,In_1160,In_956);
nand U4976 (N_4976,In_1454,In_1160);
xnor U4977 (N_4977,In_465,In_1402);
nand U4978 (N_4978,In_1387,In_1176);
or U4979 (N_4979,In_8,In_779);
xor U4980 (N_4980,In_4,In_1152);
nand U4981 (N_4981,In_454,In_1468);
and U4982 (N_4982,In_226,In_980);
nor U4983 (N_4983,In_1174,In_67);
or U4984 (N_4984,In_651,In_94);
nor U4985 (N_4985,In_886,In_1363);
nand U4986 (N_4986,In_1496,In_609);
nand U4987 (N_4987,In_792,In_1487);
xnor U4988 (N_4988,In_146,In_251);
nor U4989 (N_4989,In_675,In_642);
nor U4990 (N_4990,In_168,In_569);
nand U4991 (N_4991,In_1437,In_124);
nand U4992 (N_4992,In_1147,In_247);
nor U4993 (N_4993,In_1098,In_901);
xnor U4994 (N_4994,In_189,In_337);
nor U4995 (N_4995,In_118,In_343);
and U4996 (N_4996,In_323,In_833);
or U4997 (N_4997,In_707,In_880);
nand U4998 (N_4998,In_933,In_351);
xor U4999 (N_4999,In_788,In_765);
or U5000 (N_5000,N_3384,N_2711);
or U5001 (N_5001,N_2264,N_1090);
or U5002 (N_5002,N_3195,N_2072);
and U5003 (N_5003,N_195,N_4049);
xnor U5004 (N_5004,N_2993,N_3930);
xor U5005 (N_5005,N_429,N_2874);
xor U5006 (N_5006,N_4705,N_4568);
nor U5007 (N_5007,N_2346,N_536);
and U5008 (N_5008,N_20,N_3322);
and U5009 (N_5009,N_1037,N_4021);
or U5010 (N_5010,N_887,N_4753);
xor U5011 (N_5011,N_3943,N_2922);
nor U5012 (N_5012,N_3077,N_285);
nor U5013 (N_5013,N_4279,N_4143);
and U5014 (N_5014,N_3196,N_2706);
or U5015 (N_5015,N_317,N_315);
and U5016 (N_5016,N_2165,N_4740);
xor U5017 (N_5017,N_1135,N_1381);
or U5018 (N_5018,N_1171,N_4541);
nor U5019 (N_5019,N_2750,N_4357);
xor U5020 (N_5020,N_2998,N_4323);
and U5021 (N_5021,N_3640,N_2379);
xor U5022 (N_5022,N_2593,N_2898);
or U5023 (N_5023,N_724,N_279);
and U5024 (N_5024,N_3344,N_3897);
and U5025 (N_5025,N_2584,N_561);
or U5026 (N_5026,N_2642,N_2661);
xnor U5027 (N_5027,N_2068,N_2562);
nor U5028 (N_5028,N_3790,N_3236);
xor U5029 (N_5029,N_380,N_1344);
nor U5030 (N_5030,N_2697,N_3899);
xnor U5031 (N_5031,N_636,N_731);
and U5032 (N_5032,N_4310,N_2401);
and U5033 (N_5033,N_3405,N_218);
xor U5034 (N_5034,N_1146,N_2591);
and U5035 (N_5035,N_4627,N_4221);
and U5036 (N_5036,N_1737,N_3389);
and U5037 (N_5037,N_4561,N_3581);
nor U5038 (N_5038,N_3850,N_2933);
or U5039 (N_5039,N_3979,N_3048);
and U5040 (N_5040,N_3717,N_35);
xnor U5041 (N_5041,N_4304,N_4379);
xor U5042 (N_5042,N_314,N_600);
or U5043 (N_5043,N_1831,N_2995);
nor U5044 (N_5044,N_4138,N_2365);
and U5045 (N_5045,N_3354,N_4471);
or U5046 (N_5046,N_2159,N_4378);
xnor U5047 (N_5047,N_995,N_3295);
or U5048 (N_5048,N_1361,N_2716);
or U5049 (N_5049,N_2429,N_957);
nand U5050 (N_5050,N_2280,N_4124);
nand U5051 (N_5051,N_2219,N_2960);
and U5052 (N_5052,N_4792,N_3661);
nor U5053 (N_5053,N_1981,N_4558);
xnor U5054 (N_5054,N_1845,N_5);
nand U5055 (N_5055,N_4178,N_2534);
xnor U5056 (N_5056,N_955,N_1385);
or U5057 (N_5057,N_4983,N_1157);
nand U5058 (N_5058,N_900,N_3006);
nor U5059 (N_5059,N_2251,N_3134);
nand U5060 (N_5060,N_3728,N_333);
xor U5061 (N_5061,N_1024,N_3506);
xor U5062 (N_5062,N_2778,N_4673);
nor U5063 (N_5063,N_562,N_1996);
nor U5064 (N_5064,N_719,N_794);
nor U5065 (N_5065,N_654,N_4522);
nand U5066 (N_5066,N_3151,N_2845);
xor U5067 (N_5067,N_3992,N_4847);
and U5068 (N_5068,N_4903,N_3066);
or U5069 (N_5069,N_1322,N_1722);
nor U5070 (N_5070,N_4523,N_4490);
nor U5071 (N_5071,N_4638,N_175);
and U5072 (N_5072,N_30,N_4102);
nor U5073 (N_5073,N_2693,N_2980);
nor U5074 (N_5074,N_350,N_1680);
or U5075 (N_5075,N_4395,N_1364);
or U5076 (N_5076,N_3218,N_3181);
xnor U5077 (N_5077,N_4327,N_4537);
nor U5078 (N_5078,N_1213,N_1732);
xor U5079 (N_5079,N_2824,N_4668);
and U5080 (N_5080,N_2094,N_993);
nor U5081 (N_5081,N_786,N_1711);
xor U5082 (N_5082,N_4877,N_795);
or U5083 (N_5083,N_2924,N_1321);
and U5084 (N_5084,N_3032,N_3141);
or U5085 (N_5085,N_2905,N_868);
nand U5086 (N_5086,N_1353,N_4087);
xnor U5087 (N_5087,N_3488,N_4857);
nand U5088 (N_5088,N_3906,N_1820);
xnor U5089 (N_5089,N_3272,N_4804);
nor U5090 (N_5090,N_2830,N_2673);
nand U5091 (N_5091,N_4631,N_3783);
nand U5092 (N_5092,N_284,N_4070);
xor U5093 (N_5093,N_3241,N_2698);
and U5094 (N_5094,N_891,N_3363);
or U5095 (N_5095,N_3797,N_2321);
and U5096 (N_5096,N_158,N_1744);
or U5097 (N_5097,N_4272,N_1021);
nand U5098 (N_5098,N_730,N_3705);
and U5099 (N_5099,N_4113,N_3338);
nor U5100 (N_5100,N_3306,N_2794);
nor U5101 (N_5101,N_4636,N_163);
xor U5102 (N_5102,N_4476,N_3185);
nor U5103 (N_5103,N_1745,N_3013);
xnor U5104 (N_5104,N_2383,N_3682);
and U5105 (N_5105,N_1788,N_4012);
or U5106 (N_5106,N_3620,N_3558);
nand U5107 (N_5107,N_4534,N_601);
or U5108 (N_5108,N_1500,N_1446);
or U5109 (N_5109,N_3672,N_906);
and U5110 (N_5110,N_1221,N_2236);
nor U5111 (N_5111,N_4083,N_3975);
nand U5112 (N_5112,N_301,N_3646);
and U5113 (N_5113,N_680,N_1645);
xnor U5114 (N_5114,N_2293,N_260);
and U5115 (N_5115,N_3105,N_1257);
or U5116 (N_5116,N_3745,N_3670);
nand U5117 (N_5117,N_1931,N_381);
or U5118 (N_5118,N_4757,N_3980);
nor U5119 (N_5119,N_3974,N_963);
or U5120 (N_5120,N_366,N_1735);
xor U5121 (N_5121,N_4684,N_2532);
nand U5122 (N_5122,N_3959,N_4620);
and U5123 (N_5123,N_3978,N_119);
nor U5124 (N_5124,N_2399,N_1556);
and U5125 (N_5125,N_1856,N_1489);
or U5126 (N_5126,N_2074,N_3464);
xor U5127 (N_5127,N_2719,N_3101);
or U5128 (N_5128,N_4639,N_4502);
xor U5129 (N_5129,N_1466,N_1463);
nand U5130 (N_5130,N_1816,N_3103);
xor U5131 (N_5131,N_1461,N_4036);
nand U5132 (N_5132,N_2731,N_1895);
nor U5133 (N_5133,N_3376,N_3845);
or U5134 (N_5134,N_3886,N_3550);
xor U5135 (N_5135,N_432,N_2469);
and U5136 (N_5136,N_2690,N_2179);
xor U5137 (N_5137,N_4082,N_340);
nand U5138 (N_5138,N_2595,N_2917);
and U5139 (N_5139,N_4866,N_3518);
or U5140 (N_5140,N_2248,N_3178);
nand U5141 (N_5141,N_378,N_3860);
xnor U5142 (N_5142,N_2212,N_2783);
xnor U5143 (N_5143,N_1633,N_2678);
nor U5144 (N_5144,N_3069,N_1081);
nand U5145 (N_5145,N_4459,N_2742);
nor U5146 (N_5146,N_4403,N_1799);
or U5147 (N_5147,N_3958,N_4826);
nand U5148 (N_5148,N_3410,N_3666);
and U5149 (N_5149,N_1209,N_620);
xor U5150 (N_5150,N_4597,N_2220);
and U5151 (N_5151,N_2530,N_2686);
or U5152 (N_5152,N_1302,N_3623);
or U5153 (N_5153,N_166,N_4010);
nand U5154 (N_5154,N_2826,N_4692);
nor U5155 (N_5155,N_3075,N_759);
xnor U5156 (N_5156,N_3079,N_2700);
or U5157 (N_5157,N_4299,N_3483);
xnor U5158 (N_5158,N_4019,N_3356);
nor U5159 (N_5159,N_31,N_3380);
and U5160 (N_5160,N_421,N_1934);
and U5161 (N_5161,N_313,N_4691);
and U5162 (N_5162,N_1005,N_4090);
xor U5163 (N_5163,N_1587,N_1049);
nor U5164 (N_5164,N_1476,N_38);
and U5165 (N_5165,N_4142,N_1204);
xor U5166 (N_5166,N_2022,N_4086);
xor U5167 (N_5167,N_3276,N_836);
or U5168 (N_5168,N_1100,N_2127);
and U5169 (N_5169,N_3509,N_3005);
xnor U5170 (N_5170,N_1399,N_275);
nor U5171 (N_5171,N_3073,N_981);
nand U5172 (N_5172,N_318,N_739);
xnor U5173 (N_5173,N_170,N_1250);
or U5174 (N_5174,N_856,N_3443);
nor U5175 (N_5175,N_2345,N_2364);
and U5176 (N_5176,N_1297,N_4423);
xnor U5177 (N_5177,N_4202,N_3910);
and U5178 (N_5178,N_2134,N_2785);
xnor U5179 (N_5179,N_2173,N_977);
xor U5180 (N_5180,N_576,N_2822);
xnor U5181 (N_5181,N_3765,N_2440);
nand U5182 (N_5182,N_1042,N_2156);
and U5183 (N_5183,N_2950,N_3258);
nand U5184 (N_5184,N_1583,N_3733);
nor U5185 (N_5185,N_1129,N_4650);
nor U5186 (N_5186,N_2192,N_3251);
and U5187 (N_5187,N_2758,N_4456);
nand U5188 (N_5188,N_3018,N_1498);
nand U5189 (N_5189,N_3789,N_550);
nor U5190 (N_5190,N_2654,N_3610);
xor U5191 (N_5191,N_3952,N_3097);
nand U5192 (N_5192,N_779,N_2234);
and U5193 (N_5193,N_25,N_2491);
nand U5194 (N_5194,N_3613,N_3822);
and U5195 (N_5195,N_4210,N_1695);
xnor U5196 (N_5196,N_4472,N_3901);
xnor U5197 (N_5197,N_2850,N_2210);
nor U5198 (N_5198,N_4024,N_3222);
or U5199 (N_5199,N_2131,N_1315);
nor U5200 (N_5200,N_2827,N_4811);
xnor U5201 (N_5201,N_2232,N_1697);
nand U5202 (N_5202,N_2724,N_1442);
or U5203 (N_5203,N_2277,N_4176);
or U5204 (N_5204,N_2789,N_4418);
xnor U5205 (N_5205,N_4728,N_2615);
nor U5206 (N_5206,N_2093,N_4628);
nand U5207 (N_5207,N_2389,N_2921);
nor U5208 (N_5208,N_3233,N_3047);
and U5209 (N_5209,N_2835,N_7);
nor U5210 (N_5210,N_1174,N_3428);
nand U5211 (N_5211,N_1231,N_920);
nand U5212 (N_5212,N_3763,N_3183);
and U5213 (N_5213,N_683,N_2253);
xor U5214 (N_5214,N_396,N_2624);
and U5215 (N_5215,N_4428,N_1601);
nor U5216 (N_5216,N_1771,N_4509);
and U5217 (N_5217,N_865,N_3779);
or U5218 (N_5218,N_1626,N_2553);
and U5219 (N_5219,N_4578,N_802);
or U5220 (N_5220,N_455,N_1062);
and U5221 (N_5221,N_3283,N_3751);
and U5222 (N_5222,N_4247,N_160);
xnor U5223 (N_5223,N_3811,N_104);
or U5224 (N_5224,N_2559,N_1598);
nand U5225 (N_5225,N_477,N_3571);
or U5226 (N_5226,N_1483,N_2753);
xnor U5227 (N_5227,N_4998,N_3863);
xnor U5228 (N_5228,N_1294,N_4575);
nor U5229 (N_5229,N_3612,N_4625);
nor U5230 (N_5230,N_2167,N_354);
and U5231 (N_5231,N_2186,N_2392);
and U5232 (N_5232,N_253,N_4035);
nor U5233 (N_5233,N_1911,N_3522);
xnor U5234 (N_5234,N_1496,N_4583);
nand U5235 (N_5235,N_3089,N_4548);
and U5236 (N_5236,N_2618,N_2676);
nand U5237 (N_5237,N_659,N_4121);
xnor U5238 (N_5238,N_1909,N_126);
or U5239 (N_5239,N_94,N_1266);
nor U5240 (N_5240,N_4220,N_4413);
xnor U5241 (N_5241,N_996,N_1517);
nand U5242 (N_5242,N_488,N_1712);
xor U5243 (N_5243,N_3003,N_3374);
and U5244 (N_5244,N_1210,N_2302);
and U5245 (N_5245,N_1640,N_4164);
xnor U5246 (N_5246,N_328,N_1165);
xor U5247 (N_5247,N_2235,N_4656);
nor U5248 (N_5248,N_2291,N_596);
nor U5249 (N_5249,N_3814,N_3752);
nand U5250 (N_5250,N_2195,N_699);
or U5251 (N_5251,N_1980,N_3259);
xor U5252 (N_5252,N_2350,N_4557);
xor U5253 (N_5253,N_293,N_2701);
nand U5254 (N_5254,N_3216,N_1577);
or U5255 (N_5255,N_3228,N_70);
nor U5256 (N_5256,N_1110,N_3621);
nor U5257 (N_5257,N_3526,N_4935);
and U5258 (N_5258,N_2851,N_1958);
xor U5259 (N_5259,N_1143,N_1201);
nand U5260 (N_5260,N_2151,N_1362);
and U5261 (N_5261,N_4081,N_1020);
xnor U5262 (N_5262,N_1460,N_1904);
nor U5263 (N_5263,N_4298,N_376);
nor U5264 (N_5264,N_803,N_3207);
and U5265 (N_5265,N_619,N_4053);
nand U5266 (N_5266,N_1064,N_2437);
or U5267 (N_5267,N_4078,N_113);
and U5268 (N_5268,N_4050,N_2953);
xor U5269 (N_5269,N_608,N_2837);
xor U5270 (N_5270,N_4865,N_4189);
or U5271 (N_5271,N_4363,N_1739);
and U5272 (N_5272,N_147,N_4501);
nor U5273 (N_5273,N_2144,N_1566);
nor U5274 (N_5274,N_4590,N_2010);
nand U5275 (N_5275,N_3144,N_4308);
or U5276 (N_5276,N_1670,N_3026);
nand U5277 (N_5277,N_2986,N_2397);
nor U5278 (N_5278,N_952,N_3277);
nand U5279 (N_5279,N_3595,N_3279);
and U5280 (N_5280,N_760,N_3377);
nand U5281 (N_5281,N_2160,N_1124);
or U5282 (N_5282,N_2800,N_232);
or U5283 (N_5283,N_484,N_1096);
or U5284 (N_5284,N_1555,N_764);
nor U5285 (N_5285,N_4980,N_4514);
and U5286 (N_5286,N_983,N_1159);
or U5287 (N_5287,N_4497,N_1795);
nor U5288 (N_5288,N_3962,N_4790);
nand U5289 (N_5289,N_3677,N_1557);
xor U5290 (N_5290,N_2752,N_4201);
or U5291 (N_5291,N_2527,N_2871);
nand U5292 (N_5292,N_4416,N_4007);
and U5293 (N_5293,N_3579,N_2001);
nand U5294 (N_5294,N_2660,N_2883);
nand U5295 (N_5295,N_4856,N_4487);
nand U5296 (N_5296,N_3017,N_3611);
nor U5297 (N_5297,N_4533,N_2428);
or U5298 (N_5298,N_4169,N_801);
nor U5299 (N_5299,N_1563,N_2971);
and U5300 (N_5300,N_1436,N_2645);
xnor U5301 (N_5301,N_1793,N_583);
nor U5302 (N_5302,N_1969,N_1979);
nand U5303 (N_5303,N_4372,N_1782);
and U5304 (N_5304,N_4984,N_4799);
nand U5305 (N_5305,N_676,N_448);
or U5306 (N_5306,N_4745,N_325);
nand U5307 (N_5307,N_3656,N_2322);
and U5308 (N_5308,N_1060,N_471);
and U5309 (N_5309,N_4347,N_4491);
nand U5310 (N_5310,N_3205,N_308);
or U5311 (N_5311,N_2154,N_1593);
or U5312 (N_5312,N_3999,N_1237);
and U5313 (N_5313,N_4971,N_1681);
and U5314 (N_5314,N_1805,N_2565);
or U5315 (N_5315,N_4688,N_1083);
nand U5316 (N_5316,N_1335,N_614);
xor U5317 (N_5317,N_4311,N_1242);
nor U5318 (N_5318,N_77,N_2536);
and U5319 (N_5319,N_2882,N_2092);
nand U5320 (N_5320,N_2569,N_951);
xor U5321 (N_5321,N_3986,N_4851);
nor U5322 (N_5322,N_2393,N_1840);
nor U5323 (N_5323,N_4982,N_1740);
nor U5324 (N_5324,N_1903,N_3419);
nor U5325 (N_5325,N_1731,N_3572);
xor U5326 (N_5326,N_4239,N_280);
xor U5327 (N_5327,N_2992,N_2643);
xnor U5328 (N_5328,N_1723,N_332);
and U5329 (N_5329,N_2852,N_1669);
and U5330 (N_5330,N_224,N_986);
xor U5331 (N_5331,N_3480,N_4446);
xor U5332 (N_5332,N_4276,N_4011);
nor U5333 (N_5333,N_846,N_3415);
nor U5334 (N_5334,N_4062,N_2190);
xor U5335 (N_5335,N_2604,N_682);
xor U5336 (N_5336,N_4188,N_4879);
and U5337 (N_5337,N_978,N_3361);
or U5338 (N_5338,N_4634,N_1486);
and U5339 (N_5339,N_3747,N_2175);
xnor U5340 (N_5340,N_729,N_3099);
and U5341 (N_5341,N_2630,N_1071);
nor U5342 (N_5342,N_2290,N_3859);
nor U5343 (N_5343,N_2453,N_1419);
nand U5344 (N_5344,N_973,N_2255);
and U5345 (N_5345,N_3785,N_706);
nand U5346 (N_5346,N_3022,N_1571);
xnor U5347 (N_5347,N_3898,N_844);
nor U5348 (N_5348,N_1116,N_3395);
or U5349 (N_5349,N_3761,N_3114);
nand U5350 (N_5350,N_2132,N_1404);
nor U5351 (N_5351,N_1865,N_3867);
nand U5352 (N_5352,N_3812,N_341);
and U5353 (N_5353,N_4333,N_4251);
nor U5354 (N_5354,N_1401,N_4810);
and U5355 (N_5355,N_3176,N_3919);
nand U5356 (N_5356,N_921,N_1298);
and U5357 (N_5357,N_409,N_1727);
nor U5358 (N_5358,N_1313,N_3918);
and U5359 (N_5359,N_932,N_1445);
xnor U5360 (N_5360,N_1178,N_2537);
nand U5361 (N_5361,N_2454,N_3868);
nor U5362 (N_5362,N_2340,N_3051);
xnor U5363 (N_5363,N_2408,N_3208);
or U5364 (N_5364,N_945,N_1161);
xor U5365 (N_5365,N_511,N_3594);
or U5366 (N_5366,N_1120,N_1708);
or U5367 (N_5367,N_1869,N_1447);
or U5368 (N_5368,N_1273,N_4726);
and U5369 (N_5369,N_1539,N_4618);
nand U5370 (N_5370,N_2046,N_3976);
and U5371 (N_5371,N_2973,N_221);
or U5372 (N_5372,N_3225,N_1839);
or U5373 (N_5373,N_4889,N_1113);
nor U5374 (N_5374,N_2861,N_3448);
or U5375 (N_5375,N_3268,N_3365);
nand U5376 (N_5376,N_4848,N_2567);
nand U5377 (N_5377,N_2647,N_2841);
nor U5378 (N_5378,N_1554,N_3358);
xnor U5379 (N_5379,N_1057,N_4773);
xor U5380 (N_5380,N_2014,N_211);
nand U5381 (N_5381,N_1716,N_4965);
nor U5382 (N_5382,N_2972,N_813);
xnor U5383 (N_5383,N_3138,N_753);
or U5384 (N_5384,N_871,N_1776);
xor U5385 (N_5385,N_288,N_3062);
or U5386 (N_5386,N_3854,N_2448);
nor U5387 (N_5387,N_1785,N_2941);
and U5388 (N_5388,N_3929,N_3177);
nand U5389 (N_5389,N_2402,N_1860);
nor U5390 (N_5390,N_1179,N_884);
and U5391 (N_5391,N_3755,N_2796);
and U5392 (N_5392,N_1614,N_3346);
nand U5393 (N_5393,N_3536,N_1078);
nor U5394 (N_5394,N_1373,N_466);
and U5395 (N_5395,N_2182,N_3500);
nand U5396 (N_5396,N_4182,N_4447);
or U5397 (N_5397,N_58,N_4140);
nor U5398 (N_5398,N_3564,N_4064);
xnor U5399 (N_5399,N_1293,N_540);
xor U5400 (N_5400,N_2064,N_2418);
nor U5401 (N_5401,N_1928,N_537);
nor U5402 (N_5402,N_1874,N_4479);
or U5403 (N_5403,N_3239,N_640);
xor U5404 (N_5404,N_4316,N_524);
nand U5405 (N_5405,N_4626,N_1537);
or U5406 (N_5406,N_1147,N_2396);
xnor U5407 (N_5407,N_3645,N_2033);
nor U5408 (N_5408,N_1925,N_1278);
or U5409 (N_5409,N_2136,N_1522);
xor U5410 (N_5410,N_1764,N_1133);
and U5411 (N_5411,N_3406,N_2879);
nand U5412 (N_5412,N_343,N_176);
nand U5413 (N_5413,N_2327,N_4269);
xnor U5414 (N_5414,N_3457,N_2114);
and U5415 (N_5415,N_323,N_2400);
nand U5416 (N_5416,N_2073,N_24);
nand U5417 (N_5417,N_4351,N_3340);
nand U5418 (N_5418,N_3983,N_1248);
nor U5419 (N_5419,N_1198,N_3529);
or U5420 (N_5420,N_1365,N_3553);
nor U5421 (N_5421,N_112,N_198);
xnor U5422 (N_5422,N_2909,N_4645);
nor U5423 (N_5423,N_4813,N_252);
or U5424 (N_5424,N_1093,N_4573);
nand U5425 (N_5425,N_3997,N_1121);
and U5426 (N_5426,N_179,N_2557);
nor U5427 (N_5427,N_1249,N_2207);
and U5428 (N_5428,N_2709,N_3701);
xor U5429 (N_5429,N_4567,N_3556);
and U5430 (N_5430,N_1948,N_3709);
nand U5431 (N_5431,N_2564,N_1741);
nand U5432 (N_5432,N_1425,N_505);
or U5433 (N_5433,N_2859,N_2463);
nand U5434 (N_5434,N_2875,N_1949);
nor U5435 (N_5435,N_234,N_3189);
nor U5436 (N_5436,N_1424,N_1524);
or U5437 (N_5437,N_1913,N_3890);
and U5438 (N_5438,N_577,N_4074);
xnor U5439 (N_5439,N_1151,N_4886);
nor U5440 (N_5440,N_2482,N_2518);
and U5441 (N_5441,N_2629,N_2801);
and U5442 (N_5442,N_2413,N_2081);
nor U5443 (N_5443,N_4382,N_3209);
xor U5444 (N_5444,N_1039,N_3647);
and U5445 (N_5445,N_2158,N_4037);
nor U5446 (N_5446,N_1761,N_4766);
nand U5447 (N_5447,N_3343,N_4366);
xor U5448 (N_5448,N_4485,N_2666);
or U5449 (N_5449,N_3160,N_4655);
nor U5450 (N_5450,N_2581,N_2024);
nand U5451 (N_5451,N_3425,N_3582);
xor U5452 (N_5452,N_4966,N_4559);
nor U5453 (N_5453,N_4540,N_1503);
nor U5454 (N_5454,N_3324,N_901);
xnor U5455 (N_5455,N_4171,N_3631);
or U5456 (N_5456,N_1068,N_3896);
or U5457 (N_5457,N_1619,N_1666);
xor U5458 (N_5458,N_4819,N_656);
and U5459 (N_5459,N_1644,N_860);
or U5460 (N_5460,N_1420,N_804);
and U5461 (N_5461,N_2884,N_4274);
xor U5462 (N_5462,N_2423,N_4112);
xor U5463 (N_5463,N_4949,N_1809);
nor U5464 (N_5464,N_1216,N_3862);
nor U5465 (N_5465,N_4008,N_1907);
xor U5466 (N_5466,N_127,N_4675);
and U5467 (N_5467,N_4392,N_2942);
xor U5468 (N_5468,N_2049,N_2109);
or U5469 (N_5469,N_4929,N_1513);
nor U5470 (N_5470,N_2747,N_2237);
or U5471 (N_5471,N_3087,N_2004);
and U5472 (N_5472,N_383,N_437);
nor U5473 (N_5473,N_3262,N_10);
or U5474 (N_5474,N_1826,N_1596);
nand U5475 (N_5475,N_3155,N_387);
xnor U5476 (N_5476,N_3378,N_3469);
and U5477 (N_5477,N_4611,N_2163);
nor U5478 (N_5478,N_3815,N_4069);
or U5479 (N_5479,N_922,N_4187);
nand U5480 (N_5480,N_2620,N_3221);
xnor U5481 (N_5481,N_1218,N_1457);
and U5482 (N_5482,N_4077,N_721);
nor U5483 (N_5483,N_2477,N_1128);
xnor U5484 (N_5484,N_230,N_2543);
xnor U5485 (N_5485,N_2680,N_1898);
xor U5486 (N_5486,N_2009,N_3489);
nor U5487 (N_5487,N_2766,N_4977);
nor U5488 (N_5488,N_1599,N_3787);
nand U5489 (N_5489,N_2260,N_4619);
and U5490 (N_5490,N_2089,N_3527);
nor U5491 (N_5491,N_3038,N_2161);
or U5492 (N_5492,N_1342,N_3933);
or U5493 (N_5493,N_584,N_2560);
and U5494 (N_5494,N_1045,N_2103);
and U5495 (N_5495,N_2880,N_4324);
xnor U5496 (N_5496,N_451,N_4492);
and U5497 (N_5497,N_1127,N_3204);
nor U5498 (N_5498,N_3015,N_1794);
xor U5499 (N_5499,N_3641,N_4183);
nor U5500 (N_5500,N_4867,N_1529);
nand U5501 (N_5501,N_4224,N_3989);
or U5502 (N_5502,N_3824,N_3366);
nand U5503 (N_5503,N_2823,N_3731);
xnor U5504 (N_5504,N_60,N_1230);
nand U5505 (N_5505,N_1375,N_2672);
nand U5506 (N_5506,N_1748,N_125);
xor U5507 (N_5507,N_4772,N_2776);
xor U5508 (N_5508,N_2855,N_412);
nand U5509 (N_5509,N_3120,N_1726);
nor U5510 (N_5510,N_2897,N_3135);
xor U5511 (N_5511,N_3754,N_4834);
or U5512 (N_5512,N_3341,N_4840);
xor U5513 (N_5513,N_2863,N_33);
or U5514 (N_5514,N_3387,N_4038);
and U5515 (N_5515,N_547,N_910);
or U5516 (N_5516,N_339,N_4106);
nor U5517 (N_5517,N_2913,N_4862);
nor U5518 (N_5518,N_1070,N_1642);
xor U5519 (N_5519,N_712,N_4277);
and U5520 (N_5520,N_4881,N_4874);
or U5521 (N_5521,N_101,N_2717);
xor U5522 (N_5522,N_2026,N_1665);
nand U5523 (N_5523,N_869,N_4365);
or U5524 (N_5524,N_1651,N_183);
nand U5525 (N_5525,N_1821,N_3145);
nand U5526 (N_5526,N_1564,N_1392);
and U5527 (N_5527,N_579,N_3616);
nand U5528 (N_5528,N_306,N_4386);
nor U5529 (N_5529,N_4870,N_1547);
xor U5530 (N_5530,N_798,N_410);
or U5531 (N_5531,N_4508,N_4361);
and U5532 (N_5532,N_4669,N_2036);
nor U5533 (N_5533,N_3574,N_1183);
nand U5534 (N_5534,N_2542,N_2926);
and U5535 (N_5535,N_3441,N_1616);
or U5536 (N_5536,N_1428,N_1994);
nand U5537 (N_5537,N_1540,N_3034);
or U5538 (N_5538,N_330,N_4665);
nand U5539 (N_5539,N_2133,N_64);
or U5540 (N_5540,N_91,N_2916);
nand U5541 (N_5541,N_3994,N_2113);
nor U5542 (N_5542,N_696,N_2572);
nor U5543 (N_5543,N_4020,N_4027);
nor U5544 (N_5544,N_984,N_3095);
or U5545 (N_5545,N_1435,N_4973);
nand U5546 (N_5546,N_1960,N_2740);
and U5547 (N_5547,N_3675,N_1453);
nand U5548 (N_5548,N_4407,N_559);
or U5549 (N_5549,N_1887,N_1052);
nand U5550 (N_5550,N_3355,N_2923);
and U5551 (N_5551,N_4284,N_2746);
nand U5552 (N_5552,N_819,N_4377);
or U5553 (N_5553,N_3263,N_2244);
nand U5554 (N_5554,N_188,N_3879);
nor U5555 (N_5555,N_3800,N_1674);
nor U5556 (N_5556,N_4387,N_1199);
xor U5557 (N_5557,N_3453,N_3264);
xnor U5558 (N_5558,N_4045,N_3586);
and U5559 (N_5559,N_3117,N_1409);
xor U5560 (N_5560,N_1787,N_797);
nand U5561 (N_5561,N_3998,N_1888);
nor U5562 (N_5562,N_1940,N_1125);
or U5563 (N_5563,N_3735,N_3920);
or U5564 (N_5564,N_2869,N_778);
xor U5565 (N_5565,N_1802,N_4771);
and U5566 (N_5566,N_3080,N_3724);
nand U5567 (N_5567,N_1333,N_3833);
nand U5568 (N_5568,N_4890,N_1034);
xnor U5569 (N_5569,N_4723,N_261);
xnor U5570 (N_5570,N_4101,N_1545);
nor U5571 (N_5571,N_4996,N_2223);
and U5572 (N_5572,N_4674,N_4764);
and U5573 (N_5573,N_1170,N_1316);
nor U5574 (N_5574,N_2424,N_1007);
and U5575 (N_5575,N_1195,N_1581);
nor U5576 (N_5576,N_430,N_4593);
nor U5577 (N_5577,N_4932,N_1164);
nor U5578 (N_5578,N_2834,N_1804);
or U5579 (N_5579,N_4904,N_1610);
and U5580 (N_5580,N_3070,N_1102);
or U5581 (N_5581,N_1087,N_154);
and U5582 (N_5582,N_2813,N_4708);
nand U5583 (N_5583,N_3938,N_3700);
xor U5584 (N_5584,N_766,N_17);
and U5585 (N_5585,N_3485,N_969);
or U5586 (N_5586,N_2631,N_3068);
xor U5587 (N_5587,N_1963,N_2341);
nand U5588 (N_5588,N_1857,N_1467);
or U5589 (N_5589,N_4390,N_743);
and U5590 (N_5590,N_1526,N_4297);
nand U5591 (N_5591,N_3977,N_4408);
nor U5592 (N_5592,N_3537,N_1551);
xnor U5593 (N_5593,N_520,N_1774);
and U5594 (N_5594,N_530,N_4940);
nand U5595 (N_5595,N_3885,N_3474);
and U5596 (N_5596,N_2571,N_375);
or U5597 (N_5597,N_1779,N_4770);
or U5598 (N_5598,N_4194,N_359);
and U5599 (N_5599,N_4814,N_810);
and U5600 (N_5600,N_3315,N_4173);
xor U5601 (N_5601,N_1798,N_34);
or U5602 (N_5602,N_2445,N_3314);
and U5603 (N_5603,N_3664,N_2231);
nor U5604 (N_5604,N_3636,N_621);
or U5605 (N_5605,N_4873,N_4569);
xnor U5606 (N_5606,N_3012,N_3173);
or U5607 (N_5607,N_592,N_449);
and U5608 (N_5608,N_3072,N_1978);
or U5609 (N_5609,N_1360,N_1901);
or U5610 (N_5610,N_420,N_2355);
and U5611 (N_5611,N_2153,N_1462);
nand U5612 (N_5612,N_4913,N_1538);
xor U5613 (N_5613,N_698,N_2806);
nand U5614 (N_5614,N_472,N_1752);
or U5615 (N_5615,N_1985,N_1303);
and U5616 (N_5616,N_585,N_634);
xnor U5617 (N_5617,N_1758,N_3727);
nor U5618 (N_5618,N_4041,N_1841);
and U5619 (N_5619,N_1291,N_48);
xor U5620 (N_5620,N_2416,N_132);
or U5621 (N_5621,N_1010,N_1918);
or U5622 (N_5622,N_2005,N_799);
xnor U5623 (N_5623,N_2812,N_2649);
nand U5624 (N_5624,N_3781,N_962);
nor U5625 (N_5625,N_2318,N_3112);
xnor U5626 (N_5626,N_171,N_26);
or U5627 (N_5627,N_3227,N_4524);
nand U5628 (N_5628,N_1444,N_4464);
and U5629 (N_5629,N_2143,N_1589);
nor U5630 (N_5630,N_3866,N_4703);
nand U5631 (N_5631,N_4737,N_609);
nand U5632 (N_5632,N_2787,N_2116);
nor U5633 (N_5633,N_3940,N_839);
xnor U5634 (N_5634,N_3444,N_1699);
or U5635 (N_5635,N_2041,N_1175);
nand U5636 (N_5636,N_1878,N_4057);
nand U5637 (N_5637,N_4780,N_574);
and U5638 (N_5638,N_2390,N_2695);
nand U5639 (N_5639,N_1814,N_728);
and U5640 (N_5640,N_599,N_3285);
nor U5641 (N_5641,N_73,N_1337);
and U5642 (N_5642,N_4463,N_4901);
nand U5643 (N_5643,N_4797,N_3583);
nor U5644 (N_5644,N_1663,N_1586);
or U5645 (N_5645,N_3491,N_4046);
nor U5646 (N_5646,N_4301,N_2334);
or U5647 (N_5647,N_4678,N_1983);
and U5648 (N_5648,N_4606,N_1846);
and U5649 (N_5649,N_1079,N_2118);
xor U5650 (N_5650,N_414,N_4914);
and U5651 (N_5651,N_4717,N_2349);
xnor U5652 (N_5652,N_181,N_254);
xnor U5653 (N_5653,N_3078,N_553);
nor U5654 (N_5654,N_4504,N_4521);
xor U5655 (N_5655,N_2526,N_4450);
nor U5656 (N_5656,N_391,N_2228);
or U5657 (N_5657,N_3035,N_2045);
nand U5658 (N_5658,N_4154,N_3202);
and U5659 (N_5659,N_363,N_1267);
or U5660 (N_5660,N_3530,N_2608);
nand U5661 (N_5661,N_3364,N_3427);
nand U5662 (N_5662,N_1971,N_3764);
nor U5663 (N_5663,N_1114,N_896);
and U5664 (N_5664,N_3162,N_848);
nand U5665 (N_5665,N_2242,N_4467);
nand U5666 (N_5666,N_3465,N_961);
nand U5667 (N_5667,N_711,N_2493);
or U5668 (N_5668,N_1434,N_3308);
and U5669 (N_5669,N_2245,N_4720);
xnor U5670 (N_5670,N_3697,N_2487);
xor U5671 (N_5671,N_1270,N_1660);
nor U5672 (N_5672,N_3658,N_3806);
xnor U5673 (N_5673,N_1193,N_941);
xnor U5674 (N_5674,N_4343,N_428);
and U5675 (N_5675,N_99,N_1253);
or U5676 (N_5676,N_4591,N_4736);
nand U5677 (N_5677,N_4787,N_4871);
or U5678 (N_5678,N_4093,N_859);
or U5679 (N_5679,N_3471,N_159);
nand U5680 (N_5680,N_1286,N_3470);
xnor U5681 (N_5681,N_1459,N_4342);
or U5682 (N_5682,N_1868,N_834);
nand U5683 (N_5683,N_368,N_4535);
nand U5684 (N_5684,N_4470,N_4707);
or U5685 (N_5685,N_604,N_4952);
nor U5686 (N_5686,N_1579,N_92);
nand U5687 (N_5687,N_4796,N_2308);
and U5688 (N_5688,N_394,N_3100);
xor U5689 (N_5689,N_4912,N_668);
xnor U5690 (N_5690,N_2039,N_3242);
nand U5691 (N_5691,N_3368,N_4961);
xnor U5692 (N_5692,N_388,N_870);
and U5693 (N_5693,N_4014,N_1430);
or U5694 (N_5694,N_1449,N_55);
nand U5695 (N_5695,N_51,N_3777);
and U5696 (N_5696,N_2084,N_447);
or U5697 (N_5697,N_4257,N_2168);
xor U5698 (N_5698,N_2431,N_3401);
and U5699 (N_5699,N_2071,N_560);
and U5700 (N_5700,N_2121,N_3391);
or U5701 (N_5701,N_1251,N_4969);
nand U5702 (N_5702,N_310,N_863);
and U5703 (N_5703,N_4646,N_2959);
or U5704 (N_5704,N_1030,N_950);
nand U5705 (N_5705,N_1972,N_2889);
xor U5706 (N_5706,N_1352,N_633);
and U5707 (N_5707,N_4135,N_401);
xnor U5708 (N_5708,N_3158,N_4341);
and U5709 (N_5709,N_1631,N_1750);
or U5710 (N_5710,N_3312,N_369);
or U5711 (N_5711,N_134,N_4477);
and U5712 (N_5712,N_244,N_716);
nand U5713 (N_5713,N_4594,N_1480);
and U5714 (N_5714,N_4389,N_3882);
xor U5715 (N_5715,N_670,N_1562);
nand U5716 (N_5716,N_4507,N_1546);
and U5717 (N_5717,N_4566,N_1130);
nand U5718 (N_5718,N_2839,N_554);
nand U5719 (N_5719,N_847,N_4329);
and U5720 (N_5720,N_2965,N_605);
nand U5721 (N_5721,N_1497,N_209);
xnor U5722 (N_5722,N_2206,N_3298);
xnor U5723 (N_5723,N_4278,N_2225);
or U5724 (N_5724,N_3984,N_3149);
nor U5725 (N_5725,N_4235,N_286);
or U5726 (N_5726,N_4146,N_3157);
xor U5727 (N_5727,N_2411,N_2888);
or U5728 (N_5728,N_1525,N_1058);
and U5729 (N_5729,N_441,N_3139);
and U5730 (N_5730,N_2790,N_946);
or U5731 (N_5731,N_4908,N_2326);
or U5732 (N_5732,N_3625,N_3808);
xor U5733 (N_5733,N_3081,N_1076);
and U5734 (N_5734,N_2360,N_4123);
nand U5735 (N_5735,N_840,N_3008);
nand U5736 (N_5736,N_582,N_1172);
or U5737 (N_5737,N_4424,N_1582);
xnor U5738 (N_5738,N_954,N_1747);
nor U5739 (N_5739,N_262,N_2696);
nor U5740 (N_5740,N_3447,N_2908);
nor U5741 (N_5741,N_4044,N_3086);
xor U5742 (N_5742,N_4758,N_4640);
xor U5743 (N_5743,N_1881,N_1094);
nor U5744 (N_5744,N_3373,N_4547);
nand U5745 (N_5745,N_4098,N_3619);
and U5746 (N_5746,N_157,N_3190);
nor U5747 (N_5747,N_3907,N_3067);
and U5748 (N_5748,N_1397,N_4542);
and U5749 (N_5749,N_1542,N_3681);
nor U5750 (N_5750,N_3674,N_45);
xor U5751 (N_5751,N_548,N_4118);
nor U5752 (N_5752,N_370,N_141);
or U5753 (N_5753,N_1738,N_3495);
nand U5754 (N_5754,N_485,N_131);
and U5755 (N_5755,N_2538,N_909);
or U5756 (N_5756,N_1947,N_4777);
and U5757 (N_5757,N_2434,N_1167);
nor U5758 (N_5758,N_2828,N_1277);
or U5759 (N_5759,N_2636,N_479);
nand U5760 (N_5760,N_2927,N_3431);
and U5761 (N_5761,N_2597,N_4271);
and U5762 (N_5762,N_174,N_1031);
nand U5763 (N_5763,N_3786,N_4791);
xor U5764 (N_5764,N_3517,N_630);
nand U5765 (N_5765,N_1724,N_1823);
nand U5766 (N_5766,N_717,N_2380);
nand U5767 (N_5767,N_1639,N_122);
or U5768 (N_5768,N_2376,N_1194);
xnor U5769 (N_5769,N_75,N_593);
or U5770 (N_5770,N_1326,N_4335);
and U5771 (N_5771,N_1973,N_1935);
nor U5772 (N_5772,N_862,N_1783);
and U5773 (N_5773,N_1605,N_320);
nor U5774 (N_5774,N_3568,N_2945);
and U5775 (N_5775,N_4455,N_4944);
xnor U5776 (N_5776,N_1437,N_2309);
and U5777 (N_5777,N_4394,N_1379);
xor U5778 (N_5778,N_2205,N_3987);
nand U5779 (N_5779,N_2612,N_2996);
xor U5780 (N_5780,N_4258,N_4190);
or U5781 (N_5781,N_334,N_4400);
xnor U5782 (N_5782,N_1082,N_657);
nor U5783 (N_5783,N_4481,N_76);
and U5784 (N_5784,N_3090,N_924);
xnor U5785 (N_5785,N_1707,N_377);
and U5786 (N_5786,N_456,N_3230);
xor U5787 (N_5787,N_3423,N_3601);
nand U5788 (N_5788,N_1717,N_2540);
and U5789 (N_5789,N_4709,N_4186);
nor U5790 (N_5790,N_959,N_1970);
and U5791 (N_5791,N_4439,N_958);
xor U5792 (N_5792,N_985,N_3172);
nor U5793 (N_5793,N_1689,N_105);
and U5794 (N_5794,N_4452,N_264);
nor U5795 (N_5795,N_4992,N_3213);
nor U5796 (N_5796,N_648,N_2177);
or U5797 (N_5797,N_3759,N_1177);
or U5798 (N_5798,N_4864,N_2419);
nand U5799 (N_5799,N_3750,N_2204);
nor U5800 (N_5800,N_2216,N_1280);
xnor U5801 (N_5801,N_516,N_50);
nor U5802 (N_5802,N_2078,N_3422);
or U5803 (N_5803,N_581,N_1838);
and U5804 (N_5804,N_2359,N_4987);
xor U5805 (N_5805,N_197,N_1706);
nand U5806 (N_5806,N_1004,N_3504);
or U5807 (N_5807,N_3200,N_177);
nand U5808 (N_5808,N_4275,N_3167);
or U5809 (N_5809,N_4005,N_1661);
nor U5810 (N_5810,N_3417,N_1926);
and U5811 (N_5811,N_4930,N_602);
or U5812 (N_5812,N_4743,N_1754);
and U5813 (N_5813,N_3861,N_3317);
nand U5814 (N_5814,N_616,N_3703);
and U5815 (N_5815,N_1192,N_2034);
and U5816 (N_5816,N_3858,N_2522);
nand U5817 (N_5817,N_1097,N_3637);
or U5818 (N_5818,N_3629,N_3147);
xor U5819 (N_5819,N_889,N_4953);
nor U5820 (N_5820,N_735,N_685);
xor U5821 (N_5821,N_737,N_3836);
or U5822 (N_5822,N_2298,N_615);
xnor U5823 (N_5823,N_180,N_3928);
xnor U5824 (N_5824,N_4577,N_72);
nand U5825 (N_5825,N_1490,N_623);
xnor U5826 (N_5826,N_2925,N_2459);
or U5827 (N_5827,N_169,N_1936);
xnor U5828 (N_5828,N_164,N_2779);
nand U5829 (N_5829,N_3991,N_235);
and U5830 (N_5830,N_2887,N_2853);
or U5831 (N_5831,N_3905,N_1810);
xor U5832 (N_5832,N_2444,N_4801);
and U5833 (N_5833,N_4858,N_2713);
and U5834 (N_5834,N_2974,N_498);
or U5835 (N_5835,N_3841,N_4739);
nand U5836 (N_5836,N_3913,N_757);
nand U5837 (N_5837,N_4898,N_4896);
nor U5838 (N_5838,N_1698,N_2040);
nor U5839 (N_5839,N_1618,N_4495);
nor U5840 (N_5840,N_1650,N_415);
and U5841 (N_5841,N_3702,N_4362);
or U5842 (N_5842,N_1224,N_4126);
and U5843 (N_5843,N_220,N_2684);
and U5844 (N_5844,N_755,N_1953);
nand U5845 (N_5845,N_2432,N_4767);
and U5846 (N_5846,N_1296,N_892);
and U5847 (N_5847,N_4009,N_4152);
and U5848 (N_5848,N_3603,N_2301);
and U5849 (N_5849,N_2112,N_2233);
and U5850 (N_5850,N_645,N_3021);
xnor U5851 (N_5851,N_4550,N_982);
nor U5852 (N_5852,N_925,N_629);
nor U5853 (N_5853,N_266,N_1408);
xor U5854 (N_5854,N_2782,N_3893);
or U5855 (N_5855,N_4951,N_875);
or U5856 (N_5856,N_335,N_1786);
nor U5857 (N_5857,N_2687,N_3351);
xnor U5858 (N_5858,N_773,N_4141);
nand U5859 (N_5859,N_3288,N_3118);
nand U5860 (N_5860,N_4667,N_1567);
nand U5861 (N_5861,N_2999,N_4808);
or U5862 (N_5862,N_1696,N_1929);
xor U5863 (N_5863,N_1324,N_2635);
or U5864 (N_5864,N_2519,N_2931);
nand U5865 (N_5865,N_1521,N_2681);
nor U5866 (N_5866,N_1578,N_349);
nand U5867 (N_5867,N_3439,N_2258);
nor U5868 (N_5868,N_2733,N_210);
or U5869 (N_5869,N_678,N_874);
or U5870 (N_5870,N_3345,N_2977);
nor U5871 (N_5871,N_1622,N_213);
xnor U5872 (N_5872,N_4445,N_1332);
and U5873 (N_5873,N_3738,N_1762);
nor U5874 (N_5874,N_4199,N_236);
and U5875 (N_5875,N_3477,N_3252);
xor U5876 (N_5876,N_2670,N_2751);
xnor U5877 (N_5877,N_84,N_573);
nor U5878 (N_5878,N_2268,N_1369);
nor U5879 (N_5879,N_3714,N_139);
nor U5880 (N_5880,N_2978,N_4034);
and U5881 (N_5881,N_2060,N_1363);
nand U5882 (N_5882,N_2529,N_3589);
or U5883 (N_5883,N_1243,N_1609);
and U5884 (N_5884,N_594,N_1008);
nand U5885 (N_5885,N_1398,N_3632);
nor U5886 (N_5886,N_4066,N_713);
nor U5887 (N_5887,N_3776,N_3331);
nor U5888 (N_5888,N_3588,N_1119);
and U5889 (N_5889,N_4204,N_3798);
and U5890 (N_5890,N_1759,N_4244);
nand U5891 (N_5891,N_2633,N_1207);
nand U5892 (N_5892,N_4990,N_852);
and U5893 (N_5893,N_2743,N_756);
nor U5894 (N_5894,N_1066,N_3362);
nand U5895 (N_5895,N_942,N_3511);
xor U5896 (N_5896,N_3835,N_1828);
and U5897 (N_5897,N_145,N_2934);
xnor U5898 (N_5898,N_2172,N_2640);
and U5899 (N_5899,N_1690,N_1946);
xor U5900 (N_5900,N_549,N_873);
nand U5901 (N_5901,N_2090,N_4496);
nand U5902 (N_5902,N_586,N_3591);
nand U5903 (N_5903,N_2577,N_4104);
nor U5904 (N_5904,N_976,N_642);
nand U5905 (N_5905,N_1515,N_3916);
xor U5906 (N_5906,N_3198,N_1694);
xnor U5907 (N_5907,N_885,N_3807);
nor U5908 (N_5908,N_3502,N_3971);
nand U5909 (N_5909,N_2492,N_3523);
and U5910 (N_5910,N_4710,N_1311);
nand U5911 (N_5911,N_3020,N_2994);
nand U5912 (N_5912,N_337,N_2667);
nor U5913 (N_5913,N_2141,N_274);
xor U5914 (N_5914,N_1367,N_980);
or U5915 (N_5915,N_3609,N_686);
nor U5916 (N_5916,N_1753,N_1018);
nand U5917 (N_5917,N_3608,N_1575);
or U5918 (N_5918,N_1832,N_806);
nor U5919 (N_5919,N_3695,N_3878);
or U5920 (N_5920,N_4356,N_1149);
nor U5921 (N_5921,N_110,N_4604);
nand U5922 (N_5922,N_4779,N_3630);
and U5923 (N_5923,N_501,N_703);
and U5924 (N_5924,N_3281,N_1933);
xor U5925 (N_5925,N_2930,N_233);
or U5926 (N_5926,N_4700,N_265);
or U5927 (N_5927,N_1228,N_3237);
and U5928 (N_5928,N_2606,N_4553);
and U5929 (N_5929,N_3292,N_3721);
nor U5930 (N_5930,N_4859,N_4280);
nand U5931 (N_5931,N_1349,N_3782);
and U5932 (N_5932,N_3411,N_947);
and U5933 (N_5933,N_1044,N_641);
xnor U5934 (N_5934,N_2430,N_569);
nor U5935 (N_5935,N_3925,N_1285);
xor U5936 (N_5936,N_564,N_2969);
or U5937 (N_5937,N_133,N_989);
and U5938 (N_5938,N_4370,N_2012);
nand U5939 (N_5939,N_3060,N_4249);
or U5940 (N_5940,N_1781,N_2105);
or U5941 (N_5941,N_1069,N_1692);
or U5942 (N_5942,N_109,N_972);
or U5943 (N_5943,N_2481,N_4089);
xnor U5944 (N_5944,N_3966,N_13);
nand U5945 (N_5945,N_1643,N_3723);
xor U5946 (N_5946,N_3605,N_1181);
nor U5947 (N_5947,N_3648,N_3767);
and U5948 (N_5948,N_2023,N_161);
nand U5949 (N_5949,N_4948,N_2451);
nand U5950 (N_5950,N_116,N_0);
and U5951 (N_5951,N_662,N_1111);
nor U5952 (N_5952,N_1769,N_1872);
or U5953 (N_5953,N_4878,N_2125);
or U5954 (N_5954,N_3191,N_207);
and U5955 (N_5955,N_1939,N_3438);
nor U5956 (N_5956,N_4256,N_1089);
nand U5957 (N_5957,N_2588,N_811);
or U5958 (N_5958,N_3874,N_2668);
xnor U5959 (N_5959,N_4067,N_324);
nand U5960 (N_5960,N_3549,N_1812);
nor U5961 (N_5961,N_2951,N_1035);
or U5962 (N_5962,N_1509,N_351);
and U5963 (N_5963,N_2738,N_3956);
xor U5964 (N_5964,N_1491,N_4079);
nand U5965 (N_5965,N_2057,N_899);
nor U5966 (N_5966,N_382,N_4680);
and U5967 (N_5967,N_2868,N_913);
nand U5968 (N_5968,N_3766,N_2895);
xnor U5969 (N_5969,N_568,N_3543);
and U5970 (N_5970,N_3730,N_3704);
nand U5971 (N_5971,N_14,N_2497);
nor U5972 (N_5972,N_4240,N_16);
and U5973 (N_5973,N_1943,N_1990);
nand U5974 (N_5974,N_1319,N_2285);
nand U5975 (N_5975,N_2137,N_3418);
xnor U5976 (N_5976,N_821,N_255);
nor U5977 (N_5977,N_9,N_2138);
nand U5978 (N_5978,N_4580,N_151);
xor U5979 (N_5979,N_3041,N_3467);
or U5980 (N_5980,N_4191,N_2599);
nand U5981 (N_5981,N_289,N_3214);
or U5982 (N_5982,N_268,N_3707);
or U5983 (N_5983,N_2155,N_3840);
and U5984 (N_5984,N_4438,N_781);
nor U5985 (N_5985,N_2425,N_1047);
or U5986 (N_5986,N_2650,N_80);
nor U5987 (N_5987,N_3912,N_4883);
xor U5988 (N_5988,N_1890,N_3194);
nand U5989 (N_5989,N_1729,N_1968);
nand U5990 (N_5990,N_905,N_4412);
or U5991 (N_5991,N_2756,N_3424);
nor U5992 (N_5992,N_2730,N_953);
or U5993 (N_5993,N_2449,N_4033);
nand U5994 (N_5994,N_3995,N_3655);
or U5995 (N_5995,N_4927,N_4837);
and U5996 (N_5996,N_2979,N_628);
nor U5997 (N_5997,N_4962,N_138);
and U5998 (N_5998,N_2791,N_374);
or U5999 (N_5999,N_2110,N_4831);
nand U6000 (N_6000,N_3339,N_1988);
xnor U6001 (N_6001,N_124,N_4314);
and U6002 (N_6002,N_4170,N_3757);
nor U6003 (N_6003,N_832,N_4442);
or U6004 (N_6004,N_808,N_1701);
nand U6005 (N_6005,N_1019,N_1760);
xnor U6006 (N_6006,N_988,N_1468);
or U6007 (N_6007,N_545,N_1705);
nor U6008 (N_6008,N_1377,N_1749);
nand U6009 (N_6009,N_3049,N_2455);
nor U6010 (N_6010,N_3025,N_3302);
nor U6011 (N_6011,N_3212,N_4015);
or U6012 (N_6012,N_1028,N_1656);
xor U6013 (N_6013,N_3710,N_890);
and U6014 (N_6014,N_2734,N_1166);
or U6015 (N_6015,N_418,N_4358);
xor U6016 (N_6016,N_4159,N_1827);
nor U6017 (N_6017,N_4749,N_4262);
xnor U6018 (N_6018,N_2250,N_1684);
or U6019 (N_6019,N_3108,N_4805);
xnor U6020 (N_6020,N_1215,N_509);
nor U6021 (N_6021,N_2098,N_4933);
xnor U6022 (N_6022,N_935,N_3436);
xor U6023 (N_6023,N_2793,N_205);
xor U6024 (N_6024,N_3260,N_3659);
nand U6025 (N_6025,N_3084,N_3544);
and U6026 (N_6026,N_242,N_1641);
nor U6027 (N_6027,N_496,N_587);
and U6028 (N_6028,N_911,N_1630);
nor U6029 (N_6029,N_3736,N_677);
nand U6030 (N_6030,N_4317,N_1396);
or U6031 (N_6031,N_4512,N_4599);
nor U6032 (N_6032,N_4555,N_426);
and U6033 (N_6033,N_588,N_1534);
nand U6034 (N_6034,N_3291,N_2319);
and U6035 (N_6035,N_3033,N_1837);
xnor U6036 (N_6036,N_3856,N_4294);
and U6037 (N_6037,N_1465,N_3643);
nand U6038 (N_6038,N_3318,N_934);
or U6039 (N_6039,N_4071,N_625);
nand U6040 (N_6040,N_1386,N_4384);
nand U6041 (N_6041,N_165,N_1552);
nand U6042 (N_6042,N_2356,N_824);
nand U6043 (N_6043,N_2611,N_1849);
nor U6044 (N_6044,N_3778,N_4273);
xnor U6045 (N_6045,N_4822,N_2461);
or U6046 (N_6046,N_1919,N_2949);
nand U6047 (N_6047,N_4212,N_1471);
and U6048 (N_6048,N_4658,N_4214);
xnor U6049 (N_6049,N_468,N_3016);
or U6050 (N_6050,N_2767,N_1634);
nand U6051 (N_6051,N_782,N_2470);
nor U6052 (N_6052,N_531,N_3888);
nor U6053 (N_6053,N_103,N_1664);
xor U6054 (N_6054,N_4785,N_4465);
or U6055 (N_6055,N_2270,N_2263);
and U6056 (N_6056,N_2583,N_2435);
and U6057 (N_6057,N_785,N_3065);
nand U6058 (N_6058,N_2876,N_1388);
or U6059 (N_6059,N_3843,N_3791);
xnor U6060 (N_6060,N_1964,N_4029);
and U6061 (N_6061,N_4223,N_1505);
or U6062 (N_6062,N_2692,N_1043);
nand U6063 (N_6063,N_831,N_3142);
nor U6064 (N_6064,N_4910,N_1085);
nor U6065 (N_6065,N_4747,N_2375);
nand U6066 (N_6066,N_646,N_4028);
nand U6067 (N_6067,N_4287,N_194);
and U6068 (N_6068,N_457,N_3492);
nand U6069 (N_6069,N_517,N_1543);
nand U6070 (N_6070,N_4564,N_3098);
nand U6071 (N_6071,N_364,N_3852);
and U6072 (N_6072,N_2043,N_2374);
xnor U6073 (N_6073,N_3463,N_4443);
nor U6074 (N_6074,N_3024,N_800);
xor U6075 (N_6075,N_1766,N_4769);
or U6076 (N_6076,N_667,N_3336);
or U6077 (N_6077,N_4956,N_3644);
nand U6078 (N_6078,N_4095,N_4598);
and U6079 (N_6079,N_1115,N_4689);
or U6080 (N_6080,N_3813,N_4527);
nor U6081 (N_6081,N_2773,N_3014);
xnor U6082 (N_6082,N_1263,N_3429);
or U6083 (N_6083,N_4217,N_1654);
and U6084 (N_6084,N_2579,N_2810);
nand U6085 (N_6085,N_4653,N_1612);
and U6086 (N_6086,N_355,N_3746);
nor U6087 (N_6087,N_4572,N_1458);
nor U6088 (N_6088,N_1341,N_1632);
nand U6089 (N_6089,N_1269,N_3665);
xnor U6090 (N_6090,N_4963,N_4385);
xor U6091 (N_6091,N_256,N_386);
or U6092 (N_6092,N_3327,N_2297);
or U6093 (N_6093,N_4839,N_3156);
nor U6094 (N_6094,N_1861,N_298);
nand U6095 (N_6095,N_2708,N_2371);
nand U6096 (N_6096,N_4936,N_2191);
or U6097 (N_6097,N_990,N_2725);
nand U6098 (N_6098,N_3557,N_4084);
xnor U6099 (N_6099,N_1382,N_1108);
and U6100 (N_6100,N_3876,N_2589);
nand U6101 (N_6101,N_2832,N_2524);
xor U6102 (N_6102,N_1050,N_864);
nand U6103 (N_6103,N_2976,N_2573);
xor U6104 (N_6104,N_3210,N_2703);
or U6105 (N_6105,N_2757,N_208);
nand U6106 (N_6106,N_4894,N_3125);
or U6107 (N_6107,N_2568,N_2627);
nor U6108 (N_6108,N_714,N_1685);
or U6109 (N_6109,N_3961,N_2825);
xor U6110 (N_6110,N_200,N_2679);
or U6111 (N_6111,N_4461,N_916);
and U6112 (N_6112,N_3853,N_2104);
nor U6113 (N_6113,N_3615,N_4768);
nand U6114 (N_6114,N_4843,N_2582);
xor U6115 (N_6115,N_843,N_2140);
nand U6116 (N_6116,N_2176,N_1001);
or U6117 (N_6117,N_3040,N_3831);
xor U6118 (N_6118,N_199,N_1800);
or U6119 (N_6119,N_2550,N_3245);
or U6120 (N_6120,N_1440,N_2412);
and U6121 (N_6121,N_575,N_2803);
or U6122 (N_6122,N_4844,N_2316);
and U6123 (N_6123,N_3052,N_3635);
and U6124 (N_6124,N_1574,N_3673);
or U6125 (N_6125,N_1624,N_3768);
xnor U6126 (N_6126,N_204,N_1288);
and U6127 (N_6127,N_250,N_697);
xnor U6128 (N_6128,N_503,N_4157);
or U6129 (N_6129,N_3056,N_3240);
nand U6130 (N_6130,N_3538,N_4763);
xor U6131 (N_6131,N_1636,N_385);
and U6132 (N_6132,N_1403,N_1915);
nor U6133 (N_6133,N_2558,N_3460);
xor U6134 (N_6134,N_4698,N_2904);
and U6135 (N_6135,N_4687,N_3437);
nand U6136 (N_6136,N_2601,N_4888);
nand U6137 (N_6137,N_2625,N_3275);
or U6138 (N_6138,N_442,N_4374);
or U6139 (N_6139,N_4931,N_898);
xnor U6140 (N_6140,N_1134,N_3802);
xor U6141 (N_6141,N_2465,N_1997);
xnor U6142 (N_6142,N_904,N_1775);
nand U6143 (N_6143,N_1038,N_1173);
xnor U6144 (N_6144,N_2623,N_4884);
nor U6145 (N_6145,N_1899,N_427);
nand U6146 (N_6146,N_533,N_1314);
nor U6147 (N_6147,N_1389,N_2007);
xor U6148 (N_6148,N_3146,N_3716);
nand U6149 (N_6149,N_4198,N_3894);
and U6150 (N_6150,N_3010,N_425);
xor U6151 (N_6151,N_3973,N_23);
and U6152 (N_6152,N_2059,N_1220);
nor U6153 (N_6153,N_3039,N_2388);
nand U6154 (N_6154,N_4812,N_4116);
or U6155 (N_6155,N_1432,N_3939);
nand U6156 (N_6156,N_3743,N_1691);
xor U6157 (N_6157,N_3972,N_2146);
and U6158 (N_6158,N_758,N_49);
and U6159 (N_6159,N_4644,N_1511);
nand U6160 (N_6160,N_4326,N_4752);
xnor U6161 (N_6161,N_4696,N_3408);
nand U6162 (N_6162,N_3143,N_2377);
and U6163 (N_6163,N_3942,N_4947);
nand U6164 (N_6164,N_3685,N_4137);
and U6165 (N_6165,N_1916,N_4795);
and U6166 (N_6166,N_2174,N_1002);
or U6167 (N_6167,N_2414,N_1646);
or U6168 (N_6168,N_4635,N_4032);
and U6169 (N_6169,N_4643,N_4147);
nor U6170 (N_6170,N_2919,N_2613);
xor U6171 (N_6171,N_1667,N_2420);
and U6172 (N_6172,N_643,N_1464);
and U6173 (N_6173,N_2721,N_1422);
and U6174 (N_6174,N_512,N_3234);
xnor U6175 (N_6175,N_637,N_2018);
xnor U6176 (N_6176,N_2516,N_565);
nor U6177 (N_6177,N_854,N_649);
or U6178 (N_6178,N_2384,N_3061);
nor U6179 (N_6179,N_3838,N_815);
nor U6180 (N_6180,N_1559,N_2391);
and U6181 (N_6181,N_2117,N_939);
nor U6182 (N_6182,N_2528,N_4835);
xor U6183 (N_6183,N_3801,N_1585);
or U6184 (N_6184,N_2122,N_3985);
nor U6185 (N_6185,N_406,N_271);
xnor U6186 (N_6186,N_2123,N_11);
xnor U6187 (N_6187,N_1105,N_4727);
nor U6188 (N_6188,N_3440,N_3592);
xnor U6189 (N_6189,N_4270,N_4993);
xor U6190 (N_6190,N_502,N_541);
and U6191 (N_6191,N_4892,N_2736);
xnor U6192 (N_6192,N_1502,N_776);
or U6193 (N_6193,N_660,N_674);
nand U6194 (N_6194,N_2107,N_2139);
xor U6195 (N_6195,N_1850,N_2199);
xnor U6196 (N_6196,N_3007,N_1930);
or U6197 (N_6197,N_2514,N_4288);
nor U6198 (N_6198,N_4290,N_830);
nor U6199 (N_6199,N_3486,N_1796);
nor U6200 (N_6200,N_3548,N_1657);
nor U6201 (N_6201,N_2638,N_3934);
nor U6202 (N_6202,N_2367,N_3917);
and U6203 (N_6203,N_1256,N_3627);
xnor U6204 (N_6204,N_835,N_740);
nand U6205 (N_6205,N_360,N_4869);
nand U6206 (N_6206,N_2259,N_2292);
and U6207 (N_6207,N_4876,N_2798);
or U6208 (N_6208,N_751,N_3520);
nor U6209 (N_6209,N_1950,N_1757);
xnor U6210 (N_6210,N_4759,N_3472);
nand U6211 (N_6211,N_4722,N_3487);
or U6212 (N_6212,N_1073,N_513);
nor U6213 (N_6213,N_1427,N_489);
xnor U6214 (N_6214,N_483,N_709);
xnor U6215 (N_6215,N_4712,N_390);
or U6216 (N_6216,N_1987,N_1638);
xor U6217 (N_6217,N_307,N_1182);
or U6218 (N_6218,N_90,N_319);
or U6219 (N_6219,N_2115,N_3541);
nand U6220 (N_6220,N_1580,N_439);
nand U6221 (N_6221,N_59,N_1260);
nor U6222 (N_6222,N_1372,N_1544);
xnor U6223 (N_6223,N_1801,N_3215);
xnor U6224 (N_6224,N_1191,N_2328);
or U6225 (N_6225,N_1508,N_3036);
or U6226 (N_6226,N_2147,N_41);
nor U6227 (N_6227,N_1470,N_1494);
or U6228 (N_6228,N_3226,N_4788);
nand U6229 (N_6229,N_3169,N_1098);
xor U6230 (N_6230,N_438,N_4042);
or U6231 (N_6231,N_2311,N_4340);
nand U6232 (N_6232,N_1938,N_3769);
and U6233 (N_6233,N_2759,N_1223);
nand U6234 (N_6234,N_3296,N_1693);
and U6235 (N_6235,N_129,N_2504);
nor U6236 (N_6236,N_926,N_3403);
nand U6237 (N_6237,N_1148,N_95);
and U6238 (N_6238,N_3963,N_1011);
nand U6239 (N_6239,N_357,N_4233);
nor U6240 (N_6240,N_3186,N_1152);
xor U6241 (N_6241,N_4845,N_1107);
nor U6242 (N_6242,N_216,N_1283);
nand U6243 (N_6243,N_544,N_4715);
nand U6244 (N_6244,N_4241,N_4958);
and U6245 (N_6245,N_3909,N_2486);
and U6246 (N_6246,N_251,N_3516);
xor U6247 (N_6247,N_4733,N_2764);
nor U6248 (N_6248,N_4344,N_2067);
and U6249 (N_6249,N_2070,N_3820);
nand U6250 (N_6250,N_4510,N_3255);
xnor U6251 (N_6251,N_3638,N_1532);
and U6252 (N_6252,N_1456,N_2808);
and U6253 (N_6253,N_1905,N_2312);
or U6254 (N_6254,N_257,N_2353);
xor U6255 (N_6255,N_4552,N_1473);
xnor U6256 (N_6256,N_2739,N_790);
and U6257 (N_6257,N_1414,N_866);
xnor U6258 (N_6258,N_975,N_1227);
nand U6259 (N_6259,N_2017,N_4458);
and U6260 (N_6260,N_4832,N_3421);
xnor U6261 (N_6261,N_956,N_2421);
nand U6262 (N_6262,N_4517,N_4776);
and U6263 (N_6263,N_1235,N_4293);
nand U6264 (N_6264,N_820,N_578);
nor U6265 (N_6265,N_1479,N_1176);
and U6266 (N_6266,N_1535,N_1346);
nand U6267 (N_6267,N_2575,N_3748);
or U6268 (N_6268,N_2689,N_2718);
or U6269 (N_6269,N_3614,N_1084);
xnor U6270 (N_6270,N_1954,N_1830);
nand U6271 (N_6271,N_4565,N_3166);
and U6272 (N_6272,N_2501,N_4539);
xor U6273 (N_6273,N_3689,N_4236);
nor U6274 (N_6274,N_1883,N_407);
nor U6275 (N_6275,N_2496,N_2712);
or U6276 (N_6276,N_3501,N_1312);
nor U6277 (N_6277,N_2807,N_2552);
nor U6278 (N_6278,N_1710,N_3692);
nor U6279 (N_6279,N_2920,N_1370);
nor U6280 (N_6280,N_2438,N_2200);
xnor U6281 (N_6281,N_4144,N_4699);
xnor U6282 (N_6282,N_4694,N_3347);
or U6283 (N_6283,N_4662,N_1942);
xor U6284 (N_6284,N_4158,N_931);
and U6285 (N_6285,N_2300,N_3805);
and U6286 (N_6286,N_4821,N_1541);
nand U6287 (N_6287,N_1145,N_3326);
nor U6288 (N_6288,N_4023,N_1029);
xor U6289 (N_6289,N_222,N_1025);
nor U6290 (N_6290,N_3851,N_4318);
or U6291 (N_6291,N_1702,N_3261);
nor U6292 (N_6292,N_1649,N_1553);
nor U6293 (N_6293,N_1733,N_841);
or U6294 (N_6294,N_153,N_2289);
nand U6295 (N_6295,N_2788,N_3604);
or U6296 (N_6296,N_552,N_3617);
and U6297 (N_6297,N_1908,N_4000);
nand U6298 (N_6298,N_4145,N_4907);
xnor U6299 (N_6299,N_2013,N_2086);
nor U6300 (N_6300,N_3037,N_4360);
xnor U6301 (N_6301,N_3250,N_243);
xnor U6302 (N_6302,N_2187,N_4039);
nor U6303 (N_6303,N_2369,N_182);
xnor U6304 (N_6304,N_2626,N_880);
nor U6305 (N_6305,N_3307,N_675);
nor U6306 (N_6306,N_3902,N_4451);
or U6307 (N_6307,N_1600,N_1533);
xor U6308 (N_6308,N_1536,N_4100);
and U6309 (N_6309,N_627,N_3996);
xor U6310 (N_6310,N_4209,N_827);
nor U6311 (N_6311,N_3514,N_3397);
nor U6312 (N_6312,N_303,N_3598);
nand U6313 (N_6313,N_2710,N_861);
or U6314 (N_6314,N_1276,N_796);
and U6315 (N_6315,N_3679,N_4571);
nor U6316 (N_6316,N_1118,N_4061);
nand U6317 (N_6317,N_1617,N_237);
nand U6318 (N_6318,N_1300,N_1091);
xor U6319 (N_6319,N_1395,N_1241);
nand U6320 (N_6320,N_4131,N_4922);
xnor U6321 (N_6321,N_4605,N_2914);
or U6322 (N_6322,N_3561,N_4916);
xnor U6323 (N_6323,N_4127,N_2475);
and U6324 (N_6324,N_1867,N_4960);
or U6325 (N_6325,N_1481,N_4319);
nand U6326 (N_6326,N_1197,N_2954);
and U6327 (N_6327,N_2108,N_4798);
and U6328 (N_6328,N_4754,N_1959);
and U6329 (N_6329,N_1675,N_1519);
nand U6330 (N_6330,N_558,N_3948);
xor U6331 (N_6331,N_3982,N_4128);
nand U6332 (N_6332,N_3499,N_4824);
or U6333 (N_6333,N_2605,N_1655);
or U6334 (N_6334,N_1336,N_178);
xnor U6335 (N_6335,N_4166,N_4676);
xnor U6336 (N_6336,N_1348,N_3846);
or U6337 (N_6337,N_4995,N_2555);
or U6338 (N_6338,N_2864,N_1780);
nand U6339 (N_6339,N_1488,N_4531);
nor U6340 (N_6340,N_2603,N_3253);
xor U6341 (N_6341,N_4334,N_742);
nor U6342 (N_6342,N_644,N_2815);
nand U6343 (N_6343,N_4478,N_4111);
nor U6344 (N_6344,N_3981,N_329);
xnor U6345 (N_6345,N_2240,N_1777);
nor U6346 (N_6346,N_3203,N_1229);
nand U6347 (N_6347,N_482,N_2944);
nor U6348 (N_6348,N_2446,N_2878);
nor U6349 (N_6349,N_4134,N_3903);
nand U6350 (N_6350,N_2525,N_3667);
xor U6351 (N_6351,N_3891,N_4475);
and U6352 (N_6352,N_4762,N_476);
and U6353 (N_6353,N_1359,N_486);
nor U6354 (N_6354,N_155,N_2344);
and U6355 (N_6355,N_692,N_534);
or U6356 (N_6356,N_417,N_4954);
or U6357 (N_6357,N_812,N_1006);
nor U6358 (N_6358,N_4243,N_4367);
xnor U6359 (N_6359,N_3830,N_613);
or U6360 (N_6360,N_4373,N_4855);
and U6361 (N_6361,N_2338,N_3508);
nor U6362 (N_6362,N_2394,N_1527);
xnor U6363 (N_6363,N_4666,N_805);
xnor U6364 (N_6364,N_3310,N_3792);
and U6365 (N_6365,N_4368,N_2282);
nand U6366 (N_6366,N_3740,N_2957);
or U6367 (N_6367,N_3257,N_2570);
nor U6368 (N_6368,N_1046,N_3342);
xor U6369 (N_6369,N_1233,N_1803);
and U6370 (N_6370,N_4332,N_2313);
or U6371 (N_6371,N_1168,N_2762);
nand U6372 (N_6372,N_1000,N_2939);
and U6373 (N_6373,N_4967,N_4515);
xor U6374 (N_6374,N_2198,N_1896);
xnor U6375 (N_6375,N_3545,N_2646);
and U6376 (N_6376,N_3420,N_2306);
or U6377 (N_6377,N_1686,N_4047);
nand U6378 (N_6378,N_1523,N_4817);
and U6379 (N_6379,N_331,N_1141);
or U6380 (N_6380,N_3628,N_1126);
xnor U6381 (N_6381,N_2831,N_3562);
and U6382 (N_6382,N_1951,N_290);
nand U6383 (N_6383,N_4920,N_4793);
nand U6384 (N_6384,N_4695,N_3320);
or U6385 (N_6385,N_2019,N_4306);
nor U6386 (N_6386,N_1429,N_2988);
and U6387 (N_6387,N_4259,N_3827);
nand U6388 (N_6388,N_227,N_2769);
or U6389 (N_6389,N_4989,N_114);
nor U6390 (N_6390,N_1501,N_3136);
or U6391 (N_6391,N_2055,N_3639);
nor U6392 (N_6392,N_144,N_4383);
nor U6393 (N_6393,N_148,N_4544);
nand U6394 (N_6394,N_3106,N_3597);
xnor U6395 (N_6395,N_2847,N_918);
nor U6396 (N_6396,N_3563,N_1036);
nand U6397 (N_6397,N_1238,N_1755);
or U6398 (N_6398,N_3409,N_4543);
nor U6399 (N_6399,N_4642,N_3498);
nand U6400 (N_6400,N_2637,N_4649);
nor U6401 (N_6401,N_115,N_4266);
nor U6402 (N_6402,N_4026,N_2520);
nand U6403 (N_6403,N_356,N_4596);
xnor U6404 (N_6404,N_2037,N_1886);
and U6405 (N_6405,N_292,N_903);
and U6406 (N_6406,N_3796,N_3372);
nand U6407 (N_6407,N_3593,N_4979);
nand U6408 (N_6408,N_4938,N_4056);
nand U6409 (N_6409,N_1885,N_2768);
nand U6410 (N_6410,N_1162,N_152);
xor U6411 (N_6411,N_493,N_3402);
and U6412 (N_6412,N_3904,N_4976);
nor U6413 (N_6413,N_3780,N_1516);
nand U6414 (N_6414,N_69,N_3964);
nor U6415 (N_6415,N_1892,N_3521);
and U6416 (N_6416,N_4513,N_4457);
nor U6417 (N_6417,N_4292,N_2970);
xor U6418 (N_6418,N_1306,N_4096);
nor U6419 (N_6419,N_1982,N_2857);
xnor U6420 (N_6420,N_78,N_4554);
nand U6421 (N_6421,N_1549,N_316);
nor U6422 (N_6422,N_2848,N_3083);
or U6423 (N_6423,N_4735,N_191);
nor U6424 (N_6424,N_2088,N_784);
nor U6425 (N_6425,N_4016,N_3844);
and U6426 (N_6426,N_1131,N_3900);
or U6427 (N_6427,N_688,N_3004);
xnor U6428 (N_6428,N_506,N_1873);
and U6429 (N_6429,N_1475,N_2427);
xnor U6430 (N_6430,N_2648,N_1155);
and U6431 (N_6431,N_2533,N_2262);
or U6432 (N_6432,N_1417,N_465);
xor U6433 (N_6433,N_3414,N_597);
xor U6434 (N_6434,N_4267,N_539);
or U6435 (N_6435,N_2148,N_3955);
nor U6436 (N_6436,N_538,N_3585);
and U6437 (N_6437,N_528,N_3947);
nand U6438 (N_6438,N_2539,N_3119);
nand U6439 (N_6439,N_2664,N_987);
xnor U6440 (N_6440,N_886,N_4756);
xnor U6441 (N_6441,N_3531,N_3449);
nor U6442 (N_6442,N_3915,N_546);
xor U6443 (N_6443,N_1615,N_4846);
nor U6444 (N_6444,N_2410,N_4529);
or U6445 (N_6445,N_2407,N_283);
nor U6446 (N_6446,N_1999,N_4222);
or U6447 (N_6447,N_3580,N_3870);
nand U6448 (N_6448,N_1623,N_4346);
xnor U6449 (N_6449,N_768,N_107);
xnor U6450 (N_6450,N_1756,N_3690);
nand U6451 (N_6451,N_43,N_2900);
xor U6452 (N_6452,N_28,N_2224);
or U6453 (N_6453,N_2320,N_495);
xnor U6454 (N_6454,N_2997,N_2006);
or U6455 (N_6455,N_15,N_4964);
or U6456 (N_6456,N_653,N_1658);
nand U6457 (N_6457,N_3970,N_4928);
nand U6458 (N_6458,N_3497,N_3475);
nand U6459 (N_6459,N_4151,N_102);
nand U6460 (N_6460,N_702,N_2150);
xor U6461 (N_6461,N_4704,N_2317);
or U6462 (N_6462,N_1271,N_3269);
or U6463 (N_6463,N_1240,N_4264);
xnor U6464 (N_6464,N_3044,N_723);
and U6465 (N_6465,N_2622,N_2152);
xnor U6466 (N_6466,N_22,N_4923);
xnor U6467 (N_6467,N_1258,N_278);
nand U6468 (N_6468,N_2846,N_57);
or U6469 (N_6469,N_1190,N_1393);
or U6470 (N_6470,N_4226,N_1187);
xor U6471 (N_6471,N_3719,N_919);
or U6472 (N_6472,N_434,N_507);
and U6473 (N_6473,N_2269,N_1374);
and U6474 (N_6474,N_2490,N_2535);
nand U6475 (N_6475,N_508,N_2485);
or U6476 (N_6476,N_4614,N_4630);
or U6477 (N_6477,N_4409,N_2332);
xnor U6478 (N_6478,N_1613,N_4853);
and U6479 (N_6479,N_2,N_1132);
nand U6480 (N_6480,N_2479,N_2607);
nor U6481 (N_6481,N_1387,N_826);
and U6482 (N_6482,N_1301,N_87);
and U6483 (N_6483,N_3762,N_928);
or U6484 (N_6484,N_2464,N_2197);
and U6485 (N_6485,N_3456,N_2554);
xnor U6486 (N_6486,N_1112,N_3332);
and U6487 (N_6487,N_518,N_1514);
nand U6488 (N_6488,N_734,N_2062);
and U6489 (N_6489,N_4369,N_1441);
and U6490 (N_6490,N_1032,N_4702);
nor U6491 (N_6491,N_4441,N_2918);
xor U6492 (N_6492,N_3988,N_1818);
and U6493 (N_6493,N_1136,N_3223);
nand U6494 (N_6494,N_3450,N_2194);
nor U6495 (N_6495,N_2252,N_440);
and U6496 (N_6496,N_3494,N_3803);
and U6497 (N_6497,N_3535,N_1851);
or U6498 (N_6498,N_2844,N_2256);
or U6499 (N_6499,N_3784,N_2932);
xor U6500 (N_6500,N_4002,N_4109);
xnor U6501 (N_6501,N_1325,N_814);
xor U6502 (N_6502,N_238,N_478);
nand U6503 (N_6503,N_4677,N_3030);
nor U6504 (N_6504,N_2836,N_2513);
and U6505 (N_6505,N_4129,N_809);
nand U6506 (N_6506,N_1340,N_2940);
or U6507 (N_6507,N_4073,N_1709);
xor U6508 (N_6508,N_1714,N_4177);
nor U6509 (N_6509,N_3398,N_960);
or U6510 (N_6510,N_3505,N_2987);
and U6511 (N_6511,N_2044,N_2230);
nand U6512 (N_6512,N_872,N_1510);
nand U6513 (N_6513,N_3150,N_1400);
xnor U6514 (N_6514,N_612,N_2352);
nand U6515 (N_6515,N_3794,N_4918);
nand U6516 (N_6516,N_2433,N_137);
xor U6517 (N_6517,N_4425,N_3606);
nand U6518 (N_6518,N_4218,N_4613);
xnor U6519 (N_6519,N_1767,N_4080);
nand U6520 (N_6520,N_2129,N_1628);
nor U6521 (N_6521,N_3726,N_1679);
nor U6522 (N_6522,N_46,N_4300);
nor U6523 (N_6523,N_2531,N_2348);
and U6524 (N_6524,N_1351,N_1920);
and U6525 (N_6525,N_3742,N_3880);
and U6526 (N_6526,N_1265,N_2404);
xor U6527 (N_6527,N_2189,N_4562);
or U6528 (N_6528,N_3554,N_705);
xor U6529 (N_6529,N_1944,N_4099);
and U6530 (N_6530,N_4882,N_3753);
xnor U6531 (N_6531,N_4410,N_219);
nor U6532 (N_6532,N_373,N_3451);
nand U6533 (N_6533,N_912,N_624);
and U6534 (N_6534,N_4248,N_2048);
nor U6535 (N_6535,N_991,N_2279);
or U6536 (N_6536,N_422,N_3082);
xor U6537 (N_6537,N_1402,N_3774);
nor U6538 (N_6538,N_1558,N_4052);
xnor U6539 (N_6539,N_2471,N_572);
or U6540 (N_6540,N_4440,N_4595);
xor U6541 (N_6541,N_3729,N_2663);
xor U6542 (N_6542,N_4609,N_638);
or U6543 (N_6543,N_121,N_2860);
and U6544 (N_6544,N_535,N_3301);
and U6545 (N_6545,N_3560,N_4380);
xnor U6546 (N_6546,N_4647,N_4295);
or U6547 (N_6547,N_2457,N_571);
nand U6548 (N_6548,N_3000,N_1894);
and U6549 (N_6549,N_452,N_1443);
nand U6550 (N_6550,N_2745,N_598);
xor U6551 (N_6551,N_3388,N_2699);
and U6552 (N_6552,N_2906,N_2506);
and U6553 (N_6553,N_2744,N_4499);
xor U6554 (N_6554,N_1304,N_2907);
or U6555 (N_6555,N_3607,N_857);
and U6556 (N_6556,N_4094,N_3935);
or U6557 (N_6557,N_4629,N_4193);
and U6558 (N_6558,N_4536,N_2984);
nand U6559 (N_6559,N_1561,N_4899);
nor U6560 (N_6560,N_399,N_4484);
or U6561 (N_6561,N_4937,N_4432);
or U6562 (N_6562,N_2903,N_120);
and U6563 (N_6563,N_1854,N_2858);
nand U6564 (N_6564,N_1156,N_2047);
and U6565 (N_6565,N_2021,N_3131);
nand U6566 (N_6566,N_1611,N_2675);
nand U6567 (N_6567,N_1308,N_3367);
nor U6568 (N_6568,N_1122,N_3235);
xor U6569 (N_6569,N_4350,N_2087);
and U6570 (N_6570,N_4582,N_4909);
xnor U6571 (N_6571,N_681,N_4405);
xor U6572 (N_6572,N_4875,N_1390);
nor U6573 (N_6573,N_4991,N_4213);
nor U6574 (N_6574,N_4001,N_3446);
or U6575 (N_6575,N_2099,N_2843);
nand U6576 (N_6576,N_4683,N_326);
nand U6577 (N_6577,N_344,N_392);
nor U6578 (N_6578,N_81,N_3180);
nand U6579 (N_6579,N_693,N_3247);
xnor U6580 (N_6580,N_2082,N_791);
xnor U6581 (N_6581,N_655,N_2436);
or U6582 (N_6582,N_2484,N_3046);
and U6583 (N_6583,N_247,N_1863);
xor U6584 (N_6584,N_3140,N_2775);
and U6585 (N_6585,N_3722,N_1671);
nor U6586 (N_6586,N_3954,N_3328);
nand U6587 (N_6587,N_1394,N_3809);
nand U6588 (N_6588,N_4493,N_2447);
xor U6589 (N_6589,N_4997,N_3772);
or U6590 (N_6590,N_3187,N_761);
nor U6591 (N_6591,N_4972,N_3626);
or U6592 (N_6592,N_749,N_4549);
xnor U6593 (N_6593,N_1092,N_2315);
and U6594 (N_6594,N_3533,N_1413);
or U6595 (N_6595,N_1966,N_3570);
nor U6596 (N_6596,N_2936,N_4331);
and U6597 (N_6597,N_1784,N_1550);
or U6598 (N_6598,N_2509,N_917);
and U6599 (N_6599,N_4863,N_4838);
nand U6600 (N_6600,N_807,N_829);
and U6601 (N_6601,N_1512,N_4697);
xnor U6602 (N_6602,N_4729,N_2126);
and U6603 (N_6603,N_1703,N_4415);
and U6604 (N_6604,N_4551,N_818);
and U6605 (N_6605,N_4108,N_345);
xnor U6606 (N_6606,N_67,N_894);
nor U6607 (N_6607,N_2890,N_37);
nor U6608 (N_6608,N_3834,N_53);
nor U6609 (N_6609,N_1789,N_1808);
xnor U6610 (N_6610,N_1961,N_3478);
and U6611 (N_6611,N_2494,N_769);
and U6612 (N_6612,N_229,N_3493);
or U6613 (N_6613,N_1772,N_149);
nand U6614 (N_6614,N_2872,N_3093);
nand U6615 (N_6615,N_2854,N_893);
nand U6616 (N_6616,N_1921,N_1328);
and U6617 (N_6617,N_1259,N_4004);
or U6618 (N_6618,N_1354,N_1683);
nor U6619 (N_6619,N_444,N_851);
nand U6620 (N_6620,N_2935,N_3329);
and U6621 (N_6621,N_4800,N_4959);
and U6622 (N_6622,N_65,N_3482);
nand U6623 (N_6623,N_772,N_1763);
or U6624 (N_6624,N_4784,N_172);
or U6625 (N_6625,N_3432,N_3333);
and U6626 (N_6626,N_4724,N_3290);
nor U6627 (N_6627,N_2439,N_4352);
nor U6628 (N_6628,N_2795,N_4283);
xnor U6629 (N_6629,N_4711,N_1330);
xnor U6630 (N_6630,N_4296,N_29);
or U6631 (N_6631,N_1588,N_1290);
nand U6632 (N_6632,N_780,N_1117);
nand U6633 (N_6633,N_4716,N_2894);
nor U6634 (N_6634,N_2284,N_1687);
or U6635 (N_6635,N_2546,N_3280);
or U6636 (N_6636,N_3334,N_3164);
nor U6637 (N_6637,N_3911,N_3926);
nor U6638 (N_6638,N_3599,N_690);
nand U6639 (N_6639,N_2802,N_1196);
xnor U6640 (N_6640,N_1287,N_1573);
xnor U6641 (N_6641,N_4431,N_367);
nor U6642 (N_6642,N_2561,N_967);
or U6643 (N_6643,N_4782,N_413);
nand U6644 (N_6644,N_446,N_4781);
or U6645 (N_6645,N_2754,N_1627);
nor U6646 (N_6646,N_3576,N_4652);
or U6647 (N_6647,N_4803,N_1040);
or U6648 (N_6648,N_4924,N_4714);
nor U6649 (N_6649,N_173,N_2323);
nor U6650 (N_6650,N_86,N_3694);
xnor U6651 (N_6651,N_2466,N_4453);
and U6652 (N_6652,N_632,N_2283);
and U6653 (N_6653,N_4608,N_3968);
nand U6654 (N_6654,N_1088,N_4228);
xnor U6655 (N_6655,N_2226,N_1576);
nor U6656 (N_6656,N_3116,N_1688);
xnor U6657 (N_6657,N_2512,N_1041);
xnor U6658 (N_6658,N_4110,N_4359);
nor U6659 (N_6659,N_74,N_1202);
and U6660 (N_6660,N_551,N_4576);
nand U6661 (N_6661,N_162,N_4651);
xor U6662 (N_6662,N_2901,N_515);
nand U6663 (N_6663,N_3649,N_2286);
or U6664 (N_6664,N_694,N_3577);
xnor U6665 (N_6665,N_3872,N_3712);
nand U6666 (N_6666,N_4114,N_2726);
or U6667 (N_6667,N_2556,N_2295);
and U6668 (N_6668,N_240,N_4192);
or U6669 (N_6669,N_3547,N_4437);
nor U6670 (N_6670,N_2124,N_3111);
xnor U6671 (N_6671,N_4760,N_882);
nand U6672 (N_6672,N_4040,N_2211);
xor U6673 (N_6673,N_2029,N_1824);
or U6674 (N_6674,N_4895,N_715);
or U6675 (N_6675,N_1584,N_3575);
xnor U6676 (N_6676,N_914,N_2203);
or U6677 (N_6677,N_4474,N_2058);
and U6678 (N_6678,N_2325,N_3818);
nand U6679 (N_6679,N_1275,N_1864);
xor U6680 (N_6680,N_2600,N_3168);
xor U6681 (N_6681,N_4205,N_3669);
or U6682 (N_6682,N_4091,N_2873);
and U6683 (N_6683,N_3184,N_3951);
xnor U6684 (N_6684,N_4985,N_4738);
and U6685 (N_6685,N_2008,N_3770);
xnor U6686 (N_6686,N_4755,N_2218);
nor U6687 (N_6687,N_1380,N_2227);
and U6688 (N_6688,N_3512,N_4607);
nand U6689 (N_6689,N_4975,N_1012);
xor U6690 (N_6690,N_1897,N_3126);
nor U6691 (N_6691,N_855,N_3270);
or U6692 (N_6692,N_4232,N_1320);
nor U6693 (N_6693,N_992,N_3691);
or U6694 (N_6694,N_4433,N_4486);
xnor U6695 (N_6695,N_2142,N_4260);
and U6696 (N_6696,N_1673,N_2702);
nand U6697 (N_6697,N_1075,N_3330);
or U6698 (N_6698,N_2566,N_2964);
and U6699 (N_6699,N_750,N_296);
nor U6700 (N_6700,N_4556,N_2249);
or U6701 (N_6701,N_556,N_2705);
nor U6702 (N_6702,N_4305,N_4520);
and U6703 (N_6703,N_3965,N_3921);
nor U6704 (N_6704,N_897,N_720);
xnor U6705 (N_6705,N_664,N_4302);
and U6706 (N_6706,N_2395,N_1016);
nand U6707 (N_6707,N_117,N_1620);
xor U6708 (N_6708,N_4466,N_4179);
or U6709 (N_6709,N_3771,N_589);
and U6710 (N_6710,N_4148,N_1790);
or U6711 (N_6711,N_3064,N_2644);
or U6712 (N_6712,N_4281,N_4900);
nor U6713 (N_6713,N_1426,N_1548);
or U6714 (N_6714,N_1281,N_777);
nor U6715 (N_6715,N_3908,N_3133);
nor U6716 (N_6716,N_2056,N_2912);
nor U6717 (N_6717,N_1378,N_460);
nor U6718 (N_6718,N_933,N_752);
and U6719 (N_6719,N_521,N_4681);
and U6720 (N_6720,N_212,N_299);
or U6721 (N_6721,N_128,N_695);
xor U6722 (N_6722,N_4060,N_362);
nor U6723 (N_6723,N_3407,N_828);
and U6724 (N_6724,N_4919,N_2938);
nand U6725 (N_6725,N_402,N_3122);
and U6726 (N_6726,N_2028,N_217);
nand U6727 (N_6727,N_3211,N_1345);
nand U6728 (N_6728,N_309,N_736);
and U6729 (N_6729,N_1668,N_2652);
nor U6730 (N_6730,N_4120,N_3715);
xnor U6731 (N_6731,N_1989,N_474);
xor U6732 (N_6732,N_3857,N_2849);
nor U6733 (N_6733,N_2915,N_4943);
and U6734 (N_6734,N_1797,N_327);
or U6735 (N_6735,N_1309,N_1876);
nor U6736 (N_6736,N_4482,N_3170);
nand U6737 (N_6737,N_4219,N_2472);
nand U6738 (N_6738,N_529,N_4498);
xnor U6739 (N_6739,N_2145,N_4022);
xnor U6740 (N_6740,N_4353,N_4585);
nand U6741 (N_6741,N_663,N_2877);
or U6742 (N_6742,N_3458,N_4641);
nor U6743 (N_6743,N_2614,N_146);
xnor U6744 (N_6744,N_4388,N_1158);
xor U6745 (N_6745,N_2975,N_1478);
or U6746 (N_6746,N_56,N_746);
nand U6747 (N_6747,N_4031,N_744);
nand U6748 (N_6748,N_2720,N_4957);
nand U6749 (N_6749,N_3360,N_4511);
xor U6750 (N_6750,N_1891,N_725);
nand U6751 (N_6751,N_4054,N_2065);
nand U6752 (N_6752,N_118,N_1602);
and U6753 (N_6753,N_2838,N_404);
xnor U6754 (N_6754,N_1962,N_2990);
or U6755 (N_6755,N_372,N_1870);
xor U6756 (N_6756,N_2097,N_135);
nand U6757 (N_6757,N_2370,N_1493);
nand U6758 (N_6758,N_514,N_450);
nor U6759 (N_6759,N_1048,N_3468);
xnor U6760 (N_6760,N_837,N_1211);
nand U6761 (N_6761,N_671,N_203);
or U6762 (N_6762,N_2870,N_3528);
and U6763 (N_6763,N_4058,N_54);
nand U6764 (N_6764,N_1074,N_408);
xor U6765 (N_6765,N_1236,N_2171);
and U6766 (N_6766,N_89,N_522);
or U6767 (N_6767,N_4850,N_4115);
and U6768 (N_6768,N_1817,N_2096);
nand U6769 (N_6769,N_4661,N_19);
nor U6770 (N_6770,N_1819,N_3821);
nor U6771 (N_6771,N_1180,N_4133);
and U6772 (N_6772,N_1472,N_305);
or U6773 (N_6773,N_4312,N_1139);
and U6774 (N_6774,N_4371,N_1247);
or U6775 (N_6775,N_1859,N_1843);
nor U6776 (N_6776,N_4136,N_4117);
nand U6777 (N_6777,N_2135,N_2351);
and U6778 (N_6778,N_1065,N_4483);
xor U6779 (N_6779,N_2274,N_915);
nand U6780 (N_6780,N_3810,N_1952);
nor U6781 (N_6781,N_2659,N_4348);
or U6782 (N_6782,N_937,N_2840);
nor U6783 (N_6783,N_4946,N_747);
xor U6784 (N_6784,N_4981,N_3884);
or U6785 (N_6785,N_4375,N_1834);
nand U6786 (N_6786,N_580,N_3102);
and U6787 (N_6787,N_1967,N_4917);
nor U6788 (N_6788,N_4968,N_4603);
nor U6789 (N_6789,N_4149,N_1140);
or U6790 (N_6790,N_590,N_2331);
xnor U6791 (N_6791,N_206,N_1406);
nand U6792 (N_6792,N_4313,N_4185);
nor U6793 (N_6793,N_2829,N_1922);
or U6794 (N_6794,N_4411,N_1530);
and U6795 (N_6795,N_3110,N_1343);
nor U6796 (N_6796,N_3877,N_40);
xnor U6797 (N_6797,N_2621,N_3369);
or U6798 (N_6798,N_1974,N_2805);
or U6799 (N_6799,N_469,N_4789);
nand U6800 (N_6800,N_2966,N_4802);
nand U6801 (N_6801,N_1984,N_1884);
nand U6802 (N_6802,N_3271,N_816);
nor U6803 (N_6803,N_2149,N_2656);
or U6804 (N_6804,N_2100,N_1807);
nor U6805 (N_6805,N_1282,N_4376);
xor U6806 (N_6806,N_2257,N_463);
nand U6807 (N_6807,N_2202,N_2287);
nor U6808 (N_6808,N_2609,N_4435);
nand U6809 (N_6809,N_2770,N_2585);
nand U6810 (N_6810,N_1205,N_4701);
or U6811 (N_6811,N_423,N_1384);
and U6812 (N_6812,N_1160,N_4211);
and U6813 (N_6813,N_2102,N_3578);
and U6814 (N_6814,N_2792,N_1811);
nor U6815 (N_6815,N_3590,N_2729);
xor U6816 (N_6816,N_4468,N_3159);
xnor U6817 (N_6817,N_1366,N_100);
nand U6818 (N_6818,N_3029,N_3551);
xnor U6819 (N_6819,N_1433,N_2653);
and U6820 (N_6820,N_1806,N_3123);
nand U6821 (N_6821,N_3085,N_4017);
xor U6822 (N_6822,N_691,N_4725);
and U6823 (N_6823,N_2409,N_2943);
and U6824 (N_6824,N_4942,N_4610);
xnor U6825 (N_6825,N_3525,N_1138);
nor U6826 (N_6826,N_2201,N_2183);
or U6827 (N_6827,N_2229,N_4897);
and U6828 (N_6828,N_2503,N_1272);
and U6829 (N_6829,N_4885,N_4321);
xnor U6830 (N_6830,N_2881,N_3396);
nand U6831 (N_6831,N_2254,N_4462);
nor U6832 (N_6832,N_4828,N_248);
nand U6833 (N_6833,N_1099,N_2015);
xnor U6834 (N_6834,N_2671,N_3057);
nand U6835 (N_6835,N_4255,N_4560);
or U6836 (N_6836,N_2020,N_2368);
and U6837 (N_6837,N_3461,N_3274);
or U6838 (N_6838,N_2760,N_3266);
or U6839 (N_6839,N_4349,N_968);
nor U6840 (N_6840,N_4815,N_2456);
nand U6841 (N_6841,N_4664,N_4589);
xnor U6842 (N_6842,N_510,N_1334);
and U6843 (N_6843,N_2741,N_2510);
or U6844 (N_6844,N_2281,N_1713);
xor U6845 (N_6845,N_3028,N_4657);
or U6846 (N_6846,N_3154,N_4330);
nor U6847 (N_6847,N_348,N_4231);
nor U6848 (N_6848,N_4420,N_3321);
and U6849 (N_6849,N_2003,N_1499);
nand U6850 (N_6850,N_1591,N_527);
xnor U6851 (N_6851,N_2382,N_3484);
xor U6852 (N_6852,N_1451,N_1357);
nor U6853 (N_6853,N_3201,N_403);
or U6854 (N_6854,N_4706,N_1927);
xor U6855 (N_6855,N_793,N_1033);
xnor U6856 (N_6856,N_4208,N_1469);
or U6857 (N_6857,N_2956,N_1327);
xnor U6858 (N_6858,N_4732,N_1452);
nand U6859 (N_6859,N_168,N_4291);
and U6860 (N_6860,N_3546,N_1292);
nor U6861 (N_6861,N_1347,N_1214);
or U6862 (N_6862,N_3121,N_215);
nand U6863 (N_6863,N_1768,N_1955);
nor U6864 (N_6864,N_4868,N_4480);
or U6865 (N_6865,N_1339,N_2662);
xor U6866 (N_6866,N_1153,N_281);
nor U6867 (N_6867,N_1572,N_1880);
and U6868 (N_6868,N_3573,N_774);
or U6869 (N_6869,N_184,N_2771);
and U6870 (N_6870,N_2314,N_480);
or U6871 (N_6871,N_443,N_2213);
nand U6872 (N_6872,N_287,N_4730);
or U6873 (N_6873,N_3945,N_3379);
and U6874 (N_6874,N_902,N_1676);
or U6875 (N_6875,N_1067,N_2891);
nand U6876 (N_6876,N_4125,N_3602);
xnor U6877 (N_6877,N_2748,N_3124);
nand U6878 (N_6878,N_3058,N_500);
nand U6879 (N_6879,N_1482,N_2639);
or U6880 (N_6880,N_2657,N_1844);
nand U6881 (N_6881,N_2948,N_3325);
nand U6882 (N_6882,N_1607,N_4391);
nand U6883 (N_6883,N_888,N_4207);
nand U6884 (N_6884,N_3413,N_4854);
nor U6885 (N_6885,N_4915,N_2025);
and U6886 (N_6886,N_2085,N_3923);
xor U6887 (N_6887,N_3741,N_4417);
or U6888 (N_6888,N_3074,N_2928);
and U6889 (N_6889,N_4337,N_1682);
nor U6890 (N_6890,N_3434,N_2749);
nand U6891 (N_6891,N_4999,N_2031);
xor U6892 (N_6892,N_4364,N_3496);
nand U6893 (N_6893,N_4234,N_4097);
and U6894 (N_6894,N_2336,N_1310);
and U6895 (N_6895,N_4774,N_4809);
xor U6896 (N_6896,N_490,N_63);
xnor U6897 (N_6897,N_1232,N_1317);
nand U6898 (N_6898,N_3031,N_1200);
nand U6899 (N_6899,N_66,N_1185);
nand U6900 (N_6900,N_231,N_2480);
nand U6901 (N_6901,N_3739,N_130);
or U6902 (N_6902,N_2027,N_3305);
nand U6903 (N_6903,N_3009,N_1101);
and U6904 (N_6904,N_3660,N_4852);
xnor U6905 (N_6905,N_2694,N_1746);
nor U6906 (N_6906,N_1376,N_610);
nand U6907 (N_6907,N_2443,N_2820);
nand U6908 (N_6908,N_1637,N_2651);
xor U6909 (N_6909,N_4581,N_1154);
nand U6910 (N_6910,N_1080,N_1910);
nor U6911 (N_6911,N_4632,N_42);
nand U6912 (N_6912,N_347,N_3847);
nand U6913 (N_6913,N_4713,N_4030);
nor U6914 (N_6914,N_3220,N_1590);
nor U6915 (N_6915,N_3816,N_3848);
or U6916 (N_6916,N_2405,N_4404);
xor U6917 (N_6917,N_4238,N_4237);
nor U6918 (N_6918,N_2051,N_473);
nor U6919 (N_6919,N_3565,N_825);
nand U6920 (N_6920,N_497,N_3507);
nand U6921 (N_6921,N_4616,N_1728);
xor U6922 (N_6922,N_4172,N_2985);
nor U6923 (N_6923,N_555,N_1893);
or U6924 (N_6924,N_2052,N_661);
nand U6925 (N_6925,N_1659,N_2498);
nor U6926 (N_6926,N_3481,N_1014);
nor U6927 (N_6927,N_3229,N_3889);
nor U6928 (N_6928,N_1635,N_2276);
xor U6929 (N_6929,N_4659,N_433);
nand U6930 (N_6930,N_4623,N_1778);
nor U6931 (N_6931,N_1917,N_3206);
nand U6932 (N_6932,N_2363,N_1234);
nand U6933 (N_6933,N_3756,N_3445);
nand U6934 (N_6934,N_4197,N_258);
nand U6935 (N_6935,N_4163,N_462);
and U6936 (N_6936,N_4430,N_1730);
or U6937 (N_6937,N_689,N_4718);
and U6938 (N_6938,N_2596,N_3300);
nor U6939 (N_6939,N_4905,N_3699);
nor U6940 (N_6940,N_704,N_3937);
xnor U6941 (N_6941,N_3171,N_4950);
nand U6942 (N_6942,N_3969,N_3027);
nor U6943 (N_6943,N_701,N_2239);
nand U6944 (N_6944,N_1212,N_273);
or U6945 (N_6945,N_4518,N_62);
or U6946 (N_6946,N_1734,N_3864);
nand U6947 (N_6947,N_2910,N_1993);
nand U6948 (N_6948,N_3050,N_4018);
nand U6949 (N_6949,N_3197,N_845);
nand U6950 (N_6950,N_2337,N_3163);
or U6951 (N_6951,N_3294,N_4076);
nand U6952 (N_6952,N_416,N_3063);
nor U6953 (N_6953,N_1822,N_4048);
and U6954 (N_6954,N_4974,N_1268);
and U6955 (N_6955,N_481,N_2799);
and U6956 (N_6956,N_617,N_4836);
xor U6957 (N_6957,N_3737,N_424);
xor U6958 (N_6958,N_3400,N_4872);
xor U6959 (N_6959,N_4775,N_1391);
and U6960 (N_6960,N_3708,N_3720);
xnor U6961 (N_6961,N_1825,N_2209);
or U6962 (N_6962,N_2545,N_4601);
xor U6963 (N_6963,N_3993,N_358);
nand U6964 (N_6964,N_4617,N_943);
and U6965 (N_6965,N_239,N_3618);
nand U6966 (N_6966,N_2590,N_3043);
or U6967 (N_6967,N_2347,N_93);
nor U6968 (N_6968,N_4105,N_2765);
nand U6969 (N_6969,N_4075,N_4063);
nor U6970 (N_6970,N_277,N_3161);
and U6971 (N_6971,N_2267,N_3096);
or U6972 (N_6972,N_2106,N_3849);
or U6973 (N_6973,N_342,N_225);
nor U6974 (N_6974,N_3192,N_532);
nor U6975 (N_6975,N_2460,N_2333);
or U6976 (N_6976,N_85,N_639);
and U6977 (N_6977,N_4818,N_2587);
or U6978 (N_6978,N_2634,N_4252);
nor U6979 (N_6979,N_3352,N_2221);
xnor U6980 (N_6980,N_936,N_970);
nor U6981 (N_6981,N_397,N_226);
xor U6982 (N_6982,N_1474,N_3927);
or U6983 (N_6983,N_411,N_4778);
nand U6984 (N_6984,N_1852,N_2032);
and U6985 (N_6985,N_2217,N_1448);
nor U6986 (N_6986,N_3684,N_4393);
and U6987 (N_6987,N_202,N_246);
nand U6988 (N_6988,N_2523,N_2120);
or U6989 (N_6989,N_1855,N_1736);
nand U6990 (N_6990,N_4399,N_3224);
xor U6991 (N_6991,N_1629,N_142);
nand U6992 (N_6992,N_1721,N_2856);
and U6993 (N_6993,N_1225,N_3686);
nand U6994 (N_6994,N_321,N_3624);
nor U6995 (N_6995,N_4473,N_365);
or U6996 (N_6996,N_18,N_1652);
and U6997 (N_6997,N_1023,N_3895);
nor U6998 (N_6998,N_2947,N_3519);
xor U6999 (N_6999,N_4130,N_3130);
nor U7000 (N_7000,N_4168,N_3949);
xor U7001 (N_7001,N_4500,N_3053);
nand U7002 (N_7002,N_2342,N_1965);
and U7003 (N_7003,N_4156,N_4682);
nor U7004 (N_7004,N_4051,N_3335);
and U7005 (N_7005,N_4216,N_3869);
nor U7006 (N_7006,N_1879,N_1485);
xnor U7007 (N_7007,N_304,N_1842);
or U7008 (N_7008,N_3510,N_4721);
xnor U7009 (N_7009,N_4345,N_3390);
nor U7010 (N_7010,N_4307,N_4436);
or U7011 (N_7011,N_2288,N_3540);
xnor U7012 (N_7012,N_346,N_3148);
nand U7013 (N_7013,N_2441,N_3092);
or U7014 (N_7014,N_1013,N_4530);
nor U7015 (N_7015,N_771,N_2592);
nor U7016 (N_7016,N_618,N_3267);
or U7017 (N_7017,N_1219,N_4263);
and U7018 (N_7018,N_52,N_4354);
or U7019 (N_7019,N_2398,N_948);
nor U7020 (N_7020,N_361,N_352);
xnor U7021 (N_7021,N_71,N_1569);
nor U7022 (N_7022,N_3931,N_1338);
and U7023 (N_7023,N_3683,N_1813);
and U7024 (N_7024,N_944,N_2892);
xor U7025 (N_7025,N_2164,N_3059);
and U7026 (N_7026,N_2075,N_2011);
xnor U7027 (N_7027,N_3967,N_2450);
and U7028 (N_7028,N_4690,N_4454);
and U7029 (N_7029,N_1423,N_727);
nand U7030 (N_7030,N_3732,N_4563);
or U7031 (N_7031,N_3297,N_2682);
nand U7032 (N_7032,N_1715,N_4309);
nand U7033 (N_7033,N_2989,N_302);
or U7034 (N_7034,N_3094,N_3386);
or U7035 (N_7035,N_1371,N_1454);
nand U7036 (N_7036,N_297,N_3466);
and U7037 (N_7037,N_3476,N_3826);
nand U7038 (N_7038,N_3313,N_842);
nand U7039 (N_7039,N_4574,N_1305);
xnor U7040 (N_7040,N_143,N_1606);
or U7041 (N_7041,N_1323,N_4107);
xor U7042 (N_7042,N_2551,N_3842);
nor U7043 (N_7043,N_591,N_3678);
nor U7044 (N_7044,N_2166,N_2054);
or U7045 (N_7045,N_1975,N_519);
xnor U7046 (N_7046,N_2774,N_4902);
xnor U7047 (N_7047,N_1086,N_6);
nor U7048 (N_7048,N_523,N_652);
nor U7049 (N_7049,N_4325,N_741);
nor U7050 (N_7050,N_2885,N_338);
xnor U7051 (N_7051,N_96,N_3088);
xor U7052 (N_7052,N_2442,N_4806);
nand U7053 (N_7053,N_494,N_611);
or U7054 (N_7054,N_2214,N_3219);
nor U7055 (N_7055,N_2473,N_525);
nor U7056 (N_7056,N_3725,N_4988);
or U7057 (N_7057,N_2296,N_3823);
nand U7058 (N_7058,N_1504,N_1718);
nor U7059 (N_7059,N_3232,N_673);
or U7060 (N_7060,N_966,N_754);
and U7061 (N_7061,N_2517,N_1621);
or U7062 (N_7062,N_526,N_1009);
and U7063 (N_7063,N_47,N_475);
and U7064 (N_7064,N_2665,N_2415);
or U7065 (N_7065,N_3713,N_1792);
or U7066 (N_7066,N_4119,N_4215);
and U7067 (N_7067,N_2304,N_3001);
and U7068 (N_7068,N_606,N_3584);
and U7069 (N_7069,N_2358,N_2488);
nand U7070 (N_7070,N_878,N_2417);
and U7071 (N_7071,N_4880,N_1144);
or U7072 (N_7072,N_1889,N_2378);
and U7073 (N_7073,N_3793,N_2515);
nor U7074 (N_7074,N_3825,N_4506);
xnor U7075 (N_7075,N_2467,N_4043);
xnor U7076 (N_7076,N_1412,N_3385);
and U7077 (N_7077,N_930,N_2095);
and U7078 (N_7078,N_3113,N_2896);
nor U7079 (N_7079,N_3795,N_1383);
or U7080 (N_7080,N_3881,N_2616);
or U7081 (N_7081,N_4162,N_3883);
or U7082 (N_7082,N_1150,N_3668);
xor U7083 (N_7083,N_487,N_4338);
or U7084 (N_7084,N_4427,N_3788);
and U7085 (N_7085,N_4336,N_4230);
and U7086 (N_7086,N_4003,N_2809);
and U7087 (N_7087,N_2780,N_3357);
nor U7088 (N_7088,N_997,N_2324);
nor U7089 (N_7089,N_4315,N_4842);
xnor U7090 (N_7090,N_1307,N_767);
nand U7091 (N_7091,N_3284,N_1123);
and U7092 (N_7092,N_3152,N_2196);
nor U7093 (N_7093,N_1815,N_2576);
xor U7094 (N_7094,N_3454,N_4525);
and U7095 (N_7095,N_2541,N_3246);
or U7096 (N_7096,N_83,N_3706);
nor U7097 (N_7097,N_2674,N_1245);
or U7098 (N_7098,N_3370,N_3323);
or U7099 (N_7099,N_4820,N_2619);
nor U7100 (N_7100,N_3011,N_4679);
and U7101 (N_7101,N_4085,N_1061);
nand U7102 (N_7102,N_2222,N_789);
or U7103 (N_7103,N_2804,N_3479);
or U7104 (N_7104,N_4414,N_3076);
or U7105 (N_7105,N_1186,N_3622);
nand U7106 (N_7106,N_3657,N_2737);
and U7107 (N_7107,N_1226,N_4449);
xor U7108 (N_7108,N_877,N_3412);
nor U7109 (N_7109,N_4196,N_4906);
nand U7110 (N_7110,N_1,N_2193);
nor U7111 (N_7111,N_2111,N_1866);
and U7112 (N_7112,N_4103,N_79);
nand U7113 (N_7113,N_4528,N_4861);
nand U7114 (N_7114,N_4401,N_4088);
nand U7115 (N_7115,N_156,N_3914);
and U7116 (N_7116,N_4289,N_3394);
nand U7117 (N_7117,N_4150,N_3404);
and U7118 (N_7118,N_2842,N_1595);
xor U7119 (N_7119,N_998,N_2677);
and U7120 (N_7120,N_3950,N_745);
and U7121 (N_7121,N_4939,N_3309);
nand U7122 (N_7122,N_1017,N_965);
and U7123 (N_7123,N_3600,N_3128);
nand U7124 (N_7124,N_1410,N_849);
and U7125 (N_7125,N_4663,N_3587);
and U7126 (N_7126,N_3633,N_2547);
or U7127 (N_7127,N_4825,N_3115);
nor U7128 (N_7128,N_563,N_2502);
and U7129 (N_7129,N_1484,N_2273);
xor U7130 (N_7130,N_732,N_3381);
or U7131 (N_7131,N_4132,N_3676);
and U7132 (N_7132,N_658,N_190);
or U7133 (N_7133,N_971,N_2983);
xor U7134 (N_7134,N_2911,N_1560);
xnor U7135 (N_7135,N_3299,N_2549);
or U7136 (N_7136,N_4833,N_3256);
nor U7137 (N_7137,N_2781,N_2184);
nand U7138 (N_7138,N_267,N_4978);
xor U7139 (N_7139,N_4734,N_710);
and U7140 (N_7140,N_2357,N_4783);
or U7141 (N_7141,N_3663,N_4285);
xor U7142 (N_7142,N_2386,N_4072);
nand U7143 (N_7143,N_436,N_1355);
or U7144 (N_7144,N_4731,N_2732);
nor U7145 (N_7145,N_2246,N_2714);
or U7146 (N_7146,N_1770,N_3188);
or U7147 (N_7147,N_3375,N_2521);
nand U7148 (N_7148,N_4055,N_2867);
or U7149 (N_7149,N_2162,N_214);
xnor U7150 (N_7150,N_2991,N_2655);
or U7151 (N_7151,N_2598,N_3652);
and U7152 (N_7152,N_3711,N_4381);
and U7153 (N_7153,N_4421,N_1059);
xnor U7154 (N_7154,N_106,N_1507);
nand U7155 (N_7155,N_1986,N_2952);
nor U7156 (N_7156,N_1570,N_470);
xor U7157 (N_7157,N_2962,N_2574);
xnor U7158 (N_7158,N_3957,N_3359);
or U7159 (N_7159,N_2893,N_295);
or U7160 (N_7160,N_1912,N_4532);
and U7161 (N_7161,N_2354,N_2704);
or U7162 (N_7162,N_2902,N_3383);
nand U7163 (N_7163,N_4250,N_2343);
nand U7164 (N_7164,N_4013,N_1720);
nor U7165 (N_7165,N_4444,N_3433);
or U7166 (N_7166,N_4750,N_32);
and U7167 (N_7167,N_2495,N_193);
or U7168 (N_7168,N_3426,N_1077);
and U7169 (N_7169,N_3871,N_185);
xor U7170 (N_7170,N_2266,N_2181);
nand U7171 (N_7171,N_4654,N_3107);
xnor U7172 (N_7172,N_4429,N_1331);
or U7173 (N_7173,N_2641,N_4246);
xor U7174 (N_7174,N_1704,N_2505);
or U7175 (N_7175,N_770,N_1791);
xor U7176 (N_7176,N_4489,N_1833);
nor U7177 (N_7177,N_4786,N_1836);
nand U7178 (N_7178,N_2215,N_823);
nor U7179 (N_7179,N_4823,N_2474);
or U7180 (N_7180,N_2814,N_4426);
nor U7181 (N_7181,N_1279,N_88);
xnor U7182 (N_7182,N_2080,N_1252);
and U7183 (N_7183,N_4860,N_4229);
and U7184 (N_7184,N_687,N_3873);
nor U7185 (N_7185,N_2101,N_787);
and U7186 (N_7186,N_1592,N_4282);
nor U7187 (N_7187,N_2669,N_1875);
nand U7188 (N_7188,N_2169,N_1003);
nor U7189 (N_7189,N_4355,N_4253);
nand U7190 (N_7190,N_3567,N_249);
xor U7191 (N_7191,N_4945,N_700);
nor U7192 (N_7192,N_2691,N_3941);
xnor U7193 (N_7193,N_405,N_3248);
nor U7194 (N_7194,N_626,N_2929);
xnor U7195 (N_7195,N_3249,N_4584);
and U7196 (N_7196,N_940,N_3265);
nor U7197 (N_7197,N_1477,N_3596);
and U7198 (N_7198,N_4746,N_2091);
nand U7199 (N_7199,N_858,N_3109);
nand U7200 (N_7200,N_2967,N_2261);
or U7201 (N_7201,N_4396,N_4174);
and U7202 (N_7202,N_3311,N_3837);
and U7203 (N_7203,N_4794,N_2476);
nor U7204 (N_7204,N_1932,N_1937);
and U7205 (N_7205,N_186,N_2755);
nor U7206 (N_7206,N_4059,N_1261);
or U7207 (N_7207,N_2728,N_733);
xor U7208 (N_7208,N_371,N_2381);
nand U7209 (N_7209,N_2683,N_1264);
nor U7210 (N_7210,N_3174,N_2819);
nand U7211 (N_7211,N_2079,N_2489);
or U7212 (N_7212,N_2707,N_1072);
or U7213 (N_7213,N_2735,N_3744);
nor U7214 (N_7214,N_718,N_2544);
or U7215 (N_7215,N_1255,N_270);
xor U7216 (N_7216,N_3569,N_1991);
xor U7217 (N_7217,N_4503,N_1528);
xnor U7218 (N_7218,N_1487,N_1318);
nor U7219 (N_7219,N_2816,N_504);
xnor U7220 (N_7220,N_389,N_44);
nand U7221 (N_7221,N_3199,N_1222);
xor U7222 (N_7222,N_3304,N_2042);
and U7223 (N_7223,N_4748,N_1625);
nor U7224 (N_7224,N_1284,N_3238);
xnor U7225 (N_7225,N_1743,N_4303);
and U7226 (N_7226,N_4633,N_3179);
nand U7227 (N_7227,N_2050,N_1450);
or U7228 (N_7228,N_3071,N_2185);
nand U7229 (N_7229,N_1299,N_3865);
nor U7230 (N_7230,N_1431,N_2002);
xnor U7231 (N_7231,N_1653,N_2061);
and U7232 (N_7232,N_938,N_4893);
nor U7233 (N_7233,N_4921,N_1923);
nor U7234 (N_7234,N_4570,N_2715);
nor U7235 (N_7235,N_4494,N_419);
nand U7236 (N_7236,N_2580,N_2821);
and U7237 (N_7237,N_4955,N_4167);
nand U7238 (N_7238,N_4245,N_464);
nand U7239 (N_7239,N_3349,N_557);
or U7240 (N_7240,N_2119,N_395);
nand U7241 (N_7241,N_4741,N_2330);
xnor U7242 (N_7242,N_4488,N_679);
and U7243 (N_7243,N_1203,N_2403);
or U7244 (N_7244,N_2617,N_4615);
or U7245 (N_7245,N_4648,N_3452);
nand U7246 (N_7246,N_4829,N_4827);
nor U7247 (N_7247,N_4685,N_4592);
nor U7248 (N_7248,N_4268,N_1095);
or U7249 (N_7249,N_4184,N_36);
nand U7250 (N_7250,N_1407,N_2305);
nor U7251 (N_7251,N_4622,N_994);
or U7252 (N_7252,N_1518,N_3303);
and U7253 (N_7253,N_2063,N_1751);
and U7254 (N_7254,N_1531,N_3023);
nand U7255 (N_7255,N_3887,N_4588);
or U7256 (N_7256,N_853,N_4434);
or U7257 (N_7257,N_2275,N_3153);
and U7258 (N_7258,N_2632,N_3775);
nand U7259 (N_7259,N_907,N_2458);
nor U7260 (N_7260,N_4621,N_3350);
and U7261 (N_7261,N_3855,N_4586);
xor U7262 (N_7262,N_4065,N_2685);
nor U7263 (N_7263,N_3435,N_4165);
xor U7264 (N_7264,N_431,N_1244);
and U7265 (N_7265,N_2658,N_4660);
and U7266 (N_7266,N_2030,N_1109);
nor U7267 (N_7267,N_4744,N_1902);
or U7268 (N_7268,N_1189,N_3289);
and U7269 (N_7269,N_2862,N_1416);
xor U7270 (N_7270,N_1163,N_393);
or U7271 (N_7271,N_2817,N_2784);
nand U7272 (N_7272,N_1295,N_4587);
nand U7273 (N_7273,N_4751,N_2128);
or U7274 (N_7274,N_192,N_3337);
and U7275 (N_7275,N_1924,N_2499);
nand U7276 (N_7276,N_1871,N_4153);
xnor U7277 (N_7277,N_1608,N_276);
and U7278 (N_7278,N_2462,N_3490);
xnor U7279 (N_7279,N_2478,N_282);
xor U7280 (N_7280,N_3892,N_929);
and U7281 (N_7281,N_2786,N_763);
nor U7282 (N_7282,N_1051,N_1103);
nor U7283 (N_7283,N_4206,N_4254);
or U7284 (N_7284,N_4261,N_3653);
xor U7285 (N_7285,N_4139,N_3804);
and U7286 (N_7286,N_3278,N_2426);
nor U7287 (N_7287,N_1677,N_3165);
xnor U7288 (N_7288,N_783,N_4227);
nand U7289 (N_7289,N_4,N_2982);
or U7290 (N_7290,N_3718,N_2294);
or U7291 (N_7291,N_838,N_4200);
xnor U7292 (N_7292,N_2811,N_1206);
or U7293 (N_7293,N_2272,N_543);
and U7294 (N_7294,N_2053,N_8);
and U7295 (N_7295,N_3091,N_1439);
nor U7296 (N_7296,N_3559,N_2968);
nor U7297 (N_7297,N_2602,N_1329);
nor U7298 (N_7298,N_3319,N_3132);
xnor U7299 (N_7299,N_650,N_3137);
or U7300 (N_7300,N_566,N_927);
and U7301 (N_7301,N_595,N_3552);
xor U7302 (N_7302,N_454,N_2083);
or U7303 (N_7303,N_3534,N_4891);
or U7304 (N_7304,N_792,N_3555);
and U7305 (N_7305,N_1847,N_1246);
nand U7306 (N_7306,N_1858,N_4526);
nor U7307 (N_7307,N_2797,N_622);
nand U7308 (N_7308,N_867,N_881);
nor U7309 (N_7309,N_167,N_3019);
nand U7310 (N_7310,N_3382,N_322);
nor U7311 (N_7311,N_4122,N_123);
xor U7312 (N_7312,N_4155,N_3654);
and U7313 (N_7313,N_974,N_2385);
nand U7314 (N_7314,N_2310,N_4546);
nor U7315 (N_7315,N_570,N_3990);
or U7316 (N_7316,N_2243,N_1055);
or U7317 (N_7317,N_2955,N_4538);
xnor U7318 (N_7318,N_765,N_3348);
or U7319 (N_7319,N_3532,N_4025);
nor U7320 (N_7320,N_3819,N_822);
and U7321 (N_7321,N_2468,N_435);
nand U7322 (N_7322,N_3687,N_4849);
or U7323 (N_7323,N_259,N_4397);
or U7324 (N_7324,N_4265,N_4670);
or U7325 (N_7325,N_2563,N_3829);
and U7326 (N_7326,N_4181,N_4320);
and U7327 (N_7327,N_2937,N_39);
xor U7328 (N_7328,N_1492,N_762);
or U7329 (N_7329,N_669,N_150);
or U7330 (N_7330,N_4765,N_3459);
nand U7331 (N_7331,N_21,N_651);
nor U7332 (N_7332,N_631,N_635);
and U7333 (N_7333,N_398,N_949);
xor U7334 (N_7334,N_2307,N_1169);
or U7335 (N_7335,N_4742,N_2000);
and U7336 (N_7336,N_1765,N_1700);
or U7337 (N_7337,N_4830,N_2188);
nand U7338 (N_7338,N_748,N_1506);
or U7339 (N_7339,N_2452,N_3932);
or U7340 (N_7340,N_3042,N_4339);
xnor U7341 (N_7341,N_4671,N_3698);
nor U7342 (N_7342,N_467,N_2178);
xnor U7343 (N_7343,N_2069,N_2180);
xnor U7344 (N_7344,N_1647,N_2372);
and U7345 (N_7345,N_1678,N_2511);
nand U7346 (N_7346,N_2578,N_2366);
or U7347 (N_7347,N_3671,N_1877);
and U7348 (N_7348,N_1594,N_97);
nand U7349 (N_7349,N_3651,N_3513);
nor U7350 (N_7350,N_353,N_1998);
or U7351 (N_7351,N_4160,N_3799);
or U7352 (N_7352,N_336,N_738);
nor U7353 (N_7353,N_1405,N_3127);
nand U7354 (N_7354,N_2507,N_1142);
or U7355 (N_7355,N_4926,N_607);
and U7356 (N_7356,N_3,N_3828);
nand U7357 (N_7357,N_1356,N_4579);
nor U7358 (N_7358,N_4225,N_3734);
nor U7359 (N_7359,N_3634,N_1992);
xnor U7360 (N_7360,N_196,N_111);
and U7361 (N_7361,N_3946,N_3696);
nor U7362 (N_7362,N_3473,N_3688);
nand U7363 (N_7363,N_2038,N_1053);
nor U7364 (N_7364,N_3316,N_3371);
and U7365 (N_7365,N_458,N_2958);
nand U7366 (N_7366,N_850,N_999);
and U7367 (N_7367,N_4419,N_3430);
xnor U7368 (N_7368,N_895,N_4406);
nand U7369 (N_7369,N_1853,N_4841);
and U7370 (N_7370,N_1945,N_1015);
xnor U7371 (N_7371,N_1742,N_4672);
nand U7372 (N_7372,N_1411,N_1976);
xnor U7373 (N_7373,N_3055,N_4911);
or U7374 (N_7374,N_1520,N_979);
and U7375 (N_7375,N_2170,N_647);
xor U7376 (N_7376,N_3054,N_2688);
and U7377 (N_7377,N_2361,N_2722);
nand U7378 (N_7378,N_708,N_2373);
or U7379 (N_7379,N_3455,N_3045);
or U7380 (N_7380,N_300,N_1672);
or U7381 (N_7381,N_4816,N_2238);
nand U7382 (N_7382,N_3758,N_2247);
nand U7383 (N_7383,N_2077,N_4887);
and U7384 (N_7384,N_4986,N_964);
and U7385 (N_7385,N_4602,N_2777);
and U7386 (N_7386,N_1418,N_4807);
or U7387 (N_7387,N_2628,N_1239);
or U7388 (N_7388,N_4970,N_1289);
xor U7389 (N_7389,N_1565,N_3680);
or U7390 (N_7390,N_1773,N_311);
and U7391 (N_7391,N_1063,N_61);
and U7392 (N_7392,N_775,N_3515);
nand U7393 (N_7393,N_2066,N_1137);
nor U7394 (N_7394,N_82,N_2610);
nand U7395 (N_7395,N_4994,N_1956);
and U7396 (N_7396,N_3282,N_291);
nor U7397 (N_7397,N_2899,N_136);
and U7398 (N_7398,N_3566,N_1719);
nand U7399 (N_7399,N_4637,N_1056);
nor U7400 (N_7400,N_3442,N_1725);
xnor U7401 (N_7401,N_2763,N_12);
or U7402 (N_7402,N_4203,N_2241);
xnor U7403 (N_7403,N_3662,N_4092);
or U7404 (N_7404,N_223,N_1882);
and U7405 (N_7405,N_2157,N_3416);
and U7406 (N_7406,N_1568,N_1648);
and U7407 (N_7407,N_3503,N_1495);
or U7408 (N_7408,N_27,N_3353);
nor U7409 (N_7409,N_3953,N_4761);
and U7410 (N_7410,N_68,N_2723);
or U7411 (N_7411,N_269,N_3244);
and U7412 (N_7412,N_1022,N_4686);
or U7413 (N_7413,N_2500,N_833);
nor U7414 (N_7414,N_1848,N_4934);
and U7415 (N_7415,N_1604,N_1906);
nand U7416 (N_7416,N_499,N_2865);
nor U7417 (N_7417,N_3243,N_684);
or U7418 (N_7418,N_542,N_4328);
xnor U7419 (N_7419,N_98,N_4925);
xor U7420 (N_7420,N_1455,N_2299);
nor U7421 (N_7421,N_1184,N_4180);
nor U7422 (N_7422,N_272,N_1862);
xnor U7423 (N_7423,N_2548,N_883);
nor U7424 (N_7424,N_3399,N_3293);
nor U7425 (N_7425,N_666,N_3924);
xor U7426 (N_7426,N_1350,N_2727);
or U7427 (N_7427,N_3286,N_3524);
xor U7428 (N_7428,N_3839,N_400);
nor U7429 (N_7429,N_2208,N_1262);
and U7430 (N_7430,N_4195,N_4175);
or U7431 (N_7431,N_3922,N_2963);
and U7432 (N_7432,N_3539,N_2586);
and U7433 (N_7433,N_1900,N_379);
nor U7434 (N_7434,N_603,N_4422);
or U7435 (N_7435,N_4612,N_459);
and U7436 (N_7436,N_1995,N_4941);
and U7437 (N_7437,N_4719,N_2387);
nor U7438 (N_7438,N_2422,N_1217);
xor U7439 (N_7439,N_665,N_1026);
nand U7440 (N_7440,N_707,N_4624);
or U7441 (N_7441,N_3542,N_2278);
xnor U7442 (N_7442,N_4161,N_1274);
nand U7443 (N_7443,N_2035,N_1358);
nand U7444 (N_7444,N_4545,N_2329);
or U7445 (N_7445,N_2016,N_4322);
or U7446 (N_7446,N_1438,N_1977);
nand U7447 (N_7447,N_1208,N_263);
nand U7448 (N_7448,N_726,N_1941);
and U7449 (N_7449,N_453,N_3129);
nor U7450 (N_7450,N_228,N_879);
or U7451 (N_7451,N_2818,N_2335);
nand U7452 (N_7452,N_3944,N_312);
and U7453 (N_7453,N_1597,N_2362);
or U7454 (N_7454,N_4006,N_189);
or U7455 (N_7455,N_3393,N_3193);
and U7456 (N_7456,N_245,N_4460);
nand U7457 (N_7457,N_2866,N_2339);
nor U7458 (N_7458,N_4448,N_1188);
nor U7459 (N_7459,N_3960,N_241);
nor U7460 (N_7460,N_1603,N_923);
xnor U7461 (N_7461,N_3936,N_2130);
nor U7462 (N_7462,N_3817,N_4505);
nor U7463 (N_7463,N_3273,N_3182);
nand U7464 (N_7464,N_492,N_1368);
nor U7465 (N_7465,N_817,N_2761);
and U7466 (N_7466,N_4286,N_2271);
or U7467 (N_7467,N_3002,N_461);
nor U7468 (N_7468,N_2303,N_1054);
and U7469 (N_7469,N_3832,N_3749);
nand U7470 (N_7470,N_1835,N_788);
xor U7471 (N_7471,N_4519,N_908);
nor U7472 (N_7472,N_294,N_4516);
or U7473 (N_7473,N_4402,N_1254);
nand U7474 (N_7474,N_2833,N_1415);
and U7475 (N_7475,N_491,N_3693);
nand U7476 (N_7476,N_384,N_4469);
xor U7477 (N_7477,N_567,N_4242);
nand U7478 (N_7478,N_2076,N_2406);
and U7479 (N_7479,N_3392,N_2946);
nor U7480 (N_7480,N_1027,N_672);
or U7481 (N_7481,N_1104,N_3773);
nand U7482 (N_7482,N_1421,N_1957);
nor U7483 (N_7483,N_2886,N_3231);
nor U7484 (N_7484,N_3462,N_4600);
xnor U7485 (N_7485,N_1829,N_2265);
and U7486 (N_7486,N_140,N_2981);
or U7487 (N_7487,N_4398,N_3287);
nand U7488 (N_7488,N_2961,N_3875);
and U7489 (N_7489,N_3104,N_2594);
or U7490 (N_7490,N_876,N_3175);
nor U7491 (N_7491,N_2508,N_2772);
nand U7492 (N_7492,N_4693,N_1662);
xnor U7493 (N_7493,N_3254,N_1914);
nor U7494 (N_7494,N_108,N_722);
xnor U7495 (N_7495,N_1106,N_3760);
or U7496 (N_7496,N_187,N_201);
nand U7497 (N_7497,N_3650,N_4068);
xnor U7498 (N_7498,N_3217,N_3642);
nor U7499 (N_7499,N_2483,N_445);
or U7500 (N_7500,N_3023,N_2667);
nand U7501 (N_7501,N_1187,N_562);
xor U7502 (N_7502,N_2471,N_4901);
or U7503 (N_7503,N_2326,N_3528);
nor U7504 (N_7504,N_2104,N_649);
nor U7505 (N_7505,N_4145,N_2191);
xnor U7506 (N_7506,N_345,N_4601);
or U7507 (N_7507,N_1257,N_1637);
xor U7508 (N_7508,N_3062,N_3128);
nor U7509 (N_7509,N_2951,N_336);
nor U7510 (N_7510,N_3336,N_1213);
nand U7511 (N_7511,N_232,N_3378);
or U7512 (N_7512,N_3670,N_68);
nand U7513 (N_7513,N_3896,N_1913);
nand U7514 (N_7514,N_2695,N_2058);
and U7515 (N_7515,N_1006,N_827);
xor U7516 (N_7516,N_2122,N_4412);
nor U7517 (N_7517,N_2506,N_4464);
xor U7518 (N_7518,N_1360,N_1713);
xor U7519 (N_7519,N_1940,N_2241);
and U7520 (N_7520,N_2096,N_1322);
or U7521 (N_7521,N_4251,N_591);
nand U7522 (N_7522,N_275,N_355);
or U7523 (N_7523,N_2037,N_3359);
or U7524 (N_7524,N_3667,N_4412);
nand U7525 (N_7525,N_1919,N_1443);
nand U7526 (N_7526,N_4608,N_2382);
or U7527 (N_7527,N_4494,N_662);
or U7528 (N_7528,N_4240,N_3964);
nor U7529 (N_7529,N_4303,N_1255);
or U7530 (N_7530,N_4403,N_506);
or U7531 (N_7531,N_1404,N_2702);
and U7532 (N_7532,N_1379,N_2042);
nand U7533 (N_7533,N_2555,N_3958);
xnor U7534 (N_7534,N_4469,N_294);
or U7535 (N_7535,N_3967,N_294);
nor U7536 (N_7536,N_2582,N_3209);
nor U7537 (N_7537,N_3931,N_4026);
nor U7538 (N_7538,N_4058,N_3506);
or U7539 (N_7539,N_1007,N_4577);
and U7540 (N_7540,N_2169,N_2465);
nor U7541 (N_7541,N_3002,N_1943);
xor U7542 (N_7542,N_4384,N_2797);
nand U7543 (N_7543,N_3637,N_2247);
nand U7544 (N_7544,N_2111,N_4240);
and U7545 (N_7545,N_233,N_2723);
and U7546 (N_7546,N_1569,N_2252);
nand U7547 (N_7547,N_4980,N_444);
or U7548 (N_7548,N_3332,N_4604);
xnor U7549 (N_7549,N_4339,N_1327);
xor U7550 (N_7550,N_4342,N_572);
xnor U7551 (N_7551,N_3016,N_2029);
or U7552 (N_7552,N_556,N_72);
nor U7553 (N_7553,N_1251,N_3842);
nand U7554 (N_7554,N_3601,N_3321);
and U7555 (N_7555,N_4800,N_3391);
nand U7556 (N_7556,N_90,N_4231);
nand U7557 (N_7557,N_887,N_2166);
nor U7558 (N_7558,N_2560,N_4099);
or U7559 (N_7559,N_3279,N_2365);
nor U7560 (N_7560,N_293,N_1731);
xnor U7561 (N_7561,N_3300,N_3957);
and U7562 (N_7562,N_2444,N_1171);
xor U7563 (N_7563,N_4626,N_2454);
and U7564 (N_7564,N_2864,N_3395);
or U7565 (N_7565,N_1422,N_2056);
nand U7566 (N_7566,N_3974,N_3580);
nor U7567 (N_7567,N_976,N_4819);
nor U7568 (N_7568,N_1523,N_1299);
and U7569 (N_7569,N_774,N_4115);
nand U7570 (N_7570,N_4056,N_485);
nor U7571 (N_7571,N_3948,N_3096);
xor U7572 (N_7572,N_3582,N_4208);
xor U7573 (N_7573,N_3771,N_4611);
xnor U7574 (N_7574,N_2890,N_2625);
and U7575 (N_7575,N_4927,N_4265);
nand U7576 (N_7576,N_2905,N_4676);
and U7577 (N_7577,N_4049,N_908);
or U7578 (N_7578,N_1750,N_801);
xor U7579 (N_7579,N_1361,N_3229);
xnor U7580 (N_7580,N_4818,N_354);
nand U7581 (N_7581,N_4128,N_835);
or U7582 (N_7582,N_4780,N_4277);
nand U7583 (N_7583,N_396,N_15);
and U7584 (N_7584,N_2936,N_2979);
and U7585 (N_7585,N_3283,N_2636);
nand U7586 (N_7586,N_1249,N_3317);
or U7587 (N_7587,N_2948,N_2079);
xor U7588 (N_7588,N_2893,N_1757);
or U7589 (N_7589,N_3453,N_105);
or U7590 (N_7590,N_4877,N_441);
xnor U7591 (N_7591,N_69,N_1555);
nor U7592 (N_7592,N_3575,N_2335);
nor U7593 (N_7593,N_3226,N_220);
xnor U7594 (N_7594,N_4894,N_1532);
and U7595 (N_7595,N_3413,N_3879);
and U7596 (N_7596,N_3962,N_3125);
nand U7597 (N_7597,N_3832,N_4000);
and U7598 (N_7598,N_4455,N_2959);
and U7599 (N_7599,N_274,N_2873);
xnor U7600 (N_7600,N_3915,N_1036);
nand U7601 (N_7601,N_1468,N_2953);
xor U7602 (N_7602,N_1717,N_102);
or U7603 (N_7603,N_218,N_2820);
nand U7604 (N_7604,N_1136,N_4466);
and U7605 (N_7605,N_4913,N_4374);
or U7606 (N_7606,N_1494,N_314);
nand U7607 (N_7607,N_1869,N_1537);
nor U7608 (N_7608,N_1274,N_2672);
nand U7609 (N_7609,N_650,N_2425);
nor U7610 (N_7610,N_2830,N_3634);
and U7611 (N_7611,N_2335,N_1856);
xnor U7612 (N_7612,N_1324,N_4339);
nand U7613 (N_7613,N_725,N_1823);
nor U7614 (N_7614,N_2356,N_3291);
nand U7615 (N_7615,N_1782,N_85);
and U7616 (N_7616,N_2192,N_2762);
and U7617 (N_7617,N_701,N_922);
nand U7618 (N_7618,N_573,N_3008);
nor U7619 (N_7619,N_1484,N_1723);
nor U7620 (N_7620,N_2487,N_2231);
and U7621 (N_7621,N_1999,N_2547);
or U7622 (N_7622,N_2669,N_2418);
nor U7623 (N_7623,N_1403,N_4939);
xnor U7624 (N_7624,N_4974,N_1908);
nand U7625 (N_7625,N_686,N_4113);
and U7626 (N_7626,N_1673,N_1372);
and U7627 (N_7627,N_1671,N_364);
nand U7628 (N_7628,N_271,N_2755);
nor U7629 (N_7629,N_3167,N_1619);
xnor U7630 (N_7630,N_3872,N_727);
and U7631 (N_7631,N_3193,N_2899);
and U7632 (N_7632,N_3015,N_417);
xor U7633 (N_7633,N_3203,N_703);
or U7634 (N_7634,N_4819,N_4285);
xnor U7635 (N_7635,N_2850,N_4282);
nand U7636 (N_7636,N_4884,N_4505);
nand U7637 (N_7637,N_2620,N_4759);
nor U7638 (N_7638,N_780,N_4250);
xor U7639 (N_7639,N_127,N_2921);
or U7640 (N_7640,N_1813,N_2848);
and U7641 (N_7641,N_1419,N_2232);
or U7642 (N_7642,N_1576,N_948);
xnor U7643 (N_7643,N_3454,N_292);
nor U7644 (N_7644,N_481,N_3403);
and U7645 (N_7645,N_2272,N_927);
and U7646 (N_7646,N_38,N_1841);
xor U7647 (N_7647,N_469,N_67);
or U7648 (N_7648,N_1414,N_4996);
xnor U7649 (N_7649,N_3174,N_987);
nand U7650 (N_7650,N_2839,N_780);
nor U7651 (N_7651,N_308,N_1806);
xnor U7652 (N_7652,N_879,N_2066);
or U7653 (N_7653,N_2249,N_2375);
nor U7654 (N_7654,N_1268,N_3771);
nor U7655 (N_7655,N_248,N_975);
nor U7656 (N_7656,N_703,N_1404);
xor U7657 (N_7657,N_3350,N_4158);
nand U7658 (N_7658,N_2510,N_227);
xor U7659 (N_7659,N_4638,N_923);
nand U7660 (N_7660,N_1882,N_4190);
or U7661 (N_7661,N_4274,N_3270);
or U7662 (N_7662,N_2212,N_2196);
or U7663 (N_7663,N_1145,N_1193);
xnor U7664 (N_7664,N_1832,N_918);
or U7665 (N_7665,N_4535,N_4883);
nor U7666 (N_7666,N_4842,N_1099);
nor U7667 (N_7667,N_253,N_3210);
nor U7668 (N_7668,N_1949,N_4679);
nor U7669 (N_7669,N_2701,N_4158);
nor U7670 (N_7670,N_1029,N_804);
xnor U7671 (N_7671,N_1729,N_1627);
nor U7672 (N_7672,N_2518,N_1483);
or U7673 (N_7673,N_632,N_2676);
xor U7674 (N_7674,N_820,N_1704);
or U7675 (N_7675,N_2761,N_3262);
xnor U7676 (N_7676,N_1762,N_1782);
nand U7677 (N_7677,N_2545,N_1585);
nor U7678 (N_7678,N_4109,N_3236);
or U7679 (N_7679,N_4932,N_358);
or U7680 (N_7680,N_964,N_2955);
xnor U7681 (N_7681,N_1783,N_3197);
or U7682 (N_7682,N_3228,N_339);
nand U7683 (N_7683,N_2548,N_979);
and U7684 (N_7684,N_2138,N_2732);
nand U7685 (N_7685,N_389,N_1572);
nand U7686 (N_7686,N_4424,N_3640);
nand U7687 (N_7687,N_2189,N_495);
and U7688 (N_7688,N_3013,N_4896);
and U7689 (N_7689,N_2146,N_680);
or U7690 (N_7690,N_3409,N_275);
nor U7691 (N_7691,N_1683,N_3613);
and U7692 (N_7692,N_3979,N_4488);
xnor U7693 (N_7693,N_4674,N_4185);
xnor U7694 (N_7694,N_1301,N_279);
and U7695 (N_7695,N_4651,N_322);
nand U7696 (N_7696,N_3659,N_1525);
or U7697 (N_7697,N_3630,N_2190);
or U7698 (N_7698,N_648,N_327);
nor U7699 (N_7699,N_859,N_4931);
or U7700 (N_7700,N_4484,N_1176);
nand U7701 (N_7701,N_4256,N_4397);
nand U7702 (N_7702,N_651,N_3036);
nor U7703 (N_7703,N_1117,N_2250);
and U7704 (N_7704,N_322,N_1972);
and U7705 (N_7705,N_3068,N_1959);
nand U7706 (N_7706,N_4219,N_1900);
xor U7707 (N_7707,N_1232,N_3732);
and U7708 (N_7708,N_1602,N_3695);
nor U7709 (N_7709,N_1116,N_2315);
or U7710 (N_7710,N_612,N_347);
nor U7711 (N_7711,N_1081,N_3272);
xnor U7712 (N_7712,N_2666,N_2490);
xor U7713 (N_7713,N_2016,N_380);
and U7714 (N_7714,N_1558,N_1500);
nor U7715 (N_7715,N_4637,N_1138);
and U7716 (N_7716,N_3037,N_2493);
xor U7717 (N_7717,N_1079,N_2607);
xnor U7718 (N_7718,N_3986,N_3090);
nor U7719 (N_7719,N_3842,N_4791);
or U7720 (N_7720,N_4744,N_2723);
nor U7721 (N_7721,N_591,N_1068);
and U7722 (N_7722,N_914,N_974);
nand U7723 (N_7723,N_4192,N_4964);
nor U7724 (N_7724,N_2296,N_3976);
xnor U7725 (N_7725,N_3302,N_760);
xnor U7726 (N_7726,N_1005,N_4094);
and U7727 (N_7727,N_866,N_4919);
xor U7728 (N_7728,N_3263,N_887);
and U7729 (N_7729,N_2313,N_1288);
nand U7730 (N_7730,N_1124,N_3999);
and U7731 (N_7731,N_415,N_2152);
nand U7732 (N_7732,N_4243,N_2596);
xor U7733 (N_7733,N_4973,N_2764);
nand U7734 (N_7734,N_2158,N_3465);
and U7735 (N_7735,N_2192,N_1713);
or U7736 (N_7736,N_1543,N_2654);
nor U7737 (N_7737,N_3602,N_85);
or U7738 (N_7738,N_1865,N_2061);
and U7739 (N_7739,N_4082,N_3977);
nand U7740 (N_7740,N_327,N_375);
nor U7741 (N_7741,N_3077,N_4701);
or U7742 (N_7742,N_2271,N_635);
nand U7743 (N_7743,N_1864,N_2319);
nand U7744 (N_7744,N_818,N_1785);
and U7745 (N_7745,N_1617,N_3735);
xor U7746 (N_7746,N_1947,N_1250);
or U7747 (N_7747,N_4090,N_3148);
or U7748 (N_7748,N_438,N_2105);
or U7749 (N_7749,N_3047,N_31);
xnor U7750 (N_7750,N_1520,N_318);
or U7751 (N_7751,N_2799,N_3034);
and U7752 (N_7752,N_1752,N_1490);
or U7753 (N_7753,N_323,N_406);
or U7754 (N_7754,N_68,N_305);
nand U7755 (N_7755,N_452,N_2427);
nor U7756 (N_7756,N_2290,N_3689);
xor U7757 (N_7757,N_1542,N_1664);
nand U7758 (N_7758,N_1370,N_996);
nand U7759 (N_7759,N_528,N_1773);
nand U7760 (N_7760,N_1123,N_387);
nor U7761 (N_7761,N_3712,N_1834);
nand U7762 (N_7762,N_2023,N_2647);
or U7763 (N_7763,N_4020,N_4175);
and U7764 (N_7764,N_3205,N_68);
or U7765 (N_7765,N_4626,N_4723);
nand U7766 (N_7766,N_907,N_2596);
or U7767 (N_7767,N_1546,N_1963);
and U7768 (N_7768,N_960,N_1798);
and U7769 (N_7769,N_833,N_841);
nor U7770 (N_7770,N_3255,N_3748);
and U7771 (N_7771,N_3631,N_2936);
or U7772 (N_7772,N_3008,N_3727);
xor U7773 (N_7773,N_3984,N_2601);
nand U7774 (N_7774,N_1458,N_1865);
or U7775 (N_7775,N_4455,N_2962);
and U7776 (N_7776,N_543,N_1681);
or U7777 (N_7777,N_1302,N_879);
nand U7778 (N_7778,N_531,N_4072);
nor U7779 (N_7779,N_4730,N_1666);
or U7780 (N_7780,N_241,N_35);
and U7781 (N_7781,N_4720,N_286);
or U7782 (N_7782,N_3903,N_16);
and U7783 (N_7783,N_4205,N_1984);
and U7784 (N_7784,N_1713,N_3433);
and U7785 (N_7785,N_4236,N_959);
or U7786 (N_7786,N_2423,N_4157);
and U7787 (N_7787,N_4266,N_3503);
xnor U7788 (N_7788,N_3436,N_1452);
nand U7789 (N_7789,N_2462,N_4218);
or U7790 (N_7790,N_716,N_2505);
xnor U7791 (N_7791,N_3785,N_3119);
and U7792 (N_7792,N_3433,N_953);
xnor U7793 (N_7793,N_1963,N_1067);
and U7794 (N_7794,N_4208,N_4332);
nand U7795 (N_7795,N_162,N_3742);
or U7796 (N_7796,N_3174,N_4434);
or U7797 (N_7797,N_3925,N_732);
nand U7798 (N_7798,N_3660,N_3362);
nand U7799 (N_7799,N_1062,N_1146);
xor U7800 (N_7800,N_4028,N_928);
or U7801 (N_7801,N_4270,N_4972);
or U7802 (N_7802,N_4400,N_1755);
and U7803 (N_7803,N_3518,N_3908);
xor U7804 (N_7804,N_3852,N_382);
xnor U7805 (N_7805,N_4851,N_1689);
xnor U7806 (N_7806,N_4652,N_4956);
xor U7807 (N_7807,N_400,N_2316);
xor U7808 (N_7808,N_3369,N_4169);
or U7809 (N_7809,N_3805,N_3240);
and U7810 (N_7810,N_1290,N_3715);
xnor U7811 (N_7811,N_4426,N_4286);
nor U7812 (N_7812,N_4857,N_190);
or U7813 (N_7813,N_2645,N_4712);
xnor U7814 (N_7814,N_4231,N_4057);
nor U7815 (N_7815,N_3625,N_2062);
xnor U7816 (N_7816,N_3783,N_4940);
or U7817 (N_7817,N_3336,N_2994);
nor U7818 (N_7818,N_4458,N_2594);
nand U7819 (N_7819,N_824,N_1219);
nor U7820 (N_7820,N_1101,N_3619);
and U7821 (N_7821,N_1839,N_2376);
or U7822 (N_7822,N_894,N_399);
nor U7823 (N_7823,N_311,N_2805);
nor U7824 (N_7824,N_3140,N_1594);
nand U7825 (N_7825,N_2597,N_556);
nand U7826 (N_7826,N_881,N_1923);
and U7827 (N_7827,N_2733,N_4994);
nor U7828 (N_7828,N_1123,N_270);
nor U7829 (N_7829,N_583,N_4676);
or U7830 (N_7830,N_338,N_3518);
or U7831 (N_7831,N_3425,N_4776);
or U7832 (N_7832,N_4323,N_1276);
or U7833 (N_7833,N_4746,N_1151);
or U7834 (N_7834,N_160,N_2644);
and U7835 (N_7835,N_548,N_2371);
xor U7836 (N_7836,N_1516,N_2800);
nor U7837 (N_7837,N_795,N_263);
or U7838 (N_7838,N_4249,N_3916);
xor U7839 (N_7839,N_3648,N_4617);
and U7840 (N_7840,N_4984,N_1405);
nor U7841 (N_7841,N_3026,N_2423);
nand U7842 (N_7842,N_2547,N_756);
nor U7843 (N_7843,N_4398,N_297);
nand U7844 (N_7844,N_1025,N_2874);
xnor U7845 (N_7845,N_4508,N_961);
and U7846 (N_7846,N_3313,N_3198);
nand U7847 (N_7847,N_3258,N_1258);
or U7848 (N_7848,N_2437,N_2812);
nor U7849 (N_7849,N_330,N_4575);
nand U7850 (N_7850,N_2090,N_1639);
nand U7851 (N_7851,N_3513,N_189);
and U7852 (N_7852,N_1602,N_1803);
xor U7853 (N_7853,N_1392,N_963);
nand U7854 (N_7854,N_1310,N_368);
xor U7855 (N_7855,N_2522,N_4700);
or U7856 (N_7856,N_2853,N_4564);
or U7857 (N_7857,N_2169,N_3677);
nor U7858 (N_7858,N_2060,N_3962);
or U7859 (N_7859,N_1092,N_2024);
nand U7860 (N_7860,N_3394,N_3607);
nand U7861 (N_7861,N_2525,N_824);
and U7862 (N_7862,N_1806,N_3997);
and U7863 (N_7863,N_4238,N_3579);
nand U7864 (N_7864,N_222,N_1810);
or U7865 (N_7865,N_799,N_2521);
xor U7866 (N_7866,N_151,N_4904);
nand U7867 (N_7867,N_4019,N_947);
xnor U7868 (N_7868,N_3323,N_2897);
nor U7869 (N_7869,N_1714,N_873);
nor U7870 (N_7870,N_1226,N_4191);
nor U7871 (N_7871,N_792,N_3730);
or U7872 (N_7872,N_914,N_4544);
or U7873 (N_7873,N_1582,N_277);
nand U7874 (N_7874,N_4606,N_1691);
xnor U7875 (N_7875,N_1804,N_2761);
or U7876 (N_7876,N_2175,N_243);
and U7877 (N_7877,N_350,N_1792);
nand U7878 (N_7878,N_4280,N_236);
nand U7879 (N_7879,N_2701,N_1650);
nor U7880 (N_7880,N_2155,N_2929);
nand U7881 (N_7881,N_74,N_4789);
nor U7882 (N_7882,N_78,N_3785);
xnor U7883 (N_7883,N_3327,N_1608);
and U7884 (N_7884,N_1160,N_168);
and U7885 (N_7885,N_3208,N_1610);
nor U7886 (N_7886,N_2348,N_1496);
and U7887 (N_7887,N_911,N_1180);
nor U7888 (N_7888,N_4171,N_2651);
nand U7889 (N_7889,N_3202,N_858);
xnor U7890 (N_7890,N_1977,N_1730);
nand U7891 (N_7891,N_1444,N_1622);
or U7892 (N_7892,N_4708,N_1638);
and U7893 (N_7893,N_977,N_37);
nor U7894 (N_7894,N_2364,N_857);
nand U7895 (N_7895,N_921,N_1585);
and U7896 (N_7896,N_1623,N_2378);
nor U7897 (N_7897,N_1718,N_2634);
xor U7898 (N_7898,N_266,N_1853);
and U7899 (N_7899,N_340,N_2313);
or U7900 (N_7900,N_2254,N_2926);
xnor U7901 (N_7901,N_4997,N_287);
nor U7902 (N_7902,N_2605,N_4161);
xor U7903 (N_7903,N_3568,N_3625);
nand U7904 (N_7904,N_1447,N_4074);
nor U7905 (N_7905,N_2878,N_3463);
or U7906 (N_7906,N_2716,N_4413);
xor U7907 (N_7907,N_2009,N_617);
or U7908 (N_7908,N_1769,N_1706);
nor U7909 (N_7909,N_3589,N_3106);
or U7910 (N_7910,N_3962,N_3665);
nand U7911 (N_7911,N_4812,N_2768);
xnor U7912 (N_7912,N_1031,N_4380);
and U7913 (N_7913,N_1406,N_2703);
nand U7914 (N_7914,N_161,N_4649);
nor U7915 (N_7915,N_4279,N_664);
nor U7916 (N_7916,N_3496,N_1891);
and U7917 (N_7917,N_4104,N_3598);
and U7918 (N_7918,N_2629,N_1480);
xnor U7919 (N_7919,N_1613,N_4483);
or U7920 (N_7920,N_3334,N_2279);
and U7921 (N_7921,N_3284,N_2267);
and U7922 (N_7922,N_2879,N_289);
or U7923 (N_7923,N_3452,N_2844);
nor U7924 (N_7924,N_1186,N_727);
nand U7925 (N_7925,N_2372,N_3143);
and U7926 (N_7926,N_2052,N_1815);
and U7927 (N_7927,N_4204,N_4504);
xor U7928 (N_7928,N_3864,N_737);
xor U7929 (N_7929,N_2335,N_2921);
and U7930 (N_7930,N_919,N_4191);
and U7931 (N_7931,N_1490,N_1460);
and U7932 (N_7932,N_2782,N_2189);
or U7933 (N_7933,N_2940,N_634);
nor U7934 (N_7934,N_1580,N_4449);
xor U7935 (N_7935,N_1270,N_1394);
nand U7936 (N_7936,N_4567,N_2616);
and U7937 (N_7937,N_4220,N_1928);
and U7938 (N_7938,N_4138,N_359);
nand U7939 (N_7939,N_660,N_3266);
nand U7940 (N_7940,N_4726,N_535);
and U7941 (N_7941,N_239,N_3819);
or U7942 (N_7942,N_2015,N_3139);
nor U7943 (N_7943,N_2136,N_4290);
xnor U7944 (N_7944,N_1635,N_177);
xnor U7945 (N_7945,N_2708,N_3408);
nor U7946 (N_7946,N_4843,N_716);
nor U7947 (N_7947,N_2512,N_1513);
or U7948 (N_7948,N_4420,N_2684);
or U7949 (N_7949,N_467,N_4921);
and U7950 (N_7950,N_505,N_1704);
and U7951 (N_7951,N_4262,N_3164);
or U7952 (N_7952,N_3598,N_886);
xnor U7953 (N_7953,N_2385,N_880);
or U7954 (N_7954,N_1289,N_2799);
and U7955 (N_7955,N_2898,N_1107);
nor U7956 (N_7956,N_4999,N_2925);
nand U7957 (N_7957,N_4098,N_4666);
nand U7958 (N_7958,N_2332,N_1494);
or U7959 (N_7959,N_2921,N_2538);
nor U7960 (N_7960,N_4453,N_1255);
and U7961 (N_7961,N_164,N_1862);
nor U7962 (N_7962,N_3256,N_3000);
nor U7963 (N_7963,N_2592,N_2779);
nand U7964 (N_7964,N_3387,N_3768);
and U7965 (N_7965,N_4101,N_3994);
nor U7966 (N_7966,N_3283,N_1584);
xnor U7967 (N_7967,N_2978,N_854);
nand U7968 (N_7968,N_2943,N_4002);
nand U7969 (N_7969,N_3276,N_4758);
nor U7970 (N_7970,N_4788,N_4602);
nor U7971 (N_7971,N_4163,N_3354);
nand U7972 (N_7972,N_232,N_4496);
nor U7973 (N_7973,N_3650,N_3031);
or U7974 (N_7974,N_3677,N_2736);
or U7975 (N_7975,N_2803,N_1411);
nor U7976 (N_7976,N_3279,N_2185);
and U7977 (N_7977,N_889,N_2963);
and U7978 (N_7978,N_3720,N_1023);
or U7979 (N_7979,N_4935,N_1005);
or U7980 (N_7980,N_956,N_48);
xnor U7981 (N_7981,N_708,N_778);
and U7982 (N_7982,N_3884,N_4721);
nor U7983 (N_7983,N_2940,N_3320);
and U7984 (N_7984,N_724,N_2252);
nor U7985 (N_7985,N_1207,N_1828);
nand U7986 (N_7986,N_855,N_1764);
or U7987 (N_7987,N_2090,N_2179);
nor U7988 (N_7988,N_1412,N_947);
nand U7989 (N_7989,N_990,N_3913);
nor U7990 (N_7990,N_1352,N_3498);
or U7991 (N_7991,N_1433,N_1232);
or U7992 (N_7992,N_1227,N_3523);
and U7993 (N_7993,N_3,N_1395);
and U7994 (N_7994,N_4333,N_1513);
xnor U7995 (N_7995,N_4359,N_842);
and U7996 (N_7996,N_3261,N_3045);
and U7997 (N_7997,N_3042,N_688);
or U7998 (N_7998,N_39,N_1414);
and U7999 (N_7999,N_661,N_1014);
xor U8000 (N_8000,N_1663,N_3024);
and U8001 (N_8001,N_689,N_4672);
xnor U8002 (N_8002,N_3587,N_4234);
nor U8003 (N_8003,N_2032,N_393);
and U8004 (N_8004,N_446,N_4139);
xor U8005 (N_8005,N_496,N_2879);
xor U8006 (N_8006,N_960,N_3030);
nand U8007 (N_8007,N_3353,N_4548);
nor U8008 (N_8008,N_3023,N_2721);
nand U8009 (N_8009,N_4330,N_2880);
nor U8010 (N_8010,N_915,N_1994);
and U8011 (N_8011,N_4776,N_272);
xnor U8012 (N_8012,N_4334,N_156);
or U8013 (N_8013,N_4605,N_1814);
xnor U8014 (N_8014,N_3925,N_1977);
nand U8015 (N_8015,N_1150,N_2166);
xor U8016 (N_8016,N_4368,N_1901);
and U8017 (N_8017,N_3175,N_3909);
and U8018 (N_8018,N_4239,N_838);
nor U8019 (N_8019,N_1867,N_3292);
or U8020 (N_8020,N_3887,N_2642);
xor U8021 (N_8021,N_698,N_526);
nand U8022 (N_8022,N_4780,N_494);
nor U8023 (N_8023,N_4217,N_3909);
nand U8024 (N_8024,N_491,N_1661);
nor U8025 (N_8025,N_2189,N_4422);
nor U8026 (N_8026,N_4028,N_4985);
xnor U8027 (N_8027,N_3602,N_2065);
nor U8028 (N_8028,N_2428,N_3745);
or U8029 (N_8029,N_4842,N_4182);
nor U8030 (N_8030,N_4306,N_1633);
xnor U8031 (N_8031,N_3664,N_680);
nor U8032 (N_8032,N_1271,N_3738);
nor U8033 (N_8033,N_1884,N_2775);
or U8034 (N_8034,N_1362,N_1366);
nand U8035 (N_8035,N_1562,N_3442);
nor U8036 (N_8036,N_3937,N_2708);
xnor U8037 (N_8037,N_1101,N_3527);
nor U8038 (N_8038,N_1851,N_1475);
or U8039 (N_8039,N_4332,N_471);
xnor U8040 (N_8040,N_1510,N_1438);
nor U8041 (N_8041,N_3540,N_1253);
and U8042 (N_8042,N_3933,N_1179);
nand U8043 (N_8043,N_4155,N_4829);
xor U8044 (N_8044,N_3792,N_2277);
nand U8045 (N_8045,N_496,N_3832);
xnor U8046 (N_8046,N_917,N_3106);
nand U8047 (N_8047,N_821,N_4801);
nor U8048 (N_8048,N_2278,N_4828);
nand U8049 (N_8049,N_914,N_1129);
or U8050 (N_8050,N_2231,N_3503);
nand U8051 (N_8051,N_1978,N_551);
and U8052 (N_8052,N_2448,N_4036);
xnor U8053 (N_8053,N_242,N_2932);
xor U8054 (N_8054,N_2932,N_1004);
or U8055 (N_8055,N_4458,N_2637);
nor U8056 (N_8056,N_331,N_581);
and U8057 (N_8057,N_4220,N_1207);
or U8058 (N_8058,N_1227,N_1974);
xor U8059 (N_8059,N_4240,N_2613);
nand U8060 (N_8060,N_815,N_467);
or U8061 (N_8061,N_424,N_4174);
nand U8062 (N_8062,N_2162,N_1134);
or U8063 (N_8063,N_824,N_4438);
nor U8064 (N_8064,N_2222,N_785);
or U8065 (N_8065,N_4239,N_4848);
or U8066 (N_8066,N_2021,N_1783);
xor U8067 (N_8067,N_2562,N_3893);
nor U8068 (N_8068,N_2685,N_61);
nor U8069 (N_8069,N_4160,N_650);
xor U8070 (N_8070,N_4520,N_198);
or U8071 (N_8071,N_3772,N_11);
nand U8072 (N_8072,N_2758,N_1091);
xor U8073 (N_8073,N_4253,N_334);
nor U8074 (N_8074,N_74,N_888);
xnor U8075 (N_8075,N_2598,N_870);
xnor U8076 (N_8076,N_1514,N_4700);
nand U8077 (N_8077,N_520,N_2361);
nand U8078 (N_8078,N_1196,N_378);
or U8079 (N_8079,N_3779,N_1430);
or U8080 (N_8080,N_236,N_925);
nor U8081 (N_8081,N_1816,N_3007);
xor U8082 (N_8082,N_3811,N_480);
and U8083 (N_8083,N_4283,N_2164);
or U8084 (N_8084,N_1725,N_1675);
nor U8085 (N_8085,N_3837,N_4711);
or U8086 (N_8086,N_205,N_3043);
xnor U8087 (N_8087,N_64,N_2093);
nand U8088 (N_8088,N_2537,N_886);
xor U8089 (N_8089,N_4841,N_730);
or U8090 (N_8090,N_4444,N_1655);
and U8091 (N_8091,N_3805,N_1270);
nand U8092 (N_8092,N_4303,N_4883);
nand U8093 (N_8093,N_4171,N_150);
nand U8094 (N_8094,N_3207,N_4763);
and U8095 (N_8095,N_2819,N_826);
or U8096 (N_8096,N_301,N_2651);
and U8097 (N_8097,N_170,N_1606);
or U8098 (N_8098,N_2521,N_1114);
or U8099 (N_8099,N_902,N_983);
or U8100 (N_8100,N_3218,N_2472);
or U8101 (N_8101,N_4714,N_1568);
nor U8102 (N_8102,N_2418,N_1047);
or U8103 (N_8103,N_3561,N_827);
and U8104 (N_8104,N_3568,N_3523);
nand U8105 (N_8105,N_4748,N_3294);
xor U8106 (N_8106,N_3617,N_2417);
and U8107 (N_8107,N_1331,N_558);
and U8108 (N_8108,N_2439,N_4812);
or U8109 (N_8109,N_4687,N_1673);
and U8110 (N_8110,N_2638,N_369);
xnor U8111 (N_8111,N_1780,N_3351);
and U8112 (N_8112,N_456,N_1881);
nand U8113 (N_8113,N_2444,N_3425);
and U8114 (N_8114,N_2563,N_1525);
nor U8115 (N_8115,N_2839,N_1313);
nand U8116 (N_8116,N_2437,N_3589);
xor U8117 (N_8117,N_1013,N_3509);
or U8118 (N_8118,N_4111,N_2547);
nand U8119 (N_8119,N_1022,N_3508);
or U8120 (N_8120,N_1621,N_2859);
or U8121 (N_8121,N_3538,N_1142);
or U8122 (N_8122,N_3367,N_2613);
nor U8123 (N_8123,N_1072,N_3836);
xor U8124 (N_8124,N_2071,N_481);
and U8125 (N_8125,N_1160,N_1636);
nor U8126 (N_8126,N_4193,N_2050);
and U8127 (N_8127,N_1568,N_4174);
or U8128 (N_8128,N_730,N_600);
xor U8129 (N_8129,N_1379,N_1185);
nor U8130 (N_8130,N_671,N_4923);
nor U8131 (N_8131,N_2443,N_1274);
nor U8132 (N_8132,N_721,N_2403);
or U8133 (N_8133,N_4509,N_1130);
or U8134 (N_8134,N_958,N_56);
nor U8135 (N_8135,N_2397,N_4415);
nor U8136 (N_8136,N_4329,N_4207);
or U8137 (N_8137,N_3376,N_3239);
or U8138 (N_8138,N_455,N_228);
xor U8139 (N_8139,N_4006,N_3275);
nand U8140 (N_8140,N_4999,N_88);
xnor U8141 (N_8141,N_4931,N_902);
xnor U8142 (N_8142,N_864,N_4396);
nand U8143 (N_8143,N_3667,N_237);
nor U8144 (N_8144,N_393,N_1802);
nand U8145 (N_8145,N_3152,N_2376);
nor U8146 (N_8146,N_298,N_70);
and U8147 (N_8147,N_972,N_1988);
nor U8148 (N_8148,N_203,N_2235);
nand U8149 (N_8149,N_4863,N_3363);
nand U8150 (N_8150,N_1989,N_1992);
and U8151 (N_8151,N_457,N_4245);
xnor U8152 (N_8152,N_404,N_54);
nor U8153 (N_8153,N_1667,N_4342);
xnor U8154 (N_8154,N_3063,N_333);
or U8155 (N_8155,N_1189,N_2650);
nand U8156 (N_8156,N_1455,N_446);
and U8157 (N_8157,N_1386,N_1472);
xor U8158 (N_8158,N_3402,N_3336);
or U8159 (N_8159,N_2761,N_939);
or U8160 (N_8160,N_2209,N_1642);
or U8161 (N_8161,N_2935,N_3806);
and U8162 (N_8162,N_2021,N_724);
xnor U8163 (N_8163,N_4360,N_3621);
xor U8164 (N_8164,N_118,N_1110);
nor U8165 (N_8165,N_3547,N_2126);
xnor U8166 (N_8166,N_675,N_1051);
nand U8167 (N_8167,N_2921,N_216);
xnor U8168 (N_8168,N_1641,N_3074);
or U8169 (N_8169,N_2601,N_488);
xor U8170 (N_8170,N_2064,N_3836);
xnor U8171 (N_8171,N_2929,N_1247);
xnor U8172 (N_8172,N_649,N_906);
or U8173 (N_8173,N_2014,N_746);
nand U8174 (N_8174,N_4645,N_3645);
nor U8175 (N_8175,N_2678,N_4692);
or U8176 (N_8176,N_4473,N_2963);
nor U8177 (N_8177,N_1118,N_2955);
or U8178 (N_8178,N_1253,N_2577);
nor U8179 (N_8179,N_4512,N_732);
xnor U8180 (N_8180,N_2510,N_3809);
nor U8181 (N_8181,N_2416,N_1934);
and U8182 (N_8182,N_482,N_3906);
and U8183 (N_8183,N_4127,N_4192);
nand U8184 (N_8184,N_2040,N_2036);
or U8185 (N_8185,N_3397,N_462);
nor U8186 (N_8186,N_3470,N_2946);
and U8187 (N_8187,N_227,N_3333);
or U8188 (N_8188,N_2398,N_1171);
nand U8189 (N_8189,N_1855,N_4508);
or U8190 (N_8190,N_3686,N_2986);
xnor U8191 (N_8191,N_436,N_346);
and U8192 (N_8192,N_1789,N_2398);
nand U8193 (N_8193,N_797,N_1040);
nor U8194 (N_8194,N_4846,N_2649);
and U8195 (N_8195,N_132,N_627);
and U8196 (N_8196,N_716,N_851);
xnor U8197 (N_8197,N_492,N_1266);
or U8198 (N_8198,N_4057,N_3759);
nand U8199 (N_8199,N_2571,N_3217);
or U8200 (N_8200,N_3734,N_2368);
nor U8201 (N_8201,N_4242,N_3113);
or U8202 (N_8202,N_365,N_3437);
and U8203 (N_8203,N_3142,N_3051);
and U8204 (N_8204,N_3518,N_622);
nor U8205 (N_8205,N_2076,N_3300);
nor U8206 (N_8206,N_645,N_4643);
and U8207 (N_8207,N_1957,N_4580);
and U8208 (N_8208,N_2870,N_2757);
and U8209 (N_8209,N_3235,N_2831);
xnor U8210 (N_8210,N_635,N_4507);
xor U8211 (N_8211,N_3590,N_4234);
xnor U8212 (N_8212,N_2091,N_3096);
xor U8213 (N_8213,N_4051,N_2556);
xor U8214 (N_8214,N_347,N_3476);
nand U8215 (N_8215,N_2404,N_1591);
and U8216 (N_8216,N_678,N_2931);
or U8217 (N_8217,N_387,N_2102);
or U8218 (N_8218,N_2085,N_93);
or U8219 (N_8219,N_3078,N_2774);
nand U8220 (N_8220,N_750,N_4931);
nor U8221 (N_8221,N_1733,N_631);
nand U8222 (N_8222,N_4100,N_969);
xnor U8223 (N_8223,N_1159,N_299);
or U8224 (N_8224,N_2983,N_416);
nand U8225 (N_8225,N_1217,N_3271);
or U8226 (N_8226,N_3935,N_1656);
xnor U8227 (N_8227,N_4362,N_69);
or U8228 (N_8228,N_4591,N_1709);
nand U8229 (N_8229,N_3752,N_2417);
nor U8230 (N_8230,N_2644,N_467);
nand U8231 (N_8231,N_3428,N_3175);
or U8232 (N_8232,N_4237,N_4059);
xor U8233 (N_8233,N_2588,N_3768);
xor U8234 (N_8234,N_434,N_4142);
or U8235 (N_8235,N_150,N_4570);
nand U8236 (N_8236,N_2600,N_1373);
nor U8237 (N_8237,N_775,N_4195);
xor U8238 (N_8238,N_1908,N_4560);
nor U8239 (N_8239,N_2518,N_2478);
xnor U8240 (N_8240,N_2429,N_1142);
nand U8241 (N_8241,N_2790,N_1211);
nor U8242 (N_8242,N_2431,N_4640);
xor U8243 (N_8243,N_1757,N_1693);
nand U8244 (N_8244,N_3824,N_767);
and U8245 (N_8245,N_3134,N_4145);
nor U8246 (N_8246,N_3558,N_1785);
or U8247 (N_8247,N_2695,N_4757);
and U8248 (N_8248,N_17,N_1757);
xnor U8249 (N_8249,N_2640,N_3008);
nor U8250 (N_8250,N_2644,N_2347);
nand U8251 (N_8251,N_1980,N_1214);
nand U8252 (N_8252,N_2771,N_603);
xor U8253 (N_8253,N_1888,N_440);
or U8254 (N_8254,N_4218,N_2405);
nand U8255 (N_8255,N_1052,N_2145);
xnor U8256 (N_8256,N_4064,N_1526);
and U8257 (N_8257,N_4497,N_3490);
nor U8258 (N_8258,N_698,N_1592);
xor U8259 (N_8259,N_1723,N_3099);
and U8260 (N_8260,N_4794,N_564);
nand U8261 (N_8261,N_3272,N_4563);
nor U8262 (N_8262,N_1962,N_998);
nor U8263 (N_8263,N_1024,N_167);
xnor U8264 (N_8264,N_2224,N_3658);
xnor U8265 (N_8265,N_383,N_1630);
and U8266 (N_8266,N_4548,N_2463);
nor U8267 (N_8267,N_1073,N_1531);
nor U8268 (N_8268,N_1744,N_715);
or U8269 (N_8269,N_1968,N_3061);
and U8270 (N_8270,N_3136,N_4103);
xor U8271 (N_8271,N_813,N_2875);
or U8272 (N_8272,N_3685,N_4909);
nand U8273 (N_8273,N_4156,N_1104);
nor U8274 (N_8274,N_2201,N_937);
or U8275 (N_8275,N_3064,N_320);
nor U8276 (N_8276,N_4273,N_2415);
xor U8277 (N_8277,N_482,N_4701);
nor U8278 (N_8278,N_1532,N_2655);
nor U8279 (N_8279,N_3175,N_953);
or U8280 (N_8280,N_867,N_1249);
xor U8281 (N_8281,N_788,N_2762);
and U8282 (N_8282,N_656,N_421);
xnor U8283 (N_8283,N_1111,N_3893);
and U8284 (N_8284,N_3899,N_502);
nor U8285 (N_8285,N_803,N_2543);
nand U8286 (N_8286,N_1675,N_3171);
and U8287 (N_8287,N_3158,N_324);
xnor U8288 (N_8288,N_4030,N_1960);
xnor U8289 (N_8289,N_3225,N_2493);
nand U8290 (N_8290,N_3250,N_4724);
nor U8291 (N_8291,N_2655,N_1498);
xor U8292 (N_8292,N_3961,N_566);
nor U8293 (N_8293,N_94,N_395);
or U8294 (N_8294,N_893,N_2622);
nor U8295 (N_8295,N_2513,N_685);
and U8296 (N_8296,N_4443,N_1723);
and U8297 (N_8297,N_659,N_2863);
or U8298 (N_8298,N_3501,N_4303);
nor U8299 (N_8299,N_4306,N_4635);
xnor U8300 (N_8300,N_1302,N_4355);
and U8301 (N_8301,N_4846,N_2027);
xor U8302 (N_8302,N_4944,N_3441);
nor U8303 (N_8303,N_648,N_4940);
xnor U8304 (N_8304,N_2224,N_552);
nand U8305 (N_8305,N_3344,N_463);
xnor U8306 (N_8306,N_1218,N_180);
xor U8307 (N_8307,N_4218,N_3786);
nor U8308 (N_8308,N_3891,N_4180);
nand U8309 (N_8309,N_1404,N_3295);
nor U8310 (N_8310,N_577,N_2025);
and U8311 (N_8311,N_54,N_4151);
or U8312 (N_8312,N_3260,N_3289);
nand U8313 (N_8313,N_4485,N_3564);
and U8314 (N_8314,N_103,N_2668);
nand U8315 (N_8315,N_1855,N_1770);
and U8316 (N_8316,N_371,N_246);
and U8317 (N_8317,N_1927,N_4646);
nand U8318 (N_8318,N_4727,N_4331);
or U8319 (N_8319,N_1613,N_1752);
or U8320 (N_8320,N_105,N_872);
xor U8321 (N_8321,N_904,N_4148);
nand U8322 (N_8322,N_4974,N_3325);
nand U8323 (N_8323,N_3318,N_56);
nand U8324 (N_8324,N_154,N_940);
nor U8325 (N_8325,N_2198,N_4165);
and U8326 (N_8326,N_2975,N_838);
or U8327 (N_8327,N_2969,N_4681);
and U8328 (N_8328,N_1822,N_4138);
xnor U8329 (N_8329,N_1370,N_26);
and U8330 (N_8330,N_280,N_4629);
nor U8331 (N_8331,N_3378,N_3837);
nand U8332 (N_8332,N_61,N_4103);
xor U8333 (N_8333,N_3587,N_4724);
or U8334 (N_8334,N_55,N_1808);
nor U8335 (N_8335,N_2068,N_1753);
xor U8336 (N_8336,N_50,N_2159);
xnor U8337 (N_8337,N_4381,N_4780);
nor U8338 (N_8338,N_3617,N_3808);
nor U8339 (N_8339,N_3005,N_1027);
or U8340 (N_8340,N_3225,N_1662);
xor U8341 (N_8341,N_1300,N_1236);
or U8342 (N_8342,N_2730,N_565);
nand U8343 (N_8343,N_2158,N_1847);
and U8344 (N_8344,N_1231,N_2704);
or U8345 (N_8345,N_3254,N_2687);
nand U8346 (N_8346,N_549,N_969);
and U8347 (N_8347,N_2878,N_4648);
xnor U8348 (N_8348,N_4725,N_1774);
or U8349 (N_8349,N_4011,N_982);
and U8350 (N_8350,N_4256,N_3098);
xor U8351 (N_8351,N_2976,N_983);
nand U8352 (N_8352,N_1455,N_422);
and U8353 (N_8353,N_4837,N_2896);
and U8354 (N_8354,N_3300,N_3960);
nor U8355 (N_8355,N_32,N_3348);
xor U8356 (N_8356,N_1331,N_1224);
xnor U8357 (N_8357,N_4364,N_3426);
nand U8358 (N_8358,N_4920,N_349);
nand U8359 (N_8359,N_4493,N_430);
nor U8360 (N_8360,N_4909,N_1188);
or U8361 (N_8361,N_3980,N_2343);
or U8362 (N_8362,N_2119,N_3286);
nand U8363 (N_8363,N_4248,N_4553);
xor U8364 (N_8364,N_1910,N_715);
xor U8365 (N_8365,N_3720,N_2601);
nand U8366 (N_8366,N_68,N_1880);
or U8367 (N_8367,N_1507,N_1022);
xnor U8368 (N_8368,N_2301,N_2794);
nand U8369 (N_8369,N_1949,N_3632);
nor U8370 (N_8370,N_3641,N_186);
xnor U8371 (N_8371,N_3751,N_4733);
and U8372 (N_8372,N_2263,N_3807);
or U8373 (N_8373,N_3225,N_2932);
or U8374 (N_8374,N_2558,N_2152);
nand U8375 (N_8375,N_3284,N_4815);
xnor U8376 (N_8376,N_730,N_2754);
nor U8377 (N_8377,N_220,N_2866);
and U8378 (N_8378,N_534,N_860);
and U8379 (N_8379,N_4588,N_952);
xor U8380 (N_8380,N_2738,N_2160);
xor U8381 (N_8381,N_831,N_3634);
and U8382 (N_8382,N_4388,N_4339);
nand U8383 (N_8383,N_2332,N_4651);
and U8384 (N_8384,N_4155,N_3032);
nand U8385 (N_8385,N_412,N_580);
or U8386 (N_8386,N_3260,N_3275);
nor U8387 (N_8387,N_1600,N_255);
or U8388 (N_8388,N_3943,N_2301);
and U8389 (N_8389,N_1241,N_1456);
xnor U8390 (N_8390,N_705,N_1345);
and U8391 (N_8391,N_208,N_24);
or U8392 (N_8392,N_3945,N_4213);
and U8393 (N_8393,N_1465,N_3013);
xor U8394 (N_8394,N_4208,N_1512);
and U8395 (N_8395,N_4292,N_2493);
xnor U8396 (N_8396,N_891,N_552);
or U8397 (N_8397,N_485,N_467);
xnor U8398 (N_8398,N_4112,N_2206);
or U8399 (N_8399,N_4338,N_1825);
and U8400 (N_8400,N_4489,N_4674);
nor U8401 (N_8401,N_2110,N_1128);
and U8402 (N_8402,N_4863,N_1973);
nor U8403 (N_8403,N_2535,N_1463);
nand U8404 (N_8404,N_1053,N_2245);
nand U8405 (N_8405,N_1720,N_1232);
nor U8406 (N_8406,N_4892,N_2939);
xnor U8407 (N_8407,N_2260,N_4667);
nand U8408 (N_8408,N_139,N_2224);
nor U8409 (N_8409,N_367,N_2226);
xnor U8410 (N_8410,N_3360,N_2432);
xnor U8411 (N_8411,N_3880,N_3930);
nor U8412 (N_8412,N_2223,N_4857);
nor U8413 (N_8413,N_1532,N_4506);
nor U8414 (N_8414,N_4055,N_2724);
nor U8415 (N_8415,N_760,N_3658);
nand U8416 (N_8416,N_4713,N_77);
and U8417 (N_8417,N_2552,N_456);
or U8418 (N_8418,N_2392,N_3816);
and U8419 (N_8419,N_2127,N_134);
xnor U8420 (N_8420,N_1121,N_3057);
nand U8421 (N_8421,N_3998,N_4591);
or U8422 (N_8422,N_621,N_2883);
and U8423 (N_8423,N_331,N_4020);
and U8424 (N_8424,N_3302,N_1308);
and U8425 (N_8425,N_1492,N_4151);
and U8426 (N_8426,N_2311,N_3205);
xor U8427 (N_8427,N_4210,N_772);
xnor U8428 (N_8428,N_2973,N_15);
xnor U8429 (N_8429,N_2775,N_4366);
or U8430 (N_8430,N_1931,N_4370);
nor U8431 (N_8431,N_2615,N_2962);
nand U8432 (N_8432,N_2080,N_141);
nor U8433 (N_8433,N_4637,N_3364);
or U8434 (N_8434,N_1160,N_2472);
nand U8435 (N_8435,N_2839,N_1310);
nand U8436 (N_8436,N_4799,N_4371);
nor U8437 (N_8437,N_3598,N_4969);
or U8438 (N_8438,N_4842,N_2868);
or U8439 (N_8439,N_3567,N_4701);
nand U8440 (N_8440,N_83,N_2209);
or U8441 (N_8441,N_4976,N_749);
nor U8442 (N_8442,N_3933,N_4605);
xor U8443 (N_8443,N_198,N_4154);
nor U8444 (N_8444,N_4578,N_1305);
and U8445 (N_8445,N_2646,N_3343);
nand U8446 (N_8446,N_653,N_3268);
xor U8447 (N_8447,N_150,N_3059);
and U8448 (N_8448,N_3290,N_1038);
or U8449 (N_8449,N_2000,N_2061);
nor U8450 (N_8450,N_3958,N_954);
nand U8451 (N_8451,N_3390,N_3323);
nand U8452 (N_8452,N_584,N_1614);
nand U8453 (N_8453,N_1905,N_1504);
xor U8454 (N_8454,N_267,N_3465);
and U8455 (N_8455,N_633,N_3099);
xor U8456 (N_8456,N_4569,N_2178);
nand U8457 (N_8457,N_3328,N_1558);
or U8458 (N_8458,N_1527,N_2665);
xnor U8459 (N_8459,N_1194,N_3818);
nand U8460 (N_8460,N_3807,N_4905);
xor U8461 (N_8461,N_2967,N_4075);
xor U8462 (N_8462,N_1206,N_1121);
xnor U8463 (N_8463,N_940,N_3684);
or U8464 (N_8464,N_4978,N_1780);
or U8465 (N_8465,N_4024,N_3808);
or U8466 (N_8466,N_2096,N_762);
nand U8467 (N_8467,N_837,N_1983);
nor U8468 (N_8468,N_2349,N_1760);
xnor U8469 (N_8469,N_4535,N_1338);
or U8470 (N_8470,N_1436,N_830);
and U8471 (N_8471,N_598,N_4587);
and U8472 (N_8472,N_1866,N_3510);
xnor U8473 (N_8473,N_917,N_4609);
nor U8474 (N_8474,N_360,N_3766);
or U8475 (N_8475,N_628,N_2493);
and U8476 (N_8476,N_1258,N_2687);
nand U8477 (N_8477,N_2728,N_4783);
and U8478 (N_8478,N_2085,N_3773);
nor U8479 (N_8479,N_3719,N_3127);
nor U8480 (N_8480,N_2782,N_4875);
nor U8481 (N_8481,N_3133,N_3966);
or U8482 (N_8482,N_3105,N_777);
nor U8483 (N_8483,N_1320,N_353);
and U8484 (N_8484,N_131,N_2822);
and U8485 (N_8485,N_22,N_734);
xor U8486 (N_8486,N_2564,N_2376);
nand U8487 (N_8487,N_1558,N_2373);
nand U8488 (N_8488,N_3138,N_2819);
and U8489 (N_8489,N_3143,N_895);
xnor U8490 (N_8490,N_4910,N_1156);
xor U8491 (N_8491,N_4161,N_2770);
or U8492 (N_8492,N_933,N_3983);
nor U8493 (N_8493,N_1913,N_4399);
nand U8494 (N_8494,N_3638,N_1107);
or U8495 (N_8495,N_4094,N_2043);
xnor U8496 (N_8496,N_4079,N_3502);
nor U8497 (N_8497,N_1678,N_1235);
or U8498 (N_8498,N_3366,N_461);
xnor U8499 (N_8499,N_3253,N_4123);
nor U8500 (N_8500,N_4377,N_2311);
nand U8501 (N_8501,N_165,N_3174);
or U8502 (N_8502,N_2412,N_311);
or U8503 (N_8503,N_2032,N_139);
nand U8504 (N_8504,N_1568,N_495);
or U8505 (N_8505,N_1898,N_738);
and U8506 (N_8506,N_1158,N_1395);
nor U8507 (N_8507,N_846,N_4334);
or U8508 (N_8508,N_3746,N_2468);
and U8509 (N_8509,N_1934,N_1695);
xnor U8510 (N_8510,N_296,N_3111);
xnor U8511 (N_8511,N_975,N_2661);
and U8512 (N_8512,N_4734,N_4168);
and U8513 (N_8513,N_2760,N_2198);
and U8514 (N_8514,N_4213,N_4774);
nor U8515 (N_8515,N_1350,N_4700);
xor U8516 (N_8516,N_32,N_4952);
and U8517 (N_8517,N_2749,N_4756);
nor U8518 (N_8518,N_3525,N_4023);
nand U8519 (N_8519,N_3205,N_1655);
nand U8520 (N_8520,N_1361,N_4679);
nor U8521 (N_8521,N_1533,N_1201);
nand U8522 (N_8522,N_1313,N_769);
nand U8523 (N_8523,N_3764,N_4346);
or U8524 (N_8524,N_3790,N_2288);
or U8525 (N_8525,N_3088,N_857);
xor U8526 (N_8526,N_4130,N_2218);
nand U8527 (N_8527,N_3061,N_255);
or U8528 (N_8528,N_795,N_3691);
nor U8529 (N_8529,N_4760,N_1963);
and U8530 (N_8530,N_3037,N_1180);
or U8531 (N_8531,N_3010,N_3488);
or U8532 (N_8532,N_668,N_2280);
or U8533 (N_8533,N_4157,N_4907);
or U8534 (N_8534,N_394,N_4384);
or U8535 (N_8535,N_3290,N_2619);
nor U8536 (N_8536,N_1769,N_919);
or U8537 (N_8537,N_2459,N_4267);
xor U8538 (N_8538,N_343,N_4643);
and U8539 (N_8539,N_3002,N_1971);
xor U8540 (N_8540,N_4039,N_2296);
or U8541 (N_8541,N_3476,N_767);
or U8542 (N_8542,N_1430,N_9);
or U8543 (N_8543,N_973,N_972);
xor U8544 (N_8544,N_1984,N_1033);
nor U8545 (N_8545,N_4230,N_4670);
xor U8546 (N_8546,N_838,N_2563);
or U8547 (N_8547,N_2145,N_237);
nor U8548 (N_8548,N_4180,N_2780);
nand U8549 (N_8549,N_3835,N_902);
xnor U8550 (N_8550,N_2027,N_1306);
or U8551 (N_8551,N_2041,N_1102);
nand U8552 (N_8552,N_4403,N_679);
xor U8553 (N_8553,N_1081,N_3613);
xor U8554 (N_8554,N_3659,N_1967);
nor U8555 (N_8555,N_3793,N_4794);
or U8556 (N_8556,N_2696,N_4255);
or U8557 (N_8557,N_1860,N_25);
or U8558 (N_8558,N_1903,N_4109);
xnor U8559 (N_8559,N_1064,N_593);
nor U8560 (N_8560,N_3905,N_711);
nor U8561 (N_8561,N_390,N_1707);
or U8562 (N_8562,N_4349,N_4071);
nor U8563 (N_8563,N_604,N_4268);
nand U8564 (N_8564,N_164,N_4398);
nand U8565 (N_8565,N_803,N_3956);
nor U8566 (N_8566,N_2926,N_1352);
nor U8567 (N_8567,N_2896,N_4784);
xnor U8568 (N_8568,N_3121,N_2153);
xnor U8569 (N_8569,N_446,N_2693);
xor U8570 (N_8570,N_3151,N_4156);
and U8571 (N_8571,N_220,N_3086);
or U8572 (N_8572,N_4943,N_3704);
or U8573 (N_8573,N_3148,N_4682);
xnor U8574 (N_8574,N_307,N_1610);
nor U8575 (N_8575,N_106,N_1089);
nor U8576 (N_8576,N_1394,N_1035);
nor U8577 (N_8577,N_2476,N_4557);
or U8578 (N_8578,N_2970,N_4958);
xnor U8579 (N_8579,N_1489,N_1697);
or U8580 (N_8580,N_715,N_2074);
or U8581 (N_8581,N_1169,N_4337);
xnor U8582 (N_8582,N_810,N_2206);
xor U8583 (N_8583,N_2489,N_4472);
or U8584 (N_8584,N_2512,N_4522);
or U8585 (N_8585,N_4090,N_2301);
xor U8586 (N_8586,N_4264,N_1704);
nand U8587 (N_8587,N_2335,N_314);
nor U8588 (N_8588,N_4537,N_297);
xor U8589 (N_8589,N_4787,N_4877);
and U8590 (N_8590,N_2922,N_4251);
nor U8591 (N_8591,N_4086,N_2491);
or U8592 (N_8592,N_477,N_2024);
xnor U8593 (N_8593,N_2302,N_19);
xor U8594 (N_8594,N_1288,N_3448);
nand U8595 (N_8595,N_3489,N_1921);
xor U8596 (N_8596,N_3546,N_936);
nand U8597 (N_8597,N_31,N_104);
and U8598 (N_8598,N_2608,N_1339);
and U8599 (N_8599,N_4692,N_2260);
xnor U8600 (N_8600,N_4433,N_170);
nor U8601 (N_8601,N_587,N_3576);
and U8602 (N_8602,N_2603,N_371);
xnor U8603 (N_8603,N_4020,N_3071);
and U8604 (N_8604,N_3558,N_3122);
nand U8605 (N_8605,N_2295,N_3346);
or U8606 (N_8606,N_2079,N_1891);
nor U8607 (N_8607,N_345,N_4318);
xnor U8608 (N_8608,N_4769,N_2371);
nor U8609 (N_8609,N_1759,N_187);
nand U8610 (N_8610,N_4750,N_486);
nor U8611 (N_8611,N_4783,N_1133);
xnor U8612 (N_8612,N_2518,N_2753);
nor U8613 (N_8613,N_2000,N_1991);
xnor U8614 (N_8614,N_4429,N_2696);
nor U8615 (N_8615,N_4514,N_3872);
or U8616 (N_8616,N_638,N_3583);
xor U8617 (N_8617,N_762,N_2169);
nor U8618 (N_8618,N_4187,N_3667);
xnor U8619 (N_8619,N_1721,N_867);
nor U8620 (N_8620,N_772,N_4901);
nand U8621 (N_8621,N_728,N_992);
nor U8622 (N_8622,N_2641,N_3927);
nand U8623 (N_8623,N_4476,N_2923);
nor U8624 (N_8624,N_3166,N_3696);
nor U8625 (N_8625,N_332,N_3343);
nand U8626 (N_8626,N_3102,N_2062);
nor U8627 (N_8627,N_1123,N_54);
nor U8628 (N_8628,N_333,N_3545);
xnor U8629 (N_8629,N_358,N_3763);
nand U8630 (N_8630,N_4072,N_1293);
nor U8631 (N_8631,N_1399,N_2805);
xor U8632 (N_8632,N_322,N_3223);
and U8633 (N_8633,N_1340,N_1817);
nor U8634 (N_8634,N_3725,N_1534);
xor U8635 (N_8635,N_2048,N_519);
nor U8636 (N_8636,N_2521,N_1336);
nor U8637 (N_8637,N_2372,N_156);
xor U8638 (N_8638,N_1162,N_2533);
or U8639 (N_8639,N_693,N_3379);
nor U8640 (N_8640,N_230,N_2523);
xnor U8641 (N_8641,N_189,N_2295);
xor U8642 (N_8642,N_2445,N_4247);
and U8643 (N_8643,N_3377,N_2624);
xnor U8644 (N_8644,N_371,N_2600);
nand U8645 (N_8645,N_2462,N_1572);
xnor U8646 (N_8646,N_4570,N_3739);
nand U8647 (N_8647,N_3773,N_3050);
nand U8648 (N_8648,N_3455,N_1705);
nand U8649 (N_8649,N_3873,N_4974);
and U8650 (N_8650,N_2377,N_4186);
nor U8651 (N_8651,N_1251,N_1180);
nand U8652 (N_8652,N_1944,N_905);
nor U8653 (N_8653,N_168,N_3240);
and U8654 (N_8654,N_263,N_1616);
nor U8655 (N_8655,N_4451,N_4851);
nor U8656 (N_8656,N_2650,N_3585);
and U8657 (N_8657,N_3216,N_3086);
nor U8658 (N_8658,N_2143,N_3424);
nand U8659 (N_8659,N_650,N_1784);
nand U8660 (N_8660,N_1564,N_4812);
and U8661 (N_8661,N_684,N_2728);
nor U8662 (N_8662,N_4728,N_1273);
xnor U8663 (N_8663,N_423,N_1799);
or U8664 (N_8664,N_4058,N_2091);
nor U8665 (N_8665,N_3961,N_2315);
and U8666 (N_8666,N_1905,N_2181);
nor U8667 (N_8667,N_217,N_1006);
and U8668 (N_8668,N_1021,N_1407);
nand U8669 (N_8669,N_238,N_729);
nor U8670 (N_8670,N_2532,N_1530);
nand U8671 (N_8671,N_460,N_1131);
nor U8672 (N_8672,N_1514,N_748);
and U8673 (N_8673,N_3624,N_3114);
or U8674 (N_8674,N_4117,N_2495);
nor U8675 (N_8675,N_1726,N_4986);
nand U8676 (N_8676,N_4451,N_3123);
and U8677 (N_8677,N_3868,N_2962);
nand U8678 (N_8678,N_1065,N_3539);
nor U8679 (N_8679,N_1013,N_713);
nand U8680 (N_8680,N_886,N_3542);
and U8681 (N_8681,N_3799,N_1160);
nand U8682 (N_8682,N_623,N_1810);
nor U8683 (N_8683,N_3137,N_4550);
nor U8684 (N_8684,N_1487,N_4025);
and U8685 (N_8685,N_613,N_1590);
nor U8686 (N_8686,N_4820,N_90);
or U8687 (N_8687,N_2085,N_2335);
nor U8688 (N_8688,N_3704,N_1387);
and U8689 (N_8689,N_1938,N_4759);
nand U8690 (N_8690,N_2359,N_2358);
or U8691 (N_8691,N_2423,N_2531);
xnor U8692 (N_8692,N_4408,N_354);
nand U8693 (N_8693,N_2402,N_4222);
nor U8694 (N_8694,N_58,N_867);
nor U8695 (N_8695,N_4036,N_597);
or U8696 (N_8696,N_1751,N_3882);
or U8697 (N_8697,N_1413,N_4215);
or U8698 (N_8698,N_455,N_472);
nand U8699 (N_8699,N_1698,N_236);
nand U8700 (N_8700,N_2895,N_1503);
or U8701 (N_8701,N_298,N_3623);
nand U8702 (N_8702,N_2420,N_4239);
nor U8703 (N_8703,N_950,N_4603);
nor U8704 (N_8704,N_2087,N_3512);
nand U8705 (N_8705,N_3720,N_1727);
nor U8706 (N_8706,N_2007,N_1916);
and U8707 (N_8707,N_3603,N_3722);
xor U8708 (N_8708,N_3174,N_2438);
and U8709 (N_8709,N_937,N_4556);
or U8710 (N_8710,N_244,N_2594);
nand U8711 (N_8711,N_3955,N_4402);
or U8712 (N_8712,N_3257,N_1675);
nor U8713 (N_8713,N_4009,N_1610);
nand U8714 (N_8714,N_3720,N_117);
or U8715 (N_8715,N_1966,N_2998);
and U8716 (N_8716,N_3263,N_4008);
and U8717 (N_8717,N_3045,N_1543);
nand U8718 (N_8718,N_416,N_4757);
xnor U8719 (N_8719,N_1467,N_3152);
xor U8720 (N_8720,N_1939,N_535);
nor U8721 (N_8721,N_919,N_891);
xor U8722 (N_8722,N_1309,N_3753);
and U8723 (N_8723,N_3125,N_1062);
nand U8724 (N_8724,N_2342,N_201);
and U8725 (N_8725,N_2699,N_3655);
nand U8726 (N_8726,N_2913,N_1526);
nand U8727 (N_8727,N_3162,N_2378);
nand U8728 (N_8728,N_4518,N_2737);
nor U8729 (N_8729,N_4426,N_449);
nand U8730 (N_8730,N_933,N_2907);
and U8731 (N_8731,N_4184,N_3630);
and U8732 (N_8732,N_4144,N_842);
or U8733 (N_8733,N_4013,N_389);
or U8734 (N_8734,N_2234,N_3949);
xor U8735 (N_8735,N_732,N_1623);
and U8736 (N_8736,N_158,N_2931);
and U8737 (N_8737,N_386,N_1153);
or U8738 (N_8738,N_3552,N_403);
and U8739 (N_8739,N_2390,N_264);
or U8740 (N_8740,N_1791,N_2882);
xnor U8741 (N_8741,N_1116,N_3572);
or U8742 (N_8742,N_3148,N_1564);
nand U8743 (N_8743,N_365,N_1943);
nor U8744 (N_8744,N_870,N_2708);
and U8745 (N_8745,N_1550,N_1479);
or U8746 (N_8746,N_3497,N_2148);
xor U8747 (N_8747,N_760,N_824);
nor U8748 (N_8748,N_1111,N_2357);
xnor U8749 (N_8749,N_4833,N_2529);
and U8750 (N_8750,N_2211,N_2333);
nand U8751 (N_8751,N_2423,N_2131);
or U8752 (N_8752,N_2838,N_3456);
xor U8753 (N_8753,N_4138,N_4038);
and U8754 (N_8754,N_4707,N_2246);
xor U8755 (N_8755,N_4928,N_3908);
and U8756 (N_8756,N_3244,N_505);
or U8757 (N_8757,N_4131,N_4779);
nor U8758 (N_8758,N_3094,N_2712);
nand U8759 (N_8759,N_3187,N_4994);
nand U8760 (N_8760,N_1101,N_167);
nor U8761 (N_8761,N_2249,N_2830);
nor U8762 (N_8762,N_1636,N_3266);
and U8763 (N_8763,N_2126,N_3656);
nand U8764 (N_8764,N_3956,N_4204);
and U8765 (N_8765,N_2796,N_4735);
nor U8766 (N_8766,N_2791,N_3292);
xor U8767 (N_8767,N_1227,N_3252);
xnor U8768 (N_8768,N_491,N_3601);
or U8769 (N_8769,N_1913,N_1378);
nor U8770 (N_8770,N_3644,N_2984);
and U8771 (N_8771,N_4360,N_4747);
xnor U8772 (N_8772,N_3810,N_2404);
nand U8773 (N_8773,N_3244,N_730);
nand U8774 (N_8774,N_471,N_4677);
xor U8775 (N_8775,N_3758,N_4451);
xnor U8776 (N_8776,N_4721,N_4917);
nor U8777 (N_8777,N_2072,N_2199);
xnor U8778 (N_8778,N_26,N_1811);
nand U8779 (N_8779,N_2596,N_1051);
nor U8780 (N_8780,N_3791,N_2233);
xor U8781 (N_8781,N_3775,N_1474);
and U8782 (N_8782,N_1789,N_3520);
or U8783 (N_8783,N_541,N_4359);
xor U8784 (N_8784,N_3660,N_46);
and U8785 (N_8785,N_4486,N_4511);
nand U8786 (N_8786,N_2571,N_4253);
nand U8787 (N_8787,N_4137,N_1353);
nand U8788 (N_8788,N_2567,N_2810);
and U8789 (N_8789,N_654,N_808);
nor U8790 (N_8790,N_3684,N_1582);
nor U8791 (N_8791,N_1887,N_4807);
nor U8792 (N_8792,N_2841,N_716);
or U8793 (N_8793,N_3243,N_4039);
nor U8794 (N_8794,N_3501,N_4783);
xnor U8795 (N_8795,N_298,N_317);
nor U8796 (N_8796,N_1708,N_2222);
nor U8797 (N_8797,N_2540,N_3935);
xor U8798 (N_8798,N_3292,N_232);
nand U8799 (N_8799,N_675,N_199);
xnor U8800 (N_8800,N_3499,N_4366);
nor U8801 (N_8801,N_1507,N_2381);
and U8802 (N_8802,N_1596,N_3482);
xnor U8803 (N_8803,N_2322,N_4437);
xor U8804 (N_8804,N_4736,N_674);
nor U8805 (N_8805,N_1101,N_529);
nor U8806 (N_8806,N_4278,N_4844);
nor U8807 (N_8807,N_2880,N_1811);
nand U8808 (N_8808,N_919,N_1419);
and U8809 (N_8809,N_1376,N_3238);
nor U8810 (N_8810,N_3169,N_3637);
xor U8811 (N_8811,N_3521,N_4797);
xor U8812 (N_8812,N_2004,N_4167);
and U8813 (N_8813,N_2808,N_1732);
nand U8814 (N_8814,N_1931,N_4153);
nor U8815 (N_8815,N_1782,N_147);
xnor U8816 (N_8816,N_2982,N_2796);
xnor U8817 (N_8817,N_1093,N_1683);
or U8818 (N_8818,N_4543,N_4629);
or U8819 (N_8819,N_3833,N_4971);
and U8820 (N_8820,N_392,N_4129);
nand U8821 (N_8821,N_534,N_4654);
and U8822 (N_8822,N_2912,N_4128);
nor U8823 (N_8823,N_3345,N_2054);
and U8824 (N_8824,N_4184,N_3946);
nand U8825 (N_8825,N_3471,N_1247);
nor U8826 (N_8826,N_276,N_1935);
or U8827 (N_8827,N_3137,N_2129);
nand U8828 (N_8828,N_970,N_1678);
or U8829 (N_8829,N_3627,N_2708);
nand U8830 (N_8830,N_4965,N_1484);
xor U8831 (N_8831,N_3817,N_3209);
nand U8832 (N_8832,N_4756,N_3827);
xnor U8833 (N_8833,N_2560,N_2639);
nand U8834 (N_8834,N_726,N_4427);
nand U8835 (N_8835,N_4194,N_406);
and U8836 (N_8836,N_1146,N_3789);
nor U8837 (N_8837,N_1739,N_3724);
or U8838 (N_8838,N_225,N_2215);
xnor U8839 (N_8839,N_4637,N_3409);
nor U8840 (N_8840,N_118,N_1690);
nor U8841 (N_8841,N_1321,N_4314);
or U8842 (N_8842,N_2949,N_4269);
nor U8843 (N_8843,N_1035,N_2028);
nand U8844 (N_8844,N_2987,N_3099);
and U8845 (N_8845,N_4638,N_1148);
nor U8846 (N_8846,N_2606,N_1829);
and U8847 (N_8847,N_3245,N_4888);
nand U8848 (N_8848,N_3298,N_2613);
nor U8849 (N_8849,N_4219,N_3365);
or U8850 (N_8850,N_2012,N_4771);
or U8851 (N_8851,N_1649,N_4188);
nor U8852 (N_8852,N_3184,N_907);
or U8853 (N_8853,N_4511,N_1619);
or U8854 (N_8854,N_3002,N_1435);
xor U8855 (N_8855,N_1877,N_2584);
or U8856 (N_8856,N_3130,N_3813);
or U8857 (N_8857,N_4438,N_2932);
or U8858 (N_8858,N_4048,N_1986);
xnor U8859 (N_8859,N_2526,N_4336);
and U8860 (N_8860,N_4695,N_4268);
xor U8861 (N_8861,N_2412,N_1045);
nand U8862 (N_8862,N_1192,N_112);
xor U8863 (N_8863,N_3975,N_3194);
or U8864 (N_8864,N_1018,N_644);
and U8865 (N_8865,N_937,N_2966);
xnor U8866 (N_8866,N_1308,N_4189);
nor U8867 (N_8867,N_2680,N_3429);
nor U8868 (N_8868,N_1163,N_2336);
xnor U8869 (N_8869,N_4947,N_3897);
nand U8870 (N_8870,N_1001,N_1659);
or U8871 (N_8871,N_1500,N_4639);
nand U8872 (N_8872,N_370,N_3880);
nand U8873 (N_8873,N_1766,N_131);
nand U8874 (N_8874,N_1657,N_4204);
nand U8875 (N_8875,N_4323,N_2268);
and U8876 (N_8876,N_4186,N_3239);
xor U8877 (N_8877,N_4802,N_1435);
xnor U8878 (N_8878,N_3552,N_4955);
nand U8879 (N_8879,N_3295,N_978);
nor U8880 (N_8880,N_3718,N_1229);
or U8881 (N_8881,N_3494,N_4509);
nand U8882 (N_8882,N_87,N_2666);
nor U8883 (N_8883,N_4034,N_57);
xor U8884 (N_8884,N_2147,N_1495);
xor U8885 (N_8885,N_4848,N_4659);
nand U8886 (N_8886,N_3462,N_3919);
and U8887 (N_8887,N_4346,N_4403);
nor U8888 (N_8888,N_451,N_4222);
or U8889 (N_8889,N_4360,N_162);
nand U8890 (N_8890,N_388,N_4516);
and U8891 (N_8891,N_1301,N_308);
and U8892 (N_8892,N_191,N_362);
nand U8893 (N_8893,N_4706,N_2435);
and U8894 (N_8894,N_2353,N_3530);
nor U8895 (N_8895,N_4762,N_1474);
xor U8896 (N_8896,N_3996,N_1594);
xnor U8897 (N_8897,N_2243,N_3088);
nor U8898 (N_8898,N_3856,N_2045);
or U8899 (N_8899,N_896,N_675);
and U8900 (N_8900,N_2611,N_3580);
nand U8901 (N_8901,N_1936,N_3207);
nor U8902 (N_8902,N_2376,N_225);
or U8903 (N_8903,N_58,N_2114);
or U8904 (N_8904,N_906,N_4193);
nor U8905 (N_8905,N_1430,N_2689);
and U8906 (N_8906,N_497,N_1148);
nor U8907 (N_8907,N_971,N_426);
nand U8908 (N_8908,N_4029,N_4525);
nand U8909 (N_8909,N_3861,N_1812);
or U8910 (N_8910,N_767,N_686);
and U8911 (N_8911,N_3140,N_2190);
nand U8912 (N_8912,N_1845,N_3105);
nor U8913 (N_8913,N_2376,N_595);
nand U8914 (N_8914,N_2817,N_623);
or U8915 (N_8915,N_3372,N_2654);
and U8916 (N_8916,N_52,N_24);
xnor U8917 (N_8917,N_4600,N_4476);
nand U8918 (N_8918,N_3161,N_2255);
nor U8919 (N_8919,N_2891,N_1734);
and U8920 (N_8920,N_154,N_617);
or U8921 (N_8921,N_4654,N_1187);
and U8922 (N_8922,N_2816,N_2949);
nor U8923 (N_8923,N_4064,N_1139);
or U8924 (N_8924,N_4672,N_2292);
or U8925 (N_8925,N_4306,N_216);
and U8926 (N_8926,N_3974,N_1747);
xor U8927 (N_8927,N_3538,N_1657);
nand U8928 (N_8928,N_2306,N_4271);
xnor U8929 (N_8929,N_3064,N_4827);
or U8930 (N_8930,N_1985,N_4888);
or U8931 (N_8931,N_3732,N_1030);
nand U8932 (N_8932,N_2458,N_2259);
and U8933 (N_8933,N_4394,N_3328);
xor U8934 (N_8934,N_847,N_193);
xor U8935 (N_8935,N_4923,N_791);
or U8936 (N_8936,N_1542,N_3266);
or U8937 (N_8937,N_2630,N_3408);
xnor U8938 (N_8938,N_3988,N_139);
and U8939 (N_8939,N_3961,N_884);
and U8940 (N_8940,N_3998,N_2051);
xnor U8941 (N_8941,N_2558,N_4725);
nand U8942 (N_8942,N_3606,N_2667);
nor U8943 (N_8943,N_2292,N_3315);
xor U8944 (N_8944,N_1081,N_3232);
nand U8945 (N_8945,N_4806,N_4007);
and U8946 (N_8946,N_4683,N_1936);
xor U8947 (N_8947,N_4335,N_875);
nand U8948 (N_8948,N_532,N_277);
or U8949 (N_8949,N_2863,N_4950);
nand U8950 (N_8950,N_2219,N_1064);
and U8951 (N_8951,N_1393,N_3793);
or U8952 (N_8952,N_2748,N_3010);
nand U8953 (N_8953,N_4845,N_3389);
nand U8954 (N_8954,N_1063,N_3618);
nand U8955 (N_8955,N_164,N_4141);
nor U8956 (N_8956,N_957,N_878);
nor U8957 (N_8957,N_2247,N_2558);
nor U8958 (N_8958,N_3008,N_4625);
nor U8959 (N_8959,N_1160,N_2958);
nor U8960 (N_8960,N_3421,N_925);
or U8961 (N_8961,N_4250,N_945);
and U8962 (N_8962,N_2725,N_197);
xnor U8963 (N_8963,N_2018,N_983);
nor U8964 (N_8964,N_1637,N_333);
nor U8965 (N_8965,N_972,N_4577);
and U8966 (N_8966,N_162,N_2827);
or U8967 (N_8967,N_2109,N_252);
and U8968 (N_8968,N_4257,N_236);
nand U8969 (N_8969,N_2978,N_2501);
nor U8970 (N_8970,N_2975,N_935);
nand U8971 (N_8971,N_3010,N_3418);
nor U8972 (N_8972,N_3935,N_1732);
and U8973 (N_8973,N_1845,N_1406);
or U8974 (N_8974,N_4049,N_656);
and U8975 (N_8975,N_1107,N_1590);
xor U8976 (N_8976,N_569,N_469);
xor U8977 (N_8977,N_4531,N_2749);
or U8978 (N_8978,N_3632,N_1796);
nand U8979 (N_8979,N_374,N_810);
nand U8980 (N_8980,N_597,N_4581);
xnor U8981 (N_8981,N_2572,N_2527);
nand U8982 (N_8982,N_1474,N_813);
and U8983 (N_8983,N_3024,N_1303);
or U8984 (N_8984,N_600,N_369);
xor U8985 (N_8985,N_1073,N_2272);
nand U8986 (N_8986,N_3647,N_2636);
nand U8987 (N_8987,N_3552,N_3526);
and U8988 (N_8988,N_3796,N_3841);
xor U8989 (N_8989,N_3174,N_2148);
nor U8990 (N_8990,N_3116,N_4383);
and U8991 (N_8991,N_2964,N_4403);
xor U8992 (N_8992,N_1746,N_3772);
nand U8993 (N_8993,N_2126,N_3810);
and U8994 (N_8994,N_3750,N_1809);
and U8995 (N_8995,N_2756,N_1275);
xnor U8996 (N_8996,N_3842,N_1777);
nor U8997 (N_8997,N_1421,N_4275);
nor U8998 (N_8998,N_2249,N_2657);
xnor U8999 (N_8999,N_2869,N_610);
and U9000 (N_9000,N_1688,N_1173);
nor U9001 (N_9001,N_3634,N_3747);
xnor U9002 (N_9002,N_3586,N_711);
or U9003 (N_9003,N_3008,N_4287);
or U9004 (N_9004,N_3500,N_49);
xnor U9005 (N_9005,N_2322,N_4117);
nand U9006 (N_9006,N_1588,N_2868);
and U9007 (N_9007,N_2853,N_2222);
and U9008 (N_9008,N_4297,N_3433);
or U9009 (N_9009,N_320,N_3096);
or U9010 (N_9010,N_4565,N_2934);
or U9011 (N_9011,N_1097,N_2118);
or U9012 (N_9012,N_2347,N_4046);
nor U9013 (N_9013,N_3160,N_2080);
or U9014 (N_9014,N_2828,N_3114);
nor U9015 (N_9015,N_2884,N_1786);
nor U9016 (N_9016,N_4192,N_2483);
and U9017 (N_9017,N_1945,N_71);
and U9018 (N_9018,N_4178,N_562);
xnor U9019 (N_9019,N_4912,N_778);
and U9020 (N_9020,N_1180,N_3258);
xor U9021 (N_9021,N_516,N_2424);
nand U9022 (N_9022,N_4046,N_1475);
nor U9023 (N_9023,N_4552,N_2989);
or U9024 (N_9024,N_4984,N_543);
nor U9025 (N_9025,N_723,N_4106);
nand U9026 (N_9026,N_4036,N_1954);
xor U9027 (N_9027,N_3170,N_1053);
and U9028 (N_9028,N_4659,N_997);
nand U9029 (N_9029,N_1110,N_1862);
nor U9030 (N_9030,N_74,N_3123);
and U9031 (N_9031,N_3095,N_4097);
xor U9032 (N_9032,N_181,N_2669);
nor U9033 (N_9033,N_571,N_2898);
and U9034 (N_9034,N_4860,N_2156);
nand U9035 (N_9035,N_1473,N_2244);
nor U9036 (N_9036,N_1745,N_2557);
xnor U9037 (N_9037,N_2511,N_3005);
nor U9038 (N_9038,N_3164,N_2124);
and U9039 (N_9039,N_2872,N_3591);
xnor U9040 (N_9040,N_597,N_4821);
nand U9041 (N_9041,N_1022,N_793);
nor U9042 (N_9042,N_4638,N_2816);
xnor U9043 (N_9043,N_1829,N_677);
nor U9044 (N_9044,N_4635,N_305);
or U9045 (N_9045,N_4402,N_3350);
nand U9046 (N_9046,N_4246,N_3170);
nor U9047 (N_9047,N_2039,N_837);
xnor U9048 (N_9048,N_765,N_3782);
nand U9049 (N_9049,N_260,N_3232);
or U9050 (N_9050,N_615,N_4495);
xnor U9051 (N_9051,N_121,N_1670);
nor U9052 (N_9052,N_2794,N_2531);
nand U9053 (N_9053,N_2414,N_104);
xor U9054 (N_9054,N_4435,N_680);
xor U9055 (N_9055,N_970,N_1652);
or U9056 (N_9056,N_936,N_1981);
xor U9057 (N_9057,N_304,N_4932);
nand U9058 (N_9058,N_1975,N_231);
nand U9059 (N_9059,N_2523,N_4392);
nor U9060 (N_9060,N_2328,N_2513);
nand U9061 (N_9061,N_4817,N_2581);
xnor U9062 (N_9062,N_2393,N_2178);
nand U9063 (N_9063,N_4671,N_2342);
nor U9064 (N_9064,N_1322,N_3945);
nand U9065 (N_9065,N_4331,N_1114);
nor U9066 (N_9066,N_1845,N_136);
xor U9067 (N_9067,N_6,N_2135);
or U9068 (N_9068,N_4753,N_4370);
and U9069 (N_9069,N_1482,N_3026);
nor U9070 (N_9070,N_919,N_3691);
nor U9071 (N_9071,N_129,N_810);
and U9072 (N_9072,N_4788,N_1159);
nor U9073 (N_9073,N_2509,N_353);
nand U9074 (N_9074,N_127,N_625);
and U9075 (N_9075,N_2457,N_3568);
nor U9076 (N_9076,N_1281,N_1950);
or U9077 (N_9077,N_1249,N_1957);
or U9078 (N_9078,N_4436,N_2193);
or U9079 (N_9079,N_3408,N_2886);
nand U9080 (N_9080,N_2584,N_4892);
nor U9081 (N_9081,N_2843,N_3509);
nor U9082 (N_9082,N_2842,N_2402);
and U9083 (N_9083,N_2782,N_798);
xnor U9084 (N_9084,N_4441,N_1261);
nor U9085 (N_9085,N_4977,N_3984);
nand U9086 (N_9086,N_3878,N_2343);
and U9087 (N_9087,N_344,N_682);
nand U9088 (N_9088,N_2696,N_4515);
or U9089 (N_9089,N_3118,N_4880);
nand U9090 (N_9090,N_3340,N_1777);
nand U9091 (N_9091,N_2172,N_4025);
xor U9092 (N_9092,N_2962,N_509);
and U9093 (N_9093,N_3185,N_4695);
nor U9094 (N_9094,N_596,N_2885);
or U9095 (N_9095,N_4800,N_1511);
nor U9096 (N_9096,N_4019,N_2846);
nand U9097 (N_9097,N_520,N_590);
or U9098 (N_9098,N_4953,N_3270);
nand U9099 (N_9099,N_2139,N_4635);
nor U9100 (N_9100,N_4207,N_966);
nor U9101 (N_9101,N_4047,N_4590);
and U9102 (N_9102,N_3697,N_3110);
nand U9103 (N_9103,N_2176,N_1958);
or U9104 (N_9104,N_2074,N_3127);
and U9105 (N_9105,N_1073,N_2669);
nand U9106 (N_9106,N_220,N_447);
or U9107 (N_9107,N_4376,N_2414);
or U9108 (N_9108,N_502,N_1681);
or U9109 (N_9109,N_865,N_4340);
xor U9110 (N_9110,N_3092,N_3744);
or U9111 (N_9111,N_3514,N_1362);
xor U9112 (N_9112,N_1996,N_1183);
nor U9113 (N_9113,N_1493,N_655);
or U9114 (N_9114,N_3200,N_1715);
nand U9115 (N_9115,N_1809,N_1439);
nor U9116 (N_9116,N_3347,N_4997);
nor U9117 (N_9117,N_2284,N_217);
nor U9118 (N_9118,N_4312,N_4889);
and U9119 (N_9119,N_3201,N_2354);
or U9120 (N_9120,N_2592,N_3145);
nor U9121 (N_9121,N_3881,N_3720);
or U9122 (N_9122,N_4027,N_4072);
and U9123 (N_9123,N_3194,N_452);
and U9124 (N_9124,N_702,N_4346);
xor U9125 (N_9125,N_3668,N_3441);
or U9126 (N_9126,N_181,N_1820);
and U9127 (N_9127,N_2389,N_1547);
xnor U9128 (N_9128,N_4747,N_1598);
nand U9129 (N_9129,N_424,N_4181);
and U9130 (N_9130,N_2394,N_1317);
nand U9131 (N_9131,N_1310,N_425);
or U9132 (N_9132,N_3103,N_3611);
or U9133 (N_9133,N_3117,N_3855);
or U9134 (N_9134,N_1351,N_1278);
nand U9135 (N_9135,N_2994,N_3885);
nor U9136 (N_9136,N_261,N_2616);
xor U9137 (N_9137,N_3450,N_696);
nand U9138 (N_9138,N_1928,N_1176);
nor U9139 (N_9139,N_170,N_2394);
xor U9140 (N_9140,N_2585,N_1172);
nand U9141 (N_9141,N_3251,N_4609);
or U9142 (N_9142,N_4241,N_1484);
and U9143 (N_9143,N_271,N_3216);
xnor U9144 (N_9144,N_3180,N_679);
xor U9145 (N_9145,N_1694,N_4867);
nand U9146 (N_9146,N_1205,N_4123);
nor U9147 (N_9147,N_2814,N_2017);
xnor U9148 (N_9148,N_4479,N_1852);
or U9149 (N_9149,N_230,N_4540);
nor U9150 (N_9150,N_583,N_1439);
or U9151 (N_9151,N_362,N_192);
or U9152 (N_9152,N_1438,N_3214);
or U9153 (N_9153,N_4097,N_2175);
xor U9154 (N_9154,N_3106,N_1236);
xnor U9155 (N_9155,N_4603,N_725);
nor U9156 (N_9156,N_2427,N_1707);
or U9157 (N_9157,N_3664,N_66);
nor U9158 (N_9158,N_1777,N_3321);
nor U9159 (N_9159,N_4987,N_4561);
and U9160 (N_9160,N_3712,N_1634);
xnor U9161 (N_9161,N_3582,N_2457);
nand U9162 (N_9162,N_4926,N_2624);
and U9163 (N_9163,N_4146,N_4247);
nor U9164 (N_9164,N_854,N_3654);
and U9165 (N_9165,N_2309,N_170);
or U9166 (N_9166,N_3824,N_869);
and U9167 (N_9167,N_2827,N_7);
nor U9168 (N_9168,N_766,N_4477);
and U9169 (N_9169,N_2050,N_2872);
xnor U9170 (N_9170,N_4217,N_4703);
xnor U9171 (N_9171,N_1170,N_1484);
xor U9172 (N_9172,N_2460,N_3151);
nor U9173 (N_9173,N_1521,N_84);
nand U9174 (N_9174,N_3711,N_4332);
nand U9175 (N_9175,N_3551,N_1936);
or U9176 (N_9176,N_4822,N_4686);
nor U9177 (N_9177,N_545,N_875);
xnor U9178 (N_9178,N_1834,N_52);
or U9179 (N_9179,N_991,N_3258);
nand U9180 (N_9180,N_4952,N_2758);
nor U9181 (N_9181,N_3199,N_1294);
or U9182 (N_9182,N_3793,N_1954);
xor U9183 (N_9183,N_532,N_371);
nor U9184 (N_9184,N_3492,N_878);
xor U9185 (N_9185,N_4267,N_3375);
and U9186 (N_9186,N_4726,N_4013);
and U9187 (N_9187,N_3392,N_315);
and U9188 (N_9188,N_956,N_2731);
nor U9189 (N_9189,N_683,N_1874);
xnor U9190 (N_9190,N_3887,N_2927);
or U9191 (N_9191,N_4006,N_419);
and U9192 (N_9192,N_4825,N_200);
and U9193 (N_9193,N_620,N_4472);
nor U9194 (N_9194,N_699,N_2969);
or U9195 (N_9195,N_3043,N_2712);
xor U9196 (N_9196,N_956,N_1467);
xnor U9197 (N_9197,N_4024,N_104);
nor U9198 (N_9198,N_3856,N_907);
nor U9199 (N_9199,N_4489,N_19);
nand U9200 (N_9200,N_2558,N_3845);
or U9201 (N_9201,N_2383,N_937);
nand U9202 (N_9202,N_3242,N_1130);
or U9203 (N_9203,N_3556,N_4167);
nand U9204 (N_9204,N_1664,N_3111);
nand U9205 (N_9205,N_1521,N_12);
and U9206 (N_9206,N_4438,N_594);
or U9207 (N_9207,N_953,N_2072);
and U9208 (N_9208,N_3938,N_3834);
xor U9209 (N_9209,N_2855,N_2991);
nand U9210 (N_9210,N_115,N_1808);
and U9211 (N_9211,N_3037,N_529);
nand U9212 (N_9212,N_2133,N_1759);
xnor U9213 (N_9213,N_1337,N_4167);
xor U9214 (N_9214,N_3381,N_425);
and U9215 (N_9215,N_934,N_65);
nand U9216 (N_9216,N_4311,N_306);
xor U9217 (N_9217,N_4611,N_4182);
xnor U9218 (N_9218,N_824,N_2500);
xor U9219 (N_9219,N_297,N_3672);
nand U9220 (N_9220,N_1092,N_2633);
xor U9221 (N_9221,N_2381,N_2781);
and U9222 (N_9222,N_1699,N_1579);
nor U9223 (N_9223,N_4068,N_55);
and U9224 (N_9224,N_1582,N_2089);
xnor U9225 (N_9225,N_2304,N_1473);
and U9226 (N_9226,N_4126,N_951);
nor U9227 (N_9227,N_4254,N_3281);
xnor U9228 (N_9228,N_3540,N_4014);
or U9229 (N_9229,N_4728,N_4571);
and U9230 (N_9230,N_268,N_1136);
and U9231 (N_9231,N_1440,N_4258);
xor U9232 (N_9232,N_2372,N_2182);
nor U9233 (N_9233,N_1666,N_712);
and U9234 (N_9234,N_4600,N_2183);
and U9235 (N_9235,N_4013,N_4990);
nand U9236 (N_9236,N_2646,N_4446);
nor U9237 (N_9237,N_349,N_2651);
nand U9238 (N_9238,N_874,N_3960);
xor U9239 (N_9239,N_1930,N_894);
or U9240 (N_9240,N_3877,N_2576);
nand U9241 (N_9241,N_2681,N_4309);
nand U9242 (N_9242,N_1213,N_542);
nand U9243 (N_9243,N_3436,N_4902);
xnor U9244 (N_9244,N_2648,N_2692);
and U9245 (N_9245,N_1334,N_2401);
or U9246 (N_9246,N_2298,N_2454);
or U9247 (N_9247,N_477,N_3146);
nand U9248 (N_9248,N_1668,N_2829);
nor U9249 (N_9249,N_1263,N_3699);
nor U9250 (N_9250,N_4241,N_86);
nand U9251 (N_9251,N_3168,N_3716);
nand U9252 (N_9252,N_2612,N_2636);
nand U9253 (N_9253,N_3841,N_768);
and U9254 (N_9254,N_3131,N_470);
or U9255 (N_9255,N_1609,N_3317);
and U9256 (N_9256,N_499,N_3341);
or U9257 (N_9257,N_4083,N_4618);
nand U9258 (N_9258,N_1904,N_172);
nand U9259 (N_9259,N_2676,N_3967);
or U9260 (N_9260,N_2996,N_789);
or U9261 (N_9261,N_3446,N_1529);
or U9262 (N_9262,N_3227,N_4749);
and U9263 (N_9263,N_3707,N_194);
or U9264 (N_9264,N_1715,N_2820);
and U9265 (N_9265,N_4488,N_490);
or U9266 (N_9266,N_934,N_2877);
nand U9267 (N_9267,N_3384,N_1575);
or U9268 (N_9268,N_2775,N_1307);
nor U9269 (N_9269,N_441,N_3964);
nor U9270 (N_9270,N_3988,N_2347);
or U9271 (N_9271,N_4260,N_4245);
xor U9272 (N_9272,N_4873,N_1984);
nand U9273 (N_9273,N_4231,N_454);
nor U9274 (N_9274,N_2603,N_2092);
and U9275 (N_9275,N_499,N_3520);
and U9276 (N_9276,N_746,N_225);
nor U9277 (N_9277,N_1734,N_3241);
nand U9278 (N_9278,N_323,N_3943);
nand U9279 (N_9279,N_835,N_766);
or U9280 (N_9280,N_4535,N_2833);
and U9281 (N_9281,N_873,N_3641);
nor U9282 (N_9282,N_4818,N_3581);
nor U9283 (N_9283,N_2285,N_1984);
nand U9284 (N_9284,N_3313,N_1420);
nand U9285 (N_9285,N_1368,N_4800);
and U9286 (N_9286,N_1466,N_2271);
nor U9287 (N_9287,N_1779,N_2782);
nor U9288 (N_9288,N_3804,N_1828);
nand U9289 (N_9289,N_4272,N_4059);
and U9290 (N_9290,N_3205,N_1150);
or U9291 (N_9291,N_1217,N_2812);
and U9292 (N_9292,N_1278,N_4463);
nand U9293 (N_9293,N_4420,N_3019);
nand U9294 (N_9294,N_1214,N_2281);
nand U9295 (N_9295,N_16,N_2649);
or U9296 (N_9296,N_2779,N_1582);
or U9297 (N_9297,N_1127,N_7);
nor U9298 (N_9298,N_3466,N_470);
nor U9299 (N_9299,N_2452,N_3669);
or U9300 (N_9300,N_4071,N_4825);
or U9301 (N_9301,N_1003,N_4039);
nand U9302 (N_9302,N_3217,N_3210);
nor U9303 (N_9303,N_1776,N_4993);
and U9304 (N_9304,N_542,N_4281);
xnor U9305 (N_9305,N_2473,N_457);
and U9306 (N_9306,N_3817,N_2231);
nand U9307 (N_9307,N_879,N_1319);
nor U9308 (N_9308,N_2990,N_2195);
and U9309 (N_9309,N_1218,N_4582);
and U9310 (N_9310,N_1857,N_4041);
nand U9311 (N_9311,N_4536,N_3384);
nor U9312 (N_9312,N_4354,N_1244);
nor U9313 (N_9313,N_4696,N_468);
nand U9314 (N_9314,N_4357,N_4904);
or U9315 (N_9315,N_3769,N_1446);
nand U9316 (N_9316,N_670,N_4901);
nor U9317 (N_9317,N_1330,N_2822);
or U9318 (N_9318,N_4331,N_4873);
or U9319 (N_9319,N_1543,N_3536);
nor U9320 (N_9320,N_1617,N_2795);
nand U9321 (N_9321,N_1741,N_3654);
and U9322 (N_9322,N_3609,N_4215);
nand U9323 (N_9323,N_4989,N_2027);
or U9324 (N_9324,N_3985,N_4318);
xor U9325 (N_9325,N_987,N_1027);
nor U9326 (N_9326,N_4173,N_2390);
nand U9327 (N_9327,N_731,N_2533);
xor U9328 (N_9328,N_882,N_2478);
or U9329 (N_9329,N_3301,N_1766);
xnor U9330 (N_9330,N_1630,N_486);
nor U9331 (N_9331,N_1230,N_3346);
or U9332 (N_9332,N_2861,N_667);
and U9333 (N_9333,N_1109,N_3769);
and U9334 (N_9334,N_2412,N_2400);
xor U9335 (N_9335,N_2635,N_1309);
and U9336 (N_9336,N_198,N_4775);
xor U9337 (N_9337,N_852,N_1372);
xnor U9338 (N_9338,N_3109,N_4234);
nand U9339 (N_9339,N_1173,N_1794);
nand U9340 (N_9340,N_1026,N_2984);
nand U9341 (N_9341,N_3127,N_1548);
xnor U9342 (N_9342,N_162,N_3311);
nor U9343 (N_9343,N_3529,N_4221);
nor U9344 (N_9344,N_1650,N_3133);
nand U9345 (N_9345,N_2662,N_2221);
nor U9346 (N_9346,N_936,N_2287);
or U9347 (N_9347,N_4277,N_1199);
nor U9348 (N_9348,N_4748,N_2681);
nor U9349 (N_9349,N_4122,N_1977);
nor U9350 (N_9350,N_4633,N_3473);
nor U9351 (N_9351,N_856,N_4748);
nor U9352 (N_9352,N_254,N_121);
or U9353 (N_9353,N_2162,N_666);
xnor U9354 (N_9354,N_2502,N_4204);
xor U9355 (N_9355,N_4704,N_495);
nand U9356 (N_9356,N_4542,N_4388);
xnor U9357 (N_9357,N_4798,N_378);
nor U9358 (N_9358,N_2575,N_1989);
nor U9359 (N_9359,N_3768,N_1219);
nor U9360 (N_9360,N_4550,N_1311);
xnor U9361 (N_9361,N_1393,N_2922);
and U9362 (N_9362,N_268,N_3300);
nand U9363 (N_9363,N_2162,N_1517);
nor U9364 (N_9364,N_1950,N_3200);
or U9365 (N_9365,N_3121,N_553);
xor U9366 (N_9366,N_4743,N_1840);
xnor U9367 (N_9367,N_1947,N_1679);
nand U9368 (N_9368,N_1524,N_4719);
or U9369 (N_9369,N_3124,N_390);
nor U9370 (N_9370,N_2131,N_2055);
nand U9371 (N_9371,N_2224,N_2753);
nor U9372 (N_9372,N_2083,N_287);
or U9373 (N_9373,N_1096,N_4291);
and U9374 (N_9374,N_2897,N_142);
or U9375 (N_9375,N_1329,N_4709);
xor U9376 (N_9376,N_1846,N_1764);
and U9377 (N_9377,N_3689,N_1617);
and U9378 (N_9378,N_3406,N_4694);
or U9379 (N_9379,N_1774,N_3747);
and U9380 (N_9380,N_2447,N_2210);
nor U9381 (N_9381,N_188,N_3618);
nand U9382 (N_9382,N_661,N_3956);
nand U9383 (N_9383,N_465,N_1062);
and U9384 (N_9384,N_507,N_777);
xor U9385 (N_9385,N_908,N_1113);
or U9386 (N_9386,N_2797,N_1729);
nor U9387 (N_9387,N_3928,N_2098);
and U9388 (N_9388,N_2818,N_4053);
or U9389 (N_9389,N_4033,N_2125);
nor U9390 (N_9390,N_1393,N_1222);
nand U9391 (N_9391,N_2646,N_1272);
xnor U9392 (N_9392,N_3355,N_646);
nor U9393 (N_9393,N_1478,N_655);
nor U9394 (N_9394,N_1616,N_3885);
and U9395 (N_9395,N_1658,N_3472);
and U9396 (N_9396,N_2611,N_941);
nand U9397 (N_9397,N_4575,N_4074);
nand U9398 (N_9398,N_3239,N_3164);
or U9399 (N_9399,N_1898,N_1390);
and U9400 (N_9400,N_1609,N_3604);
nand U9401 (N_9401,N_1592,N_2463);
xor U9402 (N_9402,N_4840,N_987);
xor U9403 (N_9403,N_3867,N_3034);
nand U9404 (N_9404,N_725,N_366);
nand U9405 (N_9405,N_2805,N_349);
nand U9406 (N_9406,N_2508,N_314);
nor U9407 (N_9407,N_4395,N_2942);
xnor U9408 (N_9408,N_4750,N_4143);
nor U9409 (N_9409,N_3577,N_168);
nor U9410 (N_9410,N_2021,N_3295);
or U9411 (N_9411,N_534,N_1137);
and U9412 (N_9412,N_901,N_4847);
xor U9413 (N_9413,N_3011,N_4677);
nor U9414 (N_9414,N_4631,N_279);
and U9415 (N_9415,N_3998,N_1011);
xnor U9416 (N_9416,N_2184,N_618);
or U9417 (N_9417,N_1593,N_1370);
nor U9418 (N_9418,N_455,N_1315);
or U9419 (N_9419,N_3487,N_4537);
xor U9420 (N_9420,N_2349,N_2419);
xor U9421 (N_9421,N_4275,N_679);
or U9422 (N_9422,N_442,N_118);
nand U9423 (N_9423,N_1075,N_4048);
nand U9424 (N_9424,N_1124,N_1437);
xor U9425 (N_9425,N_4265,N_3976);
or U9426 (N_9426,N_1678,N_3515);
nor U9427 (N_9427,N_573,N_414);
or U9428 (N_9428,N_4476,N_3316);
nand U9429 (N_9429,N_1090,N_240);
xnor U9430 (N_9430,N_1291,N_3655);
or U9431 (N_9431,N_3772,N_112);
xnor U9432 (N_9432,N_3009,N_3040);
or U9433 (N_9433,N_1823,N_3300);
and U9434 (N_9434,N_1948,N_783);
nand U9435 (N_9435,N_2959,N_3866);
nand U9436 (N_9436,N_4812,N_3261);
nand U9437 (N_9437,N_4104,N_3256);
xnor U9438 (N_9438,N_3147,N_2774);
xnor U9439 (N_9439,N_3487,N_847);
and U9440 (N_9440,N_2604,N_1980);
xnor U9441 (N_9441,N_2316,N_2546);
nand U9442 (N_9442,N_2250,N_1198);
or U9443 (N_9443,N_1825,N_4184);
nor U9444 (N_9444,N_4821,N_4071);
nor U9445 (N_9445,N_4458,N_2307);
xnor U9446 (N_9446,N_1784,N_2766);
or U9447 (N_9447,N_1019,N_3538);
xor U9448 (N_9448,N_47,N_399);
or U9449 (N_9449,N_946,N_4566);
or U9450 (N_9450,N_1385,N_2960);
nor U9451 (N_9451,N_608,N_4413);
and U9452 (N_9452,N_2210,N_4645);
and U9453 (N_9453,N_2284,N_1489);
and U9454 (N_9454,N_4688,N_1043);
and U9455 (N_9455,N_907,N_4124);
xor U9456 (N_9456,N_2917,N_2128);
nor U9457 (N_9457,N_4086,N_4900);
and U9458 (N_9458,N_334,N_4917);
and U9459 (N_9459,N_1157,N_1556);
and U9460 (N_9460,N_290,N_3165);
and U9461 (N_9461,N_4103,N_3156);
and U9462 (N_9462,N_2892,N_3551);
xnor U9463 (N_9463,N_27,N_492);
or U9464 (N_9464,N_1781,N_558);
and U9465 (N_9465,N_2093,N_4303);
and U9466 (N_9466,N_4898,N_2282);
xor U9467 (N_9467,N_2821,N_2294);
xnor U9468 (N_9468,N_1379,N_2705);
nand U9469 (N_9469,N_3993,N_2776);
nand U9470 (N_9470,N_3962,N_3491);
nor U9471 (N_9471,N_4747,N_76);
nand U9472 (N_9472,N_2986,N_3821);
nor U9473 (N_9473,N_1620,N_217);
nor U9474 (N_9474,N_3739,N_1341);
nor U9475 (N_9475,N_106,N_4156);
nor U9476 (N_9476,N_1586,N_381);
nand U9477 (N_9477,N_1642,N_4518);
nor U9478 (N_9478,N_2001,N_469);
or U9479 (N_9479,N_3726,N_4260);
and U9480 (N_9480,N_732,N_156);
nand U9481 (N_9481,N_2139,N_4097);
and U9482 (N_9482,N_2052,N_631);
or U9483 (N_9483,N_952,N_1059);
nand U9484 (N_9484,N_2384,N_3539);
xor U9485 (N_9485,N_502,N_2348);
and U9486 (N_9486,N_1608,N_3068);
nand U9487 (N_9487,N_677,N_365);
and U9488 (N_9488,N_4985,N_3965);
nor U9489 (N_9489,N_231,N_3371);
or U9490 (N_9490,N_3521,N_4028);
nand U9491 (N_9491,N_4541,N_2421);
nor U9492 (N_9492,N_2661,N_4764);
nand U9493 (N_9493,N_158,N_690);
or U9494 (N_9494,N_2980,N_4707);
nand U9495 (N_9495,N_2728,N_3695);
xor U9496 (N_9496,N_3466,N_4933);
nor U9497 (N_9497,N_659,N_620);
nor U9498 (N_9498,N_3005,N_3014);
nand U9499 (N_9499,N_4785,N_2688);
nor U9500 (N_9500,N_3582,N_827);
xnor U9501 (N_9501,N_389,N_1796);
xor U9502 (N_9502,N_247,N_1258);
xor U9503 (N_9503,N_2674,N_3888);
and U9504 (N_9504,N_2020,N_1327);
nand U9505 (N_9505,N_4407,N_4608);
nand U9506 (N_9506,N_3463,N_4457);
xor U9507 (N_9507,N_4913,N_3584);
or U9508 (N_9508,N_2483,N_4921);
xor U9509 (N_9509,N_4682,N_1454);
or U9510 (N_9510,N_4693,N_4352);
and U9511 (N_9511,N_1168,N_2794);
nor U9512 (N_9512,N_2916,N_4323);
or U9513 (N_9513,N_555,N_348);
nor U9514 (N_9514,N_2218,N_49);
nand U9515 (N_9515,N_1567,N_2347);
xor U9516 (N_9516,N_4882,N_775);
nor U9517 (N_9517,N_3568,N_781);
or U9518 (N_9518,N_2410,N_841);
and U9519 (N_9519,N_1980,N_1351);
nor U9520 (N_9520,N_1652,N_167);
nand U9521 (N_9521,N_2157,N_874);
or U9522 (N_9522,N_4761,N_4880);
or U9523 (N_9523,N_4424,N_1099);
nand U9524 (N_9524,N_3843,N_3325);
nor U9525 (N_9525,N_4796,N_2660);
xnor U9526 (N_9526,N_2682,N_1557);
nand U9527 (N_9527,N_1968,N_1038);
nand U9528 (N_9528,N_454,N_1625);
nand U9529 (N_9529,N_4371,N_452);
nand U9530 (N_9530,N_2028,N_541);
xor U9531 (N_9531,N_3124,N_869);
xnor U9532 (N_9532,N_3633,N_1342);
and U9533 (N_9533,N_3872,N_181);
and U9534 (N_9534,N_2480,N_2098);
nor U9535 (N_9535,N_2098,N_850);
or U9536 (N_9536,N_4453,N_4911);
nand U9537 (N_9537,N_4342,N_526);
nor U9538 (N_9538,N_4893,N_735);
or U9539 (N_9539,N_3464,N_1824);
nand U9540 (N_9540,N_2364,N_4245);
nand U9541 (N_9541,N_4440,N_3486);
and U9542 (N_9542,N_1715,N_3125);
or U9543 (N_9543,N_3743,N_991);
or U9544 (N_9544,N_1747,N_2299);
xor U9545 (N_9545,N_2684,N_744);
or U9546 (N_9546,N_3226,N_1372);
xor U9547 (N_9547,N_4728,N_4013);
nor U9548 (N_9548,N_4571,N_653);
nand U9549 (N_9549,N_4568,N_3945);
nor U9550 (N_9550,N_2931,N_2748);
and U9551 (N_9551,N_936,N_534);
and U9552 (N_9552,N_1746,N_1143);
xor U9553 (N_9553,N_236,N_3794);
nand U9554 (N_9554,N_864,N_1547);
xnor U9555 (N_9555,N_698,N_658);
xor U9556 (N_9556,N_2935,N_2741);
nand U9557 (N_9557,N_3417,N_1509);
and U9558 (N_9558,N_3455,N_4732);
xnor U9559 (N_9559,N_744,N_1576);
or U9560 (N_9560,N_1987,N_3648);
or U9561 (N_9561,N_2167,N_836);
and U9562 (N_9562,N_2942,N_4501);
and U9563 (N_9563,N_995,N_567);
and U9564 (N_9564,N_416,N_371);
nand U9565 (N_9565,N_68,N_1864);
or U9566 (N_9566,N_2521,N_743);
and U9567 (N_9567,N_3727,N_292);
and U9568 (N_9568,N_3357,N_4133);
and U9569 (N_9569,N_2009,N_2157);
nand U9570 (N_9570,N_1762,N_4238);
or U9571 (N_9571,N_228,N_2976);
nand U9572 (N_9572,N_1393,N_893);
nor U9573 (N_9573,N_1837,N_4666);
or U9574 (N_9574,N_2131,N_3951);
and U9575 (N_9575,N_1344,N_3974);
and U9576 (N_9576,N_2976,N_2061);
and U9577 (N_9577,N_934,N_3280);
nor U9578 (N_9578,N_2620,N_1735);
and U9579 (N_9579,N_2714,N_2040);
and U9580 (N_9580,N_1930,N_4691);
and U9581 (N_9581,N_4725,N_1224);
nor U9582 (N_9582,N_4879,N_1629);
or U9583 (N_9583,N_3190,N_2364);
nor U9584 (N_9584,N_1113,N_407);
nand U9585 (N_9585,N_4780,N_3408);
or U9586 (N_9586,N_3367,N_4339);
and U9587 (N_9587,N_1209,N_3328);
or U9588 (N_9588,N_1210,N_2363);
and U9589 (N_9589,N_3069,N_4897);
nor U9590 (N_9590,N_4517,N_2040);
nor U9591 (N_9591,N_3413,N_1810);
nand U9592 (N_9592,N_1087,N_3863);
nor U9593 (N_9593,N_2788,N_1180);
xor U9594 (N_9594,N_2898,N_2775);
nand U9595 (N_9595,N_4200,N_1964);
and U9596 (N_9596,N_4831,N_34);
and U9597 (N_9597,N_3327,N_942);
and U9598 (N_9598,N_4574,N_2789);
and U9599 (N_9599,N_3892,N_450);
or U9600 (N_9600,N_4965,N_2829);
or U9601 (N_9601,N_3653,N_1999);
or U9602 (N_9602,N_2782,N_2066);
xnor U9603 (N_9603,N_4239,N_1543);
or U9604 (N_9604,N_4036,N_1018);
or U9605 (N_9605,N_1440,N_620);
and U9606 (N_9606,N_1385,N_4435);
and U9607 (N_9607,N_2195,N_4517);
or U9608 (N_9608,N_996,N_3043);
and U9609 (N_9609,N_4047,N_3494);
nand U9610 (N_9610,N_1077,N_3955);
and U9611 (N_9611,N_2370,N_1246);
nor U9612 (N_9612,N_2501,N_3151);
nor U9613 (N_9613,N_2596,N_1936);
nand U9614 (N_9614,N_3948,N_3343);
xor U9615 (N_9615,N_537,N_503);
and U9616 (N_9616,N_3552,N_124);
or U9617 (N_9617,N_776,N_4992);
nor U9618 (N_9618,N_2220,N_474);
nor U9619 (N_9619,N_895,N_3280);
nand U9620 (N_9620,N_2873,N_2607);
nor U9621 (N_9621,N_4716,N_964);
or U9622 (N_9622,N_4092,N_2701);
and U9623 (N_9623,N_1877,N_3904);
or U9624 (N_9624,N_577,N_239);
xnor U9625 (N_9625,N_4886,N_789);
and U9626 (N_9626,N_3158,N_3638);
and U9627 (N_9627,N_242,N_3557);
nand U9628 (N_9628,N_1947,N_794);
nor U9629 (N_9629,N_249,N_2731);
and U9630 (N_9630,N_1759,N_328);
xor U9631 (N_9631,N_2169,N_4350);
or U9632 (N_9632,N_4766,N_1567);
xnor U9633 (N_9633,N_605,N_4928);
or U9634 (N_9634,N_1924,N_852);
xor U9635 (N_9635,N_3469,N_3440);
nand U9636 (N_9636,N_495,N_3159);
nor U9637 (N_9637,N_2072,N_2159);
nor U9638 (N_9638,N_1217,N_1360);
nand U9639 (N_9639,N_871,N_3881);
nand U9640 (N_9640,N_1363,N_4791);
xor U9641 (N_9641,N_2848,N_2392);
or U9642 (N_9642,N_40,N_1228);
and U9643 (N_9643,N_1973,N_98);
nand U9644 (N_9644,N_1584,N_3177);
or U9645 (N_9645,N_2490,N_502);
or U9646 (N_9646,N_3162,N_499);
nand U9647 (N_9647,N_1205,N_3960);
or U9648 (N_9648,N_3496,N_4344);
nor U9649 (N_9649,N_2543,N_1552);
or U9650 (N_9650,N_2844,N_2637);
or U9651 (N_9651,N_1072,N_4062);
or U9652 (N_9652,N_4933,N_3154);
xor U9653 (N_9653,N_4878,N_2085);
and U9654 (N_9654,N_936,N_4527);
and U9655 (N_9655,N_3404,N_84);
or U9656 (N_9656,N_2122,N_4215);
xnor U9657 (N_9657,N_4306,N_446);
or U9658 (N_9658,N_1148,N_494);
and U9659 (N_9659,N_2415,N_2525);
and U9660 (N_9660,N_4034,N_2398);
xnor U9661 (N_9661,N_3173,N_1748);
and U9662 (N_9662,N_3112,N_772);
and U9663 (N_9663,N_1027,N_288);
xnor U9664 (N_9664,N_1412,N_1744);
xor U9665 (N_9665,N_1233,N_1384);
nor U9666 (N_9666,N_96,N_2593);
nand U9667 (N_9667,N_1668,N_593);
nor U9668 (N_9668,N_1164,N_3331);
and U9669 (N_9669,N_4379,N_3292);
xnor U9670 (N_9670,N_1725,N_1522);
nor U9671 (N_9671,N_985,N_3458);
xor U9672 (N_9672,N_792,N_3917);
nor U9673 (N_9673,N_1350,N_769);
xnor U9674 (N_9674,N_2130,N_3149);
and U9675 (N_9675,N_2791,N_2325);
nand U9676 (N_9676,N_459,N_4110);
and U9677 (N_9677,N_2609,N_700);
and U9678 (N_9678,N_953,N_1936);
xor U9679 (N_9679,N_1784,N_2420);
nand U9680 (N_9680,N_2479,N_3436);
nand U9681 (N_9681,N_170,N_3607);
nand U9682 (N_9682,N_139,N_3362);
xnor U9683 (N_9683,N_4936,N_1455);
xnor U9684 (N_9684,N_121,N_1530);
xor U9685 (N_9685,N_1274,N_1844);
nand U9686 (N_9686,N_395,N_4791);
nor U9687 (N_9687,N_667,N_4542);
and U9688 (N_9688,N_1572,N_3912);
and U9689 (N_9689,N_2182,N_1079);
nand U9690 (N_9690,N_101,N_3481);
and U9691 (N_9691,N_2874,N_997);
or U9692 (N_9692,N_2633,N_2707);
nor U9693 (N_9693,N_1572,N_2379);
xor U9694 (N_9694,N_4915,N_3592);
nor U9695 (N_9695,N_841,N_2959);
nor U9696 (N_9696,N_1263,N_1087);
xnor U9697 (N_9697,N_2146,N_1042);
nor U9698 (N_9698,N_2236,N_1513);
or U9699 (N_9699,N_3429,N_1052);
nor U9700 (N_9700,N_3561,N_82);
nand U9701 (N_9701,N_1870,N_479);
nand U9702 (N_9702,N_1347,N_3687);
nor U9703 (N_9703,N_1627,N_4354);
nor U9704 (N_9704,N_820,N_3885);
and U9705 (N_9705,N_1879,N_615);
nor U9706 (N_9706,N_3271,N_483);
nand U9707 (N_9707,N_1272,N_3862);
xnor U9708 (N_9708,N_1581,N_2532);
or U9709 (N_9709,N_531,N_1980);
or U9710 (N_9710,N_2648,N_770);
nor U9711 (N_9711,N_2469,N_1565);
or U9712 (N_9712,N_3288,N_2597);
or U9713 (N_9713,N_2086,N_2570);
and U9714 (N_9714,N_3457,N_1374);
nor U9715 (N_9715,N_995,N_4425);
nor U9716 (N_9716,N_1898,N_4362);
nand U9717 (N_9717,N_4946,N_1309);
and U9718 (N_9718,N_551,N_424);
and U9719 (N_9719,N_880,N_4557);
nand U9720 (N_9720,N_1197,N_613);
and U9721 (N_9721,N_4189,N_3732);
xnor U9722 (N_9722,N_721,N_550);
nand U9723 (N_9723,N_3066,N_2569);
or U9724 (N_9724,N_105,N_2726);
and U9725 (N_9725,N_4503,N_1250);
and U9726 (N_9726,N_2808,N_3369);
nor U9727 (N_9727,N_2739,N_1934);
or U9728 (N_9728,N_2600,N_394);
or U9729 (N_9729,N_1775,N_4690);
or U9730 (N_9730,N_1868,N_359);
or U9731 (N_9731,N_3302,N_242);
nand U9732 (N_9732,N_797,N_3555);
nor U9733 (N_9733,N_4217,N_107);
or U9734 (N_9734,N_4381,N_4347);
or U9735 (N_9735,N_463,N_2093);
nor U9736 (N_9736,N_1008,N_670);
nand U9737 (N_9737,N_568,N_113);
and U9738 (N_9738,N_4883,N_4316);
nand U9739 (N_9739,N_4757,N_2126);
nor U9740 (N_9740,N_2849,N_563);
xor U9741 (N_9741,N_1942,N_3027);
and U9742 (N_9742,N_1043,N_1177);
nand U9743 (N_9743,N_2525,N_3312);
or U9744 (N_9744,N_1022,N_304);
or U9745 (N_9745,N_1976,N_4376);
or U9746 (N_9746,N_1686,N_1817);
nand U9747 (N_9747,N_2987,N_3330);
or U9748 (N_9748,N_3341,N_4716);
and U9749 (N_9749,N_3675,N_2490);
or U9750 (N_9750,N_1138,N_2901);
or U9751 (N_9751,N_2456,N_1573);
nand U9752 (N_9752,N_1218,N_2700);
and U9753 (N_9753,N_1074,N_780);
and U9754 (N_9754,N_4272,N_4208);
nand U9755 (N_9755,N_337,N_3513);
nand U9756 (N_9756,N_3958,N_3122);
nand U9757 (N_9757,N_724,N_72);
and U9758 (N_9758,N_4088,N_1262);
or U9759 (N_9759,N_1312,N_4982);
or U9760 (N_9760,N_3395,N_4292);
or U9761 (N_9761,N_1276,N_3647);
and U9762 (N_9762,N_4394,N_308);
and U9763 (N_9763,N_4854,N_4381);
xnor U9764 (N_9764,N_1852,N_861);
and U9765 (N_9765,N_3189,N_4280);
and U9766 (N_9766,N_3404,N_3254);
nand U9767 (N_9767,N_2560,N_2027);
xor U9768 (N_9768,N_3764,N_3308);
and U9769 (N_9769,N_4168,N_3987);
and U9770 (N_9770,N_3414,N_4623);
xnor U9771 (N_9771,N_2291,N_2116);
or U9772 (N_9772,N_622,N_3982);
xnor U9773 (N_9773,N_2815,N_3697);
or U9774 (N_9774,N_1161,N_2395);
nand U9775 (N_9775,N_2114,N_3000);
xnor U9776 (N_9776,N_93,N_3311);
nand U9777 (N_9777,N_188,N_1463);
nand U9778 (N_9778,N_2365,N_1445);
xor U9779 (N_9779,N_2790,N_3821);
and U9780 (N_9780,N_4569,N_3603);
nor U9781 (N_9781,N_4330,N_1227);
or U9782 (N_9782,N_2946,N_735);
xor U9783 (N_9783,N_4087,N_4124);
xor U9784 (N_9784,N_4085,N_4177);
xnor U9785 (N_9785,N_2523,N_1169);
and U9786 (N_9786,N_1062,N_1221);
xnor U9787 (N_9787,N_4562,N_3043);
and U9788 (N_9788,N_3948,N_569);
nand U9789 (N_9789,N_4468,N_1024);
or U9790 (N_9790,N_3418,N_1604);
nor U9791 (N_9791,N_1822,N_3686);
nor U9792 (N_9792,N_371,N_2553);
and U9793 (N_9793,N_453,N_2289);
and U9794 (N_9794,N_4644,N_3141);
nand U9795 (N_9795,N_672,N_4482);
and U9796 (N_9796,N_762,N_4227);
xor U9797 (N_9797,N_3516,N_301);
xnor U9798 (N_9798,N_557,N_4323);
nor U9799 (N_9799,N_1406,N_1414);
nor U9800 (N_9800,N_4265,N_4029);
or U9801 (N_9801,N_3976,N_3433);
or U9802 (N_9802,N_3932,N_72);
xor U9803 (N_9803,N_4636,N_2515);
and U9804 (N_9804,N_4083,N_4574);
nor U9805 (N_9805,N_2239,N_4897);
or U9806 (N_9806,N_3718,N_661);
nor U9807 (N_9807,N_1474,N_1730);
nor U9808 (N_9808,N_718,N_2067);
xor U9809 (N_9809,N_4092,N_2274);
or U9810 (N_9810,N_4758,N_10);
and U9811 (N_9811,N_904,N_4127);
and U9812 (N_9812,N_3418,N_127);
xnor U9813 (N_9813,N_956,N_545);
and U9814 (N_9814,N_242,N_320);
xor U9815 (N_9815,N_2992,N_23);
or U9816 (N_9816,N_3421,N_1766);
nor U9817 (N_9817,N_2862,N_1374);
nand U9818 (N_9818,N_3229,N_4636);
xor U9819 (N_9819,N_1418,N_3842);
and U9820 (N_9820,N_4765,N_3854);
nor U9821 (N_9821,N_3617,N_772);
or U9822 (N_9822,N_435,N_1582);
xor U9823 (N_9823,N_3520,N_2880);
and U9824 (N_9824,N_4072,N_3828);
and U9825 (N_9825,N_4433,N_2050);
xor U9826 (N_9826,N_4253,N_3933);
nor U9827 (N_9827,N_4335,N_3896);
or U9828 (N_9828,N_915,N_924);
nor U9829 (N_9829,N_1931,N_4859);
and U9830 (N_9830,N_2191,N_470);
nor U9831 (N_9831,N_4321,N_1239);
nor U9832 (N_9832,N_4430,N_3337);
nor U9833 (N_9833,N_755,N_3747);
xnor U9834 (N_9834,N_393,N_4155);
or U9835 (N_9835,N_4569,N_3165);
and U9836 (N_9836,N_4019,N_2999);
nor U9837 (N_9837,N_4200,N_3978);
and U9838 (N_9838,N_1813,N_3220);
nor U9839 (N_9839,N_2097,N_3613);
nor U9840 (N_9840,N_4389,N_3859);
and U9841 (N_9841,N_3279,N_928);
and U9842 (N_9842,N_3199,N_3980);
or U9843 (N_9843,N_3313,N_1389);
nand U9844 (N_9844,N_4719,N_1607);
and U9845 (N_9845,N_4782,N_2537);
xor U9846 (N_9846,N_3581,N_2506);
nand U9847 (N_9847,N_4484,N_3348);
or U9848 (N_9848,N_3343,N_3893);
or U9849 (N_9849,N_4031,N_825);
or U9850 (N_9850,N_1828,N_273);
or U9851 (N_9851,N_2744,N_4487);
nor U9852 (N_9852,N_614,N_3017);
nor U9853 (N_9853,N_4708,N_3264);
nor U9854 (N_9854,N_4777,N_124);
nor U9855 (N_9855,N_534,N_3400);
and U9856 (N_9856,N_3973,N_3232);
and U9857 (N_9857,N_196,N_32);
nor U9858 (N_9858,N_2519,N_2599);
or U9859 (N_9859,N_2596,N_588);
xnor U9860 (N_9860,N_2302,N_2392);
or U9861 (N_9861,N_4970,N_2736);
xnor U9862 (N_9862,N_1045,N_3049);
xor U9863 (N_9863,N_2865,N_2323);
or U9864 (N_9864,N_1679,N_3781);
and U9865 (N_9865,N_4511,N_4390);
or U9866 (N_9866,N_404,N_19);
nand U9867 (N_9867,N_3090,N_829);
and U9868 (N_9868,N_3141,N_613);
xnor U9869 (N_9869,N_164,N_1611);
nor U9870 (N_9870,N_3370,N_2237);
xor U9871 (N_9871,N_2083,N_4682);
nand U9872 (N_9872,N_294,N_1702);
nand U9873 (N_9873,N_3613,N_4352);
and U9874 (N_9874,N_35,N_1979);
xnor U9875 (N_9875,N_2002,N_2556);
nand U9876 (N_9876,N_3601,N_990);
or U9877 (N_9877,N_21,N_550);
nand U9878 (N_9878,N_1347,N_2151);
and U9879 (N_9879,N_4615,N_3311);
and U9880 (N_9880,N_4885,N_679);
nand U9881 (N_9881,N_4761,N_1023);
and U9882 (N_9882,N_4708,N_4333);
nor U9883 (N_9883,N_2664,N_1968);
nand U9884 (N_9884,N_1703,N_4368);
or U9885 (N_9885,N_3819,N_4052);
xnor U9886 (N_9886,N_3756,N_907);
xor U9887 (N_9887,N_178,N_3392);
and U9888 (N_9888,N_779,N_4544);
and U9889 (N_9889,N_2036,N_4100);
nor U9890 (N_9890,N_4539,N_2097);
nand U9891 (N_9891,N_4404,N_4176);
nand U9892 (N_9892,N_4470,N_436);
nand U9893 (N_9893,N_50,N_927);
xor U9894 (N_9894,N_2898,N_4043);
or U9895 (N_9895,N_2703,N_182);
nand U9896 (N_9896,N_3555,N_1056);
nand U9897 (N_9897,N_3754,N_4007);
and U9898 (N_9898,N_3846,N_3707);
xor U9899 (N_9899,N_691,N_1627);
xnor U9900 (N_9900,N_2881,N_346);
or U9901 (N_9901,N_2713,N_3892);
nand U9902 (N_9902,N_3966,N_2745);
xnor U9903 (N_9903,N_2907,N_63);
and U9904 (N_9904,N_1604,N_3868);
nor U9905 (N_9905,N_2879,N_1472);
nor U9906 (N_9906,N_806,N_1259);
nor U9907 (N_9907,N_635,N_3252);
or U9908 (N_9908,N_1440,N_4959);
and U9909 (N_9909,N_2726,N_1873);
or U9910 (N_9910,N_4964,N_4106);
and U9911 (N_9911,N_1524,N_3204);
or U9912 (N_9912,N_70,N_4517);
xor U9913 (N_9913,N_2007,N_2026);
and U9914 (N_9914,N_2659,N_413);
and U9915 (N_9915,N_2449,N_3274);
xor U9916 (N_9916,N_636,N_3987);
or U9917 (N_9917,N_2630,N_1489);
and U9918 (N_9918,N_2891,N_4718);
nand U9919 (N_9919,N_681,N_4119);
nor U9920 (N_9920,N_3670,N_3134);
and U9921 (N_9921,N_1667,N_2366);
or U9922 (N_9922,N_1691,N_4556);
nand U9923 (N_9923,N_2920,N_674);
nor U9924 (N_9924,N_828,N_3851);
xnor U9925 (N_9925,N_893,N_935);
nor U9926 (N_9926,N_1408,N_1877);
or U9927 (N_9927,N_2385,N_4167);
nand U9928 (N_9928,N_1217,N_4420);
nand U9929 (N_9929,N_4684,N_4046);
nor U9930 (N_9930,N_2106,N_4356);
or U9931 (N_9931,N_3093,N_3951);
or U9932 (N_9932,N_2411,N_4658);
nor U9933 (N_9933,N_2699,N_460);
and U9934 (N_9934,N_1201,N_2225);
nor U9935 (N_9935,N_2748,N_4907);
and U9936 (N_9936,N_967,N_2836);
xnor U9937 (N_9937,N_1670,N_400);
and U9938 (N_9938,N_4071,N_3257);
or U9939 (N_9939,N_4951,N_2142);
nand U9940 (N_9940,N_190,N_1899);
or U9941 (N_9941,N_3406,N_3257);
xor U9942 (N_9942,N_4816,N_1674);
or U9943 (N_9943,N_3442,N_4697);
or U9944 (N_9944,N_1821,N_3936);
nor U9945 (N_9945,N_1167,N_152);
xnor U9946 (N_9946,N_4857,N_1220);
nand U9947 (N_9947,N_385,N_839);
or U9948 (N_9948,N_1924,N_2178);
nor U9949 (N_9949,N_682,N_1999);
nand U9950 (N_9950,N_1181,N_2322);
nor U9951 (N_9951,N_1889,N_700);
nor U9952 (N_9952,N_634,N_4961);
nand U9953 (N_9953,N_704,N_1266);
and U9954 (N_9954,N_2697,N_2153);
nor U9955 (N_9955,N_1499,N_707);
nor U9956 (N_9956,N_3838,N_4943);
nor U9957 (N_9957,N_3971,N_1211);
nand U9958 (N_9958,N_4503,N_4682);
and U9959 (N_9959,N_840,N_3902);
nand U9960 (N_9960,N_500,N_3671);
nor U9961 (N_9961,N_1563,N_2506);
or U9962 (N_9962,N_2507,N_3116);
xor U9963 (N_9963,N_1821,N_2095);
nand U9964 (N_9964,N_25,N_1855);
nor U9965 (N_9965,N_424,N_1556);
nand U9966 (N_9966,N_3271,N_2232);
xnor U9967 (N_9967,N_793,N_607);
nand U9968 (N_9968,N_4930,N_755);
xnor U9969 (N_9969,N_1884,N_520);
or U9970 (N_9970,N_2120,N_3104);
xnor U9971 (N_9971,N_1147,N_307);
nand U9972 (N_9972,N_3424,N_4354);
nand U9973 (N_9973,N_4337,N_3506);
nor U9974 (N_9974,N_2809,N_3297);
nand U9975 (N_9975,N_597,N_3941);
nor U9976 (N_9976,N_4650,N_2192);
nand U9977 (N_9977,N_540,N_1796);
xnor U9978 (N_9978,N_601,N_1294);
and U9979 (N_9979,N_2639,N_4686);
and U9980 (N_9980,N_3580,N_384);
xnor U9981 (N_9981,N_4836,N_4206);
nand U9982 (N_9982,N_99,N_2435);
nand U9983 (N_9983,N_2046,N_2082);
and U9984 (N_9984,N_386,N_362);
and U9985 (N_9985,N_3162,N_626);
and U9986 (N_9986,N_3634,N_3421);
nand U9987 (N_9987,N_2434,N_323);
nor U9988 (N_9988,N_867,N_475);
nand U9989 (N_9989,N_2400,N_2081);
and U9990 (N_9990,N_2770,N_3807);
nor U9991 (N_9991,N_734,N_1143);
and U9992 (N_9992,N_2019,N_4954);
xnor U9993 (N_9993,N_3780,N_2005);
or U9994 (N_9994,N_3320,N_836);
nand U9995 (N_9995,N_743,N_1632);
nor U9996 (N_9996,N_3295,N_629);
nand U9997 (N_9997,N_2662,N_3598);
or U9998 (N_9998,N_4190,N_1464);
and U9999 (N_9999,N_3561,N_2896);
nand U10000 (N_10000,N_8217,N_8616);
nand U10001 (N_10001,N_7603,N_7364);
and U10002 (N_10002,N_5380,N_9382);
xor U10003 (N_10003,N_7801,N_8808);
and U10004 (N_10004,N_9335,N_5997);
or U10005 (N_10005,N_8027,N_9683);
nand U10006 (N_10006,N_7892,N_7110);
or U10007 (N_10007,N_9222,N_7326);
xor U10008 (N_10008,N_8642,N_6301);
xnor U10009 (N_10009,N_5472,N_5853);
or U10010 (N_10010,N_5428,N_6872);
or U10011 (N_10011,N_6092,N_5168);
nor U10012 (N_10012,N_8116,N_6284);
xnor U10013 (N_10013,N_6730,N_6689);
or U10014 (N_10014,N_8292,N_9138);
and U10015 (N_10015,N_8493,N_6960);
nor U10016 (N_10016,N_8386,N_8419);
nor U10017 (N_10017,N_8590,N_9206);
or U10018 (N_10018,N_9331,N_9403);
nand U10019 (N_10019,N_8155,N_5872);
nor U10020 (N_10020,N_8737,N_5415);
nand U10021 (N_10021,N_6033,N_5510);
nor U10022 (N_10022,N_5118,N_9044);
or U10023 (N_10023,N_9029,N_9056);
nor U10024 (N_10024,N_6761,N_6610);
and U10025 (N_10025,N_9991,N_9534);
xor U10026 (N_10026,N_6198,N_8170);
and U10027 (N_10027,N_6004,N_5753);
xor U10028 (N_10028,N_8241,N_7732);
or U10029 (N_10029,N_8905,N_7129);
and U10030 (N_10030,N_8569,N_8499);
or U10031 (N_10031,N_7499,N_7709);
nand U10032 (N_10032,N_6785,N_6310);
xor U10033 (N_10033,N_7821,N_7758);
and U10034 (N_10034,N_6046,N_9748);
and U10035 (N_10035,N_7049,N_9633);
xor U10036 (N_10036,N_5754,N_5564);
nor U10037 (N_10037,N_9521,N_5069);
and U10038 (N_10038,N_9375,N_6285);
nor U10039 (N_10039,N_8210,N_8991);
xnor U10040 (N_10040,N_6063,N_8792);
nor U10041 (N_10041,N_7258,N_9645);
xor U10042 (N_10042,N_7459,N_5828);
xor U10043 (N_10043,N_9191,N_8346);
nor U10044 (N_10044,N_7068,N_9390);
or U10045 (N_10045,N_8188,N_7116);
nand U10046 (N_10046,N_9935,N_7570);
and U10047 (N_10047,N_6914,N_7859);
nor U10048 (N_10048,N_9372,N_8803);
or U10049 (N_10049,N_6727,N_5575);
nor U10050 (N_10050,N_8893,N_8353);
or U10051 (N_10051,N_8883,N_9198);
and U10052 (N_10052,N_9089,N_8654);
or U10053 (N_10053,N_8355,N_6748);
nand U10054 (N_10054,N_8186,N_5414);
xnor U10055 (N_10055,N_9102,N_8542);
nand U10056 (N_10056,N_7468,N_9019);
and U10057 (N_10057,N_6172,N_8361);
or U10058 (N_10058,N_8011,N_7080);
or U10059 (N_10059,N_7612,N_7653);
and U10060 (N_10060,N_5271,N_6876);
nor U10061 (N_10061,N_6850,N_6038);
nor U10062 (N_10062,N_6254,N_8403);
or U10063 (N_10063,N_9937,N_9037);
xor U10064 (N_10064,N_9563,N_9949);
xnor U10065 (N_10065,N_8388,N_7019);
and U10066 (N_10066,N_6628,N_7559);
nor U10067 (N_10067,N_9549,N_9632);
nor U10068 (N_10068,N_6188,N_6348);
nor U10069 (N_10069,N_9451,N_7903);
and U10070 (N_10070,N_8421,N_5550);
nand U10071 (N_10071,N_7022,N_5331);
nand U10072 (N_10072,N_8079,N_6179);
and U10073 (N_10073,N_9001,N_8168);
nand U10074 (N_10074,N_8836,N_8026);
nand U10075 (N_10075,N_5714,N_8600);
or U10076 (N_10076,N_6943,N_5540);
nor U10077 (N_10077,N_6679,N_8473);
xnor U10078 (N_10078,N_5335,N_8094);
nand U10079 (N_10079,N_6388,N_8567);
nor U10080 (N_10080,N_8075,N_8523);
xor U10081 (N_10081,N_6885,N_6816);
nand U10082 (N_10082,N_8598,N_6238);
nand U10083 (N_10083,N_6702,N_5966);
xor U10084 (N_10084,N_8985,N_7085);
xor U10085 (N_10085,N_6608,N_9337);
and U10086 (N_10086,N_8483,N_7523);
or U10087 (N_10087,N_7913,N_7145);
nand U10088 (N_10088,N_8220,N_5394);
xnor U10089 (N_10089,N_6669,N_7140);
and U10090 (N_10090,N_6329,N_6533);
nor U10091 (N_10091,N_6859,N_6434);
nor U10092 (N_10092,N_9893,N_5025);
xnor U10093 (N_10093,N_7392,N_5823);
and U10094 (N_10094,N_8855,N_8874);
nor U10095 (N_10095,N_8396,N_7548);
nor U10096 (N_10096,N_7641,N_8973);
or U10097 (N_10097,N_9264,N_6113);
xnor U10098 (N_10098,N_8613,N_7312);
and U10099 (N_10099,N_8514,N_7830);
nor U10100 (N_10100,N_9908,N_6911);
nand U10101 (N_10101,N_5566,N_8670);
nand U10102 (N_10102,N_8195,N_8264);
and U10103 (N_10103,N_7014,N_5653);
nor U10104 (N_10104,N_7565,N_6295);
nand U10105 (N_10105,N_8439,N_7385);
or U10106 (N_10106,N_5584,N_9237);
or U10107 (N_10107,N_8831,N_6508);
or U10108 (N_10108,N_5894,N_7157);
nand U10109 (N_10109,N_7457,N_9396);
nand U10110 (N_10110,N_7622,N_8318);
and U10111 (N_10111,N_7234,N_7490);
xnor U10112 (N_10112,N_5319,N_7374);
xor U10113 (N_10113,N_9021,N_8051);
nor U10114 (N_10114,N_5120,N_6334);
and U10115 (N_10115,N_5981,N_7763);
and U10116 (N_10116,N_6899,N_9139);
nand U10117 (N_10117,N_5212,N_6918);
and U10118 (N_10118,N_8140,N_8326);
nand U10119 (N_10119,N_9421,N_8136);
nor U10120 (N_10120,N_9689,N_5890);
or U10121 (N_10121,N_6481,N_9108);
and U10122 (N_10122,N_5225,N_8588);
and U10123 (N_10123,N_7919,N_9725);
nand U10124 (N_10124,N_9698,N_6041);
and U10125 (N_10125,N_5742,N_7505);
and U10126 (N_10126,N_8409,N_7101);
xnor U10127 (N_10127,N_7964,N_6705);
nor U10128 (N_10128,N_8391,N_9597);
nand U10129 (N_10129,N_9721,N_5778);
and U10130 (N_10130,N_6021,N_6624);
or U10131 (N_10131,N_6897,N_6668);
nand U10132 (N_10132,N_9901,N_6404);
nor U10133 (N_10133,N_5023,N_6527);
and U10134 (N_10134,N_6762,N_5869);
or U10135 (N_10135,N_7632,N_8001);
nor U10136 (N_10136,N_5868,N_5860);
xnor U10137 (N_10137,N_7183,N_9933);
or U10138 (N_10138,N_9463,N_7831);
and U10139 (N_10139,N_9718,N_7848);
and U10140 (N_10140,N_9436,N_6383);
and U10141 (N_10141,N_7788,N_9792);
or U10142 (N_10142,N_8938,N_6747);
xor U10143 (N_10143,N_5016,N_6953);
nor U10144 (N_10144,N_5343,N_8378);
nor U10145 (N_10145,N_8479,N_5052);
nand U10146 (N_10146,N_8680,N_5588);
and U10147 (N_10147,N_7290,N_6273);
xor U10148 (N_10148,N_6260,N_6696);
nand U10149 (N_10149,N_6419,N_7341);
or U10150 (N_10150,N_6180,N_7872);
nand U10151 (N_10151,N_7982,N_5810);
and U10152 (N_10152,N_6455,N_5109);
and U10153 (N_10153,N_8123,N_9464);
xor U10154 (N_10154,N_9603,N_9227);
xnor U10155 (N_10155,N_8202,N_9958);
and U10156 (N_10156,N_8731,N_5787);
xnor U10157 (N_10157,N_7450,N_8695);
xor U10158 (N_10158,N_5799,N_8247);
or U10159 (N_10159,N_9245,N_5925);
or U10160 (N_10160,N_5191,N_9615);
xnor U10161 (N_10161,N_5318,N_7617);
xnor U10162 (N_10162,N_9033,N_8748);
nand U10163 (N_10163,N_5655,N_8989);
or U10164 (N_10164,N_5492,N_9060);
nand U10165 (N_10165,N_7792,N_6479);
nand U10166 (N_10166,N_5582,N_5864);
and U10167 (N_10167,N_8314,N_5100);
nor U10168 (N_10168,N_8535,N_9739);
nor U10169 (N_10169,N_8490,N_7040);
nor U10170 (N_10170,N_9838,N_8945);
and U10171 (N_10171,N_6025,N_7091);
nor U10172 (N_10172,N_6724,N_5526);
nand U10173 (N_10173,N_9201,N_6346);
nor U10174 (N_10174,N_6871,N_8801);
and U10175 (N_10175,N_8611,N_7658);
and U10176 (N_10176,N_5350,N_6516);
nand U10177 (N_10177,N_7182,N_6358);
nand U10178 (N_10178,N_9554,N_7620);
or U10179 (N_10179,N_5610,N_7774);
nor U10180 (N_10180,N_8901,N_6621);
or U10181 (N_10181,N_8484,N_8006);
or U10182 (N_10182,N_6530,N_8764);
nor U10183 (N_10183,N_5638,N_6192);
xnor U10184 (N_10184,N_6631,N_5022);
xor U10185 (N_10185,N_5177,N_5821);
or U10186 (N_10186,N_9644,N_5920);
or U10187 (N_10187,N_9092,N_8253);
nor U10188 (N_10188,N_6903,N_8625);
and U10189 (N_10189,N_7648,N_5438);
nand U10190 (N_10190,N_9607,N_5939);
xor U10191 (N_10191,N_8390,N_5725);
xnor U10192 (N_10192,N_9118,N_9022);
xnor U10193 (N_10193,N_5771,N_6077);
or U10194 (N_10194,N_5577,N_6612);
or U10195 (N_10195,N_5161,N_9915);
and U10196 (N_10196,N_5859,N_6468);
nor U10197 (N_10197,N_6744,N_5098);
xor U10198 (N_10198,N_5258,N_9357);
xnor U10199 (N_10199,N_6096,N_8610);
or U10200 (N_10200,N_8284,N_7460);
xor U10201 (N_10201,N_5284,N_6231);
nor U10202 (N_10202,N_5358,N_6407);
nor U10203 (N_10203,N_5583,N_5163);
and U10204 (N_10204,N_6312,N_6792);
and U10205 (N_10205,N_7568,N_7199);
and U10206 (N_10206,N_5162,N_5111);
and U10207 (N_10207,N_7281,N_9459);
xor U10208 (N_10208,N_7894,N_8961);
or U10209 (N_10209,N_5571,N_7515);
nand U10210 (N_10210,N_5047,N_7125);
xnor U10211 (N_10211,N_5795,N_6952);
nor U10212 (N_10212,N_9197,N_6339);
or U10213 (N_10213,N_6580,N_7655);
or U10214 (N_10214,N_7840,N_5817);
nand U10215 (N_10215,N_7627,N_6200);
or U10216 (N_10216,N_8156,N_8227);
or U10217 (N_10217,N_8516,N_6558);
or U10218 (N_10218,N_5452,N_5707);
nand U10219 (N_10219,N_6684,N_7273);
xnor U10220 (N_10220,N_5112,N_7313);
and U10221 (N_10221,N_8614,N_9616);
and U10222 (N_10222,N_5383,N_7445);
xor U10223 (N_10223,N_5466,N_7733);
nor U10224 (N_10224,N_9565,N_5442);
nor U10225 (N_10225,N_6313,N_8142);
nand U10226 (N_10226,N_9302,N_5024);
nand U10227 (N_10227,N_7728,N_9169);
xor U10228 (N_10228,N_5700,N_5576);
nor U10229 (N_10229,N_5980,N_6995);
nand U10230 (N_10230,N_9242,N_8262);
nor U10231 (N_10231,N_7484,N_6320);
or U10232 (N_10232,N_6556,N_8312);
nand U10233 (N_10233,N_6239,N_6714);
xnor U10234 (N_10234,N_5091,N_5359);
nand U10235 (N_10235,N_8771,N_9345);
nor U10236 (N_10236,N_9086,N_6579);
nor U10237 (N_10237,N_5736,N_9048);
nand U10238 (N_10238,N_8556,N_6999);
and U10239 (N_10239,N_6435,N_6812);
or U10240 (N_10240,N_8508,N_6791);
nor U10241 (N_10241,N_9759,N_9894);
or U10242 (N_10242,N_5996,N_8908);
and U10243 (N_10243,N_6463,N_8054);
and U10244 (N_10244,N_7850,N_8971);
nor U10245 (N_10245,N_5625,N_6121);
nor U10246 (N_10246,N_5231,N_5323);
nand U10247 (N_10247,N_8848,N_6122);
xnor U10248 (N_10248,N_8699,N_9391);
and U10249 (N_10249,N_8328,N_8928);
nor U10250 (N_10250,N_8038,N_6844);
xor U10251 (N_10251,N_6736,N_6665);
xnor U10252 (N_10252,N_8622,N_9555);
nor U10253 (N_10253,N_6917,N_5171);
xnor U10254 (N_10254,N_5842,N_7710);
and U10255 (N_10255,N_7937,N_7084);
nor U10256 (N_10256,N_9047,N_7917);
nor U10257 (N_10257,N_6034,N_7926);
and U10258 (N_10258,N_6293,N_8981);
nor U10259 (N_10259,N_5900,N_5348);
nand U10260 (N_10260,N_8770,N_9000);
and U10261 (N_10261,N_9348,N_6588);
xor U10262 (N_10262,N_6742,N_7286);
nor U10263 (N_10263,N_9113,N_9909);
or U10264 (N_10264,N_6772,N_6920);
nand U10265 (N_10265,N_7093,N_6831);
or U10266 (N_10266,N_9500,N_8251);
and U10267 (N_10267,N_5006,N_8537);
xor U10268 (N_10268,N_8811,N_5322);
nand U10269 (N_10269,N_5826,N_6306);
and U10270 (N_10270,N_5246,N_7456);
xor U10271 (N_10271,N_6986,N_5355);
nand U10272 (N_10272,N_6473,N_8400);
nor U10273 (N_10273,N_7028,N_6466);
nand U10274 (N_10274,N_6622,N_6011);
xor U10275 (N_10275,N_8860,N_7675);
xnor U10276 (N_10276,N_6002,N_7253);
and U10277 (N_10277,N_8739,N_8754);
xor U10278 (N_10278,N_9276,N_9356);
nand U10279 (N_10279,N_7128,N_8609);
or U10280 (N_10280,N_9002,N_6849);
nand U10281 (N_10281,N_9685,N_7378);
xnor U10282 (N_10282,N_7931,N_8448);
nand U10283 (N_10283,N_6130,N_8549);
nand U10284 (N_10284,N_7166,N_8077);
nand U10285 (N_10285,N_8005,N_5743);
and U10286 (N_10286,N_6991,N_7349);
or U10287 (N_10287,N_5895,N_6465);
or U10288 (N_10288,N_7882,N_6270);
or U10289 (N_10289,N_5482,N_6662);
nor U10290 (N_10290,N_9746,N_6476);
nand U10291 (N_10291,N_6417,N_9185);
nand U10292 (N_10292,N_8037,N_6043);
or U10293 (N_10293,N_8198,N_8160);
nand U10294 (N_10294,N_8316,N_5059);
nor U10295 (N_10295,N_8471,N_5767);
nand U10296 (N_10296,N_8718,N_6147);
nand U10297 (N_10297,N_9052,N_5606);
or U10298 (N_10298,N_8012,N_8446);
nor U10299 (N_10299,N_8237,N_8402);
xor U10300 (N_10300,N_8095,N_6883);
nor U10301 (N_10301,N_9091,N_5659);
xnor U10302 (N_10302,N_6427,N_8231);
or U10303 (N_10303,N_5529,N_6868);
nor U10304 (N_10304,N_5568,N_8384);
or U10305 (N_10305,N_7829,N_9524);
and U10306 (N_10306,N_7358,N_9861);
nand U10307 (N_10307,N_7708,N_7910);
nand U10308 (N_10308,N_5065,N_7813);
nand U10309 (N_10309,N_9440,N_7657);
nand U10310 (N_10310,N_8106,N_6601);
nand U10311 (N_10311,N_7350,N_8641);
and U10312 (N_10312,N_6936,N_6687);
xnor U10313 (N_10313,N_7077,N_6402);
nand U10314 (N_10314,N_7549,N_9024);
nor U10315 (N_10315,N_6445,N_9338);
nand U10316 (N_10316,N_5216,N_9109);
or U10317 (N_10317,N_9659,N_6343);
nor U10318 (N_10318,N_8022,N_7000);
or U10319 (N_10319,N_8049,N_9030);
and U10320 (N_10320,N_7087,N_8169);
nand U10321 (N_10321,N_9561,N_8603);
or U10322 (N_10322,N_5850,N_7424);
nand U10323 (N_10323,N_8358,N_5494);
or U10324 (N_10324,N_6549,N_7475);
xor U10325 (N_10325,N_5833,N_7346);
or U10326 (N_10326,N_7473,N_8896);
and U10327 (N_10327,N_9434,N_6474);
nand U10328 (N_10328,N_9730,N_5757);
xor U10329 (N_10329,N_7582,N_7112);
and U10330 (N_10330,N_9919,N_7585);
nor U10331 (N_10331,N_5475,N_7525);
or U10332 (N_10332,N_8548,N_5095);
and U10333 (N_10333,N_9604,N_7644);
or U10334 (N_10334,N_9598,N_5881);
nor U10335 (N_10335,N_6766,N_7115);
or U10336 (N_10336,N_5107,N_8659);
and U10337 (N_10337,N_8302,N_5784);
nand U10338 (N_10338,N_9038,N_5789);
and U10339 (N_10339,N_5104,N_8496);
or U10340 (N_10340,N_6400,N_7833);
nand U10341 (N_10341,N_9758,N_6857);
xor U10342 (N_10342,N_7771,N_8708);
nor U10343 (N_10343,N_5669,N_9535);
and U10344 (N_10344,N_9270,N_8031);
nor U10345 (N_10345,N_9221,N_6663);
nand U10346 (N_10346,N_5619,N_9646);
nor U10347 (N_10347,N_9397,N_5621);
nand U10348 (N_10348,N_5978,N_6385);
or U10349 (N_10349,N_8452,N_7631);
or U10350 (N_10350,N_7225,N_7550);
or U10351 (N_10351,N_7396,N_9722);
nand U10352 (N_10352,N_6589,N_7008);
nor U10353 (N_10353,N_9267,N_9438);
and U10354 (N_10354,N_7185,N_9159);
nand U10355 (N_10355,N_7911,N_8107);
nand U10356 (N_10356,N_6058,N_8263);
and U10357 (N_10357,N_5197,N_7656);
nor U10358 (N_10358,N_7317,N_6478);
nor U10359 (N_10359,N_7397,N_9115);
nor U10360 (N_10360,N_5093,N_6103);
xnor U10361 (N_10361,N_7947,N_9955);
nor U10362 (N_10362,N_9333,N_9569);
and U10363 (N_10363,N_5124,N_7520);
nor U10364 (N_10364,N_8466,N_7573);
and U10365 (N_10365,N_5390,N_5697);
or U10366 (N_10366,N_8181,N_7030);
xnor U10367 (N_10367,N_5226,N_6080);
nor U10368 (N_10368,N_9114,N_6015);
or U10369 (N_10369,N_5307,N_7496);
or U10370 (N_10370,N_9230,N_8476);
nor U10371 (N_10371,N_5788,N_5051);
nor U10372 (N_10372,N_7155,N_8257);
and U10373 (N_10373,N_5422,N_5352);
nand U10374 (N_10374,N_8374,N_7767);
and U10375 (N_10375,N_5275,N_9978);
and U10376 (N_10376,N_6643,N_7070);
or U10377 (N_10377,N_9518,N_9810);
or U10378 (N_10378,N_8325,N_9970);
or U10379 (N_10379,N_8447,N_6023);
nand U10380 (N_10380,N_8392,N_9875);
xnor U10381 (N_10381,N_9508,N_5224);
nor U10382 (N_10382,N_6032,N_5173);
nand U10383 (N_10383,N_5281,N_9619);
and U10384 (N_10384,N_6839,N_8940);
and U10385 (N_10385,N_7310,N_6173);
and U10386 (N_10386,N_7347,N_6101);
nor U10387 (N_10387,N_6138,N_7980);
nor U10388 (N_10388,N_9658,N_6351);
or U10389 (N_10389,N_5096,N_7900);
and U10390 (N_10390,N_5892,N_6505);
or U10391 (N_10391,N_8131,N_6996);
nand U10392 (N_10392,N_7752,N_6604);
and U10393 (N_10393,N_9031,N_6226);
nor U10394 (N_10394,N_5076,N_9707);
or U10395 (N_10395,N_8068,N_9233);
nor U10396 (N_10396,N_6279,N_8086);
xnor U10397 (N_10397,N_9192,N_9073);
nand U10398 (N_10398,N_5694,N_6596);
nand U10399 (N_10399,N_7386,N_9918);
xnor U10400 (N_10400,N_5663,N_9769);
or U10401 (N_10401,N_8458,N_6185);
nor U10402 (N_10402,N_5070,N_5728);
nor U10403 (N_10403,N_6376,N_7990);
nand U10404 (N_10404,N_5308,N_9956);
xor U10405 (N_10405,N_9425,N_6178);
nor U10406 (N_10406,N_6289,N_5201);
and U10407 (N_10407,N_6919,N_6828);
xnor U10408 (N_10408,N_8321,N_6443);
nor U10409 (N_10409,N_6683,N_8772);
nor U10410 (N_10410,N_8778,N_9078);
nor U10411 (N_10411,N_5372,N_9843);
nor U10412 (N_10412,N_5408,N_6503);
or U10413 (N_10413,N_5692,N_5989);
nand U10414 (N_10414,N_8595,N_8551);
nand U10415 (N_10415,N_5971,N_6983);
or U10416 (N_10416,N_9187,N_7934);
or U10417 (N_10417,N_9349,N_8522);
nor U10418 (N_10418,N_7177,N_9367);
and U10419 (N_10419,N_8847,N_9116);
xnor U10420 (N_10420,N_6595,N_8952);
nor U10421 (N_10421,N_9503,N_7353);
nand U10422 (N_10422,N_9300,N_6674);
nand U10423 (N_10423,N_9015,N_7883);
or U10424 (N_10424,N_8035,N_5974);
or U10425 (N_10425,N_6545,N_5458);
xnor U10426 (N_10426,N_9481,N_9207);
nor U10427 (N_10427,N_6644,N_5252);
and U10428 (N_10428,N_9827,N_8477);
nor U10429 (N_10429,N_7005,N_8254);
or U10430 (N_10430,N_9097,N_6606);
nor U10431 (N_10431,N_9401,N_7669);
or U10432 (N_10432,N_6902,N_7092);
nand U10433 (N_10433,N_7257,N_7994);
and U10434 (N_10434,N_9283,N_7427);
and U10435 (N_10435,N_9776,N_5249);
and U10436 (N_10436,N_8041,N_6672);
or U10437 (N_10437,N_8039,N_8763);
nand U10438 (N_10438,N_8486,N_7437);
nand U10439 (N_10439,N_6378,N_8716);
and U10440 (N_10440,N_6322,N_5569);
nand U10441 (N_10441,N_8222,N_7944);
or U10442 (N_10442,N_8871,N_9393);
xnor U10443 (N_10443,N_6555,N_8751);
nand U10444 (N_10444,N_7105,N_9208);
and U10445 (N_10445,N_8583,N_9556);
and U10446 (N_10446,N_8761,N_6379);
or U10447 (N_10447,N_5046,N_9032);
nor U10448 (N_10448,N_6548,N_6682);
nor U10449 (N_10449,N_6864,N_8701);
and U10450 (N_10450,N_7551,N_5237);
xnor U10451 (N_10451,N_7516,N_5815);
and U10452 (N_10452,N_7552,N_9831);
or U10453 (N_10453,N_5469,N_5623);
nand U10454 (N_10454,N_8283,N_8621);
and U10455 (N_10455,N_6728,N_8118);
and U10456 (N_10456,N_8504,N_6887);
xor U10457 (N_10457,N_5690,N_8943);
xnor U10458 (N_10458,N_9514,N_8620);
or U10459 (N_10459,N_6553,N_6277);
or U10460 (N_10460,N_6879,N_6475);
or U10461 (N_10461,N_9580,N_8669);
xnor U10462 (N_10462,N_7635,N_8752);
nand U10463 (N_10463,N_9336,N_5726);
nand U10464 (N_10464,N_9419,N_9279);
or U10465 (N_10465,N_7731,N_6967);
or U10466 (N_10466,N_7270,N_8280);
or U10467 (N_10467,N_5506,N_8167);
or U10468 (N_10468,N_8462,N_5885);
nor U10469 (N_10469,N_9347,N_7958);
nand U10470 (N_10470,N_8032,N_9317);
nor U10471 (N_10471,N_5213,N_6733);
nand U10472 (N_10472,N_6135,N_5614);
or U10473 (N_10473,N_9506,N_5248);
nand U10474 (N_10474,N_7628,N_6982);
nand U10475 (N_10475,N_7416,N_9315);
nor U10476 (N_10476,N_9117,N_6532);
or U10477 (N_10477,N_6651,N_7454);
xnor U10478 (N_10478,N_8468,N_5187);
and U10479 (N_10479,N_9647,N_6177);
nor U10480 (N_10480,N_6607,N_7480);
or U10481 (N_10481,N_5689,N_9594);
or U10482 (N_10482,N_7064,N_5915);
nor U10483 (N_10483,N_8078,N_8015);
nand U10484 (N_10484,N_8673,N_6423);
nand U10485 (N_10485,N_7509,N_5516);
or U10486 (N_10486,N_9483,N_6645);
or U10487 (N_10487,N_9273,N_7887);
xnor U10488 (N_10488,N_8933,N_7806);
and U10489 (N_10489,N_7884,N_9751);
xor U10490 (N_10490,N_6467,N_8436);
xnor U10491 (N_10491,N_5055,N_7413);
and U10492 (N_10492,N_8105,N_9543);
and U10493 (N_10493,N_9388,N_7869);
xor U10494 (N_10494,N_7432,N_8788);
and U10495 (N_10495,N_8019,N_7609);
xnor U10496 (N_10496,N_9545,N_8776);
or U10497 (N_10497,N_8921,N_6786);
xnor U10498 (N_10498,N_9064,N_6462);
xor U10499 (N_10499,N_8794,N_9959);
nor U10500 (N_10500,N_8806,N_7151);
nand U10501 (N_10501,N_9406,N_9496);
xnor U10502 (N_10502,N_6700,N_7053);
nor U10503 (N_10503,N_5312,N_7595);
nand U10504 (N_10504,N_6323,N_9814);
and U10505 (N_10505,N_5205,N_9794);
or U10506 (N_10506,N_8780,N_9342);
and U10507 (N_10507,N_8747,N_5934);
and U10508 (N_10508,N_6894,N_8014);
nor U10509 (N_10509,N_9701,N_9035);
nand U10510 (N_10510,N_5706,N_9682);
nand U10511 (N_10511,N_5727,N_6056);
xnor U10512 (N_10512,N_8667,N_7066);
nand U10513 (N_10513,N_8927,N_5648);
and U10514 (N_10514,N_5672,N_9014);
nand U10515 (N_10515,N_7393,N_7010);
and U10516 (N_10516,N_6477,N_7498);
and U10517 (N_10517,N_8988,N_7204);
nand U10518 (N_10518,N_5528,N_8098);
or U10519 (N_10519,N_7915,N_8249);
xnor U10520 (N_10520,N_7905,N_6031);
xor U10521 (N_10521,N_6493,N_9681);
nand U10522 (N_10522,N_9850,N_5115);
nand U10523 (N_10523,N_8376,N_6124);
and U10524 (N_10524,N_6948,N_5497);
xor U10525 (N_10525,N_5518,N_9921);
nand U10526 (N_10526,N_9770,N_9103);
nor U10527 (N_10527,N_8686,N_5813);
or U10528 (N_10528,N_7012,N_7984);
nand U10529 (N_10529,N_7345,N_7287);
nand U10530 (N_10530,N_6721,N_8879);
or U10531 (N_10531,N_9250,N_9643);
or U10532 (N_10532,N_5141,N_6258);
and U10533 (N_10533,N_5188,N_6325);
nand U10534 (N_10534,N_5607,N_6502);
nor U10535 (N_10535,N_9126,N_6290);
nand U10536 (N_10536,N_8568,N_9589);
nand U10537 (N_10537,N_5878,N_5734);
or U10538 (N_10538,N_7334,N_6384);
and U10539 (N_10539,N_6895,N_6804);
or U10540 (N_10540,N_5298,N_6341);
xnor U10541 (N_10541,N_6264,N_5834);
xor U10542 (N_10542,N_6637,N_8274);
nor U10543 (N_10543,N_8862,N_9839);
xor U10544 (N_10544,N_8668,N_5473);
xnor U10545 (N_10545,N_7176,N_7781);
nor U10546 (N_10546,N_9447,N_8063);
and U10547 (N_10547,N_6541,N_7362);
or U10548 (N_10548,N_8513,N_7291);
and U10549 (N_10549,N_5914,N_5591);
and U10550 (N_10550,N_5746,N_8810);
and U10551 (N_10551,N_7328,N_5053);
xnor U10552 (N_10552,N_8852,N_9480);
and U10553 (N_10553,N_5884,N_5852);
or U10554 (N_10554,N_8197,N_8919);
nand U10555 (N_10555,N_7095,N_6382);
or U10556 (N_10556,N_8868,N_9025);
or U10557 (N_10557,N_8872,N_9194);
and U10558 (N_10558,N_7034,N_6158);
and U10559 (N_10559,N_5399,N_8999);
nor U10560 (N_10560,N_7581,N_8873);
and U10561 (N_10561,N_6878,N_6051);
or U10562 (N_10562,N_8213,N_8684);
and U10563 (N_10563,N_6935,N_5967);
nor U10564 (N_10564,N_7102,N_8219);
xnor U10565 (N_10565,N_6245,N_5656);
or U10566 (N_10566,N_8067,N_9023);
or U10567 (N_10567,N_6927,N_7662);
nand U10568 (N_10568,N_7680,N_8722);
and U10569 (N_10569,N_6756,N_9719);
nor U10570 (N_10570,N_5402,N_6515);
nand U10571 (N_10571,N_7210,N_9997);
nor U10572 (N_10572,N_8141,N_6286);
and U10573 (N_10573,N_5036,N_9835);
and U10574 (N_10574,N_8646,N_6528);
xnor U10575 (N_10575,N_6184,N_6069);
nand U10576 (N_10576,N_6019,N_5968);
or U10577 (N_10577,N_9179,N_8200);
nor U10578 (N_10578,N_8530,N_8177);
and U10579 (N_10579,N_7006,N_6016);
and U10580 (N_10580,N_6363,N_6444);
xor U10581 (N_10581,N_9596,N_8464);
xor U10582 (N_10582,N_5627,N_7200);
or U10583 (N_10583,N_7616,N_7222);
and U10584 (N_10584,N_6661,N_5363);
xor U10585 (N_10585,N_9635,N_7546);
xnor U10586 (N_10586,N_7246,N_6678);
and U10587 (N_10587,N_8698,N_8710);
and U10588 (N_10588,N_8745,N_5220);
nand U10589 (N_10589,N_5310,N_5483);
and U10590 (N_10590,N_7280,N_8586);
or U10591 (N_10591,N_7422,N_7805);
xnor U10592 (N_10592,N_7007,N_7073);
xor U10593 (N_10593,N_6636,N_6299);
or U10594 (N_10594,N_7981,N_5520);
xor U10595 (N_10595,N_7299,N_7901);
xnor U10596 (N_10596,N_5969,N_9009);
xnor U10597 (N_10597,N_8162,N_6146);
xnor U10598 (N_10598,N_6576,N_7815);
nor U10599 (N_10599,N_7108,N_5744);
xnor U10600 (N_10600,N_8666,N_7181);
xnor U10601 (N_10601,N_7404,N_8497);
and U10602 (N_10602,N_9146,N_7331);
xor U10603 (N_10603,N_7135,N_5844);
or U10604 (N_10604,N_6106,N_6115);
nand U10605 (N_10605,N_5306,N_8822);
or U10606 (N_10606,N_5956,N_7029);
and U10607 (N_10607,N_9341,N_7238);
nor U10608 (N_10608,N_7970,N_7455);
and U10609 (N_10609,N_7097,N_9974);
nand U10610 (N_10610,N_7998,N_6882);
xor U10611 (N_10611,N_5977,N_8687);
nand U10612 (N_10612,N_9591,N_7205);
or U10613 (N_10613,N_5988,N_8365);
nor U10614 (N_10614,N_5539,N_9472);
or U10615 (N_10615,N_8261,N_5048);
or U10616 (N_10616,N_7065,N_8851);
nand U10617 (N_10617,N_5870,N_6818);
nor U10618 (N_10618,N_9149,N_9100);
nand U10619 (N_10619,N_9906,N_5538);
nor U10620 (N_10620,N_9181,N_7720);
nor U10621 (N_10621,N_9482,N_5955);
or U10622 (N_10622,N_7011,N_7320);
nand U10623 (N_10623,N_5431,N_7555);
xor U10624 (N_10624,N_5077,N_6546);
nand U10625 (N_10625,N_9429,N_9405);
or U10626 (N_10626,N_5175,N_5017);
nand U10627 (N_10627,N_7082,N_5282);
or U10628 (N_10628,N_9200,N_7865);
xnor U10629 (N_10629,N_5179,N_7248);
or U10630 (N_10630,N_5798,N_5209);
xnor U10631 (N_10631,N_8090,N_7486);
or U10632 (N_10632,N_9511,N_8781);
nand U10633 (N_10633,N_8689,N_7173);
xor U10634 (N_10634,N_7757,N_6030);
and U10635 (N_10635,N_5200,N_9274);
and U10636 (N_10636,N_6437,N_7700);
nor U10637 (N_10637,N_8712,N_9319);
xor U10638 (N_10638,N_8036,N_9599);
xnor U10639 (N_10639,N_6573,N_6575);
xor U10640 (N_10640,N_7785,N_9984);
nor U10641 (N_10641,N_6688,N_8470);
xor U10642 (N_10642,N_9148,N_7873);
and U10643 (N_10643,N_5381,N_6012);
and U10644 (N_10644,N_5982,N_9387);
nand U10645 (N_10645,N_5841,N_9531);
xor U10646 (N_10646,N_5244,N_8303);
nand U10647 (N_10647,N_8120,N_7542);
nor U10648 (N_10648,N_7139,N_8114);
nor U10649 (N_10649,N_5961,N_6551);
nand U10650 (N_10650,N_6941,N_7242);
and U10651 (N_10651,N_7079,N_7907);
and U10652 (N_10652,N_5002,N_6392);
or U10653 (N_10653,N_6066,N_7239);
xnor U10654 (N_10654,N_9479,N_5041);
nand U10655 (N_10655,N_9642,N_7369);
and U10656 (N_10656,N_7985,N_5759);
and U10657 (N_10657,N_5429,N_8946);
nand U10658 (N_10658,N_9941,N_6997);
or U10659 (N_10659,N_7993,N_6020);
xor U10660 (N_10660,N_9709,N_9675);
and U10661 (N_10661,N_7466,N_8906);
xnor U10662 (N_10662,N_8649,N_8270);
nor U10663 (N_10663,N_5250,N_8252);
and U10664 (N_10664,N_5369,N_9287);
nor U10665 (N_10665,N_8733,N_5434);
nand U10666 (N_10666,N_6449,N_7111);
xnor U10667 (N_10667,N_6162,N_5802);
or U10668 (N_10668,N_9505,N_8540);
nand U10669 (N_10669,N_6214,N_9487);
or U10670 (N_10670,N_7494,N_5635);
or U10671 (N_10671,N_9147,N_6371);
and U10672 (N_10672,N_7614,N_6886);
nor U10673 (N_10673,N_5457,N_8888);
nand U10674 (N_10674,N_7808,N_7340);
nor U10675 (N_10675,N_5604,N_6869);
xnor U10676 (N_10676,N_7399,N_7948);
and U10677 (N_10677,N_9817,N_9522);
nand U10678 (N_10678,N_9856,N_6625);
and U10679 (N_10679,N_8306,N_9693);
and U10680 (N_10680,N_6068,N_9272);
or U10681 (N_10681,N_5032,N_9929);
and U10682 (N_10682,N_9848,N_8062);
nor U10683 (N_10683,N_7743,N_8313);
and U10684 (N_10684,N_8214,N_6989);
nor U10685 (N_10685,N_7613,N_8445);
and U10686 (N_10686,N_9932,N_9080);
xnor U10687 (N_10687,N_7245,N_9779);
nor U10688 (N_10688,N_7886,N_8997);
nand U10689 (N_10689,N_5855,N_5293);
xnor U10690 (N_10690,N_7724,N_9311);
nand U10691 (N_10691,N_7058,N_6175);
and U10692 (N_10692,N_8338,N_7817);
and U10693 (N_10693,N_9070,N_5292);
nor U10694 (N_10694,N_8147,N_6252);
and U10695 (N_10695,N_7895,N_5962);
nor U10696 (N_10696,N_5068,N_8267);
and U10697 (N_10697,N_7179,N_6813);
xnor U10698 (N_10698,N_9803,N_7564);
and U10699 (N_10699,N_6764,N_8559);
or U10700 (N_10700,N_9788,N_6597);
xnor U10701 (N_10701,N_7928,N_7972);
nor U10702 (N_10702,N_5143,N_9470);
and U10703 (N_10703,N_6901,N_5932);
nand U10704 (N_10704,N_6263,N_5486);
xnor U10705 (N_10705,N_8589,N_8534);
or U10706 (N_10706,N_7143,N_6364);
and U10707 (N_10707,N_6498,N_6483);
xnor U10708 (N_10708,N_7621,N_9813);
or U10709 (N_10709,N_7016,N_8688);
nor U10710 (N_10710,N_9542,N_6815);
or U10711 (N_10711,N_5018,N_5632);
or U10712 (N_10712,N_8350,N_6512);
and U10713 (N_10713,N_9628,N_6970);
and U10714 (N_10714,N_5268,N_5503);
xor U10715 (N_10715,N_6836,N_7443);
or U10716 (N_10716,N_6151,N_6854);
nor U10717 (N_10717,N_5373,N_5170);
nand U10718 (N_10718,N_6972,N_9723);
nor U10719 (N_10719,N_5658,N_6560);
nor U10720 (N_10720,N_7104,N_8009);
or U10721 (N_10721,N_7076,N_8393);
xnor U10722 (N_10722,N_8404,N_6250);
nor U10723 (N_10723,N_5637,N_7321);
xnor U10724 (N_10724,N_7150,N_8711);
or U10725 (N_10725,N_8709,N_5601);
xor U10726 (N_10726,N_9800,N_8135);
xnor U10727 (N_10727,N_6629,N_8582);
xor U10728 (N_10728,N_6397,N_9816);
nor U10729 (N_10729,N_8239,N_9416);
or U10730 (N_10730,N_5764,N_6203);
or U10731 (N_10731,N_8059,N_6617);
xor U10732 (N_10732,N_7197,N_8010);
or U10733 (N_10733,N_5157,N_8139);
and U10734 (N_10734,N_7275,N_5634);
or U10735 (N_10735,N_9055,N_9255);
and U10736 (N_10736,N_6236,N_7987);
xnor U10737 (N_10737,N_5440,N_8287);
xnor U10738 (N_10738,N_6955,N_9043);
nor U10739 (N_10739,N_7544,N_5922);
or U10740 (N_10740,N_5154,N_9783);
nand U10741 (N_10741,N_9428,N_6542);
or U10742 (N_10742,N_6968,N_6490);
xor U10743 (N_10743,N_6054,N_6880);
and U10744 (N_10744,N_5050,N_9716);
or U10745 (N_10745,N_6681,N_8876);
or U10746 (N_10746,N_9152,N_6472);
nand U10747 (N_10747,N_6840,N_9863);
or U10748 (N_10748,N_5341,N_7672);
xor U10749 (N_10749,N_8849,N_8528);
nor U10750 (N_10750,N_8902,N_7149);
or U10751 (N_10751,N_7968,N_7540);
xnor U10752 (N_10752,N_9745,N_5203);
and U10753 (N_10753,N_5297,N_8947);
and U10754 (N_10754,N_6307,N_9051);
xnor U10755 (N_10755,N_9106,N_5590);
nor U10756 (N_10756,N_8992,N_6759);
nor U10757 (N_10757,N_7963,N_7009);
xnor U10758 (N_10758,N_7495,N_7314);
nand U10759 (N_10759,N_9690,N_9677);
nor U10760 (N_10760,N_7417,N_8570);
and U10761 (N_10761,N_5504,N_8894);
or U10762 (N_10762,N_5863,N_7643);
nor U10763 (N_10763,N_5346,N_7579);
xor U10764 (N_10764,N_7419,N_7721);
nor U10765 (N_10765,N_7688,N_7405);
nand U10766 (N_10766,N_5089,N_7164);
nor U10767 (N_10767,N_8545,N_5448);
nand U10768 (N_10768,N_6737,N_7730);
or U10769 (N_10769,N_9366,N_5740);
xnor U10770 (N_10770,N_8550,N_8290);
and U10771 (N_10771,N_6050,N_9402);
and U10772 (N_10772,N_9866,N_7615);
and U10773 (N_10773,N_6915,N_9318);
xor U10774 (N_10774,N_6028,N_5031);
nor U10775 (N_10775,N_7351,N_9802);
xnor U10776 (N_10776,N_5578,N_9217);
nand U10777 (N_10777,N_5413,N_5858);
nor U10778 (N_10778,N_9968,N_8515);
or U10779 (N_10779,N_6554,N_8269);
and U10780 (N_10780,N_5138,N_9520);
and U10781 (N_10781,N_6506,N_8870);
xor U10782 (N_10782,N_9687,N_9686);
nor U10783 (N_10783,N_5896,N_8967);
or U10784 (N_10784,N_7306,N_5303);
xnor U10785 (N_10785,N_9424,N_9174);
or U10786 (N_10786,N_9972,N_8332);
or U10787 (N_10787,N_7524,N_8414);
or U10788 (N_10788,N_7381,N_9202);
nand U10789 (N_10789,N_7090,N_9963);
nor U10790 (N_10790,N_6053,N_9260);
and U10791 (N_10791,N_7663,N_5477);
nand U10792 (N_10792,N_8964,N_7256);
and U10793 (N_10793,N_6639,N_7735);
or U10794 (N_10794,N_6401,N_7786);
xnor U10795 (N_10795,N_7051,N_8560);
nand U10796 (N_10796,N_9290,N_5913);
nor U10797 (N_10797,N_5760,N_6504);
or U10798 (N_10798,N_7156,N_6297);
xnor U10799 (N_10799,N_9062,N_8972);
nand U10800 (N_10800,N_8760,N_8696);
or U10801 (N_10801,N_8637,N_8775);
and U10802 (N_10802,N_9437,N_5573);
and U10803 (N_10803,N_5768,N_7857);
and U10804 (N_10804,N_7539,N_9218);
or U10805 (N_10805,N_8839,N_5598);
nand U10806 (N_10806,N_5384,N_5276);
nor U10807 (N_10807,N_5524,N_6436);
nor U10808 (N_10808,N_9162,N_9477);
nand U10809 (N_10809,N_8243,N_9327);
and U10810 (N_10810,N_8990,N_6934);
xnor U10811 (N_10811,N_5254,N_5898);
nand U10812 (N_10812,N_7803,N_7412);
xnor U10813 (N_10813,N_9008,N_8096);
or U10814 (N_10814,N_6984,N_8797);
xor U10815 (N_10815,N_8624,N_7100);
nor U10816 (N_10816,N_8058,N_8830);
nand U10817 (N_10817,N_8970,N_9744);
or U10818 (N_10818,N_9490,N_5696);
xnor U10819 (N_10819,N_8182,N_6086);
and U10820 (N_10820,N_6585,N_8903);
and U10821 (N_10821,N_6137,N_8787);
and U10822 (N_10822,N_9266,N_7004);
nor U10823 (N_10823,N_7191,N_8364);
nand U10824 (N_10824,N_8480,N_9431);
xnor U10825 (N_10825,N_7604,N_9049);
nor U10826 (N_10826,N_8678,N_8904);
nor U10827 (N_10827,N_9811,N_5270);
nor U10828 (N_10828,N_6768,N_8969);
and U10829 (N_10829,N_9987,N_9475);
nand U10830 (N_10830,N_6183,N_6255);
nand U10831 (N_10831,N_9297,N_5792);
xor U10832 (N_10832,N_8460,N_9889);
nand U10833 (N_10833,N_8240,N_8093);
xor U10834 (N_10834,N_5454,N_9074);
nand U10835 (N_10835,N_7159,N_7694);
and U10836 (N_10836,N_5130,N_6484);
nand U10837 (N_10837,N_8727,N_5984);
nand U10838 (N_10838,N_8861,N_5416);
xor U10839 (N_10839,N_6581,N_9844);
or U10840 (N_10840,N_7611,N_5952);
nand U10841 (N_10841,N_5951,N_6957);
and U10842 (N_10842,N_7701,N_8596);
and U10843 (N_10843,N_6215,N_8679);
nand U10844 (N_10844,N_8209,N_8573);
xor U10845 (N_10845,N_5687,N_6686);
nor U10846 (N_10846,N_9111,N_6593);
and U10847 (N_10847,N_5730,N_6328);
or U10848 (N_10848,N_8260,N_5253);
and U10849 (N_10849,N_7117,N_6359);
or U10850 (N_10850,N_5688,N_8023);
and U10851 (N_10851,N_6753,N_8758);
nand U10852 (N_10852,N_5150,N_5548);
xnor U10853 (N_10853,N_5963,N_9392);
and U10854 (N_10854,N_8394,N_6451);
nand U10855 (N_10855,N_7330,N_7729);
xnor U10856 (N_10856,N_9826,N_5103);
xor U10857 (N_10857,N_9223,N_6003);
nor U10858 (N_10858,N_6300,N_8494);
xnor U10859 (N_10859,N_7168,N_6739);
or U10860 (N_10860,N_5649,N_9296);
and U10861 (N_10861,N_9741,N_6963);
or U10862 (N_10862,N_5545,N_5291);
nand U10863 (N_10863,N_7983,N_8843);
nand U10864 (N_10864,N_6234,N_7446);
nand U10865 (N_10865,N_8721,N_5586);
nor U10866 (N_10866,N_6784,N_9641);
nand U10867 (N_10867,N_9947,N_8743);
and U10868 (N_10868,N_7241,N_6735);
nand U10869 (N_10869,N_8021,N_6430);
xnor U10870 (N_10870,N_8703,N_5579);
nand U10871 (N_10871,N_5904,N_7956);
xor U10872 (N_10872,N_8527,N_6834);
nor U10873 (N_10873,N_5990,N_7832);
xor U10874 (N_10874,N_5459,N_9550);
nor U10875 (N_10875,N_9271,N_7506);
or U10876 (N_10876,N_6653,N_5152);
xor U10877 (N_10877,N_9027,N_8154);
and U10878 (N_10878,N_8518,N_8297);
and U10879 (N_10879,N_7823,N_9781);
nand U10880 (N_10880,N_7131,N_9105);
nor U10881 (N_10881,N_8615,N_5502);
nor U10882 (N_10882,N_9364,N_9457);
and U10883 (N_10883,N_8073,N_7426);
xor U10884 (N_10884,N_5449,N_6763);
nand U10885 (N_10885,N_5819,N_9629);
nor U10886 (N_10886,N_5245,N_7343);
and U10887 (N_10887,N_7629,N_9189);
nand U10888 (N_10888,N_7407,N_8858);
xnor U10889 (N_10889,N_7772,N_9328);
or U10890 (N_10890,N_5557,N_6905);
nor U10891 (N_10891,N_6534,N_9870);
or U10892 (N_10892,N_7751,N_7647);
or U10893 (N_10893,N_6061,N_6110);
or U10894 (N_10894,N_6912,N_8798);
and U10895 (N_10895,N_6893,N_5463);
nand U10896 (N_10896,N_8204,N_6779);
and U10897 (N_10897,N_8648,N_9990);
xnor U10898 (N_10898,N_9849,N_8986);
and U10899 (N_10899,N_5765,N_5661);
xor U10900 (N_10900,N_8587,N_5703);
and U10901 (N_10901,N_7361,N_5876);
xor U10902 (N_10902,N_9881,N_7429);
or U10903 (N_10903,N_6846,N_8461);
and U10904 (N_10904,N_5711,N_8960);
nand U10905 (N_10905,N_5693,N_5593);
and U10906 (N_10906,N_8430,N_7491);
nand U10907 (N_10907,N_6671,N_8604);
xor U10908 (N_10908,N_7278,N_9163);
xnor U10909 (N_10909,N_7103,N_5379);
xor U10910 (N_10910,N_9950,N_7951);
nand U10911 (N_10911,N_7556,N_5756);
xor U10912 (N_10912,N_9704,N_5919);
nor U10913 (N_10913,N_7596,N_9873);
and U10914 (N_10914,N_6738,N_8149);
or U10915 (N_10915,N_8272,N_9244);
nor U10916 (N_10916,N_9806,N_9639);
nand U10917 (N_10917,N_5329,N_6093);
xor U10918 (N_10918,N_6525,N_9636);
xor U10919 (N_10919,N_9195,N_5631);
nor U10920 (N_10920,N_9277,N_8910);
nor U10921 (N_10921,N_6396,N_5370);
and U10922 (N_10922,N_7712,N_8857);
xnor U10923 (N_10923,N_6189,N_6564);
nand U10924 (N_10924,N_5640,N_6219);
or U10925 (N_10925,N_6154,N_6412);
and U10926 (N_10926,N_6489,N_7186);
nor U10927 (N_10927,N_7687,N_5081);
or U10928 (N_10928,N_8632,N_5507);
or U10929 (N_10929,N_5094,N_9942);
xnor U10930 (N_10930,N_7044,N_9379);
xor U10931 (N_10931,N_8539,N_6222);
xor U10932 (N_10932,N_8407,N_8580);
and U10933 (N_10933,N_7284,N_8191);
or U10934 (N_10934,N_7575,N_8211);
and U10935 (N_10935,N_5255,N_8875);
nand U10936 (N_10936,N_8813,N_8046);
or U10937 (N_10937,N_8502,N_5830);
xnor U10938 (N_10938,N_7527,N_8389);
nand U10939 (N_10939,N_7229,N_9312);
nor U10940 (N_10940,N_7828,N_7677);
xor U10941 (N_10941,N_6278,N_6613);
nand U10942 (N_10942,N_5476,N_6207);
and U10943 (N_10943,N_6165,N_9020);
nor U10944 (N_10944,N_9780,N_9934);
and U10945 (N_10945,N_9453,N_6827);
and U10946 (N_10946,N_9801,N_9046);
and U10947 (N_10947,N_6916,N_9003);
or U10948 (N_10948,N_5102,N_5159);
xor U10949 (N_10949,N_8412,N_5994);
nand U10950 (N_10950,N_6079,N_9188);
and U10951 (N_10951,N_7639,N_6979);
and U10952 (N_10952,N_5537,N_5877);
and U10953 (N_10953,N_9911,N_6125);
or U10954 (N_10954,N_8658,N_6667);
or U10955 (N_10955,N_8623,N_6452);
nor U10956 (N_10956,N_7950,N_7899);
and U10957 (N_10957,N_6822,N_7220);
or U10958 (N_10958,N_9740,N_7274);
xnor U10959 (N_10959,N_6432,N_6676);
or U10960 (N_10960,N_6420,N_5704);
nor U10961 (N_10961,N_6355,N_9674);
nand U10962 (N_10962,N_8456,N_8235);
or U10963 (N_10963,N_8296,N_5534);
xnor U10964 (N_10964,N_5950,N_9167);
nand U10965 (N_10965,N_7122,N_6387);
nand U10966 (N_10966,N_7746,N_5949);
and U10967 (N_10967,N_8100,N_6108);
nand U10968 (N_10968,N_5733,N_8520);
nand U10969 (N_10969,N_8060,N_8348);
nand U10970 (N_10970,N_5460,N_5194);
and U10971 (N_10971,N_6777,N_5985);
and U10972 (N_10972,N_6283,N_5015);
xnor U10973 (N_10973,N_8702,N_7705);
nand U10974 (N_10974,N_6374,N_5556);
or U10975 (N_10975,N_9468,N_6029);
and U10976 (N_10976,N_6361,N_9624);
and U10977 (N_10977,N_6375,N_9282);
or U10978 (N_10978,N_8482,N_8594);
or U10979 (N_10979,N_6480,N_9582);
nand U10980 (N_10980,N_9867,N_8137);
and U10981 (N_10981,N_9767,N_8322);
nor U10982 (N_10982,N_5602,N_6987);
nand U10983 (N_10983,N_9606,N_6168);
nand U10984 (N_10984,N_7942,N_7927);
xnor U10985 (N_10985,N_6408,N_7787);
and U10986 (N_10986,N_9757,N_8356);
or U10987 (N_10987,N_7762,N_8951);
nand U10988 (N_10988,N_7912,N_6760);
or U10989 (N_10989,N_9966,N_6620);
and U10990 (N_10990,N_9845,N_8431);
nand U10991 (N_10991,N_8882,N_6119);
nor U10992 (N_10992,N_7973,N_9491);
and U10993 (N_10993,N_5455,N_5603);
xnor U10994 (N_10994,N_8102,N_6335);
nor U10995 (N_10995,N_9670,N_5780);
nor U10996 (N_10996,N_9137,N_9989);
nor U10997 (N_10997,N_6713,N_9666);
and U10998 (N_10998,N_8028,N_7718);
and U10999 (N_10999,N_9065,N_7736);
nor U11000 (N_11000,N_5480,N_6406);
or U11001 (N_11001,N_9011,N_6896);
or U11002 (N_11002,N_8838,N_6482);
and U11003 (N_11003,N_6819,N_5713);
xnor U11004 (N_11004,N_5565,N_7213);
nand U11005 (N_11005,N_9836,N_7794);
nor U11006 (N_11006,N_9236,N_6609);
nand U11007 (N_11007,N_6835,N_6460);
nor U11008 (N_11008,N_5643,N_5866);
xnor U11009 (N_11009,N_8704,N_5596);
or U11010 (N_11010,N_5465,N_9777);
nor U11011 (N_11011,N_9351,N_9143);
nand U11012 (N_11012,N_5468,N_5269);
and U11013 (N_11013,N_6007,N_8948);
and U11014 (N_11014,N_5389,N_7272);
nand U11015 (N_11015,N_7510,N_8127);
nand U11016 (N_11016,N_5748,N_8179);
xor U11017 (N_11017,N_9155,N_6228);
nand U11018 (N_11018,N_9763,N_5847);
or U11019 (N_11019,N_9381,N_5822);
xnor U11020 (N_11020,N_5835,N_7537);
xnor U11021 (N_11021,N_8725,N_8834);
or U11022 (N_11022,N_8956,N_9680);
xor U11023 (N_11023,N_5060,N_9072);
or U11024 (N_11024,N_6347,N_7295);
and U11025 (N_11025,N_8259,N_9868);
or U11026 (N_11026,N_5645,N_6640);
nor U11027 (N_11027,N_7974,N_9446);
or U11028 (N_11028,N_5699,N_8828);
xnor U11029 (N_11029,N_7382,N_6457);
and U11030 (N_11030,N_9940,N_6422);
or U11031 (N_11031,N_8526,N_8911);
nand U11032 (N_11032,N_7588,N_8138);
nand U11033 (N_11033,N_8438,N_7939);
nor U11034 (N_11034,N_9577,N_6531);
or U11035 (N_11035,N_8824,N_9804);
xnor U11036 (N_11036,N_5636,N_7837);
or U11037 (N_11037,N_9361,N_8399);
nor U11038 (N_11038,N_5247,N_9983);
xor U11039 (N_11039,N_5338,N_7760);
nand U11040 (N_11040,N_9782,N_9631);
and U11041 (N_11041,N_6666,N_9141);
nand U11042 (N_11042,N_9215,N_7336);
and U11043 (N_11043,N_9085,N_8311);
or U11044 (N_11044,N_5902,N_5236);
and U11045 (N_11045,N_5600,N_7933);
or U11046 (N_11046,N_9498,N_6959);
or U11047 (N_11047,N_5122,N_8744);
and U11048 (N_11048,N_5609,N_6507);
or U11049 (N_11049,N_6418,N_7262);
nand U11050 (N_11050,N_9574,N_8738);
xor U11051 (N_11051,N_6123,N_8941);
nand U11052 (N_11052,N_5407,N_7414);
or U11053 (N_11053,N_8519,N_6626);
nor U11054 (N_11054,N_5228,N_8226);
and U11055 (N_11055,N_7504,N_9013);
nor U11056 (N_11056,N_6036,N_5317);
nor U11057 (N_11057,N_7292,N_6209);
xor U11058 (N_11058,N_9652,N_7988);
xnor U11059 (N_11059,N_7690,N_7660);
or U11060 (N_11060,N_7532,N_8427);
or U11061 (N_11061,N_9442,N_7161);
xor U11062 (N_11062,N_7906,N_7188);
nand U11063 (N_11063,N_6105,N_6829);
xnor U11064 (N_11064,N_7976,N_8366);
nor U11065 (N_11065,N_9786,N_6583);
or U11066 (N_11066,N_9213,N_9088);
and U11067 (N_11067,N_9787,N_8503);
nor U11068 (N_11068,N_7914,N_9203);
xor U11069 (N_11069,N_7793,N_6909);
xor U11070 (N_11070,N_6372,N_9307);
nor U11071 (N_11071,N_9158,N_9036);
and U11072 (N_11072,N_8411,N_9637);
xor U11073 (N_11073,N_8546,N_9957);
nor U11074 (N_11074,N_6201,N_7841);
and U11075 (N_11075,N_7890,N_8925);
nand U11076 (N_11076,N_6469,N_5295);
and U11077 (N_11077,N_8337,N_8053);
and U11078 (N_11078,N_8993,N_7144);
xnor U11079 (N_11079,N_7583,N_7541);
or U11080 (N_11080,N_8432,N_6190);
xnor U11081 (N_11081,N_6240,N_5973);
or U11082 (N_11082,N_9365,N_7485);
or U11083 (N_11083,N_5263,N_7301);
xnor U11084 (N_11084,N_8726,N_7052);
nor U11085 (N_11085,N_6928,N_5144);
or U11086 (N_11086,N_8605,N_6977);
and U11087 (N_11087,N_7580,N_5646);
or U11088 (N_11088,N_6570,N_5337);
xor U11089 (N_11089,N_8998,N_9795);
nand U11090 (N_11090,N_7789,N_7236);
nand U11091 (N_11091,N_9404,N_7081);
or U11092 (N_11092,N_7363,N_7719);
nand U11093 (N_11093,N_8880,N_8184);
xor U11094 (N_11094,N_6232,N_6089);
nand U11095 (N_11095,N_5916,N_8429);
or U11096 (N_11096,N_7046,N_7659);
and U11097 (N_11097,N_6969,N_9898);
or U11098 (N_11098,N_9819,N_8024);
nand U11099 (N_11099,N_5960,N_5718);
and U11100 (N_11100,N_6715,N_6535);
and U11101 (N_11101,N_7431,N_8467);
nand U11102 (N_11102,N_7289,N_6094);
nor U11103 (N_11103,N_7896,N_6447);
nand U11104 (N_11104,N_9492,N_5239);
nor U11105 (N_11105,N_5533,N_5195);
and U11106 (N_11106,N_7447,N_8444);
nand U11107 (N_11107,N_5328,N_8317);
or U11108 (N_11108,N_6971,N_8074);
xnor U11109 (N_11109,N_8405,N_7838);
and U11110 (N_11110,N_6453,N_5814);
nor U11111 (N_11111,N_6373,N_9995);
nor U11112 (N_11112,N_5049,N_8823);
xnor U11113 (N_11113,N_7261,N_7214);
nand U11114 (N_11114,N_7325,N_7493);
or U11115 (N_11115,N_8201,N_6357);
and U11116 (N_11116,N_9252,N_6803);
or U11117 (N_11117,N_5921,N_6000);
and U11118 (N_11118,N_9509,N_5033);
and U11119 (N_11119,N_5617,N_9568);
and U11120 (N_11120,N_5652,N_6230);
and U11121 (N_11121,N_6217,N_9299);
nand U11122 (N_11122,N_8478,N_8357);
nand U11123 (N_11123,N_9454,N_7768);
or U11124 (N_11124,N_7202,N_8398);
and U11125 (N_11125,N_6981,N_6774);
nand U11126 (N_11126,N_9410,N_9449);
and U11127 (N_11127,N_8750,N_9229);
nor U11128 (N_11128,N_8779,N_9818);
nand U11129 (N_11129,N_7265,N_8640);
or U11130 (N_11130,N_5701,N_9473);
nand U11131 (N_11131,N_9981,N_5393);
xor U11132 (N_11132,N_5044,N_9075);
xor U11133 (N_11133,N_7698,N_9828);
xnor U11134 (N_11134,N_9882,N_8173);
xor U11135 (N_11135,N_9517,N_9502);
nor U11136 (N_11136,N_8635,N_6039);
nor U11137 (N_11137,N_8936,N_6590);
xnor U11138 (N_11138,N_9292,N_9812);
xnor U11139 (N_11139,N_9917,N_6337);
or U11140 (N_11140,N_6615,N_9706);
or U11141 (N_11141,N_7989,N_6142);
and U11142 (N_11142,N_6658,N_7867);
or U11143 (N_11143,N_7165,N_9558);
and U11144 (N_11144,N_7283,N_6522);
or U11145 (N_11145,N_7745,N_7966);
nor U11146 (N_11146,N_6799,N_5599);
and U11147 (N_11147,N_8189,N_9455);
nand U11148 (N_11148,N_8958,N_5781);
nor U11149 (N_11149,N_7517,N_6634);
nor U11150 (N_11150,N_7217,N_6237);
nand U11151 (N_11151,N_8422,N_7033);
and U11152 (N_11152,N_7163,N_8052);
or U11153 (N_11153,N_7623,N_5629);
xnor U11154 (N_11154,N_6074,N_5775);
nand U11155 (N_11155,N_7027,N_6370);
nor U11156 (N_11156,N_8784,N_7469);
nand U11157 (N_11157,N_9762,N_8085);
and U11158 (N_11158,N_8230,N_6875);
and U11159 (N_11159,N_5945,N_5007);
or U11160 (N_11160,N_9456,N_7127);
and U11161 (N_11161,N_9134,N_5811);
nand U11162 (N_11162,N_6129,N_9600);
xnor U11163 (N_11163,N_9145,N_6514);
xor U11164 (N_11164,N_9125,N_7231);
xnor U11165 (N_11165,N_9257,N_9124);
nand U11166 (N_11166,N_5995,N_9090);
xor U11167 (N_11167,N_9039,N_6550);
nor U11168 (N_11168,N_5397,N_6884);
nand U11169 (N_11169,N_8491,N_7571);
nand U11170 (N_11170,N_5145,N_5594);
nand U11171 (N_11171,N_7608,N_5172);
nand U11172 (N_11172,N_7420,N_5732);
and U11173 (N_11173,N_6126,N_5156);
nand U11174 (N_11174,N_5970,N_7099);
or U11175 (N_11175,N_6826,N_5267);
or U11176 (N_11176,N_8926,N_7462);
nor U11177 (N_11177,N_5905,N_5875);
nor U11178 (N_11178,N_7932,N_9789);
nand U11179 (N_11179,N_8629,N_7797);
and U11180 (N_11180,N_8360,N_8565);
nand U11181 (N_11181,N_8800,N_6732);
xnor U11182 (N_11182,N_7961,N_7816);
nor U11183 (N_11183,N_9548,N_5260);
or U11184 (N_11184,N_9953,N_7605);
and U11185 (N_11185,N_8543,N_6356);
or U11186 (N_11186,N_7713,N_5164);
or U11187 (N_11187,N_7693,N_6459);
and U11188 (N_11188,N_9977,N_5891);
nor U11189 (N_11189,N_6870,N_9923);
nor U11190 (N_11190,N_5238,N_5800);
and U11191 (N_11191,N_6616,N_8850);
nor U11192 (N_11192,N_8099,N_5535);
nand U11193 (N_11193,N_7954,N_7226);
nand U11194 (N_11194,N_6656,N_5039);
or U11195 (N_11195,N_5437,N_9012);
nand U11196 (N_11196,N_5846,N_6426);
nor U11197 (N_11197,N_5493,N_6670);
xnor U11198 (N_11198,N_9081,N_6740);
and U11199 (N_11199,N_5290,N_7133);
or U11200 (N_11200,N_5185,N_6500);
nand U11201 (N_11201,N_9332,N_7742);
nand U11202 (N_11202,N_7696,N_6133);
xnor U11203 (N_11203,N_6026,N_5897);
nand U11204 (N_11204,N_5020,N_8634);
nor U11205 (N_11205,N_5873,N_8657);
and U11206 (N_11206,N_6187,N_5613);
nand U11207 (N_11207,N_7923,N_6659);
nand U11208 (N_11208,N_6809,N_9530);
nand U11209 (N_11209,N_8369,N_5385);
or U11210 (N_11210,N_5129,N_9523);
nand U11211 (N_11211,N_9541,N_7715);
or U11212 (N_11212,N_5721,N_8833);
nor U11213 (N_11213,N_9528,N_5285);
or U11214 (N_11214,N_5735,N_7479);
xor U11215 (N_11215,N_5443,N_9576);
xnor U11216 (N_11216,N_6837,N_7825);
nand U11217 (N_11217,N_7354,N_6847);
and U11218 (N_11218,N_5752,N_9860);
nand U11219 (N_11219,N_7296,N_6599);
or U11220 (N_11220,N_8428,N_8481);
nor U11221 (N_11221,N_6958,N_5321);
xnor U11222 (N_11222,N_7722,N_5257);
and U11223 (N_11223,N_5499,N_6098);
or U11224 (N_11224,N_7482,N_6858);
and U11225 (N_11225,N_5125,N_8663);
and U11226 (N_11226,N_6773,N_5376);
nand U11227 (N_11227,N_7348,N_5641);
nor U11228 (N_11228,N_8592,N_7747);
xnor U11229 (N_11229,N_5673,N_5770);
or U11230 (N_11230,N_9247,N_7388);
and U11231 (N_11231,N_9132,N_5941);
or U11232 (N_11232,N_5057,N_5131);
and U11233 (N_11233,N_5824,N_5149);
and U11234 (N_11234,N_6083,N_6441);
nand U11235 (N_11235,N_8922,N_5597);
nor U11236 (N_11236,N_9489,N_9285);
and U11237 (N_11237,N_7379,N_7075);
and U11238 (N_11238,N_9871,N_8547);
and U11239 (N_11239,N_7249,N_9692);
nor U11240 (N_11240,N_8593,N_9077);
and U11241 (N_11241,N_8347,N_7372);
or U11242 (N_11242,N_8786,N_9688);
and U11243 (N_11243,N_7593,N_6951);
nand U11244 (N_11244,N_7986,N_5498);
nand U11245 (N_11245,N_7187,N_7259);
xnor U11246 (N_11246,N_6787,N_9669);
nand U11247 (N_11247,N_7876,N_8076);
and U11248 (N_11248,N_5751,N_6350);
or U11249 (N_11249,N_9407,N_9854);
nand U11250 (N_11250,N_5071,N_9295);
or U11251 (N_11251,N_8367,N_9067);
or U11252 (N_11252,N_7602,N_7247);
nor U11253 (N_11253,N_5058,N_8178);
xor U11254 (N_11254,N_9254,N_9862);
and U11255 (N_11255,N_9830,N_9657);
nand U11256 (N_11256,N_7279,N_5928);
nor U11257 (N_11257,N_8375,N_6697);
and U11258 (N_11258,N_9820,N_7764);
and U11259 (N_11259,N_9494,N_5277);
or U11260 (N_11260,N_6399,N_8909);
xnor U11261 (N_11261,N_7586,N_7178);
and U11262 (N_11262,N_5064,N_8749);
nor U11263 (N_11263,N_8161,N_7591);
nand U11264 (N_11264,N_6660,N_8734);
xor U11265 (N_11265,N_8965,N_8907);
and U11266 (N_11266,N_9417,N_9313);
xor U11267 (N_11267,N_8475,N_6205);
or U11268 (N_11268,N_8773,N_6169);
or U11269 (N_11269,N_5739,N_9209);
xnor U11270 (N_11270,N_6806,N_6242);
nor U11271 (N_11271,N_7601,N_6980);
xnor U11272 (N_11272,N_7403,N_6017);
and U11273 (N_11273,N_6618,N_5809);
xnor U11274 (N_11274,N_9510,N_7134);
nor U11275 (N_11275,N_9602,N_9173);
nor U11276 (N_11276,N_7670,N_9610);
or U11277 (N_11277,N_5042,N_6699);
or U11278 (N_11278,N_8185,N_5215);
nand U11279 (N_11279,N_6937,N_9121);
xnor U11280 (N_11280,N_6429,N_5063);
xnor U11281 (N_11281,N_9471,N_5940);
and U11282 (N_11282,N_7594,N_8082);
nor U11283 (N_11283,N_6778,N_9076);
xor U11284 (N_11284,N_8087,N_8083);
nor U11285 (N_11285,N_7208,N_5349);
and U11286 (N_11286,N_8183,N_6202);
xor U11287 (N_11287,N_9386,N_9588);
nor U11288 (N_11288,N_9993,N_9973);
and U11289 (N_11289,N_8275,N_5073);
nand U11290 (N_11290,N_5816,N_9224);
xor U11291 (N_11291,N_5723,N_6464);
xnor U11292 (N_11292,N_6788,N_9127);
nor U11293 (N_11293,N_5515,N_7521);
nor U11294 (N_11294,N_6073,N_5361);
and U11295 (N_11295,N_6891,N_8644);
and U11296 (N_11296,N_6204,N_6565);
xor U11297 (N_11297,N_8003,N_5505);
or U11298 (N_11298,N_6855,N_7458);
and U11299 (N_11299,N_5678,N_5999);
xor U11300 (N_11300,N_5446,N_6703);
xor U11301 (N_11301,N_6856,N_6690);
or U11302 (N_11302,N_5651,N_9493);
nor U11303 (N_11303,N_5354,N_5085);
xnor U11304 (N_11304,N_8878,N_7048);
or U11305 (N_11305,N_8453,N_8304);
and U11306 (N_11306,N_9837,N_5240);
nor U11307 (N_11307,N_6152,N_9465);
and U11308 (N_11308,N_5211,N_7309);
nand U11309 (N_11309,N_9653,N_7863);
or U11310 (N_11310,N_8425,N_8242);
nor U11311 (N_11311,N_7842,N_5430);
or U11312 (N_11312,N_5729,N_7390);
and U11313 (N_11313,N_6751,N_9432);
nand U11314 (N_11314,N_6428,N_6562);
nor U11315 (N_11315,N_6141,N_5501);
nand U11316 (N_11316,N_8672,N_8040);
nand U11317 (N_11317,N_9384,N_9028);
nand U11318 (N_11318,N_7704,N_7725);
or U11319 (N_11319,N_8529,N_8268);
nand U11320 (N_11320,N_5720,N_8664);
nor U11321 (N_11321,N_8255,N_5797);
xor U11322 (N_11322,N_7406,N_8088);
xor U11323 (N_11323,N_5899,N_9423);
nor U11324 (N_11324,N_5555,N_7471);
and U11325 (N_11325,N_5353,N_6805);
or U11326 (N_11326,N_5259,N_7338);
and U11327 (N_11327,N_9951,N_5664);
or U11328 (N_11328,N_7877,N_6635);
nand U11329 (N_11329,N_8929,N_7957);
or U11330 (N_11330,N_9123,N_7277);
and U11331 (N_11331,N_7193,N_9501);
nand U11332 (N_11332,N_9546,N_9892);
or U11333 (N_11333,N_5715,N_6719);
and U11334 (N_11334,N_6078,N_7930);
and U11335 (N_11335,N_5686,N_8975);
and U11336 (N_11336,N_9879,N_8387);
or U11337 (N_11337,N_5426,N_5347);
and U11338 (N_11338,N_5790,N_9544);
nand U11339 (N_11339,N_7809,N_9358);
and U11340 (N_11340,N_6391,N_8826);
xnor U11341 (N_11341,N_6085,N_7339);
nand U11342 (N_11342,N_9962,N_9433);
nor U11343 (N_11343,N_8571,N_8816);
and U11344 (N_11344,N_9650,N_6571);
nand U11345 (N_11345,N_9747,N_8044);
or U11346 (N_11346,N_8978,N_6398);
and U11347 (N_11347,N_7839,N_5204);
and U11348 (N_11348,N_7086,N_9765);
and U11349 (N_11349,N_9678,N_5936);
and U11350 (N_11350,N_7294,N_5930);
nor U11351 (N_11351,N_7120,N_8295);
and U11352 (N_11352,N_6369,N_7215);
xnor U11353 (N_11353,N_7652,N_7699);
nand U11354 (N_11354,N_7979,N_7487);
or U11355 (N_11355,N_8681,N_8449);
xnor U11356 (N_11356,N_7142,N_7529);
and U11357 (N_11357,N_5741,N_6225);
nor U11358 (N_11358,N_9864,N_7893);
xnor U11359 (N_11359,N_6316,N_9310);
and U11360 (N_11360,N_8150,N_7634);
and U11361 (N_11361,N_8665,N_8300);
and U11362 (N_11362,N_9370,N_6552);
xor U11363 (N_11363,N_6501,N_8163);
and U11364 (N_11364,N_6314,N_6253);
xnor U11365 (N_11365,N_8194,N_5208);
and U11366 (N_11366,N_5848,N_6830);
nor U11367 (N_11367,N_7727,N_7297);
nor U11368 (N_11368,N_6212,N_9069);
or U11369 (N_11369,N_6410,N_5670);
nor U11370 (N_11370,N_9129,N_8437);
xnor U11371 (N_11371,N_9859,N_8345);
and U11372 (N_11372,N_8351,N_7196);
and U11373 (N_11373,N_5825,N_6602);
or U11374 (N_11374,N_9907,N_8924);
or U11375 (N_11375,N_6120,N_9112);
xor U11376 (N_11376,N_5075,N_6929);
nor U11377 (N_11377,N_5758,N_6495);
nand U11378 (N_11378,N_7037,N_7599);
nand U11379 (N_11379,N_9256,N_9377);
nor U11380 (N_11380,N_6600,N_9679);
xnor U11381 (N_11381,N_9239,N_8602);
or U11382 (N_11382,N_5340,N_6461);
nand U11383 (N_11383,N_5776,N_6052);
and U11384 (N_11384,N_5137,N_8192);
nand U11385 (N_11385,N_5357,N_6537);
nand U11386 (N_11386,N_8487,N_5432);
xor U11387 (N_11387,N_8652,N_9715);
nor U11388 (N_11388,N_6881,N_6708);
xor U11389 (N_11389,N_8007,N_7691);
nor U11390 (N_11390,N_5320,N_8995);
nor U11391 (N_11391,N_6945,N_6695);
and U11392 (N_11392,N_9926,N_5773);
or U11393 (N_11393,N_7535,N_9130);
and U11394 (N_11394,N_6143,N_7844);
xnor U11395 (N_11395,N_8454,N_6145);
nor U11396 (N_11396,N_9298,N_6900);
and U11397 (N_11397,N_7697,N_7726);
nand U11398 (N_11398,N_7435,N_6303);
nand U11399 (N_11399,N_8662,N_6275);
nand U11400 (N_11400,N_7566,N_5917);
nor U11401 (N_11401,N_8047,N_9232);
nor U11402 (N_11402,N_6906,N_6424);
and U11403 (N_11403,N_5360,N_7365);
nor U11404 (N_11404,N_7389,N_6633);
and U11405 (N_11405,N_8837,N_8821);
nor U11406 (N_11406,N_7449,N_7526);
and U11407 (N_11407,N_6519,N_5078);
and U11408 (N_11408,N_6717,N_6155);
and U11409 (N_11409,N_8707,N_6492);
nor U11410 (N_11410,N_5702,N_7874);
nor U11411 (N_11411,N_5514,N_8756);
nor U11412 (N_11412,N_6923,N_8207);
nor U11413 (N_11413,N_5198,N_6470);
xnor U11414 (N_11414,N_7625,N_5622);
and U11415 (N_11415,N_6233,N_8265);
or U11416 (N_11416,N_8531,N_5479);
nor U11417 (N_11417,N_9053,N_6907);
nand U11418 (N_11418,N_6709,N_5624);
xnor U11419 (N_11419,N_7925,N_8450);
xnor U11420 (N_11420,N_8934,N_7592);
nor U11421 (N_11421,N_9343,N_8900);
xnor U11422 (N_11422,N_6752,N_9281);
xnor U11423 (N_11423,N_5034,N_7576);
nor U11424 (N_11424,N_6944,N_5519);
xor U11425 (N_11425,N_5558,N_7560);
and U11426 (N_11426,N_7025,N_7703);
and U11427 (N_11427,N_9435,N_7640);
and U11428 (N_11428,N_8853,N_9168);
or U11429 (N_11429,N_5314,N_8363);
nor U11430 (N_11430,N_9084,N_6731);
or U11431 (N_11431,N_6176,N_6305);
xnor U11432 (N_11432,N_7201,N_7513);
xor U11433 (N_11433,N_5959,N_6070);
or U11434 (N_11434,N_5769,N_5148);
nor U11435 (N_11435,N_5045,N_7999);
nand U11436 (N_11436,N_5957,N_9726);
nor U11437 (N_11437,N_9161,N_6439);
nor U11438 (N_11438,N_7866,N_5021);
or U11439 (N_11439,N_6961,N_7668);
or U11440 (N_11440,N_8579,N_8171);
xor U11441 (N_11441,N_5134,N_9992);
nand U11442 (N_11442,N_6229,N_7243);
nand U11443 (N_11443,N_5562,N_6362);
and U11444 (N_11444,N_6182,N_5222);
nand U11445 (N_11445,N_8917,N_8869);
or U11446 (N_11446,N_8769,N_7224);
nand U11447 (N_11447,N_6605,N_6800);
xor U11448 (N_11448,N_9398,N_7630);
and U11449 (N_11449,N_5513,N_5804);
nand U11450 (N_11450,N_7322,N_7748);
nor U11451 (N_11451,N_7804,N_9590);
nand U11452 (N_11452,N_8889,N_8349);
nor U11453 (N_11453,N_5944,N_7790);
nand U11454 (N_11454,N_8130,N_6913);
xor U11455 (N_11455,N_9359,N_9160);
nor U11456 (N_11456,N_8002,N_9625);
xnor U11457 (N_11457,N_7061,N_7054);
nor U11458 (N_11458,N_7749,N_8865);
nand U11459 (N_11459,N_8607,N_9474);
and U11460 (N_11460,N_6529,N_7868);
or U11461 (N_11461,N_9041,N_9154);
nand U11462 (N_11462,N_7673,N_6040);
or U11463 (N_11463,N_8457,N_5400);
nor U11464 (N_11464,N_6224,N_5662);
nor U11465 (N_11465,N_9626,N_5660);
and U11466 (N_11466,N_5874,N_5286);
or U11467 (N_11467,N_5410,N_5840);
nand U11468 (N_11468,N_5027,N_5942);
or U11469 (N_11469,N_9808,N_5280);
nand U11470 (N_11470,N_5084,N_9791);
xnor U11471 (N_11471,N_7902,N_8258);
and U11472 (N_11472,N_6795,N_9998);
and U11473 (N_11473,N_8719,N_6448);
nor U11474 (N_11474,N_6877,N_5530);
and U11475 (N_11475,N_7846,N_9790);
or U11476 (N_11476,N_8271,N_5587);
and U11477 (N_11477,N_7765,N_7410);
xnor U11478 (N_11478,N_9253,N_9980);
and U11479 (N_11479,N_9066,N_6191);
or U11480 (N_11480,N_6796,N_8489);
nor U11481 (N_11481,N_5865,N_6171);
or U11482 (N_11482,N_5750,N_7991);
nor U11483 (N_11483,N_9095,N_6440);
or U11484 (N_11484,N_6488,N_7812);
nand U11485 (N_11485,N_5508,N_9094);
nor U11486 (N_11486,N_6114,N_5683);
xor U11487 (N_11487,N_9878,N_6072);
xnor U11488 (N_11488,N_5946,N_6081);
xnor U11489 (N_11489,N_9526,N_9071);
xnor U11490 (N_11490,N_7935,N_7650);
xnor U11491 (N_11491,N_5490,N_5199);
nand U11492 (N_11492,N_5630,N_7318);
or U11493 (N_11493,N_5485,N_8286);
nor U11494 (N_11494,N_8004,N_9444);
or U11495 (N_11495,N_8291,N_9231);
nand U11496 (N_11496,N_8341,N_8216);
nor U11497 (N_11497,N_6603,N_5543);
and U11498 (N_11498,N_5542,N_7323);
xor U11499 (N_11499,N_5831,N_8661);
nand U11500 (N_11500,N_7992,N_7589);
or U11501 (N_11501,N_6274,N_6767);
nand U11502 (N_11502,N_5762,N_6368);
and U11503 (N_11503,N_6664,N_9210);
nor U11504 (N_11504,N_7955,N_6789);
nor U11505 (N_11505,N_9408,N_7285);
and U11506 (N_11506,N_8809,N_5062);
nor U11507 (N_11507,N_9891,N_8799);
xnor U11508 (N_11508,N_5926,N_6014);
and U11509 (N_11509,N_6949,N_7945);
and U11510 (N_11510,N_8380,N_5000);
nand U11511 (N_11511,N_9884,N_8512);
or U11512 (N_11512,N_5807,N_5423);
xor U11513 (N_11513,N_6450,N_9920);
nand U11514 (N_11514,N_8070,N_6824);
or U11515 (N_11515,N_9460,N_6211);
nand U11516 (N_11516,N_7711,N_5167);
xor U11517 (N_11517,N_8915,N_8511);
and U11518 (N_11518,N_5090,N_6331);
and U11519 (N_11519,N_6782,N_8996);
nand U11520 (N_11520,N_8327,N_6755);
nand U11521 (N_11521,N_6159,N_9153);
nor U11522 (N_11522,N_6271,N_8575);
xor U11523 (N_11523,N_7371,N_8335);
or U11524 (N_11524,N_8469,N_8884);
or U11525 (N_11525,N_7503,N_7098);
xor U11526 (N_11526,N_9605,N_5251);
nor U11527 (N_11527,N_8912,N_8767);
nand U11528 (N_11528,N_9399,N_5019);
and U11529 (N_11529,N_7360,N_7971);
or U11530 (N_11530,N_9778,N_8383);
or U11531 (N_11531,N_8034,N_8352);
nor U11532 (N_11532,N_7158,N_9700);
nor U11533 (N_11533,N_8340,N_7920);
nor U11534 (N_11534,N_8342,N_6327);
nand U11535 (N_11535,N_8724,N_9540);
nand U11536 (N_11536,N_7063,N_8110);
or U11537 (N_11537,N_7367,N_5722);
nor U11538 (N_11538,N_9262,N_9305);
nor U11539 (N_11539,N_9314,N_7425);
nand U11540 (N_11540,N_8675,N_5912);
xor U11541 (N_11541,N_9872,N_9761);
nor U11542 (N_11542,N_5536,N_6974);
or U11543 (N_11543,N_6704,N_8564);
xnor U11544 (N_11544,N_5827,N_7434);
and U11545 (N_11545,N_8845,N_9150);
and U11546 (N_11546,N_6720,N_9676);
nand U11547 (N_11547,N_5888,N_6851);
nor U11548 (N_11548,N_8818,N_8406);
xor U11549 (N_11549,N_6538,N_7315);
nor U11550 (N_11550,N_7035,N_9612);
nor U11551 (N_11551,N_7835,N_7714);
nor U11552 (N_11552,N_6890,N_7501);
or U11553 (N_11553,N_7607,N_6213);
xnor U11554 (N_11554,N_5387,N_7953);
xor U11555 (N_11555,N_7047,N_5708);
nor U11556 (N_11556,N_8371,N_9326);
nand U11557 (N_11557,N_9648,N_5066);
and U11558 (N_11558,N_7737,N_9466);
xnor U11559 (N_11559,N_8720,N_8923);
nand U11560 (N_11560,N_9560,N_8443);
and U11561 (N_11561,N_5296,N_7881);
xor U11562 (N_11562,N_8122,N_9960);
or U11563 (N_11563,N_6994,N_6648);
or U11564 (N_11564,N_8840,N_9822);
nand U11565 (N_11565,N_6993,N_5261);
or U11566 (N_11566,N_9241,N_5478);
and U11567 (N_11567,N_8949,N_6366);
nor U11568 (N_11568,N_9696,N_8639);
nor U11569 (N_11569,N_9570,N_5009);
nand U11570 (N_11570,N_7507,N_9199);
nand U11571 (N_11571,N_7387,N_7916);
or U11572 (N_11572,N_8959,N_9832);
and U11573 (N_11573,N_5266,N_7160);
nor U11574 (N_11574,N_7020,N_9547);
and U11575 (N_11575,N_9567,N_7587);
xor U11576 (N_11576,N_9924,N_5572);
xnor U11577 (N_11577,N_8854,N_7679);
nor U11578 (N_11578,N_5229,N_5986);
nand U11579 (N_11579,N_7062,N_5880);
and U11580 (N_11580,N_7391,N_7860);
or U11581 (N_11581,N_5893,N_5717);
and U11582 (N_11582,N_7472,N_8465);
nor U11583 (N_11583,N_7043,N_7646);
nor U11584 (N_11584,N_5030,N_9018);
nor U11585 (N_11585,N_8166,N_6692);
nor U11586 (N_11586,N_9711,N_5301);
xnor U11587 (N_11587,N_8092,N_5367);
and U11588 (N_11588,N_5453,N_7060);
nor U11589 (N_11589,N_8472,N_8308);
xnor U11590 (N_11590,N_8495,N_6216);
or U11591 (N_11591,N_8987,N_7206);
and U11592 (N_11592,N_8976,N_5230);
or U11593 (N_11593,N_9063,N_8112);
nor U11594 (N_11594,N_9754,N_9760);
or U11595 (N_11595,N_7137,N_5806);
nand U11596 (N_11596,N_5409,N_6352);
xnor U11597 (N_11597,N_8008,N_6161);
and U11598 (N_11598,N_6414,N_8305);
nor U11599 (N_11599,N_6227,N_7308);
or U11600 (N_11600,N_7235,N_5151);
nor U11601 (N_11601,N_9497,N_9734);
or U11602 (N_11602,N_9395,N_6769);
nor U11603 (N_11603,N_7436,N_7861);
nand U11604 (N_11604,N_9904,N_6308);
nand U11605 (N_11605,N_7676,N_6223);
or U11606 (N_11606,N_8723,N_7880);
or U11607 (N_11607,N_9736,N_9731);
nor U11608 (N_11608,N_5862,N_9450);
xnor U11609 (N_11609,N_8266,N_6574);
nand U11610 (N_11610,N_8124,N_9834);
nand U11611 (N_11611,N_7871,N_9573);
or U11612 (N_11612,N_7654,N_9409);
xor U11613 (N_11613,N_7453,N_9243);
or U11614 (N_11614,N_8932,N_9900);
xnor U11615 (N_11615,N_6865,N_9847);
or U11616 (N_11616,N_9785,N_6150);
and U11617 (N_11617,N_8126,N_5931);
and U11618 (N_11618,N_5424,N_7428);
nor U11619 (N_11619,N_6939,N_5227);
nor U11620 (N_11620,N_8379,N_5763);
nor U11621 (N_11621,N_8631,N_8474);
or U11622 (N_11622,N_7834,N_8119);
and U11623 (N_11623,N_7756,N_9467);
nor U11624 (N_11624,N_9412,N_7744);
nand U11625 (N_11625,N_6832,N_8152);
xnor U11626 (N_11626,N_5774,N_9608);
and U11627 (N_11627,N_6091,N_7013);
nand U11628 (N_11628,N_9664,N_6693);
nor U11629 (N_11629,N_6194,N_6062);
xnor U11630 (N_11630,N_6381,N_8705);
or U11631 (N_11631,N_7218,N_9068);
and U11632 (N_11632,N_7578,N_8842);
and U11633 (N_11633,N_7255,N_8410);
nor U11634 (N_11634,N_9059,N_5345);
nand U11635 (N_11635,N_8042,N_9323);
and U11636 (N_11636,N_7172,N_6345);
nor U11637 (N_11637,N_6904,N_9278);
nor U11638 (N_11638,N_6587,N_6324);
nand U11639 (N_11639,N_9469,N_5710);
or U11640 (N_11640,N_5235,N_8279);
nor U11641 (N_11641,N_5948,N_5867);
nor U11642 (N_11642,N_6333,N_5887);
or U11643 (N_11643,N_5371,N_5906);
and U11644 (N_11644,N_6647,N_7965);
and U11645 (N_11645,N_5560,N_5918);
or U11646 (N_11646,N_9634,N_5405);
nor U11647 (N_11647,N_5243,N_6491);
xor U11648 (N_11648,N_9922,N_8277);
and U11649 (N_11649,N_5067,N_6646);
xor U11650 (N_11650,N_7439,N_9166);
and U11651 (N_11651,N_8954,N_5160);
or U11652 (N_11652,N_8196,N_6394);
nor U11653 (N_11653,N_8740,N_7921);
nor U11654 (N_11654,N_5676,N_7154);
nor U11655 (N_11655,N_7359,N_5685);
nand U11656 (N_11656,N_9330,N_9235);
nand U11657 (N_11657,N_9093,N_6838);
and U11658 (N_11658,N_7042,N_7141);
xnor U11659 (N_11659,N_8697,N_7307);
and U11660 (N_11660,N_5072,N_9190);
or U11661 (N_11661,N_6261,N_7240);
and U11662 (N_11662,N_5684,N_7952);
nor U11663 (N_11663,N_6099,N_6317);
or U11664 (N_11664,N_6149,N_9965);
nand U11665 (N_11665,N_9905,N_6170);
and U11666 (N_11666,N_8690,N_9371);
or U11667 (N_11667,N_6598,N_5178);
nand U11668 (N_11668,N_5333,N_7264);
xnor U11669 (N_11669,N_8055,N_6001);
nand U11670 (N_11670,N_7319,N_8856);
or U11671 (N_11671,N_9764,N_5889);
xor U11672 (N_11672,N_8455,N_8887);
nand U11673 (N_11673,N_5965,N_8789);
xnor U11674 (N_11674,N_9238,N_5054);
or U11675 (N_11675,N_6336,N_7818);
nor U11676 (N_11676,N_6024,N_8581);
xor U11677 (N_11677,N_8368,N_7089);
nor U11678 (N_11678,N_5133,N_7477);
and U11679 (N_11679,N_9662,N_8759);
and U11680 (N_11680,N_6926,N_8505);
nand U11681 (N_11681,N_6793,N_5241);
nor U11682 (N_11682,N_6340,N_5766);
or U11683 (N_11683,N_6156,N_7136);
xor U11684 (N_11684,N_6281,N_8633);
nand U11685 (N_11685,N_7198,N_5958);
xor U11686 (N_11686,N_5805,N_8957);
nor U11687 (N_11687,N_8742,N_6042);
or U11688 (N_11688,N_9581,N_7545);
nor U11689 (N_11689,N_6442,N_5879);
nor U11690 (N_11690,N_8315,N_9082);
xnor U11691 (N_11691,N_9026,N_8762);
and U11692 (N_11692,N_6018,N_8606);
or U11693 (N_11693,N_8180,N_8339);
xnor U11694 (N_11694,N_7357,N_5334);
or U11695 (N_11695,N_9640,N_9258);
xnor U11696 (N_11696,N_6241,N_5496);
or U11697 (N_11697,N_7305,N_7508);
nand U11698 (N_11698,N_7474,N_9441);
nor U11699 (N_11699,N_5193,N_7686);
xnor U11700 (N_11700,N_8777,N_5854);
xnor U11701 (N_11701,N_8782,N_9735);
and U11702 (N_11702,N_7175,N_5056);
and U11703 (N_11703,N_8372,N_9655);
or U11704 (N_11704,N_6027,N_6395);
and U11705 (N_11705,N_8000,N_5279);
and U11706 (N_11706,N_8238,N_9551);
nor U11707 (N_11707,N_7798,N_6266);
or U11708 (N_11708,N_8682,N_7651);
or U11709 (N_11709,N_6431,N_7002);
nand U11710 (N_11710,N_7750,N_5305);
or U11711 (N_11711,N_6706,N_9982);
or U11712 (N_11712,N_8968,N_7784);
and U11713 (N_11713,N_8963,N_7383);
nor U11714 (N_11714,N_6783,N_7252);
nand U11715 (N_11715,N_6524,N_7522);
or U11716 (N_11716,N_5705,N_7370);
and U11717 (N_11717,N_5140,N_9728);
or U11718 (N_11718,N_7232,N_6567);
or U11719 (N_11719,N_7463,N_5169);
nor U11720 (N_11720,N_9910,N_8736);
and U11721 (N_11721,N_5487,N_5417);
and U11722 (N_11722,N_5214,N_6808);
and U11723 (N_11723,N_8628,N_8796);
xnor U11724 (N_11724,N_6010,N_8525);
xor U11725 (N_11725,N_9695,N_9420);
xor U11726 (N_11726,N_8812,N_9478);
or U11727 (N_11727,N_6365,N_6814);
and U11728 (N_11728,N_7304,N_5546);
xor U11729 (N_11729,N_9411,N_9537);
nand U11730 (N_11730,N_6691,N_9609);
or U11731 (N_11731,N_7438,N_7802);
and U11732 (N_11732,N_9622,N_8109);
xor U11733 (N_11733,N_5512,N_9887);
nand U11734 (N_11734,N_5325,N_7514);
nor U11735 (N_11735,N_9684,N_5783);
nand U11736 (N_11736,N_5608,N_8524);
and U11737 (N_11737,N_8206,N_6776);
or U11738 (N_11738,N_9798,N_8413);
nor U11739 (N_11739,N_7888,N_9912);
nand U11740 (N_11740,N_8994,N_8820);
or U11741 (N_11741,N_5462,N_9753);
nand U11742 (N_11742,N_9368,N_9986);
xor U11743 (N_11743,N_9135,N_7057);
or U11744 (N_11744,N_5605,N_5294);
or U11745 (N_11745,N_5983,N_6807);
and U11746 (N_11746,N_8236,N_9671);
or U11747 (N_11747,N_7074,N_7862);
and U11748 (N_11748,N_7118,N_8643);
and U11749 (N_11749,N_7875,N_6510);
xor U11750 (N_11750,N_8671,N_8057);
and U11751 (N_11751,N_5511,N_8498);
nor U11752 (N_11752,N_6946,N_5464);
xor U11753 (N_11753,N_6248,N_7250);
xor U11754 (N_11754,N_8030,N_5549);
nand U11755 (N_11755,N_8942,N_8844);
nor U11756 (N_11756,N_5450,N_6942);
nand U11757 (N_11757,N_9226,N_8111);
and U11758 (N_11758,N_6853,N_7113);
xnor U11759 (N_11759,N_5456,N_6649);
and U11760 (N_11760,N_8385,N_5010);
or U11761 (N_11761,N_7124,N_5302);
nor U11762 (N_11762,N_7132,N_8165);
nor U11763 (N_11763,N_8205,N_5233);
xor U11764 (N_11764,N_8805,N_9175);
xnor U11765 (N_11765,N_7855,N_7260);
xnor U11766 (N_11766,N_8501,N_6511);
xor U11767 (N_11767,N_9284,N_5412);
xor U11768 (N_11768,N_8276,N_6134);
nand U11769 (N_11769,N_5829,N_8017);
nand U11770 (N_11770,N_9857,N_9172);
xor U11771 (N_11771,N_8500,N_6750);
nor U11772 (N_11772,N_6454,N_5012);
xor U11773 (N_11773,N_7476,N_5998);
and U11774 (N_11774,N_9842,N_9883);
nand U11775 (N_11775,N_8307,N_6509);
and U11776 (N_11776,N_9228,N_9259);
xnor U11777 (N_11777,N_7233,N_5517);
nor U11778 (N_11778,N_7574,N_9595);
nand U11779 (N_11779,N_7282,N_5551);
xnor U11780 (N_11780,N_5013,N_5987);
and U11781 (N_11781,N_7619,N_8029);
nor U11782 (N_11782,N_6047,N_5299);
nand U11783 (N_11783,N_5755,N_6055);
or U11784 (N_11784,N_9961,N_8128);
and U11785 (N_11785,N_5633,N_9823);
xor U11786 (N_11786,N_9562,N_7311);
nor U11787 (N_11787,N_8660,N_9010);
nor U11788 (N_11788,N_5975,N_9975);
or U11789 (N_11789,N_8768,N_9585);
and U11790 (N_11790,N_7228,N_9855);
nand U11791 (N_11791,N_7940,N_8814);
nor U11792 (N_11792,N_5668,N_6082);
nand U11793 (N_11793,N_5849,N_8532);
or U11794 (N_11794,N_8193,N_9710);
or U11795 (N_11795,N_8343,N_5128);
nand U11796 (N_11796,N_5909,N_9799);
nor U11797 (N_11797,N_7288,N_5377);
nor U11798 (N_11798,N_5190,N_6892);
nand U11799 (N_11799,N_8433,N_9458);
nor U11800 (N_11800,N_7488,N_5615);
nand U11801 (N_11801,N_9378,N_9512);
nor U11802 (N_11802,N_7626,N_9768);
nor U11803 (N_11803,N_5650,N_5180);
and U11804 (N_11804,N_5559,N_9324);
xnor U11805 (N_11805,N_6195,N_7666);
nand U11806 (N_11806,N_9824,N_7558);
nand U11807 (N_11807,N_9994,N_6566);
nand U11808 (N_11808,N_6577,N_9613);
xnor U11809 (N_11809,N_8866,N_8146);
or U11810 (N_11810,N_8309,N_8574);
nand U11811 (N_11811,N_7373,N_9527);
and U11812 (N_11812,N_9004,N_6210);
nand U11813 (N_11813,N_5439,N_6128);
or U11814 (N_11814,N_6811,N_9702);
xnor U11815 (N_11815,N_6127,N_9611);
or U11816 (N_11816,N_7664,N_5691);
nand U11817 (N_11817,N_6139,N_6992);
and U11818 (N_11818,N_8463,N_5666);
xnor U11819 (N_11819,N_7766,N_5883);
nor U11820 (N_11820,N_5444,N_6044);
nor U11821 (N_11821,N_9720,N_6494);
and U11822 (N_11822,N_5364,N_8755);
or U11823 (N_11823,N_7531,N_8282);
and U11824 (N_11824,N_8802,N_9732);
and U11825 (N_11825,N_9529,N_9380);
or U11826 (N_11826,N_6292,N_9268);
nand U11827 (N_11827,N_8225,N_9724);
xnor U11828 (N_11828,N_8897,N_6311);
xor U11829 (N_11829,N_7441,N_9752);
and U11830 (N_11830,N_6673,N_7169);
nor U11831 (N_11831,N_7741,N_6118);
nand U11832 (N_11832,N_8097,N_7755);
nand U11833 (N_11833,N_5029,N_5882);
xor U11834 (N_11834,N_6354,N_9717);
xor U11835 (N_11835,N_8728,N_7738);
xor U11836 (N_11836,N_9519,N_8158);
nor U11837 (N_11837,N_6287,N_7300);
or U11838 (N_11838,N_8832,N_9183);
xnor U11839 (N_11839,N_7702,N_6861);
nor U11840 (N_11840,N_7684,N_5682);
and U11841 (N_11841,N_6924,N_5256);
nor U11842 (N_11842,N_6950,N_5287);
nor U11843 (N_11843,N_7126,N_7779);
xnor U11844 (N_11844,N_9663,N_6116);
xor U11845 (N_11845,N_7492,N_8859);
and U11846 (N_11846,N_6513,N_9979);
or U11847 (N_11847,N_9895,N_5038);
or U11848 (N_11848,N_9448,N_9439);
xnor U11849 (N_11849,N_7083,N_5001);
xnor U11850 (N_11850,N_9572,N_8256);
xnor U11851 (N_11851,N_5777,N_8370);
nor U11852 (N_11852,N_5011,N_6810);
nor U11853 (N_11853,N_6160,N_9316);
nand U11854 (N_11854,N_8636,N_7024);
or U11855 (N_11855,N_9251,N_6543);
and U11856 (N_11856,N_9363,N_9617);
nor U11857 (N_11857,N_6059,N_5324);
or U11858 (N_11858,N_9532,N_6908);
xor U11859 (N_11859,N_6243,N_8626);
nor U11860 (N_11860,N_8045,N_5110);
nor U11861 (N_11861,N_8071,N_7355);
xor U11862 (N_11862,N_6976,N_5121);
or U11863 (N_11863,N_8435,N_8807);
xor U11864 (N_11864,N_6064,N_7036);
nand U11865 (N_11865,N_9714,N_8706);
and U11866 (N_11866,N_9913,N_6256);
and U11867 (N_11867,N_6265,N_9971);
xnor U11868 (N_11868,N_5886,N_9703);
or U11869 (N_11869,N_5356,N_6930);
nor U11870 (N_11870,N_6107,N_5808);
xor U11871 (N_11871,N_8653,N_9566);
xor U11872 (N_11872,N_6842,N_8817);
and U11873 (N_11873,N_5105,N_8984);
nor U11874 (N_11874,N_5489,N_9815);
and U11875 (N_11875,N_5339,N_8299);
or U11876 (N_11876,N_7754,N_6022);
nor U11877 (N_11877,N_9507,N_6386);
xor U11878 (N_11878,N_8601,N_8881);
nor U11879 (N_11879,N_6627,N_6592);
or U11880 (N_11880,N_8785,N_6269);
or U11881 (N_11881,N_5035,N_5471);
or U11882 (N_11882,N_5008,N_8157);
nand U11883 (N_11883,N_5326,N_5680);
nand U11884 (N_11884,N_8117,N_8765);
xnor U11885 (N_11885,N_9925,N_7316);
nand U11886 (N_11886,N_9499,N_5411);
xnor U11887 (N_11887,N_6249,N_8521);
xor U11888 (N_11888,N_6623,N_7153);
and U11889 (N_11889,N_6095,N_5206);
nor U11890 (N_11890,N_5447,N_5836);
nor U11891 (N_11891,N_7401,N_8488);
or U11892 (N_11892,N_5642,N_5351);
or U11893 (N_11893,N_7775,N_7038);
or U11894 (N_11894,N_8359,N_6712);
nor U11895 (N_11895,N_9178,N_7577);
nand U11896 (N_11896,N_9225,N_5368);
xnor U11897 (N_11897,N_7563,N_8434);
or U11898 (N_11898,N_7685,N_9394);
nor U11899 (N_11899,N_7130,N_9874);
xor U11900 (N_11900,N_5288,N_8955);
xor U11901 (N_11901,N_7897,N_8563);
and U11902 (N_11902,N_6654,N_8746);
xor U11903 (N_11903,N_5420,N_9445);
or U11904 (N_11904,N_9733,N_8125);
or U11905 (N_11905,N_9755,N_6586);
or U11906 (N_11906,N_7908,N_9177);
nor U11907 (N_11907,N_7538,N_7039);
nand U11908 (N_11908,N_6820,N_5116);
or U11909 (N_11909,N_7184,N_9559);
xnor U11910 (N_11910,N_6794,N_6353);
xnor U11911 (N_11911,N_9584,N_6867);
or U11912 (N_11912,N_5908,N_9350);
nand U11913 (N_11913,N_6655,N_5616);
and U11914 (N_11914,N_5264,N_8066);
nor U11915 (N_11915,N_6619,N_7800);
and U11916 (N_11916,N_8694,N_8151);
xor U11917 (N_11917,N_8891,N_9775);
or U11918 (N_11918,N_8555,N_5738);
and U11919 (N_11919,N_9630,N_5667);
nand U11920 (N_11920,N_5737,N_5375);
nand U11921 (N_11921,N_6104,N_7376);
nand U11922 (N_11922,N_5611,N_5142);
nand U11923 (N_11923,N_6677,N_6998);
and U11924 (N_11924,N_5547,N_9120);
xor U11925 (N_11925,N_6221,N_7678);
and U11926 (N_11926,N_5580,N_9184);
nand U11927 (N_11927,N_8065,N_9583);
nor U11928 (N_11928,N_9749,N_7055);
nor U11929 (N_11929,N_8562,N_5181);
nor U11930 (N_11930,N_6157,N_7342);
xnor U11931 (N_11931,N_8977,N_6910);
xnor U11932 (N_11932,N_8199,N_9340);
and U11933 (N_11933,N_7106,N_9186);
and U11934 (N_11934,N_7776,N_6544);
nor U11935 (N_11935,N_9171,N_8025);
nand U11936 (N_11936,N_9007,N_7878);
xor U11937 (N_11937,N_8081,N_5761);
and U11938 (N_11938,N_6090,N_8729);
or U11939 (N_11939,N_8459,N_9944);
xor U11940 (N_11940,N_6823,N_8091);
and U11941 (N_11941,N_7380,N_8129);
xnor U11942 (N_11942,N_9320,N_7533);
xnor U11943 (N_11943,N_5278,N_5838);
nand U11944 (N_11944,N_7918,N_5541);
and U11945 (N_11945,N_9737,N_9587);
nor U11946 (N_11946,N_8885,N_9807);
nor U11947 (N_11947,N_6164,N_7266);
nor U11948 (N_11948,N_7384,N_8278);
xor U11949 (N_11949,N_6578,N_7770);
nor U11950 (N_11950,N_5418,N_7924);
or U11951 (N_11951,N_8638,N_9353);
nand U11952 (N_11952,N_6496,N_8101);
or U11953 (N_11953,N_9938,N_7207);
and U11954 (N_11954,N_6446,N_9486);
and U11955 (N_11955,N_9430,N_9946);
nand U11956 (N_11956,N_6680,N_5147);
nand U11957 (N_11957,N_7824,N_7045);
and U11958 (N_11958,N_5782,N_5232);
xnor U11959 (N_11959,N_5265,N_9833);
or U11960 (N_11960,N_8294,N_5336);
or U11961 (N_11961,N_5174,N_5626);
nand U11962 (N_11962,N_7618,N_8533);
nand U11963 (N_11963,N_9809,N_5395);
xnor U11964 (N_11964,N_5709,N_5037);
or U11965 (N_11965,N_7734,N_6975);
and U11966 (N_11966,N_7452,N_9216);
nand U11967 (N_11967,N_9400,N_5403);
nor U11968 (N_11968,N_7071,N_7889);
and U11969 (N_11969,N_6569,N_9939);
xnor U11970 (N_11970,N_5924,N_7723);
nand U11971 (N_11971,N_5153,N_5404);
xnor U11972 (N_11972,N_7059,N_5964);
nand U11973 (N_11973,N_8334,N_8783);
xor U11974 (N_11974,N_7753,N_9525);
nand U11975 (N_11975,N_9495,N_7557);
nand U11976 (N_11976,N_8172,N_8591);
nand U11977 (N_11977,N_5304,N_5189);
nand U11978 (N_11978,N_9212,N_7227);
or U11979 (N_11979,N_9571,N_9575);
or U11980 (N_11980,N_9452,N_9821);
or U11981 (N_11981,N_5522,N_8228);
or U11982 (N_11982,N_8714,N_7847);
or U11983 (N_11983,N_7411,N_8153);
xnor U11984 (N_11984,N_9756,N_6471);
and U11985 (N_11985,N_7943,N_7377);
nor U11986 (N_11986,N_6199,N_8577);
xnor U11987 (N_11987,N_5374,N_9996);
or U11988 (N_11988,N_9426,N_5488);
nand U11989 (N_11989,N_5344,N_7203);
nor U11990 (N_11990,N_5176,N_7929);
nor U11991 (N_11991,N_6852,N_8691);
nor U11992 (N_11992,N_9058,N_5933);
nor U11993 (N_11993,N_6112,N_9034);
or U11994 (N_11994,N_8715,N_8229);
nor U11995 (N_11995,N_8913,N_8863);
nor U11996 (N_11996,N_7683,N_8918);
nand U11997 (N_11997,N_7799,N_6349);
nand U11998 (N_11998,N_7195,N_5123);
or U11999 (N_11999,N_8246,N_8362);
or U12000 (N_12000,N_6652,N_8950);
nor U12001 (N_12001,N_6037,N_6280);
nand U12002 (N_12002,N_9774,N_9376);
and U12003 (N_12003,N_7023,N_9170);
nand U12004 (N_12004,N_5554,N_6758);
or U12005 (N_12005,N_5796,N_8018);
and U12006 (N_12006,N_9656,N_7219);
nor U12007 (N_12007,N_8056,N_7814);
nand U12008 (N_12008,N_7021,N_8069);
nor U12009 (N_12009,N_5196,N_5923);
xor U12010 (N_12010,N_7739,N_7001);
and U12011 (N_12011,N_5910,N_5845);
or U12012 (N_12012,N_9140,N_8164);
and U12013 (N_12013,N_8395,N_6144);
or U12014 (N_12014,N_7088,N_5087);
or U12015 (N_12015,N_7223,N_6821);
nor U12016 (N_12016,N_6075,N_6009);
nor U12017 (N_12017,N_5192,N_6780);
and U12018 (N_12018,N_5435,N_5639);
nor U12019 (N_12019,N_5445,N_9916);
nor U12020 (N_12020,N_6084,N_6196);
and U12021 (N_12021,N_8234,N_9899);
nor U12022 (N_12022,N_8330,N_6973);
and U12023 (N_12023,N_8418,N_5262);
xor U12024 (N_12024,N_9930,N_8310);
nor U12025 (N_12025,N_5857,N_7352);
xnor U12026 (N_12026,N_9045,N_8323);
and U12027 (N_12027,N_8324,N_8134);
xor U12028 (N_12028,N_9784,N_9896);
or U12029 (N_12029,N_6060,N_5953);
xor U12030 (N_12030,N_9888,N_8133);
nor U12031 (N_12031,N_6006,N_6933);
and U12032 (N_12032,N_5026,N_7467);
nor U12033 (N_12033,N_7107,N_5388);
and U12034 (N_12034,N_9321,N_5561);
xor U12035 (N_12035,N_5618,N_6594);
nand U12036 (N_12036,N_9325,N_6614);
xnor U12037 (N_12037,N_7782,N_5820);
xor U12038 (N_12038,N_8553,N_5155);
nand U12039 (N_12039,N_6848,N_8819);
nor U12040 (N_12040,N_7237,N_7395);
and U12041 (N_12041,N_5581,N_6456);
and U12042 (N_12042,N_7689,N_5427);
nand U12043 (N_12043,N_6005,N_9999);
or U12044 (N_12044,N_5221,N_6416);
and U12045 (N_12045,N_7820,N_9180);
nor U12046 (N_12046,N_5234,N_8033);
and U12047 (N_12047,N_6294,N_6344);
and U12048 (N_12048,N_6438,N_8645);
or U12049 (N_12049,N_5839,N_5943);
and U12050 (N_12050,N_7519,N_8864);
xnor U12051 (N_12051,N_9220,N_5433);
and U12052 (N_12052,N_5585,N_7642);
nor U12053 (N_12053,N_7481,N_5242);
and U12054 (N_12054,N_7221,N_5843);
xnor U12055 (N_12055,N_6726,N_6102);
nand U12056 (N_12056,N_9182,N_5014);
or U12057 (N_12057,N_7665,N_9988);
or U12058 (N_12058,N_9943,N_9931);
or U12059 (N_12059,N_8538,N_8597);
xnor U12060 (N_12060,N_5532,N_7997);
nand U12061 (N_12061,N_6749,N_6572);
or U12062 (N_12062,N_6770,N_7780);
and U12063 (N_12063,N_9691,N_8650);
nor U12064 (N_12064,N_8103,N_9729);
xnor U12065 (N_12065,N_8190,N_6131);
and U12066 (N_12066,N_7409,N_8937);
nor U12067 (N_12067,N_6377,N_8655);
xnor U12068 (N_12068,N_9005,N_8336);
nor U12069 (N_12069,N_9742,N_9385);
nor U12070 (N_12070,N_8319,N_8224);
or U12071 (N_12071,N_9793,N_7489);
xor U12072 (N_12072,N_5461,N_8795);
xnor U12073 (N_12073,N_8354,N_7483);
and U12074 (N_12074,N_6251,N_9156);
xnor U12075 (N_12075,N_8108,N_5315);
nand U12076 (N_12076,N_5061,N_9851);
or U12077 (N_12077,N_7148,N_8732);
nand U12078 (N_12078,N_8557,N_7572);
and U12079 (N_12079,N_5300,N_7796);
nand U12080 (N_12080,N_8420,N_8050);
xnor U12081 (N_12081,N_9772,N_9771);
nand U12082 (N_12082,N_7366,N_7870);
or U12083 (N_12083,N_9621,N_6862);
xor U12084 (N_12084,N_7938,N_8415);
nor U12085 (N_12085,N_5954,N_9667);
nand U12086 (N_12086,N_5567,N_6389);
and U12087 (N_12087,N_9902,N_8757);
nor U12088 (N_12088,N_7465,N_6247);
nand U12089 (N_12089,N_9301,N_5481);
nor U12090 (N_12090,N_8441,N_6765);
nand U12091 (N_12091,N_7209,N_8576);
nor U12092 (N_12092,N_8289,N_8423);
nand U12093 (N_12093,N_6409,N_8329);
nor U12094 (N_12094,N_9308,N_5436);
and U12095 (N_12095,N_8741,N_8203);
xnor U12096 (N_12096,N_5484,N_7941);
xor U12097 (N_12097,N_9618,N_6978);
nand U12098 (N_12098,N_9083,N_5544);
or U12099 (N_12099,N_9119,N_9620);
nor U12100 (N_12100,N_8618,N_6390);
or U12101 (N_12101,N_9927,N_9964);
or U12102 (N_12102,N_5731,N_7590);
xor U12103 (N_12103,N_5628,N_7067);
nand U12104 (N_12104,N_5313,N_9840);
nand U12105 (N_12105,N_7879,N_8685);
and U12106 (N_12106,N_6413,N_7674);
nor U12107 (N_12107,N_5004,N_8804);
or U12108 (N_12108,N_7706,N_9329);
nor U12109 (N_12109,N_9099,N_8585);
or U12110 (N_12110,N_5186,N_6641);
nor U12111 (N_12111,N_6925,N_6338);
nand U12112 (N_12112,N_8250,N_5794);
nor U12113 (N_12113,N_6487,N_7960);
xnor U12114 (N_12114,N_7254,N_5716);
or U12115 (N_12115,N_9373,N_6938);
xnor U12116 (N_12116,N_7553,N_6790);
and U12117 (N_12117,N_6499,N_5523);
xor U12118 (N_12118,N_5812,N_6650);
nand U12119 (N_12119,N_9697,N_5005);
nand U12120 (N_12120,N_9360,N_8674);
xor U12121 (N_12121,N_6741,N_6888);
nand U12122 (N_12122,N_6065,N_5911);
and U12123 (N_12123,N_7695,N_8293);
or U12124 (N_12124,N_7518,N_5083);
and U12125 (N_12125,N_8285,N_5695);
nand U12126 (N_12126,N_8401,N_8835);
or U12127 (N_12127,N_7356,N_9880);
xnor U12128 (N_12128,N_8382,N_6845);
and U12129 (N_12129,N_8730,N_9976);
or U12130 (N_12130,N_5671,N_8939);
xnor U12131 (N_12131,N_6966,N_6985);
xnor U12132 (N_12132,N_7909,N_6707);
nor U12133 (N_12133,N_6048,N_9016);
nand U12134 (N_12134,N_6866,N_7996);
nand U12135 (N_12135,N_7852,N_7854);
or U12136 (N_12136,N_8121,N_6962);
and U12137 (N_12137,N_6559,N_6657);
or U12138 (N_12138,N_8144,N_9914);
or U12139 (N_12139,N_7015,N_7180);
or U12140 (N_12140,N_5992,N_7303);
nor U12141 (N_12141,N_6163,N_7962);
nand U12142 (N_12142,N_8717,N_9339);
and U12143 (N_12143,N_6833,N_6380);
nor U12144 (N_12144,N_5677,N_6940);
or U12145 (N_12145,N_6685,N_7569);
or U12146 (N_12146,N_6798,N_7584);
xnor U12147 (N_12147,N_9280,N_5901);
and U12148 (N_12148,N_9773,N_7822);
nand U12149 (N_12149,N_9948,N_5470);
nand U12150 (N_12150,N_5223,N_9415);
and U12151 (N_12151,N_7162,N_7147);
nand U12152 (N_12152,N_7211,N_9128);
or U12153 (N_12153,N_5837,N_5937);
xnor U12154 (N_12154,N_7056,N_5665);
and U12155 (N_12155,N_9805,N_8281);
or U12156 (N_12156,N_5309,N_7041);
or U12157 (N_12157,N_5398,N_8554);
or U12158 (N_12158,N_7807,N_8651);
xor U12159 (N_12159,N_6743,N_6540);
nand U12160 (N_12160,N_5074,N_6136);
or U12161 (N_12161,N_5391,N_7212);
nand U12162 (N_12162,N_6825,N_9362);
xnor U12163 (N_12163,N_6087,N_9240);
nand U12164 (N_12164,N_9050,N_8416);
and U12165 (N_12165,N_5592,N_9344);
nor U12166 (N_12166,N_7904,N_6898);
and U12167 (N_12167,N_5871,N_9157);
and U12168 (N_12168,N_7332,N_7606);
xnor U12169 (N_12169,N_7967,N_8298);
or U12170 (N_12170,N_7189,N_8159);
and U12171 (N_12171,N_6956,N_7171);
and U12172 (N_12172,N_6757,N_7167);
nand U12173 (N_12173,N_6873,N_5289);
nand U12174 (N_12174,N_5207,N_5779);
and U12175 (N_12175,N_9249,N_8344);
nor U12176 (N_12176,N_5342,N_7681);
nor U12177 (N_12177,N_5218,N_8841);
or U12178 (N_12178,N_7638,N_6057);
or U12179 (N_12179,N_8301,N_7344);
nand U12180 (N_12180,N_7975,N_9061);
nor U12181 (N_12181,N_7448,N_9427);
and U12182 (N_12182,N_6526,N_5712);
nor U12183 (N_12183,N_5993,N_9533);
xnor U12184 (N_12184,N_8212,N_9750);
xor U12185 (N_12185,N_9383,N_9586);
and U12186 (N_12186,N_9306,N_8735);
or U12187 (N_12187,N_7717,N_9876);
and U12188 (N_12188,N_9104,N_8914);
xnor U12189 (N_12189,N_7119,N_6591);
or U12190 (N_12190,N_6109,N_7502);
and U12191 (N_12191,N_8898,N_7649);
nor U12192 (N_12192,N_7146,N_7791);
nand U12193 (N_12193,N_8208,N_9246);
nor U12194 (N_12194,N_9275,N_7851);
nor U12195 (N_12195,N_8793,N_6921);
or U12196 (N_12196,N_8676,N_6797);
nand U12197 (N_12197,N_7795,N_6181);
and U12198 (N_12198,N_8072,N_8143);
nor U12199 (N_12199,N_5003,N_7408);
nand U12200 (N_12200,N_6723,N_7121);
xor U12201 (N_12201,N_8377,N_9727);
or U12202 (N_12202,N_8426,N_9142);
and U12203 (N_12203,N_5832,N_5332);
nand U12204 (N_12204,N_6611,N_6922);
nor U12205 (N_12205,N_9738,N_6701);
nand U12206 (N_12206,N_7138,N_8408);
nor U12207 (N_12207,N_8485,N_5929);
and U12208 (N_12208,N_7094,N_9057);
and U12209 (N_12209,N_9536,N_9557);
and U12210 (N_12210,N_7633,N_6035);
and U12211 (N_12211,N_5082,N_9193);
nand U12212 (N_12212,N_6843,N_6186);
nor U12213 (N_12213,N_6802,N_5719);
nor U12214 (N_12214,N_8774,N_7430);
nand U12215 (N_12215,N_9354,N_8245);
nor U12216 (N_12216,N_9649,N_5040);
xor U12217 (N_12217,N_6235,N_9614);
xnor U12218 (N_12218,N_9712,N_9593);
nand U12219 (N_12219,N_8578,N_9623);
and U12220 (N_12220,N_7645,N_8982);
nand U12221 (N_12221,N_7271,N_7773);
xnor U12222 (N_12222,N_7003,N_7777);
xor U12223 (N_12223,N_9853,N_5099);
or U12224 (N_12224,N_9672,N_8656);
nand U12225 (N_12225,N_6276,N_7216);
nor U12226 (N_12226,N_7324,N_7864);
xor U12227 (N_12227,N_9985,N_6486);
nand U12228 (N_12228,N_5595,N_8612);
and U12229 (N_12229,N_8233,N_6206);
or U12230 (N_12230,N_8115,N_7811);
nand U12231 (N_12231,N_5935,N_6520);
nor U12232 (N_12232,N_7375,N_6257);
nor U12233 (N_12233,N_9651,N_9079);
xor U12234 (N_12234,N_9422,N_9578);
nand U12235 (N_12235,N_9334,N_6166);
xnor U12236 (N_12236,N_6244,N_9485);
and U12237 (N_12237,N_6296,N_8962);
or U12238 (N_12238,N_7017,N_7885);
or U12239 (N_12239,N_9743,N_9322);
xor U12240 (N_12240,N_8552,N_6947);
and U12241 (N_12241,N_9877,N_6100);
nand U12242 (N_12242,N_6304,N_8381);
nor U12243 (N_12243,N_5119,N_5382);
nand U12244 (N_12244,N_9476,N_5210);
nand U12245 (N_12245,N_8930,N_7451);
or U12246 (N_12246,N_7333,N_7251);
xor U12247 (N_12247,N_5451,N_6722);
nand U12248 (N_12248,N_7849,N_6523);
xnor U12249 (N_12249,N_6710,N_6718);
and U12250 (N_12250,N_9484,N_5441);
nand U12251 (N_12251,N_6817,N_7072);
nand U12252 (N_12252,N_7423,N_7337);
and U12253 (N_12253,N_5531,N_8979);
and U12254 (N_12254,N_8953,N_6561);
xnor U12255 (N_12255,N_5028,N_8584);
or U12256 (N_12256,N_5113,N_5219);
nand U12257 (N_12257,N_5772,N_5079);
xor U12258 (N_12258,N_9110,N_8753);
nand U12259 (N_12259,N_5927,N_5327);
and U12260 (N_12260,N_7716,N_9936);
nor U12261 (N_12261,N_9261,N_5861);
and U12262 (N_12262,N_6425,N_7554);
or U12263 (N_12263,N_9234,N_8608);
nand U12264 (N_12264,N_9708,N_9829);
nand U12265 (N_12265,N_8561,N_5366);
nor U12266 (N_12266,N_5644,N_7050);
nor U12267 (N_12267,N_9825,N_7977);
xnor U12268 (N_12268,N_7109,N_7018);
or U12269 (N_12269,N_6729,N_7843);
and U12270 (N_12270,N_7192,N_9418);
or U12271 (N_12271,N_7778,N_7536);
nor U12272 (N_12272,N_7497,N_6582);
nand U12273 (N_12273,N_6638,N_6863);
and U12274 (N_12274,N_6076,N_7534);
or U12275 (N_12275,N_8020,N_6174);
nor U12276 (N_12276,N_6698,N_8931);
xnor U12277 (N_12277,N_8713,N_6268);
or U12278 (N_12278,N_7400,N_8572);
and U12279 (N_12279,N_5674,N_8630);
and U12280 (N_12280,N_6568,N_7069);
xor U12281 (N_12281,N_5419,N_5127);
and U12282 (N_12282,N_8440,N_6367);
xor U12283 (N_12283,N_9413,N_7740);
xnor U12284 (N_12284,N_5126,N_8966);
nand U12285 (N_12285,N_7530,N_7478);
nor U12286 (N_12286,N_9133,N_8766);
and U12287 (N_12287,N_7444,N_9796);
nand U12288 (N_12288,N_8333,N_7826);
nor U12289 (N_12289,N_6291,N_6045);
xnor U12290 (N_12290,N_7898,N_9101);
nand U12291 (N_12291,N_8417,N_8064);
xnor U12292 (N_12292,N_6148,N_6841);
and U12293 (N_12293,N_9890,N_6716);
or U12294 (N_12294,N_6153,N_5681);
nor U12295 (N_12295,N_5092,N_9054);
nand U12296 (N_12296,N_7500,N_9553);
nor U12297 (N_12297,N_7853,N_5972);
or U12298 (N_12298,N_7031,N_9579);
or U12299 (N_12299,N_5139,N_7114);
and U12300 (N_12300,N_6267,N_5421);
or U12301 (N_12301,N_6088,N_7394);
nand U12302 (N_12302,N_7624,N_5401);
xor U12303 (N_12303,N_7244,N_5793);
xnor U12304 (N_12304,N_6049,N_9513);
xor U12305 (N_12305,N_8791,N_7421);
nor U12306 (N_12306,N_6132,N_8846);
or U12307 (N_12307,N_7936,N_8683);
or U12308 (N_12308,N_8886,N_8221);
and U12309 (N_12309,N_5552,N_5749);
xnor U12310 (N_12310,N_6008,N_7464);
xnor U12311 (N_12311,N_8920,N_7442);
nor U12312 (N_12312,N_5273,N_9488);
nand U12313 (N_12313,N_5991,N_6405);
nand U12314 (N_12314,N_5184,N_9564);
nand U12315 (N_12315,N_9504,N_9355);
nand U12316 (N_12316,N_5311,N_9289);
or U12317 (N_12317,N_7692,N_9205);
nand U12318 (N_12318,N_7511,N_9107);
nand U12319 (N_12319,N_7433,N_5747);
or U12320 (N_12320,N_6220,N_6298);
nor U12321 (N_12321,N_6360,N_8558);
xor U12322 (N_12322,N_7267,N_7836);
or U12323 (N_12323,N_6557,N_8442);
xnor U12324 (N_12324,N_8536,N_8043);
xor U12325 (N_12325,N_9954,N_5553);
or U12326 (N_12326,N_9694,N_5563);
xnor U12327 (N_12327,N_5136,N_6874);
nand U12328 (N_12328,N_8692,N_5146);
and U12329 (N_12329,N_9846,N_8544);
nand U12330 (N_12330,N_6332,N_7682);
nor U12331 (N_12331,N_6517,N_7276);
or U12332 (N_12332,N_6302,N_7543);
nor U12333 (N_12333,N_7418,N_8373);
or U12334 (N_12334,N_6584,N_6775);
or U12335 (N_12335,N_6259,N_7661);
xnor U12336 (N_12336,N_5365,N_8627);
nand U12337 (N_12337,N_5386,N_8867);
or U12338 (N_12338,N_8506,N_8517);
xor U12339 (N_12339,N_7636,N_5851);
nor U12340 (N_12340,N_9042,N_8273);
nor U12341 (N_12341,N_5272,N_9713);
nand U12342 (N_12342,N_7547,N_6321);
xnor U12343 (N_12343,N_6167,N_9291);
nor U12344 (N_12344,N_9841,N_7190);
and U12345 (N_12345,N_9040,N_8397);
nand U12346 (N_12346,N_9897,N_8223);
xnor U12347 (N_12347,N_5183,N_9263);
nor U12348 (N_12348,N_7230,N_5947);
and U12349 (N_12349,N_8877,N_9592);
xor U12350 (N_12350,N_9294,N_9969);
and U12351 (N_12351,N_5654,N_9952);
nand U12352 (N_12352,N_6754,N_9865);
xnor U12353 (N_12353,N_5679,N_5406);
nand U12354 (N_12354,N_9098,N_7946);
or U12355 (N_12355,N_8566,N_9885);
nor U12356 (N_12356,N_6288,N_6497);
nand U12357 (N_12357,N_6415,N_6964);
and U12358 (N_12358,N_7827,N_6071);
and U12359 (N_12359,N_8089,N_9151);
xor U12360 (N_12360,N_5657,N_7152);
nand U12361 (N_12361,N_5135,N_7600);
xnor U12362 (N_12362,N_5101,N_5803);
xnor U12363 (N_12363,N_7891,N_6315);
nand U12364 (N_12364,N_9654,N_5521);
nor U12365 (N_12365,N_9766,N_5698);
xor U12366 (N_12366,N_7528,N_8148);
and U12367 (N_12367,N_7783,N_6309);
nand U12368 (N_12368,N_7078,N_8016);
xnor U12369 (N_12369,N_5570,N_6342);
xnor U12370 (N_12370,N_5500,N_5097);
or U12371 (N_12371,N_8944,N_8061);
nand U12372 (N_12372,N_6111,N_9665);
xor U12373 (N_12373,N_5525,N_9797);
and U12374 (N_12374,N_8980,N_6932);
nand U12375 (N_12375,N_6458,N_7461);
and U12376 (N_12376,N_7194,N_6725);
nor U12377 (N_12377,N_7368,N_7026);
or U12378 (N_12378,N_6547,N_7561);
and U12379 (N_12379,N_9006,N_7032);
xnor U12380 (N_12380,N_5907,N_5202);
or U12381 (N_12381,N_6965,N_8215);
and U12382 (N_12382,N_7598,N_5392);
xnor U12383 (N_12383,N_8541,N_5396);
nor U12384 (N_12384,N_5088,N_9903);
or U12385 (N_12385,N_8244,N_6931);
nor U12386 (N_12386,N_7269,N_6990);
nor U12387 (N_12387,N_7667,N_7637);
or U12388 (N_12388,N_6421,N_9389);
and U12389 (N_12389,N_5425,N_8890);
nor U12390 (N_12390,N_6539,N_8492);
xor U12391 (N_12391,N_8080,N_7293);
or U12392 (N_12392,N_9211,N_5724);
and U12393 (N_12393,N_8700,N_9304);
nor U12394 (N_12394,N_6632,N_5330);
xor U12395 (N_12395,N_5509,N_9309);
or U12396 (N_12396,N_9462,N_8599);
nand U12397 (N_12397,N_9017,N_7327);
nand U12398 (N_12398,N_5474,N_5378);
or U12399 (N_12399,N_5158,N_6485);
nand U12400 (N_12400,N_6013,N_7949);
nand U12401 (N_12401,N_8084,N_5166);
and U12402 (N_12402,N_6117,N_6746);
nor U12403 (N_12403,N_7123,N_7398);
or U12404 (N_12404,N_7268,N_8677);
xor U12405 (N_12405,N_9552,N_8104);
nor U12406 (N_12406,N_8174,N_7470);
and U12407 (N_12407,N_9705,N_5080);
or U12408 (N_12408,N_6433,N_6771);
nand U12409 (N_12409,N_9516,N_9286);
nor U12410 (N_12410,N_5589,N_9660);
nor U12411 (N_12411,N_8935,N_9967);
and U12412 (N_12412,N_5106,N_9869);
or U12413 (N_12413,N_6318,N_7922);
xnor U12414 (N_12414,N_9627,N_6208);
xnor U12415 (N_12415,N_7819,N_8693);
and U12416 (N_12416,N_9096,N_9164);
nand U12417 (N_12417,N_9204,N_9165);
and U12418 (N_12418,N_9122,N_5976);
xor U12419 (N_12419,N_5086,N_6630);
or U12420 (N_12420,N_6781,N_5903);
nor U12421 (N_12421,N_5786,N_6518);
nand U12422 (N_12422,N_9858,N_7415);
xnor U12423 (N_12423,N_5818,N_9673);
or U12424 (N_12424,N_8320,N_8176);
xnor U12425 (N_12425,N_5283,N_5108);
nor U12426 (N_12426,N_6218,N_8827);
and U12427 (N_12427,N_6326,N_7597);
nor U12428 (N_12428,N_9668,N_9515);
xnor U12429 (N_12429,N_9886,N_5675);
nand U12430 (N_12430,N_9288,N_7978);
nand U12431 (N_12431,N_9346,N_7995);
nor U12432 (N_12432,N_5165,N_7671);
or U12433 (N_12433,N_9443,N_6675);
nor U12434 (N_12434,N_8829,N_8424);
and U12435 (N_12435,N_7759,N_6067);
or U12436 (N_12436,N_8132,N_9214);
nor U12437 (N_12437,N_9369,N_6411);
or U12438 (N_12438,N_6711,N_7856);
or U12439 (N_12439,N_9699,N_9248);
or U12440 (N_12440,N_8895,N_9131);
nand U12441 (N_12441,N_8790,N_7329);
xor U12442 (N_12442,N_8509,N_5791);
nor U12443 (N_12443,N_8288,N_8892);
xnor U12444 (N_12444,N_6988,N_6197);
nand U12445 (N_12445,N_5527,N_6860);
nand U12446 (N_12446,N_9352,N_8048);
nand U12447 (N_12447,N_6272,N_6097);
and U12448 (N_12448,N_6801,N_7512);
xnor U12449 (N_12449,N_6521,N_6246);
nor U12450 (N_12450,N_6193,N_9265);
and U12451 (N_12451,N_5801,N_7562);
xnor U12452 (N_12452,N_8113,N_8825);
and U12453 (N_12453,N_6734,N_5574);
nor U12454 (N_12454,N_8619,N_9144);
nor U12455 (N_12455,N_9136,N_7761);
and U12456 (N_12456,N_5182,N_8232);
or U12457 (N_12457,N_9293,N_5979);
or U12458 (N_12458,N_6745,N_6140);
or U12459 (N_12459,N_9303,N_8175);
nor U12460 (N_12460,N_7170,N_7402);
nand U12461 (N_12461,N_8145,N_6403);
xnor U12462 (N_12462,N_9414,N_8815);
nand U12463 (N_12463,N_9196,N_5856);
xor U12464 (N_12464,N_8451,N_7845);
and U12465 (N_12465,N_9539,N_5938);
and U12466 (N_12466,N_7969,N_7610);
nor U12467 (N_12467,N_5362,N_9928);
or U12468 (N_12468,N_8013,N_5495);
nor U12469 (N_12469,N_9219,N_6282);
xor U12470 (N_12470,N_6889,N_7174);
xnor U12471 (N_12471,N_5132,N_8983);
nand U12472 (N_12472,N_6536,N_6642);
and U12473 (N_12473,N_7769,N_7335);
nand U12474 (N_12474,N_7302,N_6319);
nand U12475 (N_12475,N_8974,N_8647);
nand U12476 (N_12476,N_6694,N_8331);
nand U12477 (N_12477,N_9461,N_8248);
nand U12478 (N_12478,N_5647,N_9269);
xor U12479 (N_12479,N_5274,N_5785);
nor U12480 (N_12480,N_5114,N_9176);
or U12481 (N_12481,N_7263,N_8510);
and U12482 (N_12482,N_8899,N_5316);
nor U12483 (N_12483,N_9538,N_8187);
and U12484 (N_12484,N_7440,N_5117);
xnor U12485 (N_12485,N_9087,N_5467);
or U12486 (N_12486,N_8916,N_6954);
nand U12487 (N_12487,N_7707,N_8617);
and U12488 (N_12488,N_7810,N_5745);
and U12489 (N_12489,N_5620,N_6262);
nor U12490 (N_12490,N_5217,N_9374);
and U12491 (N_12491,N_7567,N_5612);
xor U12492 (N_12492,N_9601,N_6563);
nor U12493 (N_12493,N_5491,N_7298);
and U12494 (N_12494,N_8218,N_9852);
nand U12495 (N_12495,N_6330,N_9661);
nand U12496 (N_12496,N_7096,N_5043);
xnor U12497 (N_12497,N_8507,N_9945);
nor U12498 (N_12498,N_7959,N_9638);
xor U12499 (N_12499,N_7858,N_6393);
xnor U12500 (N_12500,N_5126,N_7187);
xnor U12501 (N_12501,N_9381,N_7992);
nand U12502 (N_12502,N_8636,N_5398);
xnor U12503 (N_12503,N_9545,N_5127);
nand U12504 (N_12504,N_8237,N_7573);
nand U12505 (N_12505,N_9516,N_8046);
nor U12506 (N_12506,N_8515,N_7957);
xor U12507 (N_12507,N_7396,N_7987);
nor U12508 (N_12508,N_9384,N_6568);
nand U12509 (N_12509,N_8528,N_7181);
xor U12510 (N_12510,N_7250,N_8650);
xnor U12511 (N_12511,N_8003,N_6440);
and U12512 (N_12512,N_9270,N_5079);
xnor U12513 (N_12513,N_8568,N_7733);
xnor U12514 (N_12514,N_9892,N_5333);
nand U12515 (N_12515,N_5331,N_7590);
nand U12516 (N_12516,N_5315,N_6191);
nor U12517 (N_12517,N_9207,N_5894);
and U12518 (N_12518,N_7719,N_7776);
xor U12519 (N_12519,N_5045,N_7063);
nand U12520 (N_12520,N_7142,N_6445);
nand U12521 (N_12521,N_8280,N_9602);
or U12522 (N_12522,N_5134,N_5571);
or U12523 (N_12523,N_5724,N_9079);
xor U12524 (N_12524,N_6555,N_6431);
and U12525 (N_12525,N_9030,N_6346);
nor U12526 (N_12526,N_7009,N_9481);
xor U12527 (N_12527,N_7993,N_6431);
or U12528 (N_12528,N_6232,N_5919);
and U12529 (N_12529,N_6957,N_9419);
or U12530 (N_12530,N_6533,N_6843);
and U12531 (N_12531,N_8957,N_9860);
or U12532 (N_12532,N_7315,N_8361);
xor U12533 (N_12533,N_8921,N_7528);
or U12534 (N_12534,N_5352,N_7010);
or U12535 (N_12535,N_9778,N_7236);
and U12536 (N_12536,N_5550,N_6056);
nor U12537 (N_12537,N_9810,N_6176);
or U12538 (N_12538,N_7527,N_9345);
xnor U12539 (N_12539,N_9389,N_7079);
xnor U12540 (N_12540,N_5613,N_6923);
nand U12541 (N_12541,N_6685,N_7513);
xor U12542 (N_12542,N_9727,N_5719);
nand U12543 (N_12543,N_9325,N_9100);
or U12544 (N_12544,N_5054,N_9331);
and U12545 (N_12545,N_5032,N_9321);
and U12546 (N_12546,N_9252,N_9279);
or U12547 (N_12547,N_8251,N_7577);
and U12548 (N_12548,N_6568,N_7313);
nand U12549 (N_12549,N_7053,N_6515);
and U12550 (N_12550,N_8947,N_5522);
or U12551 (N_12551,N_6013,N_7050);
nor U12552 (N_12552,N_5907,N_6747);
and U12553 (N_12553,N_8125,N_8206);
and U12554 (N_12554,N_6112,N_5771);
or U12555 (N_12555,N_6304,N_9539);
xnor U12556 (N_12556,N_6153,N_7654);
nand U12557 (N_12557,N_8370,N_7912);
and U12558 (N_12558,N_7885,N_8979);
xnor U12559 (N_12559,N_7504,N_5848);
or U12560 (N_12560,N_5584,N_8776);
nand U12561 (N_12561,N_6802,N_9660);
or U12562 (N_12562,N_5483,N_9118);
nand U12563 (N_12563,N_7401,N_5915);
nor U12564 (N_12564,N_7995,N_9906);
xor U12565 (N_12565,N_7908,N_7808);
xor U12566 (N_12566,N_8705,N_7476);
nand U12567 (N_12567,N_7390,N_8782);
or U12568 (N_12568,N_8977,N_7429);
and U12569 (N_12569,N_5226,N_9508);
nor U12570 (N_12570,N_6791,N_5943);
xor U12571 (N_12571,N_6077,N_9068);
nor U12572 (N_12572,N_7732,N_5972);
nand U12573 (N_12573,N_5597,N_5484);
nand U12574 (N_12574,N_9338,N_7798);
xor U12575 (N_12575,N_5028,N_9056);
or U12576 (N_12576,N_5774,N_7837);
or U12577 (N_12577,N_7618,N_7982);
or U12578 (N_12578,N_7534,N_9428);
xnor U12579 (N_12579,N_8720,N_7275);
nand U12580 (N_12580,N_6717,N_7168);
xor U12581 (N_12581,N_9369,N_8335);
xnor U12582 (N_12582,N_7798,N_7034);
and U12583 (N_12583,N_8223,N_7481);
nor U12584 (N_12584,N_6115,N_7616);
xor U12585 (N_12585,N_8644,N_8579);
nor U12586 (N_12586,N_5548,N_9700);
nand U12587 (N_12587,N_9101,N_6430);
or U12588 (N_12588,N_9742,N_5082);
or U12589 (N_12589,N_7424,N_6726);
and U12590 (N_12590,N_6489,N_5772);
or U12591 (N_12591,N_5557,N_6997);
and U12592 (N_12592,N_5041,N_7714);
or U12593 (N_12593,N_8635,N_9066);
nand U12594 (N_12594,N_8071,N_9489);
xor U12595 (N_12595,N_6028,N_6142);
nor U12596 (N_12596,N_6538,N_8469);
nand U12597 (N_12597,N_6188,N_6400);
or U12598 (N_12598,N_9580,N_6829);
nor U12599 (N_12599,N_7537,N_5881);
and U12600 (N_12600,N_9549,N_6139);
and U12601 (N_12601,N_5956,N_5802);
nand U12602 (N_12602,N_7765,N_5639);
xnor U12603 (N_12603,N_5432,N_5463);
or U12604 (N_12604,N_6827,N_6387);
nor U12605 (N_12605,N_9233,N_7170);
xor U12606 (N_12606,N_8292,N_6343);
or U12607 (N_12607,N_6565,N_5157);
or U12608 (N_12608,N_8158,N_9376);
or U12609 (N_12609,N_7933,N_5967);
xnor U12610 (N_12610,N_6354,N_6534);
nand U12611 (N_12611,N_7385,N_6138);
nor U12612 (N_12612,N_7478,N_9265);
or U12613 (N_12613,N_5142,N_9405);
nand U12614 (N_12614,N_6604,N_7663);
or U12615 (N_12615,N_9569,N_9651);
or U12616 (N_12616,N_7759,N_5841);
or U12617 (N_12617,N_8441,N_8578);
nor U12618 (N_12618,N_8022,N_6509);
nand U12619 (N_12619,N_6397,N_5111);
nand U12620 (N_12620,N_7309,N_8050);
nand U12621 (N_12621,N_9684,N_9837);
nand U12622 (N_12622,N_9436,N_8866);
nand U12623 (N_12623,N_9839,N_6321);
nand U12624 (N_12624,N_6771,N_6135);
or U12625 (N_12625,N_7099,N_5659);
and U12626 (N_12626,N_6259,N_9456);
xnor U12627 (N_12627,N_9759,N_8255);
xor U12628 (N_12628,N_7709,N_9088);
and U12629 (N_12629,N_9351,N_5687);
nor U12630 (N_12630,N_9393,N_6767);
nand U12631 (N_12631,N_8833,N_6977);
and U12632 (N_12632,N_8353,N_8127);
and U12633 (N_12633,N_5717,N_5885);
or U12634 (N_12634,N_6683,N_9213);
and U12635 (N_12635,N_7592,N_6560);
and U12636 (N_12636,N_8461,N_6710);
or U12637 (N_12637,N_8000,N_5022);
nor U12638 (N_12638,N_7177,N_6491);
xnor U12639 (N_12639,N_5343,N_7616);
and U12640 (N_12640,N_8606,N_8052);
and U12641 (N_12641,N_7025,N_7165);
xor U12642 (N_12642,N_7029,N_6447);
or U12643 (N_12643,N_6159,N_9175);
nor U12644 (N_12644,N_5205,N_6099);
xor U12645 (N_12645,N_5720,N_7342);
and U12646 (N_12646,N_7692,N_5785);
or U12647 (N_12647,N_5436,N_7495);
nand U12648 (N_12648,N_6490,N_5830);
and U12649 (N_12649,N_6191,N_8744);
or U12650 (N_12650,N_5254,N_5919);
or U12651 (N_12651,N_9598,N_8042);
and U12652 (N_12652,N_7354,N_9918);
or U12653 (N_12653,N_5681,N_6008);
nand U12654 (N_12654,N_9948,N_9397);
or U12655 (N_12655,N_8110,N_7133);
xor U12656 (N_12656,N_5022,N_7240);
or U12657 (N_12657,N_5546,N_7704);
xor U12658 (N_12658,N_6435,N_9106);
xnor U12659 (N_12659,N_7139,N_8866);
nor U12660 (N_12660,N_8902,N_6027);
nand U12661 (N_12661,N_7504,N_7364);
xnor U12662 (N_12662,N_5119,N_6066);
nand U12663 (N_12663,N_5872,N_8142);
and U12664 (N_12664,N_6499,N_9609);
nand U12665 (N_12665,N_7233,N_7894);
or U12666 (N_12666,N_7408,N_6001);
xnor U12667 (N_12667,N_7960,N_7944);
xnor U12668 (N_12668,N_7819,N_9396);
and U12669 (N_12669,N_7962,N_9512);
xor U12670 (N_12670,N_5771,N_9126);
nand U12671 (N_12671,N_6244,N_9908);
nand U12672 (N_12672,N_7537,N_8550);
nor U12673 (N_12673,N_8634,N_6616);
or U12674 (N_12674,N_9286,N_6901);
or U12675 (N_12675,N_9124,N_6298);
xnor U12676 (N_12676,N_8415,N_5002);
xor U12677 (N_12677,N_5488,N_8251);
xnor U12678 (N_12678,N_7312,N_6976);
and U12679 (N_12679,N_5565,N_7526);
or U12680 (N_12680,N_6286,N_5321);
xnor U12681 (N_12681,N_8704,N_9343);
or U12682 (N_12682,N_7550,N_5766);
and U12683 (N_12683,N_7618,N_6715);
nor U12684 (N_12684,N_8054,N_5982);
or U12685 (N_12685,N_7079,N_5407);
nor U12686 (N_12686,N_8564,N_8645);
and U12687 (N_12687,N_5776,N_8888);
nand U12688 (N_12688,N_6428,N_5820);
nand U12689 (N_12689,N_6015,N_9395);
or U12690 (N_12690,N_9044,N_7072);
nor U12691 (N_12691,N_6313,N_7506);
xor U12692 (N_12692,N_5508,N_7819);
nor U12693 (N_12693,N_6977,N_5389);
xor U12694 (N_12694,N_7049,N_9164);
nand U12695 (N_12695,N_8820,N_6319);
nand U12696 (N_12696,N_7263,N_8533);
or U12697 (N_12697,N_8554,N_5465);
nor U12698 (N_12698,N_8318,N_7536);
nand U12699 (N_12699,N_6088,N_7919);
nor U12700 (N_12700,N_8512,N_5074);
and U12701 (N_12701,N_8959,N_7520);
xor U12702 (N_12702,N_6510,N_7321);
or U12703 (N_12703,N_6900,N_9833);
nand U12704 (N_12704,N_7851,N_8859);
and U12705 (N_12705,N_9356,N_8085);
and U12706 (N_12706,N_7865,N_8341);
nand U12707 (N_12707,N_8852,N_5938);
nand U12708 (N_12708,N_6765,N_7537);
nor U12709 (N_12709,N_8982,N_6632);
nand U12710 (N_12710,N_5856,N_5594);
and U12711 (N_12711,N_5409,N_8607);
nor U12712 (N_12712,N_9701,N_8856);
or U12713 (N_12713,N_5635,N_5092);
nor U12714 (N_12714,N_6294,N_9499);
nand U12715 (N_12715,N_5691,N_8841);
xor U12716 (N_12716,N_7520,N_8181);
nor U12717 (N_12717,N_7653,N_8700);
or U12718 (N_12718,N_9860,N_8789);
or U12719 (N_12719,N_6049,N_8850);
nand U12720 (N_12720,N_5929,N_6876);
nor U12721 (N_12721,N_7594,N_6981);
or U12722 (N_12722,N_8925,N_6425);
nor U12723 (N_12723,N_6363,N_5992);
nor U12724 (N_12724,N_9657,N_7529);
nor U12725 (N_12725,N_7414,N_8699);
nor U12726 (N_12726,N_8894,N_8202);
nand U12727 (N_12727,N_9920,N_7886);
and U12728 (N_12728,N_9222,N_6090);
nor U12729 (N_12729,N_8953,N_5745);
and U12730 (N_12730,N_5709,N_8865);
or U12731 (N_12731,N_6610,N_8527);
or U12732 (N_12732,N_8113,N_7202);
nand U12733 (N_12733,N_8017,N_6078);
nor U12734 (N_12734,N_7238,N_5701);
xor U12735 (N_12735,N_5331,N_8436);
xnor U12736 (N_12736,N_9842,N_6413);
nand U12737 (N_12737,N_7312,N_8518);
nand U12738 (N_12738,N_8026,N_7362);
and U12739 (N_12739,N_9536,N_5995);
or U12740 (N_12740,N_6554,N_8064);
and U12741 (N_12741,N_7319,N_8033);
xnor U12742 (N_12742,N_5408,N_8459);
nor U12743 (N_12743,N_9421,N_7515);
and U12744 (N_12744,N_9124,N_7334);
and U12745 (N_12745,N_9285,N_6099);
or U12746 (N_12746,N_9869,N_7453);
or U12747 (N_12747,N_5153,N_8696);
nand U12748 (N_12748,N_7601,N_5519);
nand U12749 (N_12749,N_7808,N_7903);
nand U12750 (N_12750,N_9264,N_6564);
or U12751 (N_12751,N_6813,N_6208);
or U12752 (N_12752,N_9069,N_5343);
and U12753 (N_12753,N_8011,N_7287);
and U12754 (N_12754,N_8968,N_7752);
nor U12755 (N_12755,N_8286,N_7181);
or U12756 (N_12756,N_8613,N_9634);
xnor U12757 (N_12757,N_8152,N_6650);
and U12758 (N_12758,N_7771,N_6434);
or U12759 (N_12759,N_9135,N_5192);
or U12760 (N_12760,N_6759,N_7207);
nor U12761 (N_12761,N_8809,N_6772);
or U12762 (N_12762,N_6903,N_6401);
or U12763 (N_12763,N_6639,N_7785);
nand U12764 (N_12764,N_8112,N_8886);
nand U12765 (N_12765,N_5397,N_7751);
and U12766 (N_12766,N_5199,N_9233);
or U12767 (N_12767,N_8465,N_9383);
or U12768 (N_12768,N_9592,N_5551);
or U12769 (N_12769,N_6501,N_5403);
xnor U12770 (N_12770,N_8266,N_5445);
and U12771 (N_12771,N_7618,N_9882);
xor U12772 (N_12772,N_6533,N_6761);
nand U12773 (N_12773,N_5354,N_8363);
or U12774 (N_12774,N_9333,N_8999);
or U12775 (N_12775,N_5658,N_5739);
or U12776 (N_12776,N_7911,N_8957);
or U12777 (N_12777,N_5942,N_6811);
and U12778 (N_12778,N_7418,N_6165);
or U12779 (N_12779,N_5687,N_5717);
or U12780 (N_12780,N_5254,N_6163);
nor U12781 (N_12781,N_8625,N_6391);
nor U12782 (N_12782,N_5979,N_7178);
or U12783 (N_12783,N_8117,N_5198);
or U12784 (N_12784,N_9416,N_8944);
and U12785 (N_12785,N_8525,N_9937);
or U12786 (N_12786,N_5492,N_9774);
xor U12787 (N_12787,N_9512,N_6084);
and U12788 (N_12788,N_6749,N_7491);
and U12789 (N_12789,N_7861,N_5754);
and U12790 (N_12790,N_5380,N_7298);
nand U12791 (N_12791,N_6640,N_5981);
nor U12792 (N_12792,N_9909,N_6624);
and U12793 (N_12793,N_5826,N_6663);
nand U12794 (N_12794,N_8409,N_5975);
nand U12795 (N_12795,N_5277,N_7371);
and U12796 (N_12796,N_9723,N_9040);
xnor U12797 (N_12797,N_7798,N_9011);
and U12798 (N_12798,N_9243,N_7476);
or U12799 (N_12799,N_7366,N_9149);
or U12800 (N_12800,N_7391,N_7426);
nor U12801 (N_12801,N_8063,N_7226);
or U12802 (N_12802,N_5459,N_7171);
or U12803 (N_12803,N_8470,N_6753);
nand U12804 (N_12804,N_5746,N_8684);
xnor U12805 (N_12805,N_9901,N_6734);
nand U12806 (N_12806,N_7298,N_8788);
and U12807 (N_12807,N_6153,N_7894);
nand U12808 (N_12808,N_7057,N_9358);
and U12809 (N_12809,N_6274,N_7330);
or U12810 (N_12810,N_7773,N_9012);
nor U12811 (N_12811,N_8539,N_7320);
and U12812 (N_12812,N_8843,N_7179);
or U12813 (N_12813,N_7897,N_8647);
xnor U12814 (N_12814,N_6151,N_7646);
nor U12815 (N_12815,N_6262,N_6032);
nand U12816 (N_12816,N_7230,N_7116);
or U12817 (N_12817,N_6601,N_5165);
nand U12818 (N_12818,N_7829,N_5543);
nor U12819 (N_12819,N_5755,N_7962);
and U12820 (N_12820,N_7677,N_9831);
nand U12821 (N_12821,N_7281,N_8469);
xor U12822 (N_12822,N_5385,N_9211);
and U12823 (N_12823,N_9536,N_6468);
and U12824 (N_12824,N_5560,N_7234);
or U12825 (N_12825,N_9087,N_9799);
and U12826 (N_12826,N_6048,N_7522);
nand U12827 (N_12827,N_8631,N_8368);
and U12828 (N_12828,N_9945,N_8390);
xnor U12829 (N_12829,N_6869,N_6852);
nand U12830 (N_12830,N_5539,N_5898);
xor U12831 (N_12831,N_9241,N_6044);
and U12832 (N_12832,N_9545,N_9817);
or U12833 (N_12833,N_6696,N_5924);
xnor U12834 (N_12834,N_5660,N_6875);
and U12835 (N_12835,N_6138,N_7114);
and U12836 (N_12836,N_8260,N_5589);
nand U12837 (N_12837,N_6030,N_6467);
nand U12838 (N_12838,N_6966,N_6708);
and U12839 (N_12839,N_8020,N_9648);
or U12840 (N_12840,N_5997,N_5444);
and U12841 (N_12841,N_7636,N_7563);
nor U12842 (N_12842,N_9826,N_7437);
and U12843 (N_12843,N_7948,N_7501);
and U12844 (N_12844,N_6083,N_7816);
and U12845 (N_12845,N_9164,N_6369);
or U12846 (N_12846,N_7226,N_9719);
nand U12847 (N_12847,N_7460,N_6647);
nor U12848 (N_12848,N_5921,N_7665);
or U12849 (N_12849,N_5677,N_9735);
xnor U12850 (N_12850,N_9360,N_8719);
nand U12851 (N_12851,N_8054,N_7690);
nor U12852 (N_12852,N_9724,N_6754);
xor U12853 (N_12853,N_7023,N_9319);
or U12854 (N_12854,N_8774,N_7714);
xor U12855 (N_12855,N_8031,N_8329);
and U12856 (N_12856,N_6478,N_6096);
or U12857 (N_12857,N_8177,N_6811);
xor U12858 (N_12858,N_6436,N_9075);
nor U12859 (N_12859,N_7319,N_9263);
or U12860 (N_12860,N_8573,N_5778);
nand U12861 (N_12861,N_7102,N_9148);
nand U12862 (N_12862,N_7121,N_6363);
xor U12863 (N_12863,N_7543,N_5412);
nor U12864 (N_12864,N_5266,N_5021);
xor U12865 (N_12865,N_8956,N_9262);
nor U12866 (N_12866,N_8867,N_8444);
nand U12867 (N_12867,N_6998,N_9510);
nand U12868 (N_12868,N_6628,N_9013);
nor U12869 (N_12869,N_7438,N_5006);
nand U12870 (N_12870,N_5581,N_7567);
and U12871 (N_12871,N_6356,N_9093);
and U12872 (N_12872,N_7918,N_8800);
nor U12873 (N_12873,N_7120,N_5590);
and U12874 (N_12874,N_7298,N_7136);
xnor U12875 (N_12875,N_8801,N_8207);
nor U12876 (N_12876,N_8287,N_9881);
or U12877 (N_12877,N_7167,N_6635);
nor U12878 (N_12878,N_5666,N_5771);
xor U12879 (N_12879,N_9750,N_7204);
nor U12880 (N_12880,N_8185,N_7094);
nand U12881 (N_12881,N_6000,N_5300);
nand U12882 (N_12882,N_5665,N_8203);
and U12883 (N_12883,N_9556,N_5693);
or U12884 (N_12884,N_9377,N_9411);
xor U12885 (N_12885,N_9023,N_9543);
or U12886 (N_12886,N_9191,N_8747);
and U12887 (N_12887,N_8555,N_7161);
nand U12888 (N_12888,N_7031,N_7362);
xor U12889 (N_12889,N_9224,N_5561);
nor U12890 (N_12890,N_6925,N_5825);
nand U12891 (N_12891,N_8815,N_5979);
or U12892 (N_12892,N_5394,N_9095);
nor U12893 (N_12893,N_7175,N_8022);
or U12894 (N_12894,N_9432,N_5391);
nand U12895 (N_12895,N_8872,N_9954);
nor U12896 (N_12896,N_8594,N_7831);
and U12897 (N_12897,N_8262,N_5038);
nand U12898 (N_12898,N_9246,N_9330);
nor U12899 (N_12899,N_7971,N_7769);
and U12900 (N_12900,N_9382,N_6196);
nor U12901 (N_12901,N_7007,N_6332);
or U12902 (N_12902,N_7731,N_7290);
and U12903 (N_12903,N_8073,N_6052);
and U12904 (N_12904,N_7147,N_9550);
nand U12905 (N_12905,N_7425,N_5157);
or U12906 (N_12906,N_7123,N_8566);
and U12907 (N_12907,N_5567,N_8954);
nor U12908 (N_12908,N_7407,N_8687);
xnor U12909 (N_12909,N_9763,N_5100);
and U12910 (N_12910,N_7126,N_7124);
nand U12911 (N_12911,N_9156,N_6385);
or U12912 (N_12912,N_9019,N_8833);
nand U12913 (N_12913,N_6720,N_9615);
or U12914 (N_12914,N_8659,N_8212);
nor U12915 (N_12915,N_8274,N_6018);
or U12916 (N_12916,N_6751,N_7336);
nor U12917 (N_12917,N_8221,N_8201);
nor U12918 (N_12918,N_7414,N_5560);
xor U12919 (N_12919,N_8766,N_7946);
and U12920 (N_12920,N_5934,N_5849);
nand U12921 (N_12921,N_5950,N_7322);
nor U12922 (N_12922,N_5045,N_5869);
or U12923 (N_12923,N_9735,N_5375);
xnor U12924 (N_12924,N_7151,N_6624);
nor U12925 (N_12925,N_8597,N_5290);
nor U12926 (N_12926,N_8785,N_8007);
nor U12927 (N_12927,N_7299,N_5017);
or U12928 (N_12928,N_8763,N_8251);
nand U12929 (N_12929,N_6326,N_9866);
nand U12930 (N_12930,N_9503,N_9946);
xor U12931 (N_12931,N_7016,N_5585);
and U12932 (N_12932,N_5593,N_8871);
xor U12933 (N_12933,N_5037,N_8095);
or U12934 (N_12934,N_8363,N_7734);
and U12935 (N_12935,N_8094,N_5707);
nor U12936 (N_12936,N_7106,N_5381);
xnor U12937 (N_12937,N_5660,N_9018);
or U12938 (N_12938,N_9088,N_7051);
nand U12939 (N_12939,N_8532,N_8111);
nor U12940 (N_12940,N_8039,N_7109);
and U12941 (N_12941,N_6044,N_5161);
or U12942 (N_12942,N_7021,N_5241);
and U12943 (N_12943,N_9479,N_5884);
nand U12944 (N_12944,N_5688,N_7724);
and U12945 (N_12945,N_6860,N_5149);
or U12946 (N_12946,N_5243,N_6019);
or U12947 (N_12947,N_6201,N_6994);
xor U12948 (N_12948,N_5054,N_7922);
nor U12949 (N_12949,N_5899,N_5334);
and U12950 (N_12950,N_7838,N_7784);
nor U12951 (N_12951,N_8738,N_9463);
nor U12952 (N_12952,N_9578,N_5924);
nand U12953 (N_12953,N_5374,N_7763);
nand U12954 (N_12954,N_9968,N_7940);
nand U12955 (N_12955,N_7820,N_8131);
and U12956 (N_12956,N_8572,N_5095);
nand U12957 (N_12957,N_6764,N_8226);
nor U12958 (N_12958,N_7327,N_6996);
and U12959 (N_12959,N_9424,N_7704);
or U12960 (N_12960,N_9102,N_7424);
nand U12961 (N_12961,N_7336,N_8540);
nand U12962 (N_12962,N_9962,N_7932);
and U12963 (N_12963,N_6973,N_5875);
or U12964 (N_12964,N_6043,N_6914);
and U12965 (N_12965,N_6460,N_8845);
xor U12966 (N_12966,N_7158,N_6335);
nand U12967 (N_12967,N_7418,N_9375);
xor U12968 (N_12968,N_5372,N_6164);
and U12969 (N_12969,N_9230,N_8956);
or U12970 (N_12970,N_7627,N_5872);
nor U12971 (N_12971,N_6461,N_5115);
and U12972 (N_12972,N_5267,N_8016);
or U12973 (N_12973,N_6112,N_7973);
xor U12974 (N_12974,N_8788,N_5841);
xor U12975 (N_12975,N_8631,N_9444);
or U12976 (N_12976,N_9843,N_7312);
nor U12977 (N_12977,N_8134,N_6798);
nand U12978 (N_12978,N_7052,N_7882);
nand U12979 (N_12979,N_6111,N_9819);
or U12980 (N_12980,N_9227,N_5265);
or U12981 (N_12981,N_9268,N_5215);
xor U12982 (N_12982,N_7476,N_7955);
or U12983 (N_12983,N_5607,N_8952);
xnor U12984 (N_12984,N_6969,N_5371);
xnor U12985 (N_12985,N_9988,N_9796);
nor U12986 (N_12986,N_9587,N_5079);
and U12987 (N_12987,N_9542,N_5547);
xnor U12988 (N_12988,N_7535,N_8057);
xor U12989 (N_12989,N_6244,N_5013);
xnor U12990 (N_12990,N_6005,N_5046);
xnor U12991 (N_12991,N_8185,N_5829);
xnor U12992 (N_12992,N_6442,N_5132);
nor U12993 (N_12993,N_6740,N_9890);
or U12994 (N_12994,N_9733,N_8111);
nor U12995 (N_12995,N_9932,N_5517);
and U12996 (N_12996,N_5626,N_7689);
and U12997 (N_12997,N_9227,N_8654);
nor U12998 (N_12998,N_6340,N_6706);
and U12999 (N_12999,N_8786,N_9140);
nand U13000 (N_13000,N_6283,N_5526);
or U13001 (N_13001,N_7627,N_7705);
and U13002 (N_13002,N_7006,N_5145);
or U13003 (N_13003,N_8723,N_8833);
xor U13004 (N_13004,N_8664,N_5921);
and U13005 (N_13005,N_6742,N_8464);
nor U13006 (N_13006,N_5333,N_6408);
nand U13007 (N_13007,N_7098,N_6298);
xnor U13008 (N_13008,N_9622,N_7458);
nand U13009 (N_13009,N_8548,N_9717);
nor U13010 (N_13010,N_7434,N_9367);
or U13011 (N_13011,N_9942,N_7842);
or U13012 (N_13012,N_5575,N_6470);
or U13013 (N_13013,N_6756,N_8687);
and U13014 (N_13014,N_5459,N_5918);
and U13015 (N_13015,N_9521,N_5755);
and U13016 (N_13016,N_6796,N_5395);
or U13017 (N_13017,N_8046,N_5192);
xor U13018 (N_13018,N_5999,N_6313);
nand U13019 (N_13019,N_9410,N_6619);
and U13020 (N_13020,N_8692,N_7854);
or U13021 (N_13021,N_5385,N_8926);
nand U13022 (N_13022,N_9139,N_5020);
nor U13023 (N_13023,N_5617,N_6382);
and U13024 (N_13024,N_5318,N_8332);
nand U13025 (N_13025,N_5764,N_8058);
nor U13026 (N_13026,N_7328,N_8726);
nor U13027 (N_13027,N_5841,N_5479);
nor U13028 (N_13028,N_8560,N_8991);
nand U13029 (N_13029,N_7897,N_5466);
nor U13030 (N_13030,N_8681,N_8493);
or U13031 (N_13031,N_7674,N_7923);
or U13032 (N_13032,N_7183,N_5496);
and U13033 (N_13033,N_8531,N_7070);
nand U13034 (N_13034,N_9225,N_5669);
nand U13035 (N_13035,N_8738,N_5931);
or U13036 (N_13036,N_5975,N_6559);
or U13037 (N_13037,N_8890,N_6489);
nand U13038 (N_13038,N_7839,N_8263);
xnor U13039 (N_13039,N_7711,N_9015);
xor U13040 (N_13040,N_9137,N_8096);
nor U13041 (N_13041,N_5321,N_8653);
nand U13042 (N_13042,N_9566,N_7889);
nand U13043 (N_13043,N_7501,N_6117);
xnor U13044 (N_13044,N_6562,N_8472);
nand U13045 (N_13045,N_7475,N_6147);
xor U13046 (N_13046,N_5749,N_9863);
xnor U13047 (N_13047,N_8254,N_8127);
or U13048 (N_13048,N_7813,N_6850);
xnor U13049 (N_13049,N_8666,N_8290);
and U13050 (N_13050,N_8546,N_5940);
and U13051 (N_13051,N_5559,N_5849);
nor U13052 (N_13052,N_6472,N_6575);
or U13053 (N_13053,N_9003,N_8440);
nor U13054 (N_13054,N_9054,N_7820);
and U13055 (N_13055,N_7342,N_5667);
nand U13056 (N_13056,N_8197,N_7200);
xor U13057 (N_13057,N_9953,N_7891);
xor U13058 (N_13058,N_6533,N_9864);
nor U13059 (N_13059,N_5288,N_5614);
xor U13060 (N_13060,N_8538,N_6767);
nor U13061 (N_13061,N_5614,N_7807);
xor U13062 (N_13062,N_5877,N_5600);
nand U13063 (N_13063,N_7167,N_8459);
and U13064 (N_13064,N_8371,N_7262);
and U13065 (N_13065,N_7034,N_7700);
nor U13066 (N_13066,N_7687,N_8748);
and U13067 (N_13067,N_5580,N_6967);
nor U13068 (N_13068,N_6637,N_5169);
and U13069 (N_13069,N_7897,N_5234);
or U13070 (N_13070,N_7809,N_9492);
xnor U13071 (N_13071,N_9838,N_6699);
nand U13072 (N_13072,N_8407,N_7500);
nand U13073 (N_13073,N_9467,N_5196);
and U13074 (N_13074,N_6893,N_9067);
nor U13075 (N_13075,N_9461,N_6671);
nor U13076 (N_13076,N_6473,N_6034);
and U13077 (N_13077,N_6914,N_9698);
nand U13078 (N_13078,N_6376,N_8642);
nand U13079 (N_13079,N_5412,N_5752);
or U13080 (N_13080,N_9183,N_8789);
nand U13081 (N_13081,N_8683,N_9111);
and U13082 (N_13082,N_6532,N_8046);
nand U13083 (N_13083,N_9007,N_9836);
or U13084 (N_13084,N_8625,N_9906);
or U13085 (N_13085,N_5618,N_6749);
xor U13086 (N_13086,N_6988,N_7351);
or U13087 (N_13087,N_7859,N_9074);
nor U13088 (N_13088,N_5497,N_6854);
xor U13089 (N_13089,N_7966,N_9143);
and U13090 (N_13090,N_5484,N_8673);
xnor U13091 (N_13091,N_6727,N_5371);
nand U13092 (N_13092,N_9333,N_8420);
or U13093 (N_13093,N_6198,N_5014);
xnor U13094 (N_13094,N_7051,N_8028);
or U13095 (N_13095,N_8430,N_8095);
or U13096 (N_13096,N_6419,N_6264);
and U13097 (N_13097,N_9449,N_5038);
nor U13098 (N_13098,N_8256,N_9797);
and U13099 (N_13099,N_6204,N_5654);
xor U13100 (N_13100,N_5851,N_5819);
nand U13101 (N_13101,N_7660,N_6368);
or U13102 (N_13102,N_7259,N_5455);
nand U13103 (N_13103,N_8314,N_5563);
xor U13104 (N_13104,N_5887,N_6999);
and U13105 (N_13105,N_7298,N_7776);
nand U13106 (N_13106,N_7430,N_8803);
nand U13107 (N_13107,N_5937,N_7418);
nor U13108 (N_13108,N_5918,N_6767);
nand U13109 (N_13109,N_8178,N_5006);
nand U13110 (N_13110,N_8588,N_8200);
nor U13111 (N_13111,N_9731,N_6105);
xor U13112 (N_13112,N_6612,N_8723);
nand U13113 (N_13113,N_9123,N_7316);
or U13114 (N_13114,N_6483,N_6708);
nand U13115 (N_13115,N_8576,N_9718);
nor U13116 (N_13116,N_8257,N_9170);
or U13117 (N_13117,N_9116,N_5647);
xnor U13118 (N_13118,N_7679,N_7055);
xnor U13119 (N_13119,N_9342,N_9674);
nand U13120 (N_13120,N_7179,N_7528);
xnor U13121 (N_13121,N_8407,N_5312);
or U13122 (N_13122,N_6688,N_8434);
xnor U13123 (N_13123,N_6822,N_5758);
nand U13124 (N_13124,N_5558,N_9600);
xor U13125 (N_13125,N_9296,N_5920);
xor U13126 (N_13126,N_7878,N_8568);
and U13127 (N_13127,N_8942,N_5424);
or U13128 (N_13128,N_5137,N_8155);
nand U13129 (N_13129,N_5507,N_8059);
and U13130 (N_13130,N_5622,N_9249);
xnor U13131 (N_13131,N_8231,N_6752);
and U13132 (N_13132,N_6587,N_7352);
nand U13133 (N_13133,N_9808,N_5397);
xnor U13134 (N_13134,N_5253,N_9558);
xor U13135 (N_13135,N_9642,N_9491);
or U13136 (N_13136,N_5626,N_5490);
xnor U13137 (N_13137,N_7956,N_9007);
nand U13138 (N_13138,N_8146,N_9110);
and U13139 (N_13139,N_6123,N_8130);
and U13140 (N_13140,N_8577,N_6695);
and U13141 (N_13141,N_8635,N_6692);
and U13142 (N_13142,N_9833,N_7811);
or U13143 (N_13143,N_7415,N_9353);
nand U13144 (N_13144,N_6137,N_7813);
nor U13145 (N_13145,N_8596,N_8368);
and U13146 (N_13146,N_5184,N_5069);
nor U13147 (N_13147,N_6991,N_8849);
nor U13148 (N_13148,N_8041,N_9449);
nor U13149 (N_13149,N_6872,N_5260);
xnor U13150 (N_13150,N_5744,N_9475);
or U13151 (N_13151,N_9372,N_6608);
or U13152 (N_13152,N_6091,N_9571);
or U13153 (N_13153,N_8166,N_8339);
xor U13154 (N_13154,N_9417,N_7939);
nand U13155 (N_13155,N_5820,N_6518);
nand U13156 (N_13156,N_9622,N_7428);
nand U13157 (N_13157,N_5154,N_6076);
and U13158 (N_13158,N_6906,N_5076);
xor U13159 (N_13159,N_7958,N_9208);
and U13160 (N_13160,N_6538,N_6502);
nor U13161 (N_13161,N_8548,N_7042);
or U13162 (N_13162,N_5519,N_6444);
nand U13163 (N_13163,N_6219,N_6658);
nand U13164 (N_13164,N_7451,N_7002);
and U13165 (N_13165,N_5385,N_6716);
nor U13166 (N_13166,N_6247,N_9967);
nand U13167 (N_13167,N_8580,N_7750);
nand U13168 (N_13168,N_9648,N_8789);
or U13169 (N_13169,N_8434,N_8536);
xnor U13170 (N_13170,N_7324,N_8645);
nand U13171 (N_13171,N_9615,N_9075);
or U13172 (N_13172,N_8662,N_8966);
xor U13173 (N_13173,N_5149,N_6195);
xor U13174 (N_13174,N_9602,N_9827);
nor U13175 (N_13175,N_8732,N_9184);
nand U13176 (N_13176,N_8657,N_9987);
nor U13177 (N_13177,N_7706,N_7942);
nand U13178 (N_13178,N_7970,N_5905);
nand U13179 (N_13179,N_8474,N_9715);
or U13180 (N_13180,N_8585,N_6492);
nor U13181 (N_13181,N_6759,N_9525);
or U13182 (N_13182,N_5028,N_7965);
xor U13183 (N_13183,N_7052,N_8724);
or U13184 (N_13184,N_6755,N_9726);
xnor U13185 (N_13185,N_9443,N_7546);
nand U13186 (N_13186,N_6130,N_6618);
and U13187 (N_13187,N_9352,N_6951);
xor U13188 (N_13188,N_6169,N_6801);
xnor U13189 (N_13189,N_7319,N_9522);
nor U13190 (N_13190,N_6239,N_8426);
xor U13191 (N_13191,N_6727,N_9548);
nand U13192 (N_13192,N_8726,N_6038);
nand U13193 (N_13193,N_8253,N_9126);
and U13194 (N_13194,N_7068,N_9580);
xnor U13195 (N_13195,N_6583,N_6356);
or U13196 (N_13196,N_6104,N_6700);
nor U13197 (N_13197,N_6533,N_5737);
xnor U13198 (N_13198,N_9821,N_6762);
nor U13199 (N_13199,N_9089,N_8492);
or U13200 (N_13200,N_8191,N_9404);
and U13201 (N_13201,N_8386,N_8563);
or U13202 (N_13202,N_9381,N_7273);
and U13203 (N_13203,N_6630,N_7173);
xor U13204 (N_13204,N_5127,N_8553);
nand U13205 (N_13205,N_6391,N_6230);
and U13206 (N_13206,N_5816,N_6823);
or U13207 (N_13207,N_5989,N_7879);
or U13208 (N_13208,N_9827,N_5895);
or U13209 (N_13209,N_7957,N_5876);
or U13210 (N_13210,N_6245,N_8705);
nand U13211 (N_13211,N_9956,N_7539);
nor U13212 (N_13212,N_9984,N_7230);
nor U13213 (N_13213,N_5738,N_8799);
and U13214 (N_13214,N_6501,N_7430);
nor U13215 (N_13215,N_9085,N_6386);
xnor U13216 (N_13216,N_6778,N_7492);
nor U13217 (N_13217,N_8701,N_8015);
xor U13218 (N_13218,N_7149,N_7632);
and U13219 (N_13219,N_7439,N_7137);
and U13220 (N_13220,N_7972,N_7753);
nand U13221 (N_13221,N_8942,N_8599);
or U13222 (N_13222,N_8449,N_6965);
nand U13223 (N_13223,N_6424,N_9991);
or U13224 (N_13224,N_9811,N_9248);
nor U13225 (N_13225,N_5895,N_8135);
xor U13226 (N_13226,N_6550,N_6948);
or U13227 (N_13227,N_5282,N_8772);
nand U13228 (N_13228,N_6668,N_9034);
nand U13229 (N_13229,N_5715,N_5212);
or U13230 (N_13230,N_8981,N_8286);
xnor U13231 (N_13231,N_8664,N_5806);
and U13232 (N_13232,N_5997,N_5800);
or U13233 (N_13233,N_5602,N_9764);
xor U13234 (N_13234,N_5934,N_9485);
and U13235 (N_13235,N_8597,N_7985);
nor U13236 (N_13236,N_6327,N_5416);
xnor U13237 (N_13237,N_8153,N_6294);
nor U13238 (N_13238,N_7154,N_7504);
and U13239 (N_13239,N_7386,N_5139);
nor U13240 (N_13240,N_9037,N_5210);
nor U13241 (N_13241,N_6664,N_7102);
or U13242 (N_13242,N_5407,N_8353);
and U13243 (N_13243,N_8024,N_5081);
nor U13244 (N_13244,N_9268,N_8394);
xor U13245 (N_13245,N_9220,N_9296);
and U13246 (N_13246,N_6372,N_6292);
nor U13247 (N_13247,N_6034,N_6933);
or U13248 (N_13248,N_6611,N_9607);
xnor U13249 (N_13249,N_6954,N_6976);
nor U13250 (N_13250,N_8964,N_6739);
xor U13251 (N_13251,N_6299,N_8651);
and U13252 (N_13252,N_5395,N_9558);
and U13253 (N_13253,N_9928,N_7959);
and U13254 (N_13254,N_8266,N_6997);
or U13255 (N_13255,N_6019,N_7282);
and U13256 (N_13256,N_6856,N_9209);
or U13257 (N_13257,N_5256,N_6382);
and U13258 (N_13258,N_6793,N_6102);
nand U13259 (N_13259,N_6756,N_6212);
and U13260 (N_13260,N_8251,N_8254);
and U13261 (N_13261,N_6987,N_8366);
xnor U13262 (N_13262,N_7041,N_9846);
and U13263 (N_13263,N_5300,N_7334);
and U13264 (N_13264,N_8264,N_9977);
and U13265 (N_13265,N_7246,N_5930);
xor U13266 (N_13266,N_8663,N_7710);
xnor U13267 (N_13267,N_6448,N_7979);
xor U13268 (N_13268,N_6974,N_5677);
xnor U13269 (N_13269,N_8047,N_5665);
and U13270 (N_13270,N_6679,N_6746);
xnor U13271 (N_13271,N_8931,N_7108);
or U13272 (N_13272,N_8676,N_5221);
xor U13273 (N_13273,N_8525,N_6104);
and U13274 (N_13274,N_6768,N_8040);
nor U13275 (N_13275,N_6252,N_5211);
xor U13276 (N_13276,N_9019,N_6133);
nand U13277 (N_13277,N_5315,N_5758);
and U13278 (N_13278,N_5583,N_8402);
nand U13279 (N_13279,N_7766,N_8609);
nor U13280 (N_13280,N_5256,N_7870);
nor U13281 (N_13281,N_5382,N_9090);
nor U13282 (N_13282,N_7385,N_5515);
xnor U13283 (N_13283,N_8490,N_8036);
or U13284 (N_13284,N_6001,N_5448);
nand U13285 (N_13285,N_8766,N_5109);
nor U13286 (N_13286,N_8547,N_6310);
xor U13287 (N_13287,N_9622,N_7684);
xor U13288 (N_13288,N_5155,N_9793);
nand U13289 (N_13289,N_6653,N_5654);
nand U13290 (N_13290,N_6450,N_8653);
nand U13291 (N_13291,N_8729,N_8959);
and U13292 (N_13292,N_5359,N_5868);
nor U13293 (N_13293,N_8089,N_8241);
or U13294 (N_13294,N_7771,N_7401);
and U13295 (N_13295,N_8849,N_9155);
nor U13296 (N_13296,N_9169,N_5326);
or U13297 (N_13297,N_7901,N_7054);
nand U13298 (N_13298,N_5467,N_7146);
nor U13299 (N_13299,N_5248,N_5606);
xnor U13300 (N_13300,N_6808,N_9908);
xor U13301 (N_13301,N_8895,N_9392);
nor U13302 (N_13302,N_8722,N_7837);
or U13303 (N_13303,N_6024,N_7833);
nand U13304 (N_13304,N_9092,N_9463);
xnor U13305 (N_13305,N_6976,N_7218);
and U13306 (N_13306,N_9943,N_8828);
nand U13307 (N_13307,N_6320,N_6455);
and U13308 (N_13308,N_7799,N_8359);
and U13309 (N_13309,N_6868,N_5181);
or U13310 (N_13310,N_9680,N_5758);
or U13311 (N_13311,N_5374,N_8206);
nand U13312 (N_13312,N_8238,N_7253);
and U13313 (N_13313,N_9178,N_9290);
or U13314 (N_13314,N_7530,N_6709);
nor U13315 (N_13315,N_9071,N_6987);
or U13316 (N_13316,N_7047,N_6643);
nor U13317 (N_13317,N_9075,N_5697);
and U13318 (N_13318,N_6089,N_6165);
or U13319 (N_13319,N_5899,N_6184);
nand U13320 (N_13320,N_9333,N_7896);
xnor U13321 (N_13321,N_8154,N_5896);
nor U13322 (N_13322,N_5017,N_5710);
and U13323 (N_13323,N_6818,N_9241);
nor U13324 (N_13324,N_8318,N_7458);
xnor U13325 (N_13325,N_5136,N_5402);
xor U13326 (N_13326,N_7434,N_9668);
nand U13327 (N_13327,N_7651,N_6125);
and U13328 (N_13328,N_9457,N_7431);
or U13329 (N_13329,N_9462,N_9578);
xor U13330 (N_13330,N_5271,N_7229);
and U13331 (N_13331,N_9395,N_6252);
nor U13332 (N_13332,N_9616,N_5031);
nand U13333 (N_13333,N_9595,N_6628);
and U13334 (N_13334,N_6125,N_5652);
and U13335 (N_13335,N_5522,N_5125);
or U13336 (N_13336,N_5360,N_8974);
nor U13337 (N_13337,N_5352,N_8104);
or U13338 (N_13338,N_6882,N_6814);
nor U13339 (N_13339,N_7454,N_5347);
xor U13340 (N_13340,N_8009,N_9309);
nor U13341 (N_13341,N_7848,N_7985);
xor U13342 (N_13342,N_9003,N_5751);
nand U13343 (N_13343,N_6509,N_5511);
or U13344 (N_13344,N_7765,N_8540);
or U13345 (N_13345,N_7029,N_7617);
xnor U13346 (N_13346,N_7506,N_9924);
nand U13347 (N_13347,N_8027,N_8842);
nand U13348 (N_13348,N_9020,N_8541);
xnor U13349 (N_13349,N_9858,N_8444);
xnor U13350 (N_13350,N_7026,N_5150);
nor U13351 (N_13351,N_8329,N_7904);
nor U13352 (N_13352,N_9037,N_6824);
and U13353 (N_13353,N_5642,N_7697);
xor U13354 (N_13354,N_7512,N_5069);
or U13355 (N_13355,N_7959,N_7996);
nor U13356 (N_13356,N_5430,N_5716);
xnor U13357 (N_13357,N_7125,N_5458);
and U13358 (N_13358,N_6591,N_5531);
xor U13359 (N_13359,N_5646,N_6457);
nor U13360 (N_13360,N_9515,N_6888);
xnor U13361 (N_13361,N_7446,N_9511);
or U13362 (N_13362,N_6446,N_8980);
or U13363 (N_13363,N_5262,N_9465);
and U13364 (N_13364,N_7852,N_6028);
nor U13365 (N_13365,N_8230,N_8352);
or U13366 (N_13366,N_6889,N_7095);
or U13367 (N_13367,N_5503,N_9035);
nor U13368 (N_13368,N_9611,N_6760);
nor U13369 (N_13369,N_9830,N_8087);
or U13370 (N_13370,N_5381,N_9831);
and U13371 (N_13371,N_6030,N_8052);
and U13372 (N_13372,N_5752,N_9907);
nor U13373 (N_13373,N_6442,N_5720);
or U13374 (N_13374,N_6074,N_5644);
nand U13375 (N_13375,N_6241,N_5483);
and U13376 (N_13376,N_7271,N_6000);
xnor U13377 (N_13377,N_7836,N_6668);
or U13378 (N_13378,N_8435,N_6767);
nor U13379 (N_13379,N_9533,N_8294);
nor U13380 (N_13380,N_9696,N_7914);
nor U13381 (N_13381,N_7169,N_7137);
nand U13382 (N_13382,N_8672,N_9500);
nand U13383 (N_13383,N_8245,N_8208);
nand U13384 (N_13384,N_8171,N_7241);
xnor U13385 (N_13385,N_9112,N_7523);
nand U13386 (N_13386,N_8080,N_5290);
or U13387 (N_13387,N_7832,N_7042);
nand U13388 (N_13388,N_7612,N_6076);
and U13389 (N_13389,N_8056,N_7667);
nor U13390 (N_13390,N_8255,N_7305);
and U13391 (N_13391,N_7517,N_9365);
xnor U13392 (N_13392,N_9057,N_5714);
or U13393 (N_13393,N_5375,N_7214);
xnor U13394 (N_13394,N_7157,N_7035);
nand U13395 (N_13395,N_5551,N_8439);
and U13396 (N_13396,N_8546,N_8610);
xnor U13397 (N_13397,N_6090,N_7573);
xnor U13398 (N_13398,N_9066,N_9763);
or U13399 (N_13399,N_6157,N_5443);
xnor U13400 (N_13400,N_7659,N_5104);
nand U13401 (N_13401,N_7682,N_5697);
and U13402 (N_13402,N_8417,N_8792);
and U13403 (N_13403,N_9287,N_9312);
nand U13404 (N_13404,N_7448,N_7034);
nor U13405 (N_13405,N_8066,N_5850);
nor U13406 (N_13406,N_7541,N_8544);
nand U13407 (N_13407,N_9418,N_9722);
nor U13408 (N_13408,N_9751,N_8795);
and U13409 (N_13409,N_8342,N_8417);
or U13410 (N_13410,N_8497,N_8199);
or U13411 (N_13411,N_7885,N_9536);
xor U13412 (N_13412,N_7933,N_9935);
nor U13413 (N_13413,N_5479,N_6792);
xor U13414 (N_13414,N_9446,N_5682);
nand U13415 (N_13415,N_8725,N_5450);
or U13416 (N_13416,N_6447,N_5897);
xnor U13417 (N_13417,N_6002,N_5532);
nor U13418 (N_13418,N_9151,N_6149);
xor U13419 (N_13419,N_9287,N_7456);
or U13420 (N_13420,N_7145,N_7552);
nor U13421 (N_13421,N_6524,N_9592);
xor U13422 (N_13422,N_6294,N_5474);
and U13423 (N_13423,N_7944,N_9218);
nand U13424 (N_13424,N_5354,N_6958);
or U13425 (N_13425,N_8302,N_5135);
nor U13426 (N_13426,N_8222,N_5882);
and U13427 (N_13427,N_7183,N_5222);
xnor U13428 (N_13428,N_7296,N_9132);
nand U13429 (N_13429,N_9069,N_7864);
xnor U13430 (N_13430,N_8854,N_5796);
xnor U13431 (N_13431,N_6660,N_7845);
and U13432 (N_13432,N_9408,N_8756);
and U13433 (N_13433,N_7202,N_7955);
nand U13434 (N_13434,N_5641,N_5124);
and U13435 (N_13435,N_8753,N_6573);
or U13436 (N_13436,N_9650,N_6658);
and U13437 (N_13437,N_6011,N_8244);
nor U13438 (N_13438,N_7508,N_7390);
xnor U13439 (N_13439,N_9569,N_6328);
xnor U13440 (N_13440,N_6109,N_7937);
nor U13441 (N_13441,N_6665,N_9278);
and U13442 (N_13442,N_7760,N_6487);
or U13443 (N_13443,N_9029,N_8099);
xor U13444 (N_13444,N_7500,N_7664);
xnor U13445 (N_13445,N_8506,N_5331);
nand U13446 (N_13446,N_7618,N_5754);
or U13447 (N_13447,N_9342,N_5371);
nor U13448 (N_13448,N_7232,N_6516);
nor U13449 (N_13449,N_7104,N_6778);
and U13450 (N_13450,N_9501,N_9740);
xor U13451 (N_13451,N_5940,N_9672);
and U13452 (N_13452,N_5954,N_6442);
or U13453 (N_13453,N_5255,N_8396);
or U13454 (N_13454,N_9496,N_6584);
or U13455 (N_13455,N_5587,N_8164);
nor U13456 (N_13456,N_5195,N_6615);
and U13457 (N_13457,N_9878,N_5845);
or U13458 (N_13458,N_8317,N_7326);
and U13459 (N_13459,N_8690,N_8357);
and U13460 (N_13460,N_7120,N_6643);
nor U13461 (N_13461,N_6995,N_6578);
or U13462 (N_13462,N_8317,N_8879);
nor U13463 (N_13463,N_9938,N_7668);
nand U13464 (N_13464,N_7029,N_7882);
xnor U13465 (N_13465,N_9554,N_5208);
and U13466 (N_13466,N_6464,N_6177);
nor U13467 (N_13467,N_9275,N_9390);
nand U13468 (N_13468,N_6350,N_5717);
xnor U13469 (N_13469,N_5461,N_7657);
and U13470 (N_13470,N_8430,N_8650);
xor U13471 (N_13471,N_8500,N_6348);
and U13472 (N_13472,N_7710,N_7509);
nand U13473 (N_13473,N_5562,N_8619);
nor U13474 (N_13474,N_5974,N_8540);
or U13475 (N_13475,N_7830,N_5003);
or U13476 (N_13476,N_6156,N_8138);
and U13477 (N_13477,N_5195,N_5510);
xor U13478 (N_13478,N_6241,N_9971);
and U13479 (N_13479,N_6172,N_6356);
xnor U13480 (N_13480,N_7050,N_7777);
xor U13481 (N_13481,N_9083,N_7471);
nor U13482 (N_13482,N_8088,N_8789);
and U13483 (N_13483,N_8298,N_7002);
and U13484 (N_13484,N_7650,N_6622);
or U13485 (N_13485,N_5590,N_7589);
nor U13486 (N_13486,N_9717,N_9740);
and U13487 (N_13487,N_5448,N_8878);
or U13488 (N_13488,N_5197,N_9039);
or U13489 (N_13489,N_6891,N_9278);
and U13490 (N_13490,N_8462,N_6029);
or U13491 (N_13491,N_6290,N_5710);
or U13492 (N_13492,N_6804,N_5102);
nor U13493 (N_13493,N_5213,N_8053);
xnor U13494 (N_13494,N_7987,N_5012);
xnor U13495 (N_13495,N_9226,N_5085);
nor U13496 (N_13496,N_9062,N_7449);
and U13497 (N_13497,N_7539,N_8738);
and U13498 (N_13498,N_7288,N_8389);
or U13499 (N_13499,N_5181,N_5526);
or U13500 (N_13500,N_7033,N_6898);
xor U13501 (N_13501,N_5338,N_7332);
and U13502 (N_13502,N_7330,N_9734);
and U13503 (N_13503,N_6027,N_8551);
xor U13504 (N_13504,N_8535,N_7698);
nand U13505 (N_13505,N_5864,N_5622);
and U13506 (N_13506,N_6915,N_8744);
or U13507 (N_13507,N_8378,N_5238);
or U13508 (N_13508,N_7496,N_5260);
nor U13509 (N_13509,N_6125,N_6395);
xor U13510 (N_13510,N_6363,N_9869);
nand U13511 (N_13511,N_7888,N_8198);
nand U13512 (N_13512,N_6091,N_5456);
or U13513 (N_13513,N_5137,N_8747);
xnor U13514 (N_13514,N_7684,N_8080);
nand U13515 (N_13515,N_9054,N_6776);
and U13516 (N_13516,N_8466,N_9079);
xor U13517 (N_13517,N_6973,N_8096);
nor U13518 (N_13518,N_8289,N_7260);
and U13519 (N_13519,N_5417,N_8128);
nor U13520 (N_13520,N_9264,N_6166);
or U13521 (N_13521,N_8475,N_9483);
nor U13522 (N_13522,N_6646,N_5794);
xor U13523 (N_13523,N_8142,N_7121);
or U13524 (N_13524,N_5455,N_7390);
and U13525 (N_13525,N_5235,N_7669);
nor U13526 (N_13526,N_9021,N_9675);
xnor U13527 (N_13527,N_7706,N_7672);
nor U13528 (N_13528,N_9380,N_9852);
nand U13529 (N_13529,N_7751,N_6155);
nand U13530 (N_13530,N_5098,N_9862);
xnor U13531 (N_13531,N_6835,N_6817);
xnor U13532 (N_13532,N_7631,N_6905);
and U13533 (N_13533,N_9648,N_6421);
or U13534 (N_13534,N_8962,N_5981);
and U13535 (N_13535,N_8899,N_5385);
nand U13536 (N_13536,N_7348,N_7805);
xnor U13537 (N_13537,N_6370,N_6452);
nor U13538 (N_13538,N_7542,N_9974);
or U13539 (N_13539,N_7633,N_8651);
xor U13540 (N_13540,N_9781,N_8621);
or U13541 (N_13541,N_8166,N_5058);
xor U13542 (N_13542,N_9415,N_9652);
xor U13543 (N_13543,N_9103,N_8494);
nor U13544 (N_13544,N_9945,N_9612);
and U13545 (N_13545,N_7092,N_9660);
nand U13546 (N_13546,N_5625,N_6186);
or U13547 (N_13547,N_9558,N_9190);
nand U13548 (N_13548,N_7305,N_5384);
or U13549 (N_13549,N_7707,N_8022);
or U13550 (N_13550,N_8922,N_7466);
xnor U13551 (N_13551,N_9541,N_8008);
and U13552 (N_13552,N_9213,N_7588);
xor U13553 (N_13553,N_8548,N_6104);
and U13554 (N_13554,N_7185,N_8661);
xor U13555 (N_13555,N_8779,N_7416);
and U13556 (N_13556,N_8959,N_7182);
or U13557 (N_13557,N_5532,N_6279);
nor U13558 (N_13558,N_5292,N_6204);
nor U13559 (N_13559,N_9948,N_7057);
nor U13560 (N_13560,N_6886,N_5488);
nand U13561 (N_13561,N_6000,N_7122);
nor U13562 (N_13562,N_5768,N_6471);
or U13563 (N_13563,N_8012,N_9735);
and U13564 (N_13564,N_8562,N_5661);
nand U13565 (N_13565,N_6178,N_6337);
or U13566 (N_13566,N_7296,N_5666);
xnor U13567 (N_13567,N_6226,N_6058);
xor U13568 (N_13568,N_7324,N_6084);
nor U13569 (N_13569,N_9437,N_6933);
or U13570 (N_13570,N_6575,N_9708);
and U13571 (N_13571,N_7390,N_8313);
or U13572 (N_13572,N_9991,N_9109);
or U13573 (N_13573,N_5514,N_6894);
xnor U13574 (N_13574,N_6862,N_8825);
and U13575 (N_13575,N_6271,N_7352);
and U13576 (N_13576,N_8122,N_5291);
or U13577 (N_13577,N_8307,N_6996);
nand U13578 (N_13578,N_7882,N_6433);
nand U13579 (N_13579,N_9936,N_6966);
nor U13580 (N_13580,N_5478,N_5234);
and U13581 (N_13581,N_8216,N_8603);
nor U13582 (N_13582,N_7819,N_9105);
nor U13583 (N_13583,N_5777,N_7150);
xnor U13584 (N_13584,N_9261,N_7448);
nor U13585 (N_13585,N_8218,N_8726);
or U13586 (N_13586,N_6962,N_8010);
xor U13587 (N_13587,N_8116,N_5554);
or U13588 (N_13588,N_5244,N_5816);
and U13589 (N_13589,N_5673,N_5233);
nand U13590 (N_13590,N_7448,N_9837);
or U13591 (N_13591,N_6815,N_9042);
nand U13592 (N_13592,N_7587,N_8665);
xor U13593 (N_13593,N_8315,N_5157);
xnor U13594 (N_13594,N_7548,N_5517);
nor U13595 (N_13595,N_7525,N_5029);
nand U13596 (N_13596,N_6497,N_9660);
and U13597 (N_13597,N_7712,N_9049);
or U13598 (N_13598,N_6380,N_8771);
and U13599 (N_13599,N_8934,N_6892);
xor U13600 (N_13600,N_9456,N_9656);
nor U13601 (N_13601,N_6961,N_8187);
xor U13602 (N_13602,N_8930,N_6122);
nor U13603 (N_13603,N_8976,N_7081);
or U13604 (N_13604,N_6010,N_5198);
nand U13605 (N_13605,N_8901,N_5009);
nand U13606 (N_13606,N_6416,N_9939);
or U13607 (N_13607,N_6751,N_5473);
xor U13608 (N_13608,N_6727,N_8893);
xor U13609 (N_13609,N_9740,N_5957);
nand U13610 (N_13610,N_6128,N_6928);
xor U13611 (N_13611,N_6240,N_9201);
xor U13612 (N_13612,N_7287,N_6548);
nor U13613 (N_13613,N_7035,N_9277);
or U13614 (N_13614,N_5021,N_5984);
or U13615 (N_13615,N_5494,N_6016);
and U13616 (N_13616,N_9580,N_5536);
and U13617 (N_13617,N_8235,N_7714);
and U13618 (N_13618,N_5193,N_9557);
or U13619 (N_13619,N_6651,N_5523);
nor U13620 (N_13620,N_6571,N_7474);
nor U13621 (N_13621,N_6720,N_5728);
nand U13622 (N_13622,N_7648,N_6755);
xor U13623 (N_13623,N_8302,N_9320);
or U13624 (N_13624,N_6971,N_9649);
nor U13625 (N_13625,N_6905,N_5127);
nand U13626 (N_13626,N_5394,N_5053);
nand U13627 (N_13627,N_6897,N_8110);
nand U13628 (N_13628,N_5571,N_7021);
and U13629 (N_13629,N_6133,N_7336);
xnor U13630 (N_13630,N_5761,N_7076);
nor U13631 (N_13631,N_5590,N_6863);
nand U13632 (N_13632,N_6673,N_9876);
or U13633 (N_13633,N_5331,N_8277);
nand U13634 (N_13634,N_7093,N_9641);
or U13635 (N_13635,N_9403,N_7858);
xor U13636 (N_13636,N_9281,N_8273);
nor U13637 (N_13637,N_7519,N_6542);
nand U13638 (N_13638,N_5036,N_6575);
nand U13639 (N_13639,N_8314,N_9243);
and U13640 (N_13640,N_5073,N_8458);
nand U13641 (N_13641,N_9265,N_5368);
or U13642 (N_13642,N_6273,N_7099);
nor U13643 (N_13643,N_9152,N_7023);
xnor U13644 (N_13644,N_5018,N_7194);
nand U13645 (N_13645,N_6264,N_5516);
xnor U13646 (N_13646,N_6738,N_5962);
and U13647 (N_13647,N_8096,N_7977);
and U13648 (N_13648,N_7919,N_5095);
and U13649 (N_13649,N_8178,N_6077);
and U13650 (N_13650,N_7506,N_6322);
xor U13651 (N_13651,N_9342,N_8675);
nor U13652 (N_13652,N_9633,N_7737);
or U13653 (N_13653,N_9773,N_8310);
and U13654 (N_13654,N_8063,N_8827);
xor U13655 (N_13655,N_6324,N_9303);
and U13656 (N_13656,N_7972,N_7258);
nand U13657 (N_13657,N_6363,N_5085);
or U13658 (N_13658,N_7724,N_9325);
nor U13659 (N_13659,N_9150,N_6399);
or U13660 (N_13660,N_9264,N_5317);
and U13661 (N_13661,N_7598,N_8733);
nand U13662 (N_13662,N_6618,N_9584);
and U13663 (N_13663,N_7921,N_9431);
nor U13664 (N_13664,N_7095,N_5100);
or U13665 (N_13665,N_5816,N_6400);
or U13666 (N_13666,N_6070,N_7087);
or U13667 (N_13667,N_6066,N_7082);
xnor U13668 (N_13668,N_5443,N_6150);
nand U13669 (N_13669,N_7575,N_9495);
nor U13670 (N_13670,N_5346,N_8256);
nor U13671 (N_13671,N_9286,N_8507);
and U13672 (N_13672,N_9463,N_6840);
or U13673 (N_13673,N_9115,N_5411);
nand U13674 (N_13674,N_8978,N_6713);
xor U13675 (N_13675,N_7769,N_8649);
and U13676 (N_13676,N_9959,N_7518);
nor U13677 (N_13677,N_9394,N_6952);
nor U13678 (N_13678,N_9764,N_6859);
nand U13679 (N_13679,N_7219,N_9276);
xnor U13680 (N_13680,N_5813,N_7404);
and U13681 (N_13681,N_8805,N_7784);
xnor U13682 (N_13682,N_6743,N_8851);
nor U13683 (N_13683,N_8285,N_9521);
xor U13684 (N_13684,N_5708,N_8811);
and U13685 (N_13685,N_7231,N_7712);
and U13686 (N_13686,N_8338,N_6637);
nor U13687 (N_13687,N_9145,N_7202);
nand U13688 (N_13688,N_6994,N_7993);
nor U13689 (N_13689,N_5210,N_5057);
nand U13690 (N_13690,N_6827,N_7049);
and U13691 (N_13691,N_9662,N_8283);
and U13692 (N_13692,N_6540,N_8242);
nand U13693 (N_13693,N_7725,N_7548);
nand U13694 (N_13694,N_7571,N_8104);
or U13695 (N_13695,N_7762,N_5686);
and U13696 (N_13696,N_8624,N_7976);
nor U13697 (N_13697,N_5420,N_9701);
xnor U13698 (N_13698,N_5349,N_7662);
nor U13699 (N_13699,N_6006,N_7173);
or U13700 (N_13700,N_5154,N_9028);
and U13701 (N_13701,N_9827,N_5144);
nand U13702 (N_13702,N_6135,N_5768);
nand U13703 (N_13703,N_9305,N_8290);
nand U13704 (N_13704,N_7184,N_9094);
and U13705 (N_13705,N_5690,N_9387);
xor U13706 (N_13706,N_8395,N_8131);
nand U13707 (N_13707,N_6958,N_9631);
xnor U13708 (N_13708,N_5675,N_7273);
nor U13709 (N_13709,N_7207,N_6315);
or U13710 (N_13710,N_8179,N_6947);
nor U13711 (N_13711,N_7610,N_7041);
nor U13712 (N_13712,N_6066,N_5540);
nor U13713 (N_13713,N_6524,N_9587);
or U13714 (N_13714,N_6834,N_8341);
xor U13715 (N_13715,N_9851,N_7592);
nor U13716 (N_13716,N_9580,N_8007);
and U13717 (N_13717,N_5783,N_6755);
xnor U13718 (N_13718,N_6491,N_8308);
and U13719 (N_13719,N_8257,N_7873);
xnor U13720 (N_13720,N_5183,N_6285);
and U13721 (N_13721,N_7998,N_9253);
xor U13722 (N_13722,N_5340,N_5935);
or U13723 (N_13723,N_8458,N_7419);
nor U13724 (N_13724,N_6266,N_6407);
nand U13725 (N_13725,N_7381,N_5424);
and U13726 (N_13726,N_6432,N_5239);
xor U13727 (N_13727,N_8926,N_6109);
or U13728 (N_13728,N_5603,N_9113);
nor U13729 (N_13729,N_9825,N_5540);
nor U13730 (N_13730,N_5306,N_8307);
xor U13731 (N_13731,N_5172,N_9239);
and U13732 (N_13732,N_8041,N_9535);
nor U13733 (N_13733,N_8879,N_7742);
nor U13734 (N_13734,N_8314,N_6122);
and U13735 (N_13735,N_8506,N_7459);
and U13736 (N_13736,N_9852,N_8704);
nor U13737 (N_13737,N_8192,N_6738);
nor U13738 (N_13738,N_8188,N_6932);
or U13739 (N_13739,N_9628,N_5179);
or U13740 (N_13740,N_5919,N_5170);
nand U13741 (N_13741,N_9570,N_7576);
xnor U13742 (N_13742,N_7953,N_8365);
nor U13743 (N_13743,N_7924,N_8922);
xnor U13744 (N_13744,N_9476,N_9215);
xnor U13745 (N_13745,N_9794,N_7988);
and U13746 (N_13746,N_7362,N_7063);
or U13747 (N_13747,N_9378,N_5315);
xor U13748 (N_13748,N_5069,N_7140);
nor U13749 (N_13749,N_8920,N_7975);
nand U13750 (N_13750,N_8942,N_9056);
nand U13751 (N_13751,N_6186,N_8440);
or U13752 (N_13752,N_5173,N_9748);
and U13753 (N_13753,N_8492,N_5726);
or U13754 (N_13754,N_6831,N_9127);
nand U13755 (N_13755,N_5117,N_6216);
xnor U13756 (N_13756,N_8636,N_6873);
or U13757 (N_13757,N_7680,N_5061);
or U13758 (N_13758,N_9802,N_7346);
and U13759 (N_13759,N_7372,N_5719);
nand U13760 (N_13760,N_7199,N_9710);
nand U13761 (N_13761,N_9096,N_9260);
xnor U13762 (N_13762,N_7550,N_8971);
nand U13763 (N_13763,N_7379,N_6097);
nor U13764 (N_13764,N_5016,N_8312);
nor U13765 (N_13765,N_7339,N_6877);
xor U13766 (N_13766,N_6741,N_5398);
xor U13767 (N_13767,N_7721,N_9943);
nor U13768 (N_13768,N_5023,N_9552);
nor U13769 (N_13769,N_9936,N_5439);
or U13770 (N_13770,N_5424,N_7409);
xor U13771 (N_13771,N_8754,N_6431);
nor U13772 (N_13772,N_9965,N_7865);
and U13773 (N_13773,N_6517,N_8278);
or U13774 (N_13774,N_7888,N_9203);
nor U13775 (N_13775,N_7073,N_9375);
or U13776 (N_13776,N_5560,N_9719);
nor U13777 (N_13777,N_5500,N_9758);
xnor U13778 (N_13778,N_6413,N_5281);
nor U13779 (N_13779,N_5671,N_5752);
nor U13780 (N_13780,N_8399,N_8623);
or U13781 (N_13781,N_9081,N_7825);
and U13782 (N_13782,N_8196,N_7885);
and U13783 (N_13783,N_9579,N_8937);
or U13784 (N_13784,N_7555,N_8107);
xnor U13785 (N_13785,N_7404,N_9379);
and U13786 (N_13786,N_7204,N_5450);
nor U13787 (N_13787,N_6358,N_7397);
nor U13788 (N_13788,N_6622,N_6797);
and U13789 (N_13789,N_9770,N_8392);
and U13790 (N_13790,N_5345,N_5016);
xnor U13791 (N_13791,N_8248,N_9796);
and U13792 (N_13792,N_7762,N_6343);
nand U13793 (N_13793,N_7063,N_5576);
and U13794 (N_13794,N_7541,N_7881);
and U13795 (N_13795,N_6046,N_5003);
nor U13796 (N_13796,N_9883,N_8557);
nor U13797 (N_13797,N_5904,N_6678);
xnor U13798 (N_13798,N_6753,N_5947);
or U13799 (N_13799,N_8991,N_8473);
and U13800 (N_13800,N_9323,N_6091);
and U13801 (N_13801,N_8170,N_5920);
nor U13802 (N_13802,N_7954,N_9678);
xnor U13803 (N_13803,N_9338,N_5512);
nand U13804 (N_13804,N_7176,N_9889);
nand U13805 (N_13805,N_5484,N_6854);
and U13806 (N_13806,N_7140,N_6096);
xnor U13807 (N_13807,N_8268,N_8954);
or U13808 (N_13808,N_5409,N_7567);
xor U13809 (N_13809,N_8103,N_6608);
nor U13810 (N_13810,N_5410,N_9850);
or U13811 (N_13811,N_8614,N_8635);
and U13812 (N_13812,N_6906,N_6309);
and U13813 (N_13813,N_9778,N_7388);
xnor U13814 (N_13814,N_9042,N_5183);
or U13815 (N_13815,N_9081,N_7876);
nor U13816 (N_13816,N_6551,N_6083);
nor U13817 (N_13817,N_7707,N_6201);
and U13818 (N_13818,N_6349,N_8656);
and U13819 (N_13819,N_9325,N_6951);
or U13820 (N_13820,N_8786,N_7474);
or U13821 (N_13821,N_5424,N_7267);
or U13822 (N_13822,N_9548,N_9424);
xnor U13823 (N_13823,N_9531,N_6245);
and U13824 (N_13824,N_5370,N_7320);
or U13825 (N_13825,N_7072,N_7400);
nand U13826 (N_13826,N_5995,N_7958);
or U13827 (N_13827,N_6094,N_9936);
or U13828 (N_13828,N_5289,N_9325);
nor U13829 (N_13829,N_6456,N_7689);
nand U13830 (N_13830,N_8123,N_7790);
nor U13831 (N_13831,N_9345,N_6149);
xor U13832 (N_13832,N_6547,N_9164);
or U13833 (N_13833,N_5140,N_9861);
nor U13834 (N_13834,N_5900,N_8899);
nor U13835 (N_13835,N_6510,N_7278);
nor U13836 (N_13836,N_8128,N_6332);
nor U13837 (N_13837,N_8676,N_5091);
or U13838 (N_13838,N_7585,N_5930);
xor U13839 (N_13839,N_8620,N_7874);
nor U13840 (N_13840,N_8701,N_7944);
nor U13841 (N_13841,N_8038,N_9110);
xor U13842 (N_13842,N_7770,N_6163);
or U13843 (N_13843,N_5116,N_5274);
or U13844 (N_13844,N_6453,N_6717);
nand U13845 (N_13845,N_8723,N_9487);
or U13846 (N_13846,N_6376,N_7080);
or U13847 (N_13847,N_8243,N_7836);
nand U13848 (N_13848,N_5040,N_6580);
and U13849 (N_13849,N_8226,N_8014);
nand U13850 (N_13850,N_8174,N_8125);
nand U13851 (N_13851,N_8219,N_6054);
nor U13852 (N_13852,N_8848,N_7662);
xor U13853 (N_13853,N_5011,N_7919);
nand U13854 (N_13854,N_7996,N_5942);
xnor U13855 (N_13855,N_7863,N_6791);
and U13856 (N_13856,N_7477,N_7887);
xnor U13857 (N_13857,N_5143,N_7627);
nand U13858 (N_13858,N_8659,N_6922);
nor U13859 (N_13859,N_9775,N_9387);
and U13860 (N_13860,N_6514,N_5267);
or U13861 (N_13861,N_6573,N_8401);
or U13862 (N_13862,N_5968,N_8694);
xor U13863 (N_13863,N_8295,N_9948);
or U13864 (N_13864,N_5122,N_6246);
xnor U13865 (N_13865,N_7786,N_7882);
nand U13866 (N_13866,N_9171,N_7900);
or U13867 (N_13867,N_5728,N_5067);
and U13868 (N_13868,N_7086,N_6626);
or U13869 (N_13869,N_5016,N_6939);
nor U13870 (N_13870,N_6145,N_7933);
xnor U13871 (N_13871,N_8916,N_7020);
or U13872 (N_13872,N_9767,N_9406);
and U13873 (N_13873,N_9729,N_9181);
nand U13874 (N_13874,N_9916,N_9337);
xnor U13875 (N_13875,N_7605,N_9177);
and U13876 (N_13876,N_5358,N_5013);
and U13877 (N_13877,N_8046,N_8629);
xor U13878 (N_13878,N_9716,N_7073);
nor U13879 (N_13879,N_7850,N_8806);
or U13880 (N_13880,N_7216,N_5237);
and U13881 (N_13881,N_9508,N_9835);
xnor U13882 (N_13882,N_5872,N_8922);
or U13883 (N_13883,N_5175,N_6396);
nand U13884 (N_13884,N_8756,N_9721);
and U13885 (N_13885,N_6776,N_9320);
xnor U13886 (N_13886,N_9265,N_6368);
and U13887 (N_13887,N_7295,N_8576);
nand U13888 (N_13888,N_6526,N_9472);
nand U13889 (N_13889,N_9120,N_9677);
nand U13890 (N_13890,N_6747,N_6568);
nor U13891 (N_13891,N_8221,N_9673);
or U13892 (N_13892,N_8069,N_7948);
nand U13893 (N_13893,N_5552,N_9072);
or U13894 (N_13894,N_9848,N_8682);
and U13895 (N_13895,N_8968,N_5851);
and U13896 (N_13896,N_5785,N_9205);
or U13897 (N_13897,N_8333,N_9018);
nand U13898 (N_13898,N_9411,N_6844);
or U13899 (N_13899,N_6732,N_6961);
and U13900 (N_13900,N_7515,N_6755);
nor U13901 (N_13901,N_8939,N_7301);
nand U13902 (N_13902,N_5075,N_7464);
nor U13903 (N_13903,N_6326,N_6374);
xor U13904 (N_13904,N_8174,N_8259);
nand U13905 (N_13905,N_8415,N_6545);
and U13906 (N_13906,N_8438,N_8289);
nor U13907 (N_13907,N_5867,N_9852);
nor U13908 (N_13908,N_5845,N_9573);
and U13909 (N_13909,N_6243,N_9997);
or U13910 (N_13910,N_8320,N_5739);
xor U13911 (N_13911,N_8668,N_5759);
nand U13912 (N_13912,N_7952,N_6812);
xnor U13913 (N_13913,N_9514,N_5409);
xor U13914 (N_13914,N_9421,N_9458);
or U13915 (N_13915,N_8562,N_6230);
and U13916 (N_13916,N_9563,N_7826);
nor U13917 (N_13917,N_8256,N_8543);
nor U13918 (N_13918,N_8311,N_7305);
nand U13919 (N_13919,N_8872,N_9032);
xor U13920 (N_13920,N_8480,N_5450);
nand U13921 (N_13921,N_6726,N_6176);
nand U13922 (N_13922,N_7198,N_8060);
nand U13923 (N_13923,N_5872,N_9749);
xnor U13924 (N_13924,N_7110,N_9171);
or U13925 (N_13925,N_6894,N_7080);
xnor U13926 (N_13926,N_6303,N_7942);
xor U13927 (N_13927,N_8162,N_8837);
nand U13928 (N_13928,N_9482,N_7895);
nand U13929 (N_13929,N_7995,N_9701);
xnor U13930 (N_13930,N_8262,N_5681);
xor U13931 (N_13931,N_7075,N_5687);
nand U13932 (N_13932,N_9873,N_5090);
and U13933 (N_13933,N_7212,N_5365);
nand U13934 (N_13934,N_7619,N_5268);
nand U13935 (N_13935,N_8738,N_6577);
nor U13936 (N_13936,N_9789,N_7760);
and U13937 (N_13937,N_9283,N_5198);
nor U13938 (N_13938,N_8928,N_5951);
xnor U13939 (N_13939,N_6999,N_6336);
xor U13940 (N_13940,N_5248,N_6985);
or U13941 (N_13941,N_9370,N_9774);
nor U13942 (N_13942,N_8241,N_8161);
and U13943 (N_13943,N_9860,N_9455);
nor U13944 (N_13944,N_8993,N_6263);
xor U13945 (N_13945,N_8294,N_6012);
nand U13946 (N_13946,N_8634,N_8981);
and U13947 (N_13947,N_7422,N_8123);
nor U13948 (N_13948,N_5479,N_7157);
nor U13949 (N_13949,N_9695,N_8991);
nand U13950 (N_13950,N_6603,N_9766);
nand U13951 (N_13951,N_5358,N_5669);
nand U13952 (N_13952,N_5619,N_9584);
xor U13953 (N_13953,N_6666,N_8305);
xnor U13954 (N_13954,N_8934,N_6496);
nand U13955 (N_13955,N_8218,N_5284);
and U13956 (N_13956,N_9565,N_8554);
or U13957 (N_13957,N_5291,N_9619);
xor U13958 (N_13958,N_5580,N_9078);
nand U13959 (N_13959,N_8459,N_5273);
nor U13960 (N_13960,N_9344,N_5039);
xnor U13961 (N_13961,N_9582,N_9471);
nor U13962 (N_13962,N_6110,N_8846);
and U13963 (N_13963,N_5818,N_7744);
or U13964 (N_13964,N_5912,N_6491);
and U13965 (N_13965,N_9574,N_7885);
nor U13966 (N_13966,N_9366,N_6320);
or U13967 (N_13967,N_8134,N_5581);
nand U13968 (N_13968,N_8201,N_8696);
xor U13969 (N_13969,N_8528,N_5722);
or U13970 (N_13970,N_5293,N_5345);
or U13971 (N_13971,N_5197,N_6762);
or U13972 (N_13972,N_6990,N_9581);
and U13973 (N_13973,N_7452,N_5493);
nand U13974 (N_13974,N_5968,N_7125);
nand U13975 (N_13975,N_9665,N_6563);
or U13976 (N_13976,N_6039,N_5131);
nor U13977 (N_13977,N_9060,N_7092);
nand U13978 (N_13978,N_6397,N_5536);
xor U13979 (N_13979,N_6178,N_7110);
nor U13980 (N_13980,N_7902,N_7090);
or U13981 (N_13981,N_9047,N_8620);
nor U13982 (N_13982,N_7761,N_9922);
xnor U13983 (N_13983,N_5455,N_5529);
and U13984 (N_13984,N_7770,N_9595);
or U13985 (N_13985,N_6885,N_5978);
and U13986 (N_13986,N_6780,N_7165);
or U13987 (N_13987,N_9897,N_8303);
and U13988 (N_13988,N_5737,N_7838);
nor U13989 (N_13989,N_6603,N_8696);
or U13990 (N_13990,N_7469,N_9980);
or U13991 (N_13991,N_7753,N_6168);
nand U13992 (N_13992,N_5059,N_5076);
xor U13993 (N_13993,N_7817,N_6856);
xnor U13994 (N_13994,N_6772,N_6031);
nor U13995 (N_13995,N_8274,N_5277);
nand U13996 (N_13996,N_5560,N_6835);
xnor U13997 (N_13997,N_6631,N_5189);
nor U13998 (N_13998,N_6521,N_9232);
nand U13999 (N_13999,N_6364,N_5832);
nand U14000 (N_14000,N_9441,N_7596);
nand U14001 (N_14001,N_9862,N_6550);
or U14002 (N_14002,N_9993,N_7123);
nor U14003 (N_14003,N_8200,N_5607);
nor U14004 (N_14004,N_8629,N_5904);
nand U14005 (N_14005,N_9462,N_9559);
xnor U14006 (N_14006,N_9537,N_5273);
nand U14007 (N_14007,N_7992,N_7694);
and U14008 (N_14008,N_9247,N_8945);
nand U14009 (N_14009,N_9624,N_9242);
nand U14010 (N_14010,N_6477,N_9535);
nand U14011 (N_14011,N_6059,N_9107);
nand U14012 (N_14012,N_8637,N_5600);
and U14013 (N_14013,N_5442,N_5724);
or U14014 (N_14014,N_6111,N_6534);
and U14015 (N_14015,N_8365,N_5916);
nand U14016 (N_14016,N_9708,N_9329);
or U14017 (N_14017,N_5562,N_5879);
nor U14018 (N_14018,N_9536,N_9618);
nand U14019 (N_14019,N_9824,N_9358);
xnor U14020 (N_14020,N_8904,N_8073);
or U14021 (N_14021,N_7415,N_5147);
or U14022 (N_14022,N_6431,N_9866);
or U14023 (N_14023,N_9157,N_9566);
nand U14024 (N_14024,N_5588,N_7012);
nor U14025 (N_14025,N_8507,N_5847);
xor U14026 (N_14026,N_6424,N_6322);
and U14027 (N_14027,N_8168,N_9028);
and U14028 (N_14028,N_5792,N_5942);
xor U14029 (N_14029,N_8428,N_6393);
xnor U14030 (N_14030,N_7682,N_9889);
nand U14031 (N_14031,N_8879,N_6866);
nor U14032 (N_14032,N_9104,N_7004);
and U14033 (N_14033,N_8961,N_8738);
and U14034 (N_14034,N_5124,N_8424);
xnor U14035 (N_14035,N_6882,N_5546);
nand U14036 (N_14036,N_6885,N_7221);
xnor U14037 (N_14037,N_6576,N_7049);
nor U14038 (N_14038,N_9635,N_8682);
or U14039 (N_14039,N_8038,N_5317);
xnor U14040 (N_14040,N_5900,N_7094);
or U14041 (N_14041,N_9257,N_7420);
nor U14042 (N_14042,N_8466,N_9015);
nor U14043 (N_14043,N_8261,N_7818);
xor U14044 (N_14044,N_8258,N_6957);
or U14045 (N_14045,N_9038,N_8265);
nand U14046 (N_14046,N_6160,N_7936);
nor U14047 (N_14047,N_9524,N_6867);
or U14048 (N_14048,N_9692,N_5098);
xnor U14049 (N_14049,N_7172,N_5280);
nor U14050 (N_14050,N_9349,N_9495);
nor U14051 (N_14051,N_8115,N_8746);
nor U14052 (N_14052,N_5847,N_9686);
nand U14053 (N_14053,N_5921,N_9212);
or U14054 (N_14054,N_8856,N_5014);
and U14055 (N_14055,N_5590,N_6357);
and U14056 (N_14056,N_7339,N_7235);
and U14057 (N_14057,N_9398,N_6816);
nand U14058 (N_14058,N_6691,N_6520);
nor U14059 (N_14059,N_6039,N_7040);
or U14060 (N_14060,N_8924,N_6928);
and U14061 (N_14061,N_5927,N_7432);
and U14062 (N_14062,N_5544,N_5026);
and U14063 (N_14063,N_9511,N_8473);
and U14064 (N_14064,N_9639,N_9402);
nand U14065 (N_14065,N_7366,N_8877);
xnor U14066 (N_14066,N_9953,N_7216);
and U14067 (N_14067,N_9317,N_8497);
and U14068 (N_14068,N_9679,N_9734);
xnor U14069 (N_14069,N_5377,N_5042);
xor U14070 (N_14070,N_7630,N_6168);
nor U14071 (N_14071,N_8334,N_8424);
nand U14072 (N_14072,N_7349,N_8377);
and U14073 (N_14073,N_7710,N_8683);
or U14074 (N_14074,N_6673,N_5946);
nor U14075 (N_14075,N_7666,N_5363);
and U14076 (N_14076,N_6946,N_7514);
nor U14077 (N_14077,N_9829,N_5413);
and U14078 (N_14078,N_9063,N_8437);
nand U14079 (N_14079,N_5428,N_6340);
xnor U14080 (N_14080,N_9420,N_7827);
nor U14081 (N_14081,N_8054,N_6161);
xnor U14082 (N_14082,N_5755,N_9635);
nand U14083 (N_14083,N_5169,N_9065);
nor U14084 (N_14084,N_8283,N_5772);
xnor U14085 (N_14085,N_8449,N_6129);
nor U14086 (N_14086,N_5771,N_9192);
nand U14087 (N_14087,N_9948,N_9733);
and U14088 (N_14088,N_9224,N_8068);
xnor U14089 (N_14089,N_6302,N_8025);
nand U14090 (N_14090,N_7633,N_7432);
nand U14091 (N_14091,N_8717,N_7380);
nor U14092 (N_14092,N_7836,N_7623);
and U14093 (N_14093,N_7153,N_9507);
nand U14094 (N_14094,N_8415,N_6821);
nand U14095 (N_14095,N_8767,N_7335);
nand U14096 (N_14096,N_9472,N_8636);
nand U14097 (N_14097,N_6350,N_8260);
or U14098 (N_14098,N_8380,N_7663);
xnor U14099 (N_14099,N_5910,N_5758);
xnor U14100 (N_14100,N_8777,N_6942);
nand U14101 (N_14101,N_8016,N_8698);
nand U14102 (N_14102,N_5278,N_9702);
xor U14103 (N_14103,N_6996,N_5158);
nand U14104 (N_14104,N_9257,N_8275);
or U14105 (N_14105,N_7701,N_9540);
xor U14106 (N_14106,N_6823,N_8190);
or U14107 (N_14107,N_8950,N_5580);
or U14108 (N_14108,N_7596,N_8123);
nand U14109 (N_14109,N_7847,N_8651);
or U14110 (N_14110,N_6822,N_9788);
nand U14111 (N_14111,N_7641,N_9893);
and U14112 (N_14112,N_5872,N_8427);
and U14113 (N_14113,N_6167,N_9242);
xnor U14114 (N_14114,N_5764,N_6273);
nand U14115 (N_14115,N_7579,N_8497);
nor U14116 (N_14116,N_7491,N_7192);
nand U14117 (N_14117,N_7588,N_6213);
and U14118 (N_14118,N_6051,N_5092);
nor U14119 (N_14119,N_8310,N_8593);
xor U14120 (N_14120,N_9942,N_6193);
nand U14121 (N_14121,N_8334,N_6309);
xnor U14122 (N_14122,N_6977,N_8272);
nand U14123 (N_14123,N_5850,N_5199);
nor U14124 (N_14124,N_7309,N_9626);
xnor U14125 (N_14125,N_5641,N_6491);
nand U14126 (N_14126,N_8353,N_9831);
nand U14127 (N_14127,N_7226,N_8488);
or U14128 (N_14128,N_7403,N_6631);
nor U14129 (N_14129,N_7561,N_5336);
xor U14130 (N_14130,N_7888,N_9622);
nor U14131 (N_14131,N_7259,N_9718);
nor U14132 (N_14132,N_6317,N_9071);
and U14133 (N_14133,N_5173,N_8322);
nor U14134 (N_14134,N_7737,N_6790);
and U14135 (N_14135,N_6605,N_7605);
xnor U14136 (N_14136,N_5592,N_9643);
and U14137 (N_14137,N_9153,N_6303);
nand U14138 (N_14138,N_9780,N_7728);
xor U14139 (N_14139,N_9839,N_7962);
nand U14140 (N_14140,N_5451,N_5269);
nand U14141 (N_14141,N_8136,N_5366);
and U14142 (N_14142,N_6361,N_9551);
nor U14143 (N_14143,N_6215,N_6003);
nand U14144 (N_14144,N_6562,N_5225);
and U14145 (N_14145,N_9396,N_7405);
and U14146 (N_14146,N_5334,N_7165);
nor U14147 (N_14147,N_5612,N_9395);
nand U14148 (N_14148,N_5753,N_5454);
xnor U14149 (N_14149,N_7923,N_6777);
xor U14150 (N_14150,N_7558,N_9918);
or U14151 (N_14151,N_6666,N_5271);
or U14152 (N_14152,N_8461,N_8002);
xnor U14153 (N_14153,N_5283,N_6110);
nand U14154 (N_14154,N_7943,N_5094);
nor U14155 (N_14155,N_9603,N_9595);
nand U14156 (N_14156,N_7652,N_7322);
and U14157 (N_14157,N_8893,N_9764);
nand U14158 (N_14158,N_6323,N_8031);
and U14159 (N_14159,N_7441,N_6785);
and U14160 (N_14160,N_6578,N_7679);
and U14161 (N_14161,N_7591,N_5882);
nand U14162 (N_14162,N_7715,N_9643);
nand U14163 (N_14163,N_8703,N_7088);
nand U14164 (N_14164,N_7327,N_5471);
xnor U14165 (N_14165,N_5028,N_9680);
or U14166 (N_14166,N_7343,N_6566);
nand U14167 (N_14167,N_5211,N_8127);
xnor U14168 (N_14168,N_7928,N_6362);
and U14169 (N_14169,N_7467,N_6800);
or U14170 (N_14170,N_7672,N_6682);
and U14171 (N_14171,N_5797,N_9501);
nor U14172 (N_14172,N_9102,N_9577);
and U14173 (N_14173,N_6479,N_5083);
nor U14174 (N_14174,N_8691,N_5557);
or U14175 (N_14175,N_5487,N_6680);
nand U14176 (N_14176,N_6087,N_6125);
nand U14177 (N_14177,N_9075,N_5721);
and U14178 (N_14178,N_7362,N_7841);
nor U14179 (N_14179,N_8433,N_8939);
nand U14180 (N_14180,N_9360,N_7093);
or U14181 (N_14181,N_6027,N_6581);
nor U14182 (N_14182,N_5213,N_7167);
xnor U14183 (N_14183,N_6832,N_6091);
xor U14184 (N_14184,N_6666,N_7907);
xor U14185 (N_14185,N_7736,N_8538);
nor U14186 (N_14186,N_7384,N_5334);
nor U14187 (N_14187,N_8346,N_9683);
nor U14188 (N_14188,N_5544,N_9142);
and U14189 (N_14189,N_5845,N_5948);
nand U14190 (N_14190,N_8389,N_7312);
xor U14191 (N_14191,N_5573,N_5542);
or U14192 (N_14192,N_9909,N_6389);
xnor U14193 (N_14193,N_6815,N_8180);
and U14194 (N_14194,N_8741,N_9367);
nor U14195 (N_14195,N_8152,N_6766);
or U14196 (N_14196,N_9651,N_8612);
nor U14197 (N_14197,N_5228,N_6436);
nor U14198 (N_14198,N_8080,N_5662);
and U14199 (N_14199,N_6197,N_8875);
nor U14200 (N_14200,N_9606,N_8356);
and U14201 (N_14201,N_9000,N_8785);
xor U14202 (N_14202,N_5287,N_9455);
xnor U14203 (N_14203,N_5841,N_6731);
xnor U14204 (N_14204,N_5465,N_9448);
and U14205 (N_14205,N_9078,N_6328);
and U14206 (N_14206,N_8084,N_7436);
nor U14207 (N_14207,N_8740,N_9404);
and U14208 (N_14208,N_8827,N_9835);
nand U14209 (N_14209,N_7031,N_5187);
xor U14210 (N_14210,N_9345,N_8010);
nor U14211 (N_14211,N_7790,N_9075);
xnor U14212 (N_14212,N_7894,N_7721);
or U14213 (N_14213,N_6028,N_9973);
xor U14214 (N_14214,N_7935,N_7103);
and U14215 (N_14215,N_8542,N_6299);
or U14216 (N_14216,N_7381,N_5218);
nor U14217 (N_14217,N_8966,N_5539);
or U14218 (N_14218,N_8985,N_5506);
nor U14219 (N_14219,N_9868,N_9521);
or U14220 (N_14220,N_6946,N_9177);
or U14221 (N_14221,N_5338,N_5521);
xnor U14222 (N_14222,N_8700,N_5804);
nor U14223 (N_14223,N_7478,N_8254);
xor U14224 (N_14224,N_6299,N_5981);
and U14225 (N_14225,N_5106,N_8326);
nand U14226 (N_14226,N_7112,N_6316);
or U14227 (N_14227,N_7194,N_8058);
or U14228 (N_14228,N_9943,N_5157);
nand U14229 (N_14229,N_7590,N_7160);
and U14230 (N_14230,N_9359,N_7174);
nand U14231 (N_14231,N_5133,N_8610);
nand U14232 (N_14232,N_9077,N_9461);
or U14233 (N_14233,N_9606,N_5447);
and U14234 (N_14234,N_6348,N_7141);
and U14235 (N_14235,N_7919,N_8210);
xor U14236 (N_14236,N_5277,N_9380);
nand U14237 (N_14237,N_9864,N_6840);
nand U14238 (N_14238,N_5066,N_6883);
nand U14239 (N_14239,N_7499,N_7368);
and U14240 (N_14240,N_8427,N_5141);
or U14241 (N_14241,N_7118,N_5430);
and U14242 (N_14242,N_6576,N_6807);
nor U14243 (N_14243,N_9700,N_9607);
or U14244 (N_14244,N_5975,N_7380);
nand U14245 (N_14245,N_6970,N_8512);
or U14246 (N_14246,N_6438,N_6908);
and U14247 (N_14247,N_9326,N_9185);
nand U14248 (N_14248,N_8779,N_7810);
xnor U14249 (N_14249,N_6343,N_7697);
nor U14250 (N_14250,N_5311,N_6147);
nand U14251 (N_14251,N_9970,N_8376);
nor U14252 (N_14252,N_7223,N_5757);
nand U14253 (N_14253,N_5434,N_9102);
nor U14254 (N_14254,N_6166,N_6222);
and U14255 (N_14255,N_6048,N_9081);
nor U14256 (N_14256,N_8544,N_9934);
nor U14257 (N_14257,N_7875,N_7333);
or U14258 (N_14258,N_5458,N_5833);
or U14259 (N_14259,N_8261,N_5897);
nor U14260 (N_14260,N_7267,N_7193);
nor U14261 (N_14261,N_9018,N_8058);
and U14262 (N_14262,N_5263,N_6859);
nor U14263 (N_14263,N_6640,N_8941);
xor U14264 (N_14264,N_7016,N_8576);
nand U14265 (N_14265,N_8752,N_7993);
nor U14266 (N_14266,N_7874,N_5638);
xor U14267 (N_14267,N_5447,N_9654);
or U14268 (N_14268,N_7246,N_8088);
xor U14269 (N_14269,N_9183,N_6917);
and U14270 (N_14270,N_5577,N_7324);
xor U14271 (N_14271,N_8778,N_7029);
nor U14272 (N_14272,N_5705,N_7828);
and U14273 (N_14273,N_6624,N_5570);
and U14274 (N_14274,N_9866,N_8236);
nor U14275 (N_14275,N_9249,N_9540);
nand U14276 (N_14276,N_6501,N_6937);
nand U14277 (N_14277,N_9195,N_7017);
nor U14278 (N_14278,N_6228,N_7944);
and U14279 (N_14279,N_5680,N_5452);
xnor U14280 (N_14280,N_6769,N_5460);
xnor U14281 (N_14281,N_7043,N_6826);
nand U14282 (N_14282,N_9681,N_8378);
nor U14283 (N_14283,N_9663,N_5605);
or U14284 (N_14284,N_6664,N_5307);
xor U14285 (N_14285,N_7587,N_8197);
or U14286 (N_14286,N_5957,N_6590);
or U14287 (N_14287,N_6597,N_6698);
or U14288 (N_14288,N_6782,N_6585);
or U14289 (N_14289,N_5218,N_6336);
xor U14290 (N_14290,N_5345,N_5329);
and U14291 (N_14291,N_5888,N_9381);
nor U14292 (N_14292,N_9425,N_7600);
nand U14293 (N_14293,N_8432,N_6844);
nor U14294 (N_14294,N_9521,N_8041);
nand U14295 (N_14295,N_8054,N_5333);
xnor U14296 (N_14296,N_9452,N_5577);
or U14297 (N_14297,N_9124,N_7376);
and U14298 (N_14298,N_5317,N_9493);
nand U14299 (N_14299,N_5754,N_7051);
and U14300 (N_14300,N_7537,N_9172);
xor U14301 (N_14301,N_7747,N_8857);
nand U14302 (N_14302,N_8127,N_6828);
and U14303 (N_14303,N_6716,N_9029);
nor U14304 (N_14304,N_7231,N_9714);
xor U14305 (N_14305,N_6898,N_8479);
xor U14306 (N_14306,N_7778,N_9673);
nor U14307 (N_14307,N_7650,N_5393);
and U14308 (N_14308,N_8081,N_5526);
and U14309 (N_14309,N_7052,N_8387);
and U14310 (N_14310,N_7045,N_9725);
nand U14311 (N_14311,N_5320,N_7535);
nor U14312 (N_14312,N_7391,N_9887);
or U14313 (N_14313,N_8614,N_9492);
and U14314 (N_14314,N_8500,N_5576);
and U14315 (N_14315,N_9297,N_8922);
nor U14316 (N_14316,N_6516,N_9577);
and U14317 (N_14317,N_6249,N_6518);
or U14318 (N_14318,N_8818,N_6017);
or U14319 (N_14319,N_5880,N_8064);
and U14320 (N_14320,N_8320,N_7123);
or U14321 (N_14321,N_5386,N_7737);
xor U14322 (N_14322,N_8380,N_6856);
and U14323 (N_14323,N_7524,N_8146);
xnor U14324 (N_14324,N_9541,N_9153);
and U14325 (N_14325,N_9279,N_8079);
nand U14326 (N_14326,N_7069,N_6708);
xnor U14327 (N_14327,N_8165,N_5963);
nand U14328 (N_14328,N_7140,N_5147);
and U14329 (N_14329,N_6605,N_5464);
nand U14330 (N_14330,N_9718,N_7662);
and U14331 (N_14331,N_9588,N_7930);
nand U14332 (N_14332,N_7643,N_7674);
nand U14333 (N_14333,N_8936,N_6120);
nand U14334 (N_14334,N_9786,N_9226);
and U14335 (N_14335,N_9000,N_7662);
or U14336 (N_14336,N_7322,N_8696);
and U14337 (N_14337,N_6777,N_7726);
xnor U14338 (N_14338,N_9864,N_9793);
nor U14339 (N_14339,N_9680,N_8140);
or U14340 (N_14340,N_6545,N_6619);
nor U14341 (N_14341,N_7915,N_5014);
nand U14342 (N_14342,N_7883,N_5409);
and U14343 (N_14343,N_7319,N_7337);
xnor U14344 (N_14344,N_9016,N_5145);
or U14345 (N_14345,N_6576,N_9285);
and U14346 (N_14346,N_7164,N_6850);
and U14347 (N_14347,N_9429,N_6073);
and U14348 (N_14348,N_9933,N_6741);
or U14349 (N_14349,N_7917,N_5491);
nor U14350 (N_14350,N_9671,N_6024);
nand U14351 (N_14351,N_9528,N_7390);
nand U14352 (N_14352,N_9631,N_7667);
and U14353 (N_14353,N_6072,N_9595);
xor U14354 (N_14354,N_5358,N_8618);
and U14355 (N_14355,N_6411,N_5398);
nor U14356 (N_14356,N_9355,N_9374);
nand U14357 (N_14357,N_5115,N_6441);
or U14358 (N_14358,N_6684,N_5865);
and U14359 (N_14359,N_9864,N_5315);
nor U14360 (N_14360,N_9958,N_9604);
xor U14361 (N_14361,N_6407,N_8390);
xor U14362 (N_14362,N_6795,N_9399);
nand U14363 (N_14363,N_9001,N_6099);
and U14364 (N_14364,N_5696,N_9515);
and U14365 (N_14365,N_5479,N_5111);
nor U14366 (N_14366,N_5858,N_6911);
nor U14367 (N_14367,N_9839,N_6657);
nand U14368 (N_14368,N_5494,N_7217);
xnor U14369 (N_14369,N_5931,N_5118);
and U14370 (N_14370,N_6393,N_9150);
nand U14371 (N_14371,N_9748,N_5762);
or U14372 (N_14372,N_7339,N_9898);
and U14373 (N_14373,N_5149,N_7357);
or U14374 (N_14374,N_6238,N_5888);
nand U14375 (N_14375,N_7241,N_5588);
nand U14376 (N_14376,N_8148,N_9172);
and U14377 (N_14377,N_6164,N_6510);
nor U14378 (N_14378,N_7176,N_5282);
or U14379 (N_14379,N_7251,N_7097);
and U14380 (N_14380,N_7151,N_6130);
or U14381 (N_14381,N_5353,N_8502);
or U14382 (N_14382,N_9117,N_8989);
xnor U14383 (N_14383,N_9820,N_5179);
or U14384 (N_14384,N_7112,N_5334);
and U14385 (N_14385,N_8684,N_6362);
or U14386 (N_14386,N_6937,N_6942);
nor U14387 (N_14387,N_6508,N_9972);
and U14388 (N_14388,N_9986,N_6022);
nand U14389 (N_14389,N_5086,N_8046);
or U14390 (N_14390,N_6283,N_7570);
or U14391 (N_14391,N_8375,N_9527);
xnor U14392 (N_14392,N_6811,N_6152);
nor U14393 (N_14393,N_9861,N_8951);
nand U14394 (N_14394,N_9599,N_8837);
or U14395 (N_14395,N_8473,N_8649);
nand U14396 (N_14396,N_6896,N_6081);
nor U14397 (N_14397,N_5965,N_6265);
nor U14398 (N_14398,N_5557,N_9375);
nor U14399 (N_14399,N_6139,N_6697);
or U14400 (N_14400,N_5130,N_6675);
and U14401 (N_14401,N_8401,N_5525);
nor U14402 (N_14402,N_8869,N_7392);
and U14403 (N_14403,N_9435,N_8941);
nor U14404 (N_14404,N_8116,N_8389);
or U14405 (N_14405,N_8650,N_9492);
nand U14406 (N_14406,N_6158,N_7439);
nand U14407 (N_14407,N_6154,N_7427);
or U14408 (N_14408,N_8379,N_5588);
xor U14409 (N_14409,N_7751,N_5590);
or U14410 (N_14410,N_5983,N_7762);
nor U14411 (N_14411,N_9112,N_5652);
nand U14412 (N_14412,N_5894,N_5099);
or U14413 (N_14413,N_5478,N_5387);
xor U14414 (N_14414,N_7241,N_5952);
and U14415 (N_14415,N_5960,N_6757);
nor U14416 (N_14416,N_5984,N_8189);
nand U14417 (N_14417,N_6835,N_5470);
or U14418 (N_14418,N_7574,N_8377);
or U14419 (N_14419,N_7329,N_5634);
xnor U14420 (N_14420,N_5826,N_9279);
nor U14421 (N_14421,N_8823,N_7734);
and U14422 (N_14422,N_9346,N_8048);
nand U14423 (N_14423,N_7672,N_6889);
xor U14424 (N_14424,N_5258,N_8758);
nand U14425 (N_14425,N_9243,N_6421);
xnor U14426 (N_14426,N_9857,N_6365);
xnor U14427 (N_14427,N_5235,N_5238);
or U14428 (N_14428,N_8097,N_6629);
xor U14429 (N_14429,N_5204,N_6394);
or U14430 (N_14430,N_7646,N_6116);
nor U14431 (N_14431,N_5201,N_7579);
or U14432 (N_14432,N_7893,N_9450);
and U14433 (N_14433,N_8266,N_9867);
xor U14434 (N_14434,N_8025,N_6948);
xnor U14435 (N_14435,N_5702,N_9990);
xnor U14436 (N_14436,N_8134,N_9619);
and U14437 (N_14437,N_6097,N_5834);
nand U14438 (N_14438,N_7671,N_8078);
and U14439 (N_14439,N_7996,N_6034);
xor U14440 (N_14440,N_9271,N_8883);
nor U14441 (N_14441,N_8820,N_6808);
nand U14442 (N_14442,N_8828,N_9375);
and U14443 (N_14443,N_5881,N_6976);
or U14444 (N_14444,N_6276,N_9517);
xnor U14445 (N_14445,N_8202,N_7737);
xor U14446 (N_14446,N_8875,N_5052);
nand U14447 (N_14447,N_8144,N_5588);
or U14448 (N_14448,N_8736,N_7702);
xor U14449 (N_14449,N_8787,N_6770);
and U14450 (N_14450,N_9725,N_5927);
nand U14451 (N_14451,N_6055,N_5204);
nor U14452 (N_14452,N_5836,N_6838);
nand U14453 (N_14453,N_5639,N_7524);
or U14454 (N_14454,N_9215,N_5616);
xnor U14455 (N_14455,N_6286,N_8623);
and U14456 (N_14456,N_5850,N_6595);
nand U14457 (N_14457,N_9058,N_8987);
and U14458 (N_14458,N_6767,N_9910);
xor U14459 (N_14459,N_8741,N_8033);
or U14460 (N_14460,N_8303,N_9494);
xor U14461 (N_14461,N_9762,N_6527);
xor U14462 (N_14462,N_5871,N_7238);
xnor U14463 (N_14463,N_6170,N_9892);
and U14464 (N_14464,N_9698,N_7714);
xnor U14465 (N_14465,N_9921,N_6305);
or U14466 (N_14466,N_5750,N_9156);
and U14467 (N_14467,N_7726,N_9290);
xnor U14468 (N_14468,N_6672,N_7522);
or U14469 (N_14469,N_6007,N_7541);
or U14470 (N_14470,N_6321,N_9560);
or U14471 (N_14471,N_7128,N_5465);
nand U14472 (N_14472,N_5192,N_9704);
nand U14473 (N_14473,N_8924,N_5390);
nor U14474 (N_14474,N_7941,N_5862);
or U14475 (N_14475,N_8413,N_9307);
or U14476 (N_14476,N_9223,N_9198);
and U14477 (N_14477,N_6880,N_8131);
xnor U14478 (N_14478,N_8771,N_9151);
or U14479 (N_14479,N_9078,N_5888);
nand U14480 (N_14480,N_8266,N_6710);
nor U14481 (N_14481,N_8982,N_9233);
nand U14482 (N_14482,N_7426,N_8114);
nor U14483 (N_14483,N_7111,N_5951);
or U14484 (N_14484,N_8534,N_9395);
or U14485 (N_14485,N_9073,N_7757);
xor U14486 (N_14486,N_5444,N_5669);
nor U14487 (N_14487,N_9696,N_9116);
or U14488 (N_14488,N_9163,N_6625);
nor U14489 (N_14489,N_8466,N_7927);
nor U14490 (N_14490,N_5522,N_6978);
nand U14491 (N_14491,N_5762,N_6887);
nand U14492 (N_14492,N_5754,N_9317);
nand U14493 (N_14493,N_8778,N_6369);
and U14494 (N_14494,N_8924,N_6251);
and U14495 (N_14495,N_6009,N_9397);
nor U14496 (N_14496,N_5446,N_9360);
and U14497 (N_14497,N_8693,N_9574);
or U14498 (N_14498,N_8143,N_8387);
or U14499 (N_14499,N_6522,N_5868);
nor U14500 (N_14500,N_7614,N_5293);
xnor U14501 (N_14501,N_9309,N_7822);
or U14502 (N_14502,N_5258,N_6321);
xor U14503 (N_14503,N_9649,N_9399);
and U14504 (N_14504,N_5634,N_5053);
nor U14505 (N_14505,N_9607,N_9775);
or U14506 (N_14506,N_6884,N_5027);
nand U14507 (N_14507,N_8127,N_8214);
or U14508 (N_14508,N_8572,N_8293);
nand U14509 (N_14509,N_6833,N_7073);
xor U14510 (N_14510,N_6136,N_7230);
nor U14511 (N_14511,N_5146,N_5412);
xnor U14512 (N_14512,N_8261,N_7529);
and U14513 (N_14513,N_6946,N_7775);
xnor U14514 (N_14514,N_7562,N_6341);
and U14515 (N_14515,N_7325,N_5527);
xor U14516 (N_14516,N_8123,N_5489);
and U14517 (N_14517,N_9026,N_9894);
nand U14518 (N_14518,N_5320,N_8361);
and U14519 (N_14519,N_6366,N_6163);
nand U14520 (N_14520,N_9763,N_8141);
or U14521 (N_14521,N_6623,N_8756);
or U14522 (N_14522,N_7409,N_6676);
xor U14523 (N_14523,N_6468,N_6786);
xor U14524 (N_14524,N_8638,N_7114);
xnor U14525 (N_14525,N_5898,N_9423);
nor U14526 (N_14526,N_5807,N_5944);
nand U14527 (N_14527,N_7337,N_6980);
xnor U14528 (N_14528,N_7961,N_7396);
nor U14529 (N_14529,N_9930,N_8750);
or U14530 (N_14530,N_9834,N_5188);
nor U14531 (N_14531,N_5460,N_9824);
or U14532 (N_14532,N_7351,N_5868);
and U14533 (N_14533,N_8587,N_6542);
or U14534 (N_14534,N_9437,N_9283);
and U14535 (N_14535,N_7957,N_6848);
nor U14536 (N_14536,N_7325,N_5433);
nand U14537 (N_14537,N_8026,N_7984);
nand U14538 (N_14538,N_5288,N_7165);
and U14539 (N_14539,N_9494,N_7051);
xnor U14540 (N_14540,N_5883,N_7650);
nor U14541 (N_14541,N_9541,N_7517);
nor U14542 (N_14542,N_8351,N_9170);
nand U14543 (N_14543,N_9731,N_5756);
xnor U14544 (N_14544,N_5979,N_5919);
nand U14545 (N_14545,N_7993,N_9729);
nand U14546 (N_14546,N_6410,N_5493);
or U14547 (N_14547,N_7831,N_5803);
nor U14548 (N_14548,N_7507,N_7726);
nor U14549 (N_14549,N_8054,N_6041);
nand U14550 (N_14550,N_9575,N_7999);
nor U14551 (N_14551,N_8660,N_7059);
xnor U14552 (N_14552,N_7727,N_8838);
and U14553 (N_14553,N_9610,N_6261);
and U14554 (N_14554,N_7449,N_7126);
xnor U14555 (N_14555,N_5303,N_8896);
and U14556 (N_14556,N_6922,N_6476);
nor U14557 (N_14557,N_6011,N_5305);
nand U14558 (N_14558,N_9370,N_9888);
or U14559 (N_14559,N_9665,N_7384);
nand U14560 (N_14560,N_5300,N_7161);
nor U14561 (N_14561,N_9272,N_5025);
nand U14562 (N_14562,N_6869,N_6426);
or U14563 (N_14563,N_9943,N_6576);
nor U14564 (N_14564,N_7669,N_9259);
nand U14565 (N_14565,N_6445,N_8544);
xor U14566 (N_14566,N_6372,N_5072);
xnor U14567 (N_14567,N_7386,N_5742);
nor U14568 (N_14568,N_9240,N_9122);
nor U14569 (N_14569,N_5934,N_5697);
nor U14570 (N_14570,N_7132,N_9786);
xnor U14571 (N_14571,N_9736,N_7673);
nand U14572 (N_14572,N_6052,N_9373);
nor U14573 (N_14573,N_5591,N_8616);
nor U14574 (N_14574,N_9736,N_6703);
xnor U14575 (N_14575,N_9281,N_9055);
xnor U14576 (N_14576,N_6873,N_6361);
or U14577 (N_14577,N_8964,N_8471);
and U14578 (N_14578,N_9326,N_9301);
nor U14579 (N_14579,N_7465,N_7239);
nand U14580 (N_14580,N_7529,N_5735);
or U14581 (N_14581,N_9121,N_5819);
and U14582 (N_14582,N_6566,N_8461);
xor U14583 (N_14583,N_7286,N_9525);
nand U14584 (N_14584,N_7720,N_8026);
or U14585 (N_14585,N_8466,N_6450);
and U14586 (N_14586,N_8603,N_6126);
and U14587 (N_14587,N_5292,N_5102);
nand U14588 (N_14588,N_8450,N_9191);
or U14589 (N_14589,N_8799,N_6736);
nor U14590 (N_14590,N_5631,N_8832);
or U14591 (N_14591,N_5904,N_8482);
xnor U14592 (N_14592,N_9095,N_7228);
nor U14593 (N_14593,N_5285,N_8092);
xor U14594 (N_14594,N_9540,N_8438);
or U14595 (N_14595,N_9878,N_5883);
nand U14596 (N_14596,N_7040,N_9724);
xnor U14597 (N_14597,N_9979,N_7888);
and U14598 (N_14598,N_8941,N_9900);
nand U14599 (N_14599,N_9236,N_8436);
nand U14600 (N_14600,N_7716,N_6426);
nor U14601 (N_14601,N_8775,N_6375);
xnor U14602 (N_14602,N_6085,N_7369);
xor U14603 (N_14603,N_8184,N_7020);
nand U14604 (N_14604,N_6733,N_7796);
xor U14605 (N_14605,N_5603,N_7857);
and U14606 (N_14606,N_5670,N_8676);
xnor U14607 (N_14607,N_8662,N_7000);
or U14608 (N_14608,N_5739,N_8751);
xor U14609 (N_14609,N_6576,N_5908);
xnor U14610 (N_14610,N_5537,N_8832);
or U14611 (N_14611,N_9608,N_7719);
nand U14612 (N_14612,N_5546,N_5961);
nand U14613 (N_14613,N_7273,N_8774);
nor U14614 (N_14614,N_9321,N_7030);
and U14615 (N_14615,N_6953,N_9447);
and U14616 (N_14616,N_7252,N_9402);
xor U14617 (N_14617,N_7336,N_6788);
and U14618 (N_14618,N_5351,N_6458);
nand U14619 (N_14619,N_6605,N_6339);
nor U14620 (N_14620,N_5681,N_7192);
xnor U14621 (N_14621,N_6427,N_7688);
nand U14622 (N_14622,N_8557,N_8582);
or U14623 (N_14623,N_9956,N_9950);
nand U14624 (N_14624,N_6304,N_9866);
or U14625 (N_14625,N_8874,N_9175);
xor U14626 (N_14626,N_9549,N_9894);
xor U14627 (N_14627,N_9911,N_7548);
or U14628 (N_14628,N_7831,N_7207);
or U14629 (N_14629,N_9253,N_9503);
and U14630 (N_14630,N_9738,N_9824);
xor U14631 (N_14631,N_5814,N_8117);
nand U14632 (N_14632,N_7841,N_7548);
and U14633 (N_14633,N_8979,N_9203);
or U14634 (N_14634,N_5171,N_6751);
xnor U14635 (N_14635,N_8630,N_5502);
xnor U14636 (N_14636,N_6937,N_7249);
xnor U14637 (N_14637,N_9721,N_7069);
xnor U14638 (N_14638,N_6998,N_7647);
and U14639 (N_14639,N_7597,N_6548);
xor U14640 (N_14640,N_9379,N_6676);
xor U14641 (N_14641,N_7467,N_5060);
nand U14642 (N_14642,N_8019,N_7594);
and U14643 (N_14643,N_6575,N_7927);
xor U14644 (N_14644,N_6511,N_6925);
xnor U14645 (N_14645,N_8332,N_5430);
nor U14646 (N_14646,N_7660,N_7429);
nand U14647 (N_14647,N_6759,N_7213);
nand U14648 (N_14648,N_7757,N_9965);
nand U14649 (N_14649,N_6802,N_6820);
or U14650 (N_14650,N_5191,N_7548);
xor U14651 (N_14651,N_7013,N_9482);
or U14652 (N_14652,N_7273,N_6322);
nor U14653 (N_14653,N_9396,N_6864);
nand U14654 (N_14654,N_7110,N_5657);
and U14655 (N_14655,N_6536,N_5449);
xor U14656 (N_14656,N_7554,N_8730);
and U14657 (N_14657,N_9786,N_9704);
or U14658 (N_14658,N_9715,N_8816);
and U14659 (N_14659,N_9528,N_5555);
nor U14660 (N_14660,N_5481,N_8382);
nand U14661 (N_14661,N_8366,N_7560);
and U14662 (N_14662,N_7003,N_7256);
or U14663 (N_14663,N_6362,N_5256);
nand U14664 (N_14664,N_7260,N_5100);
nand U14665 (N_14665,N_9530,N_7023);
nor U14666 (N_14666,N_5104,N_7321);
nand U14667 (N_14667,N_9954,N_5281);
nor U14668 (N_14668,N_9940,N_5126);
nor U14669 (N_14669,N_6276,N_7701);
xor U14670 (N_14670,N_7916,N_7673);
nor U14671 (N_14671,N_6042,N_5239);
nand U14672 (N_14672,N_7517,N_5559);
or U14673 (N_14673,N_8918,N_6243);
xnor U14674 (N_14674,N_6240,N_6969);
xnor U14675 (N_14675,N_7250,N_9012);
xnor U14676 (N_14676,N_6810,N_7027);
xnor U14677 (N_14677,N_6952,N_6176);
xnor U14678 (N_14678,N_5610,N_5930);
nor U14679 (N_14679,N_7879,N_5665);
xor U14680 (N_14680,N_9354,N_7043);
or U14681 (N_14681,N_8466,N_5110);
or U14682 (N_14682,N_9064,N_7931);
nand U14683 (N_14683,N_6599,N_9091);
and U14684 (N_14684,N_5896,N_7300);
nand U14685 (N_14685,N_7574,N_6354);
or U14686 (N_14686,N_9690,N_9574);
and U14687 (N_14687,N_9086,N_7755);
nor U14688 (N_14688,N_7380,N_8694);
and U14689 (N_14689,N_8883,N_9222);
xnor U14690 (N_14690,N_8713,N_5382);
or U14691 (N_14691,N_7697,N_5164);
nor U14692 (N_14692,N_6049,N_6077);
and U14693 (N_14693,N_7716,N_6863);
or U14694 (N_14694,N_6737,N_7124);
and U14695 (N_14695,N_9039,N_7750);
or U14696 (N_14696,N_6460,N_9911);
xnor U14697 (N_14697,N_8670,N_8531);
and U14698 (N_14698,N_8406,N_9120);
nor U14699 (N_14699,N_8082,N_5319);
xnor U14700 (N_14700,N_7406,N_9974);
nor U14701 (N_14701,N_7696,N_8528);
nand U14702 (N_14702,N_9610,N_7045);
and U14703 (N_14703,N_6894,N_7085);
xor U14704 (N_14704,N_7736,N_9190);
xor U14705 (N_14705,N_6335,N_5051);
or U14706 (N_14706,N_6116,N_8945);
nand U14707 (N_14707,N_5926,N_7026);
nand U14708 (N_14708,N_9702,N_6902);
nand U14709 (N_14709,N_9065,N_6748);
and U14710 (N_14710,N_5717,N_7109);
nor U14711 (N_14711,N_6028,N_9550);
or U14712 (N_14712,N_7117,N_7780);
nand U14713 (N_14713,N_5250,N_5744);
nor U14714 (N_14714,N_5073,N_5583);
or U14715 (N_14715,N_6914,N_7119);
or U14716 (N_14716,N_5263,N_7837);
or U14717 (N_14717,N_9057,N_8042);
nand U14718 (N_14718,N_7244,N_8845);
xnor U14719 (N_14719,N_5768,N_7757);
nand U14720 (N_14720,N_5977,N_7639);
and U14721 (N_14721,N_8602,N_6631);
or U14722 (N_14722,N_7951,N_8801);
nor U14723 (N_14723,N_9955,N_5399);
xnor U14724 (N_14724,N_7282,N_6037);
nand U14725 (N_14725,N_5073,N_8047);
or U14726 (N_14726,N_8471,N_9728);
and U14727 (N_14727,N_9053,N_7379);
nand U14728 (N_14728,N_5561,N_8402);
xor U14729 (N_14729,N_6799,N_7960);
xor U14730 (N_14730,N_5516,N_9151);
nand U14731 (N_14731,N_7486,N_6825);
or U14732 (N_14732,N_8614,N_9930);
or U14733 (N_14733,N_6443,N_8724);
xor U14734 (N_14734,N_8782,N_6857);
and U14735 (N_14735,N_8111,N_5223);
nor U14736 (N_14736,N_8506,N_6611);
nor U14737 (N_14737,N_8952,N_9379);
xor U14738 (N_14738,N_6690,N_7948);
nor U14739 (N_14739,N_5490,N_5470);
or U14740 (N_14740,N_9144,N_8179);
or U14741 (N_14741,N_6221,N_7899);
or U14742 (N_14742,N_7666,N_7483);
xnor U14743 (N_14743,N_8962,N_9249);
or U14744 (N_14744,N_9068,N_5794);
xor U14745 (N_14745,N_6580,N_7705);
xnor U14746 (N_14746,N_6006,N_6209);
or U14747 (N_14747,N_6764,N_6364);
nor U14748 (N_14748,N_5282,N_5185);
or U14749 (N_14749,N_8817,N_7502);
xor U14750 (N_14750,N_5740,N_9337);
and U14751 (N_14751,N_9083,N_8160);
xor U14752 (N_14752,N_6815,N_6183);
nor U14753 (N_14753,N_9130,N_6870);
or U14754 (N_14754,N_5238,N_8256);
and U14755 (N_14755,N_7613,N_8283);
and U14756 (N_14756,N_9291,N_9661);
or U14757 (N_14757,N_7278,N_9570);
xnor U14758 (N_14758,N_7020,N_9451);
xor U14759 (N_14759,N_8407,N_7681);
xor U14760 (N_14760,N_7814,N_8727);
nor U14761 (N_14761,N_8943,N_6367);
nor U14762 (N_14762,N_7233,N_6860);
nor U14763 (N_14763,N_6025,N_7464);
xnor U14764 (N_14764,N_5018,N_8471);
nand U14765 (N_14765,N_6536,N_6859);
nor U14766 (N_14766,N_6889,N_6865);
nand U14767 (N_14767,N_8214,N_9960);
nand U14768 (N_14768,N_5300,N_6046);
xnor U14769 (N_14769,N_7445,N_6505);
xnor U14770 (N_14770,N_7970,N_9972);
xnor U14771 (N_14771,N_6090,N_7158);
xor U14772 (N_14772,N_8178,N_9921);
nand U14773 (N_14773,N_6771,N_7622);
nor U14774 (N_14774,N_7204,N_9909);
nand U14775 (N_14775,N_8925,N_6818);
and U14776 (N_14776,N_8848,N_6618);
nand U14777 (N_14777,N_5758,N_5159);
xor U14778 (N_14778,N_7094,N_6556);
and U14779 (N_14779,N_5466,N_9617);
nor U14780 (N_14780,N_8183,N_5437);
and U14781 (N_14781,N_9937,N_8036);
nor U14782 (N_14782,N_8780,N_9271);
nor U14783 (N_14783,N_9600,N_8168);
or U14784 (N_14784,N_5229,N_9430);
and U14785 (N_14785,N_6732,N_5031);
or U14786 (N_14786,N_8997,N_9401);
xor U14787 (N_14787,N_7521,N_8808);
nor U14788 (N_14788,N_6061,N_6950);
nand U14789 (N_14789,N_5811,N_5846);
xor U14790 (N_14790,N_7517,N_7124);
and U14791 (N_14791,N_9041,N_6323);
nand U14792 (N_14792,N_5618,N_5298);
xnor U14793 (N_14793,N_7510,N_9595);
nor U14794 (N_14794,N_6508,N_6281);
and U14795 (N_14795,N_8341,N_6100);
nor U14796 (N_14796,N_6396,N_5410);
xnor U14797 (N_14797,N_9401,N_6883);
and U14798 (N_14798,N_6521,N_6918);
nand U14799 (N_14799,N_6787,N_9790);
and U14800 (N_14800,N_6587,N_8722);
and U14801 (N_14801,N_8797,N_7356);
xnor U14802 (N_14802,N_9690,N_6060);
nand U14803 (N_14803,N_9831,N_9611);
and U14804 (N_14804,N_6762,N_6252);
nor U14805 (N_14805,N_9432,N_7536);
and U14806 (N_14806,N_9800,N_7008);
nor U14807 (N_14807,N_8366,N_5329);
and U14808 (N_14808,N_5429,N_7856);
nand U14809 (N_14809,N_8268,N_7160);
nor U14810 (N_14810,N_7090,N_8643);
nand U14811 (N_14811,N_5259,N_5564);
xnor U14812 (N_14812,N_7236,N_8659);
nand U14813 (N_14813,N_7351,N_8875);
xor U14814 (N_14814,N_5078,N_8102);
or U14815 (N_14815,N_9739,N_6737);
nand U14816 (N_14816,N_9592,N_8190);
or U14817 (N_14817,N_9702,N_7737);
nor U14818 (N_14818,N_9035,N_5177);
nor U14819 (N_14819,N_6563,N_5211);
nand U14820 (N_14820,N_6679,N_8684);
xnor U14821 (N_14821,N_8139,N_7298);
nor U14822 (N_14822,N_9068,N_5698);
nand U14823 (N_14823,N_5713,N_8471);
and U14824 (N_14824,N_7092,N_8404);
nor U14825 (N_14825,N_9584,N_6063);
xnor U14826 (N_14826,N_8501,N_5407);
nor U14827 (N_14827,N_8132,N_8486);
or U14828 (N_14828,N_6718,N_8535);
nor U14829 (N_14829,N_9148,N_6992);
and U14830 (N_14830,N_9927,N_7651);
nand U14831 (N_14831,N_7721,N_5841);
and U14832 (N_14832,N_7961,N_6492);
nand U14833 (N_14833,N_8080,N_6697);
xor U14834 (N_14834,N_6824,N_9057);
or U14835 (N_14835,N_7549,N_8821);
xor U14836 (N_14836,N_7912,N_7018);
and U14837 (N_14837,N_5442,N_8705);
nand U14838 (N_14838,N_7954,N_5657);
and U14839 (N_14839,N_5524,N_8853);
nand U14840 (N_14840,N_8899,N_7445);
and U14841 (N_14841,N_7243,N_7013);
xor U14842 (N_14842,N_8587,N_7168);
or U14843 (N_14843,N_8092,N_6197);
nor U14844 (N_14844,N_5472,N_6123);
and U14845 (N_14845,N_5402,N_6343);
or U14846 (N_14846,N_5722,N_7572);
nor U14847 (N_14847,N_9194,N_8507);
and U14848 (N_14848,N_9884,N_8659);
nor U14849 (N_14849,N_6018,N_8450);
and U14850 (N_14850,N_8848,N_8601);
xnor U14851 (N_14851,N_8288,N_8996);
or U14852 (N_14852,N_7470,N_5918);
or U14853 (N_14853,N_7219,N_6264);
xnor U14854 (N_14854,N_7733,N_7357);
nand U14855 (N_14855,N_9911,N_8995);
and U14856 (N_14856,N_8331,N_7103);
or U14857 (N_14857,N_7863,N_9258);
nand U14858 (N_14858,N_7158,N_8703);
nor U14859 (N_14859,N_9317,N_8862);
xor U14860 (N_14860,N_6414,N_7641);
nand U14861 (N_14861,N_7666,N_5712);
nor U14862 (N_14862,N_6506,N_5197);
nand U14863 (N_14863,N_9724,N_7305);
nor U14864 (N_14864,N_9877,N_7641);
nor U14865 (N_14865,N_6505,N_8042);
nor U14866 (N_14866,N_9273,N_5803);
or U14867 (N_14867,N_9098,N_8384);
xor U14868 (N_14868,N_7075,N_8571);
xor U14869 (N_14869,N_5779,N_8328);
or U14870 (N_14870,N_9938,N_5549);
nand U14871 (N_14871,N_8669,N_5922);
or U14872 (N_14872,N_5901,N_7203);
or U14873 (N_14873,N_6220,N_5689);
nand U14874 (N_14874,N_7379,N_8457);
or U14875 (N_14875,N_9424,N_7023);
or U14876 (N_14876,N_5604,N_7443);
xnor U14877 (N_14877,N_9028,N_6148);
or U14878 (N_14878,N_9633,N_7946);
or U14879 (N_14879,N_7572,N_5069);
xnor U14880 (N_14880,N_7392,N_5029);
nor U14881 (N_14881,N_5894,N_5037);
and U14882 (N_14882,N_7334,N_5870);
and U14883 (N_14883,N_6515,N_8340);
nand U14884 (N_14884,N_9204,N_9654);
nand U14885 (N_14885,N_8321,N_9117);
or U14886 (N_14886,N_7084,N_9470);
or U14887 (N_14887,N_8415,N_6197);
and U14888 (N_14888,N_8993,N_6546);
and U14889 (N_14889,N_8888,N_8547);
or U14890 (N_14890,N_5207,N_8547);
and U14891 (N_14891,N_7020,N_9972);
or U14892 (N_14892,N_6019,N_5360);
xor U14893 (N_14893,N_6307,N_5855);
nor U14894 (N_14894,N_6177,N_8298);
and U14895 (N_14895,N_7887,N_6367);
or U14896 (N_14896,N_7662,N_9796);
nand U14897 (N_14897,N_5876,N_7764);
nor U14898 (N_14898,N_7207,N_6917);
nand U14899 (N_14899,N_6732,N_8071);
xor U14900 (N_14900,N_9645,N_7761);
and U14901 (N_14901,N_5690,N_6914);
xor U14902 (N_14902,N_8009,N_5988);
nor U14903 (N_14903,N_6706,N_7520);
nor U14904 (N_14904,N_5691,N_9384);
and U14905 (N_14905,N_9190,N_7118);
nand U14906 (N_14906,N_5599,N_5562);
xnor U14907 (N_14907,N_7055,N_6894);
nand U14908 (N_14908,N_5442,N_9327);
nand U14909 (N_14909,N_7644,N_8836);
or U14910 (N_14910,N_8682,N_9951);
or U14911 (N_14911,N_7270,N_9019);
nand U14912 (N_14912,N_6428,N_6469);
nand U14913 (N_14913,N_5439,N_7516);
xnor U14914 (N_14914,N_5465,N_6749);
or U14915 (N_14915,N_9802,N_5650);
nor U14916 (N_14916,N_7770,N_9996);
or U14917 (N_14917,N_9729,N_7620);
nand U14918 (N_14918,N_7432,N_8103);
and U14919 (N_14919,N_9266,N_6295);
or U14920 (N_14920,N_5396,N_7672);
or U14921 (N_14921,N_7420,N_8352);
nand U14922 (N_14922,N_9007,N_8567);
and U14923 (N_14923,N_7752,N_7211);
and U14924 (N_14924,N_8976,N_5701);
xnor U14925 (N_14925,N_5797,N_9585);
and U14926 (N_14926,N_5021,N_7830);
and U14927 (N_14927,N_9029,N_9499);
and U14928 (N_14928,N_5898,N_7978);
nor U14929 (N_14929,N_9744,N_9432);
and U14930 (N_14930,N_9128,N_9422);
and U14931 (N_14931,N_9544,N_9685);
nor U14932 (N_14932,N_7391,N_9402);
xor U14933 (N_14933,N_9693,N_8453);
and U14934 (N_14934,N_9133,N_8881);
and U14935 (N_14935,N_9329,N_9465);
xnor U14936 (N_14936,N_5303,N_6100);
xnor U14937 (N_14937,N_6575,N_5914);
xor U14938 (N_14938,N_8887,N_9356);
and U14939 (N_14939,N_5434,N_6367);
nor U14940 (N_14940,N_5423,N_6169);
xnor U14941 (N_14941,N_6564,N_9114);
or U14942 (N_14942,N_7060,N_8238);
or U14943 (N_14943,N_5053,N_8457);
nor U14944 (N_14944,N_9483,N_6396);
nand U14945 (N_14945,N_9995,N_7109);
nand U14946 (N_14946,N_9851,N_8021);
and U14947 (N_14947,N_6522,N_7128);
nand U14948 (N_14948,N_8352,N_5377);
or U14949 (N_14949,N_6073,N_9110);
nor U14950 (N_14950,N_5163,N_9832);
nand U14951 (N_14951,N_8442,N_9750);
nor U14952 (N_14952,N_9222,N_8418);
nand U14953 (N_14953,N_6346,N_8749);
and U14954 (N_14954,N_8814,N_7544);
or U14955 (N_14955,N_7754,N_9686);
xor U14956 (N_14956,N_6151,N_8207);
nand U14957 (N_14957,N_6447,N_6591);
xnor U14958 (N_14958,N_6318,N_7345);
xor U14959 (N_14959,N_7754,N_9366);
and U14960 (N_14960,N_6011,N_7043);
or U14961 (N_14961,N_6733,N_9456);
and U14962 (N_14962,N_9122,N_7003);
or U14963 (N_14963,N_6937,N_8045);
nand U14964 (N_14964,N_9849,N_6430);
or U14965 (N_14965,N_9748,N_8939);
xor U14966 (N_14966,N_8104,N_7215);
xor U14967 (N_14967,N_5256,N_9640);
nor U14968 (N_14968,N_5067,N_5052);
or U14969 (N_14969,N_9457,N_6148);
and U14970 (N_14970,N_8355,N_6257);
nand U14971 (N_14971,N_5311,N_8509);
nor U14972 (N_14972,N_7009,N_9881);
nor U14973 (N_14973,N_5678,N_6198);
nor U14974 (N_14974,N_5969,N_9113);
nand U14975 (N_14975,N_7621,N_8575);
and U14976 (N_14976,N_6265,N_9849);
and U14977 (N_14977,N_7378,N_8949);
nor U14978 (N_14978,N_5574,N_5672);
or U14979 (N_14979,N_6533,N_9146);
and U14980 (N_14980,N_6891,N_9698);
nand U14981 (N_14981,N_7396,N_7178);
or U14982 (N_14982,N_9631,N_6276);
or U14983 (N_14983,N_6602,N_8172);
nor U14984 (N_14984,N_6163,N_8488);
xor U14985 (N_14985,N_7792,N_6940);
nand U14986 (N_14986,N_5648,N_6151);
xor U14987 (N_14987,N_8810,N_6966);
and U14988 (N_14988,N_8303,N_5166);
and U14989 (N_14989,N_7118,N_7281);
nor U14990 (N_14990,N_9004,N_9582);
and U14991 (N_14991,N_5971,N_9650);
or U14992 (N_14992,N_8697,N_5926);
nand U14993 (N_14993,N_9917,N_8245);
nand U14994 (N_14994,N_9760,N_7434);
nor U14995 (N_14995,N_5982,N_8239);
xor U14996 (N_14996,N_6602,N_6982);
nand U14997 (N_14997,N_8752,N_7274);
or U14998 (N_14998,N_8533,N_8104);
nor U14999 (N_14999,N_6926,N_7530);
xnor UO_0 (O_0,N_11569,N_11917);
nand UO_1 (O_1,N_11904,N_12592);
nand UO_2 (O_2,N_12491,N_14436);
and UO_3 (O_3,N_13682,N_12832);
nor UO_4 (O_4,N_12850,N_11892);
and UO_5 (O_5,N_10940,N_13679);
nand UO_6 (O_6,N_10262,N_13966);
or UO_7 (O_7,N_13203,N_10395);
and UO_8 (O_8,N_12616,N_13710);
nand UO_9 (O_9,N_13736,N_11238);
xor UO_10 (O_10,N_13819,N_13111);
or UO_11 (O_11,N_12101,N_14506);
nor UO_12 (O_12,N_12293,N_10867);
xnor UO_13 (O_13,N_10035,N_11414);
and UO_14 (O_14,N_14120,N_11761);
nor UO_15 (O_15,N_14907,N_10996);
or UO_16 (O_16,N_11242,N_13668);
nand UO_17 (O_17,N_10757,N_12302);
or UO_18 (O_18,N_13512,N_11618);
nand UO_19 (O_19,N_11979,N_13505);
nor UO_20 (O_20,N_12141,N_12579);
and UO_21 (O_21,N_13055,N_11263);
nand UO_22 (O_22,N_14579,N_10082);
nand UO_23 (O_23,N_11289,N_14653);
and UO_24 (O_24,N_11161,N_13591);
xor UO_25 (O_25,N_10069,N_10010);
or UO_26 (O_26,N_10654,N_12793);
and UO_27 (O_27,N_11119,N_14466);
or UO_28 (O_28,N_13635,N_12968);
and UO_29 (O_29,N_14193,N_12905);
nand UO_30 (O_30,N_12677,N_11360);
xor UO_31 (O_31,N_14324,N_13684);
xor UO_32 (O_32,N_11304,N_10397);
xnor UO_33 (O_33,N_14530,N_10812);
and UO_34 (O_34,N_14394,N_10599);
or UO_35 (O_35,N_10085,N_14887);
nor UO_36 (O_36,N_13413,N_11902);
and UO_37 (O_37,N_10388,N_10333);
and UO_38 (O_38,N_13261,N_12947);
and UO_39 (O_39,N_10235,N_14450);
nand UO_40 (O_40,N_10206,N_11947);
and UO_41 (O_41,N_10194,N_10128);
and UO_42 (O_42,N_14238,N_13594);
nand UO_43 (O_43,N_10529,N_14137);
and UO_44 (O_44,N_11053,N_14978);
and UO_45 (O_45,N_13890,N_14667);
or UO_46 (O_46,N_13839,N_12385);
and UO_47 (O_47,N_11872,N_13030);
and UO_48 (O_48,N_14452,N_11668);
nand UO_49 (O_49,N_11122,N_11937);
or UO_50 (O_50,N_10585,N_11527);
nor UO_51 (O_51,N_11550,N_14453);
nor UO_52 (O_52,N_13639,N_12812);
or UO_53 (O_53,N_11339,N_11357);
and UO_54 (O_54,N_13297,N_14401);
and UO_55 (O_55,N_11004,N_14036);
nand UO_56 (O_56,N_10335,N_14400);
xor UO_57 (O_57,N_14379,N_13584);
and UO_58 (O_58,N_12696,N_11154);
or UO_59 (O_59,N_11028,N_14859);
nor UO_60 (O_60,N_14921,N_10287);
or UO_61 (O_61,N_12545,N_14178);
xor UO_62 (O_62,N_14589,N_12815);
or UO_63 (O_63,N_13442,N_14097);
nor UO_64 (O_64,N_11977,N_14699);
and UO_65 (O_65,N_14177,N_10848);
and UO_66 (O_66,N_14834,N_12037);
and UO_67 (O_67,N_12874,N_11852);
or UO_68 (O_68,N_11525,N_11388);
or UO_69 (O_69,N_14256,N_12719);
nand UO_70 (O_70,N_14685,N_10296);
nor UO_71 (O_71,N_13405,N_12788);
xor UO_72 (O_72,N_10248,N_11547);
nand UO_73 (O_73,N_14272,N_14486);
and UO_74 (O_74,N_11553,N_13994);
nor UO_75 (O_75,N_12589,N_13655);
nor UO_76 (O_76,N_11658,N_13555);
nor UO_77 (O_77,N_11214,N_13697);
and UO_78 (O_78,N_11196,N_14729);
xor UO_79 (O_79,N_10066,N_14337);
nor UO_80 (O_80,N_11922,N_14476);
xor UO_81 (O_81,N_12442,N_12980);
and UO_82 (O_82,N_10143,N_10096);
nor UO_83 (O_83,N_13798,N_14415);
or UO_84 (O_84,N_14388,N_12537);
or UO_85 (O_85,N_14107,N_13135);
xor UO_86 (O_86,N_14756,N_10794);
xor UO_87 (O_87,N_12889,N_13763);
or UO_88 (O_88,N_11563,N_12052);
or UO_89 (O_89,N_14084,N_11801);
and UO_90 (O_90,N_12103,N_14791);
or UO_91 (O_91,N_12391,N_10298);
nand UO_92 (O_92,N_13676,N_10034);
or UO_93 (O_93,N_14246,N_13832);
nor UO_94 (O_94,N_12048,N_14134);
and UO_95 (O_95,N_10583,N_13440);
xor UO_96 (O_96,N_10663,N_11866);
and UO_97 (O_97,N_11725,N_10134);
or UO_98 (O_98,N_13120,N_11058);
nor UO_99 (O_99,N_14396,N_10856);
nand UO_100 (O_100,N_13992,N_12483);
xnor UO_101 (O_101,N_11423,N_10191);
and UO_102 (O_102,N_14736,N_12301);
and UO_103 (O_103,N_14289,N_12256);
or UO_104 (O_104,N_10019,N_14033);
xor UO_105 (O_105,N_14469,N_11212);
nor UO_106 (O_106,N_12329,N_13772);
xnor UO_107 (O_107,N_14207,N_13737);
or UO_108 (O_108,N_11613,N_12575);
xor UO_109 (O_109,N_10293,N_10595);
and UO_110 (O_110,N_11216,N_10197);
nand UO_111 (O_111,N_10377,N_14612);
nor UO_112 (O_112,N_13378,N_14173);
nor UO_113 (O_113,N_14360,N_10324);
nand UO_114 (O_114,N_14230,N_10633);
or UO_115 (O_115,N_13127,N_12472);
nor UO_116 (O_116,N_11069,N_14763);
and UO_117 (O_117,N_12215,N_12928);
xnor UO_118 (O_118,N_10215,N_12540);
nor UO_119 (O_119,N_14815,N_14471);
nor UO_120 (O_120,N_13983,N_11452);
xor UO_121 (O_121,N_13702,N_13437);
nand UO_122 (O_122,N_12739,N_14662);
xor UO_123 (O_123,N_10227,N_11193);
and UO_124 (O_124,N_13567,N_13921);
nand UO_125 (O_125,N_11070,N_14406);
and UO_126 (O_126,N_12717,N_14595);
and UO_127 (O_127,N_14397,N_10301);
nand UO_128 (O_128,N_14239,N_12386);
nor UO_129 (O_129,N_14587,N_14100);
and UO_130 (O_130,N_10652,N_13291);
xnor UO_131 (O_131,N_11935,N_10171);
xnor UO_132 (O_132,N_14333,N_14941);
or UO_133 (O_133,N_12756,N_13404);
or UO_134 (O_134,N_11641,N_11941);
and UO_135 (O_135,N_11308,N_13428);
and UO_136 (O_136,N_11011,N_12480);
and UO_137 (O_137,N_11996,N_11392);
or UO_138 (O_138,N_14515,N_10712);
or UO_139 (O_139,N_14703,N_11634);
xor UO_140 (O_140,N_11739,N_12692);
or UO_141 (O_141,N_13875,N_10450);
or UO_142 (O_142,N_11012,N_12174);
xnor UO_143 (O_143,N_14690,N_11631);
and UO_144 (O_144,N_14484,N_13742);
nand UO_145 (O_145,N_14868,N_13731);
xor UO_146 (O_146,N_11187,N_13276);
nand UO_147 (O_147,N_10063,N_14569);
xnor UO_148 (O_148,N_11397,N_11818);
xnor UO_149 (O_149,N_13285,N_10951);
xor UO_150 (O_150,N_11967,N_13166);
or UO_151 (O_151,N_13776,N_12962);
nand UO_152 (O_152,N_13878,N_13387);
nor UO_153 (O_153,N_14660,N_10164);
nor UO_154 (O_154,N_14755,N_10681);
xor UO_155 (O_155,N_13959,N_12118);
nor UO_156 (O_156,N_14295,N_12171);
or UO_157 (O_157,N_10821,N_14762);
nor UO_158 (O_158,N_13650,N_12210);
xor UO_159 (O_159,N_14061,N_14420);
nor UO_160 (O_160,N_12789,N_12276);
nor UO_161 (O_161,N_14414,N_14386);
or UO_162 (O_162,N_10132,N_14551);
nor UO_163 (O_163,N_11176,N_12794);
or UO_164 (O_164,N_13495,N_10680);
xor UO_165 (O_165,N_11603,N_14108);
xor UO_166 (O_166,N_10793,N_12202);
nor UO_167 (O_167,N_11315,N_14204);
and UO_168 (O_168,N_12955,N_10444);
nand UO_169 (O_169,N_11548,N_11561);
or UO_170 (O_170,N_10523,N_11504);
xnor UO_171 (O_171,N_14366,N_11375);
xor UO_172 (O_172,N_13636,N_11110);
nor UO_173 (O_173,N_14816,N_10609);
nor UO_174 (O_174,N_14681,N_14540);
or UO_175 (O_175,N_12338,N_10512);
nor UO_176 (O_176,N_14116,N_12003);
or UO_177 (O_177,N_14838,N_12957);
and UO_178 (O_178,N_13333,N_14268);
or UO_179 (O_179,N_10564,N_10541);
and UO_180 (O_180,N_10543,N_11178);
xnor UO_181 (O_181,N_13546,N_13938);
and UO_182 (O_182,N_11476,N_11830);
nand UO_183 (O_183,N_14087,N_12478);
xnor UO_184 (O_184,N_12180,N_11773);
and UO_185 (O_185,N_12590,N_12194);
nor UO_186 (O_186,N_11426,N_14675);
nand UO_187 (O_187,N_14810,N_11072);
nand UO_188 (O_188,N_11073,N_10931);
or UO_189 (O_189,N_11523,N_13029);
or UO_190 (O_190,N_12969,N_11629);
nand UO_191 (O_191,N_12308,N_14898);
nor UO_192 (O_192,N_11568,N_11259);
and UO_193 (O_193,N_13849,N_13811);
nor UO_194 (O_194,N_10190,N_10698);
or UO_195 (O_195,N_14335,N_12211);
xor UO_196 (O_196,N_11298,N_14535);
and UO_197 (O_197,N_10159,N_12001);
or UO_198 (O_198,N_12148,N_11281);
or UO_199 (O_199,N_12017,N_13319);
nand UO_200 (O_200,N_14021,N_11027);
and UO_201 (O_201,N_13057,N_11016);
xnor UO_202 (O_202,N_11148,N_14732);
xor UO_203 (O_203,N_13824,N_12071);
nand UO_204 (O_204,N_11436,N_14096);
or UO_205 (O_205,N_14947,N_12383);
or UO_206 (O_206,N_10346,N_11978);
nor UO_207 (O_207,N_11457,N_11647);
or UO_208 (O_208,N_11897,N_12979);
or UO_209 (O_209,N_11555,N_11348);
nor UO_210 (O_210,N_13598,N_11177);
xnor UO_211 (O_211,N_14411,N_14646);
nor UO_212 (O_212,N_12820,N_13328);
xor UO_213 (O_213,N_11734,N_11743);
or UO_214 (O_214,N_13993,N_13916);
nor UO_215 (O_215,N_14554,N_13637);
nand UO_216 (O_216,N_11047,N_12565);
or UO_217 (O_217,N_14012,N_12923);
xor UO_218 (O_218,N_10135,N_10314);
and UO_219 (O_219,N_10524,N_11326);
xor UO_220 (O_220,N_12417,N_12636);
nand UO_221 (O_221,N_11565,N_13515);
and UO_222 (O_222,N_12411,N_12662);
nand UO_223 (O_223,N_12223,N_11080);
xor UO_224 (O_224,N_10386,N_10258);
and UO_225 (O_225,N_14369,N_14320);
or UO_226 (O_226,N_14191,N_12577);
and UO_227 (O_227,N_11284,N_11685);
nor UO_228 (O_228,N_10608,N_10003);
and UO_229 (O_229,N_10363,N_11735);
nor UO_230 (O_230,N_11522,N_14648);
nand UO_231 (O_231,N_10222,N_13686);
and UO_232 (O_232,N_10101,N_12305);
or UO_233 (O_233,N_10869,N_11919);
and UO_234 (O_234,N_14521,N_12498);
and UO_235 (O_235,N_11964,N_10038);
and UO_236 (O_236,N_11770,N_13096);
xnor UO_237 (O_237,N_13094,N_14505);
xor UO_238 (O_238,N_10705,N_10221);
nand UO_239 (O_239,N_11240,N_11573);
nand UO_240 (O_240,N_12368,N_13544);
and UO_241 (O_241,N_13420,N_12224);
and UO_242 (O_242,N_12437,N_10955);
xor UO_243 (O_243,N_11768,N_12314);
or UO_244 (O_244,N_14404,N_11994);
and UO_245 (O_245,N_12586,N_12904);
xnor UO_246 (O_246,N_13012,N_11387);
nand UO_247 (O_247,N_11912,N_12169);
or UO_248 (O_248,N_11230,N_14291);
and UO_249 (O_249,N_14070,N_11552);
xnor UO_250 (O_250,N_13603,N_10310);
xnor UO_251 (O_251,N_10774,N_13060);
nand UO_252 (O_252,N_13287,N_13517);
and UO_253 (O_253,N_10497,N_11929);
xor UO_254 (O_254,N_10274,N_11086);
and UO_255 (O_255,N_10791,N_12819);
nand UO_256 (O_256,N_11740,N_11274);
nor UO_257 (O_257,N_10023,N_11760);
and UO_258 (O_258,N_12294,N_11312);
nor UO_259 (O_259,N_11745,N_13439);
and UO_260 (O_260,N_13465,N_12233);
nand UO_261 (O_261,N_10413,N_12516);
nor UO_262 (O_262,N_13814,N_14322);
nor UO_263 (O_263,N_14429,N_11442);
nand UO_264 (O_264,N_10682,N_13690);
and UO_265 (O_265,N_10173,N_12278);
or UO_266 (O_266,N_12497,N_13043);
xor UO_267 (O_267,N_13608,N_10205);
or UO_268 (O_268,N_13251,N_14090);
nor UO_269 (O_269,N_12064,N_13454);
and UO_270 (O_270,N_11891,N_13497);
xor UO_271 (O_271,N_10138,N_10263);
nor UO_272 (O_272,N_10941,N_13854);
xor UO_273 (O_273,N_11231,N_14074);
nor UO_274 (O_274,N_14228,N_10571);
nor UO_275 (O_275,N_11421,N_14575);
nor UO_276 (O_276,N_14455,N_11393);
and UO_277 (O_277,N_10323,N_10620);
or UO_278 (O_278,N_13359,N_11959);
or UO_279 (O_279,N_12089,N_14328);
and UO_280 (O_280,N_14682,N_13260);
nor UO_281 (O_281,N_14610,N_10704);
nand UO_282 (O_282,N_11992,N_14222);
xor UO_283 (O_283,N_14444,N_14017);
or UO_284 (O_284,N_11359,N_14010);
xor UO_285 (O_285,N_12473,N_12328);
nand UO_286 (O_286,N_11621,N_13709);
xnor UO_287 (O_287,N_12614,N_10411);
and UO_288 (O_288,N_14209,N_14297);
or UO_289 (O_289,N_12273,N_10118);
and UO_290 (O_290,N_13924,N_14157);
and UO_291 (O_291,N_13503,N_12429);
or UO_292 (O_292,N_11032,N_14658);
and UO_293 (O_293,N_14919,N_13410);
nand UO_294 (O_294,N_10629,N_13228);
and UO_295 (O_295,N_11886,N_13150);
xor UO_296 (O_296,N_10611,N_13823);
or UO_297 (O_297,N_11790,N_12853);
xnor UO_298 (O_298,N_13469,N_12387);
nor UO_299 (O_299,N_14514,N_14263);
or UO_300 (O_300,N_14565,N_10784);
and UO_301 (O_301,N_10382,N_10561);
or UO_302 (O_302,N_10814,N_13519);
nand UO_303 (O_303,N_12431,N_11271);
and UO_304 (O_304,N_12045,N_14372);
nor UO_305 (O_305,N_13976,N_14812);
or UO_306 (O_306,N_14319,N_10981);
nor UO_307 (O_307,N_10691,N_11105);
xnor UO_308 (O_308,N_14309,N_11489);
or UO_309 (O_309,N_12312,N_12355);
nand UO_310 (O_310,N_13871,N_11404);
nand UO_311 (O_311,N_14303,N_10491);
nand UO_312 (O_312,N_11425,N_10475);
nand UO_313 (O_313,N_12974,N_10817);
or UO_314 (O_314,N_13990,N_14649);
xnor UO_315 (O_315,N_11144,N_14262);
and UO_316 (O_316,N_13942,N_12364);
xor UO_317 (O_317,N_11863,N_14837);
and UO_318 (O_318,N_10918,N_12861);
nand UO_319 (O_319,N_10792,N_13207);
nand UO_320 (O_320,N_14403,N_13605);
and UO_321 (O_321,N_14343,N_14765);
and UO_322 (O_322,N_12656,N_12966);
nor UO_323 (O_323,N_14820,N_11681);
nand UO_324 (O_324,N_10722,N_12270);
nand UO_325 (O_325,N_14281,N_12738);
and UO_326 (O_326,N_13210,N_13914);
and UO_327 (O_327,N_11862,N_12745);
nor UO_328 (O_328,N_12234,N_12395);
or UO_329 (O_329,N_10204,N_13642);
and UO_330 (O_330,N_10568,N_14298);
and UO_331 (O_331,N_11997,N_12988);
or UO_332 (O_332,N_13575,N_11150);
nor UO_333 (O_333,N_13504,N_12858);
and UO_334 (O_334,N_14416,N_12374);
and UO_335 (O_335,N_11273,N_12524);
nor UO_336 (O_336,N_10963,N_12639);
or UO_337 (O_337,N_11497,N_13743);
and UO_338 (O_338,N_12543,N_12941);
nor UO_339 (O_339,N_11797,N_12514);
and UO_340 (O_340,N_14916,N_10236);
nand UO_341 (O_341,N_14605,N_10037);
and UO_342 (O_342,N_12316,N_13264);
nand UO_343 (O_343,N_11462,N_14518);
nor UO_344 (O_344,N_12399,N_13196);
nor UO_345 (O_345,N_12911,N_10367);
or UO_346 (O_346,N_10690,N_11168);
nor UO_347 (O_347,N_12828,N_14311);
or UO_348 (O_348,N_13216,N_13630);
nor UO_349 (O_349,N_11249,N_10907);
nor UO_350 (O_350,N_12033,N_14677);
xor UO_351 (O_351,N_13008,N_12307);
or UO_352 (O_352,N_14233,N_13718);
nor UO_353 (O_353,N_12403,N_11502);
nor UO_354 (O_354,N_13554,N_14254);
and UO_355 (O_355,N_10107,N_11369);
xor UO_356 (O_356,N_13954,N_10348);
and UO_357 (O_357,N_12857,N_13535);
nand UO_358 (O_358,N_12207,N_14493);
and UO_359 (O_359,N_11157,N_10517);
or UO_360 (O_360,N_14744,N_11841);
xnor UO_361 (O_361,N_11976,N_13369);
xnor UO_362 (O_362,N_14079,N_14130);
or UO_363 (O_363,N_13054,N_10742);
or UO_364 (O_364,N_10695,N_13377);
and UO_365 (O_365,N_13606,N_12983);
xor UO_366 (O_366,N_12675,N_13316);
nor UO_367 (O_367,N_12534,N_13645);
nand UO_368 (O_368,N_12323,N_14781);
or UO_369 (O_369,N_13800,N_10920);
and UO_370 (O_370,N_11899,N_12153);
and UO_371 (O_371,N_12536,N_14872);
and UO_372 (O_372,N_10179,N_10841);
nand UO_373 (O_373,N_10859,N_13154);
nor UO_374 (O_374,N_14687,N_14329);
nand UO_375 (O_375,N_14590,N_13745);
or UO_376 (O_376,N_13793,N_12082);
nand UO_377 (O_377,N_12421,N_10539);
or UO_378 (O_378,N_12456,N_13388);
xnor UO_379 (O_379,N_12791,N_12769);
nand UO_380 (O_380,N_11952,N_11784);
or UO_381 (O_381,N_12352,N_10280);
and UO_382 (O_382,N_11403,N_14966);
xor UO_383 (O_383,N_11999,N_12343);
and UO_384 (O_384,N_10075,N_11116);
and UO_385 (O_385,N_10597,N_10724);
nor UO_386 (O_386,N_11849,N_12047);
and UO_387 (O_387,N_14630,N_10005);
or UO_388 (O_388,N_10637,N_13408);
xor UO_389 (O_389,N_10950,N_11903);
xor UO_390 (O_390,N_11264,N_12360);
or UO_391 (O_391,N_14014,N_11751);
xor UO_392 (O_392,N_14824,N_13320);
and UO_393 (O_393,N_12435,N_10669);
or UO_394 (O_394,N_14441,N_12022);
nand UO_395 (O_395,N_10871,N_11729);
and UO_396 (O_396,N_11700,N_10230);
and UO_397 (O_397,N_11880,N_14146);
xnor UO_398 (O_398,N_10605,N_12281);
xor UO_399 (O_399,N_10476,N_14066);
or UO_400 (O_400,N_13271,N_10477);
or UO_401 (O_401,N_11730,N_14277);
nor UO_402 (O_402,N_10777,N_11260);
and UO_403 (O_403,N_13889,N_10282);
or UO_404 (O_404,N_11083,N_10840);
xnor UO_405 (O_405,N_10699,N_12541);
or UO_406 (O_406,N_14180,N_11675);
nor UO_407 (O_407,N_11686,N_12482);
nand UO_408 (O_408,N_14785,N_14451);
xnor UO_409 (O_409,N_12196,N_14940);
xor UO_410 (O_410,N_10592,N_11821);
xor UO_411 (O_411,N_11544,N_10396);
and UO_412 (O_412,N_12887,N_12625);
xor UO_413 (O_413,N_10818,N_12382);
or UO_414 (O_414,N_14220,N_12768);
nor UO_415 (O_415,N_11950,N_11683);
nor UO_416 (O_416,N_13143,N_11516);
or UO_417 (O_417,N_14942,N_11742);
or UO_418 (O_418,N_13122,N_11310);
xnor UO_419 (O_419,N_10026,N_12372);
nor UO_420 (O_420,N_10167,N_12167);
xnor UO_421 (O_421,N_14188,N_10549);
or UO_422 (O_422,N_12304,N_13345);
and UO_423 (O_423,N_12603,N_11270);
xor UO_424 (O_424,N_12578,N_14387);
and UO_425 (O_425,N_12072,N_13748);
xnor UO_426 (O_426,N_14113,N_14546);
and UO_427 (O_427,N_13827,N_10949);
nor UO_428 (O_428,N_10487,N_10572);
xor UO_429 (O_429,N_12144,N_11542);
nand UO_430 (O_430,N_13312,N_13041);
and UO_431 (O_431,N_13020,N_11520);
nor UO_432 (O_432,N_12681,N_13592);
nor UO_433 (O_433,N_12424,N_10289);
nor UO_434 (O_434,N_13958,N_13874);
or UO_435 (O_435,N_12856,N_10671);
nand UO_436 (O_436,N_10004,N_14449);
and UO_437 (O_437,N_12197,N_12703);
and UO_438 (O_438,N_12342,N_10616);
nand UO_439 (O_439,N_11779,N_11923);
nor UO_440 (O_440,N_11973,N_11256);
nor UO_441 (O_441,N_13764,N_13835);
nand UO_442 (O_442,N_12517,N_11482);
or UO_443 (O_443,N_14608,N_11319);
xor UO_444 (O_444,N_12796,N_14206);
xnor UO_445 (O_445,N_10825,N_14098);
or UO_446 (O_446,N_14247,N_13080);
and UO_447 (O_447,N_10275,N_14234);
or UO_448 (O_448,N_14342,N_10755);
or UO_449 (O_449,N_10683,N_14778);
nand UO_450 (O_450,N_10121,N_14706);
and UO_451 (O_451,N_14242,N_10593);
and UO_452 (O_452,N_13531,N_14110);
xor UO_453 (O_453,N_12260,N_13179);
or UO_454 (O_454,N_10861,N_10375);
xor UO_455 (O_455,N_13884,N_10350);
xor UO_456 (O_456,N_14891,N_10457);
nand UO_457 (O_457,N_12783,N_13148);
nand UO_458 (O_458,N_11477,N_13181);
nand UO_459 (O_459,N_14853,N_10634);
and UO_460 (O_460,N_11223,N_11071);
and UO_461 (O_461,N_13155,N_10780);
xnor UO_462 (O_462,N_13037,N_11470);
nor UO_463 (O_463,N_12093,N_13002);
xor UO_464 (O_464,N_14544,N_11750);
nor UO_465 (O_465,N_10514,N_12805);
and UO_466 (O_466,N_10157,N_13474);
and UO_467 (O_467,N_14126,N_14592);
and UO_468 (O_468,N_10503,N_11020);
and UO_469 (O_469,N_10133,N_12347);
nor UO_470 (O_470,N_12894,N_10478);
and UO_471 (O_471,N_11194,N_10247);
and UO_472 (O_472,N_12487,N_14527);
nor UO_473 (O_473,N_13394,N_13334);
and UO_474 (O_474,N_10753,N_10974);
xor UO_475 (O_475,N_10175,N_10553);
xnor UO_476 (O_476,N_10513,N_10534);
nor UO_477 (O_477,N_13769,N_13788);
xnor UO_478 (O_478,N_14152,N_10607);
and UO_479 (O_479,N_12699,N_10606);
or UO_480 (O_480,N_13133,N_12166);
nor UO_481 (O_481,N_10218,N_14106);
nand UO_482 (O_482,N_13833,N_10988);
xor UO_483 (O_483,N_14498,N_10243);
xor UO_484 (O_484,N_13475,N_13627);
nor UO_485 (O_485,N_12407,N_10644);
nor UO_486 (O_486,N_12291,N_11748);
and UO_487 (O_487,N_13342,N_14085);
or UO_488 (O_488,N_13892,N_11126);
and UO_489 (O_489,N_13121,N_10882);
or UO_490 (O_490,N_13031,N_10701);
or UO_491 (O_491,N_10507,N_11772);
xnor UO_492 (O_492,N_10957,N_12727);
or UO_493 (O_493,N_14475,N_14772);
and UO_494 (O_494,N_14775,N_13951);
xor UO_495 (O_495,N_14390,N_10139);
or UO_496 (O_496,N_12430,N_11778);
nand UO_497 (O_497,N_12396,N_10816);
nor UO_498 (O_498,N_12035,N_14478);
nor UO_499 (O_499,N_11413,N_13840);
nor UO_500 (O_500,N_13665,N_12474);
nand UO_501 (O_501,N_14740,N_11881);
and UO_502 (O_502,N_10581,N_14140);
and UO_503 (O_503,N_13661,N_10410);
or UO_504 (O_504,N_13971,N_14748);
or UO_505 (O_505,N_10065,N_12604);
nand UO_506 (O_506,N_12890,N_11431);
nand UO_507 (O_507,N_12303,N_13202);
or UO_508 (O_508,N_11443,N_12365);
and UO_509 (O_509,N_14588,N_14895);
xnor UO_510 (O_510,N_12686,N_13629);
nand UO_511 (O_511,N_11352,N_13033);
nand UO_512 (O_512,N_12219,N_12178);
nand UO_513 (O_513,N_10405,N_14894);
nor UO_514 (O_514,N_11066,N_10112);
and UO_515 (O_515,N_12422,N_13552);
nand UO_516 (O_516,N_11924,N_10706);
and UO_517 (O_517,N_13775,N_13789);
or UO_518 (O_518,N_12615,N_14346);
xnor UO_519 (O_519,N_14040,N_12274);
nor UO_520 (O_520,N_13463,N_11672);
and UO_521 (O_521,N_12024,N_13632);
and UO_522 (O_522,N_13396,N_10783);
or UO_523 (O_523,N_13171,N_10901);
and UO_524 (O_524,N_11218,N_10312);
or UO_525 (O_525,N_14446,N_13596);
nand UO_526 (O_526,N_10060,N_10249);
nor UO_527 (O_527,N_11515,N_14259);
nand UO_528 (O_528,N_14642,N_14570);
xor UO_529 (O_529,N_13941,N_14634);
nand UO_530 (O_530,N_12557,N_10505);
nor UO_531 (O_531,N_14063,N_11677);
and UO_532 (O_532,N_14019,N_13073);
nor UO_533 (O_533,N_10071,N_12710);
nand UO_534 (O_534,N_10195,N_11637);
and UO_535 (O_535,N_11708,N_10104);
and UO_536 (O_536,N_11965,N_11430);
and UO_537 (O_537,N_12922,N_10688);
nand UO_538 (O_538,N_13872,N_13411);
xor UO_539 (O_539,N_12097,N_11054);
or UO_540 (O_540,N_10309,N_12251);
and UO_541 (O_541,N_13897,N_10315);
nand UO_542 (O_542,N_11329,N_10142);
and UO_543 (O_543,N_10053,N_12866);
and UO_544 (O_544,N_12181,N_14029);
or UO_545 (O_545,N_11471,N_11481);
xor UO_546 (O_546,N_14338,N_10741);
nor UO_547 (O_547,N_14901,N_14174);
nor UO_548 (O_548,N_13553,N_10177);
nand UO_549 (O_549,N_14023,N_10331);
nand UO_550 (O_550,N_14659,N_13356);
xnor UO_551 (O_551,N_12441,N_11318);
and UO_552 (O_552,N_13422,N_11484);
xnor UO_553 (O_553,N_13034,N_11454);
nand UO_554 (O_554,N_13447,N_10283);
xnor UO_555 (O_555,N_13604,N_11799);
nand UO_556 (O_556,N_14179,N_12976);
nor UO_557 (O_557,N_13577,N_12709);
or UO_558 (O_558,N_14926,N_10588);
or UO_559 (O_559,N_13367,N_13018);
nand UO_560 (O_560,N_14552,N_10836);
nand UO_561 (O_561,N_13142,N_11769);
nor UO_562 (O_562,N_10779,N_13610);
and UO_563 (O_563,N_14628,N_10746);
nor UO_564 (O_564,N_12933,N_13302);
nand UO_565 (O_565,N_10707,N_13644);
or UO_566 (O_566,N_14686,N_14224);
and UO_567 (O_567,N_11137,N_14026);
or UO_568 (O_568,N_14219,N_10427);
and UO_569 (O_569,N_13214,N_10909);
or UO_570 (O_570,N_14733,N_13450);
nor UO_571 (O_571,N_14918,N_12004);
or UO_572 (O_572,N_14273,N_11142);
nand UO_573 (O_573,N_13226,N_12596);
or UO_574 (O_574,N_13900,N_11014);
nor UO_575 (O_575,N_13208,N_11082);
or UO_576 (O_576,N_11018,N_14567);
xor UO_577 (O_577,N_10267,N_10694);
xor UO_578 (O_578,N_12715,N_10989);
nand UO_579 (O_579,N_14821,N_14650);
xor UO_580 (O_580,N_13085,N_13634);
xnor UO_581 (O_581,N_14643,N_11203);
nor UO_582 (O_582,N_10943,N_10985);
xnor UO_583 (O_583,N_10813,N_12561);
nor UO_584 (O_584,N_13392,N_11820);
or UO_585 (O_585,N_13158,N_10162);
and UO_586 (O_586,N_12998,N_12679);
and UO_587 (O_587,N_14500,N_11164);
xor UO_588 (O_588,N_10721,N_14313);
nor UO_589 (O_589,N_12935,N_10070);
or UO_590 (O_590,N_10991,N_12203);
and UO_591 (O_591,N_11659,N_10939);
nand UO_592 (O_592,N_11100,N_13886);
xnor UO_593 (O_593,N_12488,N_11277);
xor UO_594 (O_594,N_10045,N_12249);
xor UO_595 (O_595,N_12528,N_14915);
or UO_596 (O_596,N_12350,N_14139);
and UO_597 (O_597,N_13479,N_13873);
or UO_598 (O_598,N_10573,N_14045);
or UO_599 (O_599,N_11981,N_14694);
and UO_600 (O_600,N_13339,N_14367);
nand UO_601 (O_601,N_10300,N_14529);
or UO_602 (O_602,N_13485,N_12123);
and UO_603 (O_603,N_13834,N_13267);
nand UO_604 (O_604,N_11361,N_12716);
or UO_605 (O_605,N_11946,N_13038);
or UO_606 (O_606,N_12907,N_12122);
nand UO_607 (O_607,N_10219,N_11202);
or UO_608 (O_608,N_11958,N_12440);
nor UO_609 (O_609,N_12010,N_10202);
and UO_610 (O_610,N_13257,N_12718);
nor UO_611 (O_611,N_13213,N_13837);
nand UO_612 (O_612,N_13492,N_14048);
xor UO_613 (O_613,N_10945,N_13585);
or UO_614 (O_614,N_13866,N_11092);
and UO_615 (O_615,N_13956,N_12116);
nand UO_616 (O_616,N_13100,N_11636);
nand UO_617 (O_617,N_14892,N_12332);
nor UO_618 (O_618,N_11756,N_14864);
nor UO_619 (O_619,N_11139,N_14964);
nor UO_620 (O_620,N_14714,N_14899);
nand UO_621 (O_621,N_13801,N_11723);
nand UO_622 (O_622,N_14472,N_11588);
and UO_623 (O_623,N_10667,N_13624);
xor UO_624 (O_624,N_14599,N_11143);
and UO_625 (O_625,N_10030,N_12672);
nand UO_626 (O_626,N_11645,N_11665);
xor UO_627 (O_627,N_11458,N_13329);
nand UO_628 (O_628,N_11333,N_10054);
or UO_629 (O_629,N_11619,N_10829);
and UO_630 (O_630,N_10502,N_13344);
nor UO_631 (O_631,N_12501,N_10186);
xnor UO_632 (O_632,N_14576,N_11394);
and UO_633 (O_633,N_10966,N_11013);
nand UO_634 (O_634,N_13464,N_12817);
nor UO_635 (O_635,N_11127,N_13182);
or UO_636 (O_636,N_10891,N_13518);
xor UO_637 (O_637,N_11062,N_14199);
xnor UO_638 (O_638,N_10525,N_12978);
or UO_639 (O_639,N_12879,N_13538);
or UO_640 (O_640,N_12720,N_10431);
xnor UO_641 (O_641,N_10094,N_11009);
nand UO_642 (O_642,N_13349,N_12453);
xnor UO_643 (O_643,N_12009,N_13520);
and UO_644 (O_644,N_12100,N_10643);
and UO_645 (O_645,N_10995,N_14312);
or UO_646 (O_646,N_14361,N_10822);
nand UO_647 (O_647,N_11860,N_14347);
nor UO_648 (O_648,N_10330,N_13168);
nor UO_649 (O_649,N_14318,N_10344);
nor UO_650 (O_650,N_11048,N_14468);
xor UO_651 (O_651,N_11575,N_13581);
nand UO_652 (O_652,N_14923,N_12243);
xnor UO_653 (O_653,N_11283,N_10815);
nor UO_654 (O_654,N_10846,N_13235);
nor UO_655 (O_655,N_12628,N_14993);
or UO_656 (O_656,N_10271,N_13910);
nor UO_657 (O_657,N_13082,N_10870);
nand UO_658 (O_658,N_11755,N_10709);
or UO_659 (O_659,N_13670,N_14584);
and UO_660 (O_660,N_11480,N_12891);
nand UO_661 (O_661,N_11389,N_12521);
and UO_662 (O_662,N_14398,N_11085);
xnor UO_663 (O_663,N_11055,N_11696);
xnor UO_664 (O_664,N_12134,N_13543);
nor UO_665 (O_665,N_11622,N_13242);
or UO_666 (O_666,N_14290,N_11577);
and UO_667 (O_667,N_13759,N_12671);
nand UO_668 (O_668,N_14903,N_14060);
nor UO_669 (O_669,N_10600,N_10201);
nor UO_670 (O_670,N_12605,N_13185);
and UO_671 (O_671,N_13136,N_12201);
and UO_672 (O_672,N_14358,N_14809);
nor UO_673 (O_673,N_12337,N_12764);
xor UO_674 (O_674,N_12119,N_13138);
nor UO_675 (O_675,N_10370,N_13894);
nor UO_676 (O_676,N_14235,N_13589);
or UO_677 (O_677,N_12755,N_12067);
nor UO_678 (O_678,N_12102,N_11420);
nor UO_679 (O_679,N_12647,N_11107);
xor UO_680 (O_680,N_10584,N_14438);
nand UO_681 (O_681,N_13086,N_12925);
or UO_682 (O_682,N_13101,N_14325);
nand UO_683 (O_683,N_13131,N_10072);
and UO_684 (O_684,N_12965,N_12087);
nand UO_685 (O_685,N_10635,N_10843);
or UO_686 (O_686,N_11802,N_12707);
nand UO_687 (O_687,N_14717,N_14456);
nand UO_688 (O_688,N_13308,N_11589);
nor UO_689 (O_689,N_13974,N_12949);
and UO_690 (O_690,N_10763,N_11111);
and UO_691 (O_691,N_12873,N_11949);
or UO_692 (O_692,N_14308,N_14266);
nor UO_693 (O_693,N_13384,N_13651);
nor UO_694 (O_694,N_11845,N_11887);
and UO_695 (O_695,N_13985,N_11490);
nand UO_696 (O_696,N_13917,N_11807);
xnor UO_697 (O_697,N_11669,N_13846);
xor UO_698 (O_698,N_14125,N_12105);
and UO_699 (O_699,N_11796,N_11438);
nand UO_700 (O_700,N_10666,N_13250);
nand UO_701 (O_701,N_11512,N_14760);
xor UO_702 (O_702,N_11518,N_11330);
nor UO_703 (O_703,N_12685,N_10772);
nand UO_704 (O_704,N_11521,N_11305);
or UO_705 (O_705,N_10383,N_14621);
xor UO_706 (O_706,N_12282,N_10899);
and UO_707 (O_707,N_12868,N_11534);
nand UO_708 (O_708,N_13933,N_11455);
or UO_709 (O_709,N_14203,N_12098);
or UO_710 (O_710,N_10506,N_11380);
or UO_711 (O_711,N_11557,N_14283);
xnor UO_712 (O_712,N_12288,N_13768);
nand UO_713 (O_713,N_10318,N_12479);
and UO_714 (O_714,N_13252,N_10998);
nand UO_715 (O_715,N_12404,N_12130);
nor UO_716 (O_716,N_13314,N_12275);
and UO_717 (O_717,N_10726,N_12247);
nor UO_718 (O_718,N_13169,N_14432);
nand UO_719 (O_719,N_13472,N_11643);
nor UO_720 (O_720,N_10464,N_10481);
nor UO_721 (O_721,N_10278,N_10728);
nor UO_722 (O_722,N_14245,N_13851);
nand UO_723 (O_723,N_11101,N_11251);
xnor UO_724 (O_724,N_12975,N_11916);
nand UO_725 (O_725,N_14159,N_12080);
nor UO_726 (O_726,N_12269,N_11115);
and UO_727 (O_727,N_11098,N_14751);
or UO_728 (O_728,N_11813,N_11320);
xnor UO_729 (O_729,N_11652,N_14851);
nor UO_730 (O_730,N_12095,N_10619);
and UO_731 (O_731,N_13856,N_11081);
nand UO_732 (O_732,N_13425,N_10551);
and UO_733 (O_733,N_13300,N_11220);
nor UO_734 (O_734,N_14525,N_13152);
xnor UO_735 (O_735,N_14351,N_12272);
and UO_736 (O_736,N_13618,N_10873);
xnor UO_737 (O_737,N_14345,N_12666);
nor UO_738 (O_738,N_11889,N_10076);
nand UO_739 (O_739,N_14376,N_11342);
xnor UO_740 (O_740,N_12040,N_10785);
nor UO_741 (O_741,N_10100,N_10266);
xor UO_742 (O_742,N_11532,N_14953);
nor UO_743 (O_743,N_11870,N_10174);
xor UO_744 (O_744,N_12651,N_10912);
xor UO_745 (O_745,N_14381,N_11566);
xor UO_746 (O_746,N_11559,N_13151);
or UO_747 (O_747,N_10276,N_10868);
or UO_748 (O_748,N_14183,N_14024);
and UO_749 (O_749,N_12155,N_13303);
nand UO_750 (O_750,N_14050,N_10105);
and UO_751 (O_751,N_12051,N_13412);
nor UO_752 (O_752,N_11222,N_13327);
or UO_753 (O_753,N_14938,N_13486);
nor UO_754 (O_754,N_13968,N_12226);
and UO_755 (O_755,N_11181,N_14391);
nor UO_756 (O_756,N_13973,N_13123);
xor UO_757 (O_757,N_10659,N_13230);
nor UO_758 (O_758,N_10131,N_13195);
xnor UO_759 (O_759,N_14955,N_12570);
nand UO_760 (O_760,N_11572,N_14843);
xor UO_761 (O_761,N_13693,N_13560);
xnor UO_762 (O_762,N_13586,N_11871);
xnor UO_763 (O_763,N_13407,N_13090);
xor UO_764 (O_764,N_11355,N_14301);
xnor UO_765 (O_765,N_12286,N_13346);
nor UO_766 (O_766,N_13778,N_13313);
or UO_767 (O_767,N_10486,N_12785);
and UO_768 (O_768,N_13858,N_14069);
nand UO_769 (O_769,N_13972,N_11483);
nand UO_770 (O_770,N_13194,N_12509);
and UO_771 (O_771,N_11313,N_12790);
nand UO_772 (O_772,N_11087,N_11758);
nor UO_773 (O_773,N_14170,N_11079);
nor UO_774 (O_774,N_13671,N_11495);
nand UO_775 (O_775,N_10544,N_12864);
or UO_776 (O_776,N_11538,N_12137);
nand UO_777 (O_777,N_10787,N_14101);
or UO_778 (O_778,N_12218,N_14011);
xor UO_779 (O_779,N_10765,N_14786);
or UO_780 (O_780,N_12725,N_13614);
and UO_781 (O_781,N_11956,N_11243);
and UO_782 (O_782,N_11227,N_11350);
and UO_783 (O_783,N_10456,N_13423);
nand UO_784 (O_784,N_13337,N_12563);
nand UO_785 (O_785,N_11197,N_14025);
nor UO_786 (O_786,N_11510,N_10009);
nand UO_787 (O_787,N_14976,N_11704);
nor UO_788 (O_788,N_13817,N_13005);
or UO_789 (O_789,N_13786,N_13739);
or UO_790 (O_790,N_14925,N_11617);
nor UO_791 (O_791,N_12133,N_12648);
nor UO_792 (O_792,N_13611,N_10499);
nand UO_793 (O_793,N_13003,N_13419);
nand UO_794 (O_794,N_14623,N_12254);
nand UO_795 (O_795,N_10420,N_12549);
and UO_796 (O_796,N_10872,N_13522);
xnor UO_797 (O_797,N_11217,N_10223);
and UO_798 (O_798,N_13084,N_13461);
nor UO_799 (O_799,N_10598,N_13848);
nand UO_800 (O_800,N_10535,N_12036);
nor UO_801 (O_801,N_13831,N_13293);
or UO_802 (O_802,N_10904,N_12248);
xnor UO_803 (O_803,N_12462,N_11103);
nor UO_804 (O_804,N_12330,N_12740);
nand UO_805 (O_805,N_10508,N_10093);
nor UO_806 (O_806,N_14240,N_10930);
xnor UO_807 (O_807,N_12152,N_11247);
or UO_808 (O_808,N_12193,N_12114);
xor UO_809 (O_809,N_14243,N_14279);
or UO_810 (O_810,N_14959,N_14943);
nor UO_811 (O_811,N_14044,N_11030);
nor UO_812 (O_812,N_12849,N_11096);
or UO_813 (O_813,N_13514,N_13269);
nand UO_814 (O_814,N_11920,N_14855);
nor UO_815 (O_815,N_12232,N_11983);
nand UO_816 (O_816,N_10011,N_14216);
or UO_817 (O_817,N_11731,N_11982);
nand UO_818 (O_818,N_14483,N_14182);
nor UO_819 (O_819,N_13266,N_10567);
xnor UO_820 (O_820,N_13113,N_11590);
nand UO_821 (O_821,N_10527,N_10122);
xnor UO_822 (O_822,N_12229,N_10700);
nand UO_823 (O_823,N_13562,N_14109);
nor UO_824 (O_824,N_11529,N_10569);
nor UO_825 (O_825,N_10015,N_10849);
nand UO_826 (O_826,N_10115,N_13146);
and UO_827 (O_827,N_14032,N_10089);
xnor UO_828 (O_828,N_12060,N_13061);
nor UO_829 (O_829,N_13912,N_13716);
xor UO_830 (O_830,N_13909,N_11037);
xor UO_831 (O_831,N_13183,N_13876);
and UO_832 (O_832,N_11084,N_11466);
xor UO_833 (O_833,N_10845,N_10387);
nor UO_834 (O_834,N_14445,N_14952);
nand UO_835 (O_835,N_11783,N_10911);
or UO_836 (O_836,N_12476,N_12470);
or UO_837 (O_837,N_11592,N_12731);
nor UO_838 (O_838,N_13021,N_11167);
or UO_839 (O_839,N_12698,N_14920);
and UO_840 (O_840,N_13777,N_11491);
and UO_841 (O_841,N_11793,N_14718);
xnor UO_842 (O_842,N_10391,N_13011);
or UO_843 (O_843,N_13998,N_10485);
nor UO_844 (O_844,N_12094,N_10185);
or UO_845 (O_845,N_12402,N_10733);
xor UO_846 (O_846,N_10160,N_11049);
nor UO_847 (O_847,N_14198,N_11984);
or UO_848 (O_848,N_11511,N_12617);
and UO_849 (O_849,N_10229,N_12913);
and UO_850 (O_850,N_12613,N_12902);
and UO_851 (O_851,N_11951,N_12691);
nor UO_852 (O_852,N_12714,N_14316);
and UO_853 (O_853,N_12132,N_10268);
nor UO_854 (O_854,N_13818,N_10622);
nand UO_855 (O_855,N_13374,N_13728);
or UO_856 (O_856,N_12743,N_10184);
or UO_857 (O_857,N_14208,N_10446);
nor UO_858 (O_858,N_10664,N_12566);
nor UO_859 (O_859,N_12434,N_13448);
or UO_860 (O_860,N_11088,N_10428);
or UO_861 (O_861,N_11331,N_14094);
xor UO_862 (O_862,N_14433,N_11025);
or UO_863 (O_863,N_11609,N_12055);
nor UO_864 (O_864,N_14331,N_10442);
or UO_865 (O_865,N_12164,N_13368);
nand UO_866 (O_866,N_12505,N_10926);
xnor UO_867 (O_867,N_13687,N_10893);
and UO_868 (O_868,N_13888,N_14734);
xor UO_869 (O_869,N_13229,N_12770);
xor UO_870 (O_870,N_12580,N_13016);
xnor UO_871 (O_871,N_12622,N_13307);
or UO_872 (O_872,N_14384,N_11827);
nor UO_873 (O_873,N_11282,N_13105);
nor UO_874 (O_874,N_14984,N_11368);
xnor UO_875 (O_875,N_11288,N_13244);
and UO_876 (O_876,N_14910,N_14670);
nor UO_877 (O_877,N_13491,N_10214);
xor UO_878 (O_878,N_13784,N_12176);
nand UO_879 (O_879,N_10806,N_10878);
nand UO_880 (O_880,N_13779,N_11607);
nand UO_881 (O_881,N_10766,N_13657);
or UO_882 (O_882,N_11302,N_13205);
and UO_883 (O_883,N_10091,N_14870);
or UO_884 (O_884,N_10639,N_13108);
and UO_885 (O_885,N_14692,N_10084);
nand UO_886 (O_886,N_11753,N_11926);
or UO_887 (O_887,N_13572,N_13206);
or UO_888 (O_888,N_14399,N_10799);
or UO_889 (O_889,N_14738,N_12143);
nor UO_890 (O_890,N_11000,N_10279);
and UO_891 (O_891,N_14419,N_13376);
or UO_892 (O_892,N_12257,N_12870);
and UO_893 (O_893,N_12508,N_12208);
or UO_894 (O_894,N_13175,N_13351);
and UO_895 (O_895,N_11345,N_14163);
and UO_896 (O_896,N_11627,N_11465);
and UO_897 (O_897,N_10510,N_12573);
and UO_898 (O_898,N_14200,N_14257);
xnor UO_899 (O_899,N_10522,N_10751);
or UO_900 (O_900,N_13816,N_14720);
xnor UO_901 (O_901,N_14232,N_10355);
nand UO_902 (O_902,N_12439,N_11427);
or UO_903 (O_903,N_13401,N_11190);
nand UO_904 (O_904,N_11237,N_12826);
nand UO_905 (O_905,N_13355,N_13477);
nand UO_906 (O_906,N_11670,N_10062);
nor UO_907 (O_907,N_10956,N_11705);
xor UO_908 (O_908,N_13044,N_14671);
or UO_909 (O_909,N_14826,N_10767);
or UO_910 (O_910,N_11749,N_13826);
xor UO_911 (O_911,N_14547,N_12398);
and UO_912 (O_912,N_10018,N_12135);
xor UO_913 (O_913,N_11417,N_11549);
nand UO_914 (O_914,N_12255,N_13290);
xor UO_915 (O_915,N_10452,N_13580);
or UO_916 (O_916,N_11153,N_11562);
nand UO_917 (O_917,N_10745,N_10347);
xor UO_918 (O_918,N_12786,N_14845);
or UO_919 (O_919,N_12795,N_11189);
nor UO_920 (O_920,N_11582,N_13700);
or UO_921 (O_921,N_11701,N_10187);
and UO_922 (O_922,N_11347,N_12587);
nor UO_923 (O_923,N_11601,N_14581);
nand UO_924 (O_924,N_10027,N_12901);
xnor UO_925 (O_925,N_13695,N_14519);
nand UO_926 (O_926,N_10602,N_13681);
xnor UO_927 (O_927,N_14105,N_14031);
xor UO_928 (O_928,N_12746,N_14912);
nand UO_929 (O_929,N_10090,N_14051);
nand UO_930 (O_930,N_12469,N_13749);
xnor UO_931 (O_931,N_13680,N_11204);
nor UO_932 (O_932,N_14187,N_13631);
nand UO_933 (O_933,N_10710,N_11097);
nor UO_934 (O_934,N_10242,N_11468);
and UO_935 (O_935,N_10474,N_11335);
or UO_936 (O_936,N_13402,N_12331);
nor UO_937 (O_937,N_12781,N_14601);
nor UO_938 (O_938,N_10137,N_10906);
and UO_939 (O_939,N_10773,N_10316);
xnor UO_940 (O_940,N_10057,N_10594);
nand UO_941 (O_941,N_13511,N_11396);
or UO_942 (O_942,N_13864,N_12542);
or UO_943 (O_943,N_14035,N_12448);
or UO_944 (O_944,N_12150,N_12486);
nand UO_945 (O_945,N_11323,N_11531);
xnor UO_946 (O_946,N_14804,N_14457);
and UO_947 (O_947,N_12348,N_10358);
and UO_948 (O_948,N_14863,N_12378);
nor UO_949 (O_949,N_12690,N_11371);
nor UO_950 (O_950,N_11901,N_11174);
and UO_951 (O_951,N_14510,N_12104);
or UO_952 (O_952,N_11060,N_11576);
or UO_953 (O_953,N_14251,N_12079);
xor UO_954 (O_954,N_12766,N_11479);
or UO_955 (O_955,N_11966,N_14873);
xor UO_956 (O_956,N_11835,N_10430);
nand UO_957 (O_957,N_13761,N_10808);
xor UO_958 (O_958,N_10547,N_12723);
xor UO_959 (O_959,N_12964,N_10770);
or UO_960 (O_960,N_10371,N_11063);
xor UO_961 (O_961,N_11699,N_11022);
xor UO_962 (O_962,N_10832,N_13563);
xnor UO_963 (O_963,N_12463,N_14005);
nor UO_964 (O_964,N_14722,N_11702);
nor UO_965 (O_965,N_12994,N_13406);
nor UO_966 (O_966,N_10958,N_13982);
xor UO_967 (O_967,N_13946,N_11858);
nor UO_968 (O_968,N_12619,N_13467);
nor UO_969 (O_969,N_11583,N_11564);
or UO_970 (O_970,N_10216,N_13110);
or UO_971 (O_971,N_11324,N_14341);
xor UO_972 (O_972,N_11524,N_13616);
or UO_973 (O_973,N_14753,N_13258);
and UO_974 (O_974,N_12995,N_12800);
nand UO_975 (O_975,N_14972,N_11224);
xnor UO_976 (O_976,N_13571,N_11678);
or UO_977 (O_977,N_13935,N_13091);
or UO_978 (O_978,N_10696,N_12523);
or UO_979 (O_979,N_14593,N_10419);
xor UO_980 (O_980,N_11724,N_12477);
and UO_981 (O_981,N_12050,N_13284);
nor UO_982 (O_982,N_13698,N_14417);
nor UO_983 (O_983,N_12041,N_14792);
nand UO_984 (O_984,N_11551,N_14323);
nand UO_985 (O_985,N_10954,N_10343);
nand UO_986 (O_986,N_11044,N_13696);
or UO_987 (O_987,N_14631,N_10240);
nand UO_988 (O_988,N_14053,N_12244);
nor UO_989 (O_989,N_14627,N_13787);
nor UO_990 (O_990,N_13717,N_10288);
or UO_991 (O_991,N_10786,N_11293);
or UO_992 (O_992,N_12452,N_12688);
and UO_993 (O_993,N_11239,N_12920);
nand UO_994 (O_994,N_10123,N_13444);
and UO_995 (O_995,N_13087,N_10467);
or UO_996 (O_996,N_12190,N_10390);
nor UO_997 (O_997,N_13825,N_11123);
nor UO_998 (O_998,N_13566,N_13426);
xor UO_999 (O_999,N_10438,N_12206);
or UO_1000 (O_1000,N_12245,N_12585);
nor UO_1001 (O_1001,N_10168,N_12838);
or UO_1002 (O_1002,N_13780,N_13482);
nand UO_1003 (O_1003,N_10008,N_13615);
or UO_1004 (O_1004,N_10092,N_11822);
xnor UO_1005 (O_1005,N_14389,N_10754);
nand UO_1006 (O_1006,N_14858,N_11606);
and UO_1007 (O_1007,N_11125,N_12427);
nand UO_1008 (O_1008,N_13579,N_12775);
or UO_1009 (O_1009,N_10051,N_14315);
nor UO_1010 (O_1010,N_11219,N_10468);
or UO_1011 (O_1011,N_11121,N_10365);
nor UO_1012 (O_1012,N_12046,N_11232);
nor UO_1013 (O_1013,N_10922,N_14076);
and UO_1014 (O_1014,N_12049,N_10725);
nand UO_1015 (O_1015,N_10925,N_11541);
xor UO_1016 (O_1016,N_13438,N_10715);
nor UO_1017 (O_1017,N_14614,N_10255);
nor UO_1018 (O_1018,N_14127,N_13362);
nand UO_1019 (O_1019,N_12765,N_10254);
nand UO_1020 (O_1020,N_13187,N_10862);
or UO_1021 (O_1021,N_12236,N_14723);
nor UO_1022 (O_1022,N_12263,N_13295);
or UO_1023 (O_1023,N_13844,N_11401);
xor UO_1024 (O_1024,N_12369,N_12444);
xnor UO_1025 (O_1025,N_12915,N_10226);
nand UO_1026 (O_1026,N_14615,N_10626);
nor UO_1027 (O_1027,N_11135,N_13219);
nor UO_1028 (O_1028,N_13516,N_13542);
nand UO_1029 (O_1029,N_10141,N_14071);
or UO_1030 (O_1030,N_12327,N_10495);
xnor UO_1031 (O_1031,N_11272,N_13940);
nand UO_1032 (O_1032,N_11688,N_11854);
nand UO_1033 (O_1033,N_11410,N_10449);
xnor UO_1034 (O_1034,N_11789,N_12059);
xor UO_1035 (O_1035,N_13536,N_13762);
and UO_1036 (O_1036,N_11711,N_13275);
nor UO_1037 (O_1037,N_11390,N_14715);
xor UO_1038 (O_1038,N_14052,N_10373);
nand UO_1039 (O_1039,N_14336,N_12859);
nor UO_1040 (O_1040,N_12609,N_10781);
and UO_1041 (O_1041,N_10615,N_10515);
and UO_1042 (O_1042,N_10199,N_13891);
xnor UO_1043 (O_1043,N_13925,N_13042);
xnor UO_1044 (O_1044,N_11091,N_10326);
or UO_1045 (O_1045,N_11384,N_14168);
nand UO_1046 (O_1046,N_10579,N_11336);
xor UO_1047 (O_1047,N_11625,N_13822);
nand UO_1048 (O_1048,N_11805,N_10320);
nor UO_1049 (O_1049,N_12002,N_14181);
nor UO_1050 (O_1050,N_12267,N_13964);
xnor UO_1051 (O_1051,N_14495,N_12054);
nor UO_1052 (O_1052,N_14030,N_14278);
and UO_1053 (O_1053,N_12455,N_10250);
nand UO_1054 (O_1054,N_12464,N_13079);
nand UO_1055 (O_1055,N_13254,N_13298);
and UO_1056 (O_1056,N_12222,N_10148);
and UO_1057 (O_1057,N_10979,N_14696);
or UO_1058 (O_1058,N_12214,N_12960);
nand UO_1059 (O_1059,N_14006,N_10577);
nand UO_1060 (O_1060,N_13673,N_14931);
and UO_1061 (O_1061,N_13526,N_14509);
and UO_1062 (O_1062,N_11381,N_11833);
and UO_1063 (O_1063,N_10860,N_14730);
xnor UO_1064 (O_1064,N_13662,N_12886);
and UO_1065 (O_1065,N_11781,N_13363);
xor UO_1066 (O_1066,N_11727,N_10007);
and UO_1067 (O_1067,N_13115,N_11130);
nand UO_1068 (O_1068,N_14293,N_12379);
nor UO_1069 (O_1069,N_12831,N_11785);
nor UO_1070 (O_1070,N_12025,N_12954);
xor UO_1071 (O_1071,N_12187,N_12113);
or UO_1072 (O_1072,N_12170,N_10461);
xnor UO_1073 (O_1073,N_10417,N_12168);
or UO_1074 (O_1074,N_14077,N_14189);
nor UO_1075 (O_1075,N_11503,N_13813);
nand UO_1076 (O_1076,N_13273,N_13097);
xnor UO_1077 (O_1077,N_10604,N_11469);
nor UO_1078 (O_1078,N_11201,N_13238);
or UO_1079 (O_1079,N_14861,N_10647);
xnor UO_1080 (O_1080,N_14764,N_14392);
nand UO_1081 (O_1081,N_13068,N_12754);
nand UO_1082 (O_1082,N_10292,N_10921);
and UO_1083 (O_1083,N_10952,N_12552);
and UO_1084 (O_1084,N_13126,N_10362);
nor UO_1085 (O_1085,N_12674,N_13708);
or UO_1086 (O_1086,N_13487,N_14049);
xor UO_1087 (O_1087,N_13802,N_12450);
and UO_1088 (O_1088,N_10550,N_14896);
or UO_1089 (O_1089,N_11667,N_14683);
and UO_1090 (O_1090,N_10538,N_13928);
nor UO_1091 (O_1091,N_12673,N_12363);
and UO_1092 (O_1092,N_13927,N_14900);
and UO_1093 (O_1093,N_13989,N_13723);
nor UO_1094 (O_1094,N_11990,N_11447);
and UO_1095 (O_1095,N_10771,N_10636);
nor UO_1096 (O_1096,N_14839,N_10983);
or UO_1097 (O_1097,N_12653,N_10480);
xnor UO_1098 (O_1098,N_14086,N_10589);
xor UO_1099 (O_1099,N_10645,N_14138);
or UO_1100 (O_1100,N_10284,N_12818);
xor UO_1101 (O_1101,N_11513,N_11774);
nor UO_1102 (O_1102,N_14678,N_11626);
nor UO_1103 (O_1103,N_10389,N_10540);
nor UO_1104 (O_1104,N_14332,N_10106);
nor UO_1105 (O_1105,N_14261,N_11045);
or UO_1106 (O_1106,N_13527,N_10811);
or UO_1107 (O_1107,N_10374,N_10776);
and UO_1108 (O_1108,N_14928,N_10451);
xor UO_1109 (O_1109,N_13507,N_13231);
nand UO_1110 (O_1110,N_12595,N_11473);
nand UO_1111 (O_1111,N_12495,N_11019);
and UO_1112 (O_1112,N_13049,N_10401);
nand UO_1113 (O_1113,N_12091,N_12512);
nor UO_1114 (O_1114,N_13460,N_10730);
or UO_1115 (O_1115,N_14202,N_11975);
nand UO_1116 (O_1116,N_10482,N_10670);
xor UO_1117 (O_1117,N_13380,N_13017);
or UO_1118 (O_1118,N_12896,N_11650);
nand UO_1119 (O_1119,N_10251,N_11640);
nand UO_1120 (O_1120,N_10501,N_11744);
and UO_1121 (O_1121,N_11496,N_13607);
nor UO_1122 (O_1122,N_14988,N_14841);
nand UO_1123 (O_1123,N_14217,N_12827);
and UO_1124 (O_1124,N_13023,N_13065);
nand UO_1125 (O_1125,N_11411,N_11441);
nor UO_1126 (O_1126,N_12702,N_10161);
and UO_1127 (O_1127,N_12989,N_13256);
nor UO_1128 (O_1128,N_14657,N_14000);
xor UO_1129 (O_1129,N_14769,N_10886);
nand UO_1130 (O_1130,N_13443,N_10111);
xnor UO_1131 (O_1131,N_12416,N_11615);
or UO_1132 (O_1132,N_14965,N_14779);
and UO_1133 (O_1133,N_12844,N_14494);
and UO_1134 (O_1134,N_10775,N_11356);
and UO_1135 (O_1135,N_14930,N_12265);
nand UO_1136 (O_1136,N_12846,N_11077);
and UO_1137 (O_1137,N_13102,N_12157);
nor UO_1138 (O_1138,N_12300,N_14602);
xor UO_1139 (O_1139,N_11146,N_11112);
nand UO_1140 (O_1140,N_13957,N_11578);
nor UO_1141 (O_1141,N_10336,N_10014);
or UO_1142 (O_1142,N_14461,N_10642);
xor UO_1143 (O_1143,N_10002,N_14559);
or UO_1144 (O_1144,N_14560,N_13027);
nand UO_1145 (O_1145,N_10737,N_10220);
nand UO_1146 (O_1146,N_14171,N_14047);
nand UO_1147 (O_1147,N_12322,N_10024);
and UO_1148 (O_1148,N_14854,N_12742);
nand UO_1149 (O_1149,N_13528,N_13660);
and UO_1150 (O_1150,N_14501,N_13470);
or UO_1151 (O_1151,N_10402,N_12454);
xor UO_1152 (O_1152,N_14362,N_13587);
xor UO_1153 (O_1153,N_10914,N_11419);
nor UO_1154 (O_1154,N_14787,N_14831);
and UO_1155 (O_1155,N_12070,N_11351);
xnor UO_1156 (O_1156,N_14402,N_11875);
xor UO_1157 (O_1157,N_11233,N_14375);
nor UO_1158 (O_1158,N_12522,N_13157);
nand UO_1159 (O_1159,N_14886,N_14508);
xnor UO_1160 (O_1160,N_14226,N_12185);
xnor UO_1161 (O_1161,N_14974,N_14578);
nand UO_1162 (O_1162,N_11398,N_10119);
and UO_1163 (O_1163,N_12189,N_12938);
or UO_1164 (O_1164,N_13564,N_13052);
nor UO_1165 (O_1165,N_14624,N_14874);
nor UO_1166 (O_1166,N_10686,N_11955);
or UO_1167 (O_1167,N_13613,N_12205);
or UO_1168 (O_1168,N_10307,N_12758);
nor UO_1169 (O_1169,N_13172,N_13004);
nor UO_1170 (O_1170,N_11794,N_12973);
nand UO_1171 (O_1171,N_14585,N_13186);
nor UO_1172 (O_1172,N_14009,N_14018);
nand UO_1173 (O_1173,N_11599,N_13058);
nor UO_1174 (O_1174,N_10800,N_13898);
xnor UO_1175 (O_1175,N_12319,N_11876);
nand UO_1176 (O_1176,N_11215,N_11927);
nor UO_1177 (O_1177,N_11031,N_13842);
or UO_1178 (O_1178,N_14072,N_11211);
and UO_1179 (O_1179,N_12583,N_13576);
xor UO_1180 (O_1180,N_12042,N_11493);
and UO_1181 (O_1181,N_14860,N_11767);
and UO_1182 (O_1182,N_14489,N_14542);
and UO_1183 (O_1183,N_12780,N_14917);
nand UO_1184 (O_1184,N_12151,N_12655);
or UO_1185 (O_1185,N_12694,N_11188);
and UO_1186 (O_1186,N_14537,N_10418);
xor UO_1187 (O_1187,N_14672,N_11868);
xor UO_1188 (O_1188,N_13455,N_10033);
or UO_1189 (O_1189,N_13026,N_11391);
nand UO_1190 (O_1190,N_11033,N_11624);
or UO_1191 (O_1191,N_11341,N_10962);
and UO_1192 (O_1192,N_10587,N_13430);
nor UO_1193 (O_1193,N_12513,N_11120);
xnor UO_1194 (O_1194,N_10295,N_12564);
nand UO_1195 (O_1195,N_13215,N_14969);
or UO_1196 (O_1196,N_13481,N_11986);
and UO_1197 (O_1197,N_13225,N_10803);
or UO_1198 (O_1198,N_10150,N_10151);
nor UO_1199 (O_1199,N_14757,N_10352);
or UO_1200 (O_1200,N_13488,N_14651);
xor UO_1201 (O_1201,N_10327,N_13667);
and UO_1202 (O_1202,N_10317,N_12018);
xnor UO_1203 (O_1203,N_13991,N_13325);
nand UO_1204 (O_1204,N_12760,N_10052);
xor UO_1205 (O_1205,N_11697,N_13332);
nand UO_1206 (O_1206,N_11445,N_14819);
or UO_1207 (O_1207,N_10433,N_10228);
and UO_1208 (O_1208,N_13232,N_12177);
and UO_1209 (O_1209,N_10225,N_11679);
or UO_1210 (O_1210,N_14745,N_10651);
or UO_1211 (O_1211,N_14002,N_12892);
or UO_1212 (O_1212,N_12951,N_10864);
nand UO_1213 (O_1213,N_14710,N_11584);
xnor UO_1214 (O_1214,N_12110,N_13240);
nand UO_1215 (O_1215,N_12250,N_12237);
xor UO_1216 (O_1216,N_10416,N_14572);
and UO_1217 (O_1217,N_11970,N_13379);
nand UO_1218 (O_1218,N_10820,N_10677);
nand UO_1219 (O_1219,N_13855,N_12996);
nand UO_1220 (O_1220,N_12504,N_12683);
or UO_1221 (O_1221,N_12138,N_13808);
xor UO_1222 (O_1222,N_11253,N_10693);
xor UO_1223 (O_1223,N_12825,N_14998);
nand UO_1224 (O_1224,N_14528,N_13809);
or UO_1225 (O_1225,N_14271,N_12058);
nand UO_1226 (O_1226,N_11399,N_14711);
nor UO_1227 (O_1227,N_14823,N_13664);
or UO_1228 (O_1228,N_14511,N_14377);
nand UO_1229 (O_1229,N_14832,N_13147);
nand UO_1230 (O_1230,N_10685,N_10040);
nor UO_1231 (O_1231,N_13306,N_12680);
or UO_1232 (O_1232,N_14221,N_10050);
nor UO_1233 (O_1233,N_13619,N_11780);
or UO_1234 (O_1234,N_11432,N_12816);
xnor UO_1235 (O_1235,N_10170,N_13919);
nor UO_1236 (O_1236,N_14458,N_11693);
nand UO_1237 (O_1237,N_14205,N_10042);
xnor UO_1238 (O_1238,N_11602,N_11855);
and UO_1239 (O_1239,N_13418,N_13880);
or UO_1240 (O_1240,N_10458,N_12593);
or UO_1241 (O_1241,N_13547,N_14488);
nand UO_1242 (O_1242,N_10857,N_13570);
nand UO_1243 (O_1243,N_10429,N_10349);
nor UO_1244 (O_1244,N_12885,N_12221);
nand UO_1245 (O_1245,N_11250,N_10617);
and UO_1246 (O_1246,N_13220,N_12376);
nor UO_1247 (O_1247,N_10212,N_14789);
xor UO_1248 (O_1248,N_12390,N_10036);
nor UO_1249 (O_1249,N_12855,N_13797);
or UO_1250 (O_1250,N_12182,N_11712);
xor UO_1251 (O_1251,N_11746,N_11307);
xor UO_1252 (O_1252,N_11245,N_12345);
xor UO_1253 (O_1253,N_14693,N_14749);
nand UO_1254 (O_1254,N_14129,N_12929);
nand UO_1255 (O_1255,N_12230,N_14258);
nand UO_1256 (O_1256,N_11346,N_10108);
or UO_1257 (O_1257,N_12797,N_10233);
or UO_1258 (O_1258,N_13390,N_12953);
and UO_1259 (O_1259,N_11290,N_13223);
xor UO_1260 (O_1260,N_11236,N_12638);
nor UO_1261 (O_1261,N_14344,N_13915);
or UO_1262 (O_1262,N_14768,N_10393);
xnor UO_1263 (O_1263,N_10554,N_11003);
and UO_1264 (O_1264,N_10892,N_14808);
xor UO_1265 (O_1265,N_10500,N_11545);
xnor UO_1266 (O_1266,N_10934,N_10044);
xnor UO_1267 (O_1267,N_12493,N_13750);
nand UO_1268 (O_1268,N_13652,N_10025);
or UO_1269 (O_1269,N_14524,N_14428);
nand UO_1270 (O_1270,N_12799,N_14368);
and UO_1271 (O_1271,N_12865,N_10986);
or UO_1272 (O_1272,N_14603,N_14195);
nand UO_1273 (O_1273,N_10653,N_11580);
xnor UO_1274 (O_1274,N_12971,N_10257);
nor UO_1275 (O_1275,N_13646,N_14876);
nor UO_1276 (O_1276,N_14689,N_12326);
xnor UO_1277 (O_1277,N_11040,N_13913);
and UO_1278 (O_1278,N_14963,N_12956);
and UO_1279 (O_1279,N_11788,N_12750);
nor UO_1280 (O_1280,N_13601,N_13675);
nand UO_1281 (O_1281,N_10439,N_13272);
xnor UO_1282 (O_1282,N_11199,N_11034);
or UO_1283 (O_1283,N_13623,N_14782);
nand UO_1284 (O_1284,N_11507,N_14975);
and UO_1285 (O_1285,N_11803,N_14093);
or UO_1286 (O_1286,N_11002,N_14135);
or UO_1287 (O_1287,N_14056,N_11840);
nor UO_1288 (O_1288,N_11837,N_12627);
and UO_1289 (O_1289,N_10403,N_14265);
and UO_1290 (O_1290,N_13760,N_13109);
or UO_1291 (O_1291,N_14253,N_12977);
and UO_1292 (O_1292,N_11117,N_13358);
or UO_1293 (O_1293,N_14937,N_12425);
nor UO_1294 (O_1294,N_10632,N_11258);
or UO_1295 (O_1295,N_12841,N_14310);
xor UO_1296 (O_1296,N_12127,N_12906);
nand UO_1297 (O_1297,N_14534,N_11450);
xor UO_1298 (O_1298,N_11321,N_13104);
and UO_1299 (O_1299,N_14287,N_14990);
nand UO_1300 (O_1300,N_11989,N_12711);
or UO_1301 (O_1301,N_10437,N_11706);
nand UO_1302 (O_1302,N_13969,N_14115);
xnor UO_1303 (O_1303,N_14935,N_11673);
xor UO_1304 (O_1304,N_10022,N_14960);
nand UO_1305 (O_1305,N_10717,N_12809);
nor UO_1306 (O_1306,N_11661,N_14007);
nand UO_1307 (O_1307,N_10097,N_11737);
nor UO_1308 (O_1308,N_13274,N_12657);
or UO_1309 (O_1309,N_12801,N_12056);
and UO_1310 (O_1310,N_10454,N_12943);
or UO_1311 (O_1311,N_10244,N_11682);
nor UO_1312 (O_1312,N_14037,N_10155);
nand UO_1313 (O_1313,N_12199,N_10088);
xnor UO_1314 (O_1314,N_10166,N_13593);
xnor UO_1315 (O_1315,N_14936,N_13063);
xnor UO_1316 (O_1316,N_13862,N_12011);
nand UO_1317 (O_1317,N_14882,N_12198);
or UO_1318 (O_1318,N_11933,N_14043);
or UO_1319 (O_1319,N_13537,N_13281);
xor UO_1320 (O_1320,N_11738,N_12466);
nor UO_1321 (O_1321,N_12761,N_10964);
or UO_1322 (O_1322,N_13557,N_11133);
or UO_1323 (O_1323,N_11467,N_10927);
xnor UO_1324 (O_1324,N_12507,N_11475);
nand UO_1325 (O_1325,N_14933,N_10946);
nand UO_1326 (O_1326,N_12736,N_10145);
nor UO_1327 (O_1327,N_12888,N_12069);
and UO_1328 (O_1328,N_10738,N_10739);
and UO_1329 (O_1329,N_11151,N_12361);
nand UO_1330 (O_1330,N_13286,N_10960);
xnor UO_1331 (O_1331,N_12713,N_10353);
or UO_1332 (O_1332,N_10140,N_13249);
xor UO_1333 (O_1333,N_11657,N_13007);
nand UO_1334 (O_1334,N_12878,N_10447);
xnor UO_1335 (O_1335,N_12531,N_13550);
nor UO_1336 (O_1336,N_13204,N_13929);
nor UO_1337 (O_1337,N_12912,N_12139);
and UO_1338 (O_1338,N_13722,N_13035);
nand UO_1339 (O_1339,N_12268,N_11639);
xnor UO_1340 (O_1340,N_10731,N_14407);
nand UO_1341 (O_1341,N_13965,N_14746);
xor UO_1342 (O_1342,N_12433,N_10552);
xnor UO_1343 (O_1343,N_13046,N_11065);
or UO_1344 (O_1344,N_13590,N_11416);
nor UO_1345 (O_1345,N_13573,N_12682);
or UO_1346 (O_1346,N_13451,N_12574);
nand UO_1347 (O_1347,N_12967,N_10217);
nor UO_1348 (O_1348,N_14814,N_13643);
xor UO_1349 (O_1349,N_12432,N_14001);
or UO_1350 (O_1350,N_10824,N_13752);
and UO_1351 (O_1351,N_13500,N_10798);
xor UO_1352 (O_1352,N_14676,N_11124);
nor UO_1353 (O_1353,N_12553,N_13755);
or UO_1354 (O_1354,N_14422,N_13165);
xnor UO_1355 (O_1355,N_14747,N_14111);
or UO_1356 (O_1356,N_10077,N_14538);
xor UO_1357 (O_1357,N_14577,N_11940);
xnor UO_1358 (O_1358,N_13375,N_11651);
and UO_1359 (O_1359,N_10465,N_13794);
nor UO_1360 (O_1360,N_12999,N_12914);
or UO_1361 (O_1361,N_11791,N_10847);
nand UO_1362 (O_1362,N_13705,N_12013);
or UO_1363 (O_1363,N_12930,N_12397);
nand UO_1364 (O_1364,N_14326,N_10165);
or UO_1365 (O_1365,N_13001,N_10628);
or UO_1366 (O_1366,N_12200,N_13663);
nor UO_1367 (O_1367,N_12413,N_12843);
nand UO_1368 (O_1368,N_11228,N_14485);
and UO_1369 (O_1369,N_14777,N_10613);
and UO_1370 (O_1370,N_14015,N_10839);
nor UO_1371 (O_1371,N_12351,N_10252);
xor UO_1372 (O_1372,N_12744,N_13987);
xnor UO_1373 (O_1373,N_14218,N_13746);
nand UO_1374 (O_1374,N_12836,N_12633);
or UO_1375 (O_1375,N_12339,N_14059);
and UO_1376 (O_1376,N_11429,N_11180);
nand UO_1377 (O_1377,N_10703,N_11517);
nand UO_1378 (O_1378,N_14482,N_10188);
nand UO_1379 (O_1379,N_10519,N_13936);
nor UO_1380 (O_1380,N_13189,N_10277);
xnor UO_1381 (O_1381,N_14144,N_10421);
nand UO_1382 (O_1382,N_11676,N_12451);
xor UO_1383 (O_1383,N_10016,N_11831);
nor UO_1384 (O_1384,N_14905,N_11234);
and UO_1385 (O_1385,N_12252,N_11300);
or UO_1386 (O_1386,N_10172,N_12160);
xnor UO_1387 (O_1387,N_14999,N_11221);
xnor UO_1388 (O_1388,N_13083,N_13498);
nor UO_1389 (O_1389,N_10789,N_14827);
and UO_1390 (O_1390,N_12532,N_11536);
and UO_1391 (O_1391,N_14794,N_13860);
nand UO_1392 (O_1392,N_12544,N_12520);
nand UO_1393 (O_1393,N_12109,N_13403);
or UO_1394 (O_1394,N_12096,N_13140);
and UO_1395 (O_1395,N_12634,N_11765);
and UO_1396 (O_1396,N_10198,N_14095);
and UO_1397 (O_1397,N_13869,N_13099);
nand UO_1398 (O_1398,N_11526,N_12712);
and UO_1399 (O_1399,N_13641,N_14153);
and UO_1400 (O_1400,N_12631,N_12315);
and UO_1401 (O_1401,N_12485,N_14244);
nand UO_1402 (O_1402,N_14150,N_10650);
nand UO_1403 (O_1403,N_13340,N_14383);
and UO_1404 (O_1404,N_13807,N_10959);
nor UO_1405 (O_1405,N_12916,N_12555);
nand UO_1406 (O_1406,N_14504,N_10854);
xor UO_1407 (O_1407,N_14353,N_11373);
nor UO_1408 (O_1408,N_12950,N_14314);
xnor UO_1409 (O_1409,N_11943,N_10919);
or UO_1410 (O_1410,N_13075,N_12645);
nor UO_1411 (O_1411,N_13180,N_10532);
and UO_1412 (O_1412,N_14934,N_10660);
nand UO_1413 (O_1413,N_14704,N_12747);
nand UO_1414 (O_1414,N_13569,N_12026);
and UO_1415 (O_1415,N_10342,N_13770);
nor UO_1416 (O_1416,N_12729,N_14252);
and UO_1417 (O_1417,N_12393,N_13176);
nand UO_1418 (O_1418,N_12601,N_12882);
xor UO_1419 (O_1419,N_10910,N_13820);
xnor UO_1420 (O_1420,N_12225,N_10321);
nor UO_1421 (O_1421,N_14523,N_12120);
xor UO_1422 (O_1422,N_13735,N_14752);
xnor UO_1423 (O_1423,N_10558,N_13521);
and UO_1424 (O_1424,N_10531,N_14914);
nand UO_1425 (O_1425,N_11200,N_11367);
nor UO_1426 (O_1426,N_14477,N_12295);
nand UO_1427 (O_1427,N_13692,N_14932);
or UO_1428 (O_1428,N_14172,N_12389);
and UO_1429 (O_1429,N_14956,N_13821);
xnor UO_1430 (O_1430,N_11297,N_10448);
or UO_1431 (O_1431,N_11136,N_11424);
or UO_1432 (O_1432,N_11311,N_14867);
nand UO_1433 (O_1433,N_12598,N_13424);
xnor UO_1434 (O_1434,N_14866,N_12418);
xnor UO_1435 (O_1435,N_14967,N_14713);
nor UO_1436 (O_1436,N_14629,N_12806);
nor UO_1437 (O_1437,N_10969,N_12959);
nor UO_1438 (O_1438,N_11962,N_14637);
xnor UO_1439 (O_1439,N_14275,N_14213);
nand UO_1440 (O_1440,N_12556,N_13510);
and UO_1441 (O_1441,N_11611,N_12388);
or UO_1442 (O_1442,N_14652,N_12700);
and UO_1443 (O_1443,N_11023,N_12309);
nor UO_1444 (O_1444,N_10471,N_13393);
nand UO_1445 (O_1445,N_11102,N_13962);
xnor UO_1446 (O_1446,N_10494,N_12802);
or UO_1447 (O_1447,N_13865,N_11630);
nor UO_1448 (O_1448,N_11662,N_11574);
or UO_1449 (O_1449,N_11809,N_13977);
and UO_1450 (O_1450,N_12641,N_14716);
or UO_1451 (O_1451,N_12242,N_12635);
and UO_1452 (O_1452,N_11948,N_10687);
nor UO_1453 (O_1453,N_12654,N_10436);
nand UO_1454 (O_1454,N_10414,N_12835);
and UO_1455 (O_1455,N_10434,N_11090);
xor UO_1456 (O_1456,N_13901,N_12871);
nand UO_1457 (O_1457,N_13785,N_13177);
nand UO_1458 (O_1458,N_10624,N_13907);
nand UO_1459 (O_1459,N_14635,N_13383);
nand UO_1460 (O_1460,N_11400,N_11909);
and UO_1461 (O_1461,N_11898,N_14798);
xnor UO_1462 (O_1462,N_10511,N_10838);
nand UO_1463 (O_1463,N_12862,N_12175);
nor UO_1464 (O_1464,N_12961,N_14759);
nor UO_1465 (O_1465,N_10948,N_10672);
nand UO_1466 (O_1466,N_13089,N_14008);
or UO_1467 (O_1467,N_14811,N_11721);
or UO_1468 (O_1468,N_14878,N_11235);
and UO_1469 (O_1469,N_10905,N_13191);
nor UO_1470 (O_1470,N_12465,N_13265);
nand UO_1471 (O_1471,N_12077,N_10828);
nand UO_1472 (O_1472,N_12165,N_11717);
nand UO_1473 (O_1473,N_14973,N_10269);
nand UO_1474 (O_1474,N_10048,N_14985);
and UO_1475 (O_1475,N_10364,N_11839);
xor UO_1476 (O_1476,N_11306,N_11036);
or UO_1477 (O_1477,N_13209,N_13478);
or UO_1478 (O_1478,N_10578,N_12461);
nand UO_1479 (O_1479,N_12650,N_12792);
nand UO_1480 (O_1480,N_11365,N_14496);
or UO_1481 (O_1481,N_13125,N_12643);
or UO_1482 (O_1482,N_12090,N_14122);
nor UO_1483 (O_1483,N_14846,N_13414);
nand UO_1484 (O_1484,N_11654,N_13926);
xnor UO_1485 (O_1485,N_14229,N_10273);
nor UO_1486 (O_1486,N_11836,N_13578);
nor UO_1487 (O_1487,N_14215,N_12124);
xnor UO_1488 (O_1488,N_14997,N_12354);
xnor UO_1489 (O_1489,N_11008,N_13028);
xnor UO_1490 (O_1490,N_11192,N_12075);
nor UO_1491 (O_1491,N_10303,N_10711);
and UO_1492 (O_1492,N_10521,N_12624);
or UO_1493 (O_1493,N_14582,N_13922);
and UO_1494 (O_1494,N_14162,N_12584);
or UO_1495 (O_1495,N_10146,N_13184);
nor UO_1496 (O_1496,N_11108,N_14893);
and UO_1497 (O_1497,N_13350,N_14490);
or UO_1498 (O_1498,N_13932,N_13289);
nand UO_1499 (O_1499,N_12629,N_12186);
nor UO_1500 (O_1500,N_10158,N_11029);
or UO_1501 (O_1501,N_13850,N_11953);
xnor UO_1502 (O_1502,N_13996,N_14531);
or UO_1503 (O_1503,N_10782,N_10884);
nand UO_1504 (O_1504,N_14948,N_13796);
nor UO_1505 (O_1505,N_10736,N_14526);
nand UO_1506 (O_1506,N_14459,N_12637);
or UO_1507 (O_1507,N_14743,N_11182);
nand UO_1508 (O_1508,N_12392,N_14013);
xnor UO_1509 (O_1509,N_14549,N_10297);
or UO_1510 (O_1510,N_14836,N_11279);
nor UO_1511 (O_1511,N_13868,N_12632);
nor UO_1512 (O_1512,N_13758,N_11786);
nor UO_1513 (O_1513,N_14405,N_10290);
and UO_1514 (O_1514,N_10441,N_12726);
nor UO_1515 (O_1515,N_13633,N_13322);
nand UO_1516 (O_1516,N_11056,N_12038);
xnor UO_1517 (O_1517,N_13950,N_13879);
nand UO_1518 (O_1518,N_11828,N_10095);
nor UO_1519 (O_1519,N_10668,N_14280);
nand UO_1520 (O_1520,N_12763,N_13468);
xor UO_1521 (O_1521,N_12238,N_11719);
or UO_1522 (O_1522,N_13370,N_14994);
or UO_1523 (O_1523,N_14284,N_14374);
or UO_1524 (O_1524,N_12670,N_11407);
or UO_1525 (O_1525,N_11172,N_11067);
nand UO_1526 (O_1526,N_13721,N_14539);
and UO_1527 (O_1527,N_13930,N_12161);
nor UO_1528 (O_1528,N_11109,N_13062);
xor UO_1529 (O_1529,N_11915,N_10462);
and UO_1530 (O_1530,N_14995,N_10967);
nor UO_1531 (O_1531,N_13178,N_11914);
nand UO_1532 (O_1532,N_12283,N_10580);
or UO_1533 (O_1533,N_11957,N_12503);
or UO_1534 (O_1534,N_13647,N_11007);
nand UO_1535 (O_1535,N_10858,N_10865);
nor UO_1536 (O_1536,N_13059,N_11726);
or UO_1537 (O_1537,N_11963,N_14464);
xor UO_1538 (O_1538,N_12510,N_11896);
and UO_1539 (O_1539,N_14068,N_10422);
or UO_1540 (O_1540,N_12405,N_13162);
nor UO_1541 (O_1541,N_14822,N_14568);
or UO_1542 (O_1542,N_14776,N_10080);
nand UO_1543 (O_1543,N_11604,N_10041);
nor UO_1544 (O_1544,N_11089,N_12400);
nand UO_1545 (O_1545,N_13740,N_13640);
nor UO_1546 (O_1546,N_12909,N_13534);
nor UO_1547 (O_1547,N_11169,N_11817);
and UO_1548 (O_1548,N_14260,N_10900);
and UO_1549 (O_1549,N_10897,N_12204);
xnor UO_1550 (O_1550,N_11171,N_13751);
or UO_1551 (O_1551,N_10319,N_11041);
nor UO_1552 (O_1552,N_14175,N_13863);
nor UO_1553 (O_1553,N_14370,N_12773);
xor UO_1554 (O_1554,N_14992,N_12246);
or UO_1555 (O_1555,N_12027,N_10743);
nor UO_1556 (O_1556,N_12732,N_13237);
or UO_1557 (O_1557,N_12220,N_14481);
nand UO_1558 (O_1558,N_14793,N_10068);
nor UO_1559 (O_1559,N_14003,N_10423);
xor UO_1560 (O_1560,N_10852,N_11322);
and UO_1561 (O_1561,N_11328,N_12547);
nor UO_1562 (O_1562,N_14639,N_14197);
or UO_1563 (O_1563,N_12006,N_11764);
xor UO_1564 (O_1564,N_12380,N_13245);
xor UO_1565 (O_1565,N_13433,N_14622);
or UO_1566 (O_1566,N_11327,N_13747);
or UO_1567 (O_1567,N_12847,N_10313);
or UO_1568 (O_1568,N_14082,N_11716);
nor UO_1569 (O_1569,N_12031,N_12893);
nand UO_1570 (O_1570,N_11213,N_12362);
nand UO_1571 (O_1571,N_13236,N_12359);
nor UO_1572 (O_1572,N_10649,N_10831);
xnor UO_1573 (O_1573,N_14857,N_13417);
nor UO_1574 (O_1574,N_14062,N_12990);
nor UO_1575 (O_1575,N_12370,N_10425);
nand UO_1576 (O_1576,N_13574,N_12705);
nand UO_1577 (O_1577,N_10470,N_14462);
and UO_1578 (O_1578,N_12884,N_11179);
or UO_1579 (O_1579,N_14695,N_12771);
nor UO_1580 (O_1580,N_12810,N_12227);
xor UO_1581 (O_1581,N_10308,N_12860);
nor UO_1582 (O_1582,N_10689,N_10272);
nor UO_1583 (O_1583,N_10601,N_11995);
or UO_1584 (O_1584,N_12499,N_13315);
nor UO_1585 (O_1585,N_13141,N_13506);
and UO_1586 (O_1586,N_11038,N_13699);
nor UO_1587 (O_1587,N_10887,N_10805);
or UO_1588 (O_1588,N_11971,N_14543);
xnor UO_1589 (O_1589,N_13304,N_13173);
xnor UO_1590 (O_1590,N_11736,N_11689);
nand UO_1591 (O_1591,N_13669,N_10265);
or UO_1592 (O_1592,N_13067,N_13812);
xnor UO_1593 (O_1593,N_11906,N_14641);
xnor UO_1594 (O_1594,N_12306,N_13852);
nor UO_1595 (O_1595,N_14770,N_13565);
nor UO_1596 (O_1596,N_13103,N_12162);
xor UO_1597 (O_1597,N_10678,N_14491);
nor UO_1598 (O_1598,N_13843,N_12297);
nor UO_1599 (O_1599,N_11873,N_10727);
xnor UO_1600 (O_1600,N_11695,N_10469);
xnor UO_1601 (O_1601,N_12112,N_11015);
nor UO_1602 (O_1602,N_12554,N_11461);
or UO_1603 (O_1603,N_12753,N_13781);
nand UO_1604 (O_1604,N_13911,N_10032);
or UO_1605 (O_1605,N_10379,N_13160);
xor UO_1606 (O_1606,N_14691,N_14356);
nand UO_1607 (O_1607,N_14613,N_13294);
xnor UO_1608 (O_1608,N_12539,N_12039);
or UO_1609 (O_1609,N_11972,N_13805);
and UO_1610 (O_1610,N_10796,N_12936);
and UO_1611 (O_1611,N_14647,N_12333);
or UO_1612 (O_1612,N_12000,N_13070);
nor UO_1613 (O_1613,N_12693,N_13360);
xor UO_1614 (O_1614,N_12778,N_14795);
nor UO_1615 (O_1615,N_11804,N_10058);
nor UO_1616 (O_1616,N_14292,N_10641);
nand UO_1617 (O_1617,N_11173,N_14735);
xor UO_1618 (O_1618,N_12012,N_12401);
nand UO_1619 (O_1619,N_14889,N_14480);
nand UO_1620 (O_1620,N_10356,N_11600);
and UO_1621 (O_1621,N_10110,N_10498);
xnor UO_1622 (O_1622,N_12735,N_14166);
nand UO_1623 (O_1623,N_11763,N_13397);
or UO_1624 (O_1624,N_13545,N_13066);
xnor UO_1625 (O_1625,N_12506,N_12558);
and UO_1626 (O_1626,N_13712,N_14594);
nor UO_1627 (O_1627,N_13549,N_10154);
xnor UO_1628 (O_1628,N_13193,N_10809);
xnor UO_1629 (O_1629,N_14304,N_13395);
nand UO_1630 (O_1630,N_11415,N_11560);
and UO_1631 (O_1631,N_14702,N_13953);
nor UO_1632 (O_1632,N_11869,N_11278);
nand UO_1633 (O_1633,N_11141,N_13836);
and UO_1634 (O_1634,N_13221,N_13453);
or UO_1635 (O_1635,N_13371,N_14409);
xor UO_1636 (O_1636,N_14616,N_12546);
and UO_1637 (O_1637,N_13197,N_12346);
nor UO_1638 (O_1638,N_11379,N_13015);
nand UO_1639 (O_1639,N_13190,N_10625);
and UO_1640 (O_1640,N_12324,N_11464);
nand UO_1641 (O_1641,N_14355,N_10752);
xor UO_1642 (O_1642,N_13212,N_10833);
xor UO_1643 (O_1643,N_11593,N_12121);
nor UO_1644 (O_1644,N_10126,N_14563);
nand UO_1645 (O_1645,N_12687,N_11268);
nor UO_1646 (O_1646,N_14852,N_12652);
nand UO_1647 (O_1647,N_10562,N_14606);
or UO_1648 (O_1648,N_10714,N_10928);
xnor UO_1649 (O_1649,N_14306,N_10260);
xnor UO_1650 (O_1650,N_13595,N_12277);
nor UO_1651 (O_1651,N_12173,N_14922);
or UO_1652 (O_1652,N_12149,N_10875);
xnor UO_1653 (O_1653,N_13480,N_12076);
nor UO_1654 (O_1654,N_11530,N_13489);
nor UO_1655 (O_1655,N_14818,N_12438);
xnor UO_1656 (O_1656,N_12708,N_11710);
and UO_1657 (O_1657,N_11075,N_14725);
xnor UO_1658 (O_1658,N_14382,N_14517);
xor UO_1659 (O_1659,N_10997,N_12299);
nand UO_1660 (O_1660,N_12848,N_11301);
nand UO_1661 (O_1661,N_12829,N_14927);
xnor UO_1662 (O_1662,N_11851,N_10029);
and UO_1663 (O_1663,N_11848,N_14380);
nand UO_1664 (O_1664,N_13119,N_14731);
nand UO_1665 (O_1665,N_12667,N_11042);
xor UO_1666 (O_1666,N_10207,N_12460);
xnor UO_1667 (O_1667,N_10325,N_14871);
nor UO_1668 (O_1668,N_10181,N_10147);
nand UO_1669 (O_1669,N_10545,N_11832);
nor UO_1670 (O_1670,N_12926,N_11005);
xnor UO_1671 (O_1671,N_10339,N_13726);
xor UO_1672 (O_1672,N_10810,N_11918);
or UO_1673 (O_1673,N_12559,N_13400);
or UO_1674 (O_1674,N_13471,N_12665);
xnor UO_1675 (O_1675,N_12458,N_11824);
and UO_1676 (O_1676,N_14442,N_14664);
xor UO_1677 (O_1677,N_13733,N_10656);
and UO_1678 (O_1678,N_10933,N_14439);
or UO_1679 (O_1679,N_12621,N_12822);
nand UO_1680 (O_1680,N_13955,N_11061);
or UO_1681 (O_1681,N_12737,N_11787);
nand UO_1682 (O_1682,N_12599,N_11859);
xnor UO_1683 (O_1683,N_12373,N_14856);
nand UO_1684 (O_1684,N_11191,N_14285);
and UO_1685 (O_1685,N_10129,N_11759);
nor UO_1686 (O_1686,N_10113,N_13513);
nor UO_1687 (O_1687,N_11159,N_10493);
nand UO_1688 (O_1688,N_10340,N_12007);
xnor UO_1689 (O_1689,N_10890,N_13730);
nand UO_1690 (O_1690,N_13386,N_13078);
xor UO_1691 (O_1691,N_14561,N_13263);
and UO_1692 (O_1692,N_10729,N_10778);
xnor UO_1693 (O_1693,N_14479,N_11039);
nor UO_1694 (O_1694,N_12804,N_13139);
nand UO_1695 (O_1695,N_11276,N_13144);
or UO_1696 (O_1696,N_12787,N_12872);
and UO_1697 (O_1697,N_12279,N_11374);
nand UO_1698 (O_1698,N_12945,N_11395);
nor UO_1699 (O_1699,N_14237,N_13561);
nand UO_1700 (O_1700,N_11537,N_10264);
nor UO_1701 (O_1701,N_12777,N_12548);
and UO_1702 (O_1702,N_14571,N_13288);
nor UO_1703 (O_1703,N_14350,N_11332);
nand UO_1704 (O_1704,N_13473,N_13984);
and UO_1705 (O_1705,N_14117,N_14064);
nor UO_1706 (O_1706,N_11829,N_13753);
nor UO_1707 (O_1707,N_13499,N_14632);
nor UO_1708 (O_1708,N_11472,N_12021);
or UO_1709 (O_1709,N_11628,N_13829);
nor UO_1710 (O_1710,N_13310,N_14721);
or UO_1711 (O_1711,N_13449,N_10980);
nand UO_1712 (O_1712,N_12981,N_12985);
or UO_1713 (O_1713,N_11209,N_10103);
nand UO_1714 (O_1714,N_14663,N_13558);
xor UO_1715 (O_1715,N_14156,N_14645);
nand UO_1716 (O_1716,N_12081,N_13600);
nand UO_1717 (O_1717,N_10987,N_14212);
nor UO_1718 (O_1718,N_11378,N_11633);
xor UO_1719 (O_1719,N_13620,N_10898);
nor UO_1720 (O_1720,N_10136,N_12676);
nor UO_1721 (O_1721,N_13540,N_14712);
nand UO_1722 (O_1722,N_13771,N_11487);
and UO_1723 (O_1723,N_14708,N_12085);
nor UO_1724 (O_1724,N_12854,N_12661);
or UO_1725 (O_1725,N_13949,N_10834);
xnor UO_1726 (O_1726,N_13352,N_11186);
nand UO_1727 (O_1727,N_13098,N_12642);
nand UO_1728 (O_1728,N_11757,N_11877);
nand UO_1729 (O_1729,N_10109,N_11703);
or UO_1730 (O_1730,N_13830,N_10692);
or UO_1731 (O_1731,N_11991,N_14365);
and UO_1732 (O_1732,N_12970,N_13331);
and UO_1733 (O_1733,N_10732,N_13218);
xor UO_1734 (O_1734,N_13525,N_11776);
and UO_1735 (O_1735,N_12610,N_11707);
xor UO_1736 (O_1736,N_12751,N_14133);
nor UO_1737 (O_1737,N_11616,N_13597);
and UO_1738 (O_1738,N_10804,N_12321);
or UO_1739 (O_1739,N_13159,N_14300);
nor UO_1740 (O_1740,N_11017,N_12567);
nand UO_1741 (O_1741,N_13773,N_11078);
and UO_1742 (O_1742,N_10415,N_11433);
nor UO_1743 (O_1743,N_11074,N_11043);
nor UO_1744 (O_1744,N_13790,N_13963);
xor UO_1745 (O_1745,N_10565,N_10299);
nand UO_1746 (O_1746,N_12842,N_11128);
nor UO_1747 (O_1747,N_11292,N_11364);
nor UO_1748 (O_1748,N_14371,N_12188);
and UO_1749 (O_1749,N_12757,N_11280);
or UO_1750 (O_1750,N_12689,N_14385);
xnor UO_1751 (O_1751,N_10526,N_11338);
nor UO_1752 (O_1752,N_14556,N_10208);
nand UO_1753 (O_1753,N_12317,N_14780);
xor UO_1754 (O_1754,N_10305,N_14742);
xor UO_1755 (O_1755,N_14869,N_10061);
nor UO_1756 (O_1756,N_13689,N_14131);
or UO_1757 (O_1757,N_12630,N_11558);
and UO_1758 (O_1758,N_13920,N_10351);
and UO_1759 (O_1759,N_11296,N_12419);
xnor UO_1760 (O_1760,N_12918,N_12014);
xor UO_1761 (O_1761,N_14566,N_11052);
and UO_1762 (O_1762,N_14169,N_13881);
xnor UO_1763 (O_1763,N_10253,N_14492);
nor UO_1764 (O_1764,N_12231,N_14668);
nor UO_1765 (O_1765,N_13259,N_14507);
and UO_1766 (O_1766,N_11156,N_14016);
xnor UO_1767 (O_1767,N_14684,N_11165);
nand UO_1768 (O_1768,N_11535,N_10463);
nor UO_1769 (O_1769,N_14617,N_11106);
xnor UO_1770 (O_1770,N_14929,N_11792);
or UO_1771 (O_1771,N_12034,N_13767);
and UO_1772 (O_1772,N_14165,N_10675);
xnor UO_1773 (O_1773,N_12782,N_12919);
nand UO_1774 (O_1774,N_13895,N_14201);
or UO_1775 (O_1775,N_11754,N_10947);
xor UO_1776 (O_1776,N_10888,N_14176);
nand UO_1777 (O_1777,N_13199,N_11057);
or UO_1778 (O_1778,N_14039,N_10944);
or UO_1779 (O_1779,N_14848,N_14979);
nor UO_1780 (O_1780,N_11974,N_12074);
or UO_1781 (O_1781,N_10163,N_14296);
and UO_1782 (O_1782,N_10658,N_11932);
nand UO_1783 (O_1783,N_11501,N_14828);
xor UO_1784 (O_1784,N_11812,N_13766);
or UO_1785 (O_1785,N_14154,N_10189);
and UO_1786 (O_1786,N_10881,N_13720);
nor UO_1787 (O_1787,N_10556,N_10826);
nand UO_1788 (O_1788,N_13931,N_12767);
nand UO_1789 (O_1789,N_11035,N_10657);
xnor UO_1790 (O_1790,N_14669,N_11850);
nand UO_1791 (O_1791,N_11175,N_10392);
or UO_1792 (O_1792,N_10078,N_14463);
nand UO_1793 (O_1793,N_11428,N_13192);
xor UO_1794 (O_1794,N_14962,N_10345);
nand UO_1795 (O_1795,N_10990,N_14317);
nand UO_1796 (O_1796,N_13462,N_12020);
and UO_1797 (O_1797,N_11494,N_12086);
or UO_1798 (O_1798,N_12704,N_14460);
and UO_1799 (O_1799,N_14148,N_13970);
xor UO_1800 (O_1800,N_13628,N_10976);
or UO_1801 (O_1801,N_12128,N_12538);
or UO_1802 (O_1802,N_11114,N_13899);
nand UO_1803 (O_1803,N_11275,N_13434);
nor UO_1804 (O_1804,N_13000,N_12811);
and UO_1805 (O_1805,N_10291,N_10445);
or UO_1806 (O_1806,N_10961,N_14034);
xor UO_1807 (O_1807,N_13937,N_11382);
and UO_1808 (O_1808,N_13039,N_11671);
nor UO_1809 (O_1809,N_12511,N_10788);
nand UO_1810 (O_1810,N_11006,N_10744);
nor UO_1811 (O_1811,N_13677,N_12353);
and UO_1812 (O_1812,N_11864,N_10655);
nor UO_1813 (O_1813,N_14865,N_13804);
nor UO_1814 (O_1814,N_12107,N_14184);
and UO_1815 (O_1815,N_11026,N_13391);
or UO_1816 (O_1816,N_14267,N_14980);
nor UO_1817 (O_1817,N_12807,N_12830);
nor UO_1818 (O_1818,N_13270,N_11960);
and UO_1819 (O_1819,N_14553,N_11741);
xnor UO_1820 (O_1820,N_12721,N_13612);
or UO_1821 (O_1821,N_13979,N_13211);
xnor UO_1822 (O_1822,N_14513,N_12776);
nor UO_1823 (O_1823,N_12015,N_10718);
xnor UO_1824 (O_1824,N_10359,N_14214);
and UO_1825 (O_1825,N_12620,N_12394);
nor UO_1826 (O_1826,N_14393,N_14844);
or UO_1827 (O_1827,N_12897,N_14996);
and UO_1828 (O_1828,N_11140,N_14987);
nand UO_1829 (O_1829,N_10627,N_11608);
nand UO_1830 (O_1830,N_11908,N_10570);
nor UO_1831 (O_1831,N_14473,N_13803);
nand UO_1832 (O_1832,N_11104,N_13452);
or UO_1833 (O_1833,N_13456,N_13556);
and UO_1834 (O_1834,N_10182,N_12623);
nor UO_1835 (O_1835,N_13530,N_14989);
xor UO_1836 (O_1836,N_10582,N_13883);
xor UO_1837 (O_1837,N_10935,N_12310);
and UO_1838 (O_1838,N_10735,N_14991);
nand UO_1839 (O_1839,N_13887,N_11363);
and UO_1840 (O_1840,N_14557,N_10400);
and UO_1841 (O_1841,N_13117,N_14909);
nand UO_1842 (O_1842,N_10566,N_14211);
or UO_1843 (O_1843,N_14147,N_13129);
and UO_1844 (O_1844,N_12515,N_10281);
nor UO_1845 (O_1845,N_10169,N_10245);
xor UO_1846 (O_1846,N_10932,N_11241);
and UO_1847 (O_1847,N_11571,N_10366);
nand UO_1848 (O_1848,N_11269,N_10509);
nand UO_1849 (O_1849,N_12502,N_13621);
and UO_1850 (O_1850,N_10648,N_10338);
xor UO_1851 (O_1851,N_11987,N_14081);
or UO_1852 (O_1852,N_11944,N_14437);
and UO_1853 (O_1853,N_14945,N_11680);
nor UO_1854 (O_1854,N_13765,N_14833);
nand UO_1855 (O_1855,N_10750,N_13361);
and UO_1856 (O_1856,N_13493,N_13253);
and UO_1857 (O_1857,N_12083,N_13483);
and UO_1858 (O_1858,N_11402,N_10640);
xnor UO_1859 (O_1859,N_12924,N_10368);
and UO_1860 (O_1860,N_13859,N_11762);
or UO_1861 (O_1861,N_14558,N_14467);
and UO_1862 (O_1862,N_11434,N_11961);
or UO_1863 (O_1863,N_12869,N_12184);
and UO_1864 (O_1864,N_14850,N_14055);
or UO_1865 (O_1865,N_12239,N_12958);
xor UO_1866 (O_1866,N_14626,N_12762);
xnor UO_1867 (O_1867,N_13381,N_14448);
nor UO_1868 (O_1868,N_10394,N_12701);
xor UO_1869 (O_1869,N_13198,N_13248);
nand UO_1870 (O_1870,N_13980,N_14890);
nand UO_1871 (O_1871,N_12921,N_11094);
and UO_1872 (O_1872,N_13441,N_11093);
xnor UO_1873 (O_1873,N_13415,N_11610);
nor UO_1874 (O_1874,N_11163,N_12445);
nor UO_1875 (O_1875,N_12381,N_12292);
and UO_1876 (O_1876,N_12336,N_11691);
xnor UO_1877 (O_1877,N_13783,N_10953);
xnor UO_1878 (O_1878,N_12741,N_10992);
or UO_1879 (O_1879,N_10879,N_14089);
and UO_1880 (O_1880,N_14294,N_13024);
xor UO_1881 (O_1881,N_13694,N_13904);
xnor UO_1882 (O_1882,N_10591,N_13239);
xor UO_1883 (O_1883,N_11316,N_13988);
and UO_1884 (O_1884,N_13986,N_13343);
xor UO_1885 (O_1885,N_11684,N_14688);
and UO_1886 (O_1886,N_11299,N_12814);
and UO_1887 (O_1887,N_12349,N_12259);
nor UO_1888 (O_1888,N_11777,N_10618);
xnor UO_1889 (O_1889,N_10399,N_13952);
or UO_1890 (O_1890,N_13048,N_14004);
xor UO_1891 (O_1891,N_12481,N_13529);
nand UO_1892 (O_1892,N_14248,N_12008);
nor UO_1893 (O_1893,N_11166,N_12840);
and UO_1894 (O_1894,N_12993,N_10970);
nor UO_1895 (O_1895,N_13224,N_13092);
or UO_1896 (O_1896,N_14767,N_12784);
or UO_1897 (O_1897,N_13427,N_14754);
or UO_1898 (O_1898,N_10665,N_10576);
or UO_1899 (O_1899,N_13372,N_12063);
nor UO_1900 (O_1900,N_14801,N_12851);
nand UO_1901 (O_1901,N_14545,N_11406);
nor UO_1902 (O_1902,N_11205,N_10740);
xor UO_1903 (O_1903,N_13170,N_13945);
nor UO_1904 (O_1904,N_11255,N_10031);
nand UO_1905 (O_1905,N_11660,N_14536);
or UO_1906 (O_1906,N_12414,N_10261);
xor UO_1907 (O_1907,N_10114,N_12384);
nor UO_1908 (O_1908,N_12142,N_13799);
xor UO_1909 (O_1909,N_14636,N_12852);
or UO_1910 (O_1910,N_11825,N_10209);
and UO_1911 (O_1911,N_12944,N_11474);
xnor UO_1912 (O_1912,N_13947,N_10466);
and UO_1913 (O_1913,N_10984,N_11567);
or UO_1914 (O_1914,N_12366,N_13934);
nand UO_1915 (O_1915,N_13896,N_12290);
nand UO_1916 (O_1916,N_13975,N_12883);
xor UO_1917 (O_1917,N_13638,N_11644);
or UO_1918 (O_1918,N_10630,N_12730);
and UO_1919 (O_1919,N_14520,N_14758);
or UO_1920 (O_1920,N_10302,N_14334);
and UO_1921 (O_1921,N_11488,N_12733);
nor UO_1922 (O_1922,N_10176,N_13672);
xor UO_1923 (O_1923,N_11993,N_11895);
xor UO_1924 (O_1924,N_13795,N_10542);
nand UO_1925 (O_1925,N_11021,N_10747);
or UO_1926 (O_1926,N_11638,N_10125);
xor UO_1927 (O_1927,N_11295,N_10851);
nor UO_1928 (O_1928,N_10802,N_12172);
xnor UO_1929 (O_1929,N_14597,N_11865);
and UO_1930 (O_1930,N_11059,N_12664);
and UO_1931 (O_1931,N_13040,N_14946);
xor UO_1932 (O_1932,N_14949,N_12271);
nor UO_1933 (O_1933,N_13943,N_10412);
or UO_1934 (O_1934,N_11149,N_12500);
and UO_1935 (O_1935,N_11252,N_13445);
nand UO_1936 (O_1936,N_14143,N_12377);
xnor UO_1937 (O_1937,N_13234,N_12669);
and UO_1938 (O_1938,N_10866,N_11811);
nor UO_1939 (O_1939,N_14359,N_10231);
or UO_1940 (O_1940,N_11446,N_12984);
nand UO_1941 (O_1941,N_12163,N_11314);
and UO_1942 (O_1942,N_13163,N_12212);
nor UO_1943 (O_1943,N_10039,N_12939);
and UO_1944 (O_1944,N_13688,N_13893);
xnor UO_1945 (O_1945,N_12261,N_10354);
nor UO_1946 (O_1946,N_14227,N_13262);
xor UO_1947 (O_1947,N_11463,N_10827);
xor UO_1948 (O_1948,N_10043,N_12057);
nor UO_1949 (O_1949,N_11795,N_12910);
and UO_1950 (O_1950,N_12154,N_11492);
or UO_1951 (O_1951,N_10758,N_11635);
xor UO_1952 (O_1952,N_12572,N_11386);
xor UO_1953 (O_1953,N_13341,N_14078);
nand UO_1954 (O_1954,N_14705,N_14305);
or UO_1955 (O_1955,N_10768,N_14158);
or UO_1956 (O_1956,N_12216,N_13704);
and UO_1957 (O_1957,N_11412,N_14225);
nor UO_1958 (O_1958,N_14339,N_10533);
nor UO_1959 (O_1959,N_12313,N_10213);
and UO_1960 (O_1960,N_14620,N_11709);
nand UO_1961 (O_1961,N_12934,N_12997);
xor UO_1962 (O_1962,N_14046,N_13714);
nor UO_1963 (O_1963,N_10590,N_12496);
or UO_1964 (O_1964,N_13095,N_14065);
and UO_1965 (O_1965,N_10232,N_10064);
nor UO_1966 (O_1966,N_13188,N_13309);
xor UO_1967 (O_1967,N_11262,N_13656);
and UO_1968 (O_1968,N_11266,N_11694);
xnor UO_1969 (O_1969,N_12991,N_11674);
nand UO_1970 (O_1970,N_13853,N_14223);
nor UO_1971 (O_1971,N_10937,N_11846);
or UO_1972 (O_1972,N_14674,N_13019);
nand UO_1973 (O_1973,N_11586,N_12779);
or UO_1974 (O_1974,N_11509,N_14499);
xor UO_1975 (O_1975,N_12044,N_12183);
nand UO_1976 (O_1976,N_14057,N_12608);
or UO_1977 (O_1977,N_10702,N_10555);
or UO_1978 (O_1978,N_14349,N_14231);
or UO_1979 (O_1979,N_11422,N_14700);
or UO_1980 (O_1980,N_12358,N_13599);
and UO_1981 (O_1981,N_14196,N_14038);
xnor UO_1982 (O_1982,N_10762,N_14075);
and UO_1983 (O_1983,N_11649,N_13246);
nand UO_1984 (O_1984,N_12156,N_14327);
nor UO_1985 (O_1985,N_14877,N_13902);
and UO_1986 (O_1986,N_14364,N_11936);
or UO_1987 (O_1987,N_14724,N_11570);
nand UO_1988 (O_1988,N_14607,N_12005);
and UO_1989 (O_1989,N_13724,N_13389);
nand UO_1990 (O_1990,N_10059,N_13711);
xnor UO_1991 (O_1991,N_14583,N_14186);
nand UO_1992 (O_1992,N_11325,N_11160);
and UO_1993 (O_1993,N_10504,N_10334);
and UO_1994 (O_1994,N_12748,N_14619);
xnor UO_1995 (O_1995,N_11810,N_14982);
or UO_1996 (O_1996,N_10790,N_10200);
nand UO_1997 (O_1997,N_10889,N_11418);
nand UO_1998 (O_1998,N_14124,N_11826);
or UO_1999 (O_1999,N_10978,N_11594);
endmodule