module basic_2000_20000_2500_10_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_364,In_1750);
nor U1 (N_1,In_187,In_70);
and U2 (N_2,In_146,In_260);
and U3 (N_3,In_29,In_729);
xor U4 (N_4,In_870,In_971);
or U5 (N_5,In_1659,In_1730);
nor U6 (N_6,In_1339,In_1764);
or U7 (N_7,In_899,In_1180);
nand U8 (N_8,In_351,In_1547);
or U9 (N_9,In_393,In_1661);
nor U10 (N_10,In_341,In_1169);
nand U11 (N_11,In_771,In_409);
and U12 (N_12,In_345,In_669);
nor U13 (N_13,In_957,In_1944);
and U14 (N_14,In_1154,In_1240);
nor U15 (N_15,In_1089,In_732);
or U16 (N_16,In_1631,In_907);
nor U17 (N_17,In_542,In_1355);
or U18 (N_18,In_21,In_1682);
nor U19 (N_19,In_1598,In_1261);
and U20 (N_20,In_1504,In_1928);
or U21 (N_21,In_1331,In_1566);
nor U22 (N_22,In_338,In_989);
and U23 (N_23,In_1193,In_607);
xor U24 (N_24,In_1787,In_630);
or U25 (N_25,In_388,In_103);
and U26 (N_26,In_1250,In_502);
or U27 (N_27,In_1910,In_31);
and U28 (N_28,In_1699,In_1013);
nor U29 (N_29,In_1755,In_482);
nor U30 (N_30,In_144,In_628);
nand U31 (N_31,In_603,In_406);
xor U32 (N_32,In_1371,In_1087);
nor U33 (N_33,In_979,In_1924);
or U34 (N_34,In_1433,In_1541);
nand U35 (N_35,In_209,In_1604);
and U36 (N_36,In_1496,In_1858);
nor U37 (N_37,In_613,In_269);
or U38 (N_38,In_663,In_1563);
nor U39 (N_39,In_1579,In_253);
nand U40 (N_40,In_777,In_798);
xor U41 (N_41,In_235,In_1783);
nor U42 (N_42,In_840,In_1343);
xnor U43 (N_43,In_1701,In_498);
or U44 (N_44,In_635,In_709);
and U45 (N_45,In_195,In_1643);
and U46 (N_46,In_1825,In_1779);
nand U47 (N_47,In_311,In_951);
or U48 (N_48,In_176,In_1322);
or U49 (N_49,In_475,In_541);
nor U50 (N_50,In_1795,In_124);
and U51 (N_51,In_1065,In_1959);
or U52 (N_52,In_1006,In_740);
or U53 (N_53,In_1975,In_1562);
and U54 (N_54,In_632,In_373);
nor U55 (N_55,In_858,In_787);
xnor U56 (N_56,In_1703,In_446);
or U57 (N_57,In_1761,In_1657);
nand U58 (N_58,In_212,In_955);
nand U59 (N_59,In_539,In_401);
and U60 (N_60,In_282,In_1204);
or U61 (N_61,In_836,In_1766);
nand U62 (N_62,In_1920,In_433);
nand U63 (N_63,In_492,In_1800);
and U64 (N_64,In_1252,In_1791);
nand U65 (N_65,In_272,In_1763);
nand U66 (N_66,In_1680,In_647);
or U67 (N_67,In_1488,In_274);
nand U68 (N_68,In_166,In_268);
xnor U69 (N_69,In_1070,In_667);
nor U70 (N_70,In_1068,In_1345);
nand U71 (N_71,In_1536,In_273);
nor U72 (N_72,In_127,In_1583);
nor U73 (N_73,In_1190,In_1447);
or U74 (N_74,In_1798,In_646);
nor U75 (N_75,In_1184,In_668);
nand U76 (N_76,In_1437,In_1436);
nor U77 (N_77,In_1905,In_1704);
and U78 (N_78,In_1530,In_1112);
nor U79 (N_79,In_566,In_784);
and U80 (N_80,In_164,In_1677);
nand U81 (N_81,In_1269,In_815);
or U82 (N_82,In_1615,In_1251);
nor U83 (N_83,In_1129,In_883);
nand U84 (N_84,In_535,In_399);
or U85 (N_85,In_1757,In_417);
and U86 (N_86,In_1027,In_1652);
xor U87 (N_87,In_639,In_1569);
nor U88 (N_88,In_442,In_84);
and U89 (N_89,In_1827,In_1502);
nor U90 (N_90,In_1167,In_491);
or U91 (N_91,In_1182,In_244);
xor U92 (N_92,In_745,In_710);
nand U93 (N_93,In_1904,In_1685);
and U94 (N_94,In_1772,In_1441);
or U95 (N_95,In_69,In_389);
nand U96 (N_96,In_604,In_114);
and U97 (N_97,In_1919,In_1257);
xnor U98 (N_98,In_1951,In_856);
nor U99 (N_99,In_1277,In_137);
nand U100 (N_100,In_138,In_369);
nor U101 (N_101,In_1650,In_919);
or U102 (N_102,In_233,In_1140);
xnor U103 (N_103,In_1762,In_653);
nand U104 (N_104,In_289,In_596);
xor U105 (N_105,In_862,In_1354);
nand U106 (N_106,In_429,In_1238);
nand U107 (N_107,In_316,In_1745);
and U108 (N_108,In_1995,In_1585);
and U109 (N_109,In_1312,In_967);
nand U110 (N_110,In_193,In_1983);
nand U111 (N_111,In_1881,In_786);
and U112 (N_112,In_579,In_1876);
and U113 (N_113,In_860,In_1014);
and U114 (N_114,In_1743,In_1908);
nand U115 (N_115,In_718,In_1584);
nor U116 (N_116,In_5,In_252);
xor U117 (N_117,In_1094,In_1195);
and U118 (N_118,In_331,In_525);
nor U119 (N_119,In_1775,In_863);
nand U120 (N_120,In_1512,In_360);
nand U121 (N_121,In_271,In_1438);
nand U122 (N_122,In_1095,In_327);
nor U123 (N_123,In_145,In_404);
nand U124 (N_124,In_1047,In_1340);
or U125 (N_125,In_128,In_436);
nor U126 (N_126,In_1851,In_1024);
nand U127 (N_127,In_255,In_972);
and U128 (N_128,In_1491,In_1913);
or U129 (N_129,In_730,In_765);
and U130 (N_130,In_864,In_332);
or U131 (N_131,In_996,In_1336);
and U132 (N_132,In_1966,In_109);
xnor U133 (N_133,In_157,In_1712);
nand U134 (N_134,In_1374,In_276);
nand U135 (N_135,In_300,In_407);
nand U136 (N_136,In_82,In_270);
and U137 (N_137,In_1329,In_1553);
or U138 (N_138,In_1846,In_558);
and U139 (N_139,In_1753,In_651);
nor U140 (N_140,In_554,In_66);
nor U141 (N_141,In_1593,In_1559);
nor U142 (N_142,In_1282,In_1150);
or U143 (N_143,In_658,In_938);
nand U144 (N_144,In_733,In_825);
nor U145 (N_145,In_241,In_1359);
and U146 (N_146,In_1366,In_568);
and U147 (N_147,In_310,In_104);
nand U148 (N_148,In_1192,In_690);
nand U149 (N_149,In_246,In_1028);
xor U150 (N_150,In_843,In_1335);
nor U151 (N_151,In_1653,In_358);
nor U152 (N_152,In_918,In_547);
or U153 (N_153,In_692,In_1323);
nand U154 (N_154,In_588,In_481);
or U155 (N_155,In_655,In_159);
or U156 (N_156,In_721,In_16);
and U157 (N_157,In_529,In_1747);
or U158 (N_158,In_1855,In_1369);
nor U159 (N_159,In_1955,In_224);
nand U160 (N_160,In_1754,In_256);
and U161 (N_161,In_820,In_1759);
nor U162 (N_162,In_1271,In_984);
and U163 (N_163,In_28,In_1370);
nor U164 (N_164,In_93,In_1690);
or U165 (N_165,In_1254,In_396);
or U166 (N_166,In_203,In_323);
or U167 (N_167,In_249,In_1183);
or U168 (N_168,In_886,In_226);
or U169 (N_169,In_275,In_416);
or U170 (N_170,In_102,In_73);
nor U171 (N_171,In_656,In_1038);
nand U172 (N_172,In_123,In_940);
and U173 (N_173,In_823,In_1816);
or U174 (N_174,In_501,In_1565);
nor U175 (N_175,In_1410,In_1988);
nand U176 (N_176,In_1466,In_1211);
or U177 (N_177,In_917,In_774);
or U178 (N_178,In_457,In_1057);
nand U179 (N_179,In_594,In_1400);
nand U180 (N_180,In_1009,In_438);
or U181 (N_181,In_695,In_679);
xnor U182 (N_182,In_706,In_1073);
xor U183 (N_183,In_1160,In_291);
nand U184 (N_184,In_169,In_536);
and U185 (N_185,In_998,In_1575);
nor U186 (N_186,In_591,In_1805);
and U187 (N_187,In_200,In_910);
or U188 (N_188,In_1932,In_43);
and U189 (N_189,In_976,In_1732);
or U190 (N_190,In_1147,In_464);
nand U191 (N_191,In_1877,In_1421);
and U192 (N_192,In_804,In_1999);
xnor U193 (N_193,In_1091,In_1689);
xor U194 (N_194,In_990,In_1337);
or U195 (N_195,In_451,In_1463);
or U196 (N_196,In_179,In_1676);
or U197 (N_197,In_1596,In_754);
nand U198 (N_198,In_1085,In_26);
nor U199 (N_199,In_722,In_1746);
nand U200 (N_200,In_35,In_810);
or U201 (N_201,In_1821,In_229);
xnor U202 (N_202,In_361,In_473);
or U203 (N_203,In_1231,In_736);
and U204 (N_204,In_1061,In_1933);
or U205 (N_205,In_1036,In_428);
and U206 (N_206,In_459,In_521);
and U207 (N_207,In_325,In_315);
nor U208 (N_208,In_785,In_1208);
xor U209 (N_209,In_419,In_211);
nor U210 (N_210,In_780,In_202);
nor U211 (N_211,In_773,In_1266);
nor U212 (N_212,In_1744,In_538);
xnor U213 (N_213,In_614,In_439);
nand U214 (N_214,In_374,In_354);
and U215 (N_215,In_552,In_250);
and U216 (N_216,In_995,In_519);
nor U217 (N_217,In_1247,In_1874);
nand U218 (N_218,In_293,In_1947);
nor U219 (N_219,In_1413,In_1997);
nand U220 (N_220,In_1614,In_624);
or U221 (N_221,In_1201,In_1316);
and U222 (N_222,In_139,In_468);
nor U223 (N_223,In_671,In_363);
and U224 (N_224,In_441,In_247);
nor U225 (N_225,In_477,In_1213);
nor U226 (N_226,In_133,In_503);
nor U227 (N_227,In_1996,In_239);
and U228 (N_228,In_608,In_85);
and U229 (N_229,In_1242,In_1613);
xor U230 (N_230,In_376,In_1888);
xnor U231 (N_231,In_1313,In_56);
xor U232 (N_232,In_71,In_683);
or U233 (N_233,In_1450,In_1555);
and U234 (N_234,In_79,In_1931);
and U235 (N_235,In_1993,In_1644);
nand U236 (N_236,In_1782,In_1051);
and U237 (N_237,In_197,In_1054);
nand U238 (N_238,In_1237,In_455);
nor U239 (N_239,In_1130,In_1395);
nand U240 (N_240,In_1601,In_1980);
xnor U241 (N_241,In_696,In_403);
and U242 (N_242,In_1307,In_476);
and U243 (N_243,In_267,In_1581);
nand U244 (N_244,In_643,In_1662);
or U245 (N_245,In_962,In_472);
nand U246 (N_246,In_769,In_1222);
nor U247 (N_247,In_278,In_1673);
and U248 (N_248,In_923,In_914);
and U249 (N_249,In_116,In_466);
or U250 (N_250,In_346,In_674);
nor U251 (N_251,In_1351,In_112);
nand U252 (N_252,In_1207,In_1382);
or U253 (N_253,In_1953,In_644);
or U254 (N_254,In_1327,In_324);
and U255 (N_255,In_999,In_573);
xor U256 (N_256,In_1125,In_1170);
nor U257 (N_257,In_1573,In_704);
nand U258 (N_258,In_1317,In_198);
nand U259 (N_259,In_891,In_1696);
or U260 (N_260,In_958,In_420);
or U261 (N_261,In_609,In_953);
nand U262 (N_262,In_288,In_821);
and U263 (N_263,In_661,In_792);
and U264 (N_264,In_117,In_1640);
nor U265 (N_265,In_1939,In_1560);
nand U266 (N_266,In_33,In_1958);
xnor U267 (N_267,In_1116,In_1950);
or U268 (N_268,In_1608,In_140);
nor U269 (N_269,In_708,In_1751);
xor U270 (N_270,In_1633,In_634);
nor U271 (N_271,In_337,In_126);
xor U272 (N_272,In_177,In_1298);
nor U273 (N_273,In_1586,In_1927);
nand U274 (N_274,In_1771,In_1490);
xor U275 (N_275,In_368,In_218);
nor U276 (N_276,In_878,In_616);
or U277 (N_277,In_150,In_1119);
or U278 (N_278,In_1037,In_1287);
xor U279 (N_279,In_42,In_1268);
or U280 (N_280,In_1408,In_1402);
and U281 (N_281,In_1989,In_813);
and U282 (N_282,In_1778,In_734);
or U283 (N_283,In_453,In_892);
nor U284 (N_284,In_788,In_968);
and U285 (N_285,In_1153,In_367);
xor U286 (N_286,In_731,In_1445);
nand U287 (N_287,In_548,In_687);
or U288 (N_288,In_1734,In_1862);
and U289 (N_289,In_728,In_752);
and U290 (N_290,In_1609,In_15);
nand U291 (N_291,In_1288,In_1161);
and U292 (N_292,In_835,In_1715);
xnor U293 (N_293,In_130,In_509);
or U294 (N_294,In_672,In_1081);
and U295 (N_295,In_714,In_1998);
and U296 (N_296,In_1765,In_1926);
or U297 (N_297,In_174,In_1055);
nand U298 (N_298,In_1668,In_832);
or U299 (N_299,In_1796,In_1446);
nor U300 (N_300,In_873,In_1832);
xnor U301 (N_301,In_1811,In_1069);
and U302 (N_302,In_1058,In_750);
xor U303 (N_303,In_599,In_1056);
and U304 (N_304,In_1907,In_797);
nand U305 (N_305,In_208,In_1776);
nand U306 (N_306,In_38,In_675);
nand U307 (N_307,In_1272,In_1099);
and U308 (N_308,In_1620,In_362);
or U309 (N_309,In_762,In_355);
nand U310 (N_310,In_901,In_977);
and U311 (N_311,In_47,In_1648);
nand U312 (N_312,In_410,In_595);
or U313 (N_313,In_513,In_62);
or U314 (N_314,In_1605,In_524);
and U315 (N_315,In_236,In_850);
nor U316 (N_316,In_1546,In_186);
xnor U317 (N_317,In_950,In_631);
or U318 (N_318,In_215,In_505);
xor U319 (N_319,In_1393,In_885);
nand U320 (N_320,In_1276,In_626);
xnor U321 (N_321,In_1321,In_107);
or U322 (N_322,In_1965,In_1517);
nor U323 (N_323,In_192,In_1669);
xor U324 (N_324,In_1487,In_40);
or U325 (N_325,In_1831,In_1381);
nand U326 (N_326,In_1857,In_9);
xor U327 (N_327,In_924,In_100);
nor U328 (N_328,In_751,In_490);
xor U329 (N_329,In_340,In_1101);
nor U330 (N_330,In_1618,In_1571);
nand U331 (N_331,In_1286,In_911);
or U332 (N_332,In_592,In_279);
nand U333 (N_333,In_1952,In_386);
or U334 (N_334,In_1649,In_1155);
nand U335 (N_335,In_549,In_1628);
and U336 (N_336,In_1885,In_1552);
and U337 (N_337,In_1902,In_942);
nand U338 (N_338,In_1108,In_1976);
xor U339 (N_339,In_292,In_574);
or U340 (N_340,In_859,In_1082);
nand U341 (N_341,In_531,In_1471);
nor U342 (N_342,In_1538,In_67);
and U343 (N_343,In_75,In_1945);
nor U344 (N_344,In_263,In_1588);
or U345 (N_345,In_147,In_1300);
and U346 (N_346,In_158,In_1306);
nand U347 (N_347,In_965,In_1172);
nor U348 (N_348,In_1105,In_1171);
nor U349 (N_349,In_309,In_1672);
nor U350 (N_350,In_760,In_1258);
and U351 (N_351,In_1205,In_1405);
or U352 (N_352,In_526,In_484);
nand U353 (N_353,In_1419,In_1320);
and U354 (N_354,In_1333,In_1698);
and U355 (N_355,In_55,In_707);
nor U356 (N_356,In_90,In_474);
nand U357 (N_357,In_1539,In_3);
or U358 (N_358,In_72,In_937);
or U359 (N_359,In_1295,In_1807);
nor U360 (N_360,In_1363,In_1664);
or U361 (N_361,In_1216,In_83);
or U362 (N_362,In_1972,In_1367);
or U363 (N_363,In_1311,In_576);
or U364 (N_364,In_1706,In_589);
nand U365 (N_365,In_1387,In_1558);
or U366 (N_366,In_1721,In_1049);
and U367 (N_367,In_68,In_456);
nor U368 (N_368,In_743,In_1098);
and U369 (N_369,In_1021,In_532);
nand U370 (N_370,In_1568,In_802);
and U371 (N_371,In_264,In_1551);
and U372 (N_372,In_540,In_1937);
nor U373 (N_373,In_737,In_1378);
nor U374 (N_374,In_1325,In_666);
nand U375 (N_375,In_1886,In_1232);
nor U376 (N_376,In_143,In_1077);
or U377 (N_377,In_1603,In_1619);
nor U378 (N_378,In_500,In_1448);
nand U379 (N_379,In_1981,In_570);
or U380 (N_380,In_370,In_487);
nor U381 (N_381,In_30,In_617);
and U382 (N_382,In_32,In_1867);
or U383 (N_383,In_849,In_826);
xor U384 (N_384,In_1016,In_1506);
nor U385 (N_385,In_1425,In_232);
nor U386 (N_386,In_347,In_959);
and U387 (N_387,In_1520,In_908);
nor U388 (N_388,In_1309,In_1899);
and U389 (N_389,In_793,In_508);
and U390 (N_390,In_152,In_1864);
nand U391 (N_391,In_930,In_1814);
xor U392 (N_392,In_1849,In_583);
nor U393 (N_393,In_1592,In_183);
xor U394 (N_394,In_1641,In_806);
nor U395 (N_395,In_344,In_611);
nand U396 (N_396,In_58,In_1194);
nand U397 (N_397,In_1026,In_196);
xnor U398 (N_398,In_1632,In_783);
nor U399 (N_399,In_1522,In_1892);
nor U400 (N_400,In_1768,In_681);
xor U401 (N_401,In_1597,In_1627);
nand U402 (N_402,In_36,In_853);
nand U403 (N_403,In_1422,In_1518);
or U404 (N_404,In_1264,In_1233);
nor U405 (N_405,In_125,In_562);
or U406 (N_406,In_206,In_1812);
or U407 (N_407,In_1076,In_987);
nand U408 (N_408,In_1602,In_1185);
nor U409 (N_409,In_17,In_258);
and U410 (N_410,In_881,In_1557);
and U411 (N_411,In_1200,In_605);
nor U412 (N_412,In_1535,In_1725);
or U413 (N_413,In_449,In_96);
nor U414 (N_414,In_497,In_1912);
nand U415 (N_415,In_227,In_1681);
nand U416 (N_416,In_287,In_1564);
or U417 (N_417,In_982,In_1044);
nor U418 (N_418,In_814,In_1587);
and U419 (N_419,In_1079,In_1839);
or U420 (N_420,In_54,In_1152);
nand U421 (N_421,In_712,In_1590);
xnor U422 (N_422,In_1860,In_1507);
or U423 (N_423,In_80,In_1790);
nor U424 (N_424,In_1523,In_550);
and U425 (N_425,In_1513,In_572);
and U426 (N_426,In_865,In_398);
nor U427 (N_427,In_89,In_824);
xnor U428 (N_428,In_1942,In_766);
or U429 (N_429,In_1921,In_571);
nand U430 (N_430,In_87,In_606);
xnor U431 (N_431,In_518,In_228);
and U432 (N_432,In_929,In_900);
xor U433 (N_433,In_1900,In_1741);
and U434 (N_434,In_1255,In_1235);
and U435 (N_435,In_1015,In_1391);
nor U436 (N_436,In_776,In_855);
or U437 (N_437,In_1075,In_779);
and U438 (N_438,In_1412,In_348);
and U439 (N_439,In_171,In_1948);
and U440 (N_440,In_460,In_190);
nor U441 (N_441,In_876,In_251);
nand U442 (N_442,In_304,In_1072);
nand U443 (N_443,In_1263,In_49);
and U444 (N_444,In_567,In_470);
or U445 (N_445,In_758,In_371);
nor U446 (N_446,In_1901,In_1737);
nor U447 (N_447,In_742,In_1176);
and U448 (N_448,In_405,In_1820);
nor U449 (N_449,In_20,In_1570);
or U450 (N_450,In_1642,In_778);
nor U451 (N_451,In_1303,In_580);
or U452 (N_452,In_1967,In_1146);
or U453 (N_453,In_698,In_727);
nand U454 (N_454,In_19,In_1088);
and U455 (N_455,In_1890,In_1464);
nor U456 (N_456,In_703,In_1420);
nor U457 (N_457,In_1383,In_925);
nand U458 (N_458,In_110,In_642);
nand U459 (N_459,In_1482,In_1489);
nor U460 (N_460,In_1178,In_1660);
nand U461 (N_461,In_447,In_1457);
xor U462 (N_462,In_1930,In_1707);
and U463 (N_463,In_985,In_160);
nor U464 (N_464,In_1236,In_1990);
nor U465 (N_465,In_1050,In_1543);
nor U466 (N_466,In_1035,In_319);
or U467 (N_467,In_1493,In_1223);
and U468 (N_468,In_1005,In_1275);
xnor U469 (N_469,In_590,In_118);
or U470 (N_470,In_240,In_1357);
and U471 (N_471,In_132,In_328);
or U472 (N_472,In_1722,In_1866);
and U473 (N_473,In_504,In_191);
and U474 (N_474,In_619,In_1802);
or U475 (N_475,In_1758,In_946);
xnor U476 (N_476,In_1629,In_1709);
nor U477 (N_477,In_903,In_640);
nand U478 (N_478,In_544,In_889);
nor U479 (N_479,In_1964,In_1658);
or U480 (N_480,In_1034,In_378);
nand U481 (N_481,In_167,In_739);
xor U482 (N_482,In_1022,In_1462);
nor U483 (N_483,In_469,In_77);
or U484 (N_484,In_194,In_63);
or U485 (N_485,In_1360,In_652);
nand U486 (N_486,In_1828,In_1484);
xor U487 (N_487,In_1880,In_1683);
nand U488 (N_488,In_847,In_654);
or U489 (N_489,In_623,In_1826);
nand U490 (N_490,In_561,In_365);
or U491 (N_491,In_317,In_1505);
or U492 (N_492,In_1872,In_1040);
or U493 (N_493,In_392,In_1289);
and U494 (N_494,In_506,In_385);
nand U495 (N_495,In_1469,In_720);
or U496 (N_496,In_676,In_34);
and U497 (N_497,In_6,In_559);
or U498 (N_498,In_1884,In_1384);
nand U499 (N_499,In_1020,In_1137);
and U500 (N_500,In_136,In_1793);
or U501 (N_501,In_1453,In_99);
and U502 (N_502,In_877,In_1667);
or U503 (N_503,In_135,In_1638);
and U504 (N_504,In_1000,In_711);
and U505 (N_505,In_1949,In_902);
nor U506 (N_506,In_528,In_1149);
nand U507 (N_507,In_11,In_1624);
nor U508 (N_508,In_1914,In_1856);
xnor U509 (N_509,In_1198,In_153);
or U510 (N_510,In_1274,In_1063);
xor U511 (N_511,In_237,In_1011);
or U512 (N_512,In_1865,In_1824);
nand U513 (N_513,In_1124,In_584);
and U514 (N_514,In_717,In_1819);
and U515 (N_515,In_1285,In_1941);
or U516 (N_516,In_1465,In_1111);
nor U517 (N_517,In_1896,In_600);
and U518 (N_518,In_1002,In_575);
nor U519 (N_519,In_1053,In_872);
nand U520 (N_520,In_1519,In_1957);
and U521 (N_521,In_867,In_101);
and U522 (N_522,In_1230,In_516);
and U523 (N_523,In_95,In_1328);
nand U524 (N_524,In_1460,In_818);
nand U525 (N_525,In_1726,In_450);
or U526 (N_526,In_799,In_1647);
xnor U527 (N_527,In_1705,In_1637);
nand U528 (N_528,In_380,In_201);
xnor U529 (N_529,In_1168,In_1666);
and U530 (N_530,In_1397,In_356);
nand U531 (N_531,In_665,In_1870);
nand U532 (N_532,In_1822,In_1356);
nand U533 (N_533,In_199,In_339);
xor U534 (N_534,In_1086,In_1808);
xnor U535 (N_535,In_909,In_884);
or U536 (N_536,In_983,In_391);
and U537 (N_537,In_725,In_522);
or U538 (N_538,In_284,In_357);
or U539 (N_539,In_992,In_105);
xor U540 (N_540,In_1375,In_1334);
nand U541 (N_541,In_808,In_1749);
and U542 (N_542,In_1991,In_1938);
or U543 (N_543,In_945,In_747);
and U544 (N_544,In_45,In_812);
nand U545 (N_545,In_1476,In_1191);
or U546 (N_546,In_1612,In_222);
nand U547 (N_547,In_1777,In_155);
nor U548 (N_548,In_1107,In_4);
nor U549 (N_549,In_156,In_1424);
nor U550 (N_550,In_1362,In_1809);
nand U551 (N_551,In_699,In_845);
nand U552 (N_552,In_1936,In_1818);
nor U553 (N_553,In_1377,In_182);
and U554 (N_554,In_980,In_1968);
xor U555 (N_555,In_1361,In_308);
or U556 (N_556,In_1971,In_1164);
or U557 (N_557,In_1318,In_746);
nand U558 (N_558,In_1467,In_1946);
nor U559 (N_559,In_234,In_1248);
and U560 (N_560,In_933,In_1202);
nor U561 (N_561,In_726,In_1655);
xnor U562 (N_562,In_963,In_1157);
nor U563 (N_563,In_1935,In_1803);
nor U564 (N_564,In_724,In_1891);
nor U565 (N_565,In_1241,In_1773);
nor U566 (N_566,In_893,In_1332);
nand U567 (N_567,In_1675,In_306);
or U568 (N_568,In_796,In_1203);
or U569 (N_569,In_1041,In_91);
and U570 (N_570,In_1854,In_1815);
nand U571 (N_571,In_991,In_926);
nand U572 (N_572,In_204,In_931);
nand U573 (N_573,In_1262,In_569);
nand U574 (N_574,In_296,In_1209);
nor U575 (N_575,In_648,In_1120);
nor U576 (N_576,In_1626,In_221);
nor U577 (N_577,In_1893,In_1141);
or U578 (N_578,In_149,In_1092);
or U579 (N_579,In_1429,In_948);
nand U580 (N_580,In_621,In_1500);
nand U581 (N_581,In_59,In_1019);
or U582 (N_582,In_895,In_1830);
or U583 (N_583,In_1962,In_1394);
nand U584 (N_584,In_22,In_817);
and U585 (N_585,In_161,In_1407);
and U586 (N_586,In_1206,In_178);
nor U587 (N_587,In_693,In_350);
nor U588 (N_588,In_1510,In_1969);
nand U589 (N_589,In_1442,In_680);
or U590 (N_590,In_662,In_320);
nor U591 (N_591,In_1845,In_1740);
xnor U592 (N_592,In_94,In_912);
or U593 (N_593,In_1062,In_390);
xnor U594 (N_594,In_1310,In_641);
or U595 (N_595,In_894,In_842);
nor U596 (N_596,In_981,In_488);
or U597 (N_597,In_330,In_837);
and U598 (N_598,In_51,In_1423);
nand U599 (N_599,In_978,In_1521);
and U600 (N_600,In_1220,In_1984);
or U601 (N_601,In_1594,In_1097);
and U602 (N_602,In_1978,In_381);
and U603 (N_603,In_545,In_1227);
nand U604 (N_604,In_1396,In_1260);
nand U605 (N_605,In_297,In_1498);
nand U606 (N_606,In_587,In_1674);
nand U607 (N_607,In_1110,In_807);
nor U608 (N_608,In_1444,In_1443);
and U609 (N_609,In_431,In_1279);
nor U610 (N_610,In_1545,In_412);
and U611 (N_611,In_52,In_1039);
and U612 (N_612,In_1576,In_463);
nand U613 (N_613,In_1416,In_715);
and U614 (N_614,In_819,In_88);
nor U615 (N_615,In_830,In_1102);
nor U616 (N_616,In_1977,In_716);
and U617 (N_617,In_1308,In_44);
nor U618 (N_618,In_353,In_1799);
nand U619 (N_619,In_329,In_1302);
nand U620 (N_620,In_723,In_1385);
and U621 (N_621,In_86,In_1256);
or U622 (N_622,In_1610,In_839);
and U623 (N_623,In_1837,In_141);
nor U624 (N_624,In_283,In_254);
or U625 (N_625,In_960,In_1398);
and U626 (N_626,In_949,In_1229);
or U627 (N_627,In_586,In_921);
or U628 (N_628,In_53,In_515);
nand U629 (N_629,In_719,In_7);
or U630 (N_630,In_1373,In_1494);
and U631 (N_631,In_1386,In_479);
nor U632 (N_632,In_866,In_593);
nor U633 (N_633,In_1365,In_1481);
nand U634 (N_634,In_633,In_1514);
or U635 (N_635,In_759,In_887);
nor U636 (N_636,In_1244,In_60);
nand U637 (N_637,In_375,In_1911);
or U638 (N_638,In_1974,In_1228);
nor U639 (N_639,In_1118,In_947);
nand U640 (N_640,In_1456,In_1848);
or U641 (N_641,In_512,In_294);
and U642 (N_642,In_1894,In_1249);
or U643 (N_643,In_1616,In_1117);
nor U644 (N_644,In_1731,In_1639);
or U645 (N_645,In_851,In_700);
nor U646 (N_646,In_1449,In_424);
and U647 (N_647,In_1315,In_964);
and U648 (N_648,In_13,In_414);
xor U649 (N_649,In_1898,In_1869);
and U650 (N_650,In_1780,In_0);
or U651 (N_651,In_1029,In_1435);
xnor U652 (N_652,In_649,In_1007);
and U653 (N_653,In_1970,In_1526);
and U654 (N_654,In_1694,In_1136);
or U655 (N_655,In_514,In_1833);
or U656 (N_656,In_841,In_1003);
and U657 (N_657,In_1217,In_905);
nand U658 (N_658,In_1868,In_1817);
nand U659 (N_659,In_1199,In_1297);
and U660 (N_660,In_1064,In_831);
nor U661 (N_661,In_744,In_265);
or U662 (N_662,In_1292,In_245);
nor U663 (N_663,In_520,In_1985);
nand U664 (N_664,In_811,In_1426);
and U665 (N_665,In_1084,In_1372);
nand U666 (N_666,In_1414,In_1524);
and U667 (N_667,In_1621,In_1688);
nor U668 (N_668,In_1270,In_952);
and U669 (N_669,In_1752,In_1503);
and U670 (N_670,In_934,In_1925);
or U671 (N_671,In_1842,In_1693);
nor U672 (N_672,In_816,In_1368);
nor U673 (N_673,In_1700,In_1717);
or U674 (N_674,In_189,In_333);
nand U675 (N_675,In_702,In_465);
xnor U676 (N_676,In_684,In_1030);
or U677 (N_677,In_563,In_660);
nand U678 (N_678,In_307,In_1572);
and U679 (N_679,In_1234,In_1246);
or U680 (N_680,In_181,In_1678);
or U681 (N_681,In_184,In_629);
nand U682 (N_682,In_299,In_1364);
and U683 (N_683,In_1219,In_257);
and U684 (N_684,In_551,In_1046);
nor U685 (N_685,In_321,In_560);
nand U686 (N_686,In_1591,In_1114);
or U687 (N_687,In_185,In_64);
xor U688 (N_688,In_1411,In_678);
or U689 (N_689,In_1267,In_1113);
nand U690 (N_690,In_168,In_1540);
nand U691 (N_691,In_1353,In_523);
and U692 (N_692,In_1478,In_677);
nor U693 (N_693,In_427,In_163);
nand U694 (N_694,In_1781,In_285);
or U695 (N_695,In_352,In_1186);
nor U696 (N_696,In_303,In_343);
nand U697 (N_697,In_243,In_1187);
xnor U698 (N_698,In_205,In_1871);
and U699 (N_699,In_973,In_1728);
and U700 (N_700,In_598,In_767);
nand U701 (N_701,In_1801,In_1889);
or U702 (N_702,In_1556,In_1853);
nor U703 (N_703,In_1515,In_610);
or U704 (N_704,In_387,In_741);
or U705 (N_705,In_852,In_1511);
nor U706 (N_706,In_1278,In_738);
nand U707 (N_707,In_638,In_1346);
nand U708 (N_708,In_553,In_415);
and U709 (N_709,In_478,In_98);
and U710 (N_710,In_422,In_936);
nor U711 (N_711,In_565,In_897);
nand U712 (N_712,In_1427,In_1455);
or U713 (N_713,In_673,In_1284);
and U714 (N_714,In_1495,In_225);
or U715 (N_715,In_483,In_1440);
xnor U716 (N_716,In_78,In_939);
nand U717 (N_717,In_1516,In_430);
and U718 (N_718,In_1218,In_686);
xnor U719 (N_719,In_1106,In_115);
or U720 (N_720,In_685,In_755);
nor U721 (N_721,In_1797,In_1531);
nand U722 (N_722,In_1273,In_682);
or U723 (N_723,In_782,In_1986);
and U724 (N_724,In_1388,In_1143);
or U725 (N_725,In_691,In_537);
nor U726 (N_726,In_1646,In_688);
xor U727 (N_727,In_1083,In_615);
nand U728 (N_728,In_37,In_1174);
nand U729 (N_729,In_210,In_372);
or U730 (N_730,In_834,In_1929);
nor U731 (N_731,In_1786,In_1544);
nor U732 (N_732,In_1431,In_748);
and U733 (N_733,In_869,In_1221);
and U734 (N_734,In_1711,In_1917);
or U735 (N_735,In_434,In_1850);
or U736 (N_736,In_890,In_1473);
or U737 (N_737,In_1499,In_131);
nand U738 (N_738,In_1852,In_1829);
or U739 (N_739,In_1607,In_1923);
or U740 (N_740,In_1093,In_111);
nor U741 (N_741,In_1454,In_1043);
nand U742 (N_742,In_1134,In_875);
and U743 (N_743,In_749,In_546);
or U744 (N_744,In_46,In_1451);
and U745 (N_745,In_961,In_1080);
and U746 (N_746,In_1379,In_402);
nor U747 (N_747,In_1338,In_1165);
or U748 (N_748,In_1844,In_1600);
and U749 (N_749,In_1067,In_1380);
and U750 (N_750,In_868,In_1023);
xnor U751 (N_751,In_467,In_349);
nor U752 (N_752,In_366,In_507);
or U753 (N_753,In_1922,In_1159);
nor U754 (N_754,In_154,In_1794);
and U755 (N_755,In_1716,In_1554);
or U756 (N_756,In_1280,In_1342);
or U757 (N_757,In_906,In_879);
or U758 (N_758,In_1611,In_612);
and U759 (N_759,In_1479,In_1622);
nand U760 (N_760,In_543,In_262);
and U761 (N_761,In_1718,In_12);
nand U762 (N_762,In_493,In_1017);
nor U763 (N_763,In_993,In_1066);
and U764 (N_764,In_1774,In_1239);
or U765 (N_765,In_326,In_223);
nor U766 (N_766,In_1691,In_1580);
xnor U767 (N_767,In_1702,In_1813);
xnor U768 (N_768,In_1525,In_1529);
or U769 (N_769,In_106,In_511);
nor U770 (N_770,In_697,In_1033);
nor U771 (N_771,In_1166,In_1144);
and U772 (N_772,In_756,In_219);
or U773 (N_773,In_556,In_1785);
nand U774 (N_774,In_1403,In_1145);
nand U775 (N_775,In_170,In_1406);
nand U776 (N_776,In_379,In_828);
or U777 (N_777,In_448,In_1349);
nor U778 (N_778,In_1025,In_1756);
or U779 (N_779,In_1294,In_1534);
and U780 (N_780,In_1032,In_1769);
and U781 (N_781,In_555,In_791);
or U782 (N_782,In_1031,In_134);
and U783 (N_783,In_1840,In_932);
nand U784 (N_784,In_1909,In_1259);
nor U785 (N_785,In_1589,In_1686);
nor U786 (N_786,In_1392,In_1156);
nand U787 (N_787,In_670,In_801);
xor U788 (N_788,In_1104,In_1729);
and U789 (N_789,In_1126,In_650);
xnor U790 (N_790,In_975,In_27);
and U791 (N_791,In_1461,In_986);
nor U792 (N_792,In_1224,In_533);
and U793 (N_793,In_1501,In_180);
nand U794 (N_794,In_809,In_50);
nand U795 (N_795,In_1417,In_534);
and U796 (N_796,In_1723,In_829);
nor U797 (N_797,In_1151,In_1823);
nor U798 (N_798,In_1324,In_1253);
xor U799 (N_799,In_259,In_1430);
nand U800 (N_800,In_318,In_1173);
nor U801 (N_801,In_1100,In_1341);
nand U802 (N_802,In_622,In_1863);
or U803 (N_803,In_1916,In_1);
or U804 (N_804,In_997,In_597);
xnor U805 (N_805,In_1645,In_1226);
or U806 (N_806,In_384,In_527);
nor U807 (N_807,In_81,In_1788);
nand U808 (N_808,In_645,In_1188);
and U809 (N_809,In_1177,In_1138);
and U810 (N_810,In_1301,In_1135);
and U811 (N_811,In_838,In_454);
nand U812 (N_812,In_61,In_411);
or U813 (N_813,In_1651,In_122);
xnor U814 (N_814,In_10,In_1574);
or U815 (N_815,In_1548,In_775);
xnor U816 (N_816,In_1606,In_1181);
and U817 (N_817,In_1630,In_382);
nand U818 (N_818,In_1963,In_1389);
and U819 (N_819,In_1663,In_394);
xnor U820 (N_820,In_803,In_1838);
or U821 (N_821,In_1835,In_1671);
and U822 (N_822,In_1291,In_1142);
nor U823 (N_823,In_1595,In_1468);
or U824 (N_824,In_298,In_1128);
nand U825 (N_825,In_602,In_657);
or U826 (N_826,In_113,In_1918);
xnor U827 (N_827,In_313,In_1804);
nand U828 (N_828,In_314,In_213);
or U829 (N_829,In_1859,In_1714);
or U830 (N_830,In_1415,In_1670);
and U831 (N_831,In_1048,In_1376);
and U832 (N_832,In_1319,In_1961);
nand U833 (N_833,In_359,In_1314);
nand U834 (N_834,In_800,In_8);
or U835 (N_835,In_1458,In_1293);
nor U836 (N_836,In_1096,In_1122);
xor U837 (N_837,In_231,In_1687);
nor U838 (N_838,In_969,In_794);
nor U839 (N_839,In_1008,In_1873);
nand U840 (N_840,In_1738,In_1724);
and U841 (N_841,In_956,In_1483);
nor U842 (N_842,In_772,In_1982);
xnor U843 (N_843,In_1018,In_1748);
nand U844 (N_844,In_1225,In_395);
nand U845 (N_845,In_1189,In_882);
nor U846 (N_846,In_1492,In_1549);
nand U847 (N_847,In_1399,In_1452);
nand U848 (N_848,In_335,In_861);
nor U849 (N_849,In_301,In_768);
nor U850 (N_850,In_577,In_601);
nor U851 (N_851,In_1550,In_1304);
nand U852 (N_852,In_238,In_915);
nor U853 (N_853,In_1480,In_789);
and U854 (N_854,In_822,In_1409);
and U855 (N_855,In_1879,In_1994);
and U856 (N_856,In_1906,In_874);
nor U857 (N_857,In_627,In_286);
nor U858 (N_858,In_1895,In_1861);
nand U859 (N_859,In_142,In_480);
nor U860 (N_860,In_1634,In_1470);
or U861 (N_861,In_1834,In_1789);
and U862 (N_862,In_927,In_1132);
and U863 (N_863,In_994,In_129);
and U864 (N_864,In_1915,In_1806);
xor U865 (N_865,In_471,In_486);
and U866 (N_866,In_280,In_1767);
or U867 (N_867,In_495,In_735);
or U868 (N_868,In_928,In_581);
and U869 (N_869,In_1735,In_342);
and U870 (N_870,In_1887,In_248);
or U871 (N_871,In_1527,In_165);
or U872 (N_872,In_1577,In_935);
or U873 (N_873,In_944,In_1497);
xnor U874 (N_874,In_637,In_1348);
nor U875 (N_875,In_857,In_753);
and U876 (N_876,In_1784,In_1350);
xnor U877 (N_877,In_48,In_757);
or U878 (N_878,In_1708,In_1695);
or U879 (N_879,In_1934,In_1617);
and U880 (N_880,In_220,In_844);
or U881 (N_881,In_1528,In_1943);
or U882 (N_882,In_1636,In_620);
xnor U883 (N_883,In_120,In_1836);
nand U884 (N_884,In_790,In_1158);
nand U885 (N_885,In_175,In_1567);
or U886 (N_886,In_1401,In_443);
or U887 (N_887,In_1109,In_1352);
nor U888 (N_888,In_1770,In_1296);
or U889 (N_889,In_1212,In_920);
and U890 (N_890,In_494,In_425);
nand U891 (N_891,In_1508,In_489);
nand U892 (N_892,In_188,In_625);
xor U893 (N_893,In_1001,In_1542);
nand U894 (N_894,In_896,In_1509);
and U895 (N_895,In_1979,In_1210);
nand U896 (N_896,In_1697,In_261);
xor U897 (N_897,In_1472,In_913);
nor U898 (N_898,In_1432,In_1665);
nor U899 (N_899,In_41,In_437);
xor U900 (N_900,In_1903,In_1474);
nor U901 (N_901,In_713,In_1635);
or U902 (N_902,In_1710,In_1090);
and U903 (N_903,In_65,In_1692);
nand U904 (N_904,In_1163,In_1344);
xnor U905 (N_905,In_1954,In_1305);
or U906 (N_906,In_423,In_2);
nand U907 (N_907,In_1713,In_970);
and U908 (N_908,In_659,In_954);
nand U909 (N_909,In_1742,In_1103);
or U910 (N_910,In_1486,In_281);
xor U911 (N_911,In_1162,In_916);
nand U912 (N_912,In_1599,In_485);
nand U913 (N_913,In_458,In_1960);
and U914 (N_914,In_1197,In_1847);
and U915 (N_915,In_295,In_833);
or U916 (N_916,In_705,In_805);
nand U917 (N_917,In_1404,In_24);
nand U918 (N_918,In_418,In_1115);
and U919 (N_919,In_108,In_496);
nand U920 (N_920,In_898,In_57);
xnor U921 (N_921,In_880,In_1578);
nor U922 (N_922,In_1878,In_582);
nand U923 (N_923,In_305,In_462);
or U924 (N_924,In_1760,In_1299);
or U925 (N_925,In_1656,In_312);
nor U926 (N_926,In_1330,In_1720);
nand U927 (N_927,In_148,In_207);
nor U928 (N_928,In_557,In_1428);
nand U929 (N_929,In_413,In_1148);
xor U930 (N_930,In_1987,In_426);
nor U931 (N_931,In_694,In_1175);
nor U932 (N_932,In_1883,In_1733);
nor U933 (N_933,In_230,In_988);
and U934 (N_934,In_217,In_1139);
and U935 (N_935,In_1475,In_290);
nor U936 (N_936,In_1736,In_1123);
nand U937 (N_937,In_827,In_1347);
or U938 (N_938,In_1727,In_452);
and U939 (N_939,In_1477,In_266);
or U940 (N_940,In_764,In_517);
or U941 (N_941,In_1561,In_1679);
nor U942 (N_942,In_1326,In_618);
or U943 (N_943,In_1625,In_1071);
nand U944 (N_944,In_461,In_1052);
nand U945 (N_945,In_92,In_1843);
nor U946 (N_946,In_974,In_1004);
and U947 (N_947,In_1078,In_1179);
nand U948 (N_948,In_1739,In_1792);
nor U949 (N_949,In_336,In_97);
nor U950 (N_950,In_1042,In_445);
nor U951 (N_951,In_242,In_1956);
and U952 (N_952,In_408,In_888);
and U953 (N_953,In_1882,In_922);
nand U954 (N_954,In_322,In_400);
nand U955 (N_955,In_1265,In_1245);
nor U956 (N_956,In_636,In_1459);
nand U957 (N_957,In_1358,In_1215);
and U958 (N_958,In_302,In_1719);
nand U959 (N_959,In_1131,In_1810);
or U960 (N_960,In_1214,In_119);
nor U961 (N_961,In_121,In_1133);
and U962 (N_962,In_1060,In_1074);
and U963 (N_963,In_1533,In_1243);
nand U964 (N_964,In_1841,In_966);
nor U965 (N_965,In_781,In_689);
or U966 (N_966,In_848,In_1059);
nand U967 (N_967,In_1290,In_1012);
or U968 (N_968,In_904,In_377);
xor U969 (N_969,In_1196,In_383);
nand U970 (N_970,In_1281,In_1875);
and U971 (N_971,In_432,In_14);
nand U972 (N_972,In_770,In_564);
xnor U973 (N_973,In_530,In_585);
and U974 (N_974,In_1127,In_854);
and U975 (N_975,In_216,In_943);
and U976 (N_976,In_39,In_74);
or U977 (N_977,In_151,In_1582);
xnor U978 (N_978,In_1439,In_1623);
or U979 (N_979,In_25,In_510);
nor U980 (N_980,In_444,In_1434);
or U981 (N_981,In_1684,In_578);
or U982 (N_982,In_846,In_23);
nor U983 (N_983,In_664,In_18);
nand U984 (N_984,In_421,In_1121);
or U985 (N_985,In_440,In_334);
xnor U986 (N_986,In_397,In_761);
nor U987 (N_987,In_701,In_1992);
xor U988 (N_988,In_76,In_499);
or U989 (N_989,In_795,In_1045);
or U990 (N_990,In_1537,In_1654);
nand U991 (N_991,In_172,In_173);
nand U992 (N_992,In_1390,In_1485);
nor U993 (N_993,In_1940,In_1010);
or U994 (N_994,In_277,In_214);
or U995 (N_995,In_435,In_1973);
or U996 (N_996,In_941,In_1897);
nor U997 (N_997,In_871,In_162);
nand U998 (N_998,In_763,In_1418);
nand U999 (N_999,In_1283,In_1532);
or U1000 (N_1000,In_1657,In_849);
nand U1001 (N_1001,In_455,In_1776);
or U1002 (N_1002,In_1685,In_213);
xnor U1003 (N_1003,In_673,In_1948);
and U1004 (N_1004,In_305,In_727);
or U1005 (N_1005,In_254,In_593);
nor U1006 (N_1006,In_1794,In_123);
nand U1007 (N_1007,In_1091,In_1751);
nand U1008 (N_1008,In_569,In_1071);
or U1009 (N_1009,In_322,In_582);
and U1010 (N_1010,In_757,In_1861);
nor U1011 (N_1011,In_419,In_816);
or U1012 (N_1012,In_688,In_540);
and U1013 (N_1013,In_100,In_855);
nor U1014 (N_1014,In_1536,In_508);
and U1015 (N_1015,In_1663,In_42);
nor U1016 (N_1016,In_1360,In_832);
nor U1017 (N_1017,In_462,In_1313);
or U1018 (N_1018,In_1441,In_1893);
or U1019 (N_1019,In_1572,In_768);
and U1020 (N_1020,In_1125,In_1710);
nor U1021 (N_1021,In_1975,In_1574);
or U1022 (N_1022,In_868,In_1151);
nor U1023 (N_1023,In_882,In_442);
nand U1024 (N_1024,In_686,In_57);
nor U1025 (N_1025,In_1144,In_400);
nand U1026 (N_1026,In_636,In_1178);
or U1027 (N_1027,In_912,In_1006);
nand U1028 (N_1028,In_1191,In_1232);
xnor U1029 (N_1029,In_1142,In_724);
or U1030 (N_1030,In_255,In_867);
or U1031 (N_1031,In_1391,In_1946);
and U1032 (N_1032,In_236,In_414);
nand U1033 (N_1033,In_1008,In_1725);
nand U1034 (N_1034,In_199,In_1865);
and U1035 (N_1035,In_1902,In_563);
and U1036 (N_1036,In_1464,In_1827);
or U1037 (N_1037,In_1136,In_1459);
nand U1038 (N_1038,In_499,In_1474);
and U1039 (N_1039,In_1676,In_515);
or U1040 (N_1040,In_218,In_363);
and U1041 (N_1041,In_971,In_625);
nor U1042 (N_1042,In_998,In_544);
nand U1043 (N_1043,In_579,In_188);
or U1044 (N_1044,In_1501,In_1600);
and U1045 (N_1045,In_38,In_491);
and U1046 (N_1046,In_1526,In_560);
nor U1047 (N_1047,In_1793,In_1333);
nand U1048 (N_1048,In_522,In_1924);
nor U1049 (N_1049,In_1175,In_89);
nor U1050 (N_1050,In_709,In_163);
and U1051 (N_1051,In_1433,In_1706);
nand U1052 (N_1052,In_1479,In_770);
and U1053 (N_1053,In_1683,In_171);
and U1054 (N_1054,In_896,In_899);
and U1055 (N_1055,In_1741,In_1045);
or U1056 (N_1056,In_1957,In_451);
and U1057 (N_1057,In_352,In_831);
or U1058 (N_1058,In_1995,In_947);
or U1059 (N_1059,In_281,In_1159);
nand U1060 (N_1060,In_1266,In_810);
nand U1061 (N_1061,In_119,In_1244);
and U1062 (N_1062,In_1281,In_1000);
or U1063 (N_1063,In_152,In_1799);
and U1064 (N_1064,In_149,In_1104);
nand U1065 (N_1065,In_330,In_95);
nor U1066 (N_1066,In_648,In_549);
nand U1067 (N_1067,In_1309,In_96);
nor U1068 (N_1068,In_1259,In_1784);
nand U1069 (N_1069,In_347,In_943);
or U1070 (N_1070,In_1018,In_13);
nor U1071 (N_1071,In_1477,In_1987);
nor U1072 (N_1072,In_276,In_893);
nor U1073 (N_1073,In_1168,In_508);
or U1074 (N_1074,In_801,In_1438);
nand U1075 (N_1075,In_1372,In_1669);
and U1076 (N_1076,In_1506,In_1956);
and U1077 (N_1077,In_1689,In_717);
nand U1078 (N_1078,In_36,In_1574);
nor U1079 (N_1079,In_1657,In_1418);
nand U1080 (N_1080,In_530,In_250);
nand U1081 (N_1081,In_962,In_796);
and U1082 (N_1082,In_1358,In_450);
xor U1083 (N_1083,In_1457,In_1912);
nor U1084 (N_1084,In_774,In_731);
nor U1085 (N_1085,In_1700,In_1936);
or U1086 (N_1086,In_901,In_1636);
nand U1087 (N_1087,In_1877,In_1488);
nand U1088 (N_1088,In_1090,In_1591);
and U1089 (N_1089,In_5,In_1311);
or U1090 (N_1090,In_1840,In_451);
and U1091 (N_1091,In_1868,In_1519);
or U1092 (N_1092,In_1601,In_217);
or U1093 (N_1093,In_1269,In_1859);
and U1094 (N_1094,In_118,In_1471);
or U1095 (N_1095,In_546,In_249);
nor U1096 (N_1096,In_304,In_1339);
and U1097 (N_1097,In_611,In_1767);
or U1098 (N_1098,In_1547,In_1932);
nand U1099 (N_1099,In_1697,In_177);
xnor U1100 (N_1100,In_1317,In_1246);
nor U1101 (N_1101,In_1658,In_1471);
nand U1102 (N_1102,In_1722,In_1889);
nand U1103 (N_1103,In_1745,In_690);
or U1104 (N_1104,In_549,In_160);
xnor U1105 (N_1105,In_1576,In_1512);
nor U1106 (N_1106,In_434,In_1668);
xnor U1107 (N_1107,In_506,In_992);
nand U1108 (N_1108,In_1187,In_745);
xnor U1109 (N_1109,In_733,In_1400);
or U1110 (N_1110,In_321,In_1891);
nor U1111 (N_1111,In_1297,In_844);
nor U1112 (N_1112,In_711,In_1278);
nand U1113 (N_1113,In_1885,In_542);
nor U1114 (N_1114,In_591,In_1755);
nand U1115 (N_1115,In_84,In_34);
and U1116 (N_1116,In_1866,In_268);
nor U1117 (N_1117,In_352,In_1932);
or U1118 (N_1118,In_1588,In_88);
and U1119 (N_1119,In_411,In_1834);
or U1120 (N_1120,In_1320,In_1351);
nor U1121 (N_1121,In_1816,In_1383);
nand U1122 (N_1122,In_632,In_308);
and U1123 (N_1123,In_1536,In_1960);
or U1124 (N_1124,In_1014,In_1984);
and U1125 (N_1125,In_789,In_710);
xor U1126 (N_1126,In_1342,In_468);
or U1127 (N_1127,In_1403,In_238);
nand U1128 (N_1128,In_1800,In_39);
nor U1129 (N_1129,In_1580,In_1921);
or U1130 (N_1130,In_445,In_1818);
xnor U1131 (N_1131,In_1864,In_752);
and U1132 (N_1132,In_1517,In_1333);
xor U1133 (N_1133,In_912,In_438);
and U1134 (N_1134,In_748,In_1661);
nor U1135 (N_1135,In_731,In_1856);
or U1136 (N_1136,In_336,In_534);
nor U1137 (N_1137,In_1226,In_474);
and U1138 (N_1138,In_1635,In_728);
and U1139 (N_1139,In_864,In_719);
and U1140 (N_1140,In_1443,In_1355);
and U1141 (N_1141,In_1165,In_1016);
nand U1142 (N_1142,In_845,In_1889);
nand U1143 (N_1143,In_842,In_1627);
and U1144 (N_1144,In_112,In_187);
and U1145 (N_1145,In_1650,In_1508);
nand U1146 (N_1146,In_1028,In_993);
nor U1147 (N_1147,In_1409,In_1355);
and U1148 (N_1148,In_393,In_1312);
nor U1149 (N_1149,In_1330,In_1942);
or U1150 (N_1150,In_547,In_1221);
nor U1151 (N_1151,In_405,In_899);
nor U1152 (N_1152,In_1654,In_520);
nor U1153 (N_1153,In_1355,In_748);
or U1154 (N_1154,In_1096,In_541);
or U1155 (N_1155,In_1412,In_1067);
and U1156 (N_1156,In_1876,In_540);
xnor U1157 (N_1157,In_1218,In_1262);
nand U1158 (N_1158,In_116,In_315);
nand U1159 (N_1159,In_1384,In_970);
nand U1160 (N_1160,In_276,In_1464);
and U1161 (N_1161,In_1449,In_1501);
xor U1162 (N_1162,In_0,In_1841);
or U1163 (N_1163,In_908,In_116);
or U1164 (N_1164,In_1172,In_942);
and U1165 (N_1165,In_418,In_225);
and U1166 (N_1166,In_1083,In_273);
nand U1167 (N_1167,In_1243,In_879);
and U1168 (N_1168,In_101,In_735);
nand U1169 (N_1169,In_1415,In_230);
nand U1170 (N_1170,In_1906,In_1738);
xor U1171 (N_1171,In_982,In_828);
nand U1172 (N_1172,In_563,In_1613);
and U1173 (N_1173,In_1004,In_1138);
nand U1174 (N_1174,In_32,In_969);
nand U1175 (N_1175,In_1499,In_234);
nor U1176 (N_1176,In_827,In_291);
nand U1177 (N_1177,In_447,In_723);
or U1178 (N_1178,In_125,In_1098);
or U1179 (N_1179,In_1345,In_1639);
nand U1180 (N_1180,In_1899,In_167);
nor U1181 (N_1181,In_1542,In_218);
nor U1182 (N_1182,In_751,In_161);
nand U1183 (N_1183,In_488,In_651);
nand U1184 (N_1184,In_1441,In_1739);
nand U1185 (N_1185,In_507,In_1835);
or U1186 (N_1186,In_3,In_898);
and U1187 (N_1187,In_1920,In_115);
xor U1188 (N_1188,In_1340,In_1906);
xor U1189 (N_1189,In_1345,In_1508);
nand U1190 (N_1190,In_1340,In_886);
xnor U1191 (N_1191,In_1012,In_1582);
or U1192 (N_1192,In_840,In_1898);
or U1193 (N_1193,In_905,In_1965);
or U1194 (N_1194,In_70,In_942);
and U1195 (N_1195,In_1980,In_900);
nand U1196 (N_1196,In_1007,In_310);
nor U1197 (N_1197,In_851,In_1109);
and U1198 (N_1198,In_555,In_259);
and U1199 (N_1199,In_455,In_1286);
or U1200 (N_1200,In_1035,In_1755);
and U1201 (N_1201,In_74,In_877);
or U1202 (N_1202,In_1369,In_518);
nor U1203 (N_1203,In_1548,In_248);
or U1204 (N_1204,In_1285,In_1220);
and U1205 (N_1205,In_339,In_1948);
nor U1206 (N_1206,In_1863,In_1739);
nor U1207 (N_1207,In_1733,In_1453);
nor U1208 (N_1208,In_122,In_268);
nand U1209 (N_1209,In_763,In_127);
or U1210 (N_1210,In_691,In_89);
nand U1211 (N_1211,In_614,In_1502);
xor U1212 (N_1212,In_947,In_1011);
nor U1213 (N_1213,In_1839,In_1945);
nand U1214 (N_1214,In_871,In_1306);
nand U1215 (N_1215,In_901,In_962);
or U1216 (N_1216,In_1523,In_1242);
nand U1217 (N_1217,In_1803,In_1783);
xnor U1218 (N_1218,In_1787,In_1874);
nand U1219 (N_1219,In_1516,In_358);
nor U1220 (N_1220,In_1703,In_633);
nor U1221 (N_1221,In_576,In_1786);
nand U1222 (N_1222,In_6,In_1891);
or U1223 (N_1223,In_332,In_1410);
and U1224 (N_1224,In_1009,In_62);
or U1225 (N_1225,In_1365,In_1656);
nor U1226 (N_1226,In_1422,In_1588);
nand U1227 (N_1227,In_1954,In_766);
nand U1228 (N_1228,In_194,In_707);
nand U1229 (N_1229,In_617,In_1767);
xor U1230 (N_1230,In_688,In_1091);
nand U1231 (N_1231,In_1447,In_1970);
or U1232 (N_1232,In_763,In_292);
nor U1233 (N_1233,In_1858,In_415);
xor U1234 (N_1234,In_647,In_1601);
nor U1235 (N_1235,In_1252,In_268);
nand U1236 (N_1236,In_991,In_838);
nor U1237 (N_1237,In_1693,In_1554);
nor U1238 (N_1238,In_285,In_266);
nand U1239 (N_1239,In_1645,In_849);
or U1240 (N_1240,In_1438,In_61);
or U1241 (N_1241,In_150,In_1175);
and U1242 (N_1242,In_1255,In_1915);
or U1243 (N_1243,In_1150,In_1184);
nor U1244 (N_1244,In_1026,In_1840);
nand U1245 (N_1245,In_1334,In_1253);
nor U1246 (N_1246,In_113,In_644);
or U1247 (N_1247,In_1126,In_1583);
nand U1248 (N_1248,In_1570,In_155);
nand U1249 (N_1249,In_464,In_1835);
or U1250 (N_1250,In_1990,In_1400);
and U1251 (N_1251,In_1765,In_474);
nand U1252 (N_1252,In_1803,In_125);
and U1253 (N_1253,In_1232,In_697);
nor U1254 (N_1254,In_789,In_1369);
nand U1255 (N_1255,In_949,In_552);
or U1256 (N_1256,In_1149,In_1947);
or U1257 (N_1257,In_1698,In_411);
xor U1258 (N_1258,In_511,In_682);
or U1259 (N_1259,In_1821,In_1896);
nor U1260 (N_1260,In_479,In_1601);
nor U1261 (N_1261,In_427,In_621);
xnor U1262 (N_1262,In_971,In_1753);
or U1263 (N_1263,In_121,In_1297);
and U1264 (N_1264,In_1017,In_775);
or U1265 (N_1265,In_1846,In_944);
nor U1266 (N_1266,In_201,In_501);
nor U1267 (N_1267,In_1697,In_1354);
nor U1268 (N_1268,In_1687,In_1708);
nand U1269 (N_1269,In_1445,In_1858);
xnor U1270 (N_1270,In_349,In_295);
or U1271 (N_1271,In_1303,In_875);
nor U1272 (N_1272,In_1274,In_463);
nand U1273 (N_1273,In_1730,In_811);
nand U1274 (N_1274,In_972,In_666);
nand U1275 (N_1275,In_846,In_1744);
and U1276 (N_1276,In_37,In_801);
nand U1277 (N_1277,In_1818,In_1500);
and U1278 (N_1278,In_1550,In_1349);
or U1279 (N_1279,In_1726,In_1019);
xnor U1280 (N_1280,In_200,In_1105);
or U1281 (N_1281,In_891,In_1491);
nor U1282 (N_1282,In_1808,In_683);
and U1283 (N_1283,In_1767,In_1563);
nand U1284 (N_1284,In_739,In_1785);
xor U1285 (N_1285,In_1537,In_1054);
nor U1286 (N_1286,In_342,In_756);
or U1287 (N_1287,In_1112,In_1487);
nor U1288 (N_1288,In_850,In_532);
xnor U1289 (N_1289,In_14,In_440);
nor U1290 (N_1290,In_921,In_1286);
xnor U1291 (N_1291,In_614,In_1443);
xor U1292 (N_1292,In_1758,In_684);
and U1293 (N_1293,In_230,In_1352);
nand U1294 (N_1294,In_1403,In_702);
and U1295 (N_1295,In_1215,In_1145);
nand U1296 (N_1296,In_1195,In_838);
nor U1297 (N_1297,In_989,In_1249);
and U1298 (N_1298,In_679,In_469);
nor U1299 (N_1299,In_65,In_889);
xor U1300 (N_1300,In_241,In_1239);
or U1301 (N_1301,In_1991,In_1859);
and U1302 (N_1302,In_1303,In_1147);
nor U1303 (N_1303,In_1130,In_1805);
and U1304 (N_1304,In_919,In_1406);
nor U1305 (N_1305,In_524,In_30);
and U1306 (N_1306,In_1456,In_1953);
and U1307 (N_1307,In_940,In_821);
or U1308 (N_1308,In_1662,In_1249);
nand U1309 (N_1309,In_1022,In_188);
or U1310 (N_1310,In_479,In_1631);
xnor U1311 (N_1311,In_488,In_797);
nand U1312 (N_1312,In_678,In_1523);
xor U1313 (N_1313,In_1653,In_18);
nand U1314 (N_1314,In_1705,In_1591);
nand U1315 (N_1315,In_401,In_704);
and U1316 (N_1316,In_275,In_208);
and U1317 (N_1317,In_854,In_729);
or U1318 (N_1318,In_721,In_732);
and U1319 (N_1319,In_1005,In_135);
nor U1320 (N_1320,In_1680,In_1259);
nand U1321 (N_1321,In_797,In_1258);
and U1322 (N_1322,In_1268,In_1851);
nor U1323 (N_1323,In_1697,In_1247);
and U1324 (N_1324,In_689,In_397);
and U1325 (N_1325,In_1496,In_725);
or U1326 (N_1326,In_1778,In_1860);
nor U1327 (N_1327,In_299,In_67);
nand U1328 (N_1328,In_1005,In_612);
nand U1329 (N_1329,In_1616,In_684);
nand U1330 (N_1330,In_303,In_1027);
nor U1331 (N_1331,In_1927,In_151);
and U1332 (N_1332,In_1819,In_1602);
xor U1333 (N_1333,In_1043,In_558);
nor U1334 (N_1334,In_1059,In_453);
nand U1335 (N_1335,In_1301,In_355);
nand U1336 (N_1336,In_587,In_1145);
nand U1337 (N_1337,In_393,In_1022);
and U1338 (N_1338,In_621,In_1602);
xnor U1339 (N_1339,In_864,In_90);
nand U1340 (N_1340,In_1887,In_557);
or U1341 (N_1341,In_894,In_1877);
nor U1342 (N_1342,In_403,In_474);
or U1343 (N_1343,In_1643,In_695);
or U1344 (N_1344,In_1589,In_1285);
nand U1345 (N_1345,In_1442,In_1620);
or U1346 (N_1346,In_793,In_1786);
or U1347 (N_1347,In_989,In_687);
nor U1348 (N_1348,In_335,In_349);
nand U1349 (N_1349,In_699,In_1297);
or U1350 (N_1350,In_1084,In_331);
or U1351 (N_1351,In_1515,In_69);
or U1352 (N_1352,In_1136,In_1059);
nor U1353 (N_1353,In_1916,In_1832);
nor U1354 (N_1354,In_798,In_11);
and U1355 (N_1355,In_1463,In_1418);
xnor U1356 (N_1356,In_1717,In_731);
nor U1357 (N_1357,In_49,In_1698);
nor U1358 (N_1358,In_1979,In_304);
and U1359 (N_1359,In_670,In_388);
and U1360 (N_1360,In_640,In_887);
or U1361 (N_1361,In_866,In_1287);
xor U1362 (N_1362,In_1284,In_46);
or U1363 (N_1363,In_68,In_679);
nor U1364 (N_1364,In_1104,In_1360);
nand U1365 (N_1365,In_661,In_1206);
xor U1366 (N_1366,In_1350,In_1359);
xnor U1367 (N_1367,In_1535,In_1105);
xor U1368 (N_1368,In_1501,In_35);
nand U1369 (N_1369,In_990,In_896);
nand U1370 (N_1370,In_1507,In_972);
or U1371 (N_1371,In_742,In_1816);
or U1372 (N_1372,In_1684,In_1249);
nor U1373 (N_1373,In_556,In_731);
nor U1374 (N_1374,In_487,In_1534);
nand U1375 (N_1375,In_1397,In_1803);
and U1376 (N_1376,In_153,In_606);
or U1377 (N_1377,In_592,In_1643);
nor U1378 (N_1378,In_819,In_538);
nand U1379 (N_1379,In_1893,In_357);
nor U1380 (N_1380,In_1455,In_962);
or U1381 (N_1381,In_1884,In_210);
nor U1382 (N_1382,In_1868,In_1812);
nand U1383 (N_1383,In_1714,In_750);
and U1384 (N_1384,In_1173,In_689);
nor U1385 (N_1385,In_1967,In_420);
and U1386 (N_1386,In_728,In_991);
nor U1387 (N_1387,In_710,In_1552);
nor U1388 (N_1388,In_1200,In_1545);
nor U1389 (N_1389,In_1998,In_615);
nor U1390 (N_1390,In_1836,In_1835);
nand U1391 (N_1391,In_963,In_453);
or U1392 (N_1392,In_601,In_189);
nor U1393 (N_1393,In_1031,In_1069);
or U1394 (N_1394,In_589,In_270);
and U1395 (N_1395,In_1387,In_736);
and U1396 (N_1396,In_1207,In_1196);
nor U1397 (N_1397,In_1593,In_871);
and U1398 (N_1398,In_383,In_1201);
nor U1399 (N_1399,In_873,In_1278);
and U1400 (N_1400,In_965,In_1426);
nand U1401 (N_1401,In_1652,In_64);
nor U1402 (N_1402,In_1852,In_1605);
and U1403 (N_1403,In_1138,In_611);
and U1404 (N_1404,In_821,In_214);
nand U1405 (N_1405,In_1339,In_1793);
nand U1406 (N_1406,In_46,In_397);
nand U1407 (N_1407,In_1995,In_828);
and U1408 (N_1408,In_1685,In_1845);
and U1409 (N_1409,In_94,In_1778);
and U1410 (N_1410,In_1458,In_786);
nand U1411 (N_1411,In_700,In_1699);
nor U1412 (N_1412,In_239,In_106);
nor U1413 (N_1413,In_1320,In_1947);
xnor U1414 (N_1414,In_731,In_1518);
and U1415 (N_1415,In_72,In_396);
or U1416 (N_1416,In_1382,In_1576);
or U1417 (N_1417,In_367,In_1861);
nor U1418 (N_1418,In_1521,In_554);
and U1419 (N_1419,In_806,In_1878);
or U1420 (N_1420,In_1305,In_49);
nand U1421 (N_1421,In_1913,In_1310);
xnor U1422 (N_1422,In_1148,In_116);
nor U1423 (N_1423,In_1778,In_1389);
or U1424 (N_1424,In_418,In_1464);
xnor U1425 (N_1425,In_949,In_752);
nand U1426 (N_1426,In_365,In_785);
nor U1427 (N_1427,In_1221,In_404);
nor U1428 (N_1428,In_741,In_160);
nand U1429 (N_1429,In_1120,In_708);
nand U1430 (N_1430,In_479,In_1556);
and U1431 (N_1431,In_207,In_831);
nand U1432 (N_1432,In_1827,In_939);
nor U1433 (N_1433,In_320,In_787);
nor U1434 (N_1434,In_1644,In_600);
nand U1435 (N_1435,In_119,In_1869);
nand U1436 (N_1436,In_370,In_1985);
nand U1437 (N_1437,In_1456,In_1774);
nand U1438 (N_1438,In_849,In_404);
or U1439 (N_1439,In_46,In_1830);
xor U1440 (N_1440,In_1211,In_1234);
and U1441 (N_1441,In_1519,In_594);
nor U1442 (N_1442,In_1533,In_979);
or U1443 (N_1443,In_905,In_1074);
nand U1444 (N_1444,In_523,In_1630);
nand U1445 (N_1445,In_1272,In_1653);
xnor U1446 (N_1446,In_890,In_1811);
and U1447 (N_1447,In_551,In_376);
xor U1448 (N_1448,In_896,In_136);
and U1449 (N_1449,In_1298,In_653);
or U1450 (N_1450,In_472,In_1252);
or U1451 (N_1451,In_493,In_247);
nor U1452 (N_1452,In_1542,In_134);
and U1453 (N_1453,In_108,In_643);
or U1454 (N_1454,In_661,In_1569);
nor U1455 (N_1455,In_1718,In_1776);
and U1456 (N_1456,In_1982,In_1922);
nor U1457 (N_1457,In_304,In_1054);
or U1458 (N_1458,In_191,In_1020);
or U1459 (N_1459,In_467,In_1022);
xor U1460 (N_1460,In_1736,In_813);
or U1461 (N_1461,In_618,In_1138);
xor U1462 (N_1462,In_414,In_1722);
xor U1463 (N_1463,In_348,In_654);
or U1464 (N_1464,In_698,In_148);
or U1465 (N_1465,In_555,In_311);
or U1466 (N_1466,In_1870,In_1358);
nor U1467 (N_1467,In_647,In_912);
and U1468 (N_1468,In_20,In_103);
and U1469 (N_1469,In_1583,In_810);
nor U1470 (N_1470,In_249,In_730);
nand U1471 (N_1471,In_756,In_1646);
nor U1472 (N_1472,In_369,In_1424);
and U1473 (N_1473,In_1057,In_1863);
nand U1474 (N_1474,In_310,In_1485);
nand U1475 (N_1475,In_1359,In_290);
nor U1476 (N_1476,In_570,In_1550);
and U1477 (N_1477,In_507,In_483);
nand U1478 (N_1478,In_1499,In_1525);
nand U1479 (N_1479,In_903,In_1586);
xnor U1480 (N_1480,In_1180,In_639);
nand U1481 (N_1481,In_142,In_1374);
nor U1482 (N_1482,In_1926,In_795);
or U1483 (N_1483,In_1340,In_1955);
and U1484 (N_1484,In_1574,In_1506);
or U1485 (N_1485,In_702,In_115);
or U1486 (N_1486,In_348,In_945);
xor U1487 (N_1487,In_647,In_1982);
or U1488 (N_1488,In_1882,In_1663);
and U1489 (N_1489,In_943,In_1371);
nor U1490 (N_1490,In_353,In_833);
xnor U1491 (N_1491,In_1601,In_1984);
and U1492 (N_1492,In_1514,In_1463);
nand U1493 (N_1493,In_1903,In_181);
nor U1494 (N_1494,In_260,In_1957);
nand U1495 (N_1495,In_1519,In_1590);
or U1496 (N_1496,In_1672,In_925);
nor U1497 (N_1497,In_1247,In_1347);
nor U1498 (N_1498,In_431,In_1488);
nand U1499 (N_1499,In_1047,In_335);
and U1500 (N_1500,In_1899,In_578);
and U1501 (N_1501,In_1095,In_681);
nand U1502 (N_1502,In_1497,In_672);
or U1503 (N_1503,In_554,In_249);
nor U1504 (N_1504,In_1886,In_68);
nor U1505 (N_1505,In_1957,In_848);
xnor U1506 (N_1506,In_1576,In_1426);
nand U1507 (N_1507,In_318,In_1969);
xor U1508 (N_1508,In_468,In_326);
nand U1509 (N_1509,In_1589,In_1348);
nor U1510 (N_1510,In_529,In_1408);
nor U1511 (N_1511,In_37,In_515);
and U1512 (N_1512,In_1336,In_722);
nor U1513 (N_1513,In_458,In_1567);
and U1514 (N_1514,In_1235,In_570);
or U1515 (N_1515,In_470,In_988);
or U1516 (N_1516,In_783,In_310);
or U1517 (N_1517,In_772,In_653);
nand U1518 (N_1518,In_622,In_743);
and U1519 (N_1519,In_433,In_506);
nor U1520 (N_1520,In_498,In_1844);
xnor U1521 (N_1521,In_789,In_87);
nor U1522 (N_1522,In_1246,In_196);
nand U1523 (N_1523,In_20,In_921);
or U1524 (N_1524,In_929,In_427);
nand U1525 (N_1525,In_276,In_1896);
nand U1526 (N_1526,In_106,In_1943);
and U1527 (N_1527,In_330,In_1342);
nor U1528 (N_1528,In_14,In_1855);
nor U1529 (N_1529,In_558,In_1209);
or U1530 (N_1530,In_962,In_525);
nand U1531 (N_1531,In_1067,In_1639);
nor U1532 (N_1532,In_677,In_1259);
nor U1533 (N_1533,In_1182,In_1830);
nand U1534 (N_1534,In_1154,In_393);
xnor U1535 (N_1535,In_844,In_943);
and U1536 (N_1536,In_1370,In_1450);
nor U1537 (N_1537,In_770,In_1321);
nor U1538 (N_1538,In_320,In_1732);
or U1539 (N_1539,In_520,In_1001);
nor U1540 (N_1540,In_351,In_1984);
or U1541 (N_1541,In_124,In_1925);
or U1542 (N_1542,In_1128,In_1296);
or U1543 (N_1543,In_320,In_1115);
nand U1544 (N_1544,In_1216,In_1530);
or U1545 (N_1545,In_1190,In_540);
xor U1546 (N_1546,In_1450,In_124);
nand U1547 (N_1547,In_322,In_1802);
xnor U1548 (N_1548,In_936,In_1701);
nor U1549 (N_1549,In_374,In_1388);
nand U1550 (N_1550,In_618,In_1485);
nor U1551 (N_1551,In_20,In_1609);
and U1552 (N_1552,In_667,In_708);
or U1553 (N_1553,In_1243,In_960);
nor U1554 (N_1554,In_653,In_1548);
or U1555 (N_1555,In_1892,In_1939);
nand U1556 (N_1556,In_434,In_1950);
or U1557 (N_1557,In_1406,In_570);
nand U1558 (N_1558,In_140,In_1303);
nor U1559 (N_1559,In_1653,In_355);
nand U1560 (N_1560,In_577,In_1456);
nand U1561 (N_1561,In_274,In_749);
or U1562 (N_1562,In_404,In_797);
and U1563 (N_1563,In_98,In_937);
or U1564 (N_1564,In_1016,In_1965);
nand U1565 (N_1565,In_1599,In_1577);
nor U1566 (N_1566,In_1432,In_308);
xnor U1567 (N_1567,In_400,In_1184);
and U1568 (N_1568,In_885,In_1242);
and U1569 (N_1569,In_227,In_964);
nor U1570 (N_1570,In_1862,In_1586);
nand U1571 (N_1571,In_1692,In_706);
xnor U1572 (N_1572,In_759,In_342);
and U1573 (N_1573,In_756,In_1266);
nand U1574 (N_1574,In_1881,In_1957);
nand U1575 (N_1575,In_19,In_292);
or U1576 (N_1576,In_470,In_1761);
nand U1577 (N_1577,In_1878,In_788);
nor U1578 (N_1578,In_482,In_684);
nor U1579 (N_1579,In_105,In_1771);
xor U1580 (N_1580,In_102,In_1719);
and U1581 (N_1581,In_152,In_1174);
or U1582 (N_1582,In_1444,In_473);
and U1583 (N_1583,In_1680,In_1763);
and U1584 (N_1584,In_206,In_1846);
or U1585 (N_1585,In_1182,In_6);
and U1586 (N_1586,In_1050,In_1777);
nand U1587 (N_1587,In_841,In_20);
nor U1588 (N_1588,In_1041,In_1682);
or U1589 (N_1589,In_1033,In_461);
and U1590 (N_1590,In_292,In_676);
and U1591 (N_1591,In_894,In_795);
or U1592 (N_1592,In_719,In_526);
and U1593 (N_1593,In_1505,In_1530);
or U1594 (N_1594,In_1935,In_1812);
nor U1595 (N_1595,In_1164,In_1119);
and U1596 (N_1596,In_1467,In_385);
nor U1597 (N_1597,In_252,In_536);
nor U1598 (N_1598,In_546,In_1706);
xnor U1599 (N_1599,In_1354,In_1150);
nand U1600 (N_1600,In_1433,In_878);
or U1601 (N_1601,In_910,In_1298);
nand U1602 (N_1602,In_1357,In_1512);
nor U1603 (N_1603,In_1727,In_1869);
and U1604 (N_1604,In_1048,In_36);
or U1605 (N_1605,In_1192,In_1252);
nor U1606 (N_1606,In_132,In_1579);
nor U1607 (N_1607,In_942,In_465);
nand U1608 (N_1608,In_370,In_337);
nor U1609 (N_1609,In_1195,In_363);
nor U1610 (N_1610,In_284,In_1229);
xor U1611 (N_1611,In_1345,In_183);
nand U1612 (N_1612,In_253,In_110);
and U1613 (N_1613,In_211,In_320);
nand U1614 (N_1614,In_7,In_5);
or U1615 (N_1615,In_1994,In_1528);
and U1616 (N_1616,In_196,In_1879);
and U1617 (N_1617,In_100,In_543);
or U1618 (N_1618,In_1050,In_1998);
xor U1619 (N_1619,In_235,In_1032);
nand U1620 (N_1620,In_1960,In_1420);
or U1621 (N_1621,In_1923,In_1508);
nand U1622 (N_1622,In_8,In_1540);
nor U1623 (N_1623,In_469,In_1832);
nand U1624 (N_1624,In_784,In_1053);
or U1625 (N_1625,In_1121,In_1278);
or U1626 (N_1626,In_992,In_86);
or U1627 (N_1627,In_45,In_251);
nor U1628 (N_1628,In_1175,In_10);
and U1629 (N_1629,In_1831,In_340);
and U1630 (N_1630,In_1751,In_968);
xor U1631 (N_1631,In_142,In_1521);
nand U1632 (N_1632,In_730,In_784);
and U1633 (N_1633,In_311,In_70);
and U1634 (N_1634,In_1405,In_1399);
nor U1635 (N_1635,In_483,In_927);
nand U1636 (N_1636,In_10,In_1337);
and U1637 (N_1637,In_1713,In_1631);
nand U1638 (N_1638,In_507,In_1791);
and U1639 (N_1639,In_437,In_368);
nor U1640 (N_1640,In_627,In_819);
and U1641 (N_1641,In_353,In_441);
nand U1642 (N_1642,In_931,In_1034);
nor U1643 (N_1643,In_1485,In_623);
or U1644 (N_1644,In_262,In_751);
or U1645 (N_1645,In_119,In_1752);
xnor U1646 (N_1646,In_1475,In_1682);
xnor U1647 (N_1647,In_692,In_822);
or U1648 (N_1648,In_722,In_1617);
and U1649 (N_1649,In_877,In_1381);
or U1650 (N_1650,In_920,In_694);
nor U1651 (N_1651,In_321,In_197);
and U1652 (N_1652,In_1440,In_997);
or U1653 (N_1653,In_1308,In_629);
xnor U1654 (N_1654,In_367,In_1767);
xnor U1655 (N_1655,In_846,In_658);
nor U1656 (N_1656,In_1534,In_1773);
nor U1657 (N_1657,In_1041,In_1564);
or U1658 (N_1658,In_752,In_1256);
nor U1659 (N_1659,In_168,In_1598);
or U1660 (N_1660,In_1570,In_526);
or U1661 (N_1661,In_1418,In_1564);
or U1662 (N_1662,In_1025,In_265);
and U1663 (N_1663,In_1179,In_882);
nand U1664 (N_1664,In_1565,In_398);
nor U1665 (N_1665,In_1621,In_79);
nand U1666 (N_1666,In_763,In_975);
nand U1667 (N_1667,In_566,In_721);
nand U1668 (N_1668,In_1891,In_1538);
xor U1669 (N_1669,In_871,In_844);
and U1670 (N_1670,In_114,In_432);
nor U1671 (N_1671,In_301,In_1557);
and U1672 (N_1672,In_117,In_772);
or U1673 (N_1673,In_610,In_814);
or U1674 (N_1674,In_558,In_846);
xnor U1675 (N_1675,In_477,In_847);
or U1676 (N_1676,In_642,In_419);
and U1677 (N_1677,In_286,In_307);
xnor U1678 (N_1678,In_99,In_755);
and U1679 (N_1679,In_323,In_1569);
nand U1680 (N_1680,In_1839,In_92);
nor U1681 (N_1681,In_429,In_778);
and U1682 (N_1682,In_1611,In_1035);
xor U1683 (N_1683,In_1469,In_709);
and U1684 (N_1684,In_671,In_1290);
nand U1685 (N_1685,In_892,In_1143);
or U1686 (N_1686,In_1099,In_910);
or U1687 (N_1687,In_575,In_224);
and U1688 (N_1688,In_1066,In_143);
nor U1689 (N_1689,In_585,In_1466);
and U1690 (N_1690,In_1492,In_82);
nand U1691 (N_1691,In_901,In_23);
and U1692 (N_1692,In_1842,In_799);
and U1693 (N_1693,In_659,In_294);
and U1694 (N_1694,In_1538,In_1159);
or U1695 (N_1695,In_880,In_1117);
nand U1696 (N_1696,In_304,In_1277);
and U1697 (N_1697,In_1818,In_1909);
nor U1698 (N_1698,In_1991,In_1727);
nand U1699 (N_1699,In_218,In_30);
xor U1700 (N_1700,In_1166,In_584);
and U1701 (N_1701,In_1975,In_464);
nor U1702 (N_1702,In_1887,In_419);
nor U1703 (N_1703,In_1819,In_1522);
and U1704 (N_1704,In_1379,In_1100);
or U1705 (N_1705,In_1646,In_866);
or U1706 (N_1706,In_70,In_338);
nand U1707 (N_1707,In_1180,In_1753);
and U1708 (N_1708,In_421,In_866);
or U1709 (N_1709,In_180,In_26);
and U1710 (N_1710,In_1576,In_41);
and U1711 (N_1711,In_1158,In_126);
or U1712 (N_1712,In_1661,In_1810);
and U1713 (N_1713,In_1559,In_1975);
nor U1714 (N_1714,In_563,In_343);
or U1715 (N_1715,In_846,In_508);
and U1716 (N_1716,In_1324,In_1645);
or U1717 (N_1717,In_1310,In_208);
or U1718 (N_1718,In_246,In_928);
nor U1719 (N_1719,In_1727,In_1065);
xnor U1720 (N_1720,In_1617,In_1897);
nand U1721 (N_1721,In_1295,In_4);
or U1722 (N_1722,In_704,In_798);
nor U1723 (N_1723,In_972,In_408);
and U1724 (N_1724,In_27,In_1826);
nand U1725 (N_1725,In_380,In_1004);
or U1726 (N_1726,In_1514,In_307);
xnor U1727 (N_1727,In_166,In_1085);
or U1728 (N_1728,In_1384,In_248);
nor U1729 (N_1729,In_1590,In_1515);
and U1730 (N_1730,In_1166,In_109);
or U1731 (N_1731,In_444,In_670);
nand U1732 (N_1732,In_667,In_1994);
nor U1733 (N_1733,In_1479,In_1686);
and U1734 (N_1734,In_1277,In_1871);
nor U1735 (N_1735,In_673,In_1592);
nor U1736 (N_1736,In_372,In_602);
nor U1737 (N_1737,In_293,In_1452);
and U1738 (N_1738,In_1849,In_840);
and U1739 (N_1739,In_850,In_1599);
and U1740 (N_1740,In_1313,In_1331);
nor U1741 (N_1741,In_1799,In_1575);
nor U1742 (N_1742,In_1400,In_1533);
or U1743 (N_1743,In_826,In_729);
and U1744 (N_1744,In_1323,In_1737);
nor U1745 (N_1745,In_327,In_408);
nor U1746 (N_1746,In_1500,In_331);
or U1747 (N_1747,In_224,In_919);
nand U1748 (N_1748,In_215,In_1406);
nor U1749 (N_1749,In_651,In_726);
nand U1750 (N_1750,In_1678,In_906);
nand U1751 (N_1751,In_38,In_1405);
or U1752 (N_1752,In_929,In_431);
or U1753 (N_1753,In_271,In_140);
nor U1754 (N_1754,In_728,In_863);
nand U1755 (N_1755,In_1251,In_1392);
and U1756 (N_1756,In_926,In_1601);
or U1757 (N_1757,In_1175,In_891);
or U1758 (N_1758,In_206,In_838);
nand U1759 (N_1759,In_444,In_874);
nand U1760 (N_1760,In_132,In_855);
or U1761 (N_1761,In_546,In_1060);
and U1762 (N_1762,In_846,In_1923);
xor U1763 (N_1763,In_1601,In_366);
nor U1764 (N_1764,In_899,In_97);
or U1765 (N_1765,In_1521,In_417);
and U1766 (N_1766,In_27,In_1182);
xnor U1767 (N_1767,In_1621,In_904);
or U1768 (N_1768,In_1085,In_820);
nand U1769 (N_1769,In_1920,In_981);
and U1770 (N_1770,In_313,In_86);
nor U1771 (N_1771,In_1525,In_150);
and U1772 (N_1772,In_1837,In_568);
nand U1773 (N_1773,In_351,In_381);
nor U1774 (N_1774,In_955,In_1471);
nand U1775 (N_1775,In_1210,In_1173);
or U1776 (N_1776,In_706,In_1571);
nor U1777 (N_1777,In_593,In_1083);
nand U1778 (N_1778,In_1696,In_1627);
nor U1779 (N_1779,In_144,In_150);
nand U1780 (N_1780,In_703,In_291);
xnor U1781 (N_1781,In_631,In_684);
and U1782 (N_1782,In_1400,In_118);
or U1783 (N_1783,In_176,In_912);
or U1784 (N_1784,In_199,In_561);
or U1785 (N_1785,In_1522,In_1728);
nand U1786 (N_1786,In_98,In_1474);
and U1787 (N_1787,In_168,In_209);
nand U1788 (N_1788,In_970,In_689);
nor U1789 (N_1789,In_449,In_1198);
xor U1790 (N_1790,In_1924,In_1197);
xnor U1791 (N_1791,In_1509,In_1165);
nor U1792 (N_1792,In_395,In_1487);
xor U1793 (N_1793,In_987,In_1602);
and U1794 (N_1794,In_1487,In_733);
xor U1795 (N_1795,In_1762,In_1568);
xor U1796 (N_1796,In_1478,In_821);
or U1797 (N_1797,In_475,In_103);
nor U1798 (N_1798,In_72,In_440);
nand U1799 (N_1799,In_1484,In_1830);
nor U1800 (N_1800,In_1085,In_125);
nand U1801 (N_1801,In_1804,In_6);
nand U1802 (N_1802,In_1775,In_423);
and U1803 (N_1803,In_397,In_423);
or U1804 (N_1804,In_351,In_511);
and U1805 (N_1805,In_1922,In_371);
nand U1806 (N_1806,In_50,In_164);
nor U1807 (N_1807,In_320,In_782);
xor U1808 (N_1808,In_1865,In_1845);
and U1809 (N_1809,In_1071,In_1681);
nand U1810 (N_1810,In_1255,In_1547);
and U1811 (N_1811,In_952,In_987);
or U1812 (N_1812,In_1571,In_987);
or U1813 (N_1813,In_1602,In_843);
or U1814 (N_1814,In_1412,In_81);
nand U1815 (N_1815,In_1608,In_1234);
xor U1816 (N_1816,In_1519,In_57);
nand U1817 (N_1817,In_1690,In_121);
and U1818 (N_1818,In_261,In_1224);
and U1819 (N_1819,In_431,In_738);
and U1820 (N_1820,In_591,In_206);
nor U1821 (N_1821,In_1950,In_609);
nand U1822 (N_1822,In_709,In_804);
and U1823 (N_1823,In_219,In_696);
nor U1824 (N_1824,In_1996,In_1676);
nand U1825 (N_1825,In_983,In_801);
and U1826 (N_1826,In_973,In_533);
and U1827 (N_1827,In_108,In_865);
or U1828 (N_1828,In_700,In_1847);
and U1829 (N_1829,In_1894,In_1928);
nand U1830 (N_1830,In_274,In_648);
xnor U1831 (N_1831,In_401,In_1310);
and U1832 (N_1832,In_1905,In_1726);
nor U1833 (N_1833,In_1074,In_1867);
nand U1834 (N_1834,In_1097,In_1454);
xor U1835 (N_1835,In_276,In_1503);
nand U1836 (N_1836,In_9,In_1832);
xor U1837 (N_1837,In_1596,In_1038);
nor U1838 (N_1838,In_866,In_1294);
nor U1839 (N_1839,In_1229,In_270);
nor U1840 (N_1840,In_212,In_1368);
and U1841 (N_1841,In_399,In_792);
nor U1842 (N_1842,In_594,In_66);
nand U1843 (N_1843,In_739,In_720);
xnor U1844 (N_1844,In_679,In_1389);
nand U1845 (N_1845,In_118,In_1725);
or U1846 (N_1846,In_1232,In_1766);
and U1847 (N_1847,In_603,In_1065);
or U1848 (N_1848,In_1541,In_366);
nor U1849 (N_1849,In_931,In_235);
nand U1850 (N_1850,In_323,In_447);
and U1851 (N_1851,In_979,In_1125);
or U1852 (N_1852,In_1703,In_1874);
xor U1853 (N_1853,In_1704,In_1291);
xor U1854 (N_1854,In_699,In_1202);
nand U1855 (N_1855,In_300,In_1316);
nand U1856 (N_1856,In_239,In_1965);
or U1857 (N_1857,In_1090,In_1354);
and U1858 (N_1858,In_261,In_1871);
nand U1859 (N_1859,In_1245,In_1886);
nand U1860 (N_1860,In_503,In_625);
nand U1861 (N_1861,In_905,In_1214);
nor U1862 (N_1862,In_1127,In_1195);
or U1863 (N_1863,In_35,In_929);
or U1864 (N_1864,In_1015,In_1613);
nand U1865 (N_1865,In_1763,In_633);
and U1866 (N_1866,In_1055,In_1737);
or U1867 (N_1867,In_857,In_858);
and U1868 (N_1868,In_270,In_1013);
xnor U1869 (N_1869,In_676,In_1485);
xor U1870 (N_1870,In_989,In_706);
nand U1871 (N_1871,In_856,In_1515);
xnor U1872 (N_1872,In_1767,In_1441);
nand U1873 (N_1873,In_1268,In_1576);
and U1874 (N_1874,In_1238,In_346);
nor U1875 (N_1875,In_1221,In_1536);
nor U1876 (N_1876,In_1840,In_1587);
nor U1877 (N_1877,In_839,In_480);
xor U1878 (N_1878,In_474,In_1032);
and U1879 (N_1879,In_611,In_52);
and U1880 (N_1880,In_1184,In_231);
and U1881 (N_1881,In_1240,In_228);
nor U1882 (N_1882,In_372,In_647);
or U1883 (N_1883,In_845,In_660);
and U1884 (N_1884,In_188,In_1013);
nand U1885 (N_1885,In_127,In_1489);
and U1886 (N_1886,In_1933,In_1186);
nor U1887 (N_1887,In_1422,In_1853);
nor U1888 (N_1888,In_1779,In_1506);
xnor U1889 (N_1889,In_32,In_129);
and U1890 (N_1890,In_933,In_305);
nor U1891 (N_1891,In_1960,In_1916);
xor U1892 (N_1892,In_588,In_597);
nand U1893 (N_1893,In_1256,In_1268);
and U1894 (N_1894,In_1646,In_570);
or U1895 (N_1895,In_1266,In_116);
xor U1896 (N_1896,In_1192,In_1607);
nand U1897 (N_1897,In_1853,In_331);
and U1898 (N_1898,In_360,In_25);
or U1899 (N_1899,In_1444,In_623);
or U1900 (N_1900,In_1876,In_1219);
or U1901 (N_1901,In_530,In_254);
nor U1902 (N_1902,In_1858,In_569);
xor U1903 (N_1903,In_1529,In_692);
nor U1904 (N_1904,In_1798,In_166);
and U1905 (N_1905,In_726,In_836);
and U1906 (N_1906,In_715,In_1364);
or U1907 (N_1907,In_1025,In_1471);
xor U1908 (N_1908,In_1262,In_1742);
nor U1909 (N_1909,In_224,In_821);
or U1910 (N_1910,In_1370,In_835);
or U1911 (N_1911,In_1354,In_1981);
nor U1912 (N_1912,In_140,In_1576);
or U1913 (N_1913,In_1659,In_1453);
nor U1914 (N_1914,In_103,In_1467);
nand U1915 (N_1915,In_430,In_1580);
nand U1916 (N_1916,In_131,In_130);
nand U1917 (N_1917,In_1218,In_651);
xnor U1918 (N_1918,In_1216,In_1672);
nand U1919 (N_1919,In_624,In_829);
nor U1920 (N_1920,In_1608,In_835);
nor U1921 (N_1921,In_314,In_1385);
xor U1922 (N_1922,In_1779,In_827);
or U1923 (N_1923,In_525,In_1644);
or U1924 (N_1924,In_478,In_1924);
nand U1925 (N_1925,In_790,In_1793);
nand U1926 (N_1926,In_367,In_1181);
nand U1927 (N_1927,In_197,In_561);
and U1928 (N_1928,In_409,In_52);
xnor U1929 (N_1929,In_1778,In_1529);
and U1930 (N_1930,In_1318,In_1580);
nand U1931 (N_1931,In_1361,In_1675);
nor U1932 (N_1932,In_1031,In_1786);
nand U1933 (N_1933,In_4,In_885);
nand U1934 (N_1934,In_144,In_1961);
nand U1935 (N_1935,In_411,In_258);
or U1936 (N_1936,In_1597,In_1038);
nand U1937 (N_1937,In_910,In_457);
xor U1938 (N_1938,In_1775,In_1615);
or U1939 (N_1939,In_933,In_753);
or U1940 (N_1940,In_1555,In_611);
nor U1941 (N_1941,In_1352,In_1978);
and U1942 (N_1942,In_1790,In_1253);
and U1943 (N_1943,In_1823,In_419);
nor U1944 (N_1944,In_1274,In_920);
or U1945 (N_1945,In_514,In_886);
and U1946 (N_1946,In_1517,In_1577);
and U1947 (N_1947,In_511,In_972);
nor U1948 (N_1948,In_762,In_72);
nand U1949 (N_1949,In_1,In_1717);
or U1950 (N_1950,In_758,In_1059);
xnor U1951 (N_1951,In_393,In_144);
or U1952 (N_1952,In_1956,In_1709);
xor U1953 (N_1953,In_727,In_910);
and U1954 (N_1954,In_1068,In_1794);
nand U1955 (N_1955,In_757,In_543);
nand U1956 (N_1956,In_252,In_600);
and U1957 (N_1957,In_257,In_1081);
nand U1958 (N_1958,In_881,In_680);
and U1959 (N_1959,In_61,In_1291);
xnor U1960 (N_1960,In_1097,In_124);
nor U1961 (N_1961,In_873,In_884);
or U1962 (N_1962,In_1617,In_1141);
xnor U1963 (N_1963,In_776,In_793);
or U1964 (N_1964,In_1488,In_1968);
and U1965 (N_1965,In_2,In_1226);
xor U1966 (N_1966,In_1996,In_36);
nand U1967 (N_1967,In_689,In_194);
nor U1968 (N_1968,In_745,In_818);
nor U1969 (N_1969,In_515,In_248);
xor U1970 (N_1970,In_1437,In_1176);
and U1971 (N_1971,In_1239,In_722);
nor U1972 (N_1972,In_1199,In_873);
nand U1973 (N_1973,In_218,In_1635);
xor U1974 (N_1974,In_1405,In_1900);
nor U1975 (N_1975,In_1081,In_1533);
nand U1976 (N_1976,In_452,In_537);
or U1977 (N_1977,In_1380,In_568);
and U1978 (N_1978,In_1260,In_600);
nand U1979 (N_1979,In_1911,In_556);
and U1980 (N_1980,In_1911,In_1638);
xor U1981 (N_1981,In_178,In_592);
and U1982 (N_1982,In_540,In_1385);
nor U1983 (N_1983,In_356,In_267);
nor U1984 (N_1984,In_371,In_1242);
and U1985 (N_1985,In_408,In_1748);
and U1986 (N_1986,In_1933,In_768);
and U1987 (N_1987,In_1859,In_48);
or U1988 (N_1988,In_1636,In_1604);
nand U1989 (N_1989,In_986,In_1948);
and U1990 (N_1990,In_210,In_1731);
or U1991 (N_1991,In_112,In_1640);
nor U1992 (N_1992,In_1530,In_1840);
nor U1993 (N_1993,In_584,In_1168);
xor U1994 (N_1994,In_926,In_760);
and U1995 (N_1995,In_1147,In_1827);
and U1996 (N_1996,In_1372,In_1477);
and U1997 (N_1997,In_629,In_981);
nand U1998 (N_1998,In_1518,In_834);
or U1999 (N_1999,In_1240,In_43);
and U2000 (N_2000,N_1375,N_784);
xnor U2001 (N_2001,N_1385,N_771);
and U2002 (N_2002,N_305,N_1427);
nor U2003 (N_2003,N_1770,N_587);
and U2004 (N_2004,N_665,N_173);
and U2005 (N_2005,N_812,N_154);
nand U2006 (N_2006,N_1328,N_809);
xor U2007 (N_2007,N_75,N_1123);
nand U2008 (N_2008,N_519,N_589);
or U2009 (N_2009,N_8,N_1825);
or U2010 (N_2010,N_1312,N_1521);
nor U2011 (N_2011,N_1641,N_398);
or U2012 (N_2012,N_1971,N_1449);
xor U2013 (N_2013,N_593,N_1239);
nand U2014 (N_2014,N_1764,N_554);
and U2015 (N_2015,N_1757,N_640);
or U2016 (N_2016,N_931,N_1601);
and U2017 (N_2017,N_741,N_1915);
nor U2018 (N_2018,N_261,N_52);
or U2019 (N_2019,N_123,N_130);
and U2020 (N_2020,N_227,N_1369);
or U2021 (N_2021,N_377,N_543);
and U2022 (N_2022,N_460,N_1811);
and U2023 (N_2023,N_1076,N_687);
xor U2024 (N_2024,N_110,N_1908);
nor U2025 (N_2025,N_335,N_387);
or U2026 (N_2026,N_140,N_356);
or U2027 (N_2027,N_758,N_147);
nand U2028 (N_2028,N_1588,N_953);
or U2029 (N_2029,N_228,N_645);
nor U2030 (N_2030,N_603,N_834);
nand U2031 (N_2031,N_521,N_1736);
or U2032 (N_2032,N_1137,N_347);
nor U2033 (N_2033,N_1791,N_1384);
nor U2034 (N_2034,N_93,N_752);
nand U2035 (N_2035,N_290,N_513);
or U2036 (N_2036,N_1713,N_1780);
and U2037 (N_2037,N_1429,N_1102);
nor U2038 (N_2038,N_1262,N_82);
xor U2039 (N_2039,N_1554,N_442);
nand U2040 (N_2040,N_349,N_1927);
or U2041 (N_2041,N_1665,N_1687);
nand U2042 (N_2042,N_159,N_1335);
and U2043 (N_2043,N_1869,N_1999);
and U2044 (N_2044,N_459,N_606);
nor U2045 (N_2045,N_479,N_391);
nor U2046 (N_2046,N_974,N_57);
nor U2047 (N_2047,N_815,N_876);
nand U2048 (N_2048,N_1838,N_1723);
nor U2049 (N_2049,N_400,N_1865);
or U2050 (N_2050,N_1710,N_1593);
and U2051 (N_2051,N_1515,N_1980);
nand U2052 (N_2052,N_987,N_1500);
nor U2053 (N_2053,N_1381,N_572);
and U2054 (N_2054,N_1930,N_449);
nor U2055 (N_2055,N_1896,N_539);
and U2056 (N_2056,N_1724,N_916);
nand U2057 (N_2057,N_635,N_1735);
and U2058 (N_2058,N_1118,N_1095);
nand U2059 (N_2059,N_1964,N_1975);
nor U2060 (N_2060,N_191,N_471);
nand U2061 (N_2061,N_316,N_33);
xnor U2062 (N_2062,N_1826,N_1091);
and U2063 (N_2063,N_438,N_1018);
nand U2064 (N_2064,N_1252,N_65);
or U2065 (N_2065,N_1144,N_1456);
or U2066 (N_2066,N_1561,N_1491);
or U2067 (N_2067,N_47,N_1032);
nand U2068 (N_2068,N_1111,N_1657);
nor U2069 (N_2069,N_91,N_1510);
nand U2070 (N_2070,N_1910,N_1829);
or U2071 (N_2071,N_1273,N_1175);
or U2072 (N_2072,N_1062,N_503);
nor U2073 (N_2073,N_1636,N_1148);
nor U2074 (N_2074,N_181,N_662);
and U2075 (N_2075,N_1519,N_1858);
nor U2076 (N_2076,N_804,N_1619);
nor U2077 (N_2077,N_1991,N_41);
and U2078 (N_2078,N_249,N_745);
or U2079 (N_2079,N_274,N_168);
nor U2080 (N_2080,N_1093,N_1288);
nand U2081 (N_2081,N_294,N_1221);
nor U2082 (N_2082,N_884,N_67);
nor U2083 (N_2083,N_1926,N_1642);
or U2084 (N_2084,N_1524,N_1250);
nor U2085 (N_2085,N_1983,N_433);
and U2086 (N_2086,N_1185,N_233);
xnor U2087 (N_2087,N_1891,N_1286);
nand U2088 (N_2088,N_1443,N_1329);
and U2089 (N_2089,N_1040,N_737);
nor U2090 (N_2090,N_1614,N_145);
xnor U2091 (N_2091,N_898,N_894);
nor U2092 (N_2092,N_1270,N_11);
and U2093 (N_2093,N_1506,N_1985);
and U2094 (N_2094,N_610,N_166);
nor U2095 (N_2095,N_20,N_1338);
nor U2096 (N_2096,N_1631,N_1726);
nor U2097 (N_2097,N_772,N_1245);
nor U2098 (N_2098,N_724,N_1127);
nor U2099 (N_2099,N_155,N_1790);
or U2100 (N_2100,N_1750,N_1281);
or U2101 (N_2101,N_1502,N_1809);
nand U2102 (N_2102,N_1008,N_1581);
nor U2103 (N_2103,N_889,N_648);
and U2104 (N_2104,N_1741,N_1669);
xor U2105 (N_2105,N_656,N_1993);
nor U2106 (N_2106,N_461,N_1277);
nand U2107 (N_2107,N_259,N_415);
nand U2108 (N_2108,N_1552,N_1438);
and U2109 (N_2109,N_681,N_55);
or U2110 (N_2110,N_1104,N_1330);
and U2111 (N_2111,N_1121,N_597);
nor U2112 (N_2112,N_1487,N_310);
xor U2113 (N_2113,N_1844,N_77);
and U2114 (N_2114,N_473,N_683);
nand U2115 (N_2115,N_1535,N_295);
or U2116 (N_2116,N_1856,N_961);
nand U2117 (N_2117,N_1906,N_407);
and U2118 (N_2118,N_993,N_991);
nand U2119 (N_2119,N_776,N_1157);
nor U2120 (N_2120,N_1422,N_385);
or U2121 (N_2121,N_389,N_736);
xnor U2122 (N_2122,N_1399,N_523);
nor U2123 (N_2123,N_1358,N_1846);
nor U2124 (N_2124,N_1916,N_4);
nor U2125 (N_2125,N_1212,N_928);
or U2126 (N_2126,N_465,N_141);
or U2127 (N_2127,N_202,N_1476);
xor U2128 (N_2128,N_907,N_1717);
nor U2129 (N_2129,N_396,N_1845);
or U2130 (N_2130,N_618,N_1799);
xnor U2131 (N_2131,N_918,N_1587);
xor U2132 (N_2132,N_851,N_688);
or U2133 (N_2133,N_734,N_900);
nand U2134 (N_2134,N_1230,N_844);
nor U2135 (N_2135,N_122,N_557);
nor U2136 (N_2136,N_942,N_1536);
or U2137 (N_2137,N_873,N_210);
and U2138 (N_2138,N_667,N_1629);
nand U2139 (N_2139,N_1851,N_1932);
nor U2140 (N_2140,N_986,N_569);
nand U2141 (N_2141,N_790,N_594);
or U2142 (N_2142,N_158,N_138);
or U2143 (N_2143,N_1646,N_263);
nand U2144 (N_2144,N_518,N_1405);
nand U2145 (N_2145,N_1900,N_1549);
nand U2146 (N_2146,N_395,N_788);
nor U2147 (N_2147,N_26,N_1334);
and U2148 (N_2148,N_196,N_1508);
nor U2149 (N_2149,N_532,N_53);
nor U2150 (N_2150,N_964,N_200);
and U2151 (N_2151,N_880,N_1407);
and U2152 (N_2152,N_1672,N_397);
nand U2153 (N_2153,N_291,N_1017);
xor U2154 (N_2154,N_1603,N_983);
and U2155 (N_2155,N_810,N_1444);
nand U2156 (N_2156,N_1808,N_329);
or U2157 (N_2157,N_364,N_805);
nand U2158 (N_2158,N_56,N_800);
or U2159 (N_2159,N_1228,N_453);
nor U2160 (N_2160,N_496,N_285);
nor U2161 (N_2161,N_527,N_522);
xnor U2162 (N_2162,N_652,N_1086);
and U2163 (N_2163,N_843,N_595);
nand U2164 (N_2164,N_615,N_1386);
xor U2165 (N_2165,N_565,N_1831);
nand U2166 (N_2166,N_1174,N_949);
or U2167 (N_2167,N_1748,N_466);
and U2168 (N_2168,N_118,N_607);
nor U2169 (N_2169,N_1161,N_598);
nand U2170 (N_2170,N_1275,N_375);
and U2171 (N_2171,N_542,N_962);
and U2172 (N_2172,N_1348,N_1389);
nor U2173 (N_2173,N_629,N_1244);
or U2174 (N_2174,N_1539,N_333);
and U2175 (N_2175,N_336,N_1364);
or U2176 (N_2176,N_1708,N_1917);
xor U2177 (N_2177,N_432,N_634);
nor U2178 (N_2178,N_1716,N_1243);
or U2179 (N_2179,N_1821,N_1701);
nor U2180 (N_2180,N_911,N_1209);
nor U2181 (N_2181,N_1292,N_198);
xor U2182 (N_2182,N_677,N_1874);
nor U2183 (N_2183,N_1378,N_1314);
xnor U2184 (N_2184,N_18,N_1484);
and U2185 (N_2185,N_1450,N_863);
or U2186 (N_2186,N_1256,N_296);
nand U2187 (N_2187,N_1632,N_221);
or U2188 (N_2188,N_1024,N_478);
or U2189 (N_2189,N_908,N_897);
nor U2190 (N_2190,N_624,N_1699);
nor U2191 (N_2191,N_596,N_1666);
and U2192 (N_2192,N_1652,N_709);
or U2193 (N_2193,N_1152,N_865);
or U2194 (N_2194,N_502,N_692);
xor U2195 (N_2195,N_630,N_1238);
or U2196 (N_2196,N_787,N_1959);
nand U2197 (N_2197,N_1929,N_919);
nand U2198 (N_2198,N_1546,N_691);
and U2199 (N_2199,N_1316,N_1351);
and U2200 (N_2200,N_501,N_1379);
nor U2201 (N_2201,N_1711,N_1986);
or U2202 (N_2202,N_822,N_1191);
and U2203 (N_2203,N_457,N_701);
or U2204 (N_2204,N_94,N_1235);
nand U2205 (N_2205,N_269,N_765);
and U2206 (N_2206,N_9,N_353);
nand U2207 (N_2207,N_313,N_1637);
nor U2208 (N_2208,N_1160,N_1576);
or U2209 (N_2209,N_1278,N_1000);
xnor U2210 (N_2210,N_1297,N_1531);
nand U2211 (N_2211,N_664,N_975);
nor U2212 (N_2212,N_1530,N_488);
xor U2213 (N_2213,N_1099,N_1015);
nor U2214 (N_2214,N_782,N_872);
xor U2215 (N_2215,N_1876,N_1937);
or U2216 (N_2216,N_184,N_675);
and U2217 (N_2217,N_1967,N_1163);
nand U2218 (N_2218,N_1733,N_1568);
nand U2219 (N_2219,N_1555,N_320);
and U2220 (N_2220,N_831,N_412);
nor U2221 (N_2221,N_1225,N_1763);
or U2222 (N_2222,N_899,N_284);
and U2223 (N_2223,N_839,N_1463);
xor U2224 (N_2224,N_794,N_693);
and U2225 (N_2225,N_454,N_136);
and U2226 (N_2226,N_1433,N_1143);
or U2227 (N_2227,N_562,N_879);
or U2228 (N_2228,N_860,N_1624);
or U2229 (N_2229,N_644,N_1774);
nor U2230 (N_2230,N_1866,N_1849);
or U2231 (N_2231,N_372,N_495);
xor U2232 (N_2232,N_704,N_1756);
nand U2233 (N_2233,N_492,N_1553);
nor U2234 (N_2234,N_1705,N_1133);
nor U2235 (N_2235,N_1120,N_1534);
and U2236 (N_2236,N_1206,N_1754);
xor U2237 (N_2237,N_1216,N_1816);
and U2238 (N_2238,N_773,N_957);
nor U2239 (N_2239,N_1721,N_344);
or U2240 (N_2240,N_954,N_586);
nand U2241 (N_2241,N_278,N_1354);
nor U2242 (N_2242,N_1620,N_750);
nand U2243 (N_2243,N_514,N_1608);
nor U2244 (N_2244,N_475,N_1759);
nor U2245 (N_2245,N_1446,N_817);
nand U2246 (N_2246,N_1784,N_1651);
nor U2247 (N_2247,N_292,N_1173);
and U2248 (N_2248,N_1035,N_324);
nand U2249 (N_2249,N_1253,N_1883);
nor U2250 (N_2250,N_1300,N_161);
nand U2251 (N_2251,N_1343,N_832);
nor U2252 (N_2252,N_540,N_268);
or U2253 (N_2253,N_238,N_447);
and U2254 (N_2254,N_1566,N_666);
or U2255 (N_2255,N_1025,N_256);
nor U2256 (N_2256,N_307,N_700);
or U2257 (N_2257,N_1830,N_1394);
and U2258 (N_2258,N_1016,N_414);
nor U2259 (N_2259,N_747,N_1824);
or U2260 (N_2260,N_1541,N_711);
nor U2261 (N_2261,N_1383,N_1087);
nand U2262 (N_2262,N_760,N_64);
xor U2263 (N_2263,N_258,N_1810);
or U2264 (N_2264,N_1410,N_555);
nor U2265 (N_2265,N_1306,N_1019);
nor U2266 (N_2266,N_1049,N_558);
or U2267 (N_2267,N_152,N_1289);
nor U2268 (N_2268,N_647,N_545);
nand U2269 (N_2269,N_1951,N_1414);
nor U2270 (N_2270,N_1045,N_302);
nor U2271 (N_2271,N_1085,N_171);
or U2272 (N_2272,N_371,N_722);
and U2273 (N_2273,N_1889,N_455);
or U2274 (N_2274,N_1202,N_1526);
xnor U2275 (N_2275,N_637,N_505);
nor U2276 (N_2276,N_402,N_49);
or U2277 (N_2277,N_83,N_1890);
and U2278 (N_2278,N_1363,N_223);
nand U2279 (N_2279,N_1661,N_1565);
nor U2280 (N_2280,N_63,N_1979);
nand U2281 (N_2281,N_710,N_1728);
nor U2282 (N_2282,N_1935,N_1968);
nor U2283 (N_2283,N_759,N_1579);
or U2284 (N_2284,N_590,N_204);
nor U2285 (N_2285,N_833,N_720);
nand U2286 (N_2286,N_1153,N_823);
xnor U2287 (N_2287,N_570,N_535);
nor U2288 (N_2288,N_1956,N_1116);
or U2289 (N_2289,N_334,N_1972);
or U2290 (N_2290,N_1280,N_134);
nor U2291 (N_2291,N_1667,N_934);
or U2292 (N_2292,N_270,N_1346);
xor U2293 (N_2293,N_849,N_113);
or U2294 (N_2294,N_373,N_1633);
nor U2295 (N_2295,N_456,N_742);
or U2296 (N_2296,N_224,N_1392);
and U2297 (N_2297,N_62,N_1060);
and U2298 (N_2298,N_1324,N_1691);
xor U2299 (N_2299,N_1367,N_148);
and U2300 (N_2300,N_1279,N_1789);
nand U2301 (N_2301,N_1350,N_1695);
nor U2302 (N_2302,N_1893,N_1905);
and U2303 (N_2303,N_1490,N_1150);
nand U2304 (N_2304,N_1226,N_339);
and U2305 (N_2305,N_450,N_1697);
and U2306 (N_2306,N_1465,N_1848);
or U2307 (N_2307,N_1255,N_1479);
nand U2308 (N_2308,N_1029,N_671);
or U2309 (N_2309,N_1263,N_778);
and U2310 (N_2310,N_1042,N_1574);
nor U2311 (N_2311,N_1855,N_951);
nor U2312 (N_2312,N_408,N_1779);
or U2313 (N_2313,N_799,N_1483);
and U2314 (N_2314,N_1485,N_601);
nand U2315 (N_2315,N_28,N_1393);
nor U2316 (N_2316,N_1177,N_694);
and U2317 (N_2317,N_813,N_547);
nand U2318 (N_2318,N_1702,N_1416);
nand U2319 (N_2319,N_1237,N_0);
nor U2320 (N_2320,N_361,N_902);
nor U2321 (N_2321,N_1070,N_981);
and U2322 (N_2322,N_1658,N_128);
or U2323 (N_2323,N_904,N_1002);
nor U2324 (N_2324,N_374,N_167);
nor U2325 (N_2325,N_1220,N_685);
nor U2326 (N_2326,N_891,N_1408);
and U2327 (N_2327,N_1488,N_529);
xor U2328 (N_2328,N_1400,N_231);
nor U2329 (N_2329,N_1140,N_1992);
nor U2330 (N_2330,N_1822,N_571);
or U2331 (N_2331,N_1332,N_1545);
and U2332 (N_2332,N_1604,N_340);
nand U2333 (N_2333,N_729,N_733);
or U2334 (N_2334,N_926,N_852);
xnor U2335 (N_2335,N_1933,N_1704);
or U2336 (N_2336,N_1602,N_1006);
nand U2337 (N_2337,N_661,N_42);
nand U2338 (N_2338,N_553,N_506);
nor U2339 (N_2339,N_170,N_1788);
and U2340 (N_2340,N_1765,N_924);
nand U2341 (N_2341,N_1340,N_1327);
nand U2342 (N_2342,N_602,N_1184);
nor U2343 (N_2343,N_358,N_1714);
nor U2344 (N_2344,N_79,N_1172);
or U2345 (N_2345,N_537,N_1931);
nor U2346 (N_2346,N_1792,N_922);
nor U2347 (N_2347,N_703,N_1660);
nand U2348 (N_2348,N_1605,N_1164);
nor U2349 (N_2349,N_345,N_1974);
or U2350 (N_2350,N_1953,N_271);
nor U2351 (N_2351,N_1272,N_1492);
nand U2352 (N_2352,N_877,N_1211);
and U2353 (N_2353,N_842,N_1199);
nand U2354 (N_2354,N_1254,N_1635);
nor U2355 (N_2355,N_1195,N_573);
and U2356 (N_2356,N_668,N_578);
nand U2357 (N_2357,N_546,N_619);
nand U2358 (N_2358,N_1762,N_1204);
nor U2359 (N_2359,N_379,N_1513);
nand U2360 (N_2360,N_1639,N_1031);
nor U2361 (N_2361,N_1938,N_1613);
xnor U2362 (N_2362,N_1941,N_1377);
nor U2363 (N_2363,N_1880,N_1563);
and U2364 (N_2364,N_1946,N_489);
nor U2365 (N_2365,N_1274,N_243);
xnor U2366 (N_2366,N_753,N_72);
xor U2367 (N_2367,N_774,N_229);
xor U2368 (N_2368,N_251,N_1960);
nor U2369 (N_2369,N_699,N_1047);
and U2370 (N_2370,N_180,N_208);
nor U2371 (N_2371,N_376,N_218);
or U2372 (N_2372,N_575,N_1776);
or U2373 (N_2373,N_655,N_1740);
nor U2374 (N_2374,N_725,N_930);
nor U2375 (N_2375,N_549,N_1570);
or U2376 (N_2376,N_1615,N_1626);
or U2377 (N_2377,N_1727,N_197);
nor U2378 (N_2378,N_976,N_657);
or U2379 (N_2379,N_1976,N_840);
nor U2380 (N_2380,N_237,N_434);
and U2381 (N_2381,N_1606,N_1382);
xnor U2382 (N_2382,N_348,N_194);
nor U2383 (N_2383,N_1512,N_821);
nand U2384 (N_2384,N_1103,N_143);
xor U2385 (N_2385,N_1649,N_346);
xor U2386 (N_2386,N_568,N_1540);
nor U2387 (N_2387,N_1778,N_160);
nand U2388 (N_2388,N_1958,N_696);
and U2389 (N_2389,N_1344,N_1590);
nand U2390 (N_2390,N_989,N_1411);
and U2391 (N_2391,N_802,N_888);
nor U2392 (N_2392,N_267,N_1081);
nor U2393 (N_2393,N_1059,N_10);
and U2394 (N_2394,N_1061,N_1885);
nand U2395 (N_2395,N_1734,N_169);
or U2396 (N_2396,N_1662,N_1094);
or U2397 (N_2397,N_95,N_1374);
xor U2398 (N_2398,N_1739,N_906);
nand U2399 (N_2399,N_298,N_1168);
xnor U2400 (N_2400,N_798,N_861);
xnor U2401 (N_2401,N_70,N_1132);
or U2402 (N_2402,N_1954,N_853);
and U2403 (N_2403,N_552,N_1559);
nand U2404 (N_2404,N_621,N_1607);
and U2405 (N_2405,N_247,N_1260);
nor U2406 (N_2406,N_1621,N_507);
nor U2407 (N_2407,N_92,N_935);
nor U2408 (N_2408,N_1628,N_1773);
or U2409 (N_2409,N_674,N_201);
or U2410 (N_2410,N_1596,N_1921);
or U2411 (N_2411,N_1918,N_1547);
or U2412 (N_2412,N_1322,N_1371);
nand U2413 (N_2413,N_275,N_636);
nor U2414 (N_2414,N_1520,N_1007);
nand U2415 (N_2415,N_1949,N_1468);
nor U2416 (N_2416,N_1064,N_6);
nand U2417 (N_2417,N_528,N_207);
and U2418 (N_2418,N_1167,N_1793);
xnor U2419 (N_2419,N_628,N_971);
nor U2420 (N_2420,N_1692,N_429);
and U2421 (N_2421,N_614,N_137);
nand U2422 (N_2422,N_1850,N_164);
and U2423 (N_2423,N_1653,N_1257);
xor U2424 (N_2424,N_452,N_1224);
or U2425 (N_2425,N_585,N_1470);
or U2426 (N_2426,N_462,N_1564);
nor U2427 (N_2427,N_1413,N_1800);
nor U2428 (N_2428,N_90,N_574);
nand U2429 (N_2429,N_99,N_1843);
nor U2430 (N_2430,N_896,N_37);
nor U2431 (N_2431,N_1131,N_1112);
nand U2432 (N_2432,N_580,N_1317);
or U2433 (N_2433,N_287,N_1055);
or U2434 (N_2434,N_1857,N_1902);
or U2435 (N_2435,N_1899,N_255);
nand U2436 (N_2436,N_1482,N_1575);
nand U2437 (N_2437,N_1940,N_1920);
and U2438 (N_2438,N_723,N_1744);
nand U2439 (N_2439,N_544,N_641);
or U2440 (N_2440,N_1997,N_1690);
or U2441 (N_2441,N_317,N_119);
and U2442 (N_2442,N_1229,N_1904);
or U2443 (N_2443,N_1217,N_1580);
xor U2444 (N_2444,N_1437,N_941);
xnor U2445 (N_2445,N_244,N_1518);
nand U2446 (N_2446,N_1746,N_1677);
and U2447 (N_2447,N_477,N_1423);
or U2448 (N_2448,N_717,N_1542);
nand U2449 (N_2449,N_1768,N_150);
and U2450 (N_2450,N_959,N_117);
or U2451 (N_2451,N_40,N_1360);
or U2452 (N_2452,N_481,N_801);
and U2453 (N_2453,N_1796,N_715);
nor U2454 (N_2454,N_1988,N_1755);
and U2455 (N_2455,N_1560,N_1584);
nand U2456 (N_2456,N_1146,N_854);
and U2457 (N_2457,N_239,N_1957);
nor U2458 (N_2458,N_504,N_403);
nor U2459 (N_2459,N_1936,N_5);
nor U2460 (N_2460,N_1569,N_1315);
and U2461 (N_2461,N_1873,N_973);
nor U2462 (N_2462,N_281,N_404);
nor U2463 (N_2463,N_869,N_1514);
or U2464 (N_2464,N_866,N_1142);
and U2465 (N_2465,N_1503,N_1036);
and U2466 (N_2466,N_1511,N_943);
nand U2467 (N_2467,N_1355,N_885);
nand U2468 (N_2468,N_131,N_515);
or U2469 (N_2469,N_1170,N_222);
or U2470 (N_2470,N_1004,N_903);
or U2471 (N_2471,N_1022,N_1050);
and U2472 (N_2472,N_2,N_1135);
nand U2473 (N_2473,N_1871,N_1989);
or U2474 (N_2474,N_1777,N_1418);
nor U2475 (N_2475,N_175,N_847);
and U2476 (N_2476,N_1718,N_1679);
nor U2477 (N_2477,N_1537,N_410);
or U2478 (N_2478,N_757,N_945);
nor U2479 (N_2479,N_534,N_1339);
nand U2480 (N_2480,N_1139,N_1258);
nor U2481 (N_2481,N_678,N_526);
nor U2482 (N_2482,N_315,N_1285);
and U2483 (N_2483,N_669,N_848);
xnor U2484 (N_2484,N_1719,N_1165);
or U2485 (N_2485,N_613,N_1609);
nor U2486 (N_2486,N_818,N_1447);
and U2487 (N_2487,N_29,N_60);
xnor U2488 (N_2488,N_1373,N_1155);
or U2489 (N_2489,N_874,N_314);
or U2490 (N_2490,N_1078,N_48);
and U2491 (N_2491,N_351,N_1680);
nor U2492 (N_2492,N_424,N_1769);
or U2493 (N_2493,N_627,N_1246);
nor U2494 (N_2494,N_1558,N_413);
and U2495 (N_2495,N_474,N_102);
nor U2496 (N_2496,N_132,N_1147);
nor U2497 (N_2497,N_1516,N_516);
nand U2498 (N_2498,N_1939,N_359);
and U2499 (N_2499,N_209,N_469);
and U2500 (N_2500,N_1039,N_1234);
and U2501 (N_2501,N_135,N_1681);
nor U2502 (N_2502,N_446,N_493);
or U2503 (N_2503,N_486,N_1832);
and U2504 (N_2504,N_1010,N_14);
nor U2505 (N_2505,N_46,N_646);
or U2506 (N_2506,N_1156,N_588);
or U2507 (N_2507,N_726,N_1582);
nand U2508 (N_2508,N_1685,N_718);
and U2509 (N_2509,N_735,N_236);
nor U2510 (N_2510,N_789,N_388);
and U2511 (N_2511,N_933,N_895);
and U2512 (N_2512,N_1730,N_1391);
and U2513 (N_2513,N_841,N_406);
nor U2514 (N_2514,N_487,N_1303);
and U2515 (N_2515,N_435,N_791);
nand U2516 (N_2516,N_1337,N_875);
nor U2517 (N_2517,N_1145,N_702);
nor U2518 (N_2518,N_23,N_392);
nand U2519 (N_2519,N_1321,N_932);
nand U2520 (N_2520,N_1325,N_311);
or U2521 (N_2521,N_485,N_1638);
and U2522 (N_2522,N_368,N_103);
nor U2523 (N_2523,N_394,N_1464);
nor U2524 (N_2524,N_1761,N_25);
and U2525 (N_2525,N_61,N_1571);
nand U2526 (N_2526,N_226,N_1180);
xor U2527 (N_2527,N_520,N_1998);
or U2528 (N_2528,N_536,N_19);
or U2529 (N_2529,N_286,N_214);
or U2530 (N_2530,N_850,N_1806);
and U2531 (N_2531,N_689,N_921);
nand U2532 (N_2532,N_1406,N_13);
nor U2533 (N_2533,N_1480,N_253);
or U2534 (N_2534,N_1259,N_116);
nor U2535 (N_2535,N_441,N_524);
and U2536 (N_2536,N_1214,N_1436);
nor U2537 (N_2537,N_1640,N_1159);
and U2538 (N_2538,N_1151,N_1056);
xor U2539 (N_2539,N_1326,N_178);
nor U2540 (N_2540,N_464,N_44);
and U2541 (N_2541,N_582,N_1372);
nor U2542 (N_2542,N_80,N_1401);
nor U2543 (N_2543,N_1805,N_163);
or U2544 (N_2544,N_965,N_370);
nand U2545 (N_2545,N_497,N_1995);
or U2546 (N_2546,N_1293,N_7);
xnor U2547 (N_2547,N_1305,N_1807);
or U2548 (N_2548,N_837,N_38);
and U2549 (N_2549,N_272,N_511);
nor U2550 (N_2550,N_1737,N_1341);
nor U2551 (N_2551,N_999,N_86);
or U2552 (N_2552,N_106,N_1026);
or U2553 (N_2553,N_1556,N_139);
and U2554 (N_2554,N_1751,N_355);
or U2555 (N_2555,N_1189,N_381);
and U2556 (N_2556,N_16,N_862);
or U2557 (N_2557,N_779,N_620);
and U2558 (N_2558,N_1454,N_676);
and U2559 (N_2559,N_179,N_1474);
nor U2560 (N_2560,N_561,N_69);
and U2561 (N_2561,N_1489,N_1879);
or U2562 (N_2562,N_1493,N_1448);
or U2563 (N_2563,N_350,N_1271);
or U2564 (N_2564,N_1472,N_1694);
or U2565 (N_2565,N_1673,N_1361);
nand U2566 (N_2566,N_114,N_390);
nand U2567 (N_2567,N_1898,N_1466);
nand U2568 (N_2568,N_1706,N_1071);
nor U2569 (N_2569,N_1634,N_1440);
and U2570 (N_2570,N_1738,N_1981);
nor U2571 (N_2571,N_795,N_409);
nand U2572 (N_2572,N_984,N_1117);
or U2573 (N_2573,N_280,N_232);
and U2574 (N_2574,N_1567,N_35);
or U2575 (N_2575,N_323,N_27);
nand U2576 (N_2576,N_1894,N_1645);
nand U2577 (N_2577,N_1712,N_1075);
and U2578 (N_2578,N_1543,N_1693);
nand U2579 (N_2579,N_751,N_112);
nor U2580 (N_2580,N_230,N_909);
nor U2581 (N_2581,N_881,N_1441);
nand U2582 (N_2582,N_728,N_1925);
nand U2583 (N_2583,N_1365,N_767);
nor U2584 (N_2584,N_1668,N_380);
and U2585 (N_2585,N_1455,N_1298);
and U2586 (N_2586,N_868,N_1458);
or U2587 (N_2587,N_1884,N_354);
nand U2588 (N_2588,N_947,N_483);
xor U2589 (N_2589,N_1100,N_713);
and U2590 (N_2590,N_212,N_1471);
nand U2591 (N_2591,N_129,N_1409);
or U2592 (N_2592,N_439,N_1909);
or U2593 (N_2593,N_1241,N_1878);
nand U2594 (N_2594,N_1421,N_856);
xor U2595 (N_2595,N_1467,N_893);
or U2596 (N_2596,N_1388,N_1356);
nand U2597 (N_2597,N_855,N_1207);
nor U2598 (N_2598,N_680,N_814);
or U2599 (N_2599,N_1233,N_1417);
nand U2600 (N_2600,N_1477,N_777);
nand U2601 (N_2601,N_308,N_1052);
or U2602 (N_2602,N_257,N_857);
nor U2603 (N_2603,N_1965,N_416);
xor U2604 (N_2604,N_1218,N_225);
nor U2605 (N_2605,N_321,N_995);
or U2606 (N_2606,N_352,N_623);
nor U2607 (N_2607,N_1732,N_322);
nor U2608 (N_2608,N_592,N_886);
nor U2609 (N_2609,N_1430,N_51);
nor U2610 (N_2610,N_293,N_632);
nand U2611 (N_2611,N_1644,N_1785);
nor U2612 (N_2612,N_1190,N_1715);
nand U2613 (N_2613,N_451,N_1287);
nand U2614 (N_2614,N_743,N_1068);
or U2615 (N_2615,N_1027,N_1376);
and U2616 (N_2616,N_337,N_1767);
nor U2617 (N_2617,N_1296,N_1625);
nor U2618 (N_2618,N_531,N_420);
nor U2619 (N_2619,N_1459,N_499);
xnor U2620 (N_2620,N_1863,N_146);
nand U2621 (N_2621,N_806,N_1860);
nand U2622 (N_2622,N_1766,N_1063);
or U2623 (N_2623,N_1169,N_203);
nand U2624 (N_2624,N_1294,N_419);
and U2625 (N_2625,N_1758,N_1919);
and U2626 (N_2626,N_360,N_1439);
nor U2627 (N_2627,N_936,N_1698);
and U2628 (N_2628,N_1048,N_1188);
or U2629 (N_2629,N_1481,N_1067);
and U2630 (N_2630,N_1557,N_242);
xor U2631 (N_2631,N_276,N_331);
and U2632 (N_2632,N_1265,N_437);
and U2633 (N_2633,N_297,N_1034);
nand U2634 (N_2634,N_59,N_1962);
or U2635 (N_2635,N_405,N_1854);
or U2636 (N_2636,N_740,N_1775);
xnor U2637 (N_2637,N_183,N_125);
and U2638 (N_2638,N_1028,N_1700);
and U2639 (N_2639,N_1114,N_1397);
nor U2640 (N_2640,N_658,N_260);
or U2641 (N_2641,N_551,N_399);
nor U2642 (N_2642,N_188,N_1887);
and U2643 (N_2643,N_1181,N_98);
nor U2644 (N_2644,N_912,N_1141);
and U2645 (N_2645,N_1309,N_1676);
and U2646 (N_2646,N_384,N_783);
xnor U2647 (N_2647,N_1720,N_1053);
and U2648 (N_2648,N_1729,N_650);
nand U2649 (N_2649,N_1435,N_512);
and U2650 (N_2650,N_1772,N_1345);
or U2651 (N_2651,N_1752,N_748);
nand U2652 (N_2652,N_966,N_1310);
nand U2653 (N_2653,N_1504,N_328);
nor U2654 (N_2654,N_950,N_211);
nor U2655 (N_2655,N_187,N_1618);
nand U2656 (N_2656,N_124,N_859);
nor U2657 (N_2657,N_576,N_1186);
or U2658 (N_2658,N_567,N_1072);
nand U2659 (N_2659,N_1201,N_192);
and U2660 (N_2660,N_566,N_144);
and U2661 (N_2661,N_32,N_1840);
nand U2662 (N_2662,N_1213,N_690);
or U2663 (N_2663,N_510,N_948);
nand U2664 (N_2664,N_638,N_914);
or U2665 (N_2665,N_963,N_538);
or U2666 (N_2666,N_1158,N_1901);
and U2667 (N_2667,N_617,N_417);
or U2668 (N_2668,N_901,N_556);
nand U2669 (N_2669,N_1955,N_682);
nand U2670 (N_2670,N_1507,N_1771);
or U2671 (N_2671,N_81,N_1194);
nand U2672 (N_2672,N_463,N_927);
or U2673 (N_2673,N_1689,N_443);
xor U2674 (N_2674,N_1859,N_1794);
nor U2675 (N_2675,N_1913,N_611);
nand U2676 (N_2676,N_679,N_1731);
nor U2677 (N_2677,N_304,N_583);
and U2678 (N_2678,N_915,N_738);
nand U2679 (N_2679,N_1837,N_1795);
or U2680 (N_2680,N_1462,N_66);
and U2681 (N_2681,N_105,N_1130);
nor U2682 (N_2682,N_706,N_708);
nand U2683 (N_2683,N_796,N_1445);
and U2684 (N_2684,N_1815,N_1380);
or U2685 (N_2685,N_1627,N_480);
or U2686 (N_2686,N_1119,N_245);
nor U2687 (N_2687,N_1357,N_445);
xnor U2688 (N_2688,N_824,N_1183);
and U2689 (N_2689,N_58,N_1074);
and U2690 (N_2690,N_829,N_1599);
xnor U2691 (N_2691,N_1179,N_1115);
xor U2692 (N_2692,N_1509,N_264);
or U2693 (N_2693,N_1083,N_185);
xor U2694 (N_2694,N_104,N_1187);
nor U2695 (N_2695,N_248,N_1595);
or U2696 (N_2696,N_1077,N_246);
and U2697 (N_2697,N_517,N_1562);
or U2698 (N_2698,N_1154,N_1012);
nand U2699 (N_2699,N_1743,N_330);
nand U2700 (N_2700,N_21,N_1451);
or U2701 (N_2701,N_362,N_1760);
or U2702 (N_2702,N_1236,N_811);
nor U2703 (N_2703,N_1573,N_1005);
xor U2704 (N_2704,N_719,N_1578);
nor U2705 (N_2705,N_108,N_530);
xnor U2706 (N_2706,N_659,N_892);
and U2707 (N_2707,N_54,N_913);
or U2708 (N_2708,N_686,N_1592);
and U2709 (N_2709,N_612,N_599);
nand U2710 (N_2710,N_867,N_1109);
nand U2711 (N_2711,N_176,N_1193);
and U2712 (N_2712,N_1819,N_1420);
xor U2713 (N_2713,N_367,N_1030);
and U2714 (N_2714,N_428,N_127);
and U2715 (N_2715,N_1457,N_548);
or U2716 (N_2716,N_808,N_653);
and U2717 (N_2717,N_830,N_509);
or U2718 (N_2718,N_1432,N_1311);
and U2719 (N_2719,N_467,N_846);
or U2720 (N_2720,N_1359,N_978);
nand U2721 (N_2721,N_43,N_712);
and U2722 (N_2722,N_153,N_1912);
nand U2723 (N_2723,N_482,N_1362);
nor U2724 (N_2724,N_970,N_1970);
nor U2725 (N_2725,N_1046,N_672);
or U2726 (N_2726,N_1611,N_1396);
xor U2727 (N_2727,N_1208,N_217);
nand U2728 (N_2728,N_1090,N_946);
xor U2729 (N_2729,N_157,N_1963);
xnor U2730 (N_2730,N_1533,N_1058);
and U2731 (N_2731,N_22,N_206);
nand U2732 (N_2732,N_1428,N_1996);
xor U2733 (N_2733,N_174,N_643);
nand U2734 (N_2734,N_1594,N_649);
nor U2735 (N_2735,N_1499,N_215);
nor U2736 (N_2736,N_97,N_797);
nand U2737 (N_2737,N_177,N_235);
nand U2738 (N_2738,N_827,N_1544);
nor U2739 (N_2739,N_299,N_1261);
nor U2740 (N_2740,N_1833,N_938);
and U2741 (N_2741,N_755,N_541);
or U2742 (N_2742,N_559,N_1223);
xnor U2743 (N_2743,N_332,N_835);
nand U2744 (N_2744,N_1215,N_1065);
and U2745 (N_2745,N_418,N_1888);
xor U2746 (N_2746,N_1041,N_992);
nand U2747 (N_2747,N_1950,N_282);
or U2748 (N_2748,N_1787,N_250);
nor U2749 (N_2749,N_1283,N_622);
or U2750 (N_2750,N_1425,N_972);
or U2751 (N_2751,N_1643,N_1478);
and U2752 (N_2752,N_1136,N_45);
and U2753 (N_2753,N_920,N_807);
nor U2754 (N_2754,N_980,N_220);
and U2755 (N_2755,N_71,N_1945);
nor U2756 (N_2756,N_1276,N_195);
or U2757 (N_2757,N_1978,N_917);
or U2758 (N_2758,N_50,N_1589);
xnor U2759 (N_2759,N_1897,N_1654);
or U2760 (N_2760,N_1347,N_1101);
and U2761 (N_2761,N_24,N_1517);
nand U2762 (N_2762,N_1106,N_1934);
nor U2763 (N_2763,N_89,N_979);
nand U2764 (N_2764,N_864,N_363);
or U2765 (N_2765,N_982,N_1129);
nand U2766 (N_2766,N_1610,N_306);
nand U2767 (N_2767,N_939,N_1781);
nor U2768 (N_2768,N_944,N_1267);
nand U2769 (N_2769,N_1044,N_1387);
nand U2770 (N_2770,N_775,N_1798);
nand U2771 (N_2771,N_378,N_1994);
xor U2772 (N_2772,N_591,N_111);
or U2773 (N_2773,N_1688,N_1803);
nor U2774 (N_2774,N_716,N_1403);
and U2775 (N_2775,N_883,N_1847);
xor U2776 (N_2776,N_770,N_107);
nor U2777 (N_2777,N_357,N_1162);
or U2778 (N_2778,N_266,N_985);
nor U2779 (N_2779,N_1370,N_1987);
and U2780 (N_2780,N_186,N_393);
nor U2781 (N_2781,N_695,N_1349);
nand U2782 (N_2782,N_820,N_1525);
xor U2783 (N_2783,N_470,N_732);
nand U2784 (N_2784,N_88,N_1841);
or U2785 (N_2785,N_1961,N_910);
xnor U2786 (N_2786,N_1522,N_1037);
and U2787 (N_2787,N_730,N_560);
nand U2788 (N_2788,N_1947,N_1648);
nand U2789 (N_2789,N_342,N_1222);
or U2790 (N_2790,N_1247,N_1814);
and U2791 (N_2791,N_1886,N_1802);
nor U2792 (N_2792,N_1424,N_1054);
and U2793 (N_2793,N_1113,N_1749);
and U2794 (N_2794,N_289,N_1703);
nand U2795 (N_2795,N_468,N_609);
nand U2796 (N_2796,N_1529,N_1089);
nor U2797 (N_2797,N_115,N_1431);
nor U2798 (N_2798,N_426,N_766);
nand U2799 (N_2799,N_288,N_968);
and U2800 (N_2800,N_923,N_1862);
nand U2801 (N_2801,N_698,N_382);
and U2802 (N_2802,N_1630,N_1290);
nor U2803 (N_2803,N_967,N_1460);
nor U2804 (N_2804,N_1079,N_1586);
xnor U2805 (N_2805,N_1663,N_1682);
or U2806 (N_2806,N_1197,N_785);
nor U2807 (N_2807,N_1674,N_1683);
or U2808 (N_2808,N_193,N_1914);
or U2809 (N_2809,N_411,N_1817);
nand U2810 (N_2810,N_1496,N_484);
xor U2811 (N_2811,N_608,N_1943);
or U2812 (N_2812,N_714,N_1583);
and U2813 (N_2813,N_1323,N_793);
or U2814 (N_2814,N_977,N_120);
nand U2815 (N_2815,N_1684,N_1084);
nor U2816 (N_2816,N_325,N_670);
nor U2817 (N_2817,N_925,N_216);
and U2818 (N_2818,N_1291,N_254);
and U2819 (N_2819,N_1742,N_616);
xor U2820 (N_2820,N_1171,N_1196);
xor U2821 (N_2821,N_1538,N_819);
nand U2822 (N_2822,N_444,N_564);
and U2823 (N_2823,N_673,N_952);
nor U2824 (N_2824,N_448,N_780);
and U2825 (N_2825,N_754,N_1051);
xor U2826 (N_2826,N_151,N_427);
and U2827 (N_2827,N_162,N_1009);
nand U2828 (N_2828,N_165,N_663);
or U2829 (N_2829,N_1178,N_1532);
nand U2830 (N_2830,N_890,N_988);
and U2831 (N_2831,N_1232,N_301);
and U2832 (N_2832,N_1836,N_1722);
nand U2833 (N_2833,N_1203,N_142);
nand U2834 (N_2834,N_84,N_252);
nand U2835 (N_2835,N_1523,N_326);
xor U2836 (N_2836,N_584,N_277);
or U2837 (N_2837,N_1675,N_969);
and U2838 (N_2838,N_436,N_1585);
or U2839 (N_2839,N_219,N_838);
nor U2840 (N_2840,N_273,N_1892);
and U2841 (N_2841,N_600,N_1319);
and U2842 (N_2842,N_1498,N_1527);
nor U2843 (N_2843,N_1080,N_929);
or U2844 (N_2844,N_764,N_1868);
nor U2845 (N_2845,N_1395,N_882);
nand U2846 (N_2846,N_1877,N_1753);
and U2847 (N_2847,N_1597,N_1038);
xnor U2848 (N_2848,N_1200,N_1419);
xnor U2849 (N_2849,N_605,N_1797);
nand U2850 (N_2850,N_1043,N_660);
nand U2851 (N_2851,N_430,N_1872);
nor U2852 (N_2852,N_642,N_490);
nor U2853 (N_2853,N_1864,N_1745);
or U2854 (N_2854,N_1528,N_845);
nand U2855 (N_2855,N_1616,N_1366);
nor U2856 (N_2856,N_1249,N_1475);
nand U2857 (N_2857,N_1783,N_1108);
nand U2858 (N_2858,N_1813,N_1696);
nor U2859 (N_2859,N_78,N_1390);
or U2860 (N_2860,N_1828,N_1551);
and U2861 (N_2861,N_189,N_96);
or U2862 (N_2862,N_826,N_756);
nand U2863 (N_2863,N_631,N_401);
nor U2864 (N_2864,N_1942,N_816);
and U2865 (N_2865,N_579,N_312);
nor U2866 (N_2866,N_262,N_1623);
nor U2867 (N_2867,N_30,N_727);
nand U2868 (N_2868,N_234,N_1827);
nand U2869 (N_2869,N_172,N_1227);
and U2870 (N_2870,N_1928,N_768);
nor U2871 (N_2871,N_1747,N_563);
and U2872 (N_2872,N_749,N_1823);
nor U2873 (N_2873,N_1977,N_85);
xor U2874 (N_2874,N_383,N_1404);
nor U2875 (N_2875,N_625,N_1577);
xor U2876 (N_2876,N_1098,N_1066);
nand U2877 (N_2877,N_1318,N_300);
and U2878 (N_2878,N_15,N_1057);
xor U2879 (N_2879,N_955,N_149);
xor U2880 (N_2880,N_707,N_1505);
or U2881 (N_2881,N_1122,N_68);
nand U2882 (N_2882,N_423,N_1801);
nor U2883 (N_2883,N_990,N_533);
nand U2884 (N_2884,N_1834,N_1707);
and U2885 (N_2885,N_1368,N_878);
nor U2886 (N_2886,N_940,N_1219);
or U2887 (N_2887,N_1591,N_1990);
nor U2888 (N_2888,N_956,N_1033);
nor U2889 (N_2889,N_1282,N_1242);
nor U2890 (N_2890,N_121,N_525);
nand U2891 (N_2891,N_905,N_550);
or U2892 (N_2892,N_1023,N_1138);
xor U2893 (N_2893,N_1073,N_997);
nand U2894 (N_2894,N_109,N_1495);
nor U2895 (N_2895,N_1001,N_998);
and U2896 (N_2896,N_365,N_309);
nor U2897 (N_2897,N_639,N_1069);
nand U2898 (N_2898,N_182,N_1011);
or U2899 (N_2899,N_1852,N_1875);
xor U2900 (N_2900,N_1125,N_870);
xnor U2901 (N_2901,N_1982,N_1336);
nor U2902 (N_2902,N_836,N_1969);
nor U2903 (N_2903,N_761,N_199);
nand U2904 (N_2904,N_1304,N_1818);
xor U2905 (N_2905,N_626,N_343);
or U2906 (N_2906,N_1835,N_1205);
or U2907 (N_2907,N_762,N_476);
or U2908 (N_2908,N_828,N_431);
nand U2909 (N_2909,N_1198,N_1434);
nand U2910 (N_2910,N_1686,N_1881);
and U2911 (N_2911,N_1550,N_769);
and U2912 (N_2912,N_1097,N_803);
xnor U2913 (N_2913,N_1415,N_1812);
and U2914 (N_2914,N_421,N_386);
or U2915 (N_2915,N_279,N_156);
nor U2916 (N_2916,N_126,N_1678);
and U2917 (N_2917,N_1308,N_73);
nand U2918 (N_2918,N_500,N_1333);
nor U2919 (N_2919,N_1944,N_1182);
xnor U2920 (N_2920,N_1839,N_1398);
and U2921 (N_2921,N_786,N_498);
nor U2922 (N_2922,N_36,N_731);
nand U2923 (N_2923,N_3,N_1295);
nand U2924 (N_2924,N_746,N_1313);
nand U2925 (N_2925,N_1647,N_1870);
nor U2926 (N_2926,N_213,N_491);
nand U2927 (N_2927,N_577,N_1659);
nor U2928 (N_2928,N_1617,N_1984);
or U2929 (N_2929,N_581,N_366);
or U2930 (N_2930,N_338,N_1461);
and U2931 (N_2931,N_1664,N_472);
nand U2932 (N_2932,N_303,N_1867);
or U2933 (N_2933,N_1709,N_1782);
and U2934 (N_2934,N_369,N_1082);
nor U2935 (N_2935,N_1911,N_283);
nor U2936 (N_2936,N_1670,N_1331);
and U2937 (N_2937,N_1486,N_240);
nand U2938 (N_2938,N_1124,N_858);
nand U2939 (N_2939,N_1342,N_1107);
or U2940 (N_2940,N_1240,N_1264);
nor U2941 (N_2941,N_721,N_422);
nor U2942 (N_2942,N_1952,N_1842);
or U2943 (N_2943,N_1882,N_318);
nand U2944 (N_2944,N_1973,N_604);
or U2945 (N_2945,N_887,N_705);
or U2946 (N_2946,N_425,N_327);
or U2947 (N_2947,N_1548,N_1948);
nand U2948 (N_2948,N_1786,N_792);
and U2949 (N_2949,N_1924,N_1231);
and U2950 (N_2950,N_1353,N_651);
and U2951 (N_2951,N_1442,N_205);
nand U2952 (N_2952,N_1494,N_458);
xor U2953 (N_2953,N_1671,N_1003);
or U2954 (N_2954,N_1020,N_1861);
or U2955 (N_2955,N_1497,N_440);
and U2956 (N_2956,N_1804,N_825);
and U2957 (N_2957,N_1923,N_1210);
and U2958 (N_2958,N_1473,N_763);
or U2959 (N_2959,N_684,N_1453);
or U2960 (N_2960,N_960,N_12);
xor U2961 (N_2961,N_1903,N_494);
or U2962 (N_2962,N_319,N_996);
or U2963 (N_2963,N_1014,N_1402);
nor U2964 (N_2964,N_1656,N_87);
or U2965 (N_2965,N_1299,N_508);
or U2966 (N_2966,N_1301,N_1268);
and U2967 (N_2967,N_1320,N_1251);
nor U2968 (N_2968,N_1134,N_1248);
nand U2969 (N_2969,N_1013,N_1598);
nor U2970 (N_2970,N_34,N_1021);
nor U2971 (N_2971,N_781,N_994);
nor U2972 (N_2972,N_39,N_1284);
nand U2973 (N_2973,N_1572,N_1176);
and U2974 (N_2974,N_871,N_1622);
or U2975 (N_2975,N_341,N_31);
xor U2976 (N_2976,N_100,N_1426);
or U2977 (N_2977,N_1501,N_17);
or U2978 (N_2978,N_1966,N_265);
nor U2979 (N_2979,N_1166,N_1655);
nor U2980 (N_2980,N_1,N_1412);
or U2981 (N_2981,N_76,N_1650);
nand U2982 (N_2982,N_74,N_744);
nor U2983 (N_2983,N_1269,N_1352);
and U2984 (N_2984,N_1307,N_697);
nor U2985 (N_2985,N_1725,N_1469);
and U2986 (N_2986,N_739,N_1096);
and U2987 (N_2987,N_1266,N_1110);
or U2988 (N_2988,N_190,N_1149);
or U2989 (N_2989,N_958,N_654);
nor U2990 (N_2990,N_1126,N_1600);
and U2991 (N_2991,N_1922,N_1092);
nor U2992 (N_2992,N_1088,N_633);
or U2993 (N_2993,N_1907,N_1853);
nor U2994 (N_2994,N_1452,N_1128);
and U2995 (N_2995,N_101,N_1192);
xnor U2996 (N_2996,N_133,N_1105);
nand U2997 (N_2997,N_1302,N_1895);
and U2998 (N_2998,N_1612,N_1820);
xnor U2999 (N_2999,N_937,N_241);
or U3000 (N_3000,N_1289,N_412);
and U3001 (N_3001,N_1935,N_1213);
xnor U3002 (N_3002,N_897,N_1997);
or U3003 (N_3003,N_1228,N_1569);
or U3004 (N_3004,N_684,N_1765);
or U3005 (N_3005,N_265,N_1301);
nor U3006 (N_3006,N_1695,N_1748);
nor U3007 (N_3007,N_1417,N_706);
nand U3008 (N_3008,N_1268,N_1888);
nand U3009 (N_3009,N_415,N_1701);
nor U3010 (N_3010,N_1713,N_1243);
nor U3011 (N_3011,N_1807,N_666);
nand U3012 (N_3012,N_1097,N_1928);
and U3013 (N_3013,N_113,N_1566);
xor U3014 (N_3014,N_265,N_764);
nor U3015 (N_3015,N_520,N_345);
nand U3016 (N_3016,N_676,N_1402);
nor U3017 (N_3017,N_151,N_482);
and U3018 (N_3018,N_1199,N_1527);
or U3019 (N_3019,N_1354,N_872);
or U3020 (N_3020,N_1687,N_452);
or U3021 (N_3021,N_382,N_262);
nand U3022 (N_3022,N_1187,N_95);
and U3023 (N_3023,N_1007,N_1123);
nor U3024 (N_3024,N_1079,N_1323);
nand U3025 (N_3025,N_1296,N_407);
or U3026 (N_3026,N_1261,N_116);
nand U3027 (N_3027,N_554,N_1662);
nor U3028 (N_3028,N_384,N_1047);
and U3029 (N_3029,N_69,N_1122);
nand U3030 (N_3030,N_1748,N_869);
nor U3031 (N_3031,N_46,N_964);
nor U3032 (N_3032,N_1920,N_1944);
nand U3033 (N_3033,N_1006,N_679);
or U3034 (N_3034,N_196,N_1972);
nand U3035 (N_3035,N_1885,N_1388);
nand U3036 (N_3036,N_0,N_87);
or U3037 (N_3037,N_559,N_1523);
or U3038 (N_3038,N_983,N_1906);
nand U3039 (N_3039,N_1405,N_129);
or U3040 (N_3040,N_929,N_917);
or U3041 (N_3041,N_1710,N_328);
or U3042 (N_3042,N_1641,N_1886);
or U3043 (N_3043,N_362,N_1562);
nand U3044 (N_3044,N_271,N_1862);
nand U3045 (N_3045,N_1789,N_541);
and U3046 (N_3046,N_50,N_136);
nor U3047 (N_3047,N_179,N_1788);
and U3048 (N_3048,N_341,N_966);
or U3049 (N_3049,N_817,N_691);
nor U3050 (N_3050,N_327,N_448);
nand U3051 (N_3051,N_1239,N_219);
or U3052 (N_3052,N_274,N_1005);
nand U3053 (N_3053,N_1373,N_797);
nand U3054 (N_3054,N_984,N_804);
nor U3055 (N_3055,N_1358,N_448);
and U3056 (N_3056,N_1366,N_802);
and U3057 (N_3057,N_1691,N_813);
and U3058 (N_3058,N_1282,N_287);
nand U3059 (N_3059,N_594,N_1210);
nor U3060 (N_3060,N_742,N_620);
and U3061 (N_3061,N_1411,N_265);
and U3062 (N_3062,N_1383,N_674);
nor U3063 (N_3063,N_779,N_812);
or U3064 (N_3064,N_875,N_270);
and U3065 (N_3065,N_1102,N_1038);
and U3066 (N_3066,N_5,N_898);
nor U3067 (N_3067,N_425,N_983);
nand U3068 (N_3068,N_781,N_488);
nand U3069 (N_3069,N_1746,N_679);
xor U3070 (N_3070,N_1570,N_138);
or U3071 (N_3071,N_1996,N_1274);
nand U3072 (N_3072,N_1350,N_822);
nand U3073 (N_3073,N_1851,N_946);
nor U3074 (N_3074,N_1572,N_1256);
nand U3075 (N_3075,N_126,N_417);
xor U3076 (N_3076,N_1224,N_1880);
nand U3077 (N_3077,N_69,N_1894);
nor U3078 (N_3078,N_229,N_511);
xnor U3079 (N_3079,N_299,N_1195);
xor U3080 (N_3080,N_544,N_1943);
and U3081 (N_3081,N_1586,N_693);
and U3082 (N_3082,N_296,N_563);
or U3083 (N_3083,N_1914,N_601);
or U3084 (N_3084,N_1615,N_740);
and U3085 (N_3085,N_368,N_106);
and U3086 (N_3086,N_1860,N_974);
or U3087 (N_3087,N_1650,N_1557);
and U3088 (N_3088,N_1460,N_1994);
and U3089 (N_3089,N_1070,N_817);
nand U3090 (N_3090,N_694,N_1523);
or U3091 (N_3091,N_1572,N_1223);
or U3092 (N_3092,N_500,N_1338);
and U3093 (N_3093,N_1111,N_900);
and U3094 (N_3094,N_999,N_1043);
xnor U3095 (N_3095,N_268,N_1074);
or U3096 (N_3096,N_127,N_915);
nor U3097 (N_3097,N_1800,N_1287);
nor U3098 (N_3098,N_183,N_32);
and U3099 (N_3099,N_1044,N_1116);
or U3100 (N_3100,N_1424,N_497);
nor U3101 (N_3101,N_1800,N_84);
or U3102 (N_3102,N_66,N_553);
or U3103 (N_3103,N_1319,N_901);
or U3104 (N_3104,N_1774,N_486);
or U3105 (N_3105,N_1260,N_537);
and U3106 (N_3106,N_677,N_259);
nor U3107 (N_3107,N_363,N_1772);
nor U3108 (N_3108,N_910,N_818);
or U3109 (N_3109,N_962,N_1914);
and U3110 (N_3110,N_804,N_148);
or U3111 (N_3111,N_27,N_1026);
nand U3112 (N_3112,N_857,N_1864);
nor U3113 (N_3113,N_1901,N_824);
nand U3114 (N_3114,N_1283,N_866);
nand U3115 (N_3115,N_815,N_1452);
nor U3116 (N_3116,N_353,N_315);
and U3117 (N_3117,N_439,N_576);
xnor U3118 (N_3118,N_1555,N_1468);
nand U3119 (N_3119,N_376,N_656);
and U3120 (N_3120,N_1998,N_360);
xnor U3121 (N_3121,N_1614,N_648);
and U3122 (N_3122,N_202,N_1540);
and U3123 (N_3123,N_1447,N_1524);
xnor U3124 (N_3124,N_424,N_580);
nand U3125 (N_3125,N_730,N_1624);
or U3126 (N_3126,N_403,N_1309);
or U3127 (N_3127,N_1004,N_361);
nor U3128 (N_3128,N_1982,N_338);
or U3129 (N_3129,N_1151,N_291);
nor U3130 (N_3130,N_1488,N_792);
nor U3131 (N_3131,N_360,N_1689);
nand U3132 (N_3132,N_1478,N_1008);
and U3133 (N_3133,N_1275,N_1555);
xnor U3134 (N_3134,N_1110,N_1720);
and U3135 (N_3135,N_157,N_1324);
and U3136 (N_3136,N_1396,N_1016);
nor U3137 (N_3137,N_874,N_422);
nand U3138 (N_3138,N_1450,N_1820);
nor U3139 (N_3139,N_1811,N_609);
nor U3140 (N_3140,N_1588,N_1867);
nor U3141 (N_3141,N_1878,N_1802);
nor U3142 (N_3142,N_1098,N_1017);
nand U3143 (N_3143,N_618,N_648);
and U3144 (N_3144,N_535,N_1958);
and U3145 (N_3145,N_636,N_368);
and U3146 (N_3146,N_1723,N_1861);
xor U3147 (N_3147,N_155,N_69);
nor U3148 (N_3148,N_766,N_630);
or U3149 (N_3149,N_817,N_1852);
xnor U3150 (N_3150,N_1546,N_193);
nor U3151 (N_3151,N_701,N_1316);
nand U3152 (N_3152,N_449,N_288);
nand U3153 (N_3153,N_1897,N_74);
nor U3154 (N_3154,N_1105,N_125);
and U3155 (N_3155,N_151,N_1170);
xnor U3156 (N_3156,N_979,N_402);
nor U3157 (N_3157,N_1111,N_1032);
xnor U3158 (N_3158,N_1567,N_1825);
or U3159 (N_3159,N_1322,N_1909);
nor U3160 (N_3160,N_56,N_1822);
nand U3161 (N_3161,N_950,N_138);
nor U3162 (N_3162,N_1103,N_489);
xor U3163 (N_3163,N_1714,N_1158);
and U3164 (N_3164,N_1171,N_662);
xor U3165 (N_3165,N_1803,N_645);
nand U3166 (N_3166,N_1262,N_322);
or U3167 (N_3167,N_815,N_1426);
and U3168 (N_3168,N_1458,N_1814);
or U3169 (N_3169,N_14,N_294);
or U3170 (N_3170,N_1949,N_425);
and U3171 (N_3171,N_768,N_1285);
nand U3172 (N_3172,N_1175,N_676);
nor U3173 (N_3173,N_1673,N_1164);
or U3174 (N_3174,N_1992,N_151);
nor U3175 (N_3175,N_666,N_1046);
xnor U3176 (N_3176,N_1427,N_1783);
xnor U3177 (N_3177,N_1948,N_426);
or U3178 (N_3178,N_1857,N_1579);
nand U3179 (N_3179,N_1934,N_1618);
and U3180 (N_3180,N_586,N_967);
nand U3181 (N_3181,N_947,N_1337);
nand U3182 (N_3182,N_196,N_1218);
nand U3183 (N_3183,N_1509,N_398);
or U3184 (N_3184,N_594,N_75);
or U3185 (N_3185,N_780,N_104);
nor U3186 (N_3186,N_1665,N_1838);
nand U3187 (N_3187,N_846,N_1305);
or U3188 (N_3188,N_1001,N_301);
and U3189 (N_3189,N_256,N_894);
and U3190 (N_3190,N_632,N_1304);
nor U3191 (N_3191,N_305,N_228);
nand U3192 (N_3192,N_1015,N_471);
nand U3193 (N_3193,N_1935,N_330);
or U3194 (N_3194,N_823,N_1263);
nor U3195 (N_3195,N_203,N_920);
or U3196 (N_3196,N_1778,N_1582);
or U3197 (N_3197,N_693,N_494);
or U3198 (N_3198,N_1978,N_257);
or U3199 (N_3199,N_803,N_250);
or U3200 (N_3200,N_1254,N_1716);
or U3201 (N_3201,N_1098,N_566);
and U3202 (N_3202,N_1617,N_810);
and U3203 (N_3203,N_1367,N_1456);
or U3204 (N_3204,N_1004,N_711);
or U3205 (N_3205,N_1457,N_942);
nand U3206 (N_3206,N_1040,N_1780);
nand U3207 (N_3207,N_1016,N_559);
xor U3208 (N_3208,N_585,N_1880);
nor U3209 (N_3209,N_86,N_1842);
nand U3210 (N_3210,N_229,N_1744);
nor U3211 (N_3211,N_1111,N_928);
nand U3212 (N_3212,N_370,N_499);
and U3213 (N_3213,N_1520,N_772);
or U3214 (N_3214,N_1331,N_106);
xor U3215 (N_3215,N_629,N_1622);
or U3216 (N_3216,N_1312,N_1360);
or U3217 (N_3217,N_1581,N_1632);
and U3218 (N_3218,N_952,N_169);
and U3219 (N_3219,N_1254,N_367);
and U3220 (N_3220,N_1117,N_763);
nor U3221 (N_3221,N_1750,N_1629);
and U3222 (N_3222,N_527,N_888);
nand U3223 (N_3223,N_180,N_1985);
or U3224 (N_3224,N_528,N_540);
nand U3225 (N_3225,N_1348,N_1530);
and U3226 (N_3226,N_533,N_1098);
nand U3227 (N_3227,N_1221,N_44);
xor U3228 (N_3228,N_1263,N_752);
nand U3229 (N_3229,N_1310,N_698);
nor U3230 (N_3230,N_1635,N_803);
and U3231 (N_3231,N_1432,N_1173);
nand U3232 (N_3232,N_1601,N_425);
or U3233 (N_3233,N_131,N_1158);
nor U3234 (N_3234,N_1836,N_720);
or U3235 (N_3235,N_1538,N_1322);
or U3236 (N_3236,N_176,N_1629);
or U3237 (N_3237,N_1560,N_66);
and U3238 (N_3238,N_291,N_850);
nand U3239 (N_3239,N_426,N_385);
nor U3240 (N_3240,N_659,N_1294);
nand U3241 (N_3241,N_269,N_264);
nor U3242 (N_3242,N_1746,N_961);
nand U3243 (N_3243,N_967,N_764);
nand U3244 (N_3244,N_97,N_617);
nor U3245 (N_3245,N_1579,N_136);
nor U3246 (N_3246,N_71,N_1134);
nor U3247 (N_3247,N_1353,N_987);
or U3248 (N_3248,N_1139,N_1800);
xor U3249 (N_3249,N_1808,N_1284);
nand U3250 (N_3250,N_728,N_1941);
or U3251 (N_3251,N_468,N_497);
or U3252 (N_3252,N_1529,N_84);
and U3253 (N_3253,N_1264,N_234);
nand U3254 (N_3254,N_1175,N_441);
and U3255 (N_3255,N_1096,N_700);
or U3256 (N_3256,N_352,N_1346);
xnor U3257 (N_3257,N_752,N_342);
or U3258 (N_3258,N_20,N_29);
or U3259 (N_3259,N_667,N_560);
xor U3260 (N_3260,N_1745,N_1899);
or U3261 (N_3261,N_337,N_1957);
nand U3262 (N_3262,N_1834,N_1);
nand U3263 (N_3263,N_1331,N_678);
nor U3264 (N_3264,N_54,N_299);
and U3265 (N_3265,N_1954,N_1387);
nand U3266 (N_3266,N_464,N_1295);
nor U3267 (N_3267,N_756,N_498);
nand U3268 (N_3268,N_316,N_1047);
xnor U3269 (N_3269,N_1983,N_1773);
or U3270 (N_3270,N_1900,N_157);
nor U3271 (N_3271,N_315,N_534);
or U3272 (N_3272,N_797,N_1207);
nor U3273 (N_3273,N_1440,N_361);
or U3274 (N_3274,N_1730,N_1534);
or U3275 (N_3275,N_1742,N_111);
nand U3276 (N_3276,N_949,N_300);
nor U3277 (N_3277,N_1036,N_159);
or U3278 (N_3278,N_952,N_731);
or U3279 (N_3279,N_551,N_357);
and U3280 (N_3280,N_939,N_1881);
nor U3281 (N_3281,N_224,N_107);
nand U3282 (N_3282,N_1572,N_788);
nand U3283 (N_3283,N_1342,N_1869);
or U3284 (N_3284,N_1874,N_1414);
nor U3285 (N_3285,N_862,N_1712);
nand U3286 (N_3286,N_514,N_312);
nor U3287 (N_3287,N_220,N_173);
and U3288 (N_3288,N_895,N_239);
and U3289 (N_3289,N_1880,N_1791);
and U3290 (N_3290,N_1424,N_166);
and U3291 (N_3291,N_1991,N_101);
or U3292 (N_3292,N_1171,N_1551);
or U3293 (N_3293,N_1520,N_1806);
or U3294 (N_3294,N_1898,N_509);
nand U3295 (N_3295,N_1834,N_1304);
nand U3296 (N_3296,N_678,N_918);
nand U3297 (N_3297,N_524,N_15);
and U3298 (N_3298,N_378,N_432);
nand U3299 (N_3299,N_768,N_1035);
nand U3300 (N_3300,N_1071,N_724);
and U3301 (N_3301,N_1150,N_558);
xor U3302 (N_3302,N_1870,N_1760);
or U3303 (N_3303,N_1463,N_381);
and U3304 (N_3304,N_766,N_1555);
nand U3305 (N_3305,N_868,N_1509);
and U3306 (N_3306,N_1845,N_1774);
nand U3307 (N_3307,N_956,N_462);
or U3308 (N_3308,N_701,N_1119);
and U3309 (N_3309,N_1757,N_1400);
nand U3310 (N_3310,N_1105,N_1737);
and U3311 (N_3311,N_1714,N_618);
nor U3312 (N_3312,N_918,N_1214);
nor U3313 (N_3313,N_294,N_1700);
nor U3314 (N_3314,N_1820,N_528);
xnor U3315 (N_3315,N_188,N_338);
or U3316 (N_3316,N_766,N_354);
xnor U3317 (N_3317,N_675,N_931);
nor U3318 (N_3318,N_1829,N_631);
xnor U3319 (N_3319,N_1603,N_1971);
xor U3320 (N_3320,N_183,N_306);
or U3321 (N_3321,N_1137,N_934);
and U3322 (N_3322,N_298,N_1040);
and U3323 (N_3323,N_1059,N_938);
or U3324 (N_3324,N_1808,N_1010);
nand U3325 (N_3325,N_1675,N_1833);
nand U3326 (N_3326,N_377,N_1013);
or U3327 (N_3327,N_874,N_170);
nor U3328 (N_3328,N_38,N_1197);
nand U3329 (N_3329,N_1739,N_1909);
or U3330 (N_3330,N_1691,N_493);
or U3331 (N_3331,N_1396,N_1111);
or U3332 (N_3332,N_523,N_1598);
nand U3333 (N_3333,N_1001,N_563);
or U3334 (N_3334,N_1945,N_1940);
or U3335 (N_3335,N_1586,N_1532);
nor U3336 (N_3336,N_774,N_511);
and U3337 (N_3337,N_569,N_1060);
or U3338 (N_3338,N_929,N_1175);
nand U3339 (N_3339,N_1539,N_1046);
nor U3340 (N_3340,N_1418,N_1274);
nor U3341 (N_3341,N_1012,N_1195);
and U3342 (N_3342,N_1070,N_724);
nand U3343 (N_3343,N_955,N_1778);
nand U3344 (N_3344,N_1083,N_222);
and U3345 (N_3345,N_597,N_217);
nor U3346 (N_3346,N_420,N_1479);
and U3347 (N_3347,N_395,N_484);
nor U3348 (N_3348,N_1459,N_1374);
or U3349 (N_3349,N_1418,N_342);
nand U3350 (N_3350,N_47,N_1663);
nor U3351 (N_3351,N_1212,N_1540);
or U3352 (N_3352,N_1082,N_745);
or U3353 (N_3353,N_859,N_700);
and U3354 (N_3354,N_401,N_525);
nand U3355 (N_3355,N_525,N_1048);
and U3356 (N_3356,N_184,N_1479);
nand U3357 (N_3357,N_1482,N_1138);
or U3358 (N_3358,N_1387,N_1705);
nor U3359 (N_3359,N_1242,N_1830);
and U3360 (N_3360,N_863,N_326);
or U3361 (N_3361,N_1360,N_474);
or U3362 (N_3362,N_1293,N_1371);
or U3363 (N_3363,N_1355,N_1272);
nand U3364 (N_3364,N_545,N_39);
and U3365 (N_3365,N_1675,N_1013);
and U3366 (N_3366,N_1764,N_1628);
xor U3367 (N_3367,N_798,N_318);
nor U3368 (N_3368,N_1819,N_75);
nand U3369 (N_3369,N_239,N_1711);
and U3370 (N_3370,N_1694,N_53);
nor U3371 (N_3371,N_1603,N_595);
and U3372 (N_3372,N_683,N_1525);
nand U3373 (N_3373,N_1174,N_1197);
nor U3374 (N_3374,N_1907,N_808);
nor U3375 (N_3375,N_770,N_82);
nor U3376 (N_3376,N_706,N_1851);
nor U3377 (N_3377,N_623,N_1436);
or U3378 (N_3378,N_669,N_1055);
nand U3379 (N_3379,N_346,N_1447);
or U3380 (N_3380,N_365,N_1672);
and U3381 (N_3381,N_228,N_931);
xnor U3382 (N_3382,N_175,N_807);
or U3383 (N_3383,N_1314,N_27);
xor U3384 (N_3384,N_1560,N_1484);
xnor U3385 (N_3385,N_799,N_1519);
nand U3386 (N_3386,N_892,N_876);
nand U3387 (N_3387,N_954,N_922);
or U3388 (N_3388,N_554,N_1688);
nand U3389 (N_3389,N_1558,N_1286);
and U3390 (N_3390,N_1153,N_1500);
or U3391 (N_3391,N_229,N_1467);
xnor U3392 (N_3392,N_31,N_571);
nand U3393 (N_3393,N_1669,N_111);
nand U3394 (N_3394,N_1305,N_1845);
nand U3395 (N_3395,N_1418,N_1127);
and U3396 (N_3396,N_66,N_531);
and U3397 (N_3397,N_1857,N_1135);
xor U3398 (N_3398,N_806,N_441);
nand U3399 (N_3399,N_254,N_570);
and U3400 (N_3400,N_912,N_1047);
or U3401 (N_3401,N_1434,N_958);
nor U3402 (N_3402,N_119,N_1180);
nand U3403 (N_3403,N_1687,N_1629);
xor U3404 (N_3404,N_382,N_621);
nor U3405 (N_3405,N_1054,N_1793);
nand U3406 (N_3406,N_1824,N_960);
nand U3407 (N_3407,N_1865,N_766);
or U3408 (N_3408,N_1170,N_634);
and U3409 (N_3409,N_1967,N_1201);
nand U3410 (N_3410,N_243,N_1305);
xor U3411 (N_3411,N_913,N_94);
xor U3412 (N_3412,N_1974,N_1001);
and U3413 (N_3413,N_1612,N_1906);
nor U3414 (N_3414,N_185,N_1377);
nor U3415 (N_3415,N_303,N_413);
and U3416 (N_3416,N_979,N_1734);
and U3417 (N_3417,N_952,N_1777);
nand U3418 (N_3418,N_1057,N_23);
and U3419 (N_3419,N_655,N_1308);
nand U3420 (N_3420,N_787,N_907);
or U3421 (N_3421,N_790,N_765);
nand U3422 (N_3422,N_374,N_1963);
and U3423 (N_3423,N_784,N_1714);
and U3424 (N_3424,N_282,N_1569);
nand U3425 (N_3425,N_1604,N_749);
nand U3426 (N_3426,N_329,N_983);
and U3427 (N_3427,N_280,N_668);
or U3428 (N_3428,N_857,N_1375);
and U3429 (N_3429,N_1348,N_1005);
xnor U3430 (N_3430,N_910,N_409);
nand U3431 (N_3431,N_1084,N_904);
or U3432 (N_3432,N_1208,N_1215);
and U3433 (N_3433,N_753,N_1450);
or U3434 (N_3434,N_594,N_1316);
xor U3435 (N_3435,N_1959,N_965);
and U3436 (N_3436,N_1429,N_646);
and U3437 (N_3437,N_1123,N_1813);
nand U3438 (N_3438,N_876,N_1334);
xnor U3439 (N_3439,N_458,N_1799);
nand U3440 (N_3440,N_1966,N_175);
and U3441 (N_3441,N_1064,N_291);
and U3442 (N_3442,N_587,N_845);
nor U3443 (N_3443,N_1857,N_595);
or U3444 (N_3444,N_1867,N_918);
and U3445 (N_3445,N_1716,N_180);
nand U3446 (N_3446,N_1797,N_204);
or U3447 (N_3447,N_1975,N_302);
nand U3448 (N_3448,N_76,N_681);
or U3449 (N_3449,N_937,N_408);
or U3450 (N_3450,N_798,N_990);
nor U3451 (N_3451,N_464,N_1267);
nand U3452 (N_3452,N_826,N_1556);
and U3453 (N_3453,N_16,N_1530);
nand U3454 (N_3454,N_1520,N_1450);
nor U3455 (N_3455,N_372,N_1503);
and U3456 (N_3456,N_1769,N_750);
nand U3457 (N_3457,N_1791,N_1187);
xnor U3458 (N_3458,N_956,N_1781);
nor U3459 (N_3459,N_1775,N_1350);
or U3460 (N_3460,N_1511,N_208);
and U3461 (N_3461,N_1968,N_1104);
nor U3462 (N_3462,N_1319,N_444);
nand U3463 (N_3463,N_628,N_103);
xor U3464 (N_3464,N_1933,N_1492);
nand U3465 (N_3465,N_1533,N_1875);
and U3466 (N_3466,N_234,N_1026);
nor U3467 (N_3467,N_949,N_208);
nor U3468 (N_3468,N_860,N_1251);
nand U3469 (N_3469,N_1113,N_1985);
nor U3470 (N_3470,N_776,N_184);
or U3471 (N_3471,N_1567,N_532);
and U3472 (N_3472,N_1213,N_1912);
and U3473 (N_3473,N_1890,N_896);
and U3474 (N_3474,N_5,N_1298);
nand U3475 (N_3475,N_937,N_1452);
xor U3476 (N_3476,N_1385,N_231);
nand U3477 (N_3477,N_1190,N_853);
or U3478 (N_3478,N_1449,N_697);
and U3479 (N_3479,N_1800,N_1937);
nand U3480 (N_3480,N_1881,N_995);
nand U3481 (N_3481,N_508,N_1841);
nor U3482 (N_3482,N_1275,N_1426);
and U3483 (N_3483,N_1912,N_75);
and U3484 (N_3484,N_885,N_273);
nor U3485 (N_3485,N_639,N_634);
or U3486 (N_3486,N_91,N_12);
nor U3487 (N_3487,N_140,N_1352);
and U3488 (N_3488,N_1416,N_903);
nor U3489 (N_3489,N_1077,N_799);
nand U3490 (N_3490,N_391,N_799);
and U3491 (N_3491,N_1189,N_1399);
nand U3492 (N_3492,N_121,N_1472);
nand U3493 (N_3493,N_474,N_1366);
nor U3494 (N_3494,N_1480,N_1718);
and U3495 (N_3495,N_1867,N_683);
nand U3496 (N_3496,N_1230,N_1766);
or U3497 (N_3497,N_648,N_1137);
nor U3498 (N_3498,N_555,N_627);
and U3499 (N_3499,N_1287,N_552);
and U3500 (N_3500,N_1324,N_1402);
or U3501 (N_3501,N_842,N_495);
nor U3502 (N_3502,N_164,N_1358);
and U3503 (N_3503,N_389,N_257);
nand U3504 (N_3504,N_1619,N_453);
and U3505 (N_3505,N_1561,N_1852);
or U3506 (N_3506,N_1665,N_1478);
nor U3507 (N_3507,N_1557,N_1832);
nor U3508 (N_3508,N_485,N_339);
nand U3509 (N_3509,N_593,N_1178);
or U3510 (N_3510,N_1104,N_1900);
and U3511 (N_3511,N_1021,N_1646);
nor U3512 (N_3512,N_1015,N_1180);
nand U3513 (N_3513,N_685,N_765);
nand U3514 (N_3514,N_772,N_387);
and U3515 (N_3515,N_1478,N_436);
or U3516 (N_3516,N_1808,N_349);
nand U3517 (N_3517,N_565,N_1861);
nand U3518 (N_3518,N_1410,N_1005);
nand U3519 (N_3519,N_517,N_271);
nor U3520 (N_3520,N_1458,N_573);
nand U3521 (N_3521,N_1359,N_504);
and U3522 (N_3522,N_1495,N_985);
nor U3523 (N_3523,N_1467,N_1156);
nand U3524 (N_3524,N_312,N_1996);
or U3525 (N_3525,N_1842,N_300);
nor U3526 (N_3526,N_350,N_820);
or U3527 (N_3527,N_1257,N_9);
nand U3528 (N_3528,N_1126,N_624);
nand U3529 (N_3529,N_1813,N_80);
nand U3530 (N_3530,N_1476,N_629);
nor U3531 (N_3531,N_813,N_249);
and U3532 (N_3532,N_385,N_111);
and U3533 (N_3533,N_769,N_1723);
nand U3534 (N_3534,N_253,N_1409);
or U3535 (N_3535,N_1916,N_604);
nor U3536 (N_3536,N_650,N_1478);
nor U3537 (N_3537,N_488,N_1511);
xnor U3538 (N_3538,N_872,N_536);
xnor U3539 (N_3539,N_565,N_922);
nor U3540 (N_3540,N_391,N_1278);
nand U3541 (N_3541,N_198,N_1275);
nand U3542 (N_3542,N_1584,N_534);
nor U3543 (N_3543,N_1842,N_330);
or U3544 (N_3544,N_903,N_1061);
xor U3545 (N_3545,N_997,N_1462);
xor U3546 (N_3546,N_970,N_994);
xnor U3547 (N_3547,N_941,N_1957);
nor U3548 (N_3548,N_391,N_1268);
or U3549 (N_3549,N_138,N_646);
nand U3550 (N_3550,N_55,N_1241);
xnor U3551 (N_3551,N_1375,N_1044);
and U3552 (N_3552,N_913,N_1058);
nor U3553 (N_3553,N_1492,N_700);
xnor U3554 (N_3554,N_718,N_1197);
or U3555 (N_3555,N_1912,N_574);
or U3556 (N_3556,N_1943,N_374);
nand U3557 (N_3557,N_68,N_123);
xor U3558 (N_3558,N_1738,N_605);
or U3559 (N_3559,N_709,N_1600);
nor U3560 (N_3560,N_164,N_1775);
nand U3561 (N_3561,N_1913,N_1629);
nor U3562 (N_3562,N_1516,N_576);
nand U3563 (N_3563,N_716,N_722);
xnor U3564 (N_3564,N_995,N_750);
nor U3565 (N_3565,N_1135,N_1813);
or U3566 (N_3566,N_768,N_1036);
and U3567 (N_3567,N_1013,N_1580);
nor U3568 (N_3568,N_1544,N_1627);
xor U3569 (N_3569,N_930,N_43);
or U3570 (N_3570,N_850,N_1672);
or U3571 (N_3571,N_20,N_465);
and U3572 (N_3572,N_1093,N_856);
and U3573 (N_3573,N_1399,N_845);
nor U3574 (N_3574,N_247,N_1432);
xnor U3575 (N_3575,N_1427,N_733);
nand U3576 (N_3576,N_1729,N_1184);
or U3577 (N_3577,N_212,N_108);
and U3578 (N_3578,N_1163,N_243);
nor U3579 (N_3579,N_572,N_1759);
nor U3580 (N_3580,N_770,N_496);
nor U3581 (N_3581,N_1627,N_1117);
and U3582 (N_3582,N_92,N_135);
or U3583 (N_3583,N_1530,N_824);
nor U3584 (N_3584,N_758,N_1111);
nand U3585 (N_3585,N_633,N_249);
and U3586 (N_3586,N_1461,N_1499);
nor U3587 (N_3587,N_131,N_1701);
or U3588 (N_3588,N_476,N_1274);
nor U3589 (N_3589,N_528,N_1695);
nor U3590 (N_3590,N_281,N_1075);
nand U3591 (N_3591,N_1851,N_1710);
or U3592 (N_3592,N_1004,N_487);
or U3593 (N_3593,N_322,N_1502);
nand U3594 (N_3594,N_668,N_865);
nand U3595 (N_3595,N_1726,N_151);
and U3596 (N_3596,N_1831,N_719);
xnor U3597 (N_3597,N_27,N_1459);
or U3598 (N_3598,N_1238,N_1000);
and U3599 (N_3599,N_693,N_1138);
and U3600 (N_3600,N_1393,N_315);
and U3601 (N_3601,N_934,N_1504);
or U3602 (N_3602,N_1587,N_1838);
or U3603 (N_3603,N_1443,N_1574);
and U3604 (N_3604,N_1483,N_286);
nor U3605 (N_3605,N_1185,N_1385);
nand U3606 (N_3606,N_543,N_890);
nor U3607 (N_3607,N_553,N_988);
nand U3608 (N_3608,N_999,N_1436);
and U3609 (N_3609,N_145,N_676);
nand U3610 (N_3610,N_1157,N_402);
or U3611 (N_3611,N_382,N_1754);
and U3612 (N_3612,N_500,N_804);
nand U3613 (N_3613,N_1079,N_151);
or U3614 (N_3614,N_1705,N_1933);
nor U3615 (N_3615,N_1429,N_536);
nand U3616 (N_3616,N_1579,N_867);
and U3617 (N_3617,N_1828,N_1597);
or U3618 (N_3618,N_494,N_1979);
xor U3619 (N_3619,N_176,N_147);
and U3620 (N_3620,N_866,N_415);
nand U3621 (N_3621,N_89,N_513);
and U3622 (N_3622,N_239,N_507);
and U3623 (N_3623,N_1739,N_1394);
or U3624 (N_3624,N_1283,N_1445);
or U3625 (N_3625,N_1347,N_1021);
nand U3626 (N_3626,N_1634,N_1938);
or U3627 (N_3627,N_1439,N_1964);
or U3628 (N_3628,N_992,N_1733);
xor U3629 (N_3629,N_1534,N_650);
and U3630 (N_3630,N_1514,N_1298);
nor U3631 (N_3631,N_683,N_1577);
nor U3632 (N_3632,N_1541,N_185);
or U3633 (N_3633,N_1998,N_22);
xnor U3634 (N_3634,N_1516,N_221);
nand U3635 (N_3635,N_856,N_1388);
nand U3636 (N_3636,N_1732,N_1941);
xnor U3637 (N_3637,N_988,N_78);
nor U3638 (N_3638,N_871,N_1557);
nand U3639 (N_3639,N_1377,N_668);
and U3640 (N_3640,N_1376,N_1556);
and U3641 (N_3641,N_1806,N_264);
nor U3642 (N_3642,N_469,N_800);
nor U3643 (N_3643,N_992,N_1224);
nand U3644 (N_3644,N_1465,N_1942);
nand U3645 (N_3645,N_314,N_932);
xnor U3646 (N_3646,N_797,N_1288);
nand U3647 (N_3647,N_476,N_555);
nor U3648 (N_3648,N_1076,N_1434);
or U3649 (N_3649,N_856,N_1752);
or U3650 (N_3650,N_1976,N_296);
and U3651 (N_3651,N_567,N_1366);
nor U3652 (N_3652,N_1859,N_580);
nand U3653 (N_3653,N_1355,N_1608);
xor U3654 (N_3654,N_201,N_1443);
nor U3655 (N_3655,N_56,N_1782);
xnor U3656 (N_3656,N_1100,N_1457);
or U3657 (N_3657,N_1920,N_130);
or U3658 (N_3658,N_1488,N_1439);
or U3659 (N_3659,N_1446,N_1050);
nand U3660 (N_3660,N_810,N_1939);
nor U3661 (N_3661,N_932,N_1608);
nor U3662 (N_3662,N_484,N_1332);
or U3663 (N_3663,N_124,N_1745);
or U3664 (N_3664,N_1813,N_1130);
xnor U3665 (N_3665,N_1192,N_1629);
and U3666 (N_3666,N_1184,N_1387);
or U3667 (N_3667,N_110,N_766);
or U3668 (N_3668,N_887,N_28);
nor U3669 (N_3669,N_714,N_454);
nand U3670 (N_3670,N_148,N_984);
nor U3671 (N_3671,N_1943,N_1640);
or U3672 (N_3672,N_1333,N_403);
and U3673 (N_3673,N_556,N_1962);
nor U3674 (N_3674,N_454,N_365);
and U3675 (N_3675,N_374,N_1038);
or U3676 (N_3676,N_1329,N_535);
nor U3677 (N_3677,N_690,N_1393);
xnor U3678 (N_3678,N_101,N_1797);
nand U3679 (N_3679,N_1895,N_1655);
nor U3680 (N_3680,N_824,N_403);
or U3681 (N_3681,N_1160,N_426);
nand U3682 (N_3682,N_853,N_1913);
nand U3683 (N_3683,N_1558,N_319);
nand U3684 (N_3684,N_1776,N_68);
or U3685 (N_3685,N_1845,N_330);
and U3686 (N_3686,N_1774,N_362);
nor U3687 (N_3687,N_1098,N_1517);
or U3688 (N_3688,N_1858,N_703);
nor U3689 (N_3689,N_1666,N_1051);
nand U3690 (N_3690,N_1132,N_523);
or U3691 (N_3691,N_1884,N_1432);
nand U3692 (N_3692,N_41,N_107);
nor U3693 (N_3693,N_243,N_724);
or U3694 (N_3694,N_1452,N_398);
or U3695 (N_3695,N_1502,N_278);
nor U3696 (N_3696,N_1273,N_487);
nor U3697 (N_3697,N_1612,N_147);
xor U3698 (N_3698,N_287,N_949);
or U3699 (N_3699,N_0,N_1160);
nand U3700 (N_3700,N_1521,N_1211);
nor U3701 (N_3701,N_1058,N_760);
nand U3702 (N_3702,N_1037,N_1284);
xnor U3703 (N_3703,N_1010,N_1745);
xor U3704 (N_3704,N_1688,N_1024);
and U3705 (N_3705,N_1827,N_65);
nor U3706 (N_3706,N_1855,N_1963);
nor U3707 (N_3707,N_1865,N_757);
or U3708 (N_3708,N_203,N_618);
xor U3709 (N_3709,N_1950,N_943);
xor U3710 (N_3710,N_1423,N_957);
nor U3711 (N_3711,N_1743,N_1783);
nor U3712 (N_3712,N_445,N_1826);
or U3713 (N_3713,N_1878,N_1025);
nor U3714 (N_3714,N_123,N_581);
nor U3715 (N_3715,N_753,N_205);
or U3716 (N_3716,N_1872,N_1145);
and U3717 (N_3717,N_608,N_653);
nor U3718 (N_3718,N_1427,N_950);
or U3719 (N_3719,N_1726,N_1886);
or U3720 (N_3720,N_782,N_440);
xnor U3721 (N_3721,N_359,N_1075);
or U3722 (N_3722,N_723,N_747);
nand U3723 (N_3723,N_893,N_880);
and U3724 (N_3724,N_822,N_224);
or U3725 (N_3725,N_968,N_423);
nand U3726 (N_3726,N_1938,N_1687);
nor U3727 (N_3727,N_171,N_1727);
and U3728 (N_3728,N_298,N_1302);
and U3729 (N_3729,N_1656,N_1187);
xor U3730 (N_3730,N_1020,N_1396);
nand U3731 (N_3731,N_1500,N_573);
or U3732 (N_3732,N_1009,N_159);
xor U3733 (N_3733,N_1545,N_150);
nand U3734 (N_3734,N_702,N_1318);
nor U3735 (N_3735,N_1274,N_800);
and U3736 (N_3736,N_1716,N_1986);
nor U3737 (N_3737,N_903,N_81);
xnor U3738 (N_3738,N_1136,N_104);
and U3739 (N_3739,N_1469,N_1609);
nand U3740 (N_3740,N_863,N_1114);
or U3741 (N_3741,N_1552,N_1228);
xor U3742 (N_3742,N_84,N_1195);
or U3743 (N_3743,N_315,N_602);
nand U3744 (N_3744,N_419,N_1069);
or U3745 (N_3745,N_1099,N_993);
or U3746 (N_3746,N_445,N_1176);
xor U3747 (N_3747,N_1156,N_287);
nor U3748 (N_3748,N_1559,N_1619);
nor U3749 (N_3749,N_926,N_496);
or U3750 (N_3750,N_1529,N_985);
and U3751 (N_3751,N_149,N_1493);
nor U3752 (N_3752,N_413,N_1803);
or U3753 (N_3753,N_1045,N_1613);
and U3754 (N_3754,N_188,N_56);
nand U3755 (N_3755,N_202,N_603);
and U3756 (N_3756,N_1259,N_1187);
nand U3757 (N_3757,N_601,N_15);
and U3758 (N_3758,N_1946,N_1074);
or U3759 (N_3759,N_442,N_431);
nor U3760 (N_3760,N_1907,N_28);
nor U3761 (N_3761,N_1728,N_829);
and U3762 (N_3762,N_1262,N_1318);
nor U3763 (N_3763,N_272,N_1193);
and U3764 (N_3764,N_1079,N_297);
nor U3765 (N_3765,N_138,N_1860);
xnor U3766 (N_3766,N_1356,N_487);
nand U3767 (N_3767,N_1210,N_993);
nand U3768 (N_3768,N_1571,N_1835);
xor U3769 (N_3769,N_237,N_1094);
and U3770 (N_3770,N_1715,N_875);
or U3771 (N_3771,N_1911,N_329);
or U3772 (N_3772,N_1151,N_1229);
and U3773 (N_3773,N_1196,N_1489);
nand U3774 (N_3774,N_375,N_371);
or U3775 (N_3775,N_528,N_430);
xnor U3776 (N_3776,N_1979,N_822);
and U3777 (N_3777,N_1593,N_571);
or U3778 (N_3778,N_394,N_1731);
xnor U3779 (N_3779,N_1716,N_357);
and U3780 (N_3780,N_1209,N_380);
nand U3781 (N_3781,N_949,N_273);
nor U3782 (N_3782,N_1278,N_1823);
or U3783 (N_3783,N_1852,N_954);
nor U3784 (N_3784,N_1094,N_440);
xor U3785 (N_3785,N_1702,N_337);
or U3786 (N_3786,N_505,N_1060);
or U3787 (N_3787,N_1708,N_1234);
nor U3788 (N_3788,N_248,N_905);
nor U3789 (N_3789,N_650,N_1103);
nor U3790 (N_3790,N_1266,N_618);
xor U3791 (N_3791,N_1097,N_1085);
xor U3792 (N_3792,N_1456,N_705);
and U3793 (N_3793,N_909,N_1940);
nand U3794 (N_3794,N_587,N_1008);
and U3795 (N_3795,N_1471,N_1186);
or U3796 (N_3796,N_386,N_31);
and U3797 (N_3797,N_849,N_526);
and U3798 (N_3798,N_284,N_421);
nor U3799 (N_3799,N_1171,N_650);
nor U3800 (N_3800,N_1469,N_1464);
or U3801 (N_3801,N_1549,N_157);
nand U3802 (N_3802,N_884,N_1717);
nor U3803 (N_3803,N_1515,N_14);
nand U3804 (N_3804,N_347,N_762);
nor U3805 (N_3805,N_809,N_1486);
nor U3806 (N_3806,N_1400,N_1550);
and U3807 (N_3807,N_1323,N_1674);
nand U3808 (N_3808,N_607,N_663);
and U3809 (N_3809,N_863,N_1780);
nor U3810 (N_3810,N_743,N_934);
and U3811 (N_3811,N_1004,N_1320);
and U3812 (N_3812,N_1748,N_1369);
and U3813 (N_3813,N_864,N_1885);
nand U3814 (N_3814,N_446,N_1063);
nand U3815 (N_3815,N_1654,N_1419);
nand U3816 (N_3816,N_901,N_1117);
or U3817 (N_3817,N_360,N_1929);
and U3818 (N_3818,N_1159,N_1878);
or U3819 (N_3819,N_796,N_620);
and U3820 (N_3820,N_504,N_1449);
xor U3821 (N_3821,N_1490,N_1903);
and U3822 (N_3822,N_1093,N_1313);
xor U3823 (N_3823,N_1836,N_758);
or U3824 (N_3824,N_825,N_1549);
nor U3825 (N_3825,N_592,N_1958);
or U3826 (N_3826,N_921,N_1065);
or U3827 (N_3827,N_1895,N_1867);
nand U3828 (N_3828,N_1410,N_385);
nor U3829 (N_3829,N_929,N_936);
and U3830 (N_3830,N_935,N_978);
nand U3831 (N_3831,N_14,N_519);
nand U3832 (N_3832,N_1661,N_302);
xnor U3833 (N_3833,N_621,N_743);
and U3834 (N_3834,N_1209,N_489);
or U3835 (N_3835,N_413,N_1366);
nor U3836 (N_3836,N_1761,N_200);
and U3837 (N_3837,N_3,N_801);
and U3838 (N_3838,N_926,N_143);
nor U3839 (N_3839,N_352,N_750);
or U3840 (N_3840,N_1014,N_275);
nand U3841 (N_3841,N_1275,N_985);
xnor U3842 (N_3842,N_720,N_1310);
or U3843 (N_3843,N_971,N_1039);
or U3844 (N_3844,N_1373,N_925);
nor U3845 (N_3845,N_863,N_1142);
or U3846 (N_3846,N_1339,N_253);
nand U3847 (N_3847,N_1276,N_1496);
nor U3848 (N_3848,N_661,N_907);
nor U3849 (N_3849,N_606,N_585);
nand U3850 (N_3850,N_1921,N_890);
nor U3851 (N_3851,N_6,N_1437);
nand U3852 (N_3852,N_1254,N_1163);
and U3853 (N_3853,N_479,N_1058);
nand U3854 (N_3854,N_1681,N_1834);
nor U3855 (N_3855,N_938,N_1419);
or U3856 (N_3856,N_817,N_368);
nor U3857 (N_3857,N_1379,N_1638);
nand U3858 (N_3858,N_292,N_1194);
xor U3859 (N_3859,N_1712,N_1595);
nand U3860 (N_3860,N_1797,N_169);
or U3861 (N_3861,N_719,N_1302);
nor U3862 (N_3862,N_990,N_1883);
nand U3863 (N_3863,N_1611,N_580);
nand U3864 (N_3864,N_1156,N_1247);
or U3865 (N_3865,N_1395,N_1489);
nor U3866 (N_3866,N_158,N_1113);
xor U3867 (N_3867,N_956,N_967);
and U3868 (N_3868,N_787,N_1673);
or U3869 (N_3869,N_1852,N_396);
nand U3870 (N_3870,N_847,N_1575);
nor U3871 (N_3871,N_1169,N_564);
and U3872 (N_3872,N_1408,N_59);
nand U3873 (N_3873,N_662,N_1328);
nor U3874 (N_3874,N_1998,N_1677);
nand U3875 (N_3875,N_1357,N_1816);
and U3876 (N_3876,N_1603,N_1901);
or U3877 (N_3877,N_193,N_790);
nand U3878 (N_3878,N_1001,N_1465);
nor U3879 (N_3879,N_419,N_902);
nand U3880 (N_3880,N_367,N_476);
and U3881 (N_3881,N_893,N_1096);
or U3882 (N_3882,N_1909,N_1811);
nor U3883 (N_3883,N_594,N_1593);
and U3884 (N_3884,N_691,N_1115);
or U3885 (N_3885,N_408,N_1730);
nand U3886 (N_3886,N_398,N_1388);
nand U3887 (N_3887,N_1519,N_1819);
and U3888 (N_3888,N_1261,N_780);
nand U3889 (N_3889,N_126,N_1489);
nor U3890 (N_3890,N_1731,N_1251);
nor U3891 (N_3891,N_1503,N_1658);
nand U3892 (N_3892,N_1215,N_1493);
xor U3893 (N_3893,N_1545,N_319);
nor U3894 (N_3894,N_1464,N_519);
nand U3895 (N_3895,N_1320,N_369);
nor U3896 (N_3896,N_1179,N_805);
nor U3897 (N_3897,N_1022,N_811);
nand U3898 (N_3898,N_1703,N_381);
nand U3899 (N_3899,N_71,N_1191);
or U3900 (N_3900,N_1068,N_1517);
and U3901 (N_3901,N_1136,N_1411);
nand U3902 (N_3902,N_1639,N_1087);
nor U3903 (N_3903,N_1600,N_1850);
nand U3904 (N_3904,N_556,N_1202);
nand U3905 (N_3905,N_300,N_1532);
and U3906 (N_3906,N_780,N_346);
or U3907 (N_3907,N_1592,N_1405);
nor U3908 (N_3908,N_1883,N_1483);
and U3909 (N_3909,N_1287,N_1732);
or U3910 (N_3910,N_1198,N_725);
xor U3911 (N_3911,N_1585,N_1151);
and U3912 (N_3912,N_1355,N_1764);
xnor U3913 (N_3913,N_1444,N_1161);
or U3914 (N_3914,N_1310,N_747);
xor U3915 (N_3915,N_1913,N_1683);
or U3916 (N_3916,N_1387,N_376);
nand U3917 (N_3917,N_190,N_1242);
nor U3918 (N_3918,N_1319,N_1370);
nor U3919 (N_3919,N_1111,N_1277);
nor U3920 (N_3920,N_682,N_497);
nand U3921 (N_3921,N_1417,N_1692);
nor U3922 (N_3922,N_1638,N_1575);
xor U3923 (N_3923,N_1884,N_854);
or U3924 (N_3924,N_1693,N_326);
nand U3925 (N_3925,N_643,N_936);
and U3926 (N_3926,N_56,N_483);
or U3927 (N_3927,N_1257,N_988);
xnor U3928 (N_3928,N_1552,N_179);
nand U3929 (N_3929,N_759,N_152);
nand U3930 (N_3930,N_1005,N_1529);
or U3931 (N_3931,N_672,N_1461);
xor U3932 (N_3932,N_1358,N_98);
nand U3933 (N_3933,N_1590,N_1231);
nand U3934 (N_3934,N_1071,N_705);
or U3935 (N_3935,N_1274,N_504);
nand U3936 (N_3936,N_1835,N_895);
xor U3937 (N_3937,N_1733,N_438);
nor U3938 (N_3938,N_278,N_1809);
and U3939 (N_3939,N_333,N_1551);
nor U3940 (N_3940,N_1392,N_124);
nand U3941 (N_3941,N_275,N_369);
and U3942 (N_3942,N_302,N_661);
and U3943 (N_3943,N_1227,N_1568);
or U3944 (N_3944,N_216,N_75);
or U3945 (N_3945,N_1700,N_1084);
xnor U3946 (N_3946,N_717,N_969);
nand U3947 (N_3947,N_1777,N_827);
nor U3948 (N_3948,N_972,N_913);
nor U3949 (N_3949,N_1655,N_1427);
and U3950 (N_3950,N_1140,N_629);
nand U3951 (N_3951,N_527,N_756);
nor U3952 (N_3952,N_1913,N_1161);
and U3953 (N_3953,N_191,N_919);
nand U3954 (N_3954,N_397,N_1152);
and U3955 (N_3955,N_195,N_512);
nand U3956 (N_3956,N_1882,N_1222);
xor U3957 (N_3957,N_1337,N_567);
xnor U3958 (N_3958,N_365,N_424);
nand U3959 (N_3959,N_536,N_200);
or U3960 (N_3960,N_1148,N_1091);
nor U3961 (N_3961,N_426,N_1599);
nor U3962 (N_3962,N_247,N_1010);
or U3963 (N_3963,N_501,N_618);
nand U3964 (N_3964,N_214,N_1593);
nor U3965 (N_3965,N_216,N_1180);
nand U3966 (N_3966,N_806,N_841);
nor U3967 (N_3967,N_1007,N_491);
or U3968 (N_3968,N_1067,N_262);
or U3969 (N_3969,N_487,N_51);
or U3970 (N_3970,N_683,N_1900);
nor U3971 (N_3971,N_1870,N_1472);
nand U3972 (N_3972,N_1403,N_1183);
nor U3973 (N_3973,N_1667,N_1649);
xor U3974 (N_3974,N_1768,N_1672);
and U3975 (N_3975,N_1758,N_1878);
and U3976 (N_3976,N_1294,N_921);
nand U3977 (N_3977,N_113,N_1548);
or U3978 (N_3978,N_1636,N_235);
nand U3979 (N_3979,N_833,N_1542);
nand U3980 (N_3980,N_1724,N_1007);
and U3981 (N_3981,N_1019,N_1509);
nand U3982 (N_3982,N_116,N_552);
or U3983 (N_3983,N_1861,N_1057);
xnor U3984 (N_3984,N_876,N_1424);
nand U3985 (N_3985,N_412,N_813);
nor U3986 (N_3986,N_1951,N_640);
nor U3987 (N_3987,N_1708,N_131);
and U3988 (N_3988,N_943,N_1501);
xor U3989 (N_3989,N_431,N_863);
nor U3990 (N_3990,N_861,N_1620);
or U3991 (N_3991,N_664,N_1262);
or U3992 (N_3992,N_575,N_1610);
and U3993 (N_3993,N_603,N_1439);
and U3994 (N_3994,N_687,N_171);
or U3995 (N_3995,N_31,N_1883);
nand U3996 (N_3996,N_909,N_1609);
nand U3997 (N_3997,N_1630,N_122);
nor U3998 (N_3998,N_234,N_110);
and U3999 (N_3999,N_444,N_790);
nor U4000 (N_4000,N_3935,N_3937);
nor U4001 (N_4001,N_2823,N_2438);
or U4002 (N_4002,N_3039,N_2431);
nor U4003 (N_4003,N_3148,N_3725);
nor U4004 (N_4004,N_2597,N_2721);
nand U4005 (N_4005,N_2451,N_3470);
nand U4006 (N_4006,N_3612,N_2394);
nand U4007 (N_4007,N_3628,N_2616);
nor U4008 (N_4008,N_2379,N_2334);
or U4009 (N_4009,N_2111,N_3717);
nand U4010 (N_4010,N_2571,N_2695);
nor U4011 (N_4011,N_2024,N_2020);
nand U4012 (N_4012,N_3337,N_3237);
or U4013 (N_4013,N_2951,N_3384);
xnor U4014 (N_4014,N_3995,N_3058);
nor U4015 (N_4015,N_2796,N_2391);
and U4016 (N_4016,N_3115,N_3599);
and U4017 (N_4017,N_2384,N_2849);
nor U4018 (N_4018,N_3583,N_2484);
nand U4019 (N_4019,N_3265,N_2031);
or U4020 (N_4020,N_3909,N_2270);
and U4021 (N_4021,N_3369,N_2515);
nand U4022 (N_4022,N_3704,N_2540);
or U4023 (N_4023,N_2652,N_2522);
nand U4024 (N_4024,N_3048,N_2956);
or U4025 (N_4025,N_3318,N_3363);
nand U4026 (N_4026,N_2539,N_3343);
and U4027 (N_4027,N_3138,N_3469);
and U4028 (N_4028,N_3985,N_3947);
nor U4029 (N_4029,N_2940,N_2865);
nor U4030 (N_4030,N_3050,N_3208);
and U4031 (N_4031,N_2924,N_2328);
nand U4032 (N_4032,N_2947,N_3029);
nor U4033 (N_4033,N_2308,N_2752);
nor U4034 (N_4034,N_2845,N_2694);
or U4035 (N_4035,N_3853,N_2000);
nand U4036 (N_4036,N_3094,N_2561);
nand U4037 (N_4037,N_3388,N_3394);
or U4038 (N_4038,N_3629,N_3662);
and U4039 (N_4039,N_2079,N_3681);
nand U4040 (N_4040,N_2124,N_2266);
nand U4041 (N_4041,N_3589,N_3606);
nor U4042 (N_4042,N_3547,N_2407);
or U4043 (N_4043,N_3123,N_3705);
and U4044 (N_4044,N_2567,N_3069);
nor U4045 (N_4045,N_2954,N_3723);
and U4046 (N_4046,N_2033,N_3066);
nand U4047 (N_4047,N_3251,N_2227);
or U4048 (N_4048,N_2559,N_2758);
nor U4049 (N_4049,N_2238,N_2839);
nor U4050 (N_4050,N_2130,N_2730);
xor U4051 (N_4051,N_3966,N_2224);
nand U4052 (N_4052,N_2892,N_3800);
nand U4053 (N_4053,N_3615,N_2129);
nand U4054 (N_4054,N_2433,N_3068);
nor U4055 (N_4055,N_3358,N_3676);
nand U4056 (N_4056,N_2513,N_3409);
nor U4057 (N_4057,N_3694,N_3907);
nand U4058 (N_4058,N_2263,N_2012);
and U4059 (N_4059,N_2873,N_3750);
and U4060 (N_4060,N_2076,N_3070);
or U4061 (N_4061,N_2490,N_2307);
xor U4062 (N_4062,N_2094,N_3556);
nand U4063 (N_4063,N_2991,N_3242);
and U4064 (N_4064,N_3161,N_3010);
and U4065 (N_4065,N_2166,N_3631);
nand U4066 (N_4066,N_3128,N_2576);
and U4067 (N_4067,N_3771,N_2178);
and U4068 (N_4068,N_2792,N_3552);
nand U4069 (N_4069,N_3765,N_2748);
and U4070 (N_4070,N_2747,N_3830);
nand U4071 (N_4071,N_3801,N_2342);
nand U4072 (N_4072,N_2579,N_2908);
xnor U4073 (N_4073,N_3726,N_3913);
and U4074 (N_4074,N_2929,N_2665);
and U4075 (N_4075,N_3270,N_2708);
and U4076 (N_4076,N_3527,N_3689);
xor U4077 (N_4077,N_3938,N_2642);
nand U4078 (N_4078,N_3435,N_2900);
nor U4079 (N_4079,N_2283,N_2190);
nand U4080 (N_4080,N_3001,N_2177);
xor U4081 (N_4081,N_2282,N_2572);
and U4082 (N_4082,N_2034,N_2508);
or U4083 (N_4083,N_3328,N_2054);
and U4084 (N_4084,N_3849,N_2358);
or U4085 (N_4085,N_3829,N_3183);
or U4086 (N_4086,N_2187,N_2676);
or U4087 (N_4087,N_2301,N_3045);
nand U4088 (N_4088,N_3745,N_3475);
and U4089 (N_4089,N_3756,N_2749);
and U4090 (N_4090,N_3608,N_2493);
nor U4091 (N_4091,N_3844,N_3554);
and U4092 (N_4092,N_2740,N_2882);
nand U4093 (N_4093,N_3823,N_3570);
nand U4094 (N_4094,N_2765,N_2073);
xnor U4095 (N_4095,N_2314,N_3561);
or U4096 (N_4096,N_3092,N_3049);
xnor U4097 (N_4097,N_3540,N_3669);
nand U4098 (N_4098,N_2143,N_2797);
and U4099 (N_4099,N_3223,N_2110);
nand U4100 (N_4100,N_2953,N_3036);
or U4101 (N_4101,N_3290,N_3032);
or U4102 (N_4102,N_2085,N_3284);
and U4103 (N_4103,N_2646,N_3323);
and U4104 (N_4104,N_2174,N_2896);
or U4105 (N_4105,N_3288,N_3006);
xnor U4106 (N_4106,N_3832,N_3408);
or U4107 (N_4107,N_3338,N_2296);
nor U4108 (N_4108,N_2125,N_2372);
nor U4109 (N_4109,N_3122,N_3354);
xor U4110 (N_4110,N_2338,N_2744);
and U4111 (N_4111,N_3674,N_2479);
nor U4112 (N_4112,N_3567,N_2542);
nor U4113 (N_4113,N_2527,N_2754);
nand U4114 (N_4114,N_3763,N_3432);
or U4115 (N_4115,N_3309,N_3245);
nand U4116 (N_4116,N_2557,N_2627);
and U4117 (N_4117,N_2521,N_2969);
or U4118 (N_4118,N_2414,N_3692);
xor U4119 (N_4119,N_3142,N_2586);
or U4120 (N_4120,N_3641,N_3478);
nor U4121 (N_4121,N_3645,N_2910);
and U4122 (N_4122,N_2030,N_2002);
and U4123 (N_4123,N_3194,N_3976);
nand U4124 (N_4124,N_2331,N_2306);
nor U4125 (N_4125,N_2927,N_3224);
nand U4126 (N_4126,N_2810,N_3950);
nor U4127 (N_4127,N_2353,N_3569);
nor U4128 (N_4128,N_2651,N_3956);
nand U4129 (N_4129,N_2593,N_3678);
or U4130 (N_4130,N_3220,N_3002);
or U4131 (N_4131,N_2757,N_3346);
nand U4132 (N_4132,N_3143,N_3573);
nand U4133 (N_4133,N_2339,N_2051);
and U4134 (N_4134,N_2706,N_3162);
and U4135 (N_4135,N_3706,N_3811);
or U4136 (N_4136,N_3374,N_3412);
nor U4137 (N_4137,N_3157,N_3653);
nor U4138 (N_4138,N_2047,N_3144);
nor U4139 (N_4139,N_3794,N_2984);
nor U4140 (N_4140,N_2993,N_3775);
xnor U4141 (N_4141,N_2712,N_2366);
and U4142 (N_4142,N_3939,N_2547);
nor U4143 (N_4143,N_3498,N_3904);
nor U4144 (N_4144,N_3171,N_3361);
nand U4145 (N_4145,N_2280,N_2720);
xnor U4146 (N_4146,N_3331,N_3125);
or U4147 (N_4147,N_2454,N_2141);
nor U4148 (N_4148,N_2983,N_2554);
and U4149 (N_4149,N_3846,N_2356);
and U4150 (N_4150,N_3017,N_3177);
or U4151 (N_4151,N_3656,N_2621);
nand U4152 (N_4152,N_3781,N_3444);
nor U4153 (N_4153,N_2330,N_2977);
nand U4154 (N_4154,N_2649,N_3424);
and U4155 (N_4155,N_3782,N_3366);
nor U4156 (N_4156,N_3486,N_3111);
or U4157 (N_4157,N_2221,N_3135);
or U4158 (N_4158,N_3549,N_2423);
or U4159 (N_4159,N_3287,N_3087);
or U4160 (N_4160,N_2126,N_2251);
or U4161 (N_4161,N_3633,N_3798);
or U4162 (N_4162,N_2972,N_2589);
and U4163 (N_4163,N_3562,N_3063);
xor U4164 (N_4164,N_3743,N_2894);
and U4165 (N_4165,N_3200,N_2790);
or U4166 (N_4166,N_2236,N_3344);
nor U4167 (N_4167,N_3207,N_3004);
and U4168 (N_4168,N_3665,N_2844);
nor U4169 (N_4169,N_3341,N_2297);
or U4170 (N_4170,N_2786,N_2912);
nor U4171 (N_4171,N_3682,N_3191);
and U4172 (N_4172,N_3787,N_3600);
nand U4173 (N_4173,N_2099,N_2491);
nor U4174 (N_4174,N_3821,N_3289);
nand U4175 (N_4175,N_3500,N_3490);
nor U4176 (N_4176,N_3869,N_3373);
and U4177 (N_4177,N_3840,N_3051);
or U4178 (N_4178,N_3181,N_3532);
nor U4179 (N_4179,N_3428,N_2689);
and U4180 (N_4180,N_2478,N_2520);
and U4181 (N_4181,N_3831,N_2514);
nor U4182 (N_4182,N_2602,N_3460);
nor U4183 (N_4183,N_2058,N_3738);
xnor U4184 (N_4184,N_2874,N_2210);
and U4185 (N_4185,N_3279,N_2550);
nand U4186 (N_4186,N_3429,N_2793);
or U4187 (N_4187,N_2838,N_2499);
nand U4188 (N_4188,N_3216,N_3440);
nand U4189 (N_4189,N_3580,N_3969);
nor U4190 (N_4190,N_3778,N_3586);
nor U4191 (N_4191,N_3942,N_2544);
nand U4192 (N_4192,N_3680,N_2578);
or U4193 (N_4193,N_2074,N_2973);
nand U4194 (N_4194,N_2936,N_2619);
or U4195 (N_4195,N_2794,N_3605);
nand U4196 (N_4196,N_3859,N_3843);
nor U4197 (N_4197,N_2489,N_3613);
nor U4198 (N_4198,N_2422,N_2532);
nand U4199 (N_4199,N_3134,N_3747);
nand U4200 (N_4200,N_2137,N_3847);
or U4201 (N_4201,N_2142,N_2398);
xor U4202 (N_4202,N_3483,N_3506);
and U4203 (N_4203,N_2179,N_3912);
nor U4204 (N_4204,N_3299,N_2883);
and U4205 (N_4205,N_2165,N_3089);
nor U4206 (N_4206,N_3661,N_3825);
nand U4207 (N_4207,N_2411,N_3980);
and U4208 (N_4208,N_2080,N_3176);
nor U4209 (N_4209,N_2782,N_2937);
and U4210 (N_4210,N_3292,N_2535);
xor U4211 (N_4211,N_2851,N_3215);
nand U4212 (N_4212,N_2704,N_2502);
xor U4213 (N_4213,N_2138,N_2485);
nand U4214 (N_4214,N_2727,N_2153);
or U4215 (N_4215,N_3701,N_2897);
nand U4216 (N_4216,N_3160,N_2726);
nand U4217 (N_4217,N_3232,N_3249);
nor U4218 (N_4218,N_3489,N_3783);
or U4219 (N_4219,N_2449,N_2417);
nand U4220 (N_4220,N_3766,N_2318);
and U4221 (N_4221,N_2068,N_3710);
and U4222 (N_4222,N_2987,N_2743);
xor U4223 (N_4223,N_2320,N_3112);
xnor U4224 (N_4224,N_2536,N_3577);
and U4225 (N_4225,N_2038,N_3748);
nor U4226 (N_4226,N_2390,N_2647);
nand U4227 (N_4227,N_3899,N_2787);
or U4228 (N_4228,N_3485,N_3139);
xnor U4229 (N_4229,N_3972,N_2386);
nor U4230 (N_4230,N_2467,N_3742);
or U4231 (N_4231,N_3356,N_3865);
nor U4232 (N_4232,N_3647,N_2596);
nand U4233 (N_4233,N_2531,N_2317);
and U4234 (N_4234,N_2481,N_3262);
or U4235 (N_4235,N_2397,N_2049);
and U4236 (N_4236,N_2764,N_2418);
xnor U4237 (N_4237,N_3101,N_2276);
xnor U4238 (N_4238,N_2775,N_2673);
or U4239 (N_4239,N_2121,N_3095);
or U4240 (N_4240,N_3259,N_2884);
or U4241 (N_4241,N_2488,N_2639);
nor U4242 (N_4242,N_3990,N_3534);
nor U4243 (N_4243,N_3411,N_2373);
or U4244 (N_4244,N_2088,N_3813);
nor U4245 (N_4245,N_3601,N_3377);
nor U4246 (N_4246,N_2246,N_3749);
nand U4247 (N_4247,N_2168,N_3824);
nand U4248 (N_4248,N_2990,N_3296);
and U4249 (N_4249,N_2511,N_3838);
and U4250 (N_4250,N_2768,N_2548);
or U4251 (N_4251,N_2909,N_3278);
xor U4252 (N_4252,N_3977,N_3954);
or U4253 (N_4253,N_3997,N_2473);
xor U4254 (N_4254,N_2831,N_3150);
or U4255 (N_4255,N_2256,N_2010);
xnor U4256 (N_4256,N_3400,N_2805);
or U4257 (N_4257,N_2970,N_3974);
xnor U4258 (N_4258,N_2731,N_3281);
nor U4259 (N_4259,N_3535,N_2392);
nand U4260 (N_4260,N_3735,N_3314);
nor U4261 (N_4261,N_2861,N_3121);
nor U4262 (N_4262,N_3926,N_3867);
and U4263 (N_4263,N_3229,N_2329);
nand U4264 (N_4264,N_3236,N_3462);
and U4265 (N_4265,N_2534,N_2188);
nor U4266 (N_4266,N_3650,N_2453);
nor U4267 (N_4267,N_3467,N_2582);
and U4268 (N_4268,N_2955,N_2426);
xor U4269 (N_4269,N_3131,N_3866);
or U4270 (N_4270,N_2014,N_3345);
or U4271 (N_4271,N_2237,N_2364);
nor U4272 (N_4272,N_2618,N_3779);
or U4273 (N_4273,N_2193,N_2271);
xnor U4274 (N_4274,N_3890,N_2644);
and U4275 (N_4275,N_2875,N_2591);
nand U4276 (N_4276,N_3897,N_2506);
nand U4277 (N_4277,N_3835,N_3395);
and U4278 (N_4278,N_2273,N_3352);
nand U4279 (N_4279,N_3686,N_2286);
nand U4280 (N_4280,N_2157,N_3067);
nand U4281 (N_4281,N_2517,N_3518);
nand U4282 (N_4282,N_3520,N_2498);
nor U4283 (N_4283,N_2133,N_2396);
nor U4284 (N_4284,N_3357,N_3407);
and U4285 (N_4285,N_3419,N_3714);
or U4286 (N_4286,N_3880,N_2981);
xnor U4287 (N_4287,N_3210,N_2613);
and U4288 (N_4288,N_2464,N_3514);
nor U4289 (N_4289,N_3464,N_3127);
and U4290 (N_4290,N_2938,N_3393);
or U4291 (N_4291,N_3211,N_3250);
and U4292 (N_4292,N_3713,N_3487);
and U4293 (N_4293,N_2374,N_2570);
or U4294 (N_4294,N_2029,N_3604);
nor U4295 (N_4295,N_3350,N_2189);
and U4296 (N_4296,N_2223,N_2899);
nand U4297 (N_4297,N_2204,N_3427);
and U4298 (N_4298,N_2281,N_2555);
nand U4299 (N_4299,N_3512,N_2655);
nor U4300 (N_4300,N_2413,N_2902);
nand U4301 (N_4301,N_3334,N_2208);
and U4302 (N_4302,N_3155,N_2860);
or U4303 (N_4303,N_2163,N_2581);
nand U4304 (N_4304,N_3494,N_3221);
or U4305 (N_4305,N_2641,N_3841);
nand U4306 (N_4306,N_2978,N_2738);
nor U4307 (N_4307,N_3353,N_2933);
nor U4308 (N_4308,N_3255,N_2601);
nand U4309 (N_4309,N_3075,N_2044);
nor U4310 (N_4310,N_3433,N_3884);
nand U4311 (N_4311,N_3539,N_3167);
or U4312 (N_4312,N_3437,N_3579);
and U4313 (N_4313,N_2131,N_2350);
nand U4314 (N_4314,N_2710,N_2811);
nor U4315 (N_4315,N_3180,N_3276);
and U4316 (N_4316,N_2507,N_2018);
nor U4317 (N_4317,N_3908,N_2944);
and U4318 (N_4318,N_3193,N_3568);
or U4319 (N_4319,N_2509,N_3892);
or U4320 (N_4320,N_3626,N_2160);
or U4321 (N_4321,N_2631,N_3734);
and U4322 (N_4322,N_3348,N_2199);
nor U4323 (N_4323,N_2466,N_2463);
or U4324 (N_4324,N_3504,N_2741);
and U4325 (N_4325,N_3305,N_3584);
nand U4326 (N_4326,N_2383,N_3062);
or U4327 (N_4327,N_3531,N_3870);
nor U4328 (N_4328,N_3508,N_2290);
or U4329 (N_4329,N_3189,N_2406);
nor U4330 (N_4330,N_2568,N_2592);
or U4331 (N_4331,N_3014,N_2728);
nor U4332 (N_4332,N_3637,N_2027);
nand U4333 (N_4333,N_2922,N_2798);
nor U4334 (N_4334,N_3077,N_2055);
xnor U4335 (N_4335,N_3446,N_2421);
nor U4336 (N_4336,N_2697,N_2071);
or U4337 (N_4337,N_3591,N_3286);
or U4338 (N_4338,N_2234,N_2862);
and U4339 (N_4339,N_2197,N_2346);
or U4340 (N_4340,N_3875,N_3789);
xor U4341 (N_4341,N_3248,N_3425);
nor U4342 (N_4342,N_3736,N_3226);
nor U4343 (N_4343,N_3488,N_2368);
nor U4344 (N_4344,N_3503,N_3385);
and U4345 (N_4345,N_3716,N_3080);
and U4346 (N_4346,N_2500,N_2102);
xor U4347 (N_4347,N_2715,N_2217);
and U4348 (N_4348,N_2305,N_2767);
or U4349 (N_4349,N_3773,N_2090);
or U4350 (N_4350,N_3898,N_3380);
nor U4351 (N_4351,N_2769,N_3349);
nor U4352 (N_4352,N_3760,N_3434);
and U4353 (N_4353,N_3418,N_3911);
and U4354 (N_4354,N_2745,N_2783);
or U4355 (N_4355,N_3868,N_3302);
or U4356 (N_4356,N_2455,N_3187);
and U4357 (N_4357,N_3154,N_3666);
nand U4358 (N_4358,N_2828,N_2701);
and U4359 (N_4359,N_2289,N_3261);
xor U4360 (N_4360,N_2017,N_3040);
nand U4361 (N_4361,N_2302,N_2323);
and U4362 (N_4362,N_3836,N_3240);
and U4363 (N_4363,N_2213,N_2152);
nor U4364 (N_4364,N_3513,N_2242);
or U4365 (N_4365,N_2886,N_2195);
and U4366 (N_4366,N_3313,N_3918);
and U4367 (N_4367,N_3560,N_3205);
nor U4368 (N_4368,N_3206,N_3850);
nor U4369 (N_4369,N_3673,N_2182);
nor U4370 (N_4370,N_3636,N_2470);
nand U4371 (N_4371,N_3946,N_3657);
and U4372 (N_4372,N_3619,N_2755);
or U4373 (N_4373,N_3282,N_3978);
nor U4374 (N_4374,N_2354,N_3769);
nand U4375 (N_4375,N_3225,N_3295);
nor U4376 (N_4376,N_2316,N_3493);
and U4377 (N_4377,N_2101,N_3543);
nor U4378 (N_4378,N_3355,N_2212);
nor U4379 (N_4379,N_3117,N_2594);
nand U4380 (N_4380,N_2580,N_2169);
xor U4381 (N_4381,N_3953,N_2176);
and U4382 (N_4382,N_2920,N_3671);
nand U4383 (N_4383,N_2432,N_2226);
nand U4384 (N_4384,N_2096,N_3086);
or U4385 (N_4385,N_2265,N_2659);
and U4386 (N_4386,N_2781,N_2128);
xnor U4387 (N_4387,N_2819,N_2120);
xnor U4388 (N_4388,N_2337,N_3797);
nand U4389 (N_4389,N_3492,N_3151);
nand U4390 (N_4390,N_2148,N_3209);
nor U4391 (N_4391,N_2340,N_3664);
or U4392 (N_4392,N_3479,N_2690);
and U4393 (N_4393,N_3544,N_2636);
nand U4394 (N_4394,N_3558,N_2252);
or U4395 (N_4395,N_3304,N_3963);
and U4396 (N_4396,N_3333,N_2677);
nand U4397 (N_4397,N_2834,N_3786);
xnor U4398 (N_4398,N_3529,N_2921);
and U4399 (N_4399,N_2050,N_3234);
and U4400 (N_4400,N_3199,N_2118);
nor U4401 (N_4401,N_2240,N_3815);
or U4402 (N_4402,N_3893,N_3708);
or U4403 (N_4403,N_2159,N_2988);
or U4404 (N_4404,N_2524,N_2100);
nand U4405 (N_4405,N_3021,N_2958);
nor U4406 (N_4406,N_3351,N_2942);
nor U4407 (N_4407,N_2336,N_3381);
and U4408 (N_4408,N_2553,N_2915);
nor U4409 (N_4409,N_3239,N_3575);
nor U4410 (N_4410,N_3480,N_3550);
nor U4411 (N_4411,N_3335,N_2486);
nor U4412 (N_4412,N_3536,N_2854);
or U4413 (N_4413,N_3327,N_3930);
and U4414 (N_4414,N_2004,N_3501);
nor U4415 (N_4415,N_3389,N_3889);
or U4416 (N_4416,N_2698,N_2818);
nor U4417 (N_4417,N_3597,N_3917);
nor U4418 (N_4418,N_3858,N_3695);
xor U4419 (N_4419,N_2716,N_3784);
nor U4420 (N_4420,N_3159,N_3306);
xnor U4421 (N_4421,N_3241,N_2171);
or U4422 (N_4422,N_2345,N_2083);
and U4423 (N_4423,N_3059,N_2108);
and U4424 (N_4424,N_2615,N_2809);
nand U4425 (N_4425,N_2821,N_2122);
nor U4426 (N_4426,N_2480,N_3340);
and U4427 (N_4427,N_2161,N_3301);
or U4428 (N_4428,N_3436,N_3105);
nand U4429 (N_4429,N_3962,N_2063);
xnor U4430 (N_4430,N_2737,N_3184);
nor U4431 (N_4431,N_2742,N_3056);
nand U4432 (N_4432,N_2326,N_2430);
or U4433 (N_4433,N_2905,N_2826);
xnor U4434 (N_4434,N_3874,N_2103);
nor U4435 (N_4435,N_2191,N_2344);
and U4436 (N_4436,N_2400,N_2971);
nor U4437 (N_4437,N_2232,N_2287);
or U4438 (N_4438,N_3273,N_2925);
nand U4439 (N_4439,N_3941,N_3461);
and U4440 (N_4440,N_2552,N_2228);
nor U4441 (N_4441,N_3038,N_3826);
or U4442 (N_4442,N_3640,N_2277);
nor U4443 (N_4443,N_2763,N_2370);
nand U4444 (N_4444,N_2462,N_3108);
nor U4445 (N_4445,N_3772,N_3981);
and U4446 (N_4446,N_3906,N_2249);
or U4447 (N_4447,N_3031,N_3711);
nor U4448 (N_4448,N_3891,N_2791);
nand U4449 (N_4449,N_2078,N_3510);
nor U4450 (N_4450,N_2060,N_2445);
nor U4451 (N_4451,N_2167,N_3759);
nor U4452 (N_4452,N_3398,N_2624);
nand U4453 (N_4453,N_3257,N_3940);
and U4454 (N_4454,N_2219,N_2637);
and U4455 (N_4455,N_2546,N_2812);
nor U4456 (N_4456,N_3088,N_3195);
nand U4457 (N_4457,N_3590,N_2855);
nor U4458 (N_4458,N_2222,N_3611);
and U4459 (N_4459,N_3188,N_2450);
nor U4460 (N_4460,N_3005,N_2371);
and U4461 (N_4461,N_2268,N_2220);
and U4462 (N_4462,N_2086,N_3178);
nand U4463 (N_4463,N_3602,N_3667);
and U4464 (N_4464,N_2918,N_3422);
or U4465 (N_4465,N_2603,N_3936);
or U4466 (N_4466,N_2501,N_3126);
nand U4467 (N_4467,N_3280,N_3592);
and U4468 (N_4468,N_2587,N_3572);
xor U4469 (N_4469,N_3102,N_3574);
xnor U4470 (N_4470,N_2595,N_2399);
xor U4471 (N_4471,N_2156,N_2827);
nand U4472 (N_4472,N_3753,N_2172);
nor U4473 (N_4473,N_3203,N_2065);
nand U4474 (N_4474,N_2680,N_2804);
and U4475 (N_4475,N_2471,N_3545);
nand U4476 (N_4476,N_2341,N_2492);
or U4477 (N_4477,N_2692,N_2751);
nand U4478 (N_4478,N_3015,N_3652);
nand U4479 (N_4479,N_3438,N_3103);
nand U4480 (N_4480,N_3933,N_2871);
and U4481 (N_4481,N_3857,N_2151);
nor U4482 (N_4482,N_3378,N_2869);
nand U4483 (N_4483,N_2985,N_3466);
xor U4484 (N_4484,N_3624,N_2696);
or U4485 (N_4485,N_3202,N_3679);
nor U4486 (N_4486,N_2914,N_3372);
nand U4487 (N_4487,N_3034,N_3632);
nand U4488 (N_4488,N_2401,N_3873);
nor U4489 (N_4489,N_3727,N_2906);
or U4490 (N_4490,N_2093,N_2857);
and U4491 (N_4491,N_2255,N_2952);
nand U4492 (N_4492,N_3827,N_2476);
and U4493 (N_4493,N_3228,N_2723);
nor U4494 (N_4494,N_2359,N_3523);
nor U4495 (N_4495,N_3450,N_3994);
or U4496 (N_4496,N_3916,N_3721);
or U4497 (N_4497,N_3740,N_3528);
and U4498 (N_4498,N_3767,N_3324);
or U4499 (N_4499,N_2611,N_3312);
nand U4500 (N_4500,N_3991,N_2859);
nor U4501 (N_4501,N_3011,N_3222);
nor U4502 (N_4502,N_3975,N_2201);
or U4503 (N_4503,N_3252,N_3403);
xnor U4504 (N_4504,N_2864,N_2005);
xor U4505 (N_4505,N_2046,N_2609);
nor U4506 (N_4506,N_2519,N_3960);
nand U4507 (N_4507,N_2162,N_2230);
nand U4508 (N_4508,N_2923,N_3691);
nor U4509 (N_4509,N_2117,N_2097);
nand U4510 (N_4510,N_2526,N_2904);
xor U4511 (N_4511,N_2620,N_2678);
nor U4512 (N_4512,N_3244,N_3198);
nor U4513 (N_4513,N_2687,N_2766);
or U4514 (N_4514,N_3326,N_3339);
nor U4515 (N_4515,N_3968,N_2173);
nor U4516 (N_4516,N_3799,N_3359);
nor U4517 (N_4517,N_2267,N_2408);
nor U4518 (N_4518,N_2393,N_2997);
xor U4519 (N_4519,N_3887,N_3959);
or U4520 (N_4520,N_2750,N_3635);
and U4521 (N_4521,N_3316,N_3703);
nand U4522 (N_4522,N_3082,N_2140);
or U4523 (N_4523,N_3709,N_3928);
nor U4524 (N_4524,N_2416,N_2382);
or U4525 (N_4525,N_3596,N_2975);
xor U4526 (N_4526,N_2605,N_3668);
nor U4527 (N_4527,N_3330,N_3212);
or U4528 (N_4528,N_2203,N_3165);
nand U4529 (N_4529,N_3803,N_2614);
nand U4530 (N_4530,N_2158,N_2041);
or U4531 (N_4531,N_3585,N_2759);
nor U4532 (N_4532,N_3882,N_3511);
nand U4533 (N_4533,N_2700,N_2778);
nand U4534 (N_4534,N_3920,N_2458);
and U4535 (N_4535,N_2672,N_2107);
nor U4536 (N_4536,N_2736,N_3996);
and U4537 (N_4537,N_2019,N_2935);
nand U4538 (N_4538,N_3016,N_3406);
or U4539 (N_4539,N_3246,N_3463);
or U4540 (N_4540,N_2530,N_2709);
nand U4541 (N_4541,N_2013,N_2931);
and U4542 (N_4542,N_3943,N_3320);
and U4543 (N_4543,N_3451,N_3170);
nand U4544 (N_4544,N_2734,N_3546);
nand U4545 (N_4545,N_2056,N_2069);
and U4546 (N_4546,N_3971,N_2802);
or U4547 (N_4547,N_2891,N_3683);
and U4548 (N_4548,N_2003,N_2986);
and U4549 (N_4549,N_2911,N_3620);
and U4550 (N_4550,N_3697,N_2134);
and U4551 (N_4551,N_3751,N_2939);
nand U4552 (N_4552,N_3124,N_3837);
nand U4553 (N_4553,N_2503,N_2244);
and U4554 (N_4554,N_2833,N_2439);
nand U4555 (N_4555,N_3035,N_2718);
and U4556 (N_4556,N_3308,N_2832);
or U4557 (N_4557,N_2186,N_2945);
nor U4558 (N_4558,N_3283,N_2053);
nand U4559 (N_4559,N_3507,N_3677);
and U4560 (N_4560,N_3755,N_2684);
nor U4561 (N_4561,N_3648,N_2209);
nand U4562 (N_4562,N_2551,N_2170);
or U4563 (N_4563,N_2443,N_2584);
and U4564 (N_4564,N_2444,N_2180);
nand U4565 (N_4565,N_2773,N_3700);
nor U4566 (N_4566,N_3618,N_3399);
and U4567 (N_4567,N_2881,N_2867);
xor U4568 (N_4568,N_2739,N_3864);
xnor U4569 (N_4569,N_2761,N_2693);
nor U4570 (N_4570,N_3118,N_2992);
nor U4571 (N_4571,N_3294,N_3663);
xor U4572 (N_4572,N_3116,N_3856);
and U4573 (N_4573,N_3449,N_3496);
or U4574 (N_4574,N_2682,N_2661);
and U4575 (N_4575,N_2994,N_3744);
or U4576 (N_4576,N_3214,N_2115);
nor U4577 (N_4577,N_3013,N_2043);
xor U4578 (N_4578,N_3621,N_2842);
nor U4579 (N_4579,N_2943,N_3517);
xor U4580 (N_4580,N_3888,N_3516);
or U4581 (N_4581,N_3235,N_3819);
or U4582 (N_4582,N_2147,N_3872);
or U4583 (N_4583,N_3724,N_2062);
nand U4584 (N_4584,N_2573,N_2785);
nor U4585 (N_4585,N_2123,N_2023);
or U4586 (N_4586,N_2057,N_2288);
or U4587 (N_4587,N_3563,N_2435);
xor U4588 (N_4588,N_2327,N_3163);
and U4589 (N_4589,N_3785,N_3915);
or U4590 (N_4590,N_2367,N_2119);
nor U4591 (N_4591,N_2081,N_2868);
nand U4592 (N_4592,N_3848,N_3081);
or U4593 (N_4593,N_3622,N_3322);
or U4594 (N_4594,N_2808,N_3397);
or U4595 (N_4595,N_2852,N_3047);
nor U4596 (N_4596,N_2335,N_3458);
and U4597 (N_4597,N_2089,N_3731);
nor U4598 (N_4598,N_2760,N_2622);
nand U4599 (N_4599,N_3113,N_3812);
and U4600 (N_4600,N_3401,N_3699);
nand U4601 (N_4601,N_2235,N_2007);
nor U4602 (N_4602,N_3808,N_3603);
nor U4603 (N_4603,N_3130,N_2835);
or U4604 (N_4604,N_3147,N_3670);
and U4605 (N_4605,N_2325,N_2588);
and U4606 (N_4606,N_2380,N_3256);
xnor U4607 (N_4607,N_3595,N_3442);
or U4608 (N_4608,N_2679,N_3804);
and U4609 (N_4609,N_2529,N_3790);
nand U4610 (N_4610,N_2648,N_3957);
and U4611 (N_4611,N_3643,N_2247);
nor U4612 (N_4612,N_2295,N_2516);
and U4613 (N_4613,N_3420,N_3816);
nor U4614 (N_4614,N_2009,N_2279);
nor U4615 (N_4615,N_3988,N_3277);
nor U4616 (N_4616,N_3820,N_2930);
or U4617 (N_4617,N_2025,N_3263);
nand U4618 (N_4618,N_3519,N_3137);
nor U4619 (N_4619,N_3364,N_2989);
xor U4620 (N_4620,N_2982,N_2260);
nor U4621 (N_4621,N_3325,N_3739);
and U4622 (N_4622,N_3264,N_3522);
and U4623 (N_4623,N_3445,N_2650);
nor U4624 (N_4624,N_3598,N_2885);
or U4625 (N_4625,N_3795,N_2599);
or U4626 (N_4626,N_2813,N_2770);
nand U4627 (N_4627,N_3566,N_2298);
or U4628 (N_4628,N_2623,N_2858);
nand U4629 (N_4629,N_2104,N_2893);
nor U4630 (N_4630,N_2061,N_3146);
and U4631 (N_4631,N_2437,N_2032);
xnor U4632 (N_4632,N_2574,N_2052);
nor U4633 (N_4633,N_3541,N_2713);
or U4634 (N_4634,N_2607,N_3927);
nand U4635 (N_4635,N_2686,N_3687);
or U4636 (N_4636,N_2299,N_2066);
nor U4637 (N_4637,N_3175,N_3315);
and U4638 (N_4638,N_2261,N_3423);
xor U4639 (N_4639,N_2022,N_3649);
or U4640 (N_4640,N_3862,N_2999);
or U4641 (N_4641,N_2091,N_2436);
or U4642 (N_4642,N_3022,N_3030);
xor U4643 (N_4643,N_2275,N_3533);
and U4644 (N_4644,N_3238,N_2198);
nor U4645 (N_4645,N_3053,N_3722);
or U4646 (N_4646,N_3260,N_2045);
nor U4647 (N_4647,N_2880,N_2144);
nor U4648 (N_4648,N_2976,N_3186);
nand U4649 (N_4649,N_3967,N_2816);
nor U4650 (N_4650,N_3806,N_3387);
and U4651 (N_4651,N_2565,N_2369);
and U4652 (N_4652,N_3332,N_2556);
and U4653 (N_4653,N_2113,N_3828);
nand U4654 (N_4654,N_2830,N_3061);
nor U4655 (N_4655,N_3129,N_2448);
nand U4656 (N_4656,N_2583,N_3023);
xor U4657 (N_4657,N_3481,N_3107);
or U4658 (N_4658,N_2475,N_2889);
and U4659 (N_4659,N_3140,N_2541);
nor U4660 (N_4660,N_3120,N_3109);
nand U4661 (N_4661,N_3402,N_3564);
and U4662 (N_4662,N_3233,N_2903);
xor U4663 (N_4663,N_2294,N_2001);
and U4664 (N_4664,N_3885,N_3973);
or U4665 (N_4665,N_3149,N_3055);
xnor U4666 (N_4666,N_2960,N_2333);
xor U4667 (N_4667,N_2264,N_2866);
and U4668 (N_4668,N_3730,N_3578);
nand U4669 (N_4669,N_3658,N_2324);
or U4670 (N_4670,N_3396,N_2293);
nor U4671 (N_4671,N_3020,N_3817);
nand U4672 (N_4672,N_2634,N_3525);
and U4673 (N_4673,N_3174,N_2254);
nor U4674 (N_4674,N_3833,N_3777);
nand U4675 (N_4675,N_3473,N_3097);
or U4676 (N_4676,N_2348,N_3842);
and U4677 (N_4677,N_3521,N_3054);
nand U4678 (N_4678,N_3587,N_3623);
nor U4679 (N_4679,N_3106,N_2112);
nor U4680 (N_4680,N_2347,N_3557);
nand U4681 (N_4681,N_3274,N_2668);
or U4682 (N_4682,N_2496,N_2460);
nor U4683 (N_4683,N_3718,N_2681);
xnor U4684 (N_4684,N_3415,N_3934);
nor U4685 (N_4685,N_3537,N_2207);
nand U4686 (N_4686,N_3455,N_2262);
nor U4687 (N_4687,N_3627,N_3851);
nand U4688 (N_4688,N_2312,N_2021);
nand U4689 (N_4689,N_2724,N_2890);
nor U4690 (N_4690,N_3770,N_2926);
nor U4691 (N_4691,N_2292,N_3179);
xor U4692 (N_4692,N_2657,N_3145);
nor U4693 (N_4693,N_2913,N_3201);
nor U4694 (N_4694,N_3471,N_3368);
nand U4695 (N_4695,N_2962,N_3881);
nand U4696 (N_4696,N_2533,N_3702);
nor U4697 (N_4697,N_3336,N_2035);
nor U4698 (N_4698,N_3746,N_2803);
or U4699 (N_4699,N_2806,N_3426);
or U4700 (N_4700,N_3774,N_3696);
or U4701 (N_4701,N_3267,N_3931);
and U4702 (N_4702,N_2779,N_2116);
or U4703 (N_4703,N_2457,N_2258);
nor U4704 (N_4704,N_3414,N_2585);
nand U4705 (N_4705,N_3919,N_3929);
and U4706 (N_4706,N_2538,N_3093);
nor U4707 (N_4707,N_3609,N_3878);
and U4708 (N_4708,N_2762,N_3410);
nor U4709 (N_4709,N_2964,N_2487);
or U4710 (N_4710,N_2447,N_2351);
nor U4711 (N_4711,N_3268,N_3737);
nor U4712 (N_4712,N_3948,N_3057);
or U4713 (N_4713,N_2015,N_3698);
nor U4714 (N_4714,N_3651,N_3538);
nand U4715 (N_4715,N_2837,N_2245);
or U4716 (N_4716,N_3219,N_2352);
and U4717 (N_4717,N_2456,N_3329);
nor U4718 (N_4718,N_2363,N_2420);
nor U4719 (N_4719,N_3114,N_2563);
xnor U4720 (N_4720,N_2250,N_2545);
nor U4721 (N_4721,N_2549,N_2248);
and U4722 (N_4722,N_3104,N_3675);
nand U4723 (N_4723,N_3110,N_3900);
and U4724 (N_4724,N_2196,N_2184);
or U4725 (N_4725,N_3019,N_3074);
and U4726 (N_4726,N_3788,N_2037);
nor U4727 (N_4727,N_3099,N_2241);
xor U4728 (N_4728,N_2311,N_3382);
or U4729 (N_4729,N_2375,N_3984);
or U4730 (N_4730,N_2777,N_2863);
nor U4731 (N_4731,N_3190,N_3367);
or U4732 (N_4732,N_2872,N_3298);
or U4733 (N_4733,N_2907,N_2807);
nor U4734 (N_4734,N_3253,N_2917);
xnor U4735 (N_4735,N_3342,N_3852);
xor U4736 (N_4736,N_3970,N_2528);
and U4737 (N_4737,N_2229,N_2919);
and U4738 (N_4738,N_3477,N_3404);
nand U4739 (N_4739,N_3551,N_3639);
nand U4740 (N_4740,N_3754,N_3217);
or U4741 (N_4741,N_2355,N_2664);
and U4742 (N_4742,N_2239,N_3096);
nor U4743 (N_4743,N_3213,N_2181);
nor U4744 (N_4744,N_2776,N_3555);
nor U4745 (N_4745,N_2072,N_2799);
nand U4746 (N_4746,N_2771,N_3530);
nand U4747 (N_4747,N_3565,N_3360);
nand U4748 (N_4748,N_3390,N_2378);
nand U4749 (N_4749,N_3855,N_2495);
and U4750 (N_4750,N_3453,N_2441);
or U4751 (N_4751,N_3417,N_3983);
nand U4752 (N_4752,N_2084,N_2683);
or U4753 (N_4753,N_3729,N_2663);
or U4754 (N_4754,N_2725,N_3594);
nand U4755 (N_4755,N_2036,N_3949);
or U4756 (N_4756,N_2039,N_3168);
and U4757 (N_4757,N_2575,N_3182);
nand U4758 (N_4758,N_3505,N_3474);
nand U4759 (N_4759,N_3254,N_3204);
nor U4760 (N_4760,N_2780,N_2048);
and U4761 (N_4761,N_2941,N_2155);
xor U4762 (N_4762,N_3839,N_2154);
or U4763 (N_4763,N_2477,N_2243);
and U4764 (N_4764,N_2801,N_3482);
nor U4765 (N_4765,N_2965,N_3616);
or U4766 (N_4766,N_3559,N_2825);
or U4767 (N_4767,N_3185,N_2388);
nand U4768 (N_4768,N_3439,N_2846);
xnor U4769 (N_4769,N_3998,N_2669);
nor U4770 (N_4770,N_2092,N_2164);
nand U4771 (N_4771,N_3319,N_2959);
and U4772 (N_4772,N_2274,N_2040);
nand U4773 (N_4773,N_3158,N_3169);
or U4774 (N_4774,N_2434,N_3100);
and U4775 (N_4775,N_2139,N_3310);
and U4776 (N_4776,N_2814,N_2387);
nor U4777 (N_4777,N_2026,N_2105);
xnor U4778 (N_4778,N_2772,N_3386);
xnor U4779 (N_4779,N_2175,N_2569);
nand U4780 (N_4780,N_3275,N_3042);
nand U4781 (N_4781,N_2310,N_2200);
or U4782 (N_4782,N_2381,N_3454);
and U4783 (N_4783,N_2361,N_3132);
nand U4784 (N_4784,N_3693,N_2980);
nand U4785 (N_4785,N_2674,N_3923);
and U4786 (N_4786,N_3871,N_2214);
nand U4787 (N_4787,N_3642,N_3269);
nor U4788 (N_4788,N_2878,N_2853);
nand U4789 (N_4789,N_2629,N_2042);
nor U4790 (N_4790,N_2966,N_3796);
nand U4791 (N_4791,N_2315,N_2662);
nor U4792 (N_4792,N_3625,N_3037);
nor U4793 (N_4793,N_3922,N_3728);
nand U4794 (N_4794,N_2666,N_3818);
xnor U4795 (N_4795,N_3571,N_3365);
nand U4796 (N_4796,N_2075,N_2632);
xnor U4797 (N_4797,N_2722,N_3776);
nor U4798 (N_4798,N_3073,N_2452);
and U4799 (N_4799,N_2218,N_2389);
xor U4800 (N_4800,N_2192,N_3684);
or U4801 (N_4801,N_2968,N_3231);
nor U4802 (N_4802,N_2630,N_3499);
nand U4803 (N_4803,N_3091,N_3581);
nand U4804 (N_4804,N_2577,N_2888);
nand U4805 (N_4805,N_3654,N_2127);
or U4806 (N_4806,N_2699,N_2415);
xor U4807 (N_4807,N_3076,N_3084);
or U4808 (N_4808,N_2638,N_3293);
nand U4809 (N_4809,N_2377,N_3961);
xor U4810 (N_4810,N_2349,N_3497);
or U4811 (N_4811,N_3033,N_2967);
nor U4812 (N_4812,N_2560,N_3416);
nand U4813 (N_4813,N_3227,N_3524);
and U4814 (N_4814,N_3509,N_3894);
xor U4815 (N_4815,N_3266,N_3078);
nand U4816 (N_4816,N_3441,N_2225);
and U4817 (N_4817,N_3757,N_3297);
nor U4818 (N_4818,N_3243,N_3576);
nor U4819 (N_4819,N_2961,N_3119);
xnor U4820 (N_4820,N_2656,N_3515);
nor U4821 (N_4821,N_3166,N_2658);
and U4822 (N_4822,N_2419,N_2635);
nor U4823 (N_4823,N_2895,N_2482);
and U4824 (N_4824,N_3719,N_2403);
nand U4825 (N_4825,N_2360,N_3405);
or U4826 (N_4826,N_2512,N_2675);
or U4827 (N_4827,N_3768,N_3459);
nor U4828 (N_4828,N_3003,N_2795);
nor U4829 (N_4829,N_2667,N_3247);
or U4830 (N_4830,N_2404,N_3707);
nand U4831 (N_4831,N_2928,N_2847);
and U4832 (N_4832,N_3741,N_2343);
or U4833 (N_4833,N_2183,N_3896);
or U4834 (N_4834,N_3876,N_2505);
and U4835 (N_4835,N_2332,N_2841);
and U4836 (N_4836,N_2822,N_2876);
nand U4837 (N_4837,N_2385,N_3379);
nand U4838 (N_4838,N_2610,N_3172);
or U4839 (N_4839,N_2149,N_3685);
nor U4840 (N_4840,N_3392,N_2194);
nand U4841 (N_4841,N_3472,N_2600);
nor U4842 (N_4842,N_3071,N_2815);
nor U4843 (N_4843,N_3807,N_3614);
and U4844 (N_4844,N_3271,N_2691);
and U4845 (N_4845,N_3764,N_3098);
nand U4846 (N_4846,N_3958,N_2319);
nor U4847 (N_4847,N_2459,N_3758);
and U4848 (N_4848,N_3448,N_3845);
or U4849 (N_4849,N_2537,N_2474);
or U4850 (N_4850,N_3041,N_3307);
nor U4851 (N_4851,N_2932,N_3945);
xnor U4852 (N_4852,N_2916,N_3762);
nand U4853 (N_4853,N_3732,N_2829);
nor U4854 (N_4854,N_3007,N_2472);
and U4855 (N_4855,N_2671,N_3607);
nor U4856 (N_4856,N_2497,N_3964);
nor U4857 (N_4857,N_2109,N_2711);
nor U4858 (N_4858,N_3311,N_3834);
nand U4859 (N_4859,N_3921,N_2259);
nand U4860 (N_4860,N_3009,N_2850);
nor U4861 (N_4861,N_2257,N_3476);
or U4862 (N_4862,N_3982,N_2402);
xnor U4863 (N_4863,N_2843,N_2523);
nand U4864 (N_4864,N_2685,N_3672);
nor U4865 (N_4865,N_2995,N_3905);
nor U4866 (N_4866,N_3452,N_2948);
or U4867 (N_4867,N_3258,N_3362);
and U4868 (N_4868,N_2558,N_2395);
xnor U4869 (N_4869,N_2285,N_2145);
nor U4870 (N_4870,N_3027,N_3375);
and U4871 (N_4871,N_2114,N_2284);
nand U4872 (N_4872,N_2185,N_3993);
or U4873 (N_4873,N_2461,N_2410);
nor U4874 (N_4874,N_3914,N_2640);
nand U4875 (N_4875,N_3951,N_3761);
nand U4876 (N_4876,N_3814,N_2707);
and U4877 (N_4877,N_2705,N_2836);
nand U4878 (N_4878,N_3863,N_3955);
xnor U4879 (N_4879,N_2996,N_3376);
or U4880 (N_4880,N_2465,N_2082);
and U4881 (N_4881,N_2028,N_3924);
nor U4882 (N_4882,N_2653,N_3457);
and U4883 (N_4883,N_2132,N_2077);
nor U4884 (N_4884,N_2136,N_2934);
nand U4885 (N_4885,N_3317,N_3072);
or U4886 (N_4886,N_3456,N_2059);
nor U4887 (N_4887,N_3925,N_3979);
and U4888 (N_4888,N_2946,N_3822);
and U4889 (N_4889,N_2717,N_2733);
nor U4890 (N_4890,N_2562,N_3291);
nor U4891 (N_4891,N_3421,N_2309);
and U4892 (N_4892,N_2719,N_2703);
xnor U4893 (N_4893,N_2446,N_2714);
and U4894 (N_4894,N_2625,N_2688);
nor U4895 (N_4895,N_3164,N_2963);
and U4896 (N_4896,N_2362,N_2322);
and U4897 (N_4897,N_2321,N_2409);
nand U4898 (N_4898,N_2800,N_2784);
nor U4899 (N_4899,N_2064,N_3085);
xnor U4900 (N_4900,N_2564,N_2291);
nor U4901 (N_4901,N_3443,N_2098);
xor U4902 (N_4902,N_2879,N_2278);
xor U4903 (N_4903,N_3447,N_3079);
nor U4904 (N_4904,N_3197,N_3371);
nand U4905 (N_4905,N_3655,N_2215);
xor U4906 (N_4906,N_2702,N_2146);
nor U4907 (N_4907,N_3688,N_3141);
xnor U4908 (N_4908,N_3430,N_3230);
nor U4909 (N_4909,N_3646,N_3192);
nor U4910 (N_4910,N_2654,N_2405);
or U4911 (N_4911,N_2626,N_3465);
xor U4912 (N_4912,N_3046,N_2817);
nand U4913 (N_4913,N_3877,N_2483);
xnor U4914 (N_4914,N_2856,N_2300);
nand U4915 (N_4915,N_3660,N_3965);
nand U4916 (N_4916,N_2211,N_2606);
or U4917 (N_4917,N_3391,N_3901);
nand U4918 (N_4918,N_3752,N_2365);
nand U4919 (N_4919,N_3659,N_3638);
or U4920 (N_4920,N_2735,N_3495);
nand U4921 (N_4921,N_2898,N_2788);
nor U4922 (N_4922,N_2608,N_2412);
xnor U4923 (N_4923,N_3883,N_2440);
and U4924 (N_4924,N_3321,N_2011);
nand U4925 (N_4925,N_3952,N_2643);
or U4926 (N_4926,N_2135,N_2231);
or U4927 (N_4927,N_3588,N_2566);
nand U4928 (N_4928,N_2006,N_3526);
and U4929 (N_4929,N_3895,N_2670);
or U4930 (N_4930,N_3690,N_2303);
and U4931 (N_4931,N_2233,N_2205);
or U4932 (N_4932,N_3548,N_2753);
and U4933 (N_4933,N_2660,N_3024);
nand U4934 (N_4934,N_3012,N_2598);
or U4935 (N_4935,N_3156,N_2016);
or U4936 (N_4936,N_2425,N_3065);
nor U4937 (N_4937,N_3854,N_2840);
or U4938 (N_4938,N_2617,N_2518);
xnor U4939 (N_4939,N_3932,N_3987);
nand U4940 (N_4940,N_3593,N_3903);
nor U4941 (N_4941,N_2628,N_3044);
xnor U4942 (N_4942,N_3792,N_2732);
or U4943 (N_4943,N_3431,N_2087);
and U4944 (N_4944,N_3989,N_3793);
nor U4945 (N_4945,N_2216,N_2202);
nand U4946 (N_4946,N_2424,N_2095);
and U4947 (N_4947,N_2427,N_2067);
or U4948 (N_4948,N_3153,N_3944);
nand U4949 (N_4949,N_3791,N_3630);
and U4950 (N_4950,N_3644,N_3720);
nand U4951 (N_4951,N_2789,N_3553);
nand U4952 (N_4952,N_3000,N_3902);
and U4953 (N_4953,N_3152,N_2901);
nor U4954 (N_4954,N_3383,N_2974);
nor U4955 (N_4955,N_2645,N_3025);
or U4956 (N_4956,N_2313,N_3018);
nor U4957 (N_4957,N_2253,N_3303);
or U4958 (N_4958,N_2612,N_2870);
and U4959 (N_4959,N_3468,N_3173);
xnor U4960 (N_4960,N_3413,N_2824);
xor U4961 (N_4961,N_3285,N_2206);
nand U4962 (N_4962,N_2494,N_2304);
nand U4963 (N_4963,N_3491,N_2269);
nand U4964 (N_4964,N_2428,N_3060);
nor U4965 (N_4965,N_3043,N_3218);
nand U4966 (N_4966,N_3999,N_2070);
or U4967 (N_4967,N_2504,N_2998);
nor U4968 (N_4968,N_2957,N_3370);
nor U4969 (N_4969,N_3026,N_3028);
and U4970 (N_4970,N_2950,N_3810);
and U4971 (N_4971,N_3542,N_2543);
xnor U4972 (N_4972,N_3805,N_3008);
and U4973 (N_4973,N_3617,N_3780);
and U4974 (N_4974,N_3733,N_3083);
or U4975 (N_4975,N_2887,N_3136);
xor U4976 (N_4976,N_3886,N_3582);
nand U4977 (N_4977,N_3992,N_3090);
nand U4978 (N_4978,N_2949,N_3064);
nor U4979 (N_4979,N_2376,N_3802);
nor U4980 (N_4980,N_3484,N_2877);
nand U4981 (N_4981,N_3133,N_2633);
nand U4982 (N_4982,N_3910,N_3272);
and U4983 (N_4983,N_3634,N_3715);
and U4984 (N_4984,N_2469,N_2442);
nand U4985 (N_4985,N_2468,N_3712);
and U4986 (N_4986,N_2272,N_3196);
and U4987 (N_4987,N_2604,N_2150);
and U4988 (N_4988,N_2848,N_2357);
or U4989 (N_4989,N_2106,N_2525);
or U4990 (N_4990,N_2774,N_3860);
nor U4991 (N_4991,N_3986,N_2729);
nand U4992 (N_4992,N_2746,N_3610);
or U4993 (N_4993,N_2820,N_3052);
nor U4994 (N_4994,N_2429,N_2756);
or U4995 (N_4995,N_2590,N_3809);
or U4996 (N_4996,N_3347,N_2008);
and U4997 (N_4997,N_3502,N_3879);
nor U4998 (N_4998,N_3861,N_2979);
nand U4999 (N_4999,N_2510,N_3300);
nor U5000 (N_5000,N_3142,N_2703);
or U5001 (N_5001,N_3147,N_3032);
nor U5002 (N_5002,N_2067,N_3079);
nand U5003 (N_5003,N_3979,N_3117);
and U5004 (N_5004,N_3437,N_2009);
nand U5005 (N_5005,N_2573,N_3980);
nand U5006 (N_5006,N_3445,N_3600);
and U5007 (N_5007,N_2095,N_2006);
nand U5008 (N_5008,N_2090,N_2558);
nor U5009 (N_5009,N_3562,N_2677);
nor U5010 (N_5010,N_2497,N_2772);
and U5011 (N_5011,N_2820,N_2224);
nor U5012 (N_5012,N_2490,N_3922);
nand U5013 (N_5013,N_3375,N_3012);
nand U5014 (N_5014,N_3438,N_3756);
and U5015 (N_5015,N_2772,N_3396);
nor U5016 (N_5016,N_2613,N_2889);
or U5017 (N_5017,N_3022,N_3792);
and U5018 (N_5018,N_2680,N_3324);
nor U5019 (N_5019,N_2891,N_3592);
nor U5020 (N_5020,N_2421,N_3162);
nand U5021 (N_5021,N_2319,N_3388);
or U5022 (N_5022,N_3265,N_3592);
nor U5023 (N_5023,N_2420,N_2850);
nand U5024 (N_5024,N_3019,N_3460);
or U5025 (N_5025,N_2124,N_2676);
or U5026 (N_5026,N_3974,N_3765);
or U5027 (N_5027,N_2207,N_3191);
nand U5028 (N_5028,N_2893,N_2725);
nor U5029 (N_5029,N_3313,N_2018);
and U5030 (N_5030,N_2258,N_3358);
or U5031 (N_5031,N_3004,N_3640);
or U5032 (N_5032,N_2026,N_2403);
or U5033 (N_5033,N_2609,N_2955);
xnor U5034 (N_5034,N_2194,N_3956);
or U5035 (N_5035,N_3969,N_3306);
and U5036 (N_5036,N_3398,N_2983);
and U5037 (N_5037,N_3620,N_2074);
or U5038 (N_5038,N_2931,N_2608);
and U5039 (N_5039,N_3120,N_2685);
nand U5040 (N_5040,N_3750,N_3850);
nand U5041 (N_5041,N_3338,N_2705);
nand U5042 (N_5042,N_2014,N_2573);
nor U5043 (N_5043,N_3995,N_3575);
or U5044 (N_5044,N_2937,N_2069);
and U5045 (N_5045,N_3438,N_3684);
or U5046 (N_5046,N_2037,N_2520);
or U5047 (N_5047,N_3724,N_2556);
or U5048 (N_5048,N_2432,N_2957);
nand U5049 (N_5049,N_2847,N_3578);
or U5050 (N_5050,N_3559,N_2939);
and U5051 (N_5051,N_3550,N_2569);
nor U5052 (N_5052,N_2181,N_3230);
or U5053 (N_5053,N_2740,N_2035);
nand U5054 (N_5054,N_3884,N_2498);
and U5055 (N_5055,N_3409,N_2913);
nand U5056 (N_5056,N_3494,N_2699);
xor U5057 (N_5057,N_2225,N_2889);
xnor U5058 (N_5058,N_2738,N_2500);
nor U5059 (N_5059,N_2779,N_3267);
and U5060 (N_5060,N_2504,N_2421);
or U5061 (N_5061,N_2909,N_2322);
and U5062 (N_5062,N_2538,N_3935);
or U5063 (N_5063,N_3269,N_2642);
or U5064 (N_5064,N_2040,N_2879);
nand U5065 (N_5065,N_3070,N_2459);
and U5066 (N_5066,N_2138,N_2060);
or U5067 (N_5067,N_3389,N_2809);
nand U5068 (N_5068,N_3034,N_3755);
xnor U5069 (N_5069,N_3004,N_3487);
nor U5070 (N_5070,N_2225,N_2147);
or U5071 (N_5071,N_3160,N_2412);
or U5072 (N_5072,N_3999,N_2260);
xnor U5073 (N_5073,N_3730,N_3687);
nand U5074 (N_5074,N_3374,N_2097);
nand U5075 (N_5075,N_2949,N_3897);
and U5076 (N_5076,N_3130,N_3774);
or U5077 (N_5077,N_2797,N_3643);
or U5078 (N_5078,N_3186,N_2099);
or U5079 (N_5079,N_3216,N_3776);
nand U5080 (N_5080,N_2732,N_3789);
or U5081 (N_5081,N_2430,N_2288);
nor U5082 (N_5082,N_2765,N_3471);
nand U5083 (N_5083,N_2635,N_2329);
nor U5084 (N_5084,N_2341,N_2887);
and U5085 (N_5085,N_2751,N_3842);
nand U5086 (N_5086,N_2888,N_2557);
nand U5087 (N_5087,N_2375,N_2703);
xor U5088 (N_5088,N_2052,N_3939);
or U5089 (N_5089,N_2427,N_3692);
and U5090 (N_5090,N_2519,N_3903);
xor U5091 (N_5091,N_3612,N_2093);
or U5092 (N_5092,N_3647,N_2205);
or U5093 (N_5093,N_2723,N_2107);
xnor U5094 (N_5094,N_2190,N_3866);
nor U5095 (N_5095,N_2909,N_2410);
or U5096 (N_5096,N_2521,N_2819);
and U5097 (N_5097,N_3012,N_2954);
xor U5098 (N_5098,N_2016,N_2608);
nor U5099 (N_5099,N_2003,N_2846);
nand U5100 (N_5100,N_3162,N_2592);
and U5101 (N_5101,N_2645,N_2881);
or U5102 (N_5102,N_2983,N_3249);
nand U5103 (N_5103,N_2048,N_3179);
nor U5104 (N_5104,N_2876,N_2184);
nand U5105 (N_5105,N_3068,N_2195);
nor U5106 (N_5106,N_3919,N_2255);
nand U5107 (N_5107,N_3042,N_3664);
or U5108 (N_5108,N_3433,N_3275);
or U5109 (N_5109,N_2354,N_3653);
or U5110 (N_5110,N_3631,N_3963);
or U5111 (N_5111,N_3491,N_2356);
and U5112 (N_5112,N_3649,N_2912);
or U5113 (N_5113,N_3357,N_2476);
nand U5114 (N_5114,N_3181,N_3192);
or U5115 (N_5115,N_3257,N_3148);
and U5116 (N_5116,N_2967,N_3626);
xor U5117 (N_5117,N_2181,N_3650);
nor U5118 (N_5118,N_3554,N_3616);
or U5119 (N_5119,N_3604,N_2940);
nor U5120 (N_5120,N_3451,N_3056);
or U5121 (N_5121,N_2319,N_3686);
xnor U5122 (N_5122,N_3125,N_3409);
and U5123 (N_5123,N_3224,N_2685);
nor U5124 (N_5124,N_3504,N_3653);
nor U5125 (N_5125,N_3434,N_3577);
and U5126 (N_5126,N_3561,N_2150);
nor U5127 (N_5127,N_2553,N_2095);
nor U5128 (N_5128,N_3832,N_2109);
and U5129 (N_5129,N_3975,N_2429);
or U5130 (N_5130,N_3706,N_2769);
and U5131 (N_5131,N_2496,N_3233);
nand U5132 (N_5132,N_3019,N_2509);
xnor U5133 (N_5133,N_3045,N_2815);
xnor U5134 (N_5134,N_3283,N_2929);
nand U5135 (N_5135,N_2341,N_3299);
and U5136 (N_5136,N_3282,N_3134);
xnor U5137 (N_5137,N_3992,N_3715);
and U5138 (N_5138,N_2573,N_3557);
and U5139 (N_5139,N_2170,N_2619);
or U5140 (N_5140,N_2877,N_3146);
and U5141 (N_5141,N_3646,N_3606);
nand U5142 (N_5142,N_2020,N_3216);
nand U5143 (N_5143,N_3663,N_3371);
or U5144 (N_5144,N_2756,N_2349);
or U5145 (N_5145,N_2732,N_3834);
or U5146 (N_5146,N_2341,N_3439);
nor U5147 (N_5147,N_2085,N_3496);
nand U5148 (N_5148,N_3264,N_3969);
nor U5149 (N_5149,N_3518,N_2010);
xnor U5150 (N_5150,N_2869,N_3193);
nor U5151 (N_5151,N_2331,N_3243);
or U5152 (N_5152,N_2160,N_3704);
and U5153 (N_5153,N_2482,N_3480);
or U5154 (N_5154,N_3304,N_2570);
nand U5155 (N_5155,N_2485,N_2897);
and U5156 (N_5156,N_3027,N_2016);
and U5157 (N_5157,N_3950,N_3250);
and U5158 (N_5158,N_2268,N_3621);
or U5159 (N_5159,N_2804,N_3634);
xnor U5160 (N_5160,N_3177,N_3725);
and U5161 (N_5161,N_2290,N_3693);
or U5162 (N_5162,N_3926,N_2011);
nor U5163 (N_5163,N_3480,N_2928);
nand U5164 (N_5164,N_3040,N_3671);
nand U5165 (N_5165,N_3169,N_3763);
or U5166 (N_5166,N_3218,N_2344);
or U5167 (N_5167,N_2222,N_3838);
and U5168 (N_5168,N_2224,N_2918);
nor U5169 (N_5169,N_2785,N_3724);
and U5170 (N_5170,N_3501,N_3676);
and U5171 (N_5171,N_2098,N_2998);
or U5172 (N_5172,N_3219,N_3906);
or U5173 (N_5173,N_2425,N_3129);
nand U5174 (N_5174,N_3473,N_2951);
and U5175 (N_5175,N_2897,N_2532);
xor U5176 (N_5176,N_2796,N_2904);
nor U5177 (N_5177,N_2263,N_2551);
nor U5178 (N_5178,N_3448,N_3843);
nand U5179 (N_5179,N_2111,N_2892);
xnor U5180 (N_5180,N_3098,N_3430);
or U5181 (N_5181,N_2004,N_2802);
nand U5182 (N_5182,N_2113,N_2469);
xnor U5183 (N_5183,N_2791,N_2784);
xor U5184 (N_5184,N_3489,N_3279);
nand U5185 (N_5185,N_2229,N_3378);
xor U5186 (N_5186,N_2076,N_2539);
and U5187 (N_5187,N_2363,N_2368);
and U5188 (N_5188,N_2327,N_2369);
and U5189 (N_5189,N_2405,N_3918);
nand U5190 (N_5190,N_3065,N_3257);
nor U5191 (N_5191,N_3556,N_3179);
nand U5192 (N_5192,N_2382,N_2484);
and U5193 (N_5193,N_3349,N_3546);
nor U5194 (N_5194,N_3487,N_2664);
or U5195 (N_5195,N_2865,N_2066);
xnor U5196 (N_5196,N_2581,N_3421);
nor U5197 (N_5197,N_3749,N_3414);
nor U5198 (N_5198,N_3922,N_2969);
and U5199 (N_5199,N_3409,N_2501);
nor U5200 (N_5200,N_3970,N_3932);
or U5201 (N_5201,N_3297,N_3729);
xor U5202 (N_5202,N_2209,N_2777);
and U5203 (N_5203,N_2465,N_2583);
or U5204 (N_5204,N_2053,N_2125);
or U5205 (N_5205,N_3329,N_3896);
nor U5206 (N_5206,N_3808,N_2102);
or U5207 (N_5207,N_3846,N_3281);
or U5208 (N_5208,N_3653,N_3300);
and U5209 (N_5209,N_3595,N_3734);
nor U5210 (N_5210,N_2654,N_3698);
xor U5211 (N_5211,N_2728,N_2440);
xnor U5212 (N_5212,N_2208,N_2220);
and U5213 (N_5213,N_3232,N_2927);
or U5214 (N_5214,N_3201,N_3799);
nor U5215 (N_5215,N_3842,N_2896);
or U5216 (N_5216,N_2871,N_2003);
and U5217 (N_5217,N_2306,N_3412);
or U5218 (N_5218,N_2687,N_2396);
xor U5219 (N_5219,N_3373,N_2550);
xor U5220 (N_5220,N_3416,N_2625);
nor U5221 (N_5221,N_2510,N_3332);
nand U5222 (N_5222,N_2207,N_3459);
nor U5223 (N_5223,N_3597,N_3555);
nand U5224 (N_5224,N_2949,N_3559);
nor U5225 (N_5225,N_3667,N_2398);
and U5226 (N_5226,N_3337,N_3642);
or U5227 (N_5227,N_3793,N_2922);
and U5228 (N_5228,N_2317,N_3921);
xnor U5229 (N_5229,N_3305,N_3910);
xnor U5230 (N_5230,N_3358,N_3103);
and U5231 (N_5231,N_3317,N_2558);
nor U5232 (N_5232,N_2829,N_3773);
nor U5233 (N_5233,N_3260,N_2042);
nand U5234 (N_5234,N_2250,N_2666);
nand U5235 (N_5235,N_3753,N_3138);
nor U5236 (N_5236,N_2925,N_2220);
nand U5237 (N_5237,N_3803,N_2542);
nand U5238 (N_5238,N_2964,N_3230);
nand U5239 (N_5239,N_3379,N_2904);
nand U5240 (N_5240,N_2114,N_3803);
nand U5241 (N_5241,N_2183,N_2523);
and U5242 (N_5242,N_2075,N_3339);
nand U5243 (N_5243,N_2496,N_3427);
xnor U5244 (N_5244,N_2094,N_2069);
nor U5245 (N_5245,N_2885,N_3232);
nand U5246 (N_5246,N_3214,N_2565);
nor U5247 (N_5247,N_2986,N_3138);
and U5248 (N_5248,N_2616,N_3393);
or U5249 (N_5249,N_3633,N_2982);
or U5250 (N_5250,N_3408,N_2058);
nor U5251 (N_5251,N_3336,N_2701);
nand U5252 (N_5252,N_2494,N_3220);
nor U5253 (N_5253,N_3537,N_3165);
nor U5254 (N_5254,N_3694,N_3584);
xnor U5255 (N_5255,N_3189,N_3519);
nor U5256 (N_5256,N_2223,N_3678);
nand U5257 (N_5257,N_2627,N_3231);
xor U5258 (N_5258,N_2383,N_2961);
nand U5259 (N_5259,N_3774,N_3358);
or U5260 (N_5260,N_2448,N_3383);
or U5261 (N_5261,N_2276,N_3568);
xor U5262 (N_5262,N_2795,N_3416);
and U5263 (N_5263,N_2514,N_2534);
xnor U5264 (N_5264,N_3351,N_3031);
nand U5265 (N_5265,N_3725,N_3174);
nor U5266 (N_5266,N_3070,N_3266);
nand U5267 (N_5267,N_2083,N_3840);
and U5268 (N_5268,N_3454,N_3066);
and U5269 (N_5269,N_2577,N_3599);
and U5270 (N_5270,N_3736,N_2713);
nand U5271 (N_5271,N_3669,N_3248);
nor U5272 (N_5272,N_2043,N_3893);
nor U5273 (N_5273,N_3679,N_2218);
and U5274 (N_5274,N_2538,N_3979);
or U5275 (N_5275,N_2853,N_2902);
or U5276 (N_5276,N_2992,N_3035);
nand U5277 (N_5277,N_2333,N_2574);
xnor U5278 (N_5278,N_2354,N_2629);
and U5279 (N_5279,N_2985,N_3377);
nand U5280 (N_5280,N_3851,N_3296);
nand U5281 (N_5281,N_3770,N_2071);
nor U5282 (N_5282,N_2880,N_2694);
and U5283 (N_5283,N_2538,N_3675);
nand U5284 (N_5284,N_2643,N_3270);
or U5285 (N_5285,N_3510,N_2482);
nor U5286 (N_5286,N_3800,N_2287);
nor U5287 (N_5287,N_2165,N_2785);
or U5288 (N_5288,N_3273,N_2938);
nand U5289 (N_5289,N_3224,N_2282);
nor U5290 (N_5290,N_3806,N_3652);
nor U5291 (N_5291,N_2663,N_3604);
and U5292 (N_5292,N_3776,N_3540);
nand U5293 (N_5293,N_2370,N_2938);
or U5294 (N_5294,N_3560,N_2564);
or U5295 (N_5295,N_2368,N_3189);
and U5296 (N_5296,N_2365,N_3543);
or U5297 (N_5297,N_2623,N_3732);
nor U5298 (N_5298,N_3966,N_2978);
and U5299 (N_5299,N_3400,N_3934);
xnor U5300 (N_5300,N_2646,N_2895);
and U5301 (N_5301,N_2815,N_3042);
nand U5302 (N_5302,N_3658,N_2091);
or U5303 (N_5303,N_2859,N_2034);
and U5304 (N_5304,N_3498,N_2953);
xor U5305 (N_5305,N_3563,N_2338);
nor U5306 (N_5306,N_3451,N_3075);
xor U5307 (N_5307,N_2975,N_3558);
nand U5308 (N_5308,N_2941,N_3826);
nand U5309 (N_5309,N_2475,N_2109);
nor U5310 (N_5310,N_2911,N_3172);
or U5311 (N_5311,N_2336,N_3672);
nor U5312 (N_5312,N_2848,N_2816);
nor U5313 (N_5313,N_3577,N_2747);
nor U5314 (N_5314,N_2462,N_3250);
nor U5315 (N_5315,N_2301,N_3719);
nand U5316 (N_5316,N_2562,N_2828);
nor U5317 (N_5317,N_2502,N_3601);
and U5318 (N_5318,N_3975,N_3841);
or U5319 (N_5319,N_2175,N_2173);
or U5320 (N_5320,N_3770,N_2773);
or U5321 (N_5321,N_3341,N_2888);
nor U5322 (N_5322,N_3849,N_3384);
or U5323 (N_5323,N_2198,N_3227);
and U5324 (N_5324,N_2772,N_3304);
nor U5325 (N_5325,N_2289,N_2158);
and U5326 (N_5326,N_3072,N_3265);
nand U5327 (N_5327,N_3601,N_3457);
or U5328 (N_5328,N_3836,N_2365);
or U5329 (N_5329,N_3377,N_3044);
nor U5330 (N_5330,N_2626,N_2622);
and U5331 (N_5331,N_2688,N_2376);
or U5332 (N_5332,N_3052,N_2082);
and U5333 (N_5333,N_3697,N_3623);
or U5334 (N_5334,N_3004,N_3185);
and U5335 (N_5335,N_3884,N_3928);
and U5336 (N_5336,N_2523,N_2295);
or U5337 (N_5337,N_3385,N_2894);
or U5338 (N_5338,N_3763,N_2549);
and U5339 (N_5339,N_3569,N_3069);
nand U5340 (N_5340,N_3464,N_2669);
nor U5341 (N_5341,N_2425,N_3651);
nand U5342 (N_5342,N_3046,N_2536);
or U5343 (N_5343,N_3904,N_2116);
or U5344 (N_5344,N_3283,N_3846);
and U5345 (N_5345,N_3918,N_2966);
or U5346 (N_5346,N_2055,N_3608);
xnor U5347 (N_5347,N_3519,N_3734);
nor U5348 (N_5348,N_2142,N_2621);
nand U5349 (N_5349,N_2834,N_2258);
nor U5350 (N_5350,N_3038,N_3096);
nand U5351 (N_5351,N_3012,N_2462);
or U5352 (N_5352,N_3680,N_2698);
nor U5353 (N_5353,N_2614,N_2155);
nand U5354 (N_5354,N_2727,N_3693);
and U5355 (N_5355,N_2658,N_2963);
and U5356 (N_5356,N_3904,N_2255);
and U5357 (N_5357,N_3878,N_3923);
and U5358 (N_5358,N_3046,N_3099);
nand U5359 (N_5359,N_2572,N_2907);
nand U5360 (N_5360,N_2809,N_3972);
nor U5361 (N_5361,N_2353,N_3072);
nand U5362 (N_5362,N_3818,N_3075);
or U5363 (N_5363,N_2500,N_2468);
and U5364 (N_5364,N_3166,N_2298);
and U5365 (N_5365,N_2596,N_3042);
or U5366 (N_5366,N_2552,N_3365);
and U5367 (N_5367,N_3553,N_3947);
nor U5368 (N_5368,N_3590,N_2166);
and U5369 (N_5369,N_2937,N_2151);
nand U5370 (N_5370,N_3180,N_2979);
or U5371 (N_5371,N_3715,N_2875);
nor U5372 (N_5372,N_3742,N_3743);
nor U5373 (N_5373,N_2054,N_3994);
nor U5374 (N_5374,N_3489,N_3933);
or U5375 (N_5375,N_2389,N_3506);
or U5376 (N_5376,N_2329,N_3014);
nand U5377 (N_5377,N_3525,N_3947);
or U5378 (N_5378,N_2369,N_3864);
or U5379 (N_5379,N_2682,N_3335);
nand U5380 (N_5380,N_2771,N_2744);
nand U5381 (N_5381,N_2050,N_3882);
or U5382 (N_5382,N_2470,N_2056);
and U5383 (N_5383,N_3729,N_3953);
and U5384 (N_5384,N_3149,N_3260);
or U5385 (N_5385,N_3659,N_2788);
nor U5386 (N_5386,N_3670,N_3811);
or U5387 (N_5387,N_3922,N_2691);
or U5388 (N_5388,N_3525,N_2401);
and U5389 (N_5389,N_3896,N_3531);
nand U5390 (N_5390,N_3422,N_2497);
and U5391 (N_5391,N_3443,N_2643);
nor U5392 (N_5392,N_2126,N_2637);
xnor U5393 (N_5393,N_3240,N_2848);
or U5394 (N_5394,N_3514,N_3942);
nor U5395 (N_5395,N_2953,N_3239);
or U5396 (N_5396,N_3267,N_3061);
nand U5397 (N_5397,N_3476,N_3138);
or U5398 (N_5398,N_3225,N_2051);
nand U5399 (N_5399,N_2724,N_3216);
nor U5400 (N_5400,N_3247,N_3252);
nor U5401 (N_5401,N_2931,N_2552);
nand U5402 (N_5402,N_2557,N_2236);
or U5403 (N_5403,N_3476,N_3686);
and U5404 (N_5404,N_3220,N_2188);
and U5405 (N_5405,N_3955,N_2099);
and U5406 (N_5406,N_2587,N_3163);
and U5407 (N_5407,N_2309,N_2082);
and U5408 (N_5408,N_3879,N_2714);
and U5409 (N_5409,N_3906,N_3873);
nor U5410 (N_5410,N_3793,N_3307);
and U5411 (N_5411,N_2641,N_2703);
nand U5412 (N_5412,N_2368,N_2277);
and U5413 (N_5413,N_2949,N_3294);
and U5414 (N_5414,N_3132,N_2194);
nor U5415 (N_5415,N_3602,N_3181);
or U5416 (N_5416,N_2341,N_2506);
xnor U5417 (N_5417,N_3776,N_2571);
or U5418 (N_5418,N_2052,N_3467);
or U5419 (N_5419,N_3771,N_3827);
and U5420 (N_5420,N_3598,N_2005);
or U5421 (N_5421,N_2336,N_3729);
or U5422 (N_5422,N_2460,N_3936);
or U5423 (N_5423,N_3985,N_2408);
and U5424 (N_5424,N_2635,N_3029);
or U5425 (N_5425,N_2795,N_2488);
nand U5426 (N_5426,N_3411,N_3638);
nand U5427 (N_5427,N_3139,N_2666);
or U5428 (N_5428,N_2293,N_3830);
or U5429 (N_5429,N_3404,N_3191);
or U5430 (N_5430,N_2827,N_2626);
nor U5431 (N_5431,N_3281,N_3278);
or U5432 (N_5432,N_3885,N_3952);
xor U5433 (N_5433,N_3999,N_2419);
xnor U5434 (N_5434,N_2161,N_3656);
and U5435 (N_5435,N_2447,N_2571);
nand U5436 (N_5436,N_3390,N_3950);
xor U5437 (N_5437,N_2078,N_3141);
or U5438 (N_5438,N_3896,N_2768);
or U5439 (N_5439,N_3947,N_3458);
or U5440 (N_5440,N_2071,N_3267);
nor U5441 (N_5441,N_3706,N_2293);
and U5442 (N_5442,N_2404,N_3872);
and U5443 (N_5443,N_3676,N_3652);
nor U5444 (N_5444,N_2226,N_2812);
and U5445 (N_5445,N_3188,N_3394);
and U5446 (N_5446,N_2046,N_3956);
nor U5447 (N_5447,N_2570,N_3182);
and U5448 (N_5448,N_2295,N_3072);
and U5449 (N_5449,N_2938,N_2743);
nand U5450 (N_5450,N_2730,N_2235);
or U5451 (N_5451,N_3489,N_2647);
nand U5452 (N_5452,N_3497,N_2667);
or U5453 (N_5453,N_3728,N_3629);
nor U5454 (N_5454,N_2790,N_2605);
xor U5455 (N_5455,N_2754,N_2844);
and U5456 (N_5456,N_3301,N_3793);
nand U5457 (N_5457,N_2555,N_2141);
nor U5458 (N_5458,N_3481,N_3684);
xor U5459 (N_5459,N_3687,N_2964);
nand U5460 (N_5460,N_3274,N_2680);
xnor U5461 (N_5461,N_3081,N_3572);
or U5462 (N_5462,N_3583,N_2956);
nand U5463 (N_5463,N_3239,N_2409);
and U5464 (N_5464,N_3316,N_3577);
nand U5465 (N_5465,N_3879,N_2201);
or U5466 (N_5466,N_2215,N_3085);
nor U5467 (N_5467,N_2333,N_2705);
and U5468 (N_5468,N_3694,N_3591);
nor U5469 (N_5469,N_2925,N_3216);
nand U5470 (N_5470,N_3000,N_3369);
and U5471 (N_5471,N_3163,N_2398);
nand U5472 (N_5472,N_3244,N_3397);
nor U5473 (N_5473,N_3268,N_2230);
nand U5474 (N_5474,N_2912,N_3572);
or U5475 (N_5475,N_2753,N_2363);
or U5476 (N_5476,N_3242,N_3089);
or U5477 (N_5477,N_3113,N_2912);
nor U5478 (N_5478,N_2998,N_2599);
or U5479 (N_5479,N_2709,N_3124);
nor U5480 (N_5480,N_3271,N_3008);
nand U5481 (N_5481,N_3438,N_3661);
nor U5482 (N_5482,N_3246,N_2040);
xor U5483 (N_5483,N_3462,N_3265);
or U5484 (N_5484,N_2327,N_3122);
nand U5485 (N_5485,N_3008,N_2655);
and U5486 (N_5486,N_3173,N_3233);
nand U5487 (N_5487,N_2230,N_2365);
or U5488 (N_5488,N_2018,N_3508);
or U5489 (N_5489,N_2605,N_2310);
and U5490 (N_5490,N_3281,N_3979);
and U5491 (N_5491,N_3024,N_3148);
nand U5492 (N_5492,N_3544,N_3243);
or U5493 (N_5493,N_3514,N_2264);
nand U5494 (N_5494,N_2992,N_3122);
xor U5495 (N_5495,N_2934,N_3910);
nand U5496 (N_5496,N_3224,N_2517);
or U5497 (N_5497,N_3570,N_2644);
nand U5498 (N_5498,N_3421,N_2868);
and U5499 (N_5499,N_3562,N_2185);
nor U5500 (N_5500,N_3403,N_2423);
nor U5501 (N_5501,N_3876,N_3779);
xor U5502 (N_5502,N_2299,N_3135);
nand U5503 (N_5503,N_2464,N_2267);
nor U5504 (N_5504,N_3024,N_3732);
or U5505 (N_5505,N_2807,N_3894);
or U5506 (N_5506,N_2447,N_2610);
and U5507 (N_5507,N_3549,N_3494);
nor U5508 (N_5508,N_3844,N_2751);
or U5509 (N_5509,N_3651,N_3336);
nor U5510 (N_5510,N_2016,N_2863);
or U5511 (N_5511,N_3790,N_2740);
and U5512 (N_5512,N_3039,N_3901);
nor U5513 (N_5513,N_2192,N_2939);
nand U5514 (N_5514,N_2369,N_3233);
nor U5515 (N_5515,N_3428,N_2032);
nand U5516 (N_5516,N_2934,N_3241);
and U5517 (N_5517,N_3252,N_2627);
xnor U5518 (N_5518,N_2481,N_3507);
nand U5519 (N_5519,N_2954,N_3752);
or U5520 (N_5520,N_3563,N_3193);
nand U5521 (N_5521,N_2324,N_3002);
or U5522 (N_5522,N_3309,N_3600);
and U5523 (N_5523,N_3923,N_3454);
nand U5524 (N_5524,N_2861,N_2424);
and U5525 (N_5525,N_2940,N_2311);
nand U5526 (N_5526,N_3045,N_2702);
nor U5527 (N_5527,N_3916,N_2390);
or U5528 (N_5528,N_3846,N_3250);
and U5529 (N_5529,N_2571,N_2972);
xor U5530 (N_5530,N_3807,N_2328);
nor U5531 (N_5531,N_2014,N_3640);
and U5532 (N_5532,N_2411,N_2532);
and U5533 (N_5533,N_2530,N_3397);
nor U5534 (N_5534,N_3321,N_2308);
xor U5535 (N_5535,N_3137,N_3963);
nor U5536 (N_5536,N_2855,N_2456);
nand U5537 (N_5537,N_3976,N_2608);
or U5538 (N_5538,N_2525,N_2745);
and U5539 (N_5539,N_3455,N_3761);
nor U5540 (N_5540,N_3513,N_3844);
and U5541 (N_5541,N_3259,N_3956);
or U5542 (N_5542,N_3976,N_3439);
and U5543 (N_5543,N_2356,N_3533);
and U5544 (N_5544,N_2902,N_2145);
nand U5545 (N_5545,N_2481,N_3618);
and U5546 (N_5546,N_3453,N_2709);
or U5547 (N_5547,N_3809,N_3072);
or U5548 (N_5548,N_2569,N_3243);
nand U5549 (N_5549,N_2957,N_3653);
or U5550 (N_5550,N_2533,N_2746);
or U5551 (N_5551,N_3060,N_3636);
nand U5552 (N_5552,N_3515,N_2313);
or U5553 (N_5553,N_3732,N_3137);
nand U5554 (N_5554,N_2888,N_2327);
nand U5555 (N_5555,N_2611,N_2369);
nand U5556 (N_5556,N_3786,N_3451);
and U5557 (N_5557,N_2614,N_2299);
nor U5558 (N_5558,N_2760,N_2486);
and U5559 (N_5559,N_2233,N_2204);
nand U5560 (N_5560,N_2941,N_2015);
nand U5561 (N_5561,N_3384,N_2743);
nor U5562 (N_5562,N_2787,N_2157);
nand U5563 (N_5563,N_2060,N_2820);
nand U5564 (N_5564,N_2650,N_3586);
nand U5565 (N_5565,N_3291,N_2280);
nor U5566 (N_5566,N_3230,N_3850);
or U5567 (N_5567,N_3784,N_2136);
xnor U5568 (N_5568,N_2020,N_3546);
and U5569 (N_5569,N_2007,N_2751);
nor U5570 (N_5570,N_3191,N_3518);
nand U5571 (N_5571,N_2342,N_2078);
nand U5572 (N_5572,N_2399,N_3497);
nand U5573 (N_5573,N_2884,N_2279);
nand U5574 (N_5574,N_2860,N_3114);
xor U5575 (N_5575,N_3434,N_3123);
nand U5576 (N_5576,N_2758,N_2117);
or U5577 (N_5577,N_2981,N_3704);
or U5578 (N_5578,N_2913,N_2180);
or U5579 (N_5579,N_2035,N_3235);
or U5580 (N_5580,N_2721,N_3358);
nand U5581 (N_5581,N_2508,N_3021);
nor U5582 (N_5582,N_3294,N_2615);
and U5583 (N_5583,N_2897,N_3544);
or U5584 (N_5584,N_2340,N_3242);
nand U5585 (N_5585,N_3195,N_2151);
and U5586 (N_5586,N_2403,N_2551);
nand U5587 (N_5587,N_2637,N_2053);
nor U5588 (N_5588,N_3483,N_2609);
or U5589 (N_5589,N_2629,N_3419);
and U5590 (N_5590,N_2810,N_2514);
or U5591 (N_5591,N_2022,N_2387);
nand U5592 (N_5592,N_2834,N_2558);
and U5593 (N_5593,N_3696,N_2609);
nand U5594 (N_5594,N_2107,N_3644);
and U5595 (N_5595,N_2779,N_2651);
and U5596 (N_5596,N_3959,N_3024);
nand U5597 (N_5597,N_3281,N_2464);
and U5598 (N_5598,N_2025,N_3471);
or U5599 (N_5599,N_3651,N_3252);
and U5600 (N_5600,N_2205,N_3992);
xor U5601 (N_5601,N_3725,N_3281);
nor U5602 (N_5602,N_3409,N_2627);
xor U5603 (N_5603,N_3890,N_2360);
and U5604 (N_5604,N_2944,N_2268);
nor U5605 (N_5605,N_3571,N_3694);
or U5606 (N_5606,N_2559,N_3928);
xor U5607 (N_5607,N_3114,N_3685);
nor U5608 (N_5608,N_2023,N_3040);
nand U5609 (N_5609,N_2109,N_2286);
nand U5610 (N_5610,N_3494,N_2394);
and U5611 (N_5611,N_3004,N_2046);
nor U5612 (N_5612,N_2857,N_3470);
nor U5613 (N_5613,N_3205,N_2769);
xor U5614 (N_5614,N_3794,N_2342);
nor U5615 (N_5615,N_3792,N_3570);
and U5616 (N_5616,N_3308,N_3444);
nand U5617 (N_5617,N_2388,N_3225);
nand U5618 (N_5618,N_2569,N_2746);
and U5619 (N_5619,N_2453,N_3329);
or U5620 (N_5620,N_3867,N_2998);
nand U5621 (N_5621,N_3169,N_2792);
and U5622 (N_5622,N_3788,N_2986);
nand U5623 (N_5623,N_3428,N_3619);
nor U5624 (N_5624,N_3238,N_3882);
nand U5625 (N_5625,N_3804,N_2729);
and U5626 (N_5626,N_2460,N_3080);
or U5627 (N_5627,N_2626,N_2983);
xor U5628 (N_5628,N_2304,N_2127);
and U5629 (N_5629,N_2077,N_3638);
and U5630 (N_5630,N_2087,N_3866);
xor U5631 (N_5631,N_2074,N_3318);
nand U5632 (N_5632,N_2783,N_3778);
and U5633 (N_5633,N_3633,N_3829);
or U5634 (N_5634,N_2543,N_2053);
and U5635 (N_5635,N_3712,N_2986);
and U5636 (N_5636,N_3227,N_2617);
and U5637 (N_5637,N_3768,N_3113);
nor U5638 (N_5638,N_2073,N_3672);
or U5639 (N_5639,N_2429,N_3526);
and U5640 (N_5640,N_3075,N_3132);
nor U5641 (N_5641,N_2682,N_3010);
nor U5642 (N_5642,N_3454,N_3567);
or U5643 (N_5643,N_3553,N_3321);
or U5644 (N_5644,N_3223,N_3780);
and U5645 (N_5645,N_2911,N_3366);
nor U5646 (N_5646,N_2627,N_2203);
xnor U5647 (N_5647,N_3250,N_3055);
nand U5648 (N_5648,N_2484,N_3486);
or U5649 (N_5649,N_3541,N_3014);
or U5650 (N_5650,N_3562,N_2320);
nor U5651 (N_5651,N_3794,N_2464);
nand U5652 (N_5652,N_3560,N_2481);
and U5653 (N_5653,N_3990,N_3391);
nand U5654 (N_5654,N_2052,N_2657);
nor U5655 (N_5655,N_3414,N_2460);
nor U5656 (N_5656,N_3647,N_3891);
and U5657 (N_5657,N_3089,N_2855);
and U5658 (N_5658,N_2004,N_2578);
nor U5659 (N_5659,N_2980,N_2261);
xnor U5660 (N_5660,N_2955,N_3825);
nor U5661 (N_5661,N_2983,N_2947);
and U5662 (N_5662,N_2103,N_2292);
nor U5663 (N_5663,N_2720,N_3194);
xor U5664 (N_5664,N_2720,N_2164);
and U5665 (N_5665,N_3238,N_2946);
or U5666 (N_5666,N_2218,N_3662);
and U5667 (N_5667,N_2279,N_3580);
nand U5668 (N_5668,N_3575,N_3173);
or U5669 (N_5669,N_3067,N_2556);
nand U5670 (N_5670,N_2920,N_2140);
nand U5671 (N_5671,N_3201,N_2770);
xor U5672 (N_5672,N_3224,N_2505);
or U5673 (N_5673,N_2578,N_3499);
nor U5674 (N_5674,N_3173,N_2527);
or U5675 (N_5675,N_2517,N_2779);
nor U5676 (N_5676,N_2056,N_3693);
nand U5677 (N_5677,N_3602,N_2870);
and U5678 (N_5678,N_3070,N_3054);
and U5679 (N_5679,N_3379,N_3006);
nand U5680 (N_5680,N_3256,N_3656);
and U5681 (N_5681,N_3997,N_2438);
nor U5682 (N_5682,N_3914,N_2371);
nor U5683 (N_5683,N_2833,N_3747);
nor U5684 (N_5684,N_3550,N_2679);
or U5685 (N_5685,N_3354,N_3982);
nand U5686 (N_5686,N_3835,N_3270);
nor U5687 (N_5687,N_3245,N_2438);
nor U5688 (N_5688,N_2033,N_2281);
or U5689 (N_5689,N_2890,N_2050);
nand U5690 (N_5690,N_2715,N_3401);
nor U5691 (N_5691,N_2085,N_2963);
nor U5692 (N_5692,N_2628,N_3504);
nand U5693 (N_5693,N_2620,N_3820);
or U5694 (N_5694,N_2082,N_3519);
nor U5695 (N_5695,N_2356,N_3102);
or U5696 (N_5696,N_2140,N_3135);
nand U5697 (N_5697,N_3525,N_2983);
nor U5698 (N_5698,N_3775,N_3211);
or U5699 (N_5699,N_2703,N_2357);
nand U5700 (N_5700,N_3717,N_3942);
xnor U5701 (N_5701,N_3950,N_2191);
or U5702 (N_5702,N_3312,N_3800);
nor U5703 (N_5703,N_3860,N_3323);
nand U5704 (N_5704,N_3179,N_3132);
nor U5705 (N_5705,N_2901,N_3153);
nand U5706 (N_5706,N_2044,N_3310);
or U5707 (N_5707,N_2617,N_2071);
or U5708 (N_5708,N_3855,N_2350);
nor U5709 (N_5709,N_2619,N_3561);
nand U5710 (N_5710,N_2540,N_2822);
or U5711 (N_5711,N_2012,N_3271);
xnor U5712 (N_5712,N_2840,N_2092);
or U5713 (N_5713,N_2098,N_2411);
and U5714 (N_5714,N_3033,N_3799);
nor U5715 (N_5715,N_3070,N_3635);
and U5716 (N_5716,N_3182,N_2487);
or U5717 (N_5717,N_2807,N_2673);
nand U5718 (N_5718,N_2605,N_2987);
or U5719 (N_5719,N_3230,N_3153);
and U5720 (N_5720,N_2705,N_2079);
nor U5721 (N_5721,N_2577,N_2183);
or U5722 (N_5722,N_2304,N_3584);
nor U5723 (N_5723,N_3651,N_3160);
xnor U5724 (N_5724,N_2932,N_3172);
or U5725 (N_5725,N_3786,N_3879);
and U5726 (N_5726,N_3625,N_3414);
nor U5727 (N_5727,N_2956,N_2097);
and U5728 (N_5728,N_2719,N_2357);
or U5729 (N_5729,N_3717,N_2247);
and U5730 (N_5730,N_3533,N_2524);
or U5731 (N_5731,N_3183,N_2687);
nand U5732 (N_5732,N_3168,N_2191);
or U5733 (N_5733,N_3440,N_2866);
nand U5734 (N_5734,N_3955,N_3029);
or U5735 (N_5735,N_3793,N_2491);
nor U5736 (N_5736,N_3327,N_3147);
or U5737 (N_5737,N_2687,N_2641);
nor U5738 (N_5738,N_2369,N_2418);
or U5739 (N_5739,N_2961,N_3969);
or U5740 (N_5740,N_3313,N_3510);
or U5741 (N_5741,N_2269,N_3653);
or U5742 (N_5742,N_2702,N_2448);
nor U5743 (N_5743,N_2831,N_2301);
or U5744 (N_5744,N_3332,N_3435);
nand U5745 (N_5745,N_3080,N_2382);
nor U5746 (N_5746,N_2311,N_2393);
and U5747 (N_5747,N_3849,N_3932);
nor U5748 (N_5748,N_3148,N_2874);
xor U5749 (N_5749,N_2882,N_2158);
or U5750 (N_5750,N_2463,N_2461);
or U5751 (N_5751,N_3056,N_3888);
nand U5752 (N_5752,N_2799,N_3187);
and U5753 (N_5753,N_2147,N_3506);
xor U5754 (N_5754,N_3438,N_3883);
or U5755 (N_5755,N_2909,N_3844);
nor U5756 (N_5756,N_2511,N_3181);
nor U5757 (N_5757,N_3980,N_2058);
and U5758 (N_5758,N_3297,N_3134);
or U5759 (N_5759,N_2559,N_3219);
and U5760 (N_5760,N_3021,N_2466);
or U5761 (N_5761,N_2003,N_2028);
nor U5762 (N_5762,N_2732,N_2596);
nor U5763 (N_5763,N_2530,N_3819);
nand U5764 (N_5764,N_2109,N_2317);
nand U5765 (N_5765,N_2993,N_3013);
or U5766 (N_5766,N_3551,N_3222);
nand U5767 (N_5767,N_3570,N_3323);
nand U5768 (N_5768,N_2248,N_3987);
nand U5769 (N_5769,N_2052,N_2118);
xnor U5770 (N_5770,N_3816,N_3630);
nor U5771 (N_5771,N_2163,N_2429);
nand U5772 (N_5772,N_3484,N_3858);
or U5773 (N_5773,N_3683,N_2302);
nand U5774 (N_5774,N_3942,N_3377);
or U5775 (N_5775,N_3465,N_3069);
nor U5776 (N_5776,N_3314,N_2750);
or U5777 (N_5777,N_2665,N_2641);
and U5778 (N_5778,N_3943,N_3040);
or U5779 (N_5779,N_2900,N_3561);
or U5780 (N_5780,N_2704,N_3520);
and U5781 (N_5781,N_3712,N_3297);
or U5782 (N_5782,N_3880,N_3622);
or U5783 (N_5783,N_2975,N_2358);
xnor U5784 (N_5784,N_2251,N_2964);
and U5785 (N_5785,N_2261,N_2629);
nand U5786 (N_5786,N_3881,N_2569);
or U5787 (N_5787,N_2202,N_3587);
and U5788 (N_5788,N_3573,N_3716);
or U5789 (N_5789,N_3838,N_2502);
nand U5790 (N_5790,N_3166,N_2806);
and U5791 (N_5791,N_3918,N_2069);
or U5792 (N_5792,N_3730,N_2163);
and U5793 (N_5793,N_3909,N_2091);
and U5794 (N_5794,N_2624,N_2027);
xnor U5795 (N_5795,N_3097,N_2393);
or U5796 (N_5796,N_3071,N_3252);
and U5797 (N_5797,N_3694,N_3356);
nand U5798 (N_5798,N_2929,N_2460);
and U5799 (N_5799,N_2169,N_2111);
and U5800 (N_5800,N_3580,N_3722);
xnor U5801 (N_5801,N_3603,N_3842);
nor U5802 (N_5802,N_2920,N_2249);
xnor U5803 (N_5803,N_3388,N_2767);
nand U5804 (N_5804,N_2106,N_2386);
nor U5805 (N_5805,N_2912,N_3016);
and U5806 (N_5806,N_2020,N_3528);
and U5807 (N_5807,N_2269,N_3402);
or U5808 (N_5808,N_2822,N_2724);
and U5809 (N_5809,N_3177,N_3105);
xnor U5810 (N_5810,N_2574,N_3302);
nor U5811 (N_5811,N_3185,N_3405);
and U5812 (N_5812,N_3590,N_2642);
or U5813 (N_5813,N_3662,N_2442);
and U5814 (N_5814,N_3938,N_3231);
xnor U5815 (N_5815,N_3516,N_2825);
xor U5816 (N_5816,N_3522,N_2488);
and U5817 (N_5817,N_3491,N_3400);
xor U5818 (N_5818,N_3920,N_3653);
and U5819 (N_5819,N_3994,N_3157);
or U5820 (N_5820,N_3562,N_3873);
or U5821 (N_5821,N_2032,N_3039);
and U5822 (N_5822,N_3339,N_3550);
nand U5823 (N_5823,N_2122,N_3768);
nand U5824 (N_5824,N_2585,N_2884);
nor U5825 (N_5825,N_2346,N_3563);
and U5826 (N_5826,N_2745,N_3716);
or U5827 (N_5827,N_2906,N_2284);
xor U5828 (N_5828,N_3526,N_2244);
nor U5829 (N_5829,N_3994,N_3663);
nand U5830 (N_5830,N_2202,N_3030);
nand U5831 (N_5831,N_2080,N_2614);
and U5832 (N_5832,N_3828,N_2588);
or U5833 (N_5833,N_2778,N_3423);
nor U5834 (N_5834,N_3469,N_2361);
and U5835 (N_5835,N_3282,N_3674);
or U5836 (N_5836,N_2329,N_3077);
nor U5837 (N_5837,N_3901,N_2328);
and U5838 (N_5838,N_3575,N_2988);
and U5839 (N_5839,N_2876,N_2488);
and U5840 (N_5840,N_3353,N_2790);
nor U5841 (N_5841,N_2183,N_2252);
or U5842 (N_5842,N_3694,N_3220);
or U5843 (N_5843,N_3425,N_2586);
xor U5844 (N_5844,N_3722,N_2458);
and U5845 (N_5845,N_2922,N_2344);
nor U5846 (N_5846,N_3539,N_2836);
or U5847 (N_5847,N_2840,N_3007);
nor U5848 (N_5848,N_2448,N_2826);
and U5849 (N_5849,N_3739,N_2606);
nand U5850 (N_5850,N_3243,N_3407);
or U5851 (N_5851,N_3455,N_3954);
and U5852 (N_5852,N_3534,N_3299);
nor U5853 (N_5853,N_2180,N_2087);
or U5854 (N_5854,N_3748,N_3309);
nor U5855 (N_5855,N_3974,N_2147);
and U5856 (N_5856,N_3251,N_3117);
nor U5857 (N_5857,N_2638,N_3408);
xnor U5858 (N_5858,N_2526,N_3052);
nand U5859 (N_5859,N_3860,N_2246);
nor U5860 (N_5860,N_2994,N_3524);
or U5861 (N_5861,N_3403,N_3619);
and U5862 (N_5862,N_3136,N_3387);
and U5863 (N_5863,N_2890,N_3901);
nor U5864 (N_5864,N_2643,N_3261);
nor U5865 (N_5865,N_3008,N_2898);
xor U5866 (N_5866,N_3536,N_3335);
and U5867 (N_5867,N_3414,N_3917);
nor U5868 (N_5868,N_2178,N_3094);
nand U5869 (N_5869,N_2323,N_2373);
or U5870 (N_5870,N_3622,N_2403);
and U5871 (N_5871,N_2556,N_3398);
xor U5872 (N_5872,N_2217,N_2145);
nand U5873 (N_5873,N_2572,N_2447);
nor U5874 (N_5874,N_2920,N_2850);
or U5875 (N_5875,N_2227,N_2930);
or U5876 (N_5876,N_3658,N_3955);
nand U5877 (N_5877,N_3451,N_3106);
nor U5878 (N_5878,N_2823,N_3708);
and U5879 (N_5879,N_3881,N_3629);
nor U5880 (N_5880,N_2194,N_3352);
or U5881 (N_5881,N_3113,N_3561);
nand U5882 (N_5882,N_3345,N_2389);
xor U5883 (N_5883,N_3312,N_3215);
nand U5884 (N_5884,N_2513,N_2623);
or U5885 (N_5885,N_2855,N_3823);
nor U5886 (N_5886,N_2044,N_3889);
or U5887 (N_5887,N_2317,N_2629);
nand U5888 (N_5888,N_2690,N_2137);
nand U5889 (N_5889,N_3350,N_3209);
nand U5890 (N_5890,N_2473,N_3297);
and U5891 (N_5891,N_3065,N_3071);
or U5892 (N_5892,N_3643,N_3019);
or U5893 (N_5893,N_2467,N_2450);
nand U5894 (N_5894,N_3169,N_2561);
or U5895 (N_5895,N_3515,N_2041);
or U5896 (N_5896,N_2518,N_3002);
nand U5897 (N_5897,N_2772,N_3674);
nand U5898 (N_5898,N_3157,N_2383);
and U5899 (N_5899,N_2455,N_3653);
and U5900 (N_5900,N_3257,N_3688);
nor U5901 (N_5901,N_3042,N_3466);
xor U5902 (N_5902,N_3762,N_2328);
and U5903 (N_5903,N_2904,N_3939);
and U5904 (N_5904,N_3961,N_2635);
or U5905 (N_5905,N_2712,N_2455);
and U5906 (N_5906,N_2239,N_2751);
nor U5907 (N_5907,N_3756,N_3118);
or U5908 (N_5908,N_2135,N_3035);
and U5909 (N_5909,N_3152,N_3779);
and U5910 (N_5910,N_3164,N_2456);
or U5911 (N_5911,N_3101,N_2998);
or U5912 (N_5912,N_2308,N_3479);
or U5913 (N_5913,N_2703,N_3777);
and U5914 (N_5914,N_2921,N_2887);
nor U5915 (N_5915,N_3796,N_2909);
nand U5916 (N_5916,N_3307,N_2784);
nor U5917 (N_5917,N_2127,N_2502);
nor U5918 (N_5918,N_3142,N_2401);
xnor U5919 (N_5919,N_3928,N_3108);
nand U5920 (N_5920,N_2357,N_3440);
nand U5921 (N_5921,N_3050,N_2071);
and U5922 (N_5922,N_2624,N_2858);
xor U5923 (N_5923,N_2593,N_3390);
and U5924 (N_5924,N_2401,N_3007);
nor U5925 (N_5925,N_3433,N_3455);
nor U5926 (N_5926,N_2016,N_2681);
and U5927 (N_5927,N_2887,N_2334);
nor U5928 (N_5928,N_2303,N_2092);
and U5929 (N_5929,N_2730,N_3145);
or U5930 (N_5930,N_2752,N_2989);
nor U5931 (N_5931,N_3955,N_2399);
and U5932 (N_5932,N_3103,N_3330);
and U5933 (N_5933,N_3849,N_3642);
xor U5934 (N_5934,N_3968,N_2039);
or U5935 (N_5935,N_2321,N_2294);
and U5936 (N_5936,N_2248,N_3729);
and U5937 (N_5937,N_2841,N_3986);
nor U5938 (N_5938,N_3589,N_3187);
nor U5939 (N_5939,N_2936,N_2817);
nand U5940 (N_5940,N_2201,N_3115);
xnor U5941 (N_5941,N_3863,N_2000);
or U5942 (N_5942,N_2656,N_2879);
and U5943 (N_5943,N_2152,N_3779);
nand U5944 (N_5944,N_2343,N_2992);
xnor U5945 (N_5945,N_2022,N_2983);
nor U5946 (N_5946,N_2968,N_2538);
and U5947 (N_5947,N_2656,N_2646);
and U5948 (N_5948,N_3752,N_2415);
or U5949 (N_5949,N_3958,N_3431);
or U5950 (N_5950,N_3788,N_3482);
nand U5951 (N_5951,N_2746,N_2875);
and U5952 (N_5952,N_3319,N_3270);
and U5953 (N_5953,N_3228,N_3291);
nand U5954 (N_5954,N_2029,N_2237);
and U5955 (N_5955,N_2859,N_2435);
xnor U5956 (N_5956,N_3418,N_2150);
nand U5957 (N_5957,N_3217,N_3253);
nand U5958 (N_5958,N_3063,N_3696);
or U5959 (N_5959,N_3923,N_2808);
nor U5960 (N_5960,N_2598,N_2582);
xnor U5961 (N_5961,N_2580,N_2346);
nor U5962 (N_5962,N_2125,N_3286);
xor U5963 (N_5963,N_3233,N_3498);
or U5964 (N_5964,N_2593,N_3612);
xnor U5965 (N_5965,N_3037,N_3584);
nor U5966 (N_5966,N_2840,N_2760);
nand U5967 (N_5967,N_2976,N_3144);
nand U5968 (N_5968,N_3524,N_2165);
nand U5969 (N_5969,N_3669,N_3322);
or U5970 (N_5970,N_3155,N_3344);
nor U5971 (N_5971,N_2517,N_2579);
nand U5972 (N_5972,N_2890,N_3189);
nand U5973 (N_5973,N_2206,N_2540);
nor U5974 (N_5974,N_2320,N_3153);
xor U5975 (N_5975,N_3170,N_3448);
and U5976 (N_5976,N_3459,N_2375);
nor U5977 (N_5977,N_3078,N_2613);
xor U5978 (N_5978,N_2721,N_3184);
or U5979 (N_5979,N_3106,N_2988);
and U5980 (N_5980,N_3537,N_2591);
and U5981 (N_5981,N_2695,N_3266);
and U5982 (N_5982,N_3177,N_3590);
nand U5983 (N_5983,N_3928,N_3876);
xor U5984 (N_5984,N_2890,N_2515);
xor U5985 (N_5985,N_3278,N_2961);
or U5986 (N_5986,N_3299,N_3201);
or U5987 (N_5987,N_3470,N_2166);
or U5988 (N_5988,N_3981,N_2381);
nand U5989 (N_5989,N_3359,N_3154);
and U5990 (N_5990,N_2294,N_2789);
nand U5991 (N_5991,N_2365,N_3281);
or U5992 (N_5992,N_2690,N_2919);
and U5993 (N_5993,N_2123,N_2314);
xnor U5994 (N_5994,N_2254,N_3021);
and U5995 (N_5995,N_2195,N_3438);
and U5996 (N_5996,N_3082,N_3652);
and U5997 (N_5997,N_3391,N_3239);
xor U5998 (N_5998,N_3746,N_2696);
nand U5999 (N_5999,N_3192,N_3256);
or U6000 (N_6000,N_4374,N_5062);
nor U6001 (N_6001,N_4870,N_5203);
nor U6002 (N_6002,N_4724,N_4209);
or U6003 (N_6003,N_4442,N_4107);
nand U6004 (N_6004,N_4383,N_5059);
xnor U6005 (N_6005,N_4886,N_4037);
or U6006 (N_6006,N_5131,N_5933);
nand U6007 (N_6007,N_4660,N_5308);
nor U6008 (N_6008,N_4179,N_5068);
and U6009 (N_6009,N_4709,N_5500);
and U6010 (N_6010,N_4305,N_5527);
nand U6011 (N_6011,N_5016,N_5956);
xnor U6012 (N_6012,N_4652,N_4701);
or U6013 (N_6013,N_5344,N_5830);
nand U6014 (N_6014,N_4087,N_5389);
nand U6015 (N_6015,N_4632,N_4919);
or U6016 (N_6016,N_5113,N_5775);
or U6017 (N_6017,N_5081,N_5580);
nand U6018 (N_6018,N_4387,N_4655);
nor U6019 (N_6019,N_5869,N_4214);
or U6020 (N_6020,N_5816,N_5084);
xnor U6021 (N_6021,N_4345,N_5958);
and U6022 (N_6022,N_5616,N_5337);
nor U6023 (N_6023,N_4921,N_5388);
nand U6024 (N_6024,N_5174,N_5661);
nand U6025 (N_6025,N_5623,N_5665);
and U6026 (N_6026,N_4169,N_4472);
xor U6027 (N_6027,N_4860,N_5892);
and U6028 (N_6028,N_4876,N_4764);
and U6029 (N_6029,N_4751,N_5585);
nor U6030 (N_6030,N_4850,N_4032);
and U6031 (N_6031,N_5292,N_5626);
nand U6032 (N_6032,N_4769,N_5791);
nor U6033 (N_6033,N_5289,N_4497);
nand U6034 (N_6034,N_4903,N_4076);
xor U6035 (N_6035,N_5175,N_4829);
and U6036 (N_6036,N_4936,N_4338);
xnor U6037 (N_6037,N_5662,N_5144);
nand U6038 (N_6038,N_4201,N_4493);
and U6039 (N_6039,N_4448,N_4384);
or U6040 (N_6040,N_4450,N_4489);
nand U6041 (N_6041,N_4646,N_5087);
xor U6042 (N_6042,N_4217,N_5544);
or U6043 (N_6043,N_5558,N_5298);
nor U6044 (N_6044,N_4954,N_5032);
or U6045 (N_6045,N_4017,N_5919);
nand U6046 (N_6046,N_4015,N_4466);
and U6047 (N_6047,N_5941,N_5805);
nand U6048 (N_6048,N_5075,N_4164);
or U6049 (N_6049,N_5461,N_5227);
and U6050 (N_6050,N_4985,N_5392);
or U6051 (N_6051,N_5347,N_5149);
nand U6052 (N_6052,N_5080,N_4246);
xnor U6053 (N_6053,N_4665,N_4986);
and U6054 (N_6054,N_4331,N_5902);
nor U6055 (N_6055,N_5312,N_4651);
or U6056 (N_6056,N_5686,N_5405);
or U6057 (N_6057,N_4184,N_5287);
and U6058 (N_6058,N_5300,N_5163);
nand U6059 (N_6059,N_5364,N_4694);
and U6060 (N_6060,N_5606,N_5055);
and U6061 (N_6061,N_5443,N_4056);
nor U6062 (N_6062,N_4511,N_5969);
and U6063 (N_6063,N_4456,N_5126);
nor U6064 (N_6064,N_4647,N_4344);
nand U6065 (N_6065,N_4341,N_4046);
nand U6066 (N_6066,N_4216,N_4455);
nand U6067 (N_6067,N_4020,N_5598);
nand U6068 (N_6068,N_4594,N_5517);
and U6069 (N_6069,N_5641,N_5384);
and U6070 (N_6070,N_5744,N_4621);
nor U6071 (N_6071,N_4888,N_4162);
nor U6072 (N_6072,N_4356,N_5226);
and U6073 (N_6073,N_4950,N_4306);
and U6074 (N_6074,N_4353,N_5758);
nor U6075 (N_6075,N_5514,N_5005);
or U6076 (N_6076,N_5765,N_4396);
and U6077 (N_6077,N_5767,N_4541);
nor U6078 (N_6078,N_4153,N_4818);
or U6079 (N_6079,N_4640,N_5900);
nand U6080 (N_6080,N_5469,N_5881);
nor U6081 (N_6081,N_5414,N_4127);
nand U6082 (N_6082,N_4505,N_4639);
nand U6083 (N_6083,N_4370,N_4617);
or U6084 (N_6084,N_4776,N_4206);
nor U6085 (N_6085,N_4653,N_4117);
nand U6086 (N_6086,N_5865,N_5582);
nor U6087 (N_6087,N_4375,N_4278);
nand U6088 (N_6088,N_4218,N_5151);
xor U6089 (N_6089,N_5463,N_5245);
nand U6090 (N_6090,N_5733,N_5498);
or U6091 (N_6091,N_5138,N_4160);
and U6092 (N_6092,N_5346,N_4742);
or U6093 (N_6093,N_4309,N_5188);
nand U6094 (N_6094,N_4567,N_5966);
nand U6095 (N_6095,N_4600,N_5798);
nor U6096 (N_6096,N_5828,N_4314);
and U6097 (N_6097,N_4129,N_5330);
nand U6098 (N_6098,N_4780,N_5381);
and U6099 (N_6099,N_5189,N_4757);
or U6100 (N_6100,N_4154,N_5482);
or U6101 (N_6101,N_5655,N_5815);
nor U6102 (N_6102,N_5540,N_5372);
and U6103 (N_6103,N_4428,N_4915);
nand U6104 (N_6104,N_4502,N_5343);
or U6105 (N_6105,N_5313,N_5439);
nor U6106 (N_6106,N_5412,N_5070);
or U6107 (N_6107,N_5953,N_5596);
nand U6108 (N_6108,N_5315,N_4168);
nand U6109 (N_6109,N_4879,N_5594);
or U6110 (N_6110,N_4945,N_4235);
nand U6111 (N_6111,N_4244,N_5168);
nor U6112 (N_6112,N_4676,N_4680);
nand U6113 (N_6113,N_5581,N_4415);
or U6114 (N_6114,N_5358,N_4528);
or U6115 (N_6115,N_4102,N_5323);
or U6116 (N_6116,N_5882,N_4992);
nand U6117 (N_6117,N_4627,N_5123);
nor U6118 (N_6118,N_5438,N_5625);
or U6119 (N_6119,N_5546,N_5629);
or U6120 (N_6120,N_4398,N_5434);
nand U6121 (N_6121,N_5509,N_4385);
or U6122 (N_6122,N_4349,N_5150);
xnor U6123 (N_6123,N_5911,N_4846);
or U6124 (N_6124,N_5316,N_5489);
nand U6125 (N_6125,N_4299,N_5823);
nor U6126 (N_6126,N_4318,N_5913);
or U6127 (N_6127,N_5521,N_5810);
and U6128 (N_6128,N_5771,N_4181);
or U6129 (N_6129,N_4569,N_4796);
nor U6130 (N_6130,N_5001,N_4746);
or U6131 (N_6131,N_4626,N_4990);
and U6132 (N_6132,N_4295,N_4427);
nand U6133 (N_6133,N_4099,N_4662);
and U6134 (N_6134,N_5859,N_4265);
or U6135 (N_6135,N_5109,N_4925);
nor U6136 (N_6136,N_5355,N_5491);
xor U6137 (N_6137,N_5211,N_4559);
and U6138 (N_6138,N_4775,N_5942);
and U6139 (N_6139,N_5267,N_4351);
xor U6140 (N_6140,N_5750,N_4917);
or U6141 (N_6141,N_4530,N_4269);
or U6142 (N_6142,N_4435,N_4047);
nor U6143 (N_6143,N_4978,N_4783);
or U6144 (N_6144,N_4376,N_5831);
and U6145 (N_6145,N_4982,N_4008);
nor U6146 (N_6146,N_5992,N_4042);
nand U6147 (N_6147,N_4884,N_4750);
nand U6148 (N_6148,N_5009,N_4784);
xor U6149 (N_6149,N_4327,N_5761);
nand U6150 (N_6150,N_5687,N_5855);
nor U6151 (N_6151,N_5951,N_4744);
nor U6152 (N_6152,N_4935,N_5264);
xnor U6153 (N_6153,N_4538,N_5208);
or U6154 (N_6154,N_5564,N_5889);
xor U6155 (N_6155,N_5684,N_5967);
nor U6156 (N_6156,N_4156,N_4262);
xor U6157 (N_6157,N_4524,N_5303);
xor U6158 (N_6158,N_4219,N_4058);
nand U6159 (N_6159,N_5496,N_5664);
xnor U6160 (N_6160,N_4404,N_5813);
nor U6161 (N_6161,N_5410,N_5090);
or U6162 (N_6162,N_4968,N_5590);
and U6163 (N_6163,N_4735,N_4979);
nand U6164 (N_6164,N_4819,N_5004);
or U6165 (N_6165,N_5734,N_5879);
and U6166 (N_6166,N_5430,N_4223);
and U6167 (N_6167,N_5793,N_5507);
or U6168 (N_6168,N_5170,N_4059);
nor U6169 (N_6169,N_4555,N_4239);
or U6170 (N_6170,N_5922,N_5934);
or U6171 (N_6171,N_4820,N_5944);
nor U6172 (N_6172,N_5281,N_5587);
nor U6173 (N_6173,N_4506,N_5490);
or U6174 (N_6174,N_5112,N_4259);
or U6175 (N_6175,N_5978,N_5715);
nand U6176 (N_6176,N_5024,N_4362);
or U6177 (N_6177,N_5656,N_5547);
and U6178 (N_6178,N_4522,N_5536);
nand U6179 (N_6179,N_5039,N_4045);
xnor U6180 (N_6180,N_5860,N_4866);
nand U6181 (N_6181,N_4105,N_5111);
nand U6182 (N_6182,N_4586,N_5499);
nor U6183 (N_6183,N_5719,N_5773);
nor U6184 (N_6184,N_4789,N_5994);
and U6185 (N_6185,N_4564,N_4578);
nand U6186 (N_6186,N_4250,N_4468);
nand U6187 (N_6187,N_5965,N_4571);
nor U6188 (N_6188,N_4459,N_5578);
or U6189 (N_6189,N_4496,N_5017);
nor U6190 (N_6190,N_4650,N_4335);
nand U6191 (N_6191,N_4546,N_4411);
nor U6192 (N_6192,N_5400,N_5029);
nand U6193 (N_6193,N_5753,N_5272);
and U6194 (N_6194,N_5874,N_4738);
xnor U6195 (N_6195,N_4996,N_4109);
nand U6196 (N_6196,N_4922,N_5571);
and U6197 (N_6197,N_4342,N_5459);
and U6198 (N_6198,N_4893,N_5276);
and U6199 (N_6199,N_5095,N_5974);
or U6200 (N_6200,N_5931,N_4928);
and U6201 (N_6201,N_4963,N_5905);
nand U6202 (N_6202,N_5666,N_5345);
and U6203 (N_6203,N_5576,N_5610);
nor U6204 (N_6204,N_5319,N_4429);
nand U6205 (N_6205,N_5584,N_5853);
and U6206 (N_6206,N_4804,N_4336);
nor U6207 (N_6207,N_4609,N_4983);
nor U6208 (N_6208,N_4439,N_4720);
nor U6209 (N_6209,N_4878,N_4060);
xnor U6210 (N_6210,N_4022,N_5444);
nand U6211 (N_6211,N_5512,N_5885);
nand U6212 (N_6212,N_5339,N_4715);
and U6213 (N_6213,N_5106,N_4762);
and U6214 (N_6214,N_5652,N_5801);
or U6215 (N_6215,N_5746,N_5197);
and U6216 (N_6216,N_4659,N_5783);
or U6217 (N_6217,N_4055,N_4158);
and U6218 (N_6218,N_4712,N_5713);
or U6219 (N_6219,N_4579,N_5926);
or U6220 (N_6220,N_5711,N_4068);
and U6221 (N_6221,N_4361,N_4293);
nand U6222 (N_6222,N_5495,N_5539);
xor U6223 (N_6223,N_5895,N_5548);
nand U6224 (N_6224,N_4791,N_4705);
xor U6225 (N_6225,N_4943,N_4869);
and U6226 (N_6226,N_5550,N_5171);
nor U6227 (N_6227,N_5789,N_4551);
nor U6228 (N_6228,N_5341,N_5018);
or U6229 (N_6229,N_4215,N_5845);
or U6230 (N_6230,N_4822,N_5781);
and U6231 (N_6231,N_5252,N_4136);
and U6232 (N_6232,N_5561,N_5542);
and U6233 (N_6233,N_5759,N_4806);
or U6234 (N_6234,N_4658,N_4575);
or U6235 (N_6235,N_4389,N_4951);
nor U6236 (N_6236,N_4748,N_5140);
and U6237 (N_6237,N_5301,N_4561);
nor U6238 (N_6238,N_4061,N_4189);
or U6239 (N_6239,N_4645,N_5973);
nor U6240 (N_6240,N_4354,N_5110);
nor U6241 (N_6241,N_4298,N_5269);
or U6242 (N_6242,N_5128,N_5788);
nand U6243 (N_6243,N_5332,N_4501);
or U6244 (N_6244,N_4779,N_4119);
and U6245 (N_6245,N_4519,N_4731);
or U6246 (N_6246,N_5832,N_4337);
nor U6247 (N_6247,N_4044,N_5010);
and U6248 (N_6248,N_5136,N_5808);
or U6249 (N_6249,N_4290,N_5534);
nor U6250 (N_6250,N_4422,N_4212);
xor U6251 (N_6251,N_5821,N_5462);
xnor U6252 (N_6252,N_5254,N_5046);
and U6253 (N_6253,N_4350,N_5983);
nand U6254 (N_6254,N_4574,N_5875);
xnor U6255 (N_6255,N_4605,N_5383);
and U6256 (N_6256,N_4596,N_5446);
xnor U6257 (N_6257,N_5688,N_4155);
or U6258 (N_6258,N_4872,N_5173);
nand U6259 (N_6259,N_5555,N_4462);
nand U6260 (N_6260,N_5883,N_5708);
nor U6261 (N_6261,N_5777,N_4625);
nand U6262 (N_6262,N_5998,N_5045);
or U6263 (N_6263,N_5376,N_4090);
or U6264 (N_6264,N_5811,N_4326);
and U6265 (N_6265,N_4838,N_4348);
xor U6266 (N_6266,N_5007,N_4749);
xor U6267 (N_6267,N_5698,N_4874);
nand U6268 (N_6268,N_5871,N_4842);
nand U6269 (N_6269,N_5653,N_4438);
nand U6270 (N_6270,N_5703,N_5732);
xnor U6271 (N_6271,N_5088,N_4832);
and U6272 (N_6272,N_4294,N_5259);
xnor U6273 (N_6273,N_5402,N_5326);
or U6274 (N_6274,N_4861,N_5729);
or U6275 (N_6275,N_4133,N_5256);
nor U6276 (N_6276,N_4033,N_4110);
nor U6277 (N_6277,N_5363,N_4255);
and U6278 (N_6278,N_5371,N_4558);
nor U6279 (N_6279,N_5200,N_4853);
nand U6280 (N_6280,N_4150,N_5725);
nand U6281 (N_6281,N_4964,N_4001);
and U6282 (N_6282,N_4857,N_4587);
nor U6283 (N_6283,N_4920,N_4657);
or U6284 (N_6284,N_4260,N_4949);
nand U6285 (N_6285,N_4918,N_5949);
nor U6286 (N_6286,N_4699,N_4393);
nand U6287 (N_6287,N_5503,N_5041);
xnor U6288 (N_6288,N_5774,N_5425);
nand U6289 (N_6289,N_5685,N_5336);
or U6290 (N_6290,N_4364,N_5995);
or U6291 (N_6291,N_5689,N_5280);
nor U6292 (N_6292,N_4108,N_5844);
nand U6293 (N_6293,N_4664,N_5675);
nand U6294 (N_6294,N_5955,N_5757);
nor U6295 (N_6295,N_4431,N_5036);
nor U6296 (N_6296,N_4817,N_5671);
and U6297 (N_6297,N_5877,N_5320);
xnor U6298 (N_6298,N_4931,N_4821);
nand U6299 (N_6299,N_5103,N_4077);
nor U6300 (N_6300,N_4210,N_4135);
nand U6301 (N_6301,N_5465,N_5159);
and U6302 (N_6302,N_5178,N_4721);
or U6303 (N_6303,N_4611,N_4080);
xnor U6304 (N_6304,N_5214,N_5947);
or U6305 (N_6305,N_4892,N_5614);
nand U6306 (N_6306,N_5888,N_4906);
nor U6307 (N_6307,N_4405,N_4768);
nand U6308 (N_6308,N_5043,N_4115);
and U6309 (N_6309,N_4446,N_5360);
nand U6310 (N_6310,N_4165,N_4612);
and U6311 (N_6311,N_4677,N_4603);
nor U6312 (N_6312,N_5658,N_5195);
nor U6313 (N_6313,N_5085,N_5984);
or U6314 (N_6314,N_4036,N_4159);
or U6315 (N_6315,N_4799,N_4897);
or U6316 (N_6316,N_4321,N_5218);
xor U6317 (N_6317,N_5607,N_4713);
or U6318 (N_6318,N_5285,N_5102);
or U6319 (N_6319,N_5243,N_5894);
and U6320 (N_6320,N_5787,N_4691);
nor U6321 (N_6321,N_4220,N_5593);
nand U6322 (N_6322,N_5960,N_4395);
nand U6323 (N_6323,N_5468,N_5190);
and U6324 (N_6324,N_5851,N_5739);
nand U6325 (N_6325,N_4910,N_4794);
xnor U6326 (N_6326,N_5533,N_4436);
or U6327 (N_6327,N_4116,N_4152);
or U6328 (N_6328,N_5878,N_4771);
or U6329 (N_6329,N_4163,N_4425);
or U6330 (N_6330,N_5193,N_4868);
xnor U6331 (N_6331,N_5583,N_4955);
or U6332 (N_6332,N_5930,N_4499);
or U6333 (N_6333,N_5957,N_4078);
nand U6334 (N_6334,N_4171,N_5297);
or U6335 (N_6335,N_4743,N_5089);
nor U6336 (N_6336,N_4301,N_5311);
nand U6337 (N_6337,N_5730,N_5637);
nand U6338 (N_6338,N_5999,N_5532);
xnor U6339 (N_6339,N_4407,N_4543);
nand U6340 (N_6340,N_4018,N_5480);
or U6341 (N_6341,N_5519,N_4987);
nor U6342 (N_6342,N_5240,N_4254);
nand U6343 (N_6343,N_5266,N_4707);
nand U6344 (N_6344,N_4604,N_5597);
and U6345 (N_6345,N_5943,N_4126);
and U6346 (N_6346,N_5903,N_5620);
and U6347 (N_6347,N_4830,N_5403);
nand U6348 (N_6348,N_5391,N_5792);
and U6349 (N_6349,N_5745,N_4606);
nor U6350 (N_6350,N_5058,N_5162);
nor U6351 (N_6351,N_5954,N_4545);
nand U6352 (N_6352,N_4668,N_5317);
nor U6353 (N_6353,N_4096,N_4841);
nor U6354 (N_6354,N_4890,N_4898);
and U6355 (N_6355,N_4084,N_4113);
nand U6356 (N_6356,N_5229,N_4914);
nor U6357 (N_6357,N_5839,N_4614);
and U6358 (N_6358,N_4086,N_4121);
nand U6359 (N_6359,N_4871,N_4565);
nor U6360 (N_6360,N_4192,N_5868);
nand U6361 (N_6361,N_5492,N_4800);
nand U6362 (N_6362,N_5249,N_5856);
nor U6363 (N_6363,N_4844,N_4761);
and U6364 (N_6364,N_5707,N_5470);
or U6365 (N_6365,N_4098,N_5359);
nand U6366 (N_6366,N_5647,N_4333);
nor U6367 (N_6367,N_5985,N_4388);
nand U6368 (N_6368,N_5169,N_5820);
nand U6369 (N_6369,N_4494,N_5660);
nor U6370 (N_6370,N_5522,N_4324);
or U6371 (N_6371,N_5442,N_4225);
or U6372 (N_6372,N_5120,N_4131);
or U6373 (N_6373,N_4368,N_5023);
or U6374 (N_6374,N_4390,N_4287);
nand U6375 (N_6375,N_4881,N_4016);
xnor U6376 (N_6376,N_5104,N_4994);
xor U6377 (N_6377,N_5834,N_5731);
or U6378 (N_6378,N_5880,N_5748);
or U6379 (N_6379,N_4912,N_5204);
nand U6380 (N_6380,N_5630,N_5592);
nand U6381 (N_6381,N_5369,N_5520);
or U6382 (N_6382,N_4070,N_4803);
and U6383 (N_6383,N_4933,N_5031);
and U6384 (N_6384,N_5740,N_5460);
nor U6385 (N_6385,N_4526,N_4548);
nand U6386 (N_6386,N_5599,N_5932);
xor U6387 (N_6387,N_5663,N_5724);
or U6388 (N_6388,N_5349,N_4447);
or U6389 (N_6389,N_5318,N_5567);
xnor U6390 (N_6390,N_5270,N_4946);
and U6391 (N_6391,N_5194,N_5619);
nand U6392 (N_6392,N_5866,N_4491);
and U6393 (N_6393,N_5181,N_5968);
nor U6394 (N_6394,N_5145,N_5340);
or U6395 (N_6395,N_5065,N_5776);
and U6396 (N_6396,N_4051,N_5399);
nor U6397 (N_6397,N_5130,N_4174);
or U6398 (N_6398,N_4316,N_5146);
nand U6399 (N_6399,N_5742,N_4741);
nand U6400 (N_6400,N_4141,N_5154);
or U6401 (N_6401,N_4583,N_4905);
and U6402 (N_6402,N_5408,N_4669);
xnor U6403 (N_6403,N_4476,N_4563);
and U6404 (N_6404,N_5657,N_5044);
nand U6405 (N_6405,N_4467,N_5228);
nor U6406 (N_6406,N_4095,N_4615);
or U6407 (N_6407,N_4049,N_5231);
nand U6408 (N_6408,N_5180,N_4802);
or U6409 (N_6409,N_4207,N_4588);
xor U6410 (N_6410,N_4960,N_4371);
nand U6411 (N_6411,N_4205,N_4862);
and U6412 (N_6412,N_4975,N_5993);
or U6413 (N_6413,N_4268,N_5971);
nor U6414 (N_6414,N_5121,N_4608);
nand U6415 (N_6415,N_5604,N_5557);
nor U6416 (N_6416,N_4457,N_5196);
nand U6417 (N_6417,N_4231,N_5097);
and U6418 (N_6418,N_4852,N_5807);
nor U6419 (N_6419,N_5342,N_5806);
nand U6420 (N_6420,N_4539,N_5986);
nor U6421 (N_6421,N_4745,N_5176);
xor U6422 (N_6422,N_4509,N_4727);
and U6423 (N_6423,N_5100,N_5083);
and U6424 (N_6424,N_5271,N_4849);
and U6425 (N_6425,N_5213,N_4401);
nand U6426 (N_6426,N_4175,N_4620);
and U6427 (N_6427,N_5837,N_5948);
nor U6428 (N_6428,N_4013,N_4908);
nor U6429 (N_6429,N_5472,N_4598);
or U6430 (N_6430,N_4233,N_4417);
and U6431 (N_6431,N_5279,N_4923);
and U6432 (N_6432,N_5901,N_4666);
nand U6433 (N_6433,N_5378,N_4400);
xor U6434 (N_6434,N_4540,N_5910);
and U6435 (N_6435,N_5324,N_4125);
and U6436 (N_6436,N_4635,N_5691);
or U6437 (N_6437,N_4372,N_5861);
and U6438 (N_6438,N_5038,N_5764);
nand U6439 (N_6439,N_5432,N_5278);
xnor U6440 (N_6440,N_5386,N_4196);
and U6441 (N_6441,N_5668,N_4568);
xnor U6442 (N_6442,N_5464,N_4011);
xor U6443 (N_6443,N_5404,N_4267);
nor U6444 (N_6444,N_5235,N_5397);
and U6445 (N_6445,N_4104,N_5207);
and U6446 (N_6446,N_4824,N_4942);
xnor U6447 (N_6447,N_5466,N_4339);
nand U6448 (N_6448,N_4753,N_4232);
nand U6449 (N_6449,N_4408,N_5981);
and U6450 (N_6450,N_4440,N_5752);
or U6451 (N_6451,N_4029,N_4708);
and U6452 (N_6452,N_4026,N_4249);
and U6453 (N_6453,N_4130,N_5253);
nand U6454 (N_6454,N_4280,N_4443);
and U6455 (N_6455,N_5201,N_4788);
or U6456 (N_6456,N_4697,N_5737);
xnor U6457 (N_6457,N_5447,N_5416);
or U6458 (N_6458,N_5842,N_5401);
nand U6459 (N_6459,N_5513,N_4346);
nand U6460 (N_6460,N_5886,N_4610);
nor U6461 (N_6461,N_5426,N_5219);
nor U6462 (N_6462,N_4198,N_4685);
nand U6463 (N_6463,N_5674,N_4939);
or U6464 (N_6464,N_5223,N_5129);
nand U6465 (N_6465,N_5543,N_5644);
xor U6466 (N_6466,N_5537,N_4279);
nand U6467 (N_6467,N_5659,N_5232);
or U6468 (N_6468,N_4030,N_4334);
or U6469 (N_6469,N_4437,N_4471);
and U6470 (N_6470,N_4758,N_4865);
and U6471 (N_6471,N_5293,N_4837);
and U6472 (N_6472,N_4634,N_4369);
nand U6473 (N_6473,N_5680,N_5273);
and U6474 (N_6474,N_5348,N_5912);
and U6475 (N_6475,N_5870,N_5751);
or U6476 (N_6476,N_5803,N_4798);
nor U6477 (N_6477,N_4693,N_4756);
and U6478 (N_6478,N_5133,N_4577);
and U6479 (N_6479,N_4166,N_5328);
nor U6480 (N_6480,N_4997,N_5566);
and U6481 (N_6481,N_5251,N_5802);
xor U6482 (N_6482,N_4483,N_4969);
nand U6483 (N_6483,N_4864,N_4100);
nand U6484 (N_6484,N_4601,N_4128);
and U6485 (N_6485,N_4970,N_5064);
nand U6486 (N_6486,N_5950,N_4702);
or U6487 (N_6487,N_4325,N_4092);
nand U6488 (N_6488,N_5078,N_4106);
nor U6489 (N_6489,N_4271,N_4913);
and U6490 (N_6490,N_4726,N_4934);
nand U6491 (N_6491,N_4048,N_5457);
xor U6492 (N_6492,N_4759,N_5260);
nor U6493 (N_6493,N_4813,N_5202);
nor U6494 (N_6494,N_4760,N_4147);
nand U6495 (N_6495,N_4474,N_4887);
nand U6496 (N_6496,N_5728,N_5574);
or U6497 (N_6497,N_5862,N_4974);
nand U6498 (N_6498,N_4320,N_4747);
xnor U6499 (N_6499,N_4202,N_5858);
xor U6500 (N_6500,N_5327,N_4534);
and U6501 (N_6501,N_4302,N_4009);
or U6502 (N_6502,N_5473,N_4904);
and U6503 (N_6503,N_5538,N_5186);
nand U6504 (N_6504,N_4580,N_5257);
nor U6505 (N_6505,N_4479,N_4272);
nand U6506 (N_6506,N_5370,N_4962);
and U6507 (N_6507,N_4553,N_5559);
nand U6508 (N_6508,N_5924,N_5357);
nor U6509 (N_6509,N_5014,N_5628);
nand U6510 (N_6510,N_4291,N_5884);
and U6511 (N_6511,N_4071,N_5433);
nand U6512 (N_6512,N_4619,N_4357);
and U6513 (N_6513,N_5780,N_5701);
or U6514 (N_6514,N_4091,N_4692);
nor U6515 (N_6515,N_5822,N_5310);
nand U6516 (N_6516,N_4911,N_4552);
nor U6517 (N_6517,N_5716,N_4112);
nand U6518 (N_6518,N_4498,N_4839);
nor U6519 (N_6519,N_4204,N_4856);
nand U6520 (N_6520,N_5040,N_4241);
nand U6521 (N_6521,N_5483,N_5082);
nand U6522 (N_6522,N_5718,N_4458);
nand U6523 (N_6523,N_4286,N_4453);
and U6524 (N_6524,N_4281,N_4311);
or U6525 (N_6525,N_5720,N_5915);
nand U6526 (N_6526,N_4678,N_5541);
nand U6527 (N_6527,N_4256,N_5876);
or U6528 (N_6528,N_5939,N_5648);
nor U6529 (N_6529,N_5158,N_4211);
nand U6530 (N_6530,N_5419,N_4778);
nand U6531 (N_6531,N_5275,N_5117);
nand U6532 (N_6532,N_5937,N_5415);
or U6533 (N_6533,N_4752,N_4380);
or U6534 (N_6534,N_5945,N_4642);
and U6535 (N_6535,N_5356,N_5467);
xnor U6536 (N_6536,N_5304,N_4332);
or U6537 (N_6537,N_5451,N_5074);
or U6538 (N_6538,N_5449,N_4728);
or U6539 (N_6539,N_4485,N_5980);
and U6540 (N_6540,N_5291,N_4253);
nor U6541 (N_6541,N_5025,N_5198);
or U6542 (N_6542,N_4851,N_4649);
or U6543 (N_6543,N_5497,N_5225);
nor U6544 (N_6544,N_5051,N_5477);
or U6545 (N_6545,N_4816,N_5160);
or U6546 (N_6546,N_5636,N_5786);
and U6547 (N_6547,N_4961,N_4909);
nand U6548 (N_6548,N_4328,N_4322);
xor U6549 (N_6549,N_4283,N_4722);
and U6550 (N_6550,N_4641,N_4527);
and U6551 (N_6551,N_4674,N_5060);
nor U6552 (N_6552,N_5440,N_5769);
and U6553 (N_6553,N_5321,N_5785);
nand U6554 (N_6554,N_4394,N_4711);
nor U6555 (N_6555,N_5220,N_4433);
xor U6556 (N_6556,N_4672,N_4297);
and U6557 (N_6557,N_4319,N_4932);
or U6558 (N_6558,N_5678,N_4386);
or U6559 (N_6559,N_5215,N_5516);
nand U6560 (N_6560,N_5427,N_5772);
or U6561 (N_6561,N_5398,N_4638);
xnor U6562 (N_6562,N_4478,N_4661);
nor U6563 (N_6563,N_5002,N_4889);
xor U6564 (N_6564,N_5042,N_4191);
nor U6565 (N_6565,N_5600,N_5380);
nand U6566 (N_6566,N_4547,N_5191);
or U6567 (N_6567,N_5936,N_5172);
nand U6568 (N_6568,N_4572,N_5577);
nor U6569 (N_6569,N_4717,N_4093);
and U6570 (N_6570,N_5238,N_5056);
nand U6571 (N_6571,N_4289,N_4421);
and U6572 (N_6572,N_4593,N_5923);
nand U6573 (N_6573,N_5114,N_5143);
xor U6574 (N_6574,N_5119,N_5529);
or U6575 (N_6575,N_5799,N_5572);
nor U6576 (N_6576,N_4142,N_4732);
xnor U6577 (N_6577,N_5118,N_5935);
nor U6578 (N_6578,N_4972,N_4585);
xor U6579 (N_6579,N_4991,N_5302);
and U6580 (N_6580,N_4072,N_5366);
and U6581 (N_6581,N_4730,N_5726);
or U6582 (N_6582,N_5603,N_4793);
nor U6583 (N_6583,N_5390,N_4034);
xnor U6584 (N_6584,N_4867,N_4434);
nand U6585 (N_6585,N_5258,N_4180);
nor U6586 (N_6586,N_4807,N_4052);
nand U6587 (N_6587,N_4484,N_5568);
and U6588 (N_6588,N_4143,N_4473);
nor U6589 (N_6589,N_4197,N_4811);
and U6590 (N_6590,N_5148,N_5021);
nor U6591 (N_6591,N_5479,N_5182);
and U6592 (N_6592,N_5618,N_5155);
nand U6593 (N_6593,N_5066,N_5454);
xnor U6594 (N_6594,N_4810,N_4073);
or U6595 (N_6595,N_4024,N_4475);
nor U6596 (N_6596,N_5028,N_5283);
or U6597 (N_6597,N_5108,N_4504);
nand U6598 (N_6598,N_4203,N_4103);
and U6599 (N_6599,N_5000,N_4304);
nand U6600 (N_6600,N_5824,N_4536);
or U6601 (N_6601,N_5988,N_4140);
or U6602 (N_6602,N_5694,N_4019);
nor U6603 (N_6603,N_4976,N_5679);
or U6604 (N_6604,N_4118,N_5611);
and U6605 (N_6605,N_5209,N_4300);
nor U6606 (N_6606,N_5409,N_5161);
nor U6607 (N_6607,N_4263,N_5706);
nor U6608 (N_6608,N_5306,N_5096);
and U6609 (N_6609,N_5854,N_4226);
nand U6610 (N_6610,N_4445,N_4840);
and U6611 (N_6611,N_4465,N_5305);
nand U6612 (N_6612,N_4430,N_5699);
and U6613 (N_6613,N_5183,N_4624);
xnor U6614 (N_6614,N_4815,N_4648);
nor U6615 (N_6615,N_4377,N_4894);
or U6616 (N_6616,N_4755,N_4276);
nor U6617 (N_6617,N_5702,N_5057);
and U6618 (N_6618,N_5896,N_4151);
and U6619 (N_6619,N_5274,N_4723);
or U6620 (N_6620,N_5485,N_4602);
nor U6621 (N_6621,N_4695,N_4549);
or U6622 (N_6622,N_5812,N_4074);
nor U6623 (N_6623,N_5268,N_4929);
and U6624 (N_6624,N_5818,N_5996);
nand U6625 (N_6625,N_5448,N_4178);
nor U6626 (N_6626,N_4200,N_5333);
and U6627 (N_6627,N_4566,N_5393);
nor U6628 (N_6628,N_5990,N_4773);
and U6629 (N_6629,N_5049,N_5374);
nand U6630 (N_6630,N_5617,N_5265);
or U6631 (N_6631,N_4251,N_4737);
nor U6632 (N_6632,N_5236,N_4007);
and U6633 (N_6633,N_4329,N_4274);
nor U6634 (N_6634,N_4883,N_4958);
nand U6635 (N_6635,N_4858,N_4589);
and U6636 (N_6636,N_5420,N_4213);
or U6637 (N_6637,N_5887,N_5554);
nor U6638 (N_6638,N_5241,N_4940);
nand U6639 (N_6639,N_4463,N_5052);
nor U6640 (N_6640,N_5026,N_4835);
and U6641 (N_6641,N_4352,N_5727);
nor U6642 (N_6642,N_4616,N_5899);
xnor U6643 (N_6643,N_4628,N_4088);
nor U6644 (N_6644,N_5187,N_4183);
nor U6645 (N_6645,N_4359,N_4556);
or U6646 (N_6646,N_5250,N_5184);
nand U6647 (N_6647,N_4980,N_5179);
or U6648 (N_6648,N_4782,N_5394);
nand U6649 (N_6649,N_5621,N_4947);
and U6650 (N_6650,N_4454,N_5670);
and U6651 (N_6651,N_5749,N_4525);
and U6652 (N_6652,N_4420,N_5421);
or U6653 (N_6653,N_4512,N_5682);
and U6654 (N_6654,N_4765,N_4521);
nand U6655 (N_6655,N_4081,N_5382);
xor U6656 (N_6656,N_5681,N_5523);
nand U6657 (N_6657,N_4550,N_4264);
nand U6658 (N_6658,N_5309,N_4812);
nand U6659 (N_6659,N_4503,N_4607);
nor U6660 (N_6660,N_5705,N_4409);
nand U6661 (N_6661,N_4066,N_5925);
nor U6662 (N_6662,N_5122,N_4944);
nor U6663 (N_6663,N_5979,N_4194);
or U6664 (N_6664,N_5141,N_5505);
nor U6665 (N_6665,N_4039,N_4592);
xor U6666 (N_6666,N_5677,N_5562);
and U6667 (N_6667,N_4926,N_5212);
and U6668 (N_6668,N_4687,N_5165);
or U6669 (N_6669,N_4010,N_5224);
or U6670 (N_6670,N_5132,N_4736);
and U6671 (N_6671,N_5077,N_4423);
nor U6672 (N_6672,N_4323,N_5642);
or U6673 (N_6673,N_5569,N_5458);
nand U6674 (N_6674,N_5365,N_4989);
or U6675 (N_6675,N_5586,N_4703);
nor U6676 (N_6676,N_4003,N_4966);
nand U6677 (N_6677,N_4930,N_4719);
and U6678 (N_6678,N_4284,N_4308);
and U6679 (N_6679,N_4533,N_5262);
nand U6680 (N_6680,N_4995,N_5135);
or U6681 (N_6681,N_4770,N_5766);
xor U6682 (N_6682,N_4510,N_5697);
nand U6683 (N_6683,N_5651,N_4514);
and U6684 (N_6684,N_4317,N_4971);
or U6685 (N_6685,N_5890,N_5717);
or U6686 (N_6686,N_5814,N_4012);
nand U6687 (N_6687,N_4313,N_4005);
nor U6688 (N_6688,N_4700,N_4848);
nor U6689 (N_6689,N_4403,N_4880);
nand U6690 (N_6690,N_5137,N_5299);
nor U6691 (N_6691,N_4967,N_4444);
or U6692 (N_6692,N_4714,N_5086);
nand U6693 (N_6693,N_4688,N_5027);
nor U6694 (N_6694,N_4021,N_5247);
nand U6695 (N_6695,N_5210,N_4630);
or U6696 (N_6696,N_4781,N_5296);
and U6697 (N_6697,N_5234,N_5177);
nand U6698 (N_6698,N_5375,N_4477);
or U6699 (N_6699,N_4075,N_4242);
xor U6700 (N_6700,N_5152,N_5351);
and U6701 (N_6701,N_5589,N_5526);
nor U6702 (N_6702,N_5847,N_4834);
nand U6703 (N_6703,N_5239,N_5221);
and U6704 (N_6704,N_4613,N_4275);
nor U6705 (N_6705,N_5013,N_5205);
nand U6706 (N_6706,N_4948,N_5712);
nand U6707 (N_6707,N_5325,N_4725);
nand U6708 (N_6708,N_5242,N_4977);
nor U6709 (N_6709,N_4347,N_5991);
and U6710 (N_6710,N_4790,N_5452);
nand U6711 (N_6711,N_4690,N_5591);
nor U6712 (N_6712,N_4998,N_4988);
nand U6713 (N_6713,N_4481,N_5418);
nor U6714 (N_6714,N_5634,N_5676);
xor U6715 (N_6715,N_5329,N_5638);
xor U6716 (N_6716,N_4243,N_5331);
or U6717 (N_6717,N_5295,N_5019);
nor U6718 (N_6718,N_5531,N_5099);
or U6719 (N_6719,N_5450,N_5488);
nor U6720 (N_6720,N_4518,N_5156);
or U6721 (N_6721,N_5754,N_4441);
nand U6722 (N_6722,N_4063,N_5809);
nor U6723 (N_6723,N_4535,N_4402);
or U6724 (N_6724,N_4292,N_4307);
nand U6725 (N_6725,N_4248,N_4855);
or U6726 (N_6726,N_4079,N_5379);
or U6727 (N_6727,N_5710,N_5246);
xor U6728 (N_6728,N_4599,N_4460);
and U6729 (N_6729,N_5424,N_5997);
nor U6730 (N_6730,N_5795,N_5335);
and U6731 (N_6731,N_5487,N_4899);
nor U6732 (N_6732,N_4808,N_5825);
nand U6733 (N_6733,N_5222,N_4266);
and U6734 (N_6734,N_4684,N_4654);
nor U6735 (N_6735,N_4065,N_5307);
or U6736 (N_6736,N_4573,N_5722);
nand U6737 (N_6737,N_4973,N_4391);
nand U6738 (N_6738,N_4089,N_5700);
and U6739 (N_6739,N_4520,N_4957);
or U6740 (N_6740,N_5395,N_4787);
or U6741 (N_6741,N_5008,N_4177);
nand U6742 (N_6742,N_4706,N_5551);
or U6743 (N_6743,N_5474,N_4953);
and U6744 (N_6744,N_4378,N_5976);
or U6745 (N_6745,N_4416,N_5829);
or U6746 (N_6746,N_4671,N_5030);
xor U6747 (N_6747,N_4064,N_4792);
and U6748 (N_6748,N_5848,N_4718);
and U6749 (N_6749,N_4681,N_5445);
or U6750 (N_6750,N_5518,N_4656);
nor U6751 (N_6751,N_4959,N_4795);
nor U6752 (N_6752,N_4683,N_5595);
nor U6753 (N_6753,N_4157,N_5322);
nor U6754 (N_6754,N_5863,N_4882);
or U6755 (N_6755,N_5797,N_4902);
xnor U6756 (N_6756,N_5891,N_5841);
and U6757 (N_6757,N_5794,N_5800);
or U6758 (N_6758,N_5124,N_4190);
and U6759 (N_6759,N_4257,N_4673);
nor U6760 (N_6760,N_4067,N_4040);
or U6761 (N_6761,N_5760,N_4854);
nor U6762 (N_6762,N_5453,N_5833);
and U6763 (N_6763,N_4801,N_5940);
nand U6764 (N_6764,N_4686,N_5624);
and U6765 (N_6765,N_4675,N_4900);
nor U6766 (N_6766,N_5545,N_5779);
nand U6767 (N_6767,N_5475,N_4633);
and U6768 (N_6768,N_4513,N_5790);
nand U6769 (N_6769,N_4859,N_5092);
nor U6770 (N_6770,N_4495,N_4258);
nor U6771 (N_6771,N_5147,N_5552);
nor U6772 (N_6772,N_4480,N_4236);
nor U6773 (N_6773,N_4193,N_4689);
or U6774 (N_6774,N_4006,N_5073);
nand U6775 (N_6775,N_4123,N_4597);
nand U6776 (N_6776,N_5034,N_5050);
or U6777 (N_6777,N_4053,N_5053);
nor U6778 (N_6778,N_4831,N_5608);
nand U6779 (N_6779,N_4814,N_4195);
or U6780 (N_6780,N_5609,N_4085);
nand U6781 (N_6781,N_5139,N_5508);
and U6782 (N_6782,N_4823,N_4172);
or U6783 (N_6783,N_4896,N_4381);
xor U6784 (N_6784,N_5852,N_4907);
and U6785 (N_6785,N_4145,N_5575);
nand U6786 (N_6786,N_4228,N_4057);
nor U6787 (N_6787,N_5646,N_5015);
xor U6788 (N_6788,N_5255,N_5929);
nor U6789 (N_6789,N_5909,N_4252);
and U6790 (N_6790,N_4827,N_5481);
or U6791 (N_6791,N_4916,N_4014);
nand U6792 (N_6792,N_5107,N_5127);
or U6793 (N_6793,N_4399,N_5736);
and U6794 (N_6794,N_5964,N_4050);
and U6795 (N_6795,N_4173,N_5917);
xor U6796 (N_6796,N_4663,N_4895);
nand U6797 (N_6797,N_5282,N_4187);
or U6798 (N_6798,N_4229,N_5354);
or U6799 (N_6799,N_4488,N_5928);
and U6800 (N_6800,N_5314,N_4843);
nor U6801 (N_6801,N_5157,N_4670);
and U6802 (N_6802,N_5908,N_5601);
nor U6803 (N_6803,N_5407,N_5907);
and U6804 (N_6804,N_5116,N_5033);
nor U6805 (N_6805,N_4134,N_5762);
nor U6806 (N_6806,N_5735,N_4537);
and U6807 (N_6807,N_5836,N_4704);
or U6808 (N_6808,N_5714,N_5683);
or U6809 (N_6809,N_5826,N_4523);
or U6810 (N_6810,N_4188,N_4062);
nand U6811 (N_6811,N_5914,N_5632);
nor U6812 (N_6812,N_5835,N_5125);
and U6813 (N_6813,N_4176,N_4924);
nor U6814 (N_6814,N_4234,N_5417);
and U6815 (N_6815,N_5244,N_5206);
nand U6816 (N_6816,N_5352,N_5069);
or U6817 (N_6817,N_4885,N_4132);
nand U6818 (N_6818,N_5747,N_4097);
and U6819 (N_6819,N_4469,N_5631);
nor U6820 (N_6820,N_5367,N_4412);
and U6821 (N_6821,N_4927,N_4397);
and U6822 (N_6822,N_5334,N_4500);
xnor U6823 (N_6823,N_5756,N_5588);
or U6824 (N_6824,N_5763,N_4139);
nand U6825 (N_6825,N_4424,N_5091);
xor U6826 (N_6826,N_5549,N_5643);
xnor U6827 (N_6827,N_5920,N_5721);
nor U6828 (N_6828,N_4208,N_5864);
nand U6829 (N_6829,N_4285,N_5435);
nor U6830 (N_6830,N_5338,N_4432);
or U6831 (N_6831,N_5286,N_4636);
nor U6832 (N_6832,N_5738,N_4863);
nor U6833 (N_6833,N_5093,N_4451);
nor U6834 (N_6834,N_5411,N_4584);
nor U6835 (N_6835,N_4891,N_5872);
nand U6836 (N_6836,N_4023,N_5478);
or U6837 (N_6837,N_4114,N_5639);
nand U6838 (N_6838,N_5893,N_4590);
and U6839 (N_6839,N_5423,N_4296);
nor U6840 (N_6840,N_4414,N_4144);
nand U6841 (N_6841,N_5977,N_5167);
or U6842 (N_6842,N_5573,N_4452);
nand U6843 (N_6843,N_5047,N_4138);
or U6844 (N_6844,N_4965,N_5640);
and U6845 (N_6845,N_5105,N_5843);
or U6846 (N_6846,N_5897,N_5101);
nand U6847 (N_6847,N_4698,N_4809);
xnor U6848 (N_6848,N_4786,N_5849);
or U6849 (N_6849,N_5230,N_4875);
nand U6850 (N_6850,N_5696,N_4227);
nor U6851 (N_6851,N_5867,N_4406);
nand U6852 (N_6852,N_5770,N_4828);
nor U6853 (N_6853,N_4515,N_5563);
and U6854 (N_6854,N_4544,N_5020);
nand U6855 (N_6855,N_4043,N_5290);
nor U6856 (N_6856,N_4984,N_5406);
nand U6857 (N_6857,N_4330,N_5493);
nor U6858 (N_6858,N_5413,N_5553);
xnor U6859 (N_6859,N_4733,N_5898);
nor U6860 (N_6860,N_4581,N_4366);
nand U6861 (N_6861,N_4410,N_5962);
nor U6862 (N_6862,N_4379,N_5037);
nand U6863 (N_6863,N_4221,N_5723);
or U6864 (N_6864,N_5011,N_4027);
nand U6865 (N_6865,N_5441,N_4082);
nor U6866 (N_6866,N_4355,N_5185);
or U6867 (N_6867,N_5602,N_5649);
nor U6868 (N_6868,N_4777,N_5972);
xor U6869 (N_6869,N_4161,N_5615);
or U6870 (N_6870,N_4069,N_5063);
nand U6871 (N_6871,N_5693,N_5506);
and U6872 (N_6872,N_5248,N_5827);
nor U6873 (N_6873,N_5959,N_4766);
nor U6874 (N_6874,N_5094,N_5076);
xnor U6875 (N_6875,N_4273,N_5938);
nor U6876 (N_6876,N_4288,N_5035);
or U6877 (N_6877,N_5528,N_4938);
and U6878 (N_6878,N_5428,N_4041);
and U6879 (N_6879,N_5927,N_4237);
or U6880 (N_6880,N_4111,N_4836);
and U6881 (N_6881,N_4734,N_4261);
nor U6882 (N_6882,N_4554,N_5709);
or U6883 (N_6883,N_4182,N_4101);
or U6884 (N_6884,N_4516,N_4774);
xnor U6885 (N_6885,N_5605,N_4418);
or U6886 (N_6886,N_4631,N_4710);
xor U6887 (N_6887,N_4805,N_5022);
and U6888 (N_6888,N_4845,N_5142);
nor U6889 (N_6889,N_5741,N_4487);
nor U6890 (N_6890,N_4170,N_5819);
nand U6891 (N_6891,N_4367,N_5067);
nor U6892 (N_6892,N_5784,N_5650);
and U6893 (N_6893,N_5504,N_4618);
or U6894 (N_6894,N_4492,N_5987);
nor U6895 (N_6895,N_5422,N_5048);
and U6896 (N_6896,N_4937,N_5525);
nand U6897 (N_6897,N_5373,N_5277);
or U6898 (N_6898,N_5952,N_5054);
nor U6899 (N_6899,N_4833,N_4716);
nor U6900 (N_6900,N_4682,N_4245);
nand U6901 (N_6901,N_4363,N_5431);
or U6902 (N_6902,N_4952,N_4464);
nand U6903 (N_6903,N_5471,N_4083);
nand U6904 (N_6904,N_5061,N_5134);
nor U6905 (N_6905,N_5098,N_5635);
nand U6906 (N_6906,N_4763,N_4532);
nand U6907 (N_6907,N_5164,N_5961);
and U6908 (N_6908,N_4025,N_5362);
nand U6909 (N_6909,N_4054,N_4185);
nand U6910 (N_6910,N_5946,N_5613);
and U6911 (N_6911,N_5484,N_5502);
and U6912 (N_6912,N_5079,N_4576);
nor U6913 (N_6913,N_5840,N_5003);
nor U6914 (N_6914,N_5904,N_4637);
and U6915 (N_6915,N_4582,N_5633);
and U6916 (N_6916,N_4517,N_4343);
or U6917 (N_6917,N_4877,N_4591);
and U6918 (N_6918,N_4696,N_5115);
or U6919 (N_6919,N_5667,N_4542);
or U6920 (N_6920,N_5377,N_4767);
nor U6921 (N_6921,N_5455,N_5560);
nand U6922 (N_6922,N_5429,N_5857);
nand U6923 (N_6923,N_4981,N_4122);
nor U6924 (N_6924,N_4094,N_5817);
nand U6925 (N_6925,N_4149,N_4482);
nand U6926 (N_6926,N_4529,N_5627);
nand U6927 (N_6927,N_4508,N_5916);
nand U6928 (N_6928,N_4124,N_4629);
or U6929 (N_6929,N_5456,N_4247);
nand U6930 (N_6930,N_5350,N_5192);
nor U6931 (N_6931,N_5850,N_4426);
nand U6932 (N_6932,N_5510,N_5284);
nand U6933 (N_6933,N_4901,N_4224);
and U6934 (N_6934,N_4999,N_4360);
nor U6935 (N_6935,N_5690,N_4238);
nor U6936 (N_6936,N_4772,N_5645);
xnor U6937 (N_6937,N_5778,N_4312);
nor U6938 (N_6938,N_4167,N_5006);
xnor U6939 (N_6939,N_5166,N_5261);
nor U6940 (N_6940,N_5975,N_4754);
and U6941 (N_6941,N_5012,N_4230);
and U6942 (N_6942,N_5963,N_4557);
nor U6943 (N_6943,N_5294,N_5906);
and U6944 (N_6944,N_4199,N_4413);
and U6945 (N_6945,N_5612,N_5970);
nor U6946 (N_6946,N_5217,N_4365);
or U6947 (N_6947,N_5535,N_4595);
or U6948 (N_6948,N_4461,N_5515);
and U6949 (N_6949,N_4785,N_5288);
and U6950 (N_6950,N_5501,N_5755);
and U6951 (N_6951,N_4622,N_4340);
and U6952 (N_6952,N_4667,N_4643);
or U6953 (N_6953,N_5989,N_5368);
nand U6954 (N_6954,N_5782,N_4486);
nor U6955 (N_6955,N_4740,N_4490);
or U6956 (N_6956,N_5846,N_5511);
nor U6957 (N_6957,N_5622,N_5436);
nand U6958 (N_6958,N_5669,N_4623);
nor U6959 (N_6959,N_5385,N_4679);
and U6960 (N_6960,N_4031,N_4028);
nand U6961 (N_6961,N_4303,N_5768);
nand U6962 (N_6962,N_5072,N_4739);
nor U6963 (N_6963,N_4315,N_5873);
nand U6964 (N_6964,N_5704,N_5524);
nor U6965 (N_6965,N_4729,N_4419);
nand U6966 (N_6966,N_5387,N_4148);
or U6967 (N_6967,N_4449,N_5237);
nor U6968 (N_6968,N_5263,N_4222);
or U6969 (N_6969,N_4531,N_5396);
nand U6970 (N_6970,N_5838,N_4277);
and U6971 (N_6971,N_5233,N_5199);
nor U6972 (N_6972,N_5494,N_4470);
nor U6973 (N_6973,N_5654,N_4993);
nand U6974 (N_6974,N_5353,N_4002);
nand U6975 (N_6975,N_5216,N_4382);
nor U6976 (N_6976,N_4826,N_4146);
nor U6977 (N_6977,N_4240,N_5486);
or U6978 (N_6978,N_4847,N_4282);
and U6979 (N_6979,N_5695,N_4956);
nor U6980 (N_6980,N_5476,N_5743);
and U6981 (N_6981,N_4392,N_5361);
or U6982 (N_6982,N_4120,N_4644);
xnor U6983 (N_6983,N_5796,N_5071);
nor U6984 (N_6984,N_4941,N_4507);
and U6985 (N_6985,N_5692,N_5153);
and U6986 (N_6986,N_4004,N_5579);
nand U6987 (N_6987,N_4137,N_4825);
xnor U6988 (N_6988,N_4000,N_4560);
nor U6989 (N_6989,N_5556,N_4035);
xnor U6990 (N_6990,N_5437,N_5673);
or U6991 (N_6991,N_4797,N_5982);
nand U6992 (N_6992,N_5530,N_5570);
nand U6993 (N_6993,N_4873,N_5921);
nor U6994 (N_6994,N_4270,N_5804);
nand U6995 (N_6995,N_5918,N_5672);
or U6996 (N_6996,N_4186,N_4310);
or U6997 (N_6997,N_4358,N_4562);
nor U6998 (N_6998,N_5565,N_4570);
nand U6999 (N_6999,N_4373,N_4038);
and U7000 (N_7000,N_4023,N_4884);
and U7001 (N_7001,N_4110,N_5702);
nor U7002 (N_7002,N_5222,N_4768);
and U7003 (N_7003,N_5667,N_4265);
and U7004 (N_7004,N_4059,N_4781);
nand U7005 (N_7005,N_4566,N_4611);
nor U7006 (N_7006,N_5860,N_5190);
nor U7007 (N_7007,N_5005,N_4062);
nor U7008 (N_7008,N_4280,N_4819);
nand U7009 (N_7009,N_4357,N_5011);
xnor U7010 (N_7010,N_5856,N_5631);
or U7011 (N_7011,N_5648,N_5618);
nor U7012 (N_7012,N_4458,N_4017);
xor U7013 (N_7013,N_4998,N_4888);
nor U7014 (N_7014,N_5776,N_5573);
and U7015 (N_7015,N_4343,N_4264);
xor U7016 (N_7016,N_4394,N_4528);
and U7017 (N_7017,N_5252,N_5860);
or U7018 (N_7018,N_5889,N_4487);
or U7019 (N_7019,N_5776,N_5028);
nor U7020 (N_7020,N_5213,N_5240);
or U7021 (N_7021,N_5574,N_4770);
nor U7022 (N_7022,N_5521,N_5692);
nand U7023 (N_7023,N_4922,N_4373);
nor U7024 (N_7024,N_4475,N_4328);
and U7025 (N_7025,N_4925,N_4603);
xnor U7026 (N_7026,N_4207,N_4464);
and U7027 (N_7027,N_4808,N_5840);
and U7028 (N_7028,N_5269,N_5139);
nor U7029 (N_7029,N_4908,N_4244);
nor U7030 (N_7030,N_5322,N_5671);
nor U7031 (N_7031,N_4740,N_4946);
nand U7032 (N_7032,N_5553,N_4940);
nor U7033 (N_7033,N_4085,N_4373);
xnor U7034 (N_7034,N_4411,N_5493);
nor U7035 (N_7035,N_5550,N_5034);
nand U7036 (N_7036,N_5580,N_4889);
nand U7037 (N_7037,N_4864,N_4617);
and U7038 (N_7038,N_4940,N_4837);
nor U7039 (N_7039,N_4538,N_4984);
nor U7040 (N_7040,N_4173,N_4417);
xor U7041 (N_7041,N_4513,N_4553);
or U7042 (N_7042,N_4037,N_5257);
nand U7043 (N_7043,N_4206,N_4100);
or U7044 (N_7044,N_5304,N_5449);
nor U7045 (N_7045,N_5790,N_4560);
nand U7046 (N_7046,N_4136,N_4051);
nor U7047 (N_7047,N_5976,N_4658);
nand U7048 (N_7048,N_5184,N_5963);
or U7049 (N_7049,N_4795,N_5344);
nand U7050 (N_7050,N_5021,N_5631);
or U7051 (N_7051,N_4115,N_4327);
nand U7052 (N_7052,N_5894,N_5715);
and U7053 (N_7053,N_4995,N_5035);
nand U7054 (N_7054,N_4366,N_5165);
nor U7055 (N_7055,N_4736,N_5144);
nand U7056 (N_7056,N_4790,N_5848);
nand U7057 (N_7057,N_4756,N_5297);
nand U7058 (N_7058,N_4389,N_5841);
nor U7059 (N_7059,N_5464,N_5306);
nand U7060 (N_7060,N_5162,N_4681);
nand U7061 (N_7061,N_4014,N_5243);
nor U7062 (N_7062,N_5961,N_4944);
nand U7063 (N_7063,N_5411,N_4457);
nand U7064 (N_7064,N_4137,N_4755);
and U7065 (N_7065,N_4277,N_5824);
nand U7066 (N_7066,N_5746,N_5732);
and U7067 (N_7067,N_5715,N_4064);
and U7068 (N_7068,N_5885,N_4553);
nand U7069 (N_7069,N_4151,N_5668);
and U7070 (N_7070,N_5101,N_4037);
nand U7071 (N_7071,N_5967,N_5278);
or U7072 (N_7072,N_4451,N_5753);
nor U7073 (N_7073,N_4715,N_4286);
or U7074 (N_7074,N_5896,N_4852);
or U7075 (N_7075,N_5013,N_4306);
nand U7076 (N_7076,N_4392,N_5031);
and U7077 (N_7077,N_4555,N_4102);
and U7078 (N_7078,N_5812,N_5302);
or U7079 (N_7079,N_5284,N_4889);
xor U7080 (N_7080,N_5326,N_4737);
and U7081 (N_7081,N_5659,N_5708);
and U7082 (N_7082,N_4556,N_5946);
nand U7083 (N_7083,N_5602,N_5206);
nor U7084 (N_7084,N_4101,N_4599);
or U7085 (N_7085,N_5025,N_4390);
and U7086 (N_7086,N_4075,N_4538);
and U7087 (N_7087,N_5571,N_5799);
nor U7088 (N_7088,N_5570,N_4145);
xnor U7089 (N_7089,N_4249,N_5206);
and U7090 (N_7090,N_5119,N_5842);
xnor U7091 (N_7091,N_5439,N_4141);
or U7092 (N_7092,N_5750,N_4149);
nor U7093 (N_7093,N_5508,N_4002);
nor U7094 (N_7094,N_5321,N_4580);
and U7095 (N_7095,N_5707,N_5318);
xnor U7096 (N_7096,N_4279,N_5475);
and U7097 (N_7097,N_5658,N_5594);
and U7098 (N_7098,N_4525,N_4620);
nand U7099 (N_7099,N_4170,N_5923);
nand U7100 (N_7100,N_5380,N_5714);
and U7101 (N_7101,N_5651,N_4550);
nor U7102 (N_7102,N_4366,N_4596);
nand U7103 (N_7103,N_4865,N_4745);
nor U7104 (N_7104,N_5618,N_5382);
and U7105 (N_7105,N_5014,N_5622);
or U7106 (N_7106,N_4278,N_4318);
nand U7107 (N_7107,N_4808,N_5141);
nand U7108 (N_7108,N_4562,N_5469);
or U7109 (N_7109,N_4319,N_5480);
or U7110 (N_7110,N_4383,N_5771);
nor U7111 (N_7111,N_4795,N_5909);
nor U7112 (N_7112,N_4647,N_4722);
nor U7113 (N_7113,N_4881,N_4798);
and U7114 (N_7114,N_4058,N_5407);
nand U7115 (N_7115,N_5325,N_5144);
nor U7116 (N_7116,N_5187,N_5484);
nor U7117 (N_7117,N_5406,N_4201);
nor U7118 (N_7118,N_4993,N_4154);
or U7119 (N_7119,N_5484,N_5062);
or U7120 (N_7120,N_5865,N_5326);
or U7121 (N_7121,N_5213,N_5288);
and U7122 (N_7122,N_4641,N_4261);
or U7123 (N_7123,N_5734,N_5888);
nand U7124 (N_7124,N_4282,N_4423);
nor U7125 (N_7125,N_5766,N_5885);
nor U7126 (N_7126,N_4217,N_4214);
nand U7127 (N_7127,N_5867,N_4447);
and U7128 (N_7128,N_4624,N_5771);
nand U7129 (N_7129,N_5103,N_4893);
and U7130 (N_7130,N_5318,N_4073);
or U7131 (N_7131,N_5895,N_5549);
or U7132 (N_7132,N_4885,N_5519);
or U7133 (N_7133,N_4138,N_4975);
or U7134 (N_7134,N_5177,N_5147);
xnor U7135 (N_7135,N_5605,N_5212);
and U7136 (N_7136,N_5388,N_5003);
xnor U7137 (N_7137,N_5489,N_5118);
nand U7138 (N_7138,N_4586,N_5460);
and U7139 (N_7139,N_4801,N_4661);
and U7140 (N_7140,N_4287,N_5247);
and U7141 (N_7141,N_5365,N_4587);
nand U7142 (N_7142,N_4798,N_5057);
nor U7143 (N_7143,N_4012,N_4888);
nand U7144 (N_7144,N_4147,N_5937);
nand U7145 (N_7145,N_4666,N_5899);
or U7146 (N_7146,N_5871,N_4791);
or U7147 (N_7147,N_5197,N_5793);
nor U7148 (N_7148,N_4698,N_5259);
nand U7149 (N_7149,N_4333,N_5582);
nand U7150 (N_7150,N_5112,N_5393);
nor U7151 (N_7151,N_4712,N_5231);
nand U7152 (N_7152,N_4292,N_5377);
or U7153 (N_7153,N_4689,N_5884);
xor U7154 (N_7154,N_5066,N_4933);
and U7155 (N_7155,N_5376,N_4136);
nor U7156 (N_7156,N_4144,N_5712);
nand U7157 (N_7157,N_4644,N_5352);
xnor U7158 (N_7158,N_5681,N_4383);
xnor U7159 (N_7159,N_5399,N_5659);
nand U7160 (N_7160,N_4723,N_4773);
and U7161 (N_7161,N_5258,N_4598);
nand U7162 (N_7162,N_4705,N_4074);
nand U7163 (N_7163,N_5060,N_5091);
nor U7164 (N_7164,N_5524,N_5988);
nand U7165 (N_7165,N_4236,N_4730);
nand U7166 (N_7166,N_5296,N_5003);
nor U7167 (N_7167,N_4890,N_4937);
xnor U7168 (N_7168,N_5019,N_5777);
or U7169 (N_7169,N_5665,N_4269);
or U7170 (N_7170,N_5644,N_5734);
or U7171 (N_7171,N_4932,N_4855);
xnor U7172 (N_7172,N_5679,N_5554);
nor U7173 (N_7173,N_4317,N_4425);
nor U7174 (N_7174,N_4942,N_4960);
xnor U7175 (N_7175,N_4554,N_5330);
and U7176 (N_7176,N_4942,N_5255);
nand U7177 (N_7177,N_5300,N_4875);
nor U7178 (N_7178,N_4751,N_4600);
nor U7179 (N_7179,N_4601,N_5216);
nor U7180 (N_7180,N_5610,N_5859);
or U7181 (N_7181,N_5702,N_4338);
or U7182 (N_7182,N_4139,N_4020);
or U7183 (N_7183,N_4039,N_4438);
nand U7184 (N_7184,N_5502,N_4287);
and U7185 (N_7185,N_5785,N_4814);
nand U7186 (N_7186,N_5699,N_4981);
or U7187 (N_7187,N_5709,N_4990);
nand U7188 (N_7188,N_5897,N_5978);
nand U7189 (N_7189,N_4681,N_5819);
and U7190 (N_7190,N_5172,N_5077);
nor U7191 (N_7191,N_5271,N_5837);
nor U7192 (N_7192,N_5256,N_5078);
xor U7193 (N_7193,N_4661,N_5893);
nor U7194 (N_7194,N_4914,N_4801);
or U7195 (N_7195,N_4747,N_4627);
and U7196 (N_7196,N_5510,N_4269);
or U7197 (N_7197,N_4031,N_4700);
nor U7198 (N_7198,N_5766,N_4859);
and U7199 (N_7199,N_5795,N_5481);
or U7200 (N_7200,N_5649,N_4473);
and U7201 (N_7201,N_4892,N_4455);
nor U7202 (N_7202,N_4091,N_4536);
and U7203 (N_7203,N_4634,N_4969);
and U7204 (N_7204,N_5802,N_4868);
and U7205 (N_7205,N_4869,N_5429);
and U7206 (N_7206,N_4412,N_4702);
nor U7207 (N_7207,N_5918,N_5716);
and U7208 (N_7208,N_5141,N_5215);
xnor U7209 (N_7209,N_5788,N_5911);
and U7210 (N_7210,N_5085,N_4274);
and U7211 (N_7211,N_5233,N_4915);
and U7212 (N_7212,N_5835,N_5106);
nand U7213 (N_7213,N_5812,N_4475);
nand U7214 (N_7214,N_5674,N_5584);
nand U7215 (N_7215,N_5763,N_5256);
nand U7216 (N_7216,N_5074,N_4841);
nor U7217 (N_7217,N_4062,N_5548);
xor U7218 (N_7218,N_5954,N_5119);
and U7219 (N_7219,N_5548,N_4946);
or U7220 (N_7220,N_4719,N_5441);
or U7221 (N_7221,N_5356,N_5919);
nand U7222 (N_7222,N_5963,N_4072);
nor U7223 (N_7223,N_4605,N_5533);
or U7224 (N_7224,N_5175,N_4314);
nor U7225 (N_7225,N_5658,N_5460);
and U7226 (N_7226,N_4739,N_5168);
nand U7227 (N_7227,N_4986,N_4209);
xor U7228 (N_7228,N_5385,N_5746);
nand U7229 (N_7229,N_5528,N_4840);
and U7230 (N_7230,N_4868,N_4291);
nand U7231 (N_7231,N_4083,N_5853);
xnor U7232 (N_7232,N_5107,N_5725);
nand U7233 (N_7233,N_4958,N_4222);
or U7234 (N_7234,N_5503,N_5435);
and U7235 (N_7235,N_4520,N_4272);
or U7236 (N_7236,N_5511,N_4080);
nand U7237 (N_7237,N_5011,N_4713);
xnor U7238 (N_7238,N_5968,N_5972);
nand U7239 (N_7239,N_5890,N_5519);
nor U7240 (N_7240,N_5046,N_4715);
and U7241 (N_7241,N_5263,N_5388);
nand U7242 (N_7242,N_4274,N_4319);
xnor U7243 (N_7243,N_4988,N_4435);
or U7244 (N_7244,N_4963,N_5251);
and U7245 (N_7245,N_5509,N_5360);
nand U7246 (N_7246,N_5315,N_5585);
nor U7247 (N_7247,N_5527,N_4999);
or U7248 (N_7248,N_5137,N_5594);
nor U7249 (N_7249,N_4001,N_4921);
or U7250 (N_7250,N_4573,N_5684);
and U7251 (N_7251,N_5518,N_5541);
nor U7252 (N_7252,N_5610,N_5337);
nand U7253 (N_7253,N_5050,N_5476);
nand U7254 (N_7254,N_4685,N_5223);
or U7255 (N_7255,N_4214,N_4283);
nand U7256 (N_7256,N_5047,N_4526);
or U7257 (N_7257,N_5633,N_5236);
and U7258 (N_7258,N_4512,N_5265);
nor U7259 (N_7259,N_4179,N_5413);
nand U7260 (N_7260,N_5574,N_4277);
nand U7261 (N_7261,N_5822,N_4539);
and U7262 (N_7262,N_5112,N_4483);
or U7263 (N_7263,N_4050,N_5732);
and U7264 (N_7264,N_4966,N_4266);
and U7265 (N_7265,N_4304,N_5761);
or U7266 (N_7266,N_4747,N_4197);
xor U7267 (N_7267,N_4746,N_5469);
and U7268 (N_7268,N_4751,N_4731);
nand U7269 (N_7269,N_4457,N_4488);
and U7270 (N_7270,N_4078,N_5485);
xor U7271 (N_7271,N_4713,N_5589);
and U7272 (N_7272,N_4964,N_4917);
nand U7273 (N_7273,N_5437,N_4712);
and U7274 (N_7274,N_5394,N_4161);
xnor U7275 (N_7275,N_5861,N_4181);
and U7276 (N_7276,N_4041,N_5534);
and U7277 (N_7277,N_5303,N_4460);
xor U7278 (N_7278,N_5841,N_5236);
xor U7279 (N_7279,N_5029,N_4817);
and U7280 (N_7280,N_4280,N_4071);
nand U7281 (N_7281,N_4417,N_4304);
and U7282 (N_7282,N_5785,N_4919);
nand U7283 (N_7283,N_4710,N_4958);
nand U7284 (N_7284,N_5428,N_5730);
nand U7285 (N_7285,N_5356,N_4169);
and U7286 (N_7286,N_4877,N_4331);
or U7287 (N_7287,N_5953,N_5246);
or U7288 (N_7288,N_5250,N_5522);
and U7289 (N_7289,N_4077,N_5915);
or U7290 (N_7290,N_5492,N_5430);
or U7291 (N_7291,N_5083,N_5268);
nor U7292 (N_7292,N_4013,N_4797);
or U7293 (N_7293,N_5792,N_4865);
and U7294 (N_7294,N_5922,N_5317);
nor U7295 (N_7295,N_4382,N_5564);
and U7296 (N_7296,N_4865,N_5891);
or U7297 (N_7297,N_5149,N_5321);
and U7298 (N_7298,N_4089,N_5694);
nand U7299 (N_7299,N_5932,N_4627);
or U7300 (N_7300,N_5240,N_5493);
and U7301 (N_7301,N_5357,N_4762);
xnor U7302 (N_7302,N_5127,N_4340);
and U7303 (N_7303,N_5592,N_5936);
nor U7304 (N_7304,N_4471,N_5914);
nor U7305 (N_7305,N_5175,N_4827);
nand U7306 (N_7306,N_4897,N_5014);
nand U7307 (N_7307,N_4850,N_5106);
xnor U7308 (N_7308,N_5054,N_5588);
nand U7309 (N_7309,N_4717,N_4927);
or U7310 (N_7310,N_5453,N_4652);
or U7311 (N_7311,N_5221,N_4802);
nor U7312 (N_7312,N_5315,N_4181);
xor U7313 (N_7313,N_4272,N_4997);
and U7314 (N_7314,N_4169,N_4087);
nor U7315 (N_7315,N_5336,N_4080);
nand U7316 (N_7316,N_5227,N_5774);
nor U7317 (N_7317,N_5767,N_5480);
and U7318 (N_7318,N_4937,N_5904);
nor U7319 (N_7319,N_4906,N_5471);
xor U7320 (N_7320,N_4959,N_5052);
nor U7321 (N_7321,N_5759,N_4236);
nand U7322 (N_7322,N_5169,N_4470);
xnor U7323 (N_7323,N_4689,N_5867);
nand U7324 (N_7324,N_4298,N_4621);
or U7325 (N_7325,N_4060,N_4409);
nand U7326 (N_7326,N_4096,N_5526);
nor U7327 (N_7327,N_4690,N_5462);
xnor U7328 (N_7328,N_5039,N_5484);
and U7329 (N_7329,N_4858,N_4347);
xnor U7330 (N_7330,N_5511,N_4307);
xnor U7331 (N_7331,N_4536,N_4836);
xor U7332 (N_7332,N_4659,N_4225);
and U7333 (N_7333,N_5638,N_4408);
and U7334 (N_7334,N_5955,N_4365);
nand U7335 (N_7335,N_4161,N_5322);
and U7336 (N_7336,N_5381,N_5669);
or U7337 (N_7337,N_5723,N_4088);
nor U7338 (N_7338,N_5526,N_4830);
nor U7339 (N_7339,N_5268,N_4020);
nand U7340 (N_7340,N_4446,N_4485);
xor U7341 (N_7341,N_4182,N_4020);
nand U7342 (N_7342,N_5841,N_5822);
or U7343 (N_7343,N_5868,N_4818);
and U7344 (N_7344,N_4692,N_5546);
xnor U7345 (N_7345,N_5376,N_4528);
nand U7346 (N_7346,N_4976,N_4767);
or U7347 (N_7347,N_5006,N_4311);
nand U7348 (N_7348,N_5099,N_4872);
nor U7349 (N_7349,N_4891,N_5256);
and U7350 (N_7350,N_4415,N_5656);
or U7351 (N_7351,N_4387,N_4880);
xnor U7352 (N_7352,N_4641,N_5651);
and U7353 (N_7353,N_5197,N_4242);
and U7354 (N_7354,N_4799,N_4357);
or U7355 (N_7355,N_5440,N_5422);
and U7356 (N_7356,N_4014,N_4901);
nand U7357 (N_7357,N_5569,N_4866);
nand U7358 (N_7358,N_5028,N_4463);
nor U7359 (N_7359,N_5674,N_4579);
and U7360 (N_7360,N_4195,N_5364);
and U7361 (N_7361,N_5998,N_5614);
or U7362 (N_7362,N_5608,N_5001);
nand U7363 (N_7363,N_4418,N_4185);
or U7364 (N_7364,N_4430,N_5638);
and U7365 (N_7365,N_5147,N_5335);
nor U7366 (N_7366,N_4591,N_5426);
or U7367 (N_7367,N_4282,N_5201);
or U7368 (N_7368,N_4500,N_4692);
and U7369 (N_7369,N_5090,N_5172);
and U7370 (N_7370,N_5786,N_4843);
or U7371 (N_7371,N_4296,N_5844);
and U7372 (N_7372,N_4891,N_5259);
nor U7373 (N_7373,N_4975,N_5818);
or U7374 (N_7374,N_4963,N_5549);
nand U7375 (N_7375,N_5905,N_5318);
and U7376 (N_7376,N_5685,N_5355);
or U7377 (N_7377,N_4225,N_5914);
or U7378 (N_7378,N_4077,N_4581);
and U7379 (N_7379,N_4565,N_4080);
and U7380 (N_7380,N_5311,N_5991);
nor U7381 (N_7381,N_4465,N_4147);
nor U7382 (N_7382,N_4500,N_4569);
xor U7383 (N_7383,N_5820,N_4292);
nand U7384 (N_7384,N_4601,N_5246);
nor U7385 (N_7385,N_4353,N_4974);
nand U7386 (N_7386,N_5168,N_5365);
nor U7387 (N_7387,N_5645,N_5771);
and U7388 (N_7388,N_5641,N_4510);
nor U7389 (N_7389,N_4427,N_5724);
or U7390 (N_7390,N_4077,N_5138);
nor U7391 (N_7391,N_4705,N_4962);
nor U7392 (N_7392,N_5300,N_5972);
nand U7393 (N_7393,N_4698,N_5519);
and U7394 (N_7394,N_4294,N_4301);
nor U7395 (N_7395,N_4182,N_5146);
and U7396 (N_7396,N_4967,N_4961);
nor U7397 (N_7397,N_5391,N_5927);
nand U7398 (N_7398,N_4503,N_4237);
or U7399 (N_7399,N_5044,N_4968);
or U7400 (N_7400,N_4954,N_5272);
and U7401 (N_7401,N_5468,N_5955);
and U7402 (N_7402,N_4298,N_4970);
nand U7403 (N_7403,N_5484,N_5756);
nand U7404 (N_7404,N_5442,N_5520);
nor U7405 (N_7405,N_4217,N_5227);
nand U7406 (N_7406,N_5769,N_5341);
and U7407 (N_7407,N_5969,N_5960);
and U7408 (N_7408,N_5487,N_4460);
and U7409 (N_7409,N_5669,N_4206);
or U7410 (N_7410,N_5744,N_5522);
and U7411 (N_7411,N_4498,N_5867);
nor U7412 (N_7412,N_5241,N_4073);
nor U7413 (N_7413,N_4926,N_5699);
and U7414 (N_7414,N_4937,N_5087);
nor U7415 (N_7415,N_4128,N_4468);
and U7416 (N_7416,N_5685,N_4087);
or U7417 (N_7417,N_5827,N_5903);
and U7418 (N_7418,N_5427,N_5347);
and U7419 (N_7419,N_4523,N_4862);
or U7420 (N_7420,N_5530,N_4947);
nor U7421 (N_7421,N_5099,N_5742);
nor U7422 (N_7422,N_4444,N_4697);
or U7423 (N_7423,N_4972,N_5957);
xor U7424 (N_7424,N_4436,N_4071);
nor U7425 (N_7425,N_5028,N_4121);
nor U7426 (N_7426,N_4655,N_5612);
nor U7427 (N_7427,N_5933,N_4262);
xor U7428 (N_7428,N_5630,N_4927);
nor U7429 (N_7429,N_4383,N_5412);
or U7430 (N_7430,N_4443,N_5178);
nor U7431 (N_7431,N_4047,N_4744);
or U7432 (N_7432,N_4030,N_4408);
nor U7433 (N_7433,N_5917,N_4493);
or U7434 (N_7434,N_4351,N_5413);
nor U7435 (N_7435,N_5800,N_4473);
xor U7436 (N_7436,N_4944,N_5893);
or U7437 (N_7437,N_5769,N_4389);
and U7438 (N_7438,N_5629,N_5161);
nor U7439 (N_7439,N_4042,N_5537);
nor U7440 (N_7440,N_4690,N_4022);
nor U7441 (N_7441,N_5662,N_5143);
and U7442 (N_7442,N_4080,N_5764);
or U7443 (N_7443,N_5950,N_4625);
or U7444 (N_7444,N_5644,N_5118);
and U7445 (N_7445,N_5182,N_4066);
nor U7446 (N_7446,N_5361,N_4731);
nor U7447 (N_7447,N_4808,N_4151);
nand U7448 (N_7448,N_4786,N_5778);
xnor U7449 (N_7449,N_4710,N_5795);
nor U7450 (N_7450,N_5462,N_5125);
and U7451 (N_7451,N_4515,N_5578);
nand U7452 (N_7452,N_5181,N_5938);
and U7453 (N_7453,N_5126,N_5350);
and U7454 (N_7454,N_5866,N_5015);
nor U7455 (N_7455,N_5095,N_5180);
nand U7456 (N_7456,N_4675,N_5296);
nand U7457 (N_7457,N_5831,N_4468);
nand U7458 (N_7458,N_4978,N_5741);
and U7459 (N_7459,N_4794,N_4453);
and U7460 (N_7460,N_4321,N_4971);
nor U7461 (N_7461,N_4939,N_5662);
nor U7462 (N_7462,N_4207,N_4577);
nor U7463 (N_7463,N_4486,N_4751);
and U7464 (N_7464,N_5514,N_5281);
and U7465 (N_7465,N_4179,N_5491);
xor U7466 (N_7466,N_5124,N_4997);
or U7467 (N_7467,N_4211,N_4070);
nor U7468 (N_7468,N_5439,N_5743);
nand U7469 (N_7469,N_5863,N_4542);
nand U7470 (N_7470,N_4562,N_5715);
or U7471 (N_7471,N_5687,N_5466);
and U7472 (N_7472,N_4243,N_5011);
nor U7473 (N_7473,N_5388,N_5904);
nor U7474 (N_7474,N_5861,N_5792);
nand U7475 (N_7475,N_5798,N_5096);
xnor U7476 (N_7476,N_5216,N_4109);
nand U7477 (N_7477,N_5503,N_5418);
or U7478 (N_7478,N_4351,N_5226);
or U7479 (N_7479,N_5334,N_5261);
and U7480 (N_7480,N_5442,N_5719);
nand U7481 (N_7481,N_5752,N_4753);
nand U7482 (N_7482,N_4173,N_4692);
or U7483 (N_7483,N_4908,N_4182);
nor U7484 (N_7484,N_5506,N_5994);
nand U7485 (N_7485,N_5522,N_4425);
or U7486 (N_7486,N_4579,N_4078);
and U7487 (N_7487,N_5805,N_5494);
and U7488 (N_7488,N_4017,N_4833);
xnor U7489 (N_7489,N_4805,N_5156);
and U7490 (N_7490,N_4013,N_5884);
nor U7491 (N_7491,N_4560,N_4771);
and U7492 (N_7492,N_4635,N_5955);
nand U7493 (N_7493,N_5553,N_5451);
nor U7494 (N_7494,N_4984,N_4924);
or U7495 (N_7495,N_4706,N_5276);
and U7496 (N_7496,N_4767,N_5297);
and U7497 (N_7497,N_5433,N_4151);
or U7498 (N_7498,N_5238,N_5418);
nor U7499 (N_7499,N_4102,N_4240);
nand U7500 (N_7500,N_5602,N_4489);
xnor U7501 (N_7501,N_5368,N_4929);
or U7502 (N_7502,N_4423,N_4571);
nor U7503 (N_7503,N_5878,N_4151);
or U7504 (N_7504,N_4764,N_4940);
nor U7505 (N_7505,N_4822,N_4718);
or U7506 (N_7506,N_5724,N_5202);
and U7507 (N_7507,N_5871,N_4026);
and U7508 (N_7508,N_5442,N_5610);
or U7509 (N_7509,N_5212,N_5228);
or U7510 (N_7510,N_5610,N_5690);
and U7511 (N_7511,N_4246,N_5772);
nand U7512 (N_7512,N_4646,N_4801);
nor U7513 (N_7513,N_4826,N_5870);
xnor U7514 (N_7514,N_5943,N_5046);
nor U7515 (N_7515,N_5271,N_4142);
or U7516 (N_7516,N_4900,N_4509);
or U7517 (N_7517,N_4806,N_4555);
or U7518 (N_7518,N_4496,N_5947);
nand U7519 (N_7519,N_5513,N_5229);
and U7520 (N_7520,N_4993,N_4756);
nand U7521 (N_7521,N_5518,N_5841);
or U7522 (N_7522,N_5209,N_5567);
and U7523 (N_7523,N_4191,N_5991);
xnor U7524 (N_7524,N_4687,N_4038);
nand U7525 (N_7525,N_5559,N_4985);
nand U7526 (N_7526,N_5258,N_4517);
nor U7527 (N_7527,N_5698,N_4407);
or U7528 (N_7528,N_5648,N_4534);
and U7529 (N_7529,N_4740,N_5837);
nor U7530 (N_7530,N_4002,N_4942);
nor U7531 (N_7531,N_4102,N_4583);
nor U7532 (N_7532,N_4295,N_5515);
or U7533 (N_7533,N_5395,N_5668);
nor U7534 (N_7534,N_5302,N_4960);
or U7535 (N_7535,N_5990,N_5881);
nor U7536 (N_7536,N_5177,N_5618);
and U7537 (N_7537,N_4277,N_4989);
xor U7538 (N_7538,N_5294,N_4786);
nand U7539 (N_7539,N_5168,N_5385);
and U7540 (N_7540,N_5266,N_5228);
nand U7541 (N_7541,N_4160,N_5614);
xor U7542 (N_7542,N_4476,N_4668);
and U7543 (N_7543,N_5060,N_5323);
and U7544 (N_7544,N_5401,N_5840);
and U7545 (N_7545,N_5237,N_5383);
xor U7546 (N_7546,N_4999,N_5088);
nor U7547 (N_7547,N_5923,N_4320);
xor U7548 (N_7548,N_5520,N_4883);
or U7549 (N_7549,N_4739,N_5263);
or U7550 (N_7550,N_4936,N_5152);
nor U7551 (N_7551,N_4409,N_4843);
and U7552 (N_7552,N_4492,N_5610);
nor U7553 (N_7553,N_4748,N_5916);
and U7554 (N_7554,N_4302,N_5072);
and U7555 (N_7555,N_4962,N_5681);
nor U7556 (N_7556,N_5300,N_4837);
or U7557 (N_7557,N_5101,N_4562);
nand U7558 (N_7558,N_4272,N_4229);
or U7559 (N_7559,N_4054,N_5616);
and U7560 (N_7560,N_4518,N_4987);
nand U7561 (N_7561,N_4140,N_4425);
or U7562 (N_7562,N_5395,N_5921);
and U7563 (N_7563,N_4178,N_4199);
or U7564 (N_7564,N_5688,N_4226);
xor U7565 (N_7565,N_5623,N_5394);
xnor U7566 (N_7566,N_5747,N_4132);
and U7567 (N_7567,N_5409,N_5115);
nor U7568 (N_7568,N_5441,N_4468);
xnor U7569 (N_7569,N_5236,N_5421);
or U7570 (N_7570,N_5056,N_5120);
and U7571 (N_7571,N_5981,N_5445);
and U7572 (N_7572,N_4047,N_5580);
nor U7573 (N_7573,N_4671,N_4892);
nor U7574 (N_7574,N_5517,N_5860);
nor U7575 (N_7575,N_4587,N_4834);
and U7576 (N_7576,N_4804,N_5670);
and U7577 (N_7577,N_5235,N_5211);
and U7578 (N_7578,N_5328,N_4263);
and U7579 (N_7579,N_4640,N_4155);
and U7580 (N_7580,N_5548,N_5221);
or U7581 (N_7581,N_5873,N_4662);
or U7582 (N_7582,N_4627,N_5899);
or U7583 (N_7583,N_5471,N_5582);
nor U7584 (N_7584,N_4033,N_5147);
or U7585 (N_7585,N_5890,N_4071);
and U7586 (N_7586,N_5708,N_4231);
nor U7587 (N_7587,N_4875,N_4465);
nand U7588 (N_7588,N_5525,N_4232);
nand U7589 (N_7589,N_5930,N_5093);
or U7590 (N_7590,N_5748,N_4284);
or U7591 (N_7591,N_4111,N_4436);
nor U7592 (N_7592,N_5817,N_4741);
and U7593 (N_7593,N_4416,N_5731);
or U7594 (N_7594,N_4023,N_5123);
or U7595 (N_7595,N_4804,N_5561);
nand U7596 (N_7596,N_5559,N_5042);
and U7597 (N_7597,N_5502,N_4499);
nor U7598 (N_7598,N_4042,N_4698);
nor U7599 (N_7599,N_5549,N_5825);
nor U7600 (N_7600,N_5878,N_5160);
nand U7601 (N_7601,N_5914,N_4903);
nand U7602 (N_7602,N_5972,N_5215);
nand U7603 (N_7603,N_5075,N_5388);
nand U7604 (N_7604,N_5844,N_5505);
and U7605 (N_7605,N_5207,N_5401);
nand U7606 (N_7606,N_5609,N_4089);
or U7607 (N_7607,N_4779,N_5291);
xor U7608 (N_7608,N_4827,N_5809);
nor U7609 (N_7609,N_4131,N_4737);
nor U7610 (N_7610,N_4098,N_5956);
or U7611 (N_7611,N_4041,N_4095);
and U7612 (N_7612,N_5131,N_4214);
nor U7613 (N_7613,N_4321,N_4246);
nand U7614 (N_7614,N_4760,N_4285);
or U7615 (N_7615,N_5915,N_5641);
nor U7616 (N_7616,N_4262,N_5225);
nor U7617 (N_7617,N_4676,N_4394);
nor U7618 (N_7618,N_5833,N_4165);
nand U7619 (N_7619,N_5554,N_4525);
nor U7620 (N_7620,N_5045,N_4179);
nor U7621 (N_7621,N_4324,N_4076);
nor U7622 (N_7622,N_4597,N_4088);
nor U7623 (N_7623,N_4994,N_4693);
nand U7624 (N_7624,N_5325,N_4994);
nor U7625 (N_7625,N_4331,N_4695);
nor U7626 (N_7626,N_5682,N_4147);
nand U7627 (N_7627,N_5297,N_5712);
and U7628 (N_7628,N_5161,N_5277);
and U7629 (N_7629,N_5039,N_5365);
or U7630 (N_7630,N_5423,N_4364);
or U7631 (N_7631,N_4830,N_5091);
nor U7632 (N_7632,N_4182,N_5873);
nor U7633 (N_7633,N_5467,N_5698);
nor U7634 (N_7634,N_4878,N_4388);
or U7635 (N_7635,N_5834,N_4230);
xnor U7636 (N_7636,N_5526,N_5864);
nor U7637 (N_7637,N_4475,N_4937);
nand U7638 (N_7638,N_4405,N_4757);
nand U7639 (N_7639,N_5230,N_5827);
and U7640 (N_7640,N_5223,N_5482);
nand U7641 (N_7641,N_4790,N_5673);
xor U7642 (N_7642,N_5193,N_4232);
and U7643 (N_7643,N_5470,N_5203);
and U7644 (N_7644,N_4114,N_5611);
and U7645 (N_7645,N_4745,N_4844);
or U7646 (N_7646,N_5313,N_4934);
nand U7647 (N_7647,N_4072,N_5321);
nor U7648 (N_7648,N_5164,N_4511);
nand U7649 (N_7649,N_5381,N_4478);
xnor U7650 (N_7650,N_4383,N_5714);
and U7651 (N_7651,N_4784,N_5194);
or U7652 (N_7652,N_4645,N_4825);
nor U7653 (N_7653,N_5518,N_5990);
and U7654 (N_7654,N_5115,N_5932);
nor U7655 (N_7655,N_5539,N_5830);
nand U7656 (N_7656,N_5522,N_5823);
and U7657 (N_7657,N_4382,N_5045);
or U7658 (N_7658,N_5625,N_5650);
nand U7659 (N_7659,N_5155,N_4151);
or U7660 (N_7660,N_4027,N_5964);
nand U7661 (N_7661,N_4574,N_4859);
or U7662 (N_7662,N_4596,N_4759);
nand U7663 (N_7663,N_4688,N_5620);
nor U7664 (N_7664,N_5169,N_4541);
nand U7665 (N_7665,N_4666,N_5492);
nor U7666 (N_7666,N_4074,N_4337);
nand U7667 (N_7667,N_4940,N_5970);
or U7668 (N_7668,N_4143,N_5377);
nor U7669 (N_7669,N_4734,N_4460);
and U7670 (N_7670,N_4885,N_4140);
nand U7671 (N_7671,N_4905,N_5148);
nand U7672 (N_7672,N_4988,N_4841);
and U7673 (N_7673,N_4241,N_5177);
or U7674 (N_7674,N_5063,N_5419);
or U7675 (N_7675,N_4199,N_4344);
or U7676 (N_7676,N_5670,N_4717);
nor U7677 (N_7677,N_5158,N_5825);
or U7678 (N_7678,N_5414,N_5021);
or U7679 (N_7679,N_5085,N_5188);
and U7680 (N_7680,N_5047,N_5273);
or U7681 (N_7681,N_4574,N_4395);
or U7682 (N_7682,N_5523,N_4738);
nand U7683 (N_7683,N_5891,N_5954);
or U7684 (N_7684,N_4826,N_4299);
nor U7685 (N_7685,N_5683,N_4440);
or U7686 (N_7686,N_4051,N_4139);
nor U7687 (N_7687,N_4296,N_4680);
or U7688 (N_7688,N_4950,N_4863);
and U7689 (N_7689,N_4727,N_4856);
nand U7690 (N_7690,N_4410,N_4658);
or U7691 (N_7691,N_4173,N_4206);
or U7692 (N_7692,N_5494,N_5632);
nand U7693 (N_7693,N_5841,N_5193);
nor U7694 (N_7694,N_4348,N_4501);
nand U7695 (N_7695,N_4739,N_5687);
xnor U7696 (N_7696,N_5573,N_4416);
and U7697 (N_7697,N_5644,N_5773);
nand U7698 (N_7698,N_4705,N_5397);
nor U7699 (N_7699,N_4659,N_5101);
nor U7700 (N_7700,N_4474,N_5468);
nand U7701 (N_7701,N_5332,N_4870);
or U7702 (N_7702,N_5592,N_5825);
nand U7703 (N_7703,N_5965,N_5279);
or U7704 (N_7704,N_5820,N_4719);
nand U7705 (N_7705,N_4399,N_5612);
or U7706 (N_7706,N_5534,N_5759);
xor U7707 (N_7707,N_4307,N_4644);
nand U7708 (N_7708,N_4600,N_4759);
or U7709 (N_7709,N_4533,N_5349);
xor U7710 (N_7710,N_4160,N_5541);
or U7711 (N_7711,N_5876,N_5870);
nor U7712 (N_7712,N_5206,N_4866);
and U7713 (N_7713,N_4042,N_4238);
nand U7714 (N_7714,N_5328,N_5508);
nand U7715 (N_7715,N_5874,N_5227);
nor U7716 (N_7716,N_5469,N_4386);
nor U7717 (N_7717,N_4364,N_5118);
nor U7718 (N_7718,N_4929,N_5614);
and U7719 (N_7719,N_4089,N_5380);
and U7720 (N_7720,N_4245,N_5952);
or U7721 (N_7721,N_5745,N_4397);
and U7722 (N_7722,N_5248,N_5395);
nand U7723 (N_7723,N_5297,N_5219);
and U7724 (N_7724,N_4973,N_5992);
or U7725 (N_7725,N_5868,N_4627);
xor U7726 (N_7726,N_5315,N_4034);
or U7727 (N_7727,N_4684,N_5806);
or U7728 (N_7728,N_5076,N_4878);
nor U7729 (N_7729,N_5395,N_5779);
nor U7730 (N_7730,N_4901,N_5346);
or U7731 (N_7731,N_4661,N_4491);
nor U7732 (N_7732,N_4658,N_4197);
or U7733 (N_7733,N_5509,N_4541);
nand U7734 (N_7734,N_5703,N_5358);
nor U7735 (N_7735,N_5113,N_4500);
nand U7736 (N_7736,N_5887,N_5965);
nand U7737 (N_7737,N_4530,N_5760);
nand U7738 (N_7738,N_5308,N_5370);
and U7739 (N_7739,N_4856,N_4125);
nand U7740 (N_7740,N_4536,N_4820);
or U7741 (N_7741,N_5702,N_4745);
or U7742 (N_7742,N_5057,N_4766);
nand U7743 (N_7743,N_5619,N_4676);
nand U7744 (N_7744,N_4500,N_4702);
nand U7745 (N_7745,N_5823,N_5561);
or U7746 (N_7746,N_4826,N_5583);
nand U7747 (N_7747,N_4395,N_5267);
and U7748 (N_7748,N_5806,N_5355);
nand U7749 (N_7749,N_4554,N_4165);
or U7750 (N_7750,N_5850,N_5566);
nor U7751 (N_7751,N_5662,N_5723);
nand U7752 (N_7752,N_5883,N_4241);
nand U7753 (N_7753,N_4654,N_5379);
nor U7754 (N_7754,N_5409,N_5401);
or U7755 (N_7755,N_5671,N_4160);
nand U7756 (N_7756,N_4028,N_4125);
nand U7757 (N_7757,N_4797,N_4282);
and U7758 (N_7758,N_4445,N_5675);
or U7759 (N_7759,N_4869,N_5312);
and U7760 (N_7760,N_4087,N_4362);
and U7761 (N_7761,N_4224,N_5308);
and U7762 (N_7762,N_5024,N_4574);
nor U7763 (N_7763,N_4538,N_5548);
nand U7764 (N_7764,N_5634,N_5932);
xnor U7765 (N_7765,N_5482,N_4290);
nor U7766 (N_7766,N_5006,N_5788);
or U7767 (N_7767,N_5318,N_4173);
nand U7768 (N_7768,N_4157,N_5769);
or U7769 (N_7769,N_5821,N_5950);
nand U7770 (N_7770,N_5401,N_4254);
nand U7771 (N_7771,N_5901,N_5775);
and U7772 (N_7772,N_5186,N_5210);
nor U7773 (N_7773,N_4611,N_5125);
or U7774 (N_7774,N_5889,N_4507);
xnor U7775 (N_7775,N_5222,N_5342);
and U7776 (N_7776,N_5894,N_5733);
nand U7777 (N_7777,N_4908,N_4053);
nor U7778 (N_7778,N_5289,N_4593);
nand U7779 (N_7779,N_4118,N_4578);
nand U7780 (N_7780,N_5522,N_4058);
or U7781 (N_7781,N_5063,N_4348);
nand U7782 (N_7782,N_5081,N_4067);
or U7783 (N_7783,N_5757,N_4391);
nor U7784 (N_7784,N_4070,N_5943);
and U7785 (N_7785,N_4949,N_5601);
nand U7786 (N_7786,N_5620,N_5403);
nor U7787 (N_7787,N_5475,N_4362);
or U7788 (N_7788,N_5427,N_5139);
and U7789 (N_7789,N_4009,N_4892);
nor U7790 (N_7790,N_5222,N_5150);
nor U7791 (N_7791,N_4093,N_5612);
nand U7792 (N_7792,N_5765,N_4816);
xnor U7793 (N_7793,N_5076,N_5852);
nor U7794 (N_7794,N_4935,N_5643);
nor U7795 (N_7795,N_4227,N_5178);
or U7796 (N_7796,N_5420,N_5307);
and U7797 (N_7797,N_5812,N_5670);
and U7798 (N_7798,N_5654,N_5868);
xor U7799 (N_7799,N_4260,N_4200);
nor U7800 (N_7800,N_4626,N_5130);
and U7801 (N_7801,N_5398,N_5443);
nand U7802 (N_7802,N_5607,N_4767);
nor U7803 (N_7803,N_5986,N_5014);
or U7804 (N_7804,N_5997,N_4527);
and U7805 (N_7805,N_4993,N_5086);
nand U7806 (N_7806,N_5371,N_5151);
and U7807 (N_7807,N_5807,N_4829);
nor U7808 (N_7808,N_4368,N_5868);
and U7809 (N_7809,N_4968,N_5026);
xnor U7810 (N_7810,N_4371,N_4574);
nand U7811 (N_7811,N_4380,N_5709);
and U7812 (N_7812,N_4112,N_5600);
nand U7813 (N_7813,N_5660,N_5126);
nor U7814 (N_7814,N_5206,N_5251);
nor U7815 (N_7815,N_4309,N_4120);
xor U7816 (N_7816,N_4625,N_5521);
nand U7817 (N_7817,N_4534,N_5421);
nand U7818 (N_7818,N_5846,N_5907);
or U7819 (N_7819,N_5510,N_5662);
and U7820 (N_7820,N_4261,N_5624);
xnor U7821 (N_7821,N_5107,N_4954);
nand U7822 (N_7822,N_5556,N_5826);
nand U7823 (N_7823,N_5798,N_4794);
and U7824 (N_7824,N_4668,N_5023);
nand U7825 (N_7825,N_5290,N_4409);
and U7826 (N_7826,N_5291,N_5227);
and U7827 (N_7827,N_4654,N_4143);
nor U7828 (N_7828,N_5292,N_4169);
nor U7829 (N_7829,N_5991,N_5225);
nor U7830 (N_7830,N_4182,N_5283);
and U7831 (N_7831,N_5595,N_5772);
or U7832 (N_7832,N_4701,N_5877);
or U7833 (N_7833,N_5260,N_5471);
or U7834 (N_7834,N_4258,N_4097);
or U7835 (N_7835,N_5952,N_5296);
and U7836 (N_7836,N_5764,N_5454);
and U7837 (N_7837,N_4723,N_5086);
nor U7838 (N_7838,N_5374,N_4535);
and U7839 (N_7839,N_4903,N_4504);
or U7840 (N_7840,N_5654,N_4171);
xnor U7841 (N_7841,N_4245,N_4342);
and U7842 (N_7842,N_5542,N_5103);
and U7843 (N_7843,N_5635,N_5365);
nor U7844 (N_7844,N_5616,N_5279);
nand U7845 (N_7845,N_5798,N_4070);
nand U7846 (N_7846,N_5655,N_5316);
or U7847 (N_7847,N_4001,N_4183);
xor U7848 (N_7848,N_5633,N_5040);
nor U7849 (N_7849,N_5356,N_4915);
nor U7850 (N_7850,N_4403,N_4041);
nand U7851 (N_7851,N_5494,N_4995);
xor U7852 (N_7852,N_5431,N_5550);
nand U7853 (N_7853,N_4588,N_5945);
nor U7854 (N_7854,N_4154,N_4155);
or U7855 (N_7855,N_4795,N_5043);
xnor U7856 (N_7856,N_4046,N_4062);
or U7857 (N_7857,N_5506,N_5993);
and U7858 (N_7858,N_4508,N_5372);
nand U7859 (N_7859,N_5940,N_4904);
nor U7860 (N_7860,N_4976,N_4562);
xnor U7861 (N_7861,N_4293,N_4453);
and U7862 (N_7862,N_5831,N_4638);
nand U7863 (N_7863,N_4973,N_5709);
and U7864 (N_7864,N_4518,N_4799);
or U7865 (N_7865,N_5914,N_5815);
nand U7866 (N_7866,N_5111,N_5575);
xor U7867 (N_7867,N_5504,N_4881);
and U7868 (N_7868,N_5910,N_4819);
and U7869 (N_7869,N_4830,N_5049);
or U7870 (N_7870,N_4467,N_4125);
nand U7871 (N_7871,N_4390,N_4168);
nor U7872 (N_7872,N_4492,N_5228);
nor U7873 (N_7873,N_5716,N_5643);
nor U7874 (N_7874,N_4607,N_4723);
or U7875 (N_7875,N_4538,N_4817);
and U7876 (N_7876,N_4497,N_5560);
and U7877 (N_7877,N_5571,N_4860);
or U7878 (N_7878,N_4338,N_5001);
or U7879 (N_7879,N_5744,N_5480);
or U7880 (N_7880,N_5155,N_4848);
and U7881 (N_7881,N_4966,N_4321);
and U7882 (N_7882,N_5262,N_4408);
and U7883 (N_7883,N_4359,N_5422);
xor U7884 (N_7884,N_4803,N_4767);
and U7885 (N_7885,N_4713,N_4216);
nand U7886 (N_7886,N_4443,N_5076);
nor U7887 (N_7887,N_4102,N_5519);
nand U7888 (N_7888,N_5036,N_5804);
nor U7889 (N_7889,N_4503,N_4957);
or U7890 (N_7890,N_4863,N_4944);
or U7891 (N_7891,N_4905,N_5431);
nor U7892 (N_7892,N_5126,N_5940);
and U7893 (N_7893,N_5199,N_5660);
nor U7894 (N_7894,N_4128,N_4607);
or U7895 (N_7895,N_4804,N_4698);
and U7896 (N_7896,N_5201,N_4281);
or U7897 (N_7897,N_4685,N_4536);
nand U7898 (N_7898,N_4871,N_5364);
or U7899 (N_7899,N_5992,N_5677);
nand U7900 (N_7900,N_5761,N_5694);
xor U7901 (N_7901,N_4126,N_5633);
and U7902 (N_7902,N_5831,N_4431);
nand U7903 (N_7903,N_5898,N_5235);
nand U7904 (N_7904,N_4641,N_4233);
and U7905 (N_7905,N_4573,N_5889);
or U7906 (N_7906,N_4253,N_5047);
and U7907 (N_7907,N_4929,N_5837);
or U7908 (N_7908,N_5509,N_4553);
xnor U7909 (N_7909,N_4750,N_4622);
and U7910 (N_7910,N_4474,N_4461);
xnor U7911 (N_7911,N_5434,N_4044);
and U7912 (N_7912,N_5705,N_5179);
nor U7913 (N_7913,N_4972,N_4075);
nand U7914 (N_7914,N_4218,N_4594);
and U7915 (N_7915,N_4162,N_4737);
nand U7916 (N_7916,N_4348,N_5219);
or U7917 (N_7917,N_5579,N_4993);
and U7918 (N_7918,N_5755,N_4082);
nor U7919 (N_7919,N_5585,N_5184);
nor U7920 (N_7920,N_5176,N_4891);
nor U7921 (N_7921,N_5649,N_5819);
nand U7922 (N_7922,N_4680,N_5559);
or U7923 (N_7923,N_5312,N_4683);
nand U7924 (N_7924,N_4615,N_5584);
and U7925 (N_7925,N_5963,N_4060);
or U7926 (N_7926,N_4333,N_4622);
and U7927 (N_7927,N_5045,N_4541);
and U7928 (N_7928,N_4781,N_4408);
nor U7929 (N_7929,N_4802,N_4944);
xor U7930 (N_7930,N_5774,N_4359);
or U7931 (N_7931,N_4010,N_5205);
or U7932 (N_7932,N_4410,N_5289);
or U7933 (N_7933,N_5044,N_4873);
and U7934 (N_7934,N_4956,N_4563);
nand U7935 (N_7935,N_5732,N_5967);
nor U7936 (N_7936,N_4029,N_4902);
or U7937 (N_7937,N_5435,N_4418);
nand U7938 (N_7938,N_4833,N_4291);
and U7939 (N_7939,N_4883,N_4361);
nor U7940 (N_7940,N_4509,N_4402);
or U7941 (N_7941,N_5289,N_4380);
or U7942 (N_7942,N_4779,N_4924);
nand U7943 (N_7943,N_5921,N_4988);
and U7944 (N_7944,N_4748,N_4971);
and U7945 (N_7945,N_5704,N_4936);
or U7946 (N_7946,N_4264,N_5689);
or U7947 (N_7947,N_4703,N_5742);
nand U7948 (N_7948,N_4907,N_4094);
and U7949 (N_7949,N_5270,N_4747);
nor U7950 (N_7950,N_4214,N_4025);
and U7951 (N_7951,N_4596,N_5632);
and U7952 (N_7952,N_4286,N_4954);
and U7953 (N_7953,N_4230,N_4040);
and U7954 (N_7954,N_4548,N_4961);
nor U7955 (N_7955,N_4671,N_4039);
nand U7956 (N_7956,N_4295,N_4939);
xor U7957 (N_7957,N_4975,N_5347);
xnor U7958 (N_7958,N_4655,N_4962);
or U7959 (N_7959,N_4946,N_5723);
and U7960 (N_7960,N_4745,N_5324);
and U7961 (N_7961,N_4101,N_4308);
nand U7962 (N_7962,N_4867,N_4768);
nor U7963 (N_7963,N_5653,N_5595);
or U7964 (N_7964,N_4970,N_5217);
and U7965 (N_7965,N_4609,N_4921);
or U7966 (N_7966,N_5724,N_4669);
and U7967 (N_7967,N_4683,N_4796);
or U7968 (N_7968,N_4098,N_5733);
nand U7969 (N_7969,N_5762,N_5425);
nand U7970 (N_7970,N_4312,N_4620);
and U7971 (N_7971,N_4257,N_4576);
xnor U7972 (N_7972,N_4712,N_4877);
nand U7973 (N_7973,N_4308,N_5343);
nor U7974 (N_7974,N_4273,N_4517);
and U7975 (N_7975,N_5229,N_5608);
and U7976 (N_7976,N_4490,N_5397);
nand U7977 (N_7977,N_5583,N_4058);
and U7978 (N_7978,N_5587,N_5555);
or U7979 (N_7979,N_5225,N_5234);
xor U7980 (N_7980,N_4883,N_5214);
nor U7981 (N_7981,N_4313,N_4357);
or U7982 (N_7982,N_5983,N_4957);
xor U7983 (N_7983,N_5374,N_5863);
and U7984 (N_7984,N_5596,N_5412);
and U7985 (N_7985,N_4446,N_4824);
and U7986 (N_7986,N_5239,N_5795);
nand U7987 (N_7987,N_5842,N_4361);
nor U7988 (N_7988,N_5707,N_4887);
and U7989 (N_7989,N_4500,N_5905);
xor U7990 (N_7990,N_5058,N_5341);
nor U7991 (N_7991,N_4124,N_5185);
or U7992 (N_7992,N_4001,N_5361);
and U7993 (N_7993,N_4194,N_5821);
nand U7994 (N_7994,N_4575,N_5327);
nor U7995 (N_7995,N_5617,N_5181);
nor U7996 (N_7996,N_4583,N_4049);
nor U7997 (N_7997,N_4015,N_5654);
and U7998 (N_7998,N_4342,N_5219);
xnor U7999 (N_7999,N_4524,N_5799);
nand U8000 (N_8000,N_6607,N_6089);
and U8001 (N_8001,N_7872,N_6101);
or U8002 (N_8002,N_6361,N_6469);
or U8003 (N_8003,N_7418,N_7640);
or U8004 (N_8004,N_6477,N_7396);
and U8005 (N_8005,N_6969,N_7860);
nand U8006 (N_8006,N_7850,N_7447);
nand U8007 (N_8007,N_7730,N_7903);
or U8008 (N_8008,N_7681,N_7463);
or U8009 (N_8009,N_6524,N_6783);
nor U8010 (N_8010,N_7653,N_7778);
and U8011 (N_8011,N_7987,N_6757);
xor U8012 (N_8012,N_7928,N_6127);
and U8013 (N_8013,N_6136,N_7289);
and U8014 (N_8014,N_7702,N_6146);
and U8015 (N_8015,N_6784,N_7094);
and U8016 (N_8016,N_7774,N_7971);
or U8017 (N_8017,N_6055,N_7646);
nor U8018 (N_8018,N_7602,N_7853);
nor U8019 (N_8019,N_7397,N_6228);
nand U8020 (N_8020,N_7726,N_7487);
nor U8021 (N_8021,N_6486,N_6043);
nor U8022 (N_8022,N_7376,N_6384);
or U8023 (N_8023,N_7632,N_6370);
nand U8024 (N_8024,N_7331,N_7773);
and U8025 (N_8025,N_7270,N_7758);
or U8026 (N_8026,N_6295,N_7312);
nand U8027 (N_8027,N_6404,N_6603);
nor U8028 (N_8028,N_7931,N_6674);
nand U8029 (N_8029,N_7859,N_6706);
nor U8030 (N_8030,N_7349,N_6391);
and U8031 (N_8031,N_7736,N_6655);
nor U8032 (N_8032,N_7658,N_7122);
nor U8033 (N_8033,N_6693,N_6464);
xor U8034 (N_8034,N_6004,N_6258);
nand U8035 (N_8035,N_6418,N_7033);
nand U8036 (N_8036,N_7454,N_6651);
or U8037 (N_8037,N_7152,N_7252);
nor U8038 (N_8038,N_6183,N_7556);
nand U8039 (N_8039,N_6664,N_6601);
and U8040 (N_8040,N_6402,N_6897);
and U8041 (N_8041,N_7827,N_6102);
and U8042 (N_8042,N_7406,N_7886);
and U8043 (N_8043,N_6881,N_7919);
or U8044 (N_8044,N_7916,N_7108);
nand U8045 (N_8045,N_7683,N_7475);
and U8046 (N_8046,N_7223,N_7912);
nand U8047 (N_8047,N_7274,N_6491);
xnor U8048 (N_8048,N_6821,N_7548);
nor U8049 (N_8049,N_6452,N_6448);
nor U8050 (N_8050,N_7044,N_7842);
and U8051 (N_8051,N_7756,N_7442);
xnor U8052 (N_8052,N_6993,N_6346);
nor U8053 (N_8053,N_6538,N_7911);
or U8054 (N_8054,N_6846,N_7216);
or U8055 (N_8055,N_6378,N_6949);
nor U8056 (N_8056,N_7114,N_6744);
or U8057 (N_8057,N_6720,N_7573);
xor U8058 (N_8058,N_7455,N_7298);
nand U8059 (N_8059,N_7932,N_7608);
and U8060 (N_8060,N_7539,N_6454);
nor U8061 (N_8061,N_7569,N_6581);
nand U8062 (N_8062,N_7205,N_6342);
xor U8063 (N_8063,N_6044,N_6589);
and U8064 (N_8064,N_7106,N_6755);
or U8065 (N_8065,N_6040,N_7494);
or U8066 (N_8066,N_7235,N_7535);
or U8067 (N_8067,N_7023,N_6272);
or U8068 (N_8068,N_7765,N_6928);
and U8069 (N_8069,N_7124,N_6809);
nor U8070 (N_8070,N_7170,N_7846);
nor U8071 (N_8071,N_6833,N_6773);
or U8072 (N_8072,N_7669,N_6215);
nor U8073 (N_8073,N_6910,N_6944);
nor U8074 (N_8074,N_7924,N_7220);
and U8075 (N_8075,N_6147,N_6943);
and U8076 (N_8076,N_7137,N_6261);
or U8077 (N_8077,N_6165,N_6340);
or U8078 (N_8078,N_6734,N_6294);
xor U8079 (N_8079,N_7028,N_7690);
nor U8080 (N_8080,N_7670,N_7282);
nor U8081 (N_8081,N_7481,N_6758);
and U8082 (N_8082,N_7510,N_7682);
nand U8083 (N_8083,N_6770,N_6523);
and U8084 (N_8084,N_6826,N_7404);
nor U8085 (N_8085,N_6775,N_6869);
and U8086 (N_8086,N_6593,N_6729);
and U8087 (N_8087,N_7657,N_7322);
nor U8088 (N_8088,N_7836,N_6592);
or U8089 (N_8089,N_7930,N_7389);
or U8090 (N_8090,N_7361,N_7750);
or U8091 (N_8091,N_6798,N_7874);
nand U8092 (N_8092,N_6386,N_7807);
nand U8093 (N_8093,N_6439,N_6108);
or U8094 (N_8094,N_7590,N_7526);
xor U8095 (N_8095,N_7787,N_7645);
and U8096 (N_8096,N_7966,N_6400);
nor U8097 (N_8097,N_7741,N_7667);
or U8098 (N_8098,N_6360,N_6266);
or U8099 (N_8099,N_6742,N_7009);
nor U8100 (N_8100,N_7808,N_6345);
or U8101 (N_8101,N_7259,N_7474);
or U8102 (N_8102,N_6210,N_7528);
nand U8103 (N_8103,N_6575,N_6251);
xor U8104 (N_8104,N_6242,N_7062);
nand U8105 (N_8105,N_6181,N_7275);
or U8106 (N_8106,N_6236,N_7473);
and U8107 (N_8107,N_6564,N_7049);
nand U8108 (N_8108,N_7105,N_6283);
nand U8109 (N_8109,N_7140,N_7003);
nand U8110 (N_8110,N_7277,N_7985);
xor U8111 (N_8111,N_7878,N_6190);
nor U8112 (N_8112,N_7844,N_7079);
nand U8113 (N_8113,N_6313,N_7318);
and U8114 (N_8114,N_6791,N_7231);
or U8115 (N_8115,N_6895,N_6768);
nand U8116 (N_8116,N_6098,N_7438);
nor U8117 (N_8117,N_7253,N_7129);
and U8118 (N_8118,N_7156,N_6354);
xnor U8119 (N_8119,N_6094,N_6740);
and U8120 (N_8120,N_7477,N_7663);
xor U8121 (N_8121,N_6460,N_6647);
nand U8122 (N_8122,N_7221,N_7939);
nor U8123 (N_8123,N_7629,N_6657);
and U8124 (N_8124,N_7247,N_6233);
and U8125 (N_8125,N_6492,N_6580);
and U8126 (N_8126,N_7290,N_6224);
nand U8127 (N_8127,N_7697,N_7999);
nand U8128 (N_8128,N_7772,N_6608);
nand U8129 (N_8129,N_7135,N_7570);
nand U8130 (N_8130,N_7696,N_7190);
or U8131 (N_8131,N_6972,N_7305);
nand U8132 (N_8132,N_6625,N_7525);
xor U8133 (N_8133,N_7278,N_7695);
or U8134 (N_8134,N_7990,N_6894);
nand U8135 (N_8135,N_7013,N_7864);
nor U8136 (N_8136,N_7032,N_6296);
nand U8137 (N_8137,N_7411,N_7965);
and U8138 (N_8138,N_6304,N_6597);
nor U8139 (N_8139,N_7926,N_6079);
xor U8140 (N_8140,N_6663,N_7934);
or U8141 (N_8141,N_7018,N_6947);
nor U8142 (N_8142,N_6551,N_7245);
nand U8143 (N_8143,N_7465,N_7011);
and U8144 (N_8144,N_6925,N_7962);
or U8145 (N_8145,N_6095,N_7008);
or U8146 (N_8146,N_7947,N_7536);
or U8147 (N_8147,N_7288,N_6462);
or U8148 (N_8148,N_7858,N_6186);
and U8149 (N_8149,N_6899,N_6029);
nor U8150 (N_8150,N_7036,N_7350);
nand U8151 (N_8151,N_7359,N_6362);
nor U8152 (N_8152,N_6927,N_6543);
nand U8153 (N_8153,N_6868,N_6844);
and U8154 (N_8154,N_7711,N_6009);
nor U8155 (N_8155,N_6479,N_7056);
or U8156 (N_8156,N_7542,N_6828);
and U8157 (N_8157,N_6010,N_7345);
or U8158 (N_8158,N_6811,N_6907);
and U8159 (N_8159,N_6694,N_7889);
nor U8160 (N_8160,N_6877,N_6099);
nand U8161 (N_8161,N_6222,N_6167);
nor U8162 (N_8162,N_7642,N_6013);
and U8163 (N_8163,N_7800,N_6633);
or U8164 (N_8164,N_6748,N_7311);
nand U8165 (N_8165,N_6053,N_7577);
and U8166 (N_8166,N_7978,N_6586);
or U8167 (N_8167,N_6987,N_6964);
and U8168 (N_8168,N_7565,N_7347);
or U8169 (N_8169,N_6379,N_6428);
xor U8170 (N_8170,N_7552,N_7019);
or U8171 (N_8171,N_6105,N_7664);
nor U8172 (N_8172,N_6217,N_6561);
nand U8173 (N_8173,N_6414,N_7143);
or U8174 (N_8174,N_7904,N_6872);
nand U8175 (N_8175,N_7177,N_7784);
or U8176 (N_8176,N_6025,N_7902);
and U8177 (N_8177,N_7740,N_6364);
or U8178 (N_8178,N_7202,N_7944);
and U8179 (N_8179,N_6245,N_6387);
or U8180 (N_8180,N_6137,N_7405);
and U8181 (N_8181,N_7352,N_6471);
and U8182 (N_8182,N_7224,N_7964);
nand U8183 (N_8183,N_6014,N_7401);
or U8184 (N_8184,N_6918,N_6435);
and U8185 (N_8185,N_7716,N_7644);
nand U8186 (N_8186,N_6810,N_7203);
and U8187 (N_8187,N_7309,N_6749);
nor U8188 (N_8188,N_7641,N_7792);
nand U8189 (N_8189,N_7899,N_7377);
nor U8190 (N_8190,N_6500,N_6307);
xor U8191 (N_8191,N_6198,N_6312);
nor U8192 (N_8192,N_6660,N_6801);
xor U8193 (N_8193,N_6047,N_7648);
nor U8194 (N_8194,N_6549,N_6206);
and U8195 (N_8195,N_7634,N_7849);
nand U8196 (N_8196,N_6638,N_7768);
nor U8197 (N_8197,N_7212,N_7483);
or U8198 (N_8198,N_6271,N_6830);
and U8199 (N_8199,N_7597,N_6725);
nor U8200 (N_8200,N_7561,N_6743);
or U8201 (N_8201,N_7575,N_6730);
nor U8202 (N_8202,N_6466,N_7456);
nand U8203 (N_8203,N_6503,N_6106);
and U8204 (N_8204,N_7698,N_6936);
and U8205 (N_8205,N_6531,N_7144);
or U8206 (N_8206,N_7211,N_7102);
or U8207 (N_8207,N_6838,N_6789);
nand U8208 (N_8208,N_6957,N_6058);
xor U8209 (N_8209,N_7954,N_6498);
nand U8210 (N_8210,N_7166,N_7790);
or U8211 (N_8211,N_7898,N_7650);
or U8212 (N_8212,N_6401,N_7198);
nor U8213 (N_8213,N_6124,N_6259);
nand U8214 (N_8214,N_6445,N_7433);
xor U8215 (N_8215,N_7169,N_6546);
xor U8216 (N_8216,N_7559,N_7611);
nand U8217 (N_8217,N_7625,N_6036);
nand U8218 (N_8218,N_6563,N_6287);
or U8219 (N_8219,N_6336,N_7533);
nand U8220 (N_8220,N_6458,N_7328);
and U8221 (N_8221,N_6028,N_7386);
nor U8222 (N_8222,N_7714,N_7250);
or U8223 (N_8223,N_6722,N_6558);
xor U8224 (N_8224,N_6858,N_7039);
xnor U8225 (N_8225,N_7598,N_7030);
or U8226 (N_8226,N_7724,N_7233);
or U8227 (N_8227,N_7436,N_6178);
or U8228 (N_8228,N_6268,N_6686);
nand U8229 (N_8229,N_7343,N_7004);
and U8230 (N_8230,N_7489,N_7427);
and U8231 (N_8231,N_7178,N_7199);
or U8232 (N_8232,N_6082,N_7668);
or U8233 (N_8233,N_6472,N_6637);
nor U8234 (N_8234,N_7785,N_6073);
nor U8235 (N_8235,N_6999,N_6382);
or U8236 (N_8236,N_7313,N_7006);
nand U8237 (N_8237,N_7603,N_6548);
or U8238 (N_8238,N_6049,N_7638);
nand U8239 (N_8239,N_6166,N_6335);
and U8240 (N_8240,N_6065,N_6118);
xnor U8241 (N_8241,N_7676,N_7053);
nand U8242 (N_8242,N_6220,N_7010);
xor U8243 (N_8243,N_6041,N_7993);
nand U8244 (N_8244,N_6156,N_7496);
nand U8245 (N_8245,N_7449,N_7434);
nor U8246 (N_8246,N_6636,N_7339);
nand U8247 (N_8247,N_7720,N_6171);
or U8248 (N_8248,N_7798,N_7234);
and U8249 (N_8249,N_6642,N_6254);
nor U8250 (N_8250,N_7459,N_6062);
nor U8251 (N_8251,N_6022,N_7895);
nand U8252 (N_8252,N_6656,N_7867);
nand U8253 (N_8253,N_6679,N_6015);
and U8254 (N_8254,N_7751,N_7795);
xnor U8255 (N_8255,N_7174,N_6978);
or U8256 (N_8256,N_6527,N_6483);
or U8257 (N_8257,N_6953,N_6511);
or U8258 (N_8258,N_6349,N_6727);
xnor U8259 (N_8259,N_6455,N_7677);
nor U8260 (N_8260,N_6060,N_7194);
nor U8261 (N_8261,N_7977,N_7315);
nand U8262 (N_8262,N_6199,N_7117);
nand U8263 (N_8263,N_7232,N_6680);
nand U8264 (N_8264,N_6504,N_7478);
nor U8265 (N_8265,N_7165,N_6780);
and U8266 (N_8266,N_6805,N_7617);
nor U8267 (N_8267,N_7090,N_7107);
and U8268 (N_8268,N_6322,N_6032);
xor U8269 (N_8269,N_6115,N_6356);
nor U8270 (N_8270,N_7951,N_6068);
or U8271 (N_8271,N_7593,N_6735);
xor U8272 (N_8272,N_7420,N_7066);
and U8273 (N_8273,N_7953,N_7430);
and U8274 (N_8274,N_7596,N_7703);
and U8275 (N_8275,N_6061,N_7024);
nor U8276 (N_8276,N_7186,N_6717);
nand U8277 (N_8277,N_7471,N_6209);
and U8278 (N_8278,N_7851,N_7722);
nand U8279 (N_8279,N_6884,N_6473);
nor U8280 (N_8280,N_7257,N_7995);
nand U8281 (N_8281,N_6457,N_6248);
nand U8282 (N_8282,N_6176,N_6667);
xor U8283 (N_8283,N_7337,N_6359);
or U8284 (N_8284,N_6157,N_6970);
and U8285 (N_8285,N_7422,N_6232);
and U8286 (N_8286,N_7627,N_6684);
and U8287 (N_8287,N_7885,N_7545);
nor U8288 (N_8288,N_6870,N_6474);
nor U8289 (N_8289,N_7745,N_7937);
nand U8290 (N_8290,N_7656,N_7390);
nand U8291 (N_8291,N_6604,N_7378);
nor U8292 (N_8292,N_6343,N_6395);
nor U8293 (N_8293,N_6624,N_6393);
nor U8294 (N_8294,N_7151,N_7530);
or U8295 (N_8295,N_7109,N_6977);
nand U8296 (N_8296,N_7310,N_7027);
or U8297 (N_8297,N_6622,N_6290);
and U8298 (N_8298,N_6196,N_6595);
xnor U8299 (N_8299,N_7128,N_7414);
nor U8300 (N_8300,N_6974,N_7168);
xnor U8301 (N_8301,N_6929,N_7067);
nand U8302 (N_8302,N_7779,N_7097);
and U8303 (N_8303,N_6066,N_7409);
or U8304 (N_8304,N_7078,N_6606);
and U8305 (N_8305,N_7208,N_7585);
nand U8306 (N_8306,N_6279,N_6247);
xor U8307 (N_8307,N_7149,N_7909);
xnor U8308 (N_8308,N_7821,N_7729);
nor U8309 (N_8309,N_6415,N_7891);
nand U8310 (N_8310,N_7723,N_6021);
nand U8311 (N_8311,N_6540,N_6634);
and U8312 (N_8312,N_6886,N_6467);
or U8313 (N_8313,N_7046,N_7896);
nand U8314 (N_8314,N_7517,N_6797);
or U8315 (N_8315,N_7111,N_6229);
and U8316 (N_8316,N_6713,N_6839);
nand U8317 (N_8317,N_6803,N_7863);
and U8318 (N_8318,N_6726,N_6644);
nor U8319 (N_8319,N_7957,N_7982);
and U8320 (N_8320,N_7016,N_7666);
xnor U8321 (N_8321,N_6705,N_7193);
nor U8322 (N_8322,N_6933,N_6611);
and U8323 (N_8323,N_6623,N_7907);
nor U8324 (N_8324,N_7141,N_7292);
or U8325 (N_8325,N_7468,N_6935);
or U8326 (N_8326,N_7267,N_7484);
and U8327 (N_8327,N_6760,N_6308);
nor U8328 (N_8328,N_7370,N_7497);
and U8329 (N_8329,N_7823,N_7647);
or U8330 (N_8330,N_6630,N_6596);
xor U8331 (N_8331,N_7412,N_6373);
nand U8332 (N_8332,N_6912,N_6003);
nor U8333 (N_8333,N_6085,N_6747);
and U8334 (N_8334,N_7197,N_7413);
nand U8335 (N_8335,N_7960,N_7635);
or U8336 (N_8336,N_6024,N_7848);
or U8337 (N_8337,N_7622,N_6175);
and U8338 (N_8338,N_7678,N_6100);
xnor U8339 (N_8339,N_6390,N_7334);
or U8340 (N_8340,N_7123,N_7240);
xnor U8341 (N_8341,N_6450,N_6554);
and U8342 (N_8342,N_7520,N_6121);
or U8343 (N_8343,N_6347,N_6109);
nor U8344 (N_8344,N_6613,N_6012);
nand U8345 (N_8345,N_7938,N_6185);
or U8346 (N_8346,N_6582,N_7881);
xnor U8347 (N_8347,N_7341,N_7540);
and U8348 (N_8348,N_6239,N_6505);
or U8349 (N_8349,N_6182,N_6513);
nor U8350 (N_8350,N_6357,N_6218);
nor U8351 (N_8351,N_7824,N_7665);
and U8352 (N_8352,N_6767,N_6535);
nor U8353 (N_8353,N_6406,N_6148);
xor U8354 (N_8354,N_7900,N_6501);
and U8355 (N_8355,N_6337,N_7158);
nor U8356 (N_8356,N_7748,N_7776);
nand U8357 (N_8357,N_6752,N_7184);
nand U8358 (N_8358,N_7618,N_6643);
and U8359 (N_8359,N_7777,N_7280);
or U8360 (N_8360,N_7811,N_6681);
or U8361 (N_8361,N_6097,N_6380);
xnor U8362 (N_8362,N_7616,N_7547);
or U8363 (N_8363,N_7155,N_6880);
xor U8364 (N_8364,N_6698,N_7271);
xor U8365 (N_8365,N_6204,N_7639);
nand U8366 (N_8366,N_7572,N_7351);
or U8367 (N_8367,N_6184,N_6096);
nand U8368 (N_8368,N_6434,N_7883);
nor U8369 (N_8369,N_7069,N_7366);
nand U8370 (N_8370,N_7188,N_6541);
nand U8371 (N_8371,N_7374,N_7794);
xor U8372 (N_8372,N_7191,N_6806);
or U8373 (N_8373,N_6116,N_7762);
xor U8374 (N_8374,N_7380,N_7061);
or U8375 (N_8375,N_6619,N_7356);
nand U8376 (N_8376,N_6235,N_6265);
nand U8377 (N_8377,N_7451,N_6676);
and U8378 (N_8378,N_6280,N_7324);
and U8379 (N_8379,N_7687,N_6800);
and U8380 (N_8380,N_7710,N_7956);
and U8381 (N_8381,N_6733,N_7981);
or U8382 (N_8382,N_7104,N_7052);
or U8383 (N_8383,N_6288,N_7708);
or U8384 (N_8384,N_7375,N_6971);
xnor U8385 (N_8385,N_7148,N_7335);
or U8386 (N_8386,N_7237,N_7012);
and U8387 (N_8387,N_7415,N_6901);
or U8388 (N_8388,N_7888,N_6348);
and U8389 (N_8389,N_6609,N_7828);
and U8390 (N_8390,N_6352,N_7537);
nand U8391 (N_8391,N_7834,N_6632);
nand U8392 (N_8392,N_7908,N_6497);
nand U8393 (N_8393,N_6107,N_6782);
nand U8394 (N_8394,N_6263,N_6951);
and U8395 (N_8395,N_6162,N_6990);
nor U8396 (N_8396,N_6793,N_6699);
and U8397 (N_8397,N_6994,N_6134);
or U8398 (N_8398,N_7945,N_7467);
nor U8399 (N_8399,N_6916,N_6711);
or U8400 (N_8400,N_6695,N_7336);
nor U8401 (N_8401,N_6570,N_7684);
xnor U8402 (N_8402,N_7796,N_6986);
xor U8403 (N_8403,N_6683,N_6834);
and U8404 (N_8404,N_7501,N_7991);
nor U8405 (N_8405,N_6804,N_6104);
nand U8406 (N_8406,N_7073,N_6188);
or U8407 (N_8407,N_6143,N_6598);
nand U8408 (N_8408,N_6984,N_7273);
nand U8409 (N_8409,N_7970,N_7180);
or U8410 (N_8410,N_6366,N_7580);
or U8411 (N_8411,N_6154,N_6052);
or U8412 (N_8412,N_6090,N_7486);
nand U8413 (N_8413,N_6753,N_6367);
or U8414 (N_8414,N_7544,N_7431);
nand U8415 (N_8415,N_6072,N_6700);
nor U8416 (N_8416,N_7428,N_6653);
xnor U8417 (N_8417,N_7865,N_7880);
xnor U8418 (N_8418,N_7226,N_7862);
nand U8419 (N_8419,N_7890,N_7940);
and U8420 (N_8420,N_6552,N_6103);
or U8421 (N_8421,N_7228,N_7959);
xnor U8422 (N_8422,N_7379,N_7814);
and U8423 (N_8423,N_6620,N_7717);
nand U8424 (N_8424,N_7949,N_6835);
or U8425 (N_8425,N_6305,N_7769);
nor U8426 (N_8426,N_7727,N_7980);
and U8427 (N_8427,N_6256,N_6075);
or U8428 (N_8428,N_7296,N_7571);
xnor U8429 (N_8429,N_6091,N_6216);
and U8430 (N_8430,N_7239,N_6076);
and U8431 (N_8431,N_7464,N_6904);
or U8432 (N_8432,N_7020,N_7164);
and U8433 (N_8433,N_6955,N_6278);
and U8434 (N_8434,N_6276,N_6763);
and U8435 (N_8435,N_6692,N_7157);
or U8436 (N_8436,N_6484,N_6771);
or U8437 (N_8437,N_7421,N_6422);
xor U8438 (N_8438,N_7576,N_6341);
xnor U8439 (N_8439,N_7000,N_6855);
nand U8440 (N_8440,N_7996,N_7913);
nor U8441 (N_8441,N_7014,N_6539);
nand U8442 (N_8442,N_7917,N_6081);
nand U8443 (N_8443,N_7813,N_6602);
nand U8444 (N_8444,N_7905,N_6463);
nand U8445 (N_8445,N_7163,N_6030);
nand U8446 (N_8446,N_7134,N_7251);
and U8447 (N_8447,N_6584,N_7096);
nand U8448 (N_8448,N_7568,N_6954);
nand U8449 (N_8449,N_7815,N_7495);
xor U8450 (N_8450,N_6790,N_7532);
nor U8451 (N_8451,N_6908,N_7457);
nand U8452 (N_8452,N_6646,N_6225);
nor U8453 (N_8453,N_7192,N_7870);
and U8454 (N_8454,N_7272,N_6197);
and U8455 (N_8455,N_6291,N_6723);
nor U8456 (N_8456,N_7115,N_7812);
and U8457 (N_8457,N_6662,N_6120);
nand U8458 (N_8458,N_7387,N_7215);
nand U8459 (N_8459,N_7975,N_7749);
nand U8460 (N_8460,N_6392,N_7589);
and U8461 (N_8461,N_7498,N_6863);
or U8462 (N_8462,N_7038,N_7839);
nor U8463 (N_8463,N_7121,N_7643);
or U8464 (N_8464,N_7534,N_6201);
or U8465 (N_8465,N_6368,N_7175);
nand U8466 (N_8466,N_6119,N_6528);
xor U8467 (N_8467,N_6310,N_7118);
and U8468 (N_8468,N_7265,N_6436);
and U8469 (N_8469,N_7424,N_7743);
or U8470 (N_8470,N_6817,N_6111);
nand U8471 (N_8471,N_6802,N_7967);
or U8472 (N_8472,N_6475,N_6145);
nor U8473 (N_8473,N_6149,N_7041);
nor U8474 (N_8474,N_7021,N_7920);
nand U8475 (N_8475,N_6051,N_7139);
or U8476 (N_8476,N_7725,N_7040);
nor U8477 (N_8477,N_7417,N_7225);
nor U8478 (N_8478,N_7286,N_6982);
nor U8479 (N_8479,N_7515,N_6084);
xnor U8480 (N_8480,N_6150,N_6856);
and U8481 (N_8481,N_7416,N_6932);
and U8482 (N_8482,N_6244,N_7935);
and U8483 (N_8483,N_7789,N_6441);
xnor U8484 (N_8484,N_7269,N_6117);
and U8485 (N_8485,N_6728,N_6572);
and U8486 (N_8486,N_6113,N_6226);
nand U8487 (N_8487,N_6764,N_6732);
nor U8488 (N_8488,N_6442,N_6691);
nand U8489 (N_8489,N_6665,N_7113);
and U8490 (N_8490,N_6187,N_7302);
and U8491 (N_8491,N_7142,N_6427);
or U8492 (N_8492,N_7599,N_6861);
and U8493 (N_8493,N_6666,N_6125);
and U8494 (N_8494,N_6945,N_7739);
and U8495 (N_8495,N_6419,N_6823);
and U8496 (N_8496,N_7372,N_7029);
nor U8497 (N_8497,N_6520,N_6917);
nand U8498 (N_8498,N_6281,N_7894);
nor U8499 (N_8499,N_7488,N_6779);
and U8500 (N_8500,N_6652,N_7974);
and U8501 (N_8501,N_6286,N_6840);
nor U8502 (N_8502,N_7918,N_7804);
nor U8503 (N_8503,N_7847,N_6416);
nand U8504 (N_8504,N_7555,N_7402);
or U8505 (N_8505,N_7747,N_6237);
nor U8506 (N_8506,N_7963,N_6542);
xnor U8507 (N_8507,N_6578,N_6567);
nor U8508 (N_8508,N_7213,N_6083);
or U8509 (N_8509,N_6514,N_6566);
nor U8510 (N_8510,N_7476,N_7043);
nor U8511 (N_8511,N_7173,N_7531);
nand U8512 (N_8512,N_6616,N_6939);
nor U8513 (N_8513,N_7660,N_7448);
or U8514 (N_8514,N_6997,N_7435);
xor U8515 (N_8515,N_6292,N_7493);
or U8516 (N_8516,N_6064,N_6948);
nor U8517 (N_8517,N_6142,N_6736);
nor U8518 (N_8518,N_7901,N_6942);
xor U8519 (N_8519,N_6574,N_6319);
nand U8520 (N_8520,N_7994,N_7089);
nand U8521 (N_8521,N_6983,N_6715);
nand U8522 (N_8522,N_7988,N_6063);
nand U8523 (N_8523,N_6299,N_6410);
nor U8524 (N_8524,N_7976,N_6923);
and U8525 (N_8525,N_6853,N_7673);
xor U8526 (N_8526,N_7461,N_7160);
or U8527 (N_8527,N_7080,N_6144);
and U8528 (N_8528,N_6007,N_6996);
nand U8529 (N_8529,N_6848,N_6866);
and U8530 (N_8530,N_7521,N_6708);
xnor U8531 (N_8531,N_6635,N_6260);
and U8532 (N_8532,N_7299,N_7450);
or U8533 (N_8533,N_7636,N_6913);
nor U8534 (N_8534,N_7574,N_7992);
or U8535 (N_8535,N_6885,N_6980);
xnor U8536 (N_8536,N_6252,N_7230);
or U8537 (N_8537,N_7588,N_6685);
nand U8538 (N_8538,N_7783,N_7838);
nand U8539 (N_8539,N_6191,N_6650);
nand U8540 (N_8540,N_6078,N_6394);
xnor U8541 (N_8541,N_6122,N_7432);
or U8542 (N_8542,N_7738,N_6326);
nor U8543 (N_8543,N_6363,N_7466);
or U8544 (N_8544,N_7519,N_7301);
nor U8545 (N_8545,N_6591,N_7718);
and U8546 (N_8546,N_7958,N_7055);
or U8547 (N_8547,N_6960,N_7159);
and U8548 (N_8548,N_6898,N_7112);
or U8549 (N_8549,N_7822,N_6417);
and U8550 (N_8550,N_7624,N_6493);
or U8551 (N_8551,N_6069,N_6027);
or U8552 (N_8552,N_6938,N_7172);
and U8553 (N_8553,N_7546,N_7983);
or U8554 (N_8554,N_7835,N_6536);
and U8555 (N_8555,N_7754,N_6837);
and U8556 (N_8556,N_6243,N_6140);
nand U8557 (N_8557,N_6214,N_7470);
nor U8558 (N_8558,N_6000,N_6461);
and U8559 (N_8559,N_7527,N_7293);
nor U8560 (N_8560,N_7241,N_7554);
or U8561 (N_8561,N_7605,N_7025);
or U8562 (N_8562,N_7026,N_6440);
and U8563 (N_8563,N_6555,N_7699);
xnor U8564 (N_8564,N_7780,N_6219);
and U8565 (N_8565,N_7482,N_6019);
and U8566 (N_8566,N_7353,N_6559);
and U8567 (N_8567,N_7070,N_6696);
and U8568 (N_8568,N_7419,N_6544);
and U8569 (N_8569,N_7941,N_7766);
nor U8570 (N_8570,N_6277,N_6822);
nor U8571 (N_8571,N_7704,N_7759);
nor U8572 (N_8572,N_6883,N_7054);
nor U8573 (N_8573,N_7162,N_6327);
nor U8574 (N_8574,N_6480,N_7408);
or U8575 (N_8575,N_7098,N_7381);
nor U8576 (N_8576,N_6878,N_7692);
or U8577 (N_8577,N_7264,N_7887);
and U8578 (N_8578,N_7176,N_7972);
xnor U8579 (N_8579,N_7831,N_6697);
and U8580 (N_8580,N_7358,N_7303);
nand U8581 (N_8581,N_6172,N_6533);
nand U8582 (N_8582,N_7179,N_7788);
or U8583 (N_8583,N_6914,N_6961);
xnor U8584 (N_8584,N_6842,N_6323);
nor U8585 (N_8585,N_7391,N_6282);
xor U8586 (N_8586,N_6815,N_7437);
nand U8587 (N_8587,N_7833,N_7746);
and U8588 (N_8588,N_7065,N_7150);
and U8589 (N_8589,N_7136,N_7426);
or U8590 (N_8590,N_6718,N_6832);
nor U8591 (N_8591,N_6042,N_7187);
xnor U8592 (N_8592,N_7562,N_7087);
nor U8593 (N_8593,N_6179,N_7384);
and U8594 (N_8594,N_6565,N_7626);
xor U8595 (N_8595,N_6016,N_7512);
or U8596 (N_8596,N_6375,N_6139);
nor U8597 (N_8597,N_6930,N_7587);
and U8598 (N_8598,N_7857,N_7120);
nand U8599 (N_8599,N_6864,N_7204);
nor U8600 (N_8600,N_7505,N_7342);
nand U8601 (N_8601,N_6412,N_7705);
and U8602 (N_8602,N_7266,N_7440);
and U8603 (N_8603,N_6114,N_6151);
nand U8604 (N_8604,N_7445,N_6774);
and U8605 (N_8605,N_7781,N_7227);
nand U8606 (N_8606,N_6888,N_6739);
or U8607 (N_8607,N_7316,N_7592);
xnor U8608 (N_8608,N_6919,N_6046);
nor U8609 (N_8609,N_6639,N_6130);
nor U8610 (N_8610,N_7731,N_6459);
nand U8611 (N_8611,N_6673,N_7291);
and U8612 (N_8612,N_6270,N_7661);
and U8613 (N_8613,N_6485,N_7679);
nor U8614 (N_8614,N_6751,N_7915);
and U8615 (N_8615,N_7877,N_6425);
nand U8616 (N_8616,N_6397,N_7385);
or U8617 (N_8617,N_7154,N_7258);
or U8618 (N_8618,N_7734,N_6355);
nor U8619 (N_8619,N_6577,N_7146);
or U8620 (N_8620,N_7686,N_6035);
and U8621 (N_8621,N_6794,N_6973);
or U8622 (N_8622,N_6034,N_6194);
nor U8623 (N_8623,N_7817,N_7897);
nand U8624 (N_8624,N_7671,N_6795);
or U8625 (N_8625,N_6212,N_6257);
or U8626 (N_8626,N_6583,N_7764);
nor U8627 (N_8627,N_7701,N_6138);
and U8628 (N_8628,N_6262,N_7394);
or U8629 (N_8629,N_6631,N_6998);
nor U8630 (N_8630,N_7085,N_6807);
or U8631 (N_8631,N_6371,N_7238);
or U8632 (N_8632,N_6174,N_7492);
nor U8633 (N_8633,N_7852,N_7145);
nor U8634 (N_8634,N_7832,N_6617);
nand U8635 (N_8635,N_6020,N_7619);
nor U8636 (N_8636,N_7961,N_6829);
nand U8637 (N_8637,N_6813,N_6776);
nor U8638 (N_8638,N_6429,N_7500);
nor U8639 (N_8639,N_6761,N_6495);
and U8640 (N_8640,N_7218,N_7595);
or U8641 (N_8641,N_7508,N_6135);
nand U8642 (N_8642,N_7893,N_6001);
and U8643 (N_8643,N_7214,N_7383);
and U8644 (N_8644,N_6850,N_7007);
and U8645 (N_8645,N_7399,N_7805);
nand U8646 (N_8646,N_6873,N_7869);
or U8647 (N_8647,N_6508,N_7441);
nand U8648 (N_8648,N_6300,N_7538);
or U8649 (N_8649,N_7200,N_6274);
or U8650 (N_8650,N_7300,N_7952);
nor U8651 (N_8651,N_6374,N_7392);
and U8652 (N_8652,N_7630,N_7721);
nand U8653 (N_8653,N_7855,N_6211);
nor U8654 (N_8654,N_7942,N_6796);
and U8655 (N_8655,N_6859,N_7771);
and U8656 (N_8656,N_6153,N_7873);
xor U8657 (N_8657,N_6437,N_6376);
nand U8658 (N_8658,N_7210,N_6490);
or U8659 (N_8659,N_6926,N_6309);
nand U8660 (N_8660,N_6321,N_6267);
or U8661 (N_8661,N_6470,N_6170);
nand U8662 (N_8662,N_6339,N_6965);
nand U8663 (N_8663,N_6967,N_7001);
nand U8664 (N_8664,N_6077,N_6478);
nor U8665 (N_8665,N_6519,N_7304);
and U8666 (N_8666,N_7084,N_6372);
xnor U8667 (N_8667,N_7925,N_7446);
and U8668 (N_8668,N_7943,N_7439);
nor U8669 (N_8669,N_6887,N_6906);
or U8670 (N_8670,N_6093,N_7306);
or U8671 (N_8671,N_6334,N_6909);
and U8672 (N_8672,N_6671,N_6875);
xnor U8673 (N_8673,N_6921,N_6857);
nor U8674 (N_8674,N_6369,N_7255);
or U8675 (N_8675,N_7830,N_7308);
and U8676 (N_8676,N_6314,N_7936);
nand U8677 (N_8677,N_6365,N_7551);
nand U8678 (N_8678,N_7791,N_7601);
nor U8679 (N_8679,N_6737,N_7479);
nor U8680 (N_8680,N_7816,N_7884);
or U8681 (N_8681,N_7591,N_7005);
nor U8682 (N_8682,N_6284,N_7034);
nand U8683 (N_8683,N_7284,N_7077);
nand U8684 (N_8684,N_6891,N_7649);
nand U8685 (N_8685,N_6521,N_7153);
nor U8686 (N_8686,N_7083,N_7075);
nand U8687 (N_8687,N_7509,N_6195);
or U8688 (N_8688,N_7071,N_6958);
nand U8689 (N_8689,N_6273,N_6628);
xor U8690 (N_8690,N_6668,N_6388);
nor U8691 (N_8691,N_7689,N_7058);
or U8692 (N_8692,N_6594,N_6731);
or U8693 (N_8693,N_6344,N_7367);
or U8694 (N_8694,N_6302,N_6297);
and U8695 (N_8695,N_7933,N_6351);
or U8696 (N_8696,N_6550,N_6023);
and U8697 (N_8697,N_7579,N_7183);
nor U8698 (N_8698,N_6092,N_6039);
and U8699 (N_8699,N_6221,N_7969);
nand U8700 (N_8700,N_6433,N_7979);
nand U8701 (N_8701,N_6843,N_6289);
nand U8702 (N_8702,N_7680,N_6956);
nand U8703 (N_8703,N_6738,N_6488);
nand U8704 (N_8704,N_7543,N_7057);
or U8705 (N_8705,N_6621,N_7797);
or U8706 (N_8706,N_7841,N_6529);
and U8707 (N_8707,N_7346,N_6750);
nand U8708 (N_8708,N_6230,N_7125);
and U8709 (N_8709,N_6446,N_6408);
xor U8710 (N_8710,N_7922,N_6976);
and U8711 (N_8711,N_6223,N_6385);
nor U8712 (N_8712,N_7499,N_7567);
nor U8713 (N_8713,N_6205,N_7048);
nor U8714 (N_8714,N_7578,N_6516);
xor U8715 (N_8715,N_6088,N_7189);
and U8716 (N_8716,N_7693,N_7480);
or U8717 (N_8717,N_6754,N_6002);
xor U8718 (N_8718,N_7081,N_6865);
nor U8719 (N_8719,N_7244,N_7209);
nand U8720 (N_8720,N_6250,N_7843);
nor U8721 (N_8721,N_7845,N_6610);
nand U8722 (N_8722,N_6778,N_7610);
and U8723 (N_8723,N_7329,N_6502);
or U8724 (N_8724,N_7330,N_7829);
and U8725 (N_8725,N_6557,N_6048);
nand U8726 (N_8726,N_7452,N_6963);
xnor U8727 (N_8727,N_6645,N_6241);
or U8728 (N_8728,N_7360,N_6534);
nor U8729 (N_8729,N_6164,N_7037);
and U8730 (N_8730,N_6413,N_7606);
or U8731 (N_8731,N_6189,N_6054);
xor U8732 (N_8732,N_6383,N_7806);
and U8733 (N_8733,N_6525,N_6011);
nand U8734 (N_8734,N_7042,N_6249);
xor U8735 (N_8735,N_6537,N_7604);
nand U8736 (N_8736,N_7719,N_7088);
and U8737 (N_8737,N_6545,N_6661);
xnor U8738 (N_8738,N_7130,N_7167);
and U8739 (N_8739,N_7735,N_7672);
xnor U8740 (N_8740,N_7256,N_6759);
xnor U8741 (N_8741,N_7249,N_7325);
nor U8742 (N_8742,N_6772,N_6315);
nand U8743 (N_8743,N_6903,N_7760);
and U8744 (N_8744,N_6820,N_7490);
or U8745 (N_8745,N_7217,N_6426);
nor U8746 (N_8746,N_7327,N_6614);
nor U8747 (N_8747,N_6173,N_7091);
xnor U8748 (N_8748,N_7820,N_7263);
and U8749 (N_8749,N_7246,N_6553);
nand U8750 (N_8750,N_6332,N_6507);
and U8751 (N_8751,N_6481,N_7314);
nand U8752 (N_8752,N_6799,N_6227);
or U8753 (N_8753,N_6882,N_6407);
nand U8754 (N_8754,N_7685,N_7229);
nor U8755 (N_8755,N_7694,N_7986);
or U8756 (N_8756,N_6396,N_7400);
nand U8757 (N_8757,N_6159,N_7876);
or U8758 (N_8758,N_6968,N_6818);
nor U8759 (N_8759,N_6423,N_6569);
nand U8760 (N_8760,N_6285,N_6871);
and U8761 (N_8761,N_6152,N_7594);
or U8762 (N_8762,N_6985,N_7276);
nand U8763 (N_8763,N_6133,N_6132);
or U8764 (N_8764,N_6629,N_7927);
or U8765 (N_8765,N_7775,N_7799);
and U8766 (N_8766,N_7333,N_6975);
and U8767 (N_8767,N_6449,N_6006);
nor U8768 (N_8768,N_7132,N_7388);
and U8769 (N_8769,N_7092,N_7652);
nand U8770 (N_8770,N_7837,N_6465);
or U8771 (N_8771,N_7818,N_7294);
and U8772 (N_8772,N_6432,N_7782);
xor U8773 (N_8773,N_7371,N_7068);
nand U8774 (N_8774,N_7453,N_7260);
or U8775 (N_8775,N_6381,N_6745);
nor U8776 (N_8776,N_7803,N_7713);
xnor U8777 (N_8777,N_7875,N_7553);
or U8778 (N_8778,N_7131,N_7196);
or U8779 (N_8779,N_6889,N_7691);
nand U8780 (N_8780,N_6071,N_6716);
and U8781 (N_8781,N_7733,N_7522);
and U8782 (N_8782,N_7138,N_6687);
nor U8783 (N_8783,N_6707,N_6057);
nor U8784 (N_8784,N_6721,N_7307);
nand U8785 (N_8785,N_6177,N_6163);
and U8786 (N_8786,N_7744,N_6991);
or U8787 (N_8787,N_6893,N_6605);
nor U8788 (N_8788,N_7326,N_6812);
nand U8789 (N_8789,N_7093,N_6403);
nor U8790 (N_8790,N_6128,N_6325);
or U8791 (N_8791,N_7279,N_7063);
nand U8792 (N_8792,N_7767,N_7395);
nand U8793 (N_8793,N_7929,N_6518);
and U8794 (N_8794,N_6788,N_7655);
and U8795 (N_8795,N_6316,N_7059);
nand U8796 (N_8796,N_7524,N_6688);
or U8797 (N_8797,N_7035,N_6330);
and U8798 (N_8798,N_6056,N_6482);
or U8799 (N_8799,N_6599,N_6141);
or U8800 (N_8800,N_7600,N_6087);
and U8801 (N_8801,N_6293,N_6424);
nor U8802 (N_8802,N_6847,N_6438);
and U8803 (N_8803,N_7126,N_6420);
or U8804 (N_8804,N_6627,N_6431);
xnor U8805 (N_8805,N_7051,N_7110);
and U8806 (N_8806,N_7968,N_6208);
or U8807 (N_8807,N_6358,N_6409);
nand U8808 (N_8808,N_7628,N_7050);
and U8809 (N_8809,N_6618,N_6831);
nand U8810 (N_8810,N_6499,N_6940);
nand U8811 (N_8811,N_6981,N_7633);
or U8812 (N_8812,N_6905,N_6568);
nand U8813 (N_8813,N_6649,N_6444);
nor U8814 (N_8814,N_7566,N_7770);
nand U8815 (N_8815,N_7506,N_6306);
and U8816 (N_8816,N_7523,N_6086);
nor U8817 (N_8817,N_6701,N_7674);
or U8818 (N_8818,N_6867,N_7340);
or U8819 (N_8819,N_6640,N_7856);
and U8820 (N_8820,N_6769,N_6234);
nand U8821 (N_8821,N_7923,N_6050);
and U8822 (N_8822,N_7398,N_6301);
or U8823 (N_8823,N_7786,N_7243);
or U8824 (N_8824,N_7047,N_7423);
nor U8825 (N_8825,N_7583,N_6924);
or U8826 (N_8826,N_7882,N_7997);
xnor U8827 (N_8827,N_7613,N_7802);
xnor U8828 (N_8828,N_7171,N_7541);
xor U8829 (N_8829,N_6017,N_7761);
nand U8830 (N_8830,N_6193,N_6328);
or U8831 (N_8831,N_6659,N_7403);
and U8832 (N_8832,N_6045,N_6587);
xnor U8833 (N_8833,N_6792,N_7871);
nand U8834 (N_8834,N_6892,N_7826);
nand U8835 (N_8835,N_7868,N_6678);
or U8836 (N_8836,N_7368,N_6712);
nand U8837 (N_8837,N_7550,N_6389);
nor U8838 (N_8838,N_7507,N_6112);
or U8839 (N_8839,N_7317,N_7950);
or U8840 (N_8840,N_7295,N_7757);
or U8841 (N_8841,N_7728,N_7181);
and U8842 (N_8842,N_7659,N_7906);
or U8843 (N_8843,N_7443,N_7323);
nand U8844 (N_8844,N_7262,N_7364);
or U8845 (N_8845,N_6246,N_7623);
and U8846 (N_8846,N_6059,N_6922);
nand U8847 (N_8847,N_6192,N_7031);
xor U8848 (N_8848,N_7354,N_6765);
nand U8849 (N_8849,N_6168,N_6129);
nor U8850 (N_8850,N_6920,N_7879);
and U8851 (N_8851,N_7809,N_7116);
nand U8852 (N_8852,N_6202,N_6238);
nor U8853 (N_8853,N_6786,N_7504);
xnor U8854 (N_8854,N_7460,N_6709);
nand U8855 (N_8855,N_6231,N_6160);
nor U8856 (N_8856,N_7620,N_7637);
nand U8857 (N_8857,N_6762,N_6275);
nor U8858 (N_8858,N_7369,N_7086);
or U8859 (N_8859,N_7973,N_7100);
or U8860 (N_8860,N_6874,N_6399);
nand U8861 (N_8861,N_7854,N_6704);
nor U8862 (N_8862,N_6562,N_7563);
and U8863 (N_8863,N_7737,N_6453);
nand U8864 (N_8864,N_6200,N_6213);
xnor U8865 (N_8865,N_7514,N_7281);
or U8866 (N_8866,N_6318,N_6814);
or U8867 (N_8867,N_7755,N_7582);
nand U8868 (N_8868,N_6854,N_7362);
and U8869 (N_8869,N_7753,N_6487);
nor U8870 (N_8870,N_7763,N_6031);
nor U8871 (N_8871,N_6626,N_7614);
xor U8872 (N_8872,N_6825,N_6600);
nand U8873 (N_8873,N_7248,N_7529);
xnor U8874 (N_8874,N_6746,N_7076);
nor U8875 (N_8875,N_6298,N_6515);
nand U8876 (N_8876,N_6979,N_7045);
or U8877 (N_8877,N_7810,N_7182);
nand U8878 (N_8878,N_7348,N_7607);
nor U8879 (N_8879,N_6677,N_7261);
and U8880 (N_8880,N_7103,N_7201);
nand U8881 (N_8881,N_7715,N_6126);
or U8882 (N_8882,N_7612,N_6123);
nand U8883 (N_8883,N_7382,N_6074);
xnor U8884 (N_8884,N_6522,N_7344);
or U8885 (N_8885,N_7320,N_6353);
and U8886 (N_8886,N_6934,N_7662);
and U8887 (N_8887,N_7793,N_6849);
or U8888 (N_8888,N_6988,N_7195);
and U8889 (N_8889,N_7675,N_6331);
nand U8890 (N_8890,N_6714,N_6785);
and U8891 (N_8891,N_6377,N_7363);
and U8892 (N_8892,N_7357,N_7892);
nor U8893 (N_8893,N_7984,N_7503);
and U8894 (N_8894,N_6560,N_6952);
and U8895 (N_8895,N_7219,N_6902);
or U8896 (N_8896,N_6494,N_6931);
nor U8897 (N_8897,N_6819,N_6995);
and U8898 (N_8898,N_7242,N_6615);
nand U8899 (N_8899,N_6512,N_6303);
xnor U8900 (N_8900,N_6824,N_7491);
nor U8901 (N_8901,N_6468,N_7022);
and U8902 (N_8902,N_7485,N_7921);
nor U8903 (N_8903,N_6547,N_6959);
nor U8904 (N_8904,N_7074,N_6682);
xnor U8905 (N_8905,N_6756,N_6526);
or U8906 (N_8906,N_6588,N_6532);
or U8907 (N_8907,N_7429,N_6851);
nand U8908 (N_8908,N_6862,N_6317);
or U8909 (N_8909,N_6510,N_7355);
nand U8910 (N_8910,N_6161,N_7948);
nor U8911 (N_8911,N_6398,N_7584);
and U8912 (N_8912,N_6451,N_6937);
or U8913 (N_8913,N_7732,N_6324);
or U8914 (N_8914,N_6430,N_6506);
or U8915 (N_8915,N_6808,N_6879);
nand U8916 (N_8916,N_7462,N_6033);
nor U8917 (N_8917,N_7015,N_6255);
xor U8918 (N_8918,N_7268,N_6670);
xnor U8919 (N_8919,N_6405,N_6571);
and U8920 (N_8920,N_6320,N_6777);
nor U8921 (N_8921,N_6860,N_7549);
nor U8922 (N_8922,N_6158,N_6689);
nand U8923 (N_8923,N_7127,N_6658);
nor U8924 (N_8924,N_7207,N_7095);
nor U8925 (N_8925,N_6110,N_6067);
or U8926 (N_8926,N_6329,N_7444);
nor U8927 (N_8927,N_7518,N_6155);
xor U8928 (N_8928,N_6946,N_7700);
nor U8929 (N_8929,N_6654,N_6333);
and U8930 (N_8930,N_7621,N_7365);
and U8931 (N_8931,N_6018,N_6675);
or U8932 (N_8932,N_7825,N_6845);
nand U8933 (N_8933,N_6509,N_7319);
or U8934 (N_8934,N_7502,N_6590);
or U8935 (N_8935,N_7338,N_7099);
nor U8936 (N_8936,N_7133,N_7564);
and U8937 (N_8937,N_7989,N_6579);
xor U8938 (N_8938,N_6573,N_6966);
or U8939 (N_8939,N_7819,N_7161);
nor U8940 (N_8940,N_6037,N_6941);
and U8941 (N_8941,N_6264,N_7283);
xnor U8942 (N_8942,N_7516,N_7631);
and U8943 (N_8943,N_6781,N_7101);
and U8944 (N_8944,N_6008,N_6080);
and U8945 (N_8945,N_6576,N_6530);
nand U8946 (N_8946,N_6350,N_7752);
and U8947 (N_8947,N_6672,N_6070);
xnor U8948 (N_8948,N_7254,N_7840);
nor U8949 (N_8949,N_7998,N_7707);
and U8950 (N_8950,N_6703,N_7458);
and U8951 (N_8951,N_7706,N_7688);
and U8952 (N_8952,N_7560,N_7119);
and U8953 (N_8953,N_7206,N_7064);
nor U8954 (N_8954,N_7946,N_6890);
or U8955 (N_8955,N_6517,N_6992);
or U8956 (N_8956,N_7407,N_7002);
nor U8957 (N_8957,N_7082,N_6989);
and U8958 (N_8958,N_6648,N_6836);
and U8959 (N_8959,N_6741,N_6476);
nand U8960 (N_8960,N_6710,N_7914);
or U8961 (N_8961,N_7581,N_6816);
or U8962 (N_8962,N_6496,N_6841);
and U8963 (N_8963,N_7651,N_6719);
and U8964 (N_8964,N_7513,N_6180);
nor U8965 (N_8965,N_6338,N_6456);
xor U8966 (N_8966,N_6962,N_7586);
or U8967 (N_8967,N_6421,N_7185);
or U8968 (N_8968,N_6612,N_6766);
nor U8969 (N_8969,N_7393,N_6787);
nor U8970 (N_8970,N_7147,N_6203);
nand U8971 (N_8971,N_6207,N_6915);
nor U8972 (N_8972,N_6447,N_6253);
nor U8973 (N_8973,N_7709,N_6038);
nor U8974 (N_8974,N_6827,N_6724);
nor U8975 (N_8975,N_6169,N_6585);
and U8976 (N_8976,N_7801,N_6852);
nor U8977 (N_8977,N_7287,N_7017);
or U8978 (N_8978,N_7469,N_7615);
nand U8979 (N_8979,N_6005,N_7472);
xnor U8980 (N_8980,N_7297,N_7321);
nand U8981 (N_8981,N_6641,N_7410);
nand U8982 (N_8982,N_7285,N_6489);
nor U8983 (N_8983,N_6702,N_7712);
and U8984 (N_8984,N_6269,N_6669);
nor U8985 (N_8985,N_7557,N_6911);
nor U8986 (N_8986,N_7861,N_7060);
and U8987 (N_8987,N_7558,N_6896);
and U8988 (N_8988,N_7609,N_6311);
xnor U8989 (N_8989,N_7332,N_6900);
nand U8990 (N_8990,N_6556,N_6690);
nand U8991 (N_8991,N_6411,N_7866);
nand U8992 (N_8992,N_6950,N_6876);
and U8993 (N_8993,N_6131,N_7955);
or U8994 (N_8994,N_7222,N_7654);
and U8995 (N_8995,N_6240,N_7072);
or U8996 (N_8996,N_7425,N_7511);
or U8997 (N_8997,N_7373,N_7910);
and U8998 (N_8998,N_7236,N_6443);
and U8999 (N_8999,N_6026,N_7742);
nor U9000 (N_9000,N_6841,N_6405);
nor U9001 (N_9001,N_7705,N_6655);
and U9002 (N_9002,N_7219,N_7388);
nand U9003 (N_9003,N_6971,N_7034);
nand U9004 (N_9004,N_6925,N_6263);
xnor U9005 (N_9005,N_7395,N_7448);
nor U9006 (N_9006,N_7808,N_6409);
nor U9007 (N_9007,N_6737,N_7454);
or U9008 (N_9008,N_7171,N_6087);
nand U9009 (N_9009,N_6693,N_7491);
nor U9010 (N_9010,N_6422,N_7420);
nand U9011 (N_9011,N_6817,N_6438);
nand U9012 (N_9012,N_6630,N_6351);
nand U9013 (N_9013,N_6007,N_6067);
and U9014 (N_9014,N_7199,N_7457);
and U9015 (N_9015,N_6842,N_6005);
nand U9016 (N_9016,N_7400,N_6399);
nand U9017 (N_9017,N_6180,N_7617);
nand U9018 (N_9018,N_7792,N_7128);
nand U9019 (N_9019,N_6922,N_7725);
and U9020 (N_9020,N_6922,N_6420);
nor U9021 (N_9021,N_7101,N_6329);
nor U9022 (N_9022,N_7177,N_6519);
nand U9023 (N_9023,N_7142,N_6846);
or U9024 (N_9024,N_6946,N_6417);
xor U9025 (N_9025,N_6479,N_7646);
nand U9026 (N_9026,N_7842,N_7640);
and U9027 (N_9027,N_7797,N_7260);
and U9028 (N_9028,N_6672,N_6605);
nand U9029 (N_9029,N_6572,N_7313);
and U9030 (N_9030,N_6484,N_7280);
nor U9031 (N_9031,N_6627,N_6379);
or U9032 (N_9032,N_6543,N_7110);
or U9033 (N_9033,N_7836,N_7061);
and U9034 (N_9034,N_7554,N_7789);
xor U9035 (N_9035,N_7173,N_6382);
or U9036 (N_9036,N_6927,N_7363);
and U9037 (N_9037,N_6132,N_7021);
or U9038 (N_9038,N_6197,N_7689);
nand U9039 (N_9039,N_7466,N_6417);
and U9040 (N_9040,N_6985,N_7205);
xnor U9041 (N_9041,N_6812,N_7933);
or U9042 (N_9042,N_7369,N_7991);
nand U9043 (N_9043,N_7980,N_6367);
or U9044 (N_9044,N_6408,N_7671);
or U9045 (N_9045,N_6464,N_7117);
xnor U9046 (N_9046,N_7919,N_7345);
and U9047 (N_9047,N_6429,N_7974);
nor U9048 (N_9048,N_7639,N_7544);
and U9049 (N_9049,N_6539,N_6748);
nand U9050 (N_9050,N_7005,N_6389);
nand U9051 (N_9051,N_6896,N_6003);
nor U9052 (N_9052,N_6052,N_6464);
xnor U9053 (N_9053,N_7059,N_6971);
nor U9054 (N_9054,N_7666,N_7890);
nor U9055 (N_9055,N_6015,N_6496);
xnor U9056 (N_9056,N_7972,N_7023);
nand U9057 (N_9057,N_6933,N_7643);
nand U9058 (N_9058,N_7232,N_6299);
or U9059 (N_9059,N_6088,N_6689);
or U9060 (N_9060,N_7195,N_6781);
xnor U9061 (N_9061,N_7836,N_7148);
nand U9062 (N_9062,N_7273,N_7301);
or U9063 (N_9063,N_7968,N_6837);
and U9064 (N_9064,N_7342,N_7232);
or U9065 (N_9065,N_6939,N_7083);
nand U9066 (N_9066,N_6032,N_6811);
and U9067 (N_9067,N_7323,N_6064);
and U9068 (N_9068,N_6616,N_7504);
or U9069 (N_9069,N_6344,N_7402);
and U9070 (N_9070,N_7849,N_7669);
and U9071 (N_9071,N_6807,N_7124);
nor U9072 (N_9072,N_7441,N_6908);
xnor U9073 (N_9073,N_6172,N_6366);
nand U9074 (N_9074,N_7004,N_7066);
nand U9075 (N_9075,N_6583,N_6208);
nand U9076 (N_9076,N_7673,N_6926);
nor U9077 (N_9077,N_7441,N_6862);
and U9078 (N_9078,N_7129,N_6673);
and U9079 (N_9079,N_6300,N_7694);
nor U9080 (N_9080,N_6854,N_6939);
or U9081 (N_9081,N_6035,N_6586);
and U9082 (N_9082,N_6943,N_7426);
and U9083 (N_9083,N_6585,N_6871);
xor U9084 (N_9084,N_7790,N_7891);
or U9085 (N_9085,N_7659,N_6989);
nor U9086 (N_9086,N_6774,N_7840);
nand U9087 (N_9087,N_7839,N_7133);
nor U9088 (N_9088,N_6344,N_7781);
nand U9089 (N_9089,N_7828,N_7837);
or U9090 (N_9090,N_6416,N_6715);
nor U9091 (N_9091,N_7607,N_6345);
and U9092 (N_9092,N_7406,N_7370);
or U9093 (N_9093,N_7654,N_6068);
or U9094 (N_9094,N_6639,N_6164);
and U9095 (N_9095,N_6982,N_7330);
nor U9096 (N_9096,N_6882,N_6369);
nand U9097 (N_9097,N_7469,N_7172);
nand U9098 (N_9098,N_6694,N_6740);
nor U9099 (N_9099,N_6368,N_7705);
nand U9100 (N_9100,N_7992,N_7395);
and U9101 (N_9101,N_6878,N_6693);
and U9102 (N_9102,N_7049,N_6274);
nand U9103 (N_9103,N_6063,N_7569);
or U9104 (N_9104,N_6295,N_6336);
nor U9105 (N_9105,N_7132,N_7220);
or U9106 (N_9106,N_6136,N_7763);
nor U9107 (N_9107,N_6631,N_7719);
nand U9108 (N_9108,N_6190,N_7044);
nor U9109 (N_9109,N_7539,N_7051);
nand U9110 (N_9110,N_6202,N_6827);
nor U9111 (N_9111,N_6471,N_7731);
nor U9112 (N_9112,N_7774,N_6873);
nand U9113 (N_9113,N_7468,N_7604);
and U9114 (N_9114,N_7395,N_7898);
nor U9115 (N_9115,N_7604,N_6501);
nor U9116 (N_9116,N_6727,N_7569);
nor U9117 (N_9117,N_7230,N_6857);
and U9118 (N_9118,N_6884,N_6513);
nor U9119 (N_9119,N_7879,N_6692);
and U9120 (N_9120,N_6623,N_7226);
xnor U9121 (N_9121,N_7959,N_6729);
xnor U9122 (N_9122,N_7407,N_6231);
xnor U9123 (N_9123,N_6782,N_7618);
nand U9124 (N_9124,N_6465,N_7769);
and U9125 (N_9125,N_7479,N_7210);
nand U9126 (N_9126,N_7076,N_6661);
or U9127 (N_9127,N_6022,N_6829);
and U9128 (N_9128,N_7717,N_6883);
or U9129 (N_9129,N_7910,N_7770);
xor U9130 (N_9130,N_7881,N_7809);
nor U9131 (N_9131,N_7460,N_6726);
nor U9132 (N_9132,N_6808,N_6088);
nand U9133 (N_9133,N_6593,N_7608);
or U9134 (N_9134,N_6497,N_7414);
nor U9135 (N_9135,N_6629,N_6231);
nand U9136 (N_9136,N_6803,N_6886);
or U9137 (N_9137,N_7365,N_7818);
nor U9138 (N_9138,N_6277,N_7624);
nor U9139 (N_9139,N_6308,N_6088);
nor U9140 (N_9140,N_6042,N_7867);
xor U9141 (N_9141,N_7416,N_6757);
or U9142 (N_9142,N_6771,N_7889);
and U9143 (N_9143,N_6938,N_7730);
or U9144 (N_9144,N_7766,N_6977);
and U9145 (N_9145,N_6750,N_6090);
and U9146 (N_9146,N_7684,N_7353);
nand U9147 (N_9147,N_6686,N_6705);
nor U9148 (N_9148,N_6811,N_7610);
or U9149 (N_9149,N_6483,N_6362);
nor U9150 (N_9150,N_7969,N_6645);
or U9151 (N_9151,N_7149,N_6903);
or U9152 (N_9152,N_6579,N_6025);
and U9153 (N_9153,N_6783,N_7325);
nand U9154 (N_9154,N_7373,N_7197);
or U9155 (N_9155,N_6607,N_6416);
nand U9156 (N_9156,N_6944,N_7539);
xor U9157 (N_9157,N_6100,N_7545);
and U9158 (N_9158,N_6017,N_7437);
and U9159 (N_9159,N_7881,N_7584);
xor U9160 (N_9160,N_6447,N_7170);
nor U9161 (N_9161,N_7194,N_7099);
nand U9162 (N_9162,N_6012,N_6320);
and U9163 (N_9163,N_7557,N_7777);
and U9164 (N_9164,N_7042,N_7420);
and U9165 (N_9165,N_7564,N_6573);
nand U9166 (N_9166,N_7383,N_7060);
nor U9167 (N_9167,N_7707,N_6747);
nor U9168 (N_9168,N_7041,N_7634);
xor U9169 (N_9169,N_7535,N_6937);
xor U9170 (N_9170,N_6032,N_6810);
nor U9171 (N_9171,N_7685,N_6666);
or U9172 (N_9172,N_6945,N_7759);
or U9173 (N_9173,N_7151,N_7145);
nand U9174 (N_9174,N_6510,N_6300);
nand U9175 (N_9175,N_7997,N_7473);
nor U9176 (N_9176,N_6677,N_6875);
nand U9177 (N_9177,N_6229,N_7675);
nand U9178 (N_9178,N_6669,N_7185);
or U9179 (N_9179,N_6748,N_7524);
and U9180 (N_9180,N_7008,N_6698);
nor U9181 (N_9181,N_7361,N_6953);
nand U9182 (N_9182,N_6617,N_6586);
nor U9183 (N_9183,N_6470,N_6664);
nand U9184 (N_9184,N_7111,N_7427);
xor U9185 (N_9185,N_7096,N_7964);
or U9186 (N_9186,N_7000,N_7044);
or U9187 (N_9187,N_6488,N_7716);
xnor U9188 (N_9188,N_6093,N_6418);
or U9189 (N_9189,N_6845,N_6187);
or U9190 (N_9190,N_6486,N_6784);
xor U9191 (N_9191,N_7845,N_7121);
nand U9192 (N_9192,N_6496,N_7627);
or U9193 (N_9193,N_6613,N_7656);
and U9194 (N_9194,N_7541,N_6286);
nand U9195 (N_9195,N_7064,N_7114);
nand U9196 (N_9196,N_6817,N_6687);
nand U9197 (N_9197,N_6320,N_7505);
and U9198 (N_9198,N_7150,N_7607);
and U9199 (N_9199,N_7217,N_6183);
nor U9200 (N_9200,N_7430,N_6395);
nor U9201 (N_9201,N_7390,N_7018);
nor U9202 (N_9202,N_6647,N_6136);
and U9203 (N_9203,N_6110,N_6475);
nor U9204 (N_9204,N_6951,N_6741);
nand U9205 (N_9205,N_6778,N_7726);
nor U9206 (N_9206,N_7744,N_6887);
and U9207 (N_9207,N_6544,N_7152);
xor U9208 (N_9208,N_6490,N_6276);
xnor U9209 (N_9209,N_7836,N_7598);
nor U9210 (N_9210,N_7356,N_7800);
nand U9211 (N_9211,N_7230,N_7566);
or U9212 (N_9212,N_7485,N_6606);
xor U9213 (N_9213,N_6658,N_7903);
or U9214 (N_9214,N_6257,N_6333);
nand U9215 (N_9215,N_6793,N_7980);
and U9216 (N_9216,N_6065,N_7297);
nand U9217 (N_9217,N_6239,N_6335);
nor U9218 (N_9218,N_6518,N_7072);
nor U9219 (N_9219,N_7840,N_7512);
or U9220 (N_9220,N_7393,N_7038);
nor U9221 (N_9221,N_7360,N_7624);
nand U9222 (N_9222,N_7912,N_6369);
nand U9223 (N_9223,N_7468,N_7620);
nor U9224 (N_9224,N_6303,N_7284);
nor U9225 (N_9225,N_6040,N_6810);
nand U9226 (N_9226,N_7811,N_6082);
nor U9227 (N_9227,N_7084,N_7027);
or U9228 (N_9228,N_7682,N_6846);
or U9229 (N_9229,N_7033,N_6479);
nand U9230 (N_9230,N_7231,N_7728);
and U9231 (N_9231,N_7213,N_7619);
nor U9232 (N_9232,N_6216,N_7114);
nor U9233 (N_9233,N_6276,N_7864);
nand U9234 (N_9234,N_7252,N_6359);
nand U9235 (N_9235,N_7197,N_7771);
and U9236 (N_9236,N_7544,N_7229);
or U9237 (N_9237,N_6630,N_6869);
and U9238 (N_9238,N_6795,N_7429);
nand U9239 (N_9239,N_6676,N_7248);
or U9240 (N_9240,N_7677,N_6158);
nor U9241 (N_9241,N_6883,N_6466);
and U9242 (N_9242,N_6730,N_6107);
and U9243 (N_9243,N_7176,N_6295);
nor U9244 (N_9244,N_7209,N_6923);
and U9245 (N_9245,N_6697,N_6006);
nor U9246 (N_9246,N_6829,N_6767);
nand U9247 (N_9247,N_6111,N_7019);
nor U9248 (N_9248,N_7328,N_7815);
and U9249 (N_9249,N_7626,N_7165);
nand U9250 (N_9250,N_7247,N_7472);
or U9251 (N_9251,N_6052,N_6910);
nand U9252 (N_9252,N_6903,N_6470);
nand U9253 (N_9253,N_6567,N_7541);
xnor U9254 (N_9254,N_6221,N_7093);
nand U9255 (N_9255,N_6319,N_6683);
or U9256 (N_9256,N_6561,N_6921);
and U9257 (N_9257,N_6742,N_7507);
nor U9258 (N_9258,N_6498,N_6183);
nand U9259 (N_9259,N_6543,N_7901);
or U9260 (N_9260,N_7980,N_7223);
and U9261 (N_9261,N_6681,N_7409);
and U9262 (N_9262,N_6544,N_7267);
nor U9263 (N_9263,N_7590,N_7338);
nor U9264 (N_9264,N_7696,N_6704);
nand U9265 (N_9265,N_7344,N_6279);
or U9266 (N_9266,N_7879,N_6653);
nor U9267 (N_9267,N_7173,N_6680);
nand U9268 (N_9268,N_6484,N_7681);
nand U9269 (N_9269,N_6695,N_6385);
and U9270 (N_9270,N_6739,N_7065);
and U9271 (N_9271,N_6319,N_7618);
nor U9272 (N_9272,N_7936,N_6683);
nor U9273 (N_9273,N_6936,N_6013);
nand U9274 (N_9274,N_7254,N_7782);
nand U9275 (N_9275,N_6134,N_6892);
and U9276 (N_9276,N_6049,N_7145);
and U9277 (N_9277,N_7047,N_6332);
or U9278 (N_9278,N_7654,N_6810);
nand U9279 (N_9279,N_6331,N_7120);
and U9280 (N_9280,N_6857,N_6030);
or U9281 (N_9281,N_6995,N_6676);
or U9282 (N_9282,N_7477,N_6132);
and U9283 (N_9283,N_7414,N_6399);
nor U9284 (N_9284,N_6918,N_7018);
and U9285 (N_9285,N_6809,N_6628);
or U9286 (N_9286,N_6933,N_7822);
xor U9287 (N_9287,N_6862,N_7563);
xnor U9288 (N_9288,N_6102,N_6687);
or U9289 (N_9289,N_6102,N_7589);
nor U9290 (N_9290,N_6036,N_7643);
and U9291 (N_9291,N_6201,N_6084);
nor U9292 (N_9292,N_7504,N_6797);
and U9293 (N_9293,N_7547,N_7427);
and U9294 (N_9294,N_6381,N_6860);
xor U9295 (N_9295,N_6134,N_6975);
and U9296 (N_9296,N_7959,N_6733);
or U9297 (N_9297,N_6715,N_7097);
nand U9298 (N_9298,N_7824,N_6156);
nor U9299 (N_9299,N_7260,N_6381);
or U9300 (N_9300,N_7085,N_7224);
nor U9301 (N_9301,N_6818,N_6120);
or U9302 (N_9302,N_7440,N_6359);
nor U9303 (N_9303,N_7122,N_7397);
nand U9304 (N_9304,N_6881,N_7580);
nor U9305 (N_9305,N_6548,N_6971);
and U9306 (N_9306,N_7740,N_7268);
or U9307 (N_9307,N_6971,N_6145);
nand U9308 (N_9308,N_7046,N_6058);
nand U9309 (N_9309,N_7547,N_7166);
nand U9310 (N_9310,N_6263,N_7900);
nor U9311 (N_9311,N_7454,N_6992);
or U9312 (N_9312,N_7705,N_7644);
nor U9313 (N_9313,N_6891,N_6141);
nor U9314 (N_9314,N_7232,N_6242);
nand U9315 (N_9315,N_7819,N_6934);
and U9316 (N_9316,N_7749,N_7976);
and U9317 (N_9317,N_6243,N_6031);
and U9318 (N_9318,N_7456,N_6145);
xor U9319 (N_9319,N_7364,N_6045);
nand U9320 (N_9320,N_7268,N_7686);
or U9321 (N_9321,N_6223,N_7041);
nand U9322 (N_9322,N_6500,N_7884);
nor U9323 (N_9323,N_6509,N_6008);
or U9324 (N_9324,N_7639,N_7981);
nor U9325 (N_9325,N_6517,N_7702);
nand U9326 (N_9326,N_6228,N_7075);
nand U9327 (N_9327,N_6914,N_6828);
xnor U9328 (N_9328,N_6892,N_7808);
or U9329 (N_9329,N_7693,N_7329);
or U9330 (N_9330,N_6536,N_6324);
nor U9331 (N_9331,N_6188,N_6330);
nand U9332 (N_9332,N_6826,N_6060);
nand U9333 (N_9333,N_7929,N_7585);
xor U9334 (N_9334,N_7071,N_6662);
nor U9335 (N_9335,N_7467,N_6078);
nor U9336 (N_9336,N_7232,N_7786);
nand U9337 (N_9337,N_6162,N_6509);
or U9338 (N_9338,N_6510,N_6474);
or U9339 (N_9339,N_7228,N_7121);
and U9340 (N_9340,N_7045,N_7781);
or U9341 (N_9341,N_6122,N_7547);
nor U9342 (N_9342,N_6983,N_6701);
nor U9343 (N_9343,N_6750,N_6319);
nand U9344 (N_9344,N_7081,N_7112);
xor U9345 (N_9345,N_6800,N_7823);
or U9346 (N_9346,N_6865,N_7452);
nor U9347 (N_9347,N_6585,N_6035);
nor U9348 (N_9348,N_7991,N_7188);
or U9349 (N_9349,N_7876,N_7255);
nor U9350 (N_9350,N_7122,N_7059);
nand U9351 (N_9351,N_7902,N_7046);
nand U9352 (N_9352,N_7517,N_7839);
and U9353 (N_9353,N_7424,N_6616);
and U9354 (N_9354,N_7523,N_6873);
xor U9355 (N_9355,N_7231,N_7919);
nor U9356 (N_9356,N_7291,N_7273);
nor U9357 (N_9357,N_6679,N_6300);
or U9358 (N_9358,N_6077,N_7033);
nand U9359 (N_9359,N_6725,N_7999);
nor U9360 (N_9360,N_7338,N_6279);
or U9361 (N_9361,N_6055,N_6276);
or U9362 (N_9362,N_6053,N_7193);
nand U9363 (N_9363,N_6746,N_6584);
nand U9364 (N_9364,N_7500,N_6924);
nand U9365 (N_9365,N_7479,N_6040);
or U9366 (N_9366,N_7055,N_6732);
xor U9367 (N_9367,N_6262,N_7336);
nor U9368 (N_9368,N_6251,N_7147);
or U9369 (N_9369,N_6036,N_6423);
nand U9370 (N_9370,N_6018,N_6425);
and U9371 (N_9371,N_6405,N_7819);
nor U9372 (N_9372,N_7299,N_7729);
or U9373 (N_9373,N_6972,N_6768);
or U9374 (N_9374,N_6479,N_7809);
nor U9375 (N_9375,N_7579,N_6230);
or U9376 (N_9376,N_6349,N_7345);
nand U9377 (N_9377,N_6727,N_7503);
or U9378 (N_9378,N_7779,N_7289);
and U9379 (N_9379,N_7593,N_7709);
xor U9380 (N_9380,N_7871,N_6496);
and U9381 (N_9381,N_7957,N_6624);
or U9382 (N_9382,N_6165,N_6693);
nor U9383 (N_9383,N_6807,N_7616);
nor U9384 (N_9384,N_6619,N_7151);
nor U9385 (N_9385,N_6403,N_6563);
xnor U9386 (N_9386,N_7527,N_7337);
and U9387 (N_9387,N_7487,N_7322);
and U9388 (N_9388,N_6486,N_6177);
nand U9389 (N_9389,N_6360,N_7989);
nor U9390 (N_9390,N_7244,N_7825);
and U9391 (N_9391,N_6218,N_7483);
nor U9392 (N_9392,N_6640,N_7838);
nand U9393 (N_9393,N_7384,N_7359);
nand U9394 (N_9394,N_7053,N_6104);
nor U9395 (N_9395,N_7717,N_6698);
nand U9396 (N_9396,N_7444,N_7828);
nor U9397 (N_9397,N_6750,N_7325);
nand U9398 (N_9398,N_7402,N_6780);
nor U9399 (N_9399,N_7101,N_6661);
or U9400 (N_9400,N_7838,N_7468);
and U9401 (N_9401,N_6889,N_6816);
xor U9402 (N_9402,N_7555,N_7272);
and U9403 (N_9403,N_7693,N_7834);
and U9404 (N_9404,N_7714,N_6079);
or U9405 (N_9405,N_7119,N_6411);
or U9406 (N_9406,N_6850,N_7350);
and U9407 (N_9407,N_7761,N_6417);
nor U9408 (N_9408,N_6550,N_7861);
nor U9409 (N_9409,N_6877,N_6816);
nand U9410 (N_9410,N_6401,N_7374);
and U9411 (N_9411,N_6280,N_7013);
nor U9412 (N_9412,N_6493,N_6962);
and U9413 (N_9413,N_7320,N_7348);
nor U9414 (N_9414,N_7791,N_7020);
xnor U9415 (N_9415,N_6751,N_7872);
and U9416 (N_9416,N_7485,N_6727);
or U9417 (N_9417,N_6956,N_7937);
and U9418 (N_9418,N_7345,N_7611);
or U9419 (N_9419,N_6656,N_7924);
or U9420 (N_9420,N_7269,N_6835);
xnor U9421 (N_9421,N_6244,N_7878);
and U9422 (N_9422,N_7542,N_6128);
nor U9423 (N_9423,N_6014,N_6217);
or U9424 (N_9424,N_6094,N_7564);
nand U9425 (N_9425,N_6491,N_7491);
nand U9426 (N_9426,N_7549,N_7554);
nand U9427 (N_9427,N_7585,N_6991);
nor U9428 (N_9428,N_6083,N_6512);
and U9429 (N_9429,N_7519,N_6225);
and U9430 (N_9430,N_7482,N_7643);
nand U9431 (N_9431,N_7375,N_6745);
nor U9432 (N_9432,N_7573,N_7875);
nor U9433 (N_9433,N_7915,N_6265);
and U9434 (N_9434,N_7421,N_7678);
nor U9435 (N_9435,N_6800,N_7637);
or U9436 (N_9436,N_6906,N_6230);
nand U9437 (N_9437,N_6418,N_7936);
xnor U9438 (N_9438,N_6138,N_6150);
nand U9439 (N_9439,N_6963,N_7817);
nand U9440 (N_9440,N_6326,N_6997);
nand U9441 (N_9441,N_7895,N_7607);
nand U9442 (N_9442,N_6362,N_7788);
nor U9443 (N_9443,N_6160,N_6659);
and U9444 (N_9444,N_7961,N_7862);
and U9445 (N_9445,N_7806,N_6547);
nor U9446 (N_9446,N_6086,N_7616);
and U9447 (N_9447,N_6321,N_7178);
nand U9448 (N_9448,N_7206,N_7831);
and U9449 (N_9449,N_7976,N_6466);
or U9450 (N_9450,N_6457,N_6247);
xor U9451 (N_9451,N_6971,N_7138);
nor U9452 (N_9452,N_6201,N_6607);
nor U9453 (N_9453,N_7412,N_7338);
nand U9454 (N_9454,N_6286,N_7649);
and U9455 (N_9455,N_6930,N_7067);
nand U9456 (N_9456,N_7634,N_7471);
or U9457 (N_9457,N_6504,N_6953);
or U9458 (N_9458,N_6683,N_6276);
or U9459 (N_9459,N_6301,N_7667);
nand U9460 (N_9460,N_6872,N_7038);
xor U9461 (N_9461,N_7709,N_6549);
or U9462 (N_9462,N_6891,N_6211);
or U9463 (N_9463,N_7487,N_7833);
or U9464 (N_9464,N_7058,N_7017);
xnor U9465 (N_9465,N_7441,N_7177);
nand U9466 (N_9466,N_6125,N_7608);
nor U9467 (N_9467,N_6507,N_7895);
nor U9468 (N_9468,N_7094,N_7307);
xnor U9469 (N_9469,N_7159,N_7584);
nand U9470 (N_9470,N_7300,N_6833);
nor U9471 (N_9471,N_6496,N_6569);
nand U9472 (N_9472,N_7618,N_7334);
nand U9473 (N_9473,N_7956,N_6362);
or U9474 (N_9474,N_7959,N_7497);
nor U9475 (N_9475,N_6600,N_7082);
nand U9476 (N_9476,N_7888,N_7180);
nand U9477 (N_9477,N_6097,N_6537);
nand U9478 (N_9478,N_7109,N_7269);
nor U9479 (N_9479,N_7286,N_7472);
nand U9480 (N_9480,N_7571,N_6975);
and U9481 (N_9481,N_6515,N_6909);
xor U9482 (N_9482,N_6698,N_6838);
or U9483 (N_9483,N_7180,N_7812);
nor U9484 (N_9484,N_7782,N_6679);
and U9485 (N_9485,N_6729,N_7993);
nand U9486 (N_9486,N_6787,N_7259);
or U9487 (N_9487,N_6024,N_7260);
and U9488 (N_9488,N_6304,N_7083);
and U9489 (N_9489,N_7425,N_6467);
nand U9490 (N_9490,N_6751,N_7606);
or U9491 (N_9491,N_6999,N_7130);
xor U9492 (N_9492,N_7596,N_7569);
and U9493 (N_9493,N_6973,N_6535);
nand U9494 (N_9494,N_7504,N_6784);
xnor U9495 (N_9495,N_7633,N_7730);
and U9496 (N_9496,N_7041,N_6986);
nand U9497 (N_9497,N_7379,N_7443);
and U9498 (N_9498,N_7915,N_6929);
or U9499 (N_9499,N_7543,N_6838);
nand U9500 (N_9500,N_6601,N_7845);
nand U9501 (N_9501,N_6172,N_6584);
nor U9502 (N_9502,N_7162,N_7514);
or U9503 (N_9503,N_6091,N_7934);
or U9504 (N_9504,N_6157,N_7254);
nand U9505 (N_9505,N_7709,N_6507);
nand U9506 (N_9506,N_6615,N_6389);
or U9507 (N_9507,N_7374,N_6960);
xor U9508 (N_9508,N_6111,N_7172);
or U9509 (N_9509,N_6884,N_7847);
xnor U9510 (N_9510,N_7363,N_6685);
and U9511 (N_9511,N_6697,N_7654);
nand U9512 (N_9512,N_7010,N_6108);
nand U9513 (N_9513,N_6838,N_6304);
or U9514 (N_9514,N_7844,N_7774);
or U9515 (N_9515,N_7819,N_7441);
or U9516 (N_9516,N_7495,N_7264);
nor U9517 (N_9517,N_7015,N_6666);
or U9518 (N_9518,N_6620,N_6881);
xor U9519 (N_9519,N_6061,N_6869);
nor U9520 (N_9520,N_7878,N_6223);
and U9521 (N_9521,N_7541,N_6143);
or U9522 (N_9522,N_7866,N_7360);
nand U9523 (N_9523,N_6766,N_7996);
nand U9524 (N_9524,N_7023,N_6948);
nand U9525 (N_9525,N_6559,N_7494);
nor U9526 (N_9526,N_7891,N_7230);
and U9527 (N_9527,N_7497,N_7019);
nand U9528 (N_9528,N_6907,N_6662);
and U9529 (N_9529,N_6240,N_7419);
and U9530 (N_9530,N_6595,N_7490);
xnor U9531 (N_9531,N_7111,N_7800);
and U9532 (N_9532,N_6057,N_7247);
and U9533 (N_9533,N_7703,N_6704);
and U9534 (N_9534,N_6086,N_6219);
xnor U9535 (N_9535,N_7923,N_7757);
nor U9536 (N_9536,N_7807,N_7888);
and U9537 (N_9537,N_7729,N_6198);
xnor U9538 (N_9538,N_7715,N_6263);
or U9539 (N_9539,N_7331,N_6473);
nor U9540 (N_9540,N_6479,N_6204);
xor U9541 (N_9541,N_6062,N_7269);
or U9542 (N_9542,N_6806,N_6734);
and U9543 (N_9543,N_7638,N_7364);
nand U9544 (N_9544,N_6200,N_6430);
nor U9545 (N_9545,N_6539,N_7723);
or U9546 (N_9546,N_7700,N_7261);
xor U9547 (N_9547,N_7143,N_6638);
nor U9548 (N_9548,N_6127,N_6457);
and U9549 (N_9549,N_7566,N_7140);
and U9550 (N_9550,N_7901,N_6157);
or U9551 (N_9551,N_7584,N_7255);
nor U9552 (N_9552,N_7437,N_6034);
and U9553 (N_9553,N_6639,N_7751);
xor U9554 (N_9554,N_7618,N_7379);
nand U9555 (N_9555,N_7127,N_7739);
nand U9556 (N_9556,N_6696,N_7674);
and U9557 (N_9557,N_7156,N_7647);
and U9558 (N_9558,N_7389,N_7128);
nand U9559 (N_9559,N_6260,N_6871);
and U9560 (N_9560,N_7635,N_6588);
or U9561 (N_9561,N_6380,N_6608);
or U9562 (N_9562,N_7745,N_7483);
and U9563 (N_9563,N_7394,N_6838);
and U9564 (N_9564,N_6121,N_7569);
and U9565 (N_9565,N_6029,N_6983);
xnor U9566 (N_9566,N_7651,N_7985);
or U9567 (N_9567,N_6414,N_7210);
nand U9568 (N_9568,N_7681,N_6299);
nor U9569 (N_9569,N_7417,N_7870);
and U9570 (N_9570,N_6913,N_6647);
nor U9571 (N_9571,N_7563,N_7300);
nand U9572 (N_9572,N_6942,N_6346);
xor U9573 (N_9573,N_6917,N_6092);
or U9574 (N_9574,N_7947,N_7742);
nor U9575 (N_9575,N_7651,N_6901);
or U9576 (N_9576,N_7068,N_7047);
nor U9577 (N_9577,N_7410,N_7527);
nor U9578 (N_9578,N_7624,N_7927);
and U9579 (N_9579,N_6789,N_7518);
nand U9580 (N_9580,N_6362,N_7669);
or U9581 (N_9581,N_7755,N_7168);
nor U9582 (N_9582,N_6249,N_7811);
or U9583 (N_9583,N_7712,N_7083);
xnor U9584 (N_9584,N_6604,N_6145);
xor U9585 (N_9585,N_7484,N_7462);
or U9586 (N_9586,N_7268,N_7786);
nor U9587 (N_9587,N_6200,N_7295);
and U9588 (N_9588,N_7195,N_6436);
nor U9589 (N_9589,N_6604,N_6901);
and U9590 (N_9590,N_6278,N_7782);
or U9591 (N_9591,N_6429,N_6825);
or U9592 (N_9592,N_6310,N_7806);
nand U9593 (N_9593,N_7849,N_6690);
and U9594 (N_9594,N_7019,N_6268);
or U9595 (N_9595,N_7900,N_7247);
nand U9596 (N_9596,N_7725,N_7091);
and U9597 (N_9597,N_7206,N_7656);
or U9598 (N_9598,N_6379,N_6078);
nand U9599 (N_9599,N_7962,N_6136);
xor U9600 (N_9600,N_6841,N_7744);
or U9601 (N_9601,N_6340,N_6555);
and U9602 (N_9602,N_6218,N_6149);
or U9603 (N_9603,N_7925,N_7590);
and U9604 (N_9604,N_7774,N_7306);
xor U9605 (N_9605,N_6323,N_6574);
xnor U9606 (N_9606,N_7847,N_6140);
or U9607 (N_9607,N_7378,N_6018);
nor U9608 (N_9608,N_6368,N_7876);
nand U9609 (N_9609,N_7417,N_7093);
and U9610 (N_9610,N_7240,N_7783);
nand U9611 (N_9611,N_7505,N_6856);
nand U9612 (N_9612,N_6016,N_6259);
or U9613 (N_9613,N_7471,N_7760);
nor U9614 (N_9614,N_7861,N_7192);
and U9615 (N_9615,N_7855,N_7017);
or U9616 (N_9616,N_6334,N_6912);
xor U9617 (N_9617,N_6158,N_7019);
xor U9618 (N_9618,N_7228,N_6360);
nand U9619 (N_9619,N_6286,N_6430);
nand U9620 (N_9620,N_6230,N_7800);
xnor U9621 (N_9621,N_7885,N_7944);
and U9622 (N_9622,N_6050,N_7767);
and U9623 (N_9623,N_7520,N_7747);
and U9624 (N_9624,N_6897,N_7898);
and U9625 (N_9625,N_7538,N_6237);
nor U9626 (N_9626,N_7363,N_6439);
nand U9627 (N_9627,N_7684,N_6149);
or U9628 (N_9628,N_6467,N_7638);
nor U9629 (N_9629,N_6936,N_7511);
and U9630 (N_9630,N_7996,N_7923);
and U9631 (N_9631,N_7508,N_7022);
nand U9632 (N_9632,N_7240,N_6701);
nand U9633 (N_9633,N_7976,N_6275);
nor U9634 (N_9634,N_7206,N_7191);
and U9635 (N_9635,N_6917,N_7772);
nor U9636 (N_9636,N_7474,N_7017);
nand U9637 (N_9637,N_7789,N_6035);
xnor U9638 (N_9638,N_6459,N_7115);
nor U9639 (N_9639,N_6725,N_6338);
nand U9640 (N_9640,N_6706,N_7458);
nor U9641 (N_9641,N_7591,N_7022);
or U9642 (N_9642,N_6829,N_6525);
and U9643 (N_9643,N_6198,N_7852);
or U9644 (N_9644,N_7828,N_7080);
xor U9645 (N_9645,N_7226,N_7522);
nor U9646 (N_9646,N_6808,N_6485);
and U9647 (N_9647,N_7454,N_7209);
xor U9648 (N_9648,N_6012,N_6591);
and U9649 (N_9649,N_6109,N_6094);
or U9650 (N_9650,N_6016,N_7805);
or U9651 (N_9651,N_7993,N_7318);
and U9652 (N_9652,N_7782,N_7371);
nor U9653 (N_9653,N_6913,N_7218);
nand U9654 (N_9654,N_7691,N_7034);
and U9655 (N_9655,N_7612,N_7321);
and U9656 (N_9656,N_7377,N_7869);
nor U9657 (N_9657,N_6686,N_7994);
nand U9658 (N_9658,N_7833,N_6236);
nor U9659 (N_9659,N_7896,N_7167);
or U9660 (N_9660,N_7550,N_6747);
nand U9661 (N_9661,N_6554,N_6013);
nor U9662 (N_9662,N_6457,N_6700);
or U9663 (N_9663,N_6569,N_6902);
nor U9664 (N_9664,N_7475,N_7743);
or U9665 (N_9665,N_7442,N_6416);
or U9666 (N_9666,N_7927,N_7511);
or U9667 (N_9667,N_7981,N_7587);
nand U9668 (N_9668,N_7465,N_6937);
and U9669 (N_9669,N_7782,N_6099);
nor U9670 (N_9670,N_7222,N_7215);
nor U9671 (N_9671,N_7224,N_6633);
or U9672 (N_9672,N_6421,N_7032);
xnor U9673 (N_9673,N_7384,N_7467);
nor U9674 (N_9674,N_7859,N_7857);
nor U9675 (N_9675,N_7705,N_7574);
nor U9676 (N_9676,N_6299,N_7723);
and U9677 (N_9677,N_7109,N_6793);
xor U9678 (N_9678,N_6086,N_6601);
nand U9679 (N_9679,N_6571,N_6795);
and U9680 (N_9680,N_6282,N_6738);
and U9681 (N_9681,N_6623,N_6774);
or U9682 (N_9682,N_6258,N_6240);
and U9683 (N_9683,N_7795,N_7900);
nor U9684 (N_9684,N_7483,N_6868);
nor U9685 (N_9685,N_7017,N_6869);
nand U9686 (N_9686,N_7415,N_7214);
or U9687 (N_9687,N_6587,N_7975);
nand U9688 (N_9688,N_6832,N_6738);
and U9689 (N_9689,N_7114,N_7360);
and U9690 (N_9690,N_6781,N_7227);
nand U9691 (N_9691,N_7526,N_7853);
and U9692 (N_9692,N_6013,N_7463);
xor U9693 (N_9693,N_7012,N_7757);
xor U9694 (N_9694,N_7915,N_7239);
and U9695 (N_9695,N_6833,N_6360);
nand U9696 (N_9696,N_7270,N_6494);
or U9697 (N_9697,N_7110,N_7421);
nand U9698 (N_9698,N_7589,N_6825);
nor U9699 (N_9699,N_7528,N_6356);
and U9700 (N_9700,N_6887,N_7474);
nand U9701 (N_9701,N_7722,N_6574);
nand U9702 (N_9702,N_7986,N_7975);
and U9703 (N_9703,N_6994,N_6158);
nor U9704 (N_9704,N_6547,N_6347);
nand U9705 (N_9705,N_7910,N_6788);
nor U9706 (N_9706,N_6284,N_6021);
nor U9707 (N_9707,N_7514,N_6730);
nand U9708 (N_9708,N_6646,N_7459);
and U9709 (N_9709,N_7401,N_7017);
nor U9710 (N_9710,N_6693,N_7448);
nand U9711 (N_9711,N_6536,N_6939);
nor U9712 (N_9712,N_7793,N_7414);
or U9713 (N_9713,N_6052,N_6609);
xor U9714 (N_9714,N_6110,N_7382);
or U9715 (N_9715,N_6330,N_7288);
or U9716 (N_9716,N_6068,N_7648);
nand U9717 (N_9717,N_7635,N_6151);
nand U9718 (N_9718,N_7505,N_6551);
and U9719 (N_9719,N_7319,N_6868);
nand U9720 (N_9720,N_6069,N_7469);
nor U9721 (N_9721,N_7522,N_7915);
nor U9722 (N_9722,N_7953,N_7611);
nor U9723 (N_9723,N_6347,N_6298);
nor U9724 (N_9724,N_7234,N_7707);
or U9725 (N_9725,N_7223,N_7102);
and U9726 (N_9726,N_7793,N_6567);
and U9727 (N_9727,N_7902,N_6020);
nor U9728 (N_9728,N_6204,N_7511);
and U9729 (N_9729,N_7480,N_7995);
or U9730 (N_9730,N_7266,N_6604);
nor U9731 (N_9731,N_6633,N_7232);
xnor U9732 (N_9732,N_7130,N_7721);
or U9733 (N_9733,N_6387,N_6512);
or U9734 (N_9734,N_6717,N_7737);
and U9735 (N_9735,N_7675,N_6880);
or U9736 (N_9736,N_7335,N_7790);
nand U9737 (N_9737,N_6966,N_7232);
nand U9738 (N_9738,N_7328,N_6541);
or U9739 (N_9739,N_6278,N_6171);
nand U9740 (N_9740,N_7018,N_7373);
and U9741 (N_9741,N_7537,N_7515);
nor U9742 (N_9742,N_7187,N_7997);
or U9743 (N_9743,N_7983,N_7425);
and U9744 (N_9744,N_6357,N_6976);
xnor U9745 (N_9745,N_7272,N_7064);
and U9746 (N_9746,N_6774,N_7643);
nor U9747 (N_9747,N_6099,N_6533);
or U9748 (N_9748,N_7473,N_7965);
nor U9749 (N_9749,N_7822,N_6116);
xnor U9750 (N_9750,N_7147,N_6108);
or U9751 (N_9751,N_7329,N_6159);
nor U9752 (N_9752,N_7804,N_6855);
or U9753 (N_9753,N_7009,N_7812);
and U9754 (N_9754,N_7225,N_6568);
or U9755 (N_9755,N_6449,N_7547);
nand U9756 (N_9756,N_7875,N_7219);
nor U9757 (N_9757,N_7168,N_6517);
or U9758 (N_9758,N_6881,N_7178);
and U9759 (N_9759,N_6600,N_7908);
nand U9760 (N_9760,N_7796,N_7865);
or U9761 (N_9761,N_6448,N_7948);
and U9762 (N_9762,N_6992,N_7274);
and U9763 (N_9763,N_6312,N_7419);
or U9764 (N_9764,N_6359,N_7345);
nand U9765 (N_9765,N_6816,N_7705);
or U9766 (N_9766,N_6519,N_6370);
nor U9767 (N_9767,N_7179,N_7807);
or U9768 (N_9768,N_6772,N_6342);
nor U9769 (N_9769,N_6445,N_6488);
and U9770 (N_9770,N_6112,N_7997);
nand U9771 (N_9771,N_7386,N_6869);
or U9772 (N_9772,N_6959,N_7175);
nor U9773 (N_9773,N_6706,N_6477);
or U9774 (N_9774,N_6258,N_7942);
and U9775 (N_9775,N_6484,N_7859);
or U9776 (N_9776,N_6609,N_6716);
and U9777 (N_9777,N_7006,N_6151);
or U9778 (N_9778,N_6500,N_7883);
nor U9779 (N_9779,N_6261,N_7791);
and U9780 (N_9780,N_7719,N_7667);
and U9781 (N_9781,N_7849,N_7334);
nor U9782 (N_9782,N_7133,N_6337);
nand U9783 (N_9783,N_7297,N_7210);
and U9784 (N_9784,N_6402,N_7086);
or U9785 (N_9785,N_7580,N_6946);
nand U9786 (N_9786,N_7250,N_6974);
and U9787 (N_9787,N_7131,N_6558);
and U9788 (N_9788,N_6461,N_7846);
nand U9789 (N_9789,N_7005,N_7238);
xor U9790 (N_9790,N_7640,N_7525);
or U9791 (N_9791,N_7603,N_7287);
xor U9792 (N_9792,N_6773,N_7402);
nor U9793 (N_9793,N_6804,N_7163);
nand U9794 (N_9794,N_7605,N_6761);
or U9795 (N_9795,N_6247,N_6392);
and U9796 (N_9796,N_6073,N_6185);
nor U9797 (N_9797,N_6354,N_7394);
nand U9798 (N_9798,N_7727,N_6830);
nor U9799 (N_9799,N_6030,N_6049);
and U9800 (N_9800,N_6215,N_7268);
nand U9801 (N_9801,N_7728,N_7346);
nand U9802 (N_9802,N_6752,N_7535);
or U9803 (N_9803,N_6418,N_6311);
or U9804 (N_9804,N_6244,N_7969);
nor U9805 (N_9805,N_6923,N_6150);
nand U9806 (N_9806,N_7266,N_7269);
nand U9807 (N_9807,N_6477,N_6762);
or U9808 (N_9808,N_7360,N_6783);
or U9809 (N_9809,N_7482,N_6090);
or U9810 (N_9810,N_7052,N_7224);
and U9811 (N_9811,N_7241,N_6861);
and U9812 (N_9812,N_7789,N_7880);
nand U9813 (N_9813,N_7582,N_7514);
or U9814 (N_9814,N_6075,N_7137);
and U9815 (N_9815,N_6939,N_7484);
or U9816 (N_9816,N_6020,N_6386);
or U9817 (N_9817,N_7839,N_6979);
or U9818 (N_9818,N_6469,N_7926);
nand U9819 (N_9819,N_7250,N_7596);
or U9820 (N_9820,N_6784,N_6475);
and U9821 (N_9821,N_6389,N_6537);
and U9822 (N_9822,N_6673,N_7425);
nor U9823 (N_9823,N_7530,N_6573);
nor U9824 (N_9824,N_7912,N_6064);
or U9825 (N_9825,N_6042,N_7146);
nor U9826 (N_9826,N_7988,N_7040);
nor U9827 (N_9827,N_6829,N_7157);
and U9828 (N_9828,N_6914,N_6709);
and U9829 (N_9829,N_6108,N_7452);
nand U9830 (N_9830,N_6254,N_7676);
and U9831 (N_9831,N_6839,N_6072);
xnor U9832 (N_9832,N_6859,N_7809);
or U9833 (N_9833,N_7043,N_7066);
or U9834 (N_9834,N_7563,N_7959);
nand U9835 (N_9835,N_6403,N_7618);
nor U9836 (N_9836,N_6487,N_7592);
nor U9837 (N_9837,N_6556,N_6345);
nand U9838 (N_9838,N_7320,N_6460);
nor U9839 (N_9839,N_7724,N_7582);
nand U9840 (N_9840,N_7127,N_7774);
or U9841 (N_9841,N_6120,N_6093);
or U9842 (N_9842,N_6683,N_7122);
nor U9843 (N_9843,N_7695,N_7026);
xnor U9844 (N_9844,N_7235,N_7091);
and U9845 (N_9845,N_7278,N_6100);
nor U9846 (N_9846,N_7037,N_6932);
nor U9847 (N_9847,N_6998,N_7757);
nor U9848 (N_9848,N_7337,N_6731);
or U9849 (N_9849,N_6662,N_7821);
xor U9850 (N_9850,N_6398,N_7043);
and U9851 (N_9851,N_7267,N_7545);
nor U9852 (N_9852,N_6018,N_6337);
or U9853 (N_9853,N_6042,N_7440);
nor U9854 (N_9854,N_6964,N_6854);
and U9855 (N_9855,N_7133,N_7983);
nand U9856 (N_9856,N_7735,N_6149);
or U9857 (N_9857,N_6372,N_7896);
or U9858 (N_9858,N_6096,N_6669);
nor U9859 (N_9859,N_6818,N_7537);
or U9860 (N_9860,N_6849,N_7227);
xnor U9861 (N_9861,N_7302,N_6071);
or U9862 (N_9862,N_6847,N_7017);
nand U9863 (N_9863,N_6456,N_7112);
or U9864 (N_9864,N_6362,N_7872);
nand U9865 (N_9865,N_7037,N_6944);
and U9866 (N_9866,N_7016,N_6447);
nand U9867 (N_9867,N_6854,N_7242);
nand U9868 (N_9868,N_6730,N_6383);
nor U9869 (N_9869,N_6956,N_6634);
and U9870 (N_9870,N_6555,N_6225);
and U9871 (N_9871,N_6876,N_7147);
or U9872 (N_9872,N_7402,N_6261);
or U9873 (N_9873,N_6388,N_7288);
nand U9874 (N_9874,N_7079,N_6825);
or U9875 (N_9875,N_6352,N_6577);
and U9876 (N_9876,N_7098,N_6833);
nand U9877 (N_9877,N_7838,N_6802);
and U9878 (N_9878,N_7851,N_6392);
and U9879 (N_9879,N_7760,N_7366);
and U9880 (N_9880,N_6301,N_6731);
xnor U9881 (N_9881,N_7747,N_6302);
or U9882 (N_9882,N_6162,N_7437);
and U9883 (N_9883,N_7477,N_6618);
nand U9884 (N_9884,N_6182,N_7983);
nand U9885 (N_9885,N_6575,N_7564);
and U9886 (N_9886,N_7397,N_7018);
nor U9887 (N_9887,N_7931,N_6676);
or U9888 (N_9888,N_6989,N_7931);
nor U9889 (N_9889,N_6861,N_7235);
and U9890 (N_9890,N_6188,N_6947);
nand U9891 (N_9891,N_6334,N_6052);
nor U9892 (N_9892,N_6569,N_7293);
nor U9893 (N_9893,N_6076,N_7431);
nand U9894 (N_9894,N_7597,N_7086);
nand U9895 (N_9895,N_7232,N_6902);
or U9896 (N_9896,N_7775,N_6900);
nor U9897 (N_9897,N_7379,N_6706);
nor U9898 (N_9898,N_6985,N_7076);
nor U9899 (N_9899,N_6156,N_7025);
and U9900 (N_9900,N_7767,N_7801);
nand U9901 (N_9901,N_6694,N_6060);
and U9902 (N_9902,N_6542,N_6511);
or U9903 (N_9903,N_6957,N_6453);
or U9904 (N_9904,N_7892,N_6828);
nor U9905 (N_9905,N_6669,N_6876);
and U9906 (N_9906,N_6467,N_6554);
nand U9907 (N_9907,N_7218,N_7924);
or U9908 (N_9908,N_7738,N_7190);
nor U9909 (N_9909,N_6073,N_6656);
nand U9910 (N_9910,N_6322,N_7166);
xnor U9911 (N_9911,N_7571,N_7498);
or U9912 (N_9912,N_6824,N_6490);
nor U9913 (N_9913,N_6514,N_7034);
nand U9914 (N_9914,N_7282,N_7443);
or U9915 (N_9915,N_6460,N_7388);
xor U9916 (N_9916,N_7690,N_6350);
nand U9917 (N_9917,N_7711,N_6699);
xnor U9918 (N_9918,N_7758,N_6950);
and U9919 (N_9919,N_7833,N_6554);
and U9920 (N_9920,N_7022,N_6450);
nor U9921 (N_9921,N_7365,N_6496);
and U9922 (N_9922,N_7683,N_6440);
or U9923 (N_9923,N_7471,N_7289);
nand U9924 (N_9924,N_6223,N_6642);
nor U9925 (N_9925,N_7977,N_7855);
and U9926 (N_9926,N_6123,N_6926);
nor U9927 (N_9927,N_6271,N_7772);
and U9928 (N_9928,N_7685,N_7687);
nor U9929 (N_9929,N_6260,N_7016);
xor U9930 (N_9930,N_7350,N_6909);
xnor U9931 (N_9931,N_6794,N_6999);
and U9932 (N_9932,N_7350,N_7010);
nand U9933 (N_9933,N_7777,N_7642);
or U9934 (N_9934,N_6174,N_7500);
and U9935 (N_9935,N_6590,N_6136);
nor U9936 (N_9936,N_7038,N_6983);
nor U9937 (N_9937,N_7750,N_6625);
or U9938 (N_9938,N_6107,N_7962);
nor U9939 (N_9939,N_7449,N_7682);
or U9940 (N_9940,N_7581,N_7066);
nor U9941 (N_9941,N_6500,N_7126);
nand U9942 (N_9942,N_7223,N_6033);
nand U9943 (N_9943,N_6337,N_6962);
and U9944 (N_9944,N_6852,N_7775);
xor U9945 (N_9945,N_6010,N_7024);
or U9946 (N_9946,N_6042,N_7984);
and U9947 (N_9947,N_6992,N_7044);
nor U9948 (N_9948,N_7555,N_7362);
or U9949 (N_9949,N_6819,N_6837);
nor U9950 (N_9950,N_6224,N_7570);
nor U9951 (N_9951,N_6364,N_6331);
and U9952 (N_9952,N_6279,N_6511);
nor U9953 (N_9953,N_7011,N_7219);
or U9954 (N_9954,N_7645,N_7907);
and U9955 (N_9955,N_7654,N_6598);
and U9956 (N_9956,N_6770,N_6500);
nand U9957 (N_9957,N_7130,N_6095);
nand U9958 (N_9958,N_6077,N_6025);
nor U9959 (N_9959,N_6877,N_7103);
nand U9960 (N_9960,N_6909,N_7094);
nor U9961 (N_9961,N_6476,N_6824);
nand U9962 (N_9962,N_7105,N_6892);
nand U9963 (N_9963,N_7312,N_6414);
and U9964 (N_9964,N_7153,N_6769);
or U9965 (N_9965,N_7585,N_7942);
xnor U9966 (N_9966,N_6067,N_7885);
or U9967 (N_9967,N_7846,N_6041);
nor U9968 (N_9968,N_6350,N_6200);
or U9969 (N_9969,N_7598,N_6290);
and U9970 (N_9970,N_7804,N_7046);
nand U9971 (N_9971,N_6748,N_7567);
nor U9972 (N_9972,N_7378,N_6788);
or U9973 (N_9973,N_6939,N_7774);
and U9974 (N_9974,N_6876,N_6957);
nand U9975 (N_9975,N_7313,N_6476);
nor U9976 (N_9976,N_6483,N_6809);
or U9977 (N_9977,N_6596,N_6413);
or U9978 (N_9978,N_7288,N_7043);
nand U9979 (N_9979,N_7829,N_6503);
nand U9980 (N_9980,N_6473,N_6757);
xor U9981 (N_9981,N_7635,N_7556);
nand U9982 (N_9982,N_6807,N_7795);
or U9983 (N_9983,N_6762,N_6938);
nor U9984 (N_9984,N_7992,N_7133);
and U9985 (N_9985,N_7157,N_7395);
or U9986 (N_9986,N_6541,N_7391);
nor U9987 (N_9987,N_6518,N_7243);
and U9988 (N_9988,N_7451,N_7898);
nand U9989 (N_9989,N_7650,N_7900);
nand U9990 (N_9990,N_7755,N_6106);
or U9991 (N_9991,N_6054,N_6374);
or U9992 (N_9992,N_7330,N_6848);
nand U9993 (N_9993,N_6253,N_6109);
nand U9994 (N_9994,N_7114,N_7544);
nor U9995 (N_9995,N_7329,N_6987);
nand U9996 (N_9996,N_6811,N_6234);
xor U9997 (N_9997,N_6896,N_7030);
or U9998 (N_9998,N_7888,N_7366);
or U9999 (N_9999,N_6455,N_6580);
xnor U10000 (N_10000,N_9036,N_9374);
nand U10001 (N_10001,N_9411,N_8873);
nor U10002 (N_10002,N_8303,N_8182);
nor U10003 (N_10003,N_8386,N_8753);
and U10004 (N_10004,N_9730,N_9475);
xnor U10005 (N_10005,N_9797,N_9071);
xor U10006 (N_10006,N_8148,N_8054);
xnor U10007 (N_10007,N_8991,N_8890);
xnor U10008 (N_10008,N_9487,N_9093);
nor U10009 (N_10009,N_9329,N_9896);
nand U10010 (N_10010,N_8381,N_9554);
nor U10011 (N_10011,N_8447,N_8319);
nor U10012 (N_10012,N_9553,N_9031);
and U10013 (N_10013,N_8704,N_8814);
and U10014 (N_10014,N_8894,N_9306);
nand U10015 (N_10015,N_9027,N_9178);
or U10016 (N_10016,N_9349,N_8389);
nor U10017 (N_10017,N_9160,N_8938);
and U10018 (N_10018,N_8458,N_8237);
and U10019 (N_10019,N_9425,N_8837);
nand U10020 (N_10020,N_8394,N_8732);
and U10021 (N_10021,N_8106,N_8820);
nand U10022 (N_10022,N_9701,N_8209);
nand U10023 (N_10023,N_8642,N_9422);
or U10024 (N_10024,N_9972,N_9074);
or U10025 (N_10025,N_8507,N_8798);
nor U10026 (N_10026,N_9585,N_8758);
and U10027 (N_10027,N_9398,N_8183);
nor U10028 (N_10028,N_9895,N_9853);
nor U10029 (N_10029,N_9357,N_9571);
xor U10030 (N_10030,N_8214,N_9700);
and U10031 (N_10031,N_9076,N_9614);
nand U10032 (N_10032,N_9932,N_8002);
nand U10033 (N_10033,N_8055,N_9898);
and U10034 (N_10034,N_9302,N_8573);
and U10035 (N_10035,N_8752,N_9197);
and U10036 (N_10036,N_9156,N_9819);
xor U10037 (N_10037,N_9780,N_9207);
and U10038 (N_10038,N_8360,N_8056);
nor U10039 (N_10039,N_8454,N_8527);
nand U10040 (N_10040,N_9957,N_8526);
nand U10041 (N_10041,N_9118,N_9698);
nand U10042 (N_10042,N_8062,N_9865);
or U10043 (N_10043,N_8750,N_9666);
xnor U10044 (N_10044,N_8039,N_8441);
nand U10045 (N_10045,N_9758,N_9619);
or U10046 (N_10046,N_9460,N_9454);
xor U10047 (N_10047,N_8504,N_8057);
nand U10048 (N_10048,N_9963,N_9172);
and U10049 (N_10049,N_9401,N_9053);
or U10050 (N_10050,N_8627,N_8866);
nand U10051 (N_10051,N_8726,N_8302);
nor U10052 (N_10052,N_8058,N_9580);
xor U10053 (N_10053,N_8396,N_8265);
nor U10054 (N_10054,N_9991,N_9163);
nand U10055 (N_10055,N_8013,N_9385);
or U10056 (N_10056,N_8023,N_9908);
nand U10057 (N_10057,N_9808,N_9511);
and U10058 (N_10058,N_9778,N_9362);
and U10059 (N_10059,N_8180,N_8179);
xor U10060 (N_10060,N_9826,N_8562);
nor U10061 (N_10061,N_9912,N_9843);
and U10062 (N_10062,N_8595,N_8286);
or U10063 (N_10063,N_9337,N_9540);
and U10064 (N_10064,N_9065,N_8287);
and U10065 (N_10065,N_9890,N_9879);
nor U10066 (N_10066,N_8468,N_9674);
or U10067 (N_10067,N_9442,N_8639);
nor U10068 (N_10068,N_9413,N_8564);
or U10069 (N_10069,N_9380,N_9870);
or U10070 (N_10070,N_9873,N_9276);
nor U10071 (N_10071,N_9951,N_8486);
nand U10072 (N_10072,N_8212,N_9564);
or U10073 (N_10073,N_8865,N_9849);
and U10074 (N_10074,N_9394,N_9145);
nor U10075 (N_10075,N_9303,N_8030);
or U10076 (N_10076,N_8082,N_8397);
or U10077 (N_10077,N_9747,N_8464);
or U10078 (N_10078,N_9596,N_8083);
nor U10079 (N_10079,N_9222,N_8554);
or U10080 (N_10080,N_8605,N_9250);
and U10081 (N_10081,N_9646,N_8980);
nand U10082 (N_10082,N_9805,N_8843);
nor U10083 (N_10083,N_9907,N_8177);
or U10084 (N_10084,N_8952,N_9673);
nand U10085 (N_10085,N_9625,N_9419);
nor U10086 (N_10086,N_9948,N_8232);
xnor U10087 (N_10087,N_9950,N_8090);
or U10088 (N_10088,N_8757,N_9760);
or U10089 (N_10089,N_9902,N_9939);
nand U10090 (N_10090,N_8384,N_8373);
and U10091 (N_10091,N_9520,N_8835);
or U10092 (N_10092,N_9059,N_9347);
xor U10093 (N_10093,N_9204,N_9359);
and U10094 (N_10094,N_8707,N_8939);
or U10095 (N_10095,N_9886,N_8742);
nor U10096 (N_10096,N_8300,N_9878);
nand U10097 (N_10097,N_8785,N_9954);
nand U10098 (N_10098,N_8216,N_8594);
nand U10099 (N_10099,N_9196,N_9308);
nand U10100 (N_10100,N_8660,N_8724);
nand U10101 (N_10101,N_9952,N_8816);
nor U10102 (N_10102,N_8471,N_8080);
or U10103 (N_10103,N_8756,N_8987);
and U10104 (N_10104,N_9899,N_9874);
and U10105 (N_10105,N_8599,N_9693);
xor U10106 (N_10106,N_8277,N_9180);
and U10107 (N_10107,N_8824,N_9785);
nor U10108 (N_10108,N_8141,N_9736);
and U10109 (N_10109,N_9533,N_8734);
nand U10110 (N_10110,N_8174,N_9927);
nor U10111 (N_10111,N_9705,N_8221);
and U10112 (N_10112,N_9630,N_9566);
xnor U10113 (N_10113,N_8637,N_9535);
nand U10114 (N_10114,N_9491,N_9035);
and U10115 (N_10115,N_8646,N_8689);
xor U10116 (N_10116,N_9561,N_9288);
and U10117 (N_10117,N_9488,N_8235);
or U10118 (N_10118,N_8603,N_9299);
and U10119 (N_10119,N_9942,N_8040);
nand U10120 (N_10120,N_8923,N_8936);
nor U10121 (N_10121,N_9236,N_9775);
or U10122 (N_10122,N_9828,N_9706);
or U10123 (N_10123,N_9749,N_9690);
nand U10124 (N_10124,N_9502,N_8391);
nand U10125 (N_10125,N_9721,N_9193);
and U10126 (N_10126,N_9549,N_8518);
nor U10127 (N_10127,N_8268,N_8898);
or U10128 (N_10128,N_9798,N_9530);
or U10129 (N_10129,N_9993,N_9528);
xnor U10130 (N_10130,N_9212,N_8499);
and U10131 (N_10131,N_8596,N_9069);
or U10132 (N_10132,N_8116,N_8585);
and U10133 (N_10133,N_9113,N_8781);
and U10134 (N_10134,N_8679,N_8297);
nor U10135 (N_10135,N_9218,N_8826);
nand U10136 (N_10136,N_8383,N_8634);
nor U10137 (N_10137,N_8238,N_8537);
nor U10138 (N_10138,N_8289,N_8570);
or U10139 (N_10139,N_9296,N_8694);
xor U10140 (N_10140,N_8111,N_9396);
xnor U10141 (N_10141,N_9844,N_8004);
xor U10142 (N_10142,N_8661,N_8893);
nand U10143 (N_10143,N_9365,N_9788);
nor U10144 (N_10144,N_8399,N_9022);
or U10145 (N_10145,N_8346,N_9096);
nand U10146 (N_10146,N_8986,N_8509);
nor U10147 (N_10147,N_9930,N_8130);
nor U10148 (N_10148,N_8043,N_9161);
and U10149 (N_10149,N_9921,N_9311);
or U10150 (N_10150,N_9806,N_8012);
nand U10151 (N_10151,N_9301,N_8444);
or U10152 (N_10152,N_9710,N_8198);
or U10153 (N_10153,N_9709,N_8892);
or U10154 (N_10154,N_8610,N_8985);
or U10155 (N_10155,N_8476,N_9718);
or U10156 (N_10156,N_8768,N_8071);
and U10157 (N_10157,N_8921,N_8547);
nand U10158 (N_10158,N_9838,N_9327);
or U10159 (N_10159,N_9143,N_9795);
and U10160 (N_10160,N_8204,N_8871);
nand U10161 (N_10161,N_8484,N_8717);
xor U10162 (N_10162,N_9132,N_9312);
nor U10163 (N_10163,N_9195,N_9015);
xor U10164 (N_10164,N_8850,N_9485);
and U10165 (N_10165,N_8560,N_9041);
nor U10166 (N_10166,N_9771,N_9624);
and U10167 (N_10167,N_8127,N_9174);
and U10168 (N_10168,N_9068,N_9131);
or U10169 (N_10169,N_8548,N_8510);
nand U10170 (N_10170,N_8928,N_9050);
and U10171 (N_10171,N_9964,N_9432);
nor U10172 (N_10172,N_8948,N_9547);
or U10173 (N_10173,N_9237,N_8167);
and U10174 (N_10174,N_9078,N_8354);
and U10175 (N_10175,N_8010,N_9555);
nor U10176 (N_10176,N_8147,N_9228);
nand U10177 (N_10177,N_8641,N_8613);
nor U10178 (N_10178,N_8940,N_9338);
nand U10179 (N_10179,N_8431,N_8736);
nor U10180 (N_10180,N_8579,N_9756);
or U10181 (N_10181,N_8188,N_8359);
nand U10182 (N_10182,N_8625,N_8546);
and U10183 (N_10183,N_8173,N_9522);
nor U10184 (N_10184,N_8291,N_8496);
nand U10185 (N_10185,N_8981,N_8203);
or U10186 (N_10186,N_9043,N_8154);
nor U10187 (N_10187,N_8839,N_8448);
nor U10188 (N_10188,N_8440,N_8999);
nor U10189 (N_10189,N_8908,N_8869);
nand U10190 (N_10190,N_8979,N_8421);
and U10191 (N_10191,N_8022,N_9184);
and U10192 (N_10192,N_9017,N_9375);
nand U10193 (N_10193,N_9591,N_8954);
and U10194 (N_10194,N_8915,N_8793);
xor U10195 (N_10195,N_8126,N_8746);
nand U10196 (N_10196,N_9168,N_8701);
and U10197 (N_10197,N_8305,N_9428);
and U10198 (N_10198,N_9602,N_9367);
and U10199 (N_10199,N_8900,N_9594);
and U10200 (N_10200,N_9650,N_9998);
and U10201 (N_10201,N_8483,N_8868);
or U10202 (N_10202,N_9242,N_8118);
nor U10203 (N_10203,N_9965,N_8153);
and U10204 (N_10204,N_8827,N_8025);
or U10205 (N_10205,N_8419,N_9608);
xnor U10206 (N_10206,N_9309,N_9020);
and U10207 (N_10207,N_9514,N_8345);
xor U10208 (N_10208,N_9983,N_8593);
or U10209 (N_10209,N_9493,N_9344);
or U10210 (N_10210,N_9711,N_9012);
nand U10211 (N_10211,N_8787,N_8206);
and U10212 (N_10212,N_9929,N_9019);
and U10213 (N_10213,N_9298,N_9370);
and U10214 (N_10214,N_8145,N_8912);
nand U10215 (N_10215,N_9975,N_9745);
nor U10216 (N_10216,N_9509,N_9264);
nand U10217 (N_10217,N_9453,N_8129);
and U10218 (N_10218,N_9351,N_8122);
nor U10219 (N_10219,N_8505,N_8103);
or U10220 (N_10220,N_8965,N_8133);
nand U10221 (N_10221,N_9960,N_9979);
and U10222 (N_10222,N_9284,N_9007);
nor U10223 (N_10223,N_8571,N_9823);
or U10224 (N_10224,N_8971,N_9784);
or U10225 (N_10225,N_9616,N_8308);
and U10226 (N_10226,N_8748,N_8765);
nor U10227 (N_10227,N_9787,N_9770);
or U10228 (N_10228,N_8540,N_9116);
nor U10229 (N_10229,N_9044,N_8864);
or U10230 (N_10230,N_8121,N_8407);
and U10231 (N_10231,N_8503,N_9618);
and U10232 (N_10232,N_8693,N_9513);
nand U10233 (N_10233,N_8318,N_9025);
nor U10234 (N_10234,N_9166,N_8060);
nor U10235 (N_10235,N_8759,N_8513);
xnor U10236 (N_10236,N_9424,N_9829);
or U10237 (N_10237,N_9595,N_9791);
and U10238 (N_10238,N_8353,N_8333);
nand U10239 (N_10239,N_9063,N_8716);
or U10240 (N_10240,N_9361,N_9822);
nor U10241 (N_10241,N_8463,N_9437);
nand U10242 (N_10242,N_9576,N_9371);
nor U10243 (N_10243,N_8805,N_8493);
nand U10244 (N_10244,N_9271,N_8737);
nor U10245 (N_10245,N_8490,N_8810);
or U10246 (N_10246,N_9497,N_8261);
nor U10247 (N_10247,N_9639,N_8208);
nor U10248 (N_10248,N_9407,N_8451);
nand U10249 (N_10249,N_8671,N_8608);
and U10250 (N_10250,N_9740,N_9702);
xnor U10251 (N_10251,N_8973,N_8684);
nor U10252 (N_10252,N_8115,N_8280);
and U10253 (N_10253,N_8164,N_8534);
nor U10254 (N_10254,N_8522,N_9042);
or U10255 (N_10255,N_8352,N_8229);
xnor U10256 (N_10256,N_8446,N_9423);
or U10257 (N_10257,N_8320,N_8310);
and U10258 (N_10258,N_9275,N_9612);
or U10259 (N_10259,N_8665,N_8512);
nand U10260 (N_10260,N_9542,N_8783);
nand U10261 (N_10261,N_9794,N_9274);
and U10262 (N_10262,N_9056,N_8970);
xnor U10263 (N_10263,N_9606,N_9003);
and U10264 (N_10264,N_8993,N_9691);
or U10265 (N_10265,N_8770,N_9974);
nor U10266 (N_10266,N_9130,N_8663);
nand U10267 (N_10267,N_8744,N_9609);
or U10268 (N_10268,N_9776,N_8977);
nor U10269 (N_10269,N_9915,N_9820);
or U10270 (N_10270,N_8779,N_8213);
nand U10271 (N_10271,N_8323,N_8623);
and U10272 (N_10272,N_9656,N_9928);
nand U10273 (N_10273,N_8844,N_9845);
nand U10274 (N_10274,N_8687,N_8713);
and U10275 (N_10275,N_9482,N_9583);
nand U10276 (N_10276,N_8363,N_9897);
nor U10277 (N_10277,N_9165,N_9343);
nand U10278 (N_10278,N_8508,N_9953);
xor U10279 (N_10279,N_9047,N_8371);
nand U10280 (N_10280,N_9457,N_8053);
or U10281 (N_10281,N_9456,N_9668);
nand U10282 (N_10282,N_8739,N_9500);
and U10283 (N_10283,N_9431,N_9144);
xor U10284 (N_10284,N_9640,N_9499);
nor U10285 (N_10285,N_9107,N_9969);
nand U10286 (N_10286,N_8574,N_9722);
nand U10287 (N_10287,N_8190,N_8307);
nand U10288 (N_10288,N_9598,N_8215);
and U10289 (N_10289,N_9438,N_9280);
nand U10290 (N_10290,N_9120,N_9647);
or U10291 (N_10291,N_8852,N_9529);
nor U10292 (N_10292,N_9094,N_9725);
xor U10293 (N_10293,N_9089,N_9436);
and U10294 (N_10294,N_9379,N_9495);
xor U10295 (N_10295,N_9082,N_9100);
xnor U10296 (N_10296,N_9333,N_8601);
nor U10297 (N_10297,N_8523,N_8664);
nand U10298 (N_10298,N_9988,N_8897);
xnor U10299 (N_10299,N_8450,N_9133);
nor U10300 (N_10300,N_8643,N_8604);
and U10301 (N_10301,N_9956,N_8968);
or U10302 (N_10302,N_9038,N_8920);
and U10303 (N_10303,N_9779,N_9006);
nand U10304 (N_10304,N_8259,N_9449);
or U10305 (N_10305,N_8566,N_8740);
nand U10306 (N_10306,N_9016,N_8628);
nor U10307 (N_10307,N_8249,N_9317);
and U10308 (N_10308,N_9512,N_8761);
or U10309 (N_10309,N_8146,N_8851);
nand U10310 (N_10310,N_8943,N_8715);
nand U10311 (N_10311,N_9090,N_8926);
or U10312 (N_10312,N_8647,N_8015);
nand U10313 (N_10313,N_8581,N_8831);
nand U10314 (N_10314,N_9860,N_8568);
or U10315 (N_10315,N_9119,N_9814);
xnor U10316 (N_10316,N_8413,N_8000);
xnor U10317 (N_10317,N_9737,N_9137);
xnor U10318 (N_10318,N_8963,N_8166);
or U10319 (N_10319,N_8863,N_8036);
or U10320 (N_10320,N_8804,N_8150);
or U10321 (N_10321,N_9395,N_8364);
and U10322 (N_10322,N_9416,N_8487);
nor U10323 (N_10323,N_9507,N_8078);
xnor U10324 (N_10324,N_9384,N_9005);
or U10325 (N_10325,N_9281,N_8836);
nand U10326 (N_10326,N_9240,N_8005);
or U10327 (N_10327,N_9238,N_9732);
nor U10328 (N_10328,N_8370,N_8161);
nor U10329 (N_10329,N_9225,N_8872);
and U10330 (N_10330,N_8224,N_8369);
and U10331 (N_10331,N_8932,N_8408);
nand U10332 (N_10332,N_9523,N_8008);
or U10333 (N_10333,N_9996,N_8372);
nand U10334 (N_10334,N_8191,N_9095);
nor U10335 (N_10335,N_8230,N_9962);
nand U10336 (N_10336,N_8218,N_8640);
and U10337 (N_10337,N_8442,N_9318);
nor U10338 (N_10338,N_9961,N_9628);
nand U10339 (N_10339,N_9526,N_8387);
or U10340 (N_10340,N_8223,N_9662);
and U10341 (N_10341,N_8561,N_8632);
or U10342 (N_10342,N_8226,N_9182);
xor U10343 (N_10343,N_8652,N_9154);
nor U10344 (N_10344,N_9105,N_8176);
xnor U10345 (N_10345,N_9450,N_9903);
nand U10346 (N_10346,N_9735,N_8375);
or U10347 (N_10347,N_8855,N_8849);
or U10348 (N_10348,N_8047,N_9092);
or U10349 (N_10349,N_8806,N_9048);
and U10350 (N_10350,N_8847,N_8211);
and U10351 (N_10351,N_8031,N_8418);
or U10352 (N_10352,N_9479,N_9346);
nand U10353 (N_10353,N_9088,N_8611);
nand U10354 (N_10354,N_8482,N_9943);
and U10355 (N_10355,N_9273,N_8065);
nand U10356 (N_10356,N_8813,N_9136);
nand U10357 (N_10357,N_9660,N_9014);
and U10358 (N_10358,N_8735,N_8254);
nor U10359 (N_10359,N_9834,N_8983);
or U10360 (N_10360,N_9590,N_8492);
nand U10361 (N_10361,N_8324,N_8175);
and U10362 (N_10362,N_8901,N_9128);
nand U10363 (N_10363,N_9049,N_9739);
nor U10364 (N_10364,N_8747,N_9231);
and U10365 (N_10365,N_8003,N_8317);
and U10366 (N_10366,N_9905,N_8829);
xor U10367 (N_10367,N_8631,N_8279);
or U10368 (N_10368,N_9987,N_8157);
or U10369 (N_10369,N_8449,N_9148);
nor U10370 (N_10370,N_8621,N_8690);
and U10371 (N_10371,N_8168,N_8457);
xor U10372 (N_10372,N_9075,N_8020);
or U10373 (N_10373,N_8197,N_8135);
nor U10374 (N_10374,N_9773,N_9310);
nand U10375 (N_10375,N_8597,N_9170);
nor U10376 (N_10376,N_9233,N_8911);
nor U10377 (N_10377,N_8799,N_8234);
or U10378 (N_10378,N_8772,N_9358);
or U10379 (N_10379,N_9919,N_9187);
and U10380 (N_10380,N_8348,N_9813);
nor U10381 (N_10381,N_8019,N_8244);
and U10382 (N_10382,N_9129,N_8142);
and U10383 (N_10383,N_9633,N_8536);
nand U10384 (N_10384,N_8087,N_9435);
xnor U10385 (N_10385,N_9984,N_9415);
xnor U10386 (N_10386,N_8958,N_9750);
nand U10387 (N_10387,N_9629,N_8972);
or U10388 (N_10388,N_8708,N_9510);
and U10389 (N_10389,N_9536,N_9752);
and U10390 (N_10390,N_9832,N_9186);
nand U10391 (N_10391,N_8430,N_8434);
nor U10392 (N_10392,N_9597,N_8933);
or U10393 (N_10393,N_8606,N_9686);
and U10394 (N_10394,N_8124,N_9469);
nor U10395 (N_10395,N_8411,N_9888);
xor U10396 (N_10396,N_9158,N_9642);
or U10397 (N_10397,N_9652,N_9386);
xnor U10398 (N_10398,N_8098,N_9517);
or U10399 (N_10399,N_8825,N_9966);
or U10400 (N_10400,N_8170,N_8755);
and U10401 (N_10401,N_9149,N_9657);
and U10402 (N_10402,N_9173,N_9470);
and U10403 (N_10403,N_9191,N_8644);
nor U10404 (N_10404,N_9570,N_8709);
nand U10405 (N_10405,N_8455,N_9489);
nand U10406 (N_10406,N_8338,N_8158);
nor U10407 (N_10407,N_9644,N_9257);
nor U10408 (N_10408,N_9150,N_8169);
or U10409 (N_10409,N_8361,N_9188);
xnor U10410 (N_10410,N_8720,N_8366);
nand U10411 (N_10411,N_8104,N_9326);
xnor U10412 (N_10412,N_9887,N_8882);
or U10413 (N_10413,N_9104,N_9671);
xor U10414 (N_10414,N_8994,N_9029);
and U10415 (N_10415,N_9334,N_8883);
or U10416 (N_10416,N_8151,N_8710);
xor U10417 (N_10417,N_9356,N_9541);
and U10418 (N_10418,N_8041,N_8842);
nand U10419 (N_10419,N_9408,N_8559);
and U10420 (N_10420,N_8018,N_9947);
nand U10421 (N_10421,N_9655,N_8809);
nor U10422 (N_10422,N_9263,N_8329);
and U10423 (N_10423,N_9505,N_9039);
or U10424 (N_10424,N_9377,N_9654);
and U10425 (N_10425,N_9283,N_9402);
nor U10426 (N_10426,N_9861,N_9588);
and U10427 (N_10427,N_9492,N_9224);
nor U10428 (N_10428,N_8026,N_9913);
nand U10429 (N_10429,N_8341,N_8501);
and U10430 (N_10430,N_9501,N_8967);
nand U10431 (N_10431,N_8269,N_9243);
nand U10432 (N_10432,N_9474,N_9252);
nand U10433 (N_10433,N_9971,N_9748);
nand U10434 (N_10434,N_9325,N_9751);
xor U10435 (N_10435,N_9831,N_9297);
nand U10436 (N_10436,N_9840,N_9692);
or U10437 (N_10437,N_8674,N_8475);
and U10438 (N_10438,N_9884,N_9316);
nor U10439 (N_10439,N_9680,N_9645);
and U10440 (N_10440,N_9909,N_9430);
or U10441 (N_10441,N_9551,N_9232);
nand U10442 (N_10442,N_9269,N_9615);
xor U10443 (N_10443,N_9171,N_8095);
or U10444 (N_10444,N_8405,N_8472);
nand U10445 (N_10445,N_9743,N_8944);
and U10446 (N_10446,N_8001,N_8480);
and U10447 (N_10447,N_9135,N_9285);
nand U10448 (N_10448,N_8466,N_8706);
xor U10449 (N_10449,N_9997,N_9889);
and U10450 (N_10450,N_8243,N_9990);
nand U10451 (N_10451,N_9578,N_9060);
nand U10452 (N_10452,N_9175,N_8807);
or U10453 (N_10453,N_8347,N_9382);
nand U10454 (N_10454,N_8281,N_8273);
and U10455 (N_10455,N_8990,N_8395);
nand U10456 (N_10456,N_9550,N_9759);
nand U10457 (N_10457,N_8553,N_9681);
or U10458 (N_10458,N_8262,N_9933);
or U10459 (N_10459,N_9314,N_8042);
or U10460 (N_10460,N_9841,N_9409);
or U10461 (N_10461,N_8006,N_8903);
nor U10462 (N_10462,N_9894,N_9804);
and U10463 (N_10463,N_8888,N_8946);
nor U10464 (N_10464,N_8766,N_8107);
nand U10465 (N_10465,N_8196,N_8439);
nor U10466 (N_10466,N_8034,N_8859);
nor U10467 (N_10467,N_9321,N_9295);
xor U10468 (N_10468,N_9605,N_8296);
and U10469 (N_10469,N_9342,N_8648);
and U10470 (N_10470,N_9286,N_8511);
or U10471 (N_10471,N_8741,N_9123);
nor U10472 (N_10472,N_9600,N_8830);
nor U10473 (N_10473,N_9293,N_9440);
nor U10474 (N_10474,N_9715,N_8557);
nor U10475 (N_10475,N_9223,N_8077);
or U10476 (N_10476,N_9230,N_9028);
nand U10477 (N_10477,N_9072,N_9484);
nor U10478 (N_10478,N_8743,N_9376);
and U10479 (N_10479,N_9976,N_8245);
nand U10480 (N_10480,N_9676,N_8725);
nand U10481 (N_10481,N_8295,N_9253);
and U10482 (N_10482,N_9247,N_9684);
and U10483 (N_10483,N_8343,N_9266);
or U10484 (N_10484,N_9292,N_9087);
or U10485 (N_10485,N_9373,N_9799);
nor U10486 (N_10486,N_8294,N_8853);
nand U10487 (N_10487,N_8021,N_9938);
and U10488 (N_10488,N_8425,N_9926);
and U10489 (N_10489,N_9443,N_8616);
nand U10490 (N_10490,N_9821,N_9871);
nor U10491 (N_10491,N_8988,N_8282);
xor U10492 (N_10492,N_8791,N_8283);
xnor U10493 (N_10493,N_8780,N_9613);
nor U10494 (N_10494,N_9839,N_8241);
or U10495 (N_10495,N_9139,N_9918);
nand U10496 (N_10496,N_8120,N_8957);
nor U10497 (N_10497,N_8822,N_9290);
and U10498 (N_10498,N_8955,N_9836);
nand U10499 (N_10499,N_9635,N_8795);
and U10500 (N_10500,N_9000,N_8917);
or U10501 (N_10501,N_8941,N_8178);
and U10502 (N_10502,N_9458,N_8666);
and U10503 (N_10503,N_9515,N_8091);
nor U10504 (N_10504,N_9587,N_8698);
or U10505 (N_10505,N_9863,N_9875);
or U10506 (N_10506,N_8867,N_9368);
or U10507 (N_10507,N_8144,N_9842);
nand U10508 (N_10508,N_9392,N_8073);
and U10509 (N_10509,N_8081,N_9768);
xnor U10510 (N_10510,N_9864,N_9112);
and U10511 (N_10511,N_9155,N_9862);
nand U10512 (N_10512,N_8550,N_9716);
or U10513 (N_10513,N_9858,N_9181);
xor U10514 (N_10514,N_9847,N_8551);
nand U10515 (N_10515,N_9226,N_8678);
or U10516 (N_10516,N_8443,N_8239);
nor U10517 (N_10517,N_9968,N_9677);
and U10518 (N_10518,N_9573,N_8420);
nand U10519 (N_10519,N_9925,N_9661);
nand U10520 (N_10520,N_8876,N_8626);
or U10521 (N_10521,N_9754,N_9708);
nor U10522 (N_10522,N_8491,N_9304);
nand U10523 (N_10523,N_9727,N_9563);
and U10524 (N_10524,N_8764,N_9763);
nand U10525 (N_10525,N_8801,N_8293);
xnor U10526 (N_10526,N_9366,N_9081);
nand U10527 (N_10527,N_8879,N_9506);
and U10528 (N_10528,N_8086,N_9552);
nor U10529 (N_10529,N_9627,N_9345);
and U10530 (N_10530,N_8192,N_9868);
nor U10531 (N_10531,N_9177,N_8252);
and U10532 (N_10532,N_8668,N_8379);
xnor U10533 (N_10533,N_8231,N_8521);
and U10534 (N_10534,N_8050,N_9742);
or U10535 (N_10535,N_8334,N_8201);
nand U10536 (N_10536,N_8870,N_9891);
and U10537 (N_10537,N_9448,N_9405);
nor U10538 (N_10538,N_9807,N_9620);
or U10539 (N_10539,N_9265,N_9589);
or U10540 (N_10540,N_9881,N_8592);
nor U10541 (N_10541,N_9970,N_8075);
nand U10542 (N_10542,N_8271,N_9320);
nor U10543 (N_10543,N_9641,N_9877);
and U10544 (N_10544,N_8588,N_9789);
or U10545 (N_10545,N_8532,N_9221);
and U10546 (N_10546,N_9481,N_8422);
nand U10547 (N_10547,N_9427,N_9211);
and U10548 (N_10548,N_8502,N_9811);
and U10549 (N_10549,N_8428,N_9117);
xor U10550 (N_10550,N_8914,N_9855);
nor U10551 (N_10551,N_9623,N_8974);
and U10552 (N_10552,N_9593,N_9248);
nor U10553 (N_10553,N_9167,N_8467);
nor U10554 (N_10554,N_9546,N_8712);
xor U10555 (N_10555,N_9021,N_9340);
nor U10556 (N_10556,N_8885,N_8949);
nor U10557 (N_10557,N_8702,N_8821);
and U10558 (N_10558,N_9203,N_9336);
or U10559 (N_10559,N_8889,N_8675);
and U10560 (N_10560,N_8680,N_9282);
nor U10561 (N_10561,N_9518,N_9219);
and U10562 (N_10562,N_8961,N_8834);
nand U10563 (N_10563,N_9201,N_8108);
nand U10564 (N_10564,N_9707,N_9892);
and U10565 (N_10565,N_8011,N_9461);
and U10566 (N_10566,N_9127,N_8790);
xnor U10567 (N_10567,N_9073,N_9185);
nor U10568 (N_10568,N_8385,N_8028);
nor U10569 (N_10569,N_9946,N_9086);
nand U10570 (N_10570,N_8860,N_8895);
nor U10571 (N_10571,N_8817,N_9648);
and U10572 (N_10572,N_8886,N_9802);
nand U10573 (N_10573,N_8270,N_9872);
and U10574 (N_10574,N_9508,N_8033);
and U10575 (N_10575,N_9369,N_8909);
or U10576 (N_10576,N_8545,N_9592);
nor U10577 (N_10577,N_8638,N_8014);
xnor U10578 (N_10578,N_9746,N_8881);
xor U10579 (N_10579,N_8189,N_8929);
nand U10580 (N_10580,N_9246,N_9904);
nor U10581 (N_10581,N_8255,N_8667);
or U10582 (N_10582,N_9331,N_9348);
nand U10583 (N_10583,N_8984,N_8276);
and U10584 (N_10584,N_8344,N_8066);
and U10585 (N_10585,N_9192,N_9986);
and U10586 (N_10586,N_8220,N_9611);
nand U10587 (N_10587,N_8953,N_9256);
or U10588 (N_10588,N_8131,N_9313);
and U10589 (N_10589,N_8771,N_8913);
or U10590 (N_10590,N_8749,N_8199);
xnor U10591 (N_10591,N_8427,N_9162);
or U10592 (N_10592,N_9433,N_9315);
and U10593 (N_10593,N_8769,N_8848);
and U10594 (N_10594,N_8722,N_9729);
nor U10595 (N_10595,N_9287,N_9557);
or U10596 (N_10596,N_8410,N_9451);
and U10597 (N_10597,N_8495,N_8808);
or U10598 (N_10598,N_9978,N_8695);
or U10599 (N_10599,N_8089,N_8541);
and U10600 (N_10600,N_8960,N_8519);
and U10601 (N_10601,N_8219,N_8478);
nand U10602 (N_10602,N_9857,N_9208);
nand U10603 (N_10603,N_9410,N_8904);
and U10604 (N_10604,N_8275,N_8533);
xnor U10605 (N_10605,N_9607,N_9268);
and U10606 (N_10606,N_8782,N_9944);
nor U10607 (N_10607,N_8465,N_8838);
nor U10608 (N_10608,N_8576,N_8653);
nand U10609 (N_10609,N_9270,N_8723);
xor U10610 (N_10610,N_8937,N_9544);
xnor U10611 (N_10611,N_8048,N_8210);
nor U10612 (N_10612,N_9023,N_8462);
nor U10613 (N_10613,N_8325,N_8845);
and U10614 (N_10614,N_8811,N_9803);
and U10615 (N_10615,N_9766,N_9663);
and U10616 (N_10616,N_8143,N_8681);
or U10617 (N_10617,N_8423,N_8922);
or U10618 (N_10618,N_9330,N_9694);
and U10619 (N_10619,N_8544,N_9617);
nand U10620 (N_10620,N_8964,N_9824);
nand U10621 (N_10621,N_9328,N_9404);
and U10622 (N_10622,N_9955,N_8773);
and U10623 (N_10623,N_8812,N_8718);
nand U10624 (N_10624,N_8246,N_8284);
nor U10625 (N_10625,N_8200,N_8589);
and U10626 (N_10626,N_8840,N_9478);
or U10627 (N_10627,N_8760,N_9352);
and U10628 (N_10628,N_8163,N_8473);
nor U10629 (N_10629,N_9378,N_8024);
or U10630 (N_10630,N_8332,N_8587);
nand U10631 (N_10631,N_9397,N_9121);
and U10632 (N_10632,N_8676,N_8035);
nor U10633 (N_10633,N_9621,N_8950);
or U10634 (N_10634,N_8670,N_9685);
nand U10635 (N_10635,N_9471,N_9900);
nand U10636 (N_10636,N_8645,N_8064);
and U10637 (N_10637,N_8858,N_8292);
nand U10638 (N_10638,N_9414,N_8339);
or U10639 (N_10639,N_8538,N_9767);
nor U10640 (N_10640,N_9636,N_9504);
nor U10641 (N_10641,N_8272,N_9917);
and U10642 (N_10642,N_9856,N_9741);
and U10643 (N_10643,N_8721,N_8539);
nor U10644 (N_10644,N_9305,N_9261);
nand U10645 (N_10645,N_9244,N_8128);
or U10646 (N_10646,N_9920,N_8110);
and U10647 (N_10647,N_8682,N_8524);
or U10648 (N_10648,N_9558,N_9537);
xnor U10649 (N_10649,N_9525,N_8222);
nand U10650 (N_10650,N_9704,N_8942);
or U10651 (N_10651,N_8930,N_8902);
nand U10652 (N_10652,N_8401,N_9055);
and U10653 (N_10653,N_9360,N_8337);
or U10654 (N_10654,N_8891,N_9880);
nor U10655 (N_10655,N_9810,N_8152);
nor U10656 (N_10656,N_8326,N_9202);
and U10657 (N_10657,N_9455,N_8575);
and U10658 (N_10658,N_8435,N_9388);
or U10659 (N_10659,N_8092,N_9323);
or U10660 (N_10660,N_9653,N_8045);
and U10661 (N_10661,N_9817,N_8094);
and U10662 (N_10662,N_9937,N_9575);
and U10663 (N_10663,N_8290,N_8796);
or U10664 (N_10664,N_8651,N_9164);
nand U10665 (N_10665,N_8322,N_9294);
and U10666 (N_10666,N_9572,N_8461);
or U10667 (N_10667,N_9601,N_9901);
nand U10668 (N_10668,N_8029,N_9109);
or U10669 (N_10669,N_8777,N_9278);
xor U10670 (N_10670,N_8683,N_8624);
xor U10671 (N_10671,N_9809,N_8311);
nand U10672 (N_10672,N_9111,N_8113);
or U10673 (N_10673,N_8935,N_9783);
nand U10674 (N_10674,N_8417,N_9169);
nand U10675 (N_10675,N_8635,N_9723);
and U10676 (N_10676,N_9476,N_9949);
or U10677 (N_10677,N_8436,N_8350);
nor U10678 (N_10678,N_8500,N_8531);
and U10679 (N_10679,N_8017,N_8377);
xnor U10680 (N_10680,N_8727,N_9054);
or U10681 (N_10681,N_8351,N_8037);
nand U10682 (N_10682,N_9008,N_8880);
nand U10683 (N_10683,N_9234,N_8433);
nor U10684 (N_10684,N_9339,N_9866);
xnor U10685 (N_10685,N_9494,N_8497);
nand U10686 (N_10686,N_8172,N_8068);
xor U10687 (N_10687,N_8485,N_9643);
nor U10688 (N_10688,N_8543,N_9126);
and U10689 (N_10689,N_8378,N_9769);
nor U10690 (N_10690,N_9473,N_8567);
and U10691 (N_10691,N_9665,N_9846);
or U10692 (N_10692,N_9189,N_9134);
nand U10693 (N_10693,N_9157,N_9973);
and U10694 (N_10694,N_9307,N_9159);
or U10695 (N_10695,N_9695,N_9548);
or U10696 (N_10696,N_8584,N_9568);
and U10697 (N_10697,N_8577,N_8096);
and U10698 (N_10698,N_9830,N_8392);
nand U10699 (N_10699,N_9141,N_8730);
nor U10700 (N_10700,N_8312,N_9786);
xnor U10701 (N_10701,N_8117,N_9216);
nor U10702 (N_10702,N_8376,N_9324);
and U10703 (N_10703,N_9277,N_9459);
and U10704 (N_10704,N_9559,N_9638);
nand U10705 (N_10705,N_9183,N_8887);
nand U10706 (N_10706,N_9393,N_8404);
or U10707 (N_10707,N_9389,N_9387);
nor U10708 (N_10708,N_9670,N_9774);
nand U10709 (N_10709,N_8194,N_9516);
and U10710 (N_10710,N_8951,N_9077);
nor U10711 (N_10711,N_8382,N_9210);
nor U10712 (N_10712,N_8959,N_9581);
xnor U10713 (N_10713,N_8819,N_9527);
and U10714 (N_10714,N_8357,N_9319);
nor U10715 (N_10715,N_8818,N_9792);
nor U10716 (N_10716,N_9400,N_9790);
and U10717 (N_10717,N_8602,N_8125);
or U10718 (N_10718,N_9883,N_9032);
nor U10719 (N_10719,N_9934,N_9772);
nand U10720 (N_10720,N_9827,N_9796);
nand U10721 (N_10721,N_8393,N_9982);
nand U10722 (N_10722,N_9194,N_8815);
or U10723 (N_10723,N_8966,N_9179);
nor U10724 (N_10724,N_8250,N_9057);
xor U10725 (N_10725,N_9200,N_8784);
nand U10726 (N_10726,N_9124,N_8861);
nand U10727 (N_10727,N_8257,N_8506);
nor U10728 (N_10728,N_9697,N_9959);
or U10729 (N_10729,N_9782,N_9279);
nor U10730 (N_10730,N_9703,N_9757);
nand U10731 (N_10731,N_9815,N_9220);
and U10732 (N_10732,N_9018,N_9140);
or U10733 (N_10733,N_9106,N_9239);
nor U10734 (N_10734,N_8899,N_8658);
nor U10735 (N_10735,N_8070,N_9801);
or U10736 (N_10736,N_9444,N_9101);
and U10737 (N_10737,N_9914,N_8049);
nand U10738 (N_10738,N_9447,N_8833);
nand U10739 (N_10739,N_9659,N_9565);
nand U10740 (N_10740,N_9399,N_8225);
xnor U10741 (N_10741,N_8931,N_8477);
and U10742 (N_10742,N_8456,N_8656);
and U10743 (N_10743,N_8202,N_8380);
or U10744 (N_10744,N_8969,N_9924);
or U10745 (N_10745,N_9876,N_9724);
nor U10746 (N_10746,N_8155,N_8649);
and U10747 (N_10747,N_9793,N_9151);
nor U10748 (N_10748,N_8774,N_9562);
nand U10749 (N_10749,N_9906,N_8236);
or U10750 (N_10750,N_8100,N_9229);
nand U10751 (N_10751,N_9682,N_8615);
and U10752 (N_10752,N_8079,N_9052);
nand U10753 (N_10753,N_8630,N_9755);
nor U10754 (N_10754,N_8288,N_8857);
nand U10755 (N_10755,N_9604,N_8136);
nor U10756 (N_10756,N_9922,N_8688);
nor U10757 (N_10757,N_9464,N_9851);
or U10758 (N_10758,N_8514,N_8109);
nand U10759 (N_10759,N_8569,N_9556);
and U10760 (N_10760,N_9699,N_9045);
nor U10761 (N_10761,N_9622,N_8327);
and U10762 (N_10762,N_8802,N_9885);
nand U10763 (N_10763,N_9584,N_8494);
nor U10764 (N_10764,N_8517,N_8657);
nand U10765 (N_10765,N_8171,N_8591);
nor U10766 (N_10766,N_8685,N_9272);
nand U10767 (N_10767,N_8400,N_8185);
and U10768 (N_10768,N_8906,N_9353);
nor U10769 (N_10769,N_9062,N_9262);
nor U10770 (N_10770,N_8331,N_9446);
xor U10771 (N_10771,N_8612,N_9854);
nand U10772 (N_10772,N_8260,N_8956);
or U10773 (N_10773,N_9848,N_9255);
or U10774 (N_10774,N_8578,N_8149);
or U10775 (N_10775,N_8530,N_8520);
nor U10776 (N_10776,N_8247,N_9483);
and U10777 (N_10777,N_9009,N_9672);
xnor U10778 (N_10778,N_9217,N_9445);
and U10779 (N_10779,N_9439,N_8429);
nor U10780 (N_10780,N_9138,N_8132);
nor U10781 (N_10781,N_8388,N_9235);
nand U10782 (N_10782,N_8874,N_8355);
xnor U10783 (N_10783,N_9762,N_8614);
or U10784 (N_10784,N_8763,N_8875);
nor U10785 (N_10785,N_8406,N_9577);
nor U10786 (N_10786,N_8659,N_8059);
or U10787 (N_10787,N_8995,N_8797);
nand U10788 (N_10788,N_8669,N_8498);
nor U10789 (N_10789,N_8481,N_9215);
xor U10790 (N_10790,N_8134,N_8556);
or U10791 (N_10791,N_9486,N_9738);
xnor U10792 (N_10792,N_8617,N_9452);
or U10793 (N_10793,N_8620,N_8349);
nor U10794 (N_10794,N_9679,N_9372);
and U10795 (N_10795,N_9258,N_9066);
and U10796 (N_10796,N_8445,N_9726);
or U10797 (N_10797,N_8762,N_9835);
nand U10798 (N_10798,N_8982,N_9582);
nand U10799 (N_10799,N_9429,N_8607);
nor U10800 (N_10800,N_8138,N_8778);
or U10801 (N_10801,N_8925,N_8976);
or U10802 (N_10802,N_9403,N_9994);
nand U10803 (N_10803,N_8069,N_9999);
nor U10804 (N_10804,N_8934,N_9480);
or U10805 (N_10805,N_8085,N_8046);
and U10806 (N_10806,N_9152,N_8217);
or U10807 (N_10807,N_8084,N_8193);
and U10808 (N_10808,N_9083,N_9046);
nand U10809 (N_10809,N_9753,N_9002);
and U10810 (N_10810,N_8195,N_8119);
or U10811 (N_10811,N_8846,N_8992);
or U10812 (N_10812,N_9989,N_9935);
nand U10813 (N_10813,N_9030,N_9632);
or U10814 (N_10814,N_8424,N_8598);
and U10815 (N_10815,N_9869,N_8776);
and U10816 (N_10816,N_8662,N_9667);
nor U10817 (N_10817,N_9004,N_9260);
nand U10818 (N_10818,N_8622,N_9355);
xnor U10819 (N_10819,N_8714,N_8905);
and U10820 (N_10820,N_9719,N_8711);
or U10821 (N_10821,N_8535,N_8565);
nand U10822 (N_10822,N_9967,N_9931);
xor U10823 (N_10823,N_8016,N_8572);
nor U10824 (N_10824,N_8093,N_9241);
nor U10825 (N_10825,N_8728,N_9717);
nand U10826 (N_10826,N_8123,N_8074);
nor U10827 (N_10827,N_8655,N_9146);
or U10828 (N_10828,N_9206,N_9381);
and U10829 (N_10829,N_8403,N_8745);
or U10830 (N_10830,N_8800,N_9011);
nand U10831 (N_10831,N_8854,N_8156);
or U10832 (N_10832,N_8488,N_9472);
nor U10833 (N_10833,N_8285,N_8453);
nand U10834 (N_10834,N_9103,N_9322);
nand U10835 (N_10835,N_9420,N_9496);
nand U10836 (N_10836,N_9675,N_9761);
nor U10837 (N_10837,N_9061,N_9916);
nor U10838 (N_10838,N_8691,N_8673);
and U10839 (N_10839,N_8555,N_9777);
or U10840 (N_10840,N_8947,N_9728);
and U10841 (N_10841,N_9532,N_8253);
nand U10842 (N_10842,N_8549,N_8832);
nor U10843 (N_10843,N_8751,N_8924);
nand U10844 (N_10844,N_9102,N_9421);
nand U10845 (N_10845,N_8775,N_9812);
nand U10846 (N_10846,N_8978,N_8398);
and U10847 (N_10847,N_8945,N_8910);
xnor U10848 (N_10848,N_8242,N_9958);
or U10849 (N_10849,N_9574,N_9744);
nand U10850 (N_10850,N_8650,N_9995);
nand U10851 (N_10851,N_9941,N_8516);
nor U10852 (N_10852,N_8731,N_8618);
nand U10853 (N_10853,N_8390,N_8582);
nor U10854 (N_10854,N_8884,N_8729);
nor U10855 (N_10855,N_8313,N_8692);
or U10856 (N_10856,N_8139,N_8061);
and U10857 (N_10857,N_9251,N_8470);
nand U10858 (N_10858,N_8927,N_8633);
nand U10859 (N_10859,N_8437,N_8896);
and U10860 (N_10860,N_9816,N_8459);
nor U10861 (N_10861,N_8101,N_8705);
or U10862 (N_10862,N_9010,N_9098);
nand U10863 (N_10863,N_8340,N_9291);
or U10864 (N_10864,N_8580,N_8140);
or U10865 (N_10865,N_9543,N_9545);
and U10866 (N_10866,N_8841,N_9800);
or U10867 (N_10867,N_9249,N_9923);
nor U10868 (N_10868,N_9467,N_9466);
xor U10869 (N_10869,N_9142,N_8330);
or U10870 (N_10870,N_9412,N_9867);
xor U10871 (N_10871,N_8186,N_9837);
nor U10872 (N_10872,N_8583,N_9524);
xor U10873 (N_10873,N_8160,N_8460);
or U10874 (N_10874,N_9462,N_8794);
nand U10875 (N_10875,N_9013,N_8563);
nand U10876 (N_10876,N_9634,N_9531);
or U10877 (N_10877,N_8088,N_8362);
or U10878 (N_10878,N_9825,N_9209);
or U10879 (N_10879,N_8105,N_9833);
nand U10880 (N_10880,N_9733,N_9040);
or U10881 (N_10881,N_9108,N_8558);
nor U10882 (N_10882,N_8998,N_9859);
and U10883 (N_10883,N_8067,N_9981);
nor U10884 (N_10884,N_9213,N_9153);
or U10885 (N_10885,N_8063,N_8919);
and U10886 (N_10886,N_9689,N_9110);
and U10887 (N_10887,N_9688,N_8733);
nand U10888 (N_10888,N_8314,N_9350);
and U10889 (N_10889,N_9024,N_9115);
nor U10890 (N_10890,N_9534,N_9712);
or U10891 (N_10891,N_8165,N_9091);
nor U10892 (N_10892,N_8856,N_8696);
nor U10893 (N_10893,N_8828,N_9214);
nand U10894 (N_10894,N_9037,N_8489);
or U10895 (N_10895,N_8256,N_9390);
and U10896 (N_10896,N_9696,N_8258);
nand U10897 (N_10897,N_8789,N_9434);
nor U10898 (N_10898,N_9678,N_8032);
or U10899 (N_10899,N_9058,N_9521);
xnor U10900 (N_10900,N_9765,N_9567);
nor U10901 (N_10901,N_8416,N_8099);
or U10902 (N_10902,N_8414,N_8479);
or U10903 (N_10903,N_9714,N_8962);
nor U10904 (N_10904,N_8989,N_9498);
nand U10905 (N_10905,N_8205,N_9936);
and U10906 (N_10906,N_9539,N_9122);
nand U10907 (N_10907,N_9850,N_9992);
nor U10908 (N_10908,N_9332,N_8309);
or U10909 (N_10909,N_9579,N_8686);
and U10910 (N_10910,N_8412,N_8754);
nor U10911 (N_10911,N_8719,N_9669);
xnor U10912 (N_10912,N_8469,N_9364);
xnor U10913 (N_10913,N_8044,N_9300);
or U10914 (N_10914,N_9079,N_8248);
and U10915 (N_10915,N_9490,N_8997);
nor U10916 (N_10916,N_8316,N_8738);
or U10917 (N_10917,N_9205,N_8038);
nand U10918 (N_10918,N_9734,N_8336);
nand U10919 (N_10919,N_8102,N_8452);
and U10920 (N_10920,N_8823,N_8321);
nor U10921 (N_10921,N_9259,N_8298);
and U10922 (N_10922,N_8009,N_8700);
nor U10923 (N_10923,N_9034,N_8918);
xnor U10924 (N_10924,N_9147,N_8438);
and U10925 (N_10925,N_8076,N_8877);
and U10926 (N_10926,N_9468,N_8996);
and U10927 (N_10927,N_8788,N_9341);
or U10928 (N_10928,N_9354,N_8097);
xnor U10929 (N_10929,N_9067,N_8052);
xor U10930 (N_10930,N_8792,N_9940);
or U10931 (N_10931,N_9781,N_9335);
or U10932 (N_10932,N_9503,N_9626);
or U10933 (N_10933,N_8803,N_8278);
or U10934 (N_10934,N_8368,N_9519);
or U10935 (N_10935,N_9603,N_9911);
or U10936 (N_10936,N_8051,N_8306);
xor U10937 (N_10937,N_8228,N_9977);
or U10938 (N_10938,N_8335,N_9267);
xor U10939 (N_10939,N_8263,N_8027);
nor U10940 (N_10940,N_8636,N_8703);
nor U10941 (N_10941,N_9560,N_8137);
nand U10942 (N_10942,N_9051,N_9064);
or U10943 (N_10943,N_8274,N_9599);
or U10944 (N_10944,N_8315,N_9198);
nand U10945 (N_10945,N_8552,N_8878);
nor U10946 (N_10946,N_8328,N_9085);
or U10947 (N_10947,N_9818,N_9658);
or U10948 (N_10948,N_9569,N_8356);
nor U10949 (N_10949,N_9687,N_9610);
or U10950 (N_10950,N_9651,N_8251);
and U10951 (N_10951,N_8402,N_9980);
nor U10952 (N_10952,N_8975,N_9254);
nor U10953 (N_10953,N_9477,N_8304);
or U10954 (N_10954,N_9637,N_9114);
and U10955 (N_10955,N_9586,N_8266);
and U10956 (N_10956,N_8654,N_8862);
or U10957 (N_10957,N_8528,N_9245);
nand U10958 (N_10958,N_9099,N_9882);
nor U10959 (N_10959,N_8159,N_9664);
nor U10960 (N_10960,N_8184,N_9391);
nand U10961 (N_10961,N_9893,N_8767);
nor U10962 (N_10962,N_9001,N_9176);
and U10963 (N_10963,N_9463,N_8240);
nor U10964 (N_10964,N_8114,N_8677);
xnor U10965 (N_10965,N_9683,N_8907);
nor U10966 (N_10966,N_8367,N_9097);
or U10967 (N_10967,N_9125,N_9731);
or U10968 (N_10968,N_8786,N_8474);
or U10969 (N_10969,N_8542,N_8365);
nand U10970 (N_10970,N_9190,N_9080);
or U10971 (N_10971,N_9426,N_8181);
nor U10972 (N_10972,N_9289,N_8629);
or U10973 (N_10973,N_9383,N_8515);
nand U10974 (N_10974,N_8358,N_8609);
nor U10975 (N_10975,N_8112,N_9070);
nor U10976 (N_10976,N_8162,N_9033);
nand U10977 (N_10977,N_8600,N_9985);
or U10978 (N_10978,N_8267,N_9363);
or U10979 (N_10979,N_9465,N_8432);
and U10980 (N_10980,N_8590,N_8586);
nand U10981 (N_10981,N_8697,N_9713);
nand U10982 (N_10982,N_9418,N_8415);
or U10983 (N_10983,N_8207,N_8409);
nor U10984 (N_10984,N_8233,N_9538);
nand U10985 (N_10985,N_8374,N_8342);
and U10986 (N_10986,N_9631,N_9084);
and U10987 (N_10987,N_9720,N_8227);
nand U10988 (N_10988,N_9852,N_8525);
nand U10989 (N_10989,N_9441,N_9417);
or U10990 (N_10990,N_9945,N_8699);
nor U10991 (N_10991,N_8007,N_8529);
and U10992 (N_10992,N_9910,N_9406);
nand U10993 (N_10993,N_9026,N_8072);
nor U10994 (N_10994,N_8301,N_8187);
and U10995 (N_10995,N_8264,N_9649);
or U10996 (N_10996,N_9764,N_8426);
nor U10997 (N_10997,N_9199,N_8672);
and U10998 (N_10998,N_8299,N_8916);
nor U10999 (N_10999,N_8619,N_9227);
and U11000 (N_11000,N_9888,N_9126);
nand U11001 (N_11001,N_9194,N_9238);
nand U11002 (N_11002,N_9401,N_8158);
or U11003 (N_11003,N_9974,N_8458);
nand U11004 (N_11004,N_9218,N_9905);
and U11005 (N_11005,N_9556,N_9684);
nand U11006 (N_11006,N_9300,N_8883);
and U11007 (N_11007,N_9423,N_8523);
nor U11008 (N_11008,N_9009,N_9378);
nand U11009 (N_11009,N_8320,N_8544);
or U11010 (N_11010,N_9953,N_8556);
nand U11011 (N_11011,N_8140,N_8615);
and U11012 (N_11012,N_8926,N_8528);
nor U11013 (N_11013,N_8698,N_9624);
nand U11014 (N_11014,N_8705,N_9462);
nand U11015 (N_11015,N_8396,N_8535);
or U11016 (N_11016,N_9686,N_9721);
nand U11017 (N_11017,N_8545,N_8041);
and U11018 (N_11018,N_8988,N_8787);
nor U11019 (N_11019,N_9207,N_9318);
nand U11020 (N_11020,N_8356,N_9535);
nor U11021 (N_11021,N_9185,N_8699);
nor U11022 (N_11022,N_8670,N_8037);
or U11023 (N_11023,N_8615,N_8961);
nor U11024 (N_11024,N_8424,N_8619);
nor U11025 (N_11025,N_8469,N_9426);
nor U11026 (N_11026,N_8441,N_9365);
and U11027 (N_11027,N_8354,N_9540);
and U11028 (N_11028,N_8158,N_9944);
or U11029 (N_11029,N_9567,N_8595);
nand U11030 (N_11030,N_8208,N_8947);
nor U11031 (N_11031,N_8554,N_8881);
and U11032 (N_11032,N_8617,N_8862);
or U11033 (N_11033,N_8122,N_9577);
and U11034 (N_11034,N_8022,N_8111);
xnor U11035 (N_11035,N_9491,N_8210);
or U11036 (N_11036,N_8311,N_8039);
and U11037 (N_11037,N_8306,N_8448);
nor U11038 (N_11038,N_9255,N_8231);
and U11039 (N_11039,N_9143,N_8070);
and U11040 (N_11040,N_8110,N_9238);
or U11041 (N_11041,N_9024,N_9973);
and U11042 (N_11042,N_9336,N_9784);
and U11043 (N_11043,N_8476,N_9830);
and U11044 (N_11044,N_9544,N_8261);
and U11045 (N_11045,N_9904,N_9255);
nor U11046 (N_11046,N_8110,N_9643);
nor U11047 (N_11047,N_9320,N_8716);
nand U11048 (N_11048,N_8245,N_8456);
xor U11049 (N_11049,N_8531,N_8097);
or U11050 (N_11050,N_8624,N_9416);
nor U11051 (N_11051,N_9338,N_8705);
nand U11052 (N_11052,N_9461,N_9512);
and U11053 (N_11053,N_9384,N_9415);
nand U11054 (N_11054,N_8330,N_9532);
or U11055 (N_11055,N_9999,N_9062);
or U11056 (N_11056,N_9953,N_9089);
and U11057 (N_11057,N_8218,N_9427);
xor U11058 (N_11058,N_9248,N_8962);
nor U11059 (N_11059,N_8471,N_8845);
nand U11060 (N_11060,N_9092,N_9667);
nor U11061 (N_11061,N_9261,N_8059);
or U11062 (N_11062,N_8190,N_8682);
and U11063 (N_11063,N_9942,N_9504);
nand U11064 (N_11064,N_9930,N_9469);
xnor U11065 (N_11065,N_8525,N_8615);
nand U11066 (N_11066,N_8578,N_8998);
xor U11067 (N_11067,N_8424,N_9506);
and U11068 (N_11068,N_9544,N_9561);
xnor U11069 (N_11069,N_9967,N_9563);
or U11070 (N_11070,N_8617,N_8711);
nor U11071 (N_11071,N_8395,N_8418);
xnor U11072 (N_11072,N_9194,N_9306);
and U11073 (N_11073,N_9850,N_8213);
nand U11074 (N_11074,N_9018,N_9431);
nor U11075 (N_11075,N_9229,N_8724);
nor U11076 (N_11076,N_8275,N_9682);
and U11077 (N_11077,N_8780,N_9256);
nand U11078 (N_11078,N_9141,N_9737);
nor U11079 (N_11079,N_8908,N_9651);
or U11080 (N_11080,N_8731,N_8457);
xnor U11081 (N_11081,N_8562,N_9227);
and U11082 (N_11082,N_9138,N_9030);
nor U11083 (N_11083,N_9225,N_8085);
nor U11084 (N_11084,N_9667,N_9369);
nand U11085 (N_11085,N_9239,N_9402);
nor U11086 (N_11086,N_9817,N_8710);
xnor U11087 (N_11087,N_8943,N_8155);
nor U11088 (N_11088,N_8642,N_9307);
or U11089 (N_11089,N_8757,N_9611);
and U11090 (N_11090,N_8353,N_9006);
nor U11091 (N_11091,N_8378,N_9078);
nand U11092 (N_11092,N_9526,N_9722);
nand U11093 (N_11093,N_9750,N_9265);
or U11094 (N_11094,N_8483,N_9760);
nor U11095 (N_11095,N_9628,N_9177);
and U11096 (N_11096,N_8806,N_8069);
nand U11097 (N_11097,N_9535,N_9521);
nor U11098 (N_11098,N_9081,N_9532);
or U11099 (N_11099,N_9580,N_8003);
and U11100 (N_11100,N_9784,N_8206);
or U11101 (N_11101,N_9774,N_9059);
xnor U11102 (N_11102,N_9593,N_9390);
or U11103 (N_11103,N_9480,N_9315);
and U11104 (N_11104,N_9326,N_8935);
and U11105 (N_11105,N_8247,N_9672);
or U11106 (N_11106,N_9669,N_8880);
or U11107 (N_11107,N_9277,N_8894);
nand U11108 (N_11108,N_9343,N_9589);
nor U11109 (N_11109,N_8696,N_9219);
xnor U11110 (N_11110,N_8688,N_9962);
nor U11111 (N_11111,N_9035,N_8996);
or U11112 (N_11112,N_9189,N_8360);
nor U11113 (N_11113,N_9243,N_9788);
and U11114 (N_11114,N_9043,N_8803);
and U11115 (N_11115,N_8262,N_8476);
and U11116 (N_11116,N_9084,N_8828);
and U11117 (N_11117,N_8332,N_8754);
nor U11118 (N_11118,N_9400,N_9044);
nor U11119 (N_11119,N_8683,N_9703);
nor U11120 (N_11120,N_8446,N_9351);
nand U11121 (N_11121,N_8403,N_8028);
nand U11122 (N_11122,N_8256,N_8054);
nand U11123 (N_11123,N_8898,N_8966);
nand U11124 (N_11124,N_9163,N_8741);
or U11125 (N_11125,N_8872,N_8960);
nor U11126 (N_11126,N_9980,N_9801);
nor U11127 (N_11127,N_9409,N_8410);
or U11128 (N_11128,N_8786,N_8075);
nand U11129 (N_11129,N_8397,N_8979);
nor U11130 (N_11130,N_8174,N_9007);
nand U11131 (N_11131,N_9252,N_8062);
nor U11132 (N_11132,N_9604,N_9685);
or U11133 (N_11133,N_9424,N_8616);
and U11134 (N_11134,N_9010,N_9758);
nor U11135 (N_11135,N_9824,N_9122);
xor U11136 (N_11136,N_8840,N_8992);
or U11137 (N_11137,N_8258,N_9151);
and U11138 (N_11138,N_9163,N_8775);
and U11139 (N_11139,N_9090,N_9934);
and U11140 (N_11140,N_9139,N_8604);
and U11141 (N_11141,N_8170,N_9600);
or U11142 (N_11142,N_9866,N_8947);
nand U11143 (N_11143,N_8673,N_8682);
or U11144 (N_11144,N_9884,N_8581);
nor U11145 (N_11145,N_9462,N_9912);
xor U11146 (N_11146,N_8542,N_8346);
nor U11147 (N_11147,N_8959,N_8141);
or U11148 (N_11148,N_8381,N_8533);
or U11149 (N_11149,N_8608,N_9501);
nand U11150 (N_11150,N_9859,N_9620);
or U11151 (N_11151,N_9275,N_8176);
or U11152 (N_11152,N_9947,N_8227);
and U11153 (N_11153,N_8797,N_9912);
and U11154 (N_11154,N_8305,N_9171);
or U11155 (N_11155,N_8444,N_8161);
nor U11156 (N_11156,N_8571,N_9256);
nor U11157 (N_11157,N_8878,N_9879);
xor U11158 (N_11158,N_9631,N_9598);
nor U11159 (N_11159,N_9868,N_9021);
nor U11160 (N_11160,N_9635,N_8028);
nor U11161 (N_11161,N_9870,N_8200);
and U11162 (N_11162,N_8857,N_9729);
xnor U11163 (N_11163,N_8982,N_8506);
nor U11164 (N_11164,N_9318,N_8176);
or U11165 (N_11165,N_8580,N_9754);
or U11166 (N_11166,N_8716,N_8510);
or U11167 (N_11167,N_8171,N_9110);
xor U11168 (N_11168,N_9258,N_8641);
xor U11169 (N_11169,N_8362,N_9858);
nand U11170 (N_11170,N_8497,N_8059);
xor U11171 (N_11171,N_9152,N_8686);
and U11172 (N_11172,N_9904,N_9715);
and U11173 (N_11173,N_9854,N_9363);
nor U11174 (N_11174,N_8719,N_9613);
or U11175 (N_11175,N_8496,N_9319);
and U11176 (N_11176,N_8938,N_8031);
or U11177 (N_11177,N_9622,N_9327);
or U11178 (N_11178,N_9666,N_8209);
nor U11179 (N_11179,N_8143,N_8164);
xnor U11180 (N_11180,N_9862,N_9480);
and U11181 (N_11181,N_8112,N_9288);
and U11182 (N_11182,N_9195,N_9056);
nor U11183 (N_11183,N_8516,N_8408);
nor U11184 (N_11184,N_9066,N_8869);
or U11185 (N_11185,N_8216,N_9803);
or U11186 (N_11186,N_9118,N_8640);
or U11187 (N_11187,N_8903,N_8740);
nor U11188 (N_11188,N_8434,N_8987);
or U11189 (N_11189,N_8021,N_8653);
xor U11190 (N_11190,N_8069,N_8900);
and U11191 (N_11191,N_9951,N_8057);
xor U11192 (N_11192,N_9548,N_8962);
and U11193 (N_11193,N_8288,N_9406);
or U11194 (N_11194,N_8990,N_9635);
nor U11195 (N_11195,N_8984,N_8319);
and U11196 (N_11196,N_9402,N_8684);
nor U11197 (N_11197,N_9302,N_8109);
nand U11198 (N_11198,N_9754,N_8721);
and U11199 (N_11199,N_9838,N_9152);
and U11200 (N_11200,N_9650,N_9063);
and U11201 (N_11201,N_9575,N_8333);
nand U11202 (N_11202,N_9177,N_9659);
and U11203 (N_11203,N_9155,N_8898);
and U11204 (N_11204,N_8008,N_8850);
and U11205 (N_11205,N_8419,N_9331);
nand U11206 (N_11206,N_8674,N_9751);
nor U11207 (N_11207,N_9488,N_8195);
and U11208 (N_11208,N_8345,N_9942);
nor U11209 (N_11209,N_8313,N_8277);
xnor U11210 (N_11210,N_9269,N_8032);
nand U11211 (N_11211,N_8907,N_9254);
xnor U11212 (N_11212,N_9104,N_9114);
nand U11213 (N_11213,N_8395,N_9312);
nand U11214 (N_11214,N_8192,N_9693);
or U11215 (N_11215,N_9007,N_9436);
or U11216 (N_11216,N_8027,N_9789);
or U11217 (N_11217,N_9078,N_8298);
or U11218 (N_11218,N_8852,N_8683);
nor U11219 (N_11219,N_9562,N_9139);
nor U11220 (N_11220,N_8400,N_8342);
and U11221 (N_11221,N_8597,N_8901);
nand U11222 (N_11222,N_8005,N_8549);
and U11223 (N_11223,N_9232,N_9610);
xor U11224 (N_11224,N_8931,N_9765);
or U11225 (N_11225,N_8500,N_8026);
nor U11226 (N_11226,N_8366,N_9684);
or U11227 (N_11227,N_9017,N_8949);
nand U11228 (N_11228,N_9201,N_8515);
or U11229 (N_11229,N_8180,N_9033);
and U11230 (N_11230,N_9672,N_9108);
nor U11231 (N_11231,N_9069,N_8696);
xor U11232 (N_11232,N_8904,N_9626);
nand U11233 (N_11233,N_9669,N_9805);
xor U11234 (N_11234,N_9797,N_8401);
or U11235 (N_11235,N_8546,N_9673);
or U11236 (N_11236,N_8279,N_8499);
or U11237 (N_11237,N_9809,N_8447);
or U11238 (N_11238,N_8868,N_8127);
or U11239 (N_11239,N_8808,N_8552);
or U11240 (N_11240,N_8644,N_9429);
and U11241 (N_11241,N_8481,N_9498);
nor U11242 (N_11242,N_8551,N_9155);
or U11243 (N_11243,N_8749,N_8461);
nor U11244 (N_11244,N_8233,N_8180);
nor U11245 (N_11245,N_9581,N_8229);
or U11246 (N_11246,N_9163,N_8672);
nand U11247 (N_11247,N_9157,N_9092);
and U11248 (N_11248,N_9915,N_8424);
nor U11249 (N_11249,N_9850,N_8346);
and U11250 (N_11250,N_8610,N_9553);
or U11251 (N_11251,N_9109,N_8318);
or U11252 (N_11252,N_9480,N_9207);
nor U11253 (N_11253,N_8183,N_8286);
or U11254 (N_11254,N_8037,N_8786);
nand U11255 (N_11255,N_9042,N_8683);
xnor U11256 (N_11256,N_9346,N_8680);
nand U11257 (N_11257,N_8008,N_9828);
nor U11258 (N_11258,N_9595,N_8199);
and U11259 (N_11259,N_9323,N_9185);
nor U11260 (N_11260,N_9233,N_8528);
or U11261 (N_11261,N_8047,N_8143);
nor U11262 (N_11262,N_8534,N_9578);
or U11263 (N_11263,N_9412,N_9353);
or U11264 (N_11264,N_8835,N_9125);
or U11265 (N_11265,N_9001,N_8353);
nand U11266 (N_11266,N_9365,N_9993);
nand U11267 (N_11267,N_9078,N_9786);
xor U11268 (N_11268,N_9569,N_9976);
or U11269 (N_11269,N_8869,N_8274);
nor U11270 (N_11270,N_9084,N_8724);
and U11271 (N_11271,N_8558,N_8265);
nor U11272 (N_11272,N_8544,N_8271);
and U11273 (N_11273,N_9435,N_8698);
and U11274 (N_11274,N_8079,N_9013);
and U11275 (N_11275,N_9468,N_9062);
xnor U11276 (N_11276,N_9202,N_8019);
nor U11277 (N_11277,N_8526,N_8070);
and U11278 (N_11278,N_9274,N_9085);
nand U11279 (N_11279,N_9408,N_9363);
nand U11280 (N_11280,N_8830,N_8395);
and U11281 (N_11281,N_8290,N_9810);
nand U11282 (N_11282,N_8808,N_8710);
and U11283 (N_11283,N_8294,N_9432);
xor U11284 (N_11284,N_8054,N_8914);
nor U11285 (N_11285,N_9751,N_8806);
nor U11286 (N_11286,N_8730,N_8382);
nor U11287 (N_11287,N_9346,N_8903);
nor U11288 (N_11288,N_8823,N_9591);
and U11289 (N_11289,N_9788,N_9463);
and U11290 (N_11290,N_8528,N_8369);
and U11291 (N_11291,N_9242,N_9950);
nor U11292 (N_11292,N_8564,N_8088);
nand U11293 (N_11293,N_8426,N_8568);
nand U11294 (N_11294,N_8558,N_9230);
nor U11295 (N_11295,N_9674,N_8176);
nor U11296 (N_11296,N_8514,N_8263);
or U11297 (N_11297,N_9934,N_8688);
or U11298 (N_11298,N_9693,N_9159);
or U11299 (N_11299,N_9024,N_9766);
nand U11300 (N_11300,N_9821,N_9327);
nand U11301 (N_11301,N_8872,N_9863);
nand U11302 (N_11302,N_8321,N_9486);
or U11303 (N_11303,N_9187,N_8095);
nor U11304 (N_11304,N_8270,N_9628);
and U11305 (N_11305,N_8141,N_8633);
and U11306 (N_11306,N_8328,N_9087);
nor U11307 (N_11307,N_9936,N_8410);
or U11308 (N_11308,N_9457,N_9166);
xor U11309 (N_11309,N_8801,N_8915);
nor U11310 (N_11310,N_9714,N_8397);
and U11311 (N_11311,N_9904,N_9685);
nor U11312 (N_11312,N_8809,N_8841);
and U11313 (N_11313,N_9835,N_8331);
or U11314 (N_11314,N_8678,N_9997);
and U11315 (N_11315,N_9294,N_9083);
nor U11316 (N_11316,N_9548,N_9598);
nand U11317 (N_11317,N_9117,N_8997);
or U11318 (N_11318,N_9543,N_9172);
nand U11319 (N_11319,N_8941,N_8310);
xnor U11320 (N_11320,N_8237,N_8002);
nand U11321 (N_11321,N_8069,N_9596);
nor U11322 (N_11322,N_8052,N_8920);
or U11323 (N_11323,N_9223,N_8961);
nand U11324 (N_11324,N_8181,N_8277);
nand U11325 (N_11325,N_8941,N_9685);
or U11326 (N_11326,N_9064,N_9864);
and U11327 (N_11327,N_8001,N_9243);
or U11328 (N_11328,N_9578,N_8824);
or U11329 (N_11329,N_8609,N_9346);
or U11330 (N_11330,N_9757,N_8878);
and U11331 (N_11331,N_9736,N_8571);
nor U11332 (N_11332,N_8145,N_9551);
xor U11333 (N_11333,N_8314,N_8503);
and U11334 (N_11334,N_8195,N_9361);
or U11335 (N_11335,N_8342,N_8198);
nor U11336 (N_11336,N_8907,N_8726);
nor U11337 (N_11337,N_9957,N_9829);
nor U11338 (N_11338,N_8204,N_9930);
and U11339 (N_11339,N_9485,N_9715);
and U11340 (N_11340,N_8167,N_8321);
and U11341 (N_11341,N_8324,N_9778);
or U11342 (N_11342,N_9430,N_9953);
xnor U11343 (N_11343,N_9171,N_8942);
nand U11344 (N_11344,N_8039,N_8307);
or U11345 (N_11345,N_9928,N_9046);
nand U11346 (N_11346,N_9000,N_9515);
and U11347 (N_11347,N_9657,N_9020);
and U11348 (N_11348,N_9480,N_9761);
and U11349 (N_11349,N_9763,N_8059);
and U11350 (N_11350,N_9416,N_8232);
nor U11351 (N_11351,N_8763,N_8068);
or U11352 (N_11352,N_9885,N_9435);
and U11353 (N_11353,N_8713,N_9519);
or U11354 (N_11354,N_8421,N_8876);
nor U11355 (N_11355,N_8242,N_8461);
nor U11356 (N_11356,N_8273,N_8578);
nand U11357 (N_11357,N_9260,N_9114);
xnor U11358 (N_11358,N_9606,N_8769);
xnor U11359 (N_11359,N_8770,N_9291);
and U11360 (N_11360,N_9798,N_8781);
and U11361 (N_11361,N_9396,N_8275);
and U11362 (N_11362,N_8479,N_8659);
nand U11363 (N_11363,N_9692,N_9005);
nor U11364 (N_11364,N_8503,N_9746);
and U11365 (N_11365,N_9989,N_8231);
xor U11366 (N_11366,N_9959,N_8172);
xor U11367 (N_11367,N_8774,N_9256);
nor U11368 (N_11368,N_9193,N_9360);
or U11369 (N_11369,N_8949,N_9294);
and U11370 (N_11370,N_8333,N_8459);
nor U11371 (N_11371,N_9070,N_8332);
nand U11372 (N_11372,N_9278,N_9184);
nand U11373 (N_11373,N_8377,N_9294);
nand U11374 (N_11374,N_9676,N_9735);
nor U11375 (N_11375,N_8622,N_8048);
nand U11376 (N_11376,N_9356,N_9228);
nand U11377 (N_11377,N_8948,N_9772);
nor U11378 (N_11378,N_8017,N_9963);
and U11379 (N_11379,N_8629,N_9898);
or U11380 (N_11380,N_9657,N_9124);
nor U11381 (N_11381,N_9127,N_9938);
and U11382 (N_11382,N_8172,N_8428);
nor U11383 (N_11383,N_9500,N_9540);
or U11384 (N_11384,N_8330,N_8455);
nand U11385 (N_11385,N_8975,N_9036);
xor U11386 (N_11386,N_9018,N_8351);
xnor U11387 (N_11387,N_8438,N_9407);
and U11388 (N_11388,N_8396,N_8080);
nand U11389 (N_11389,N_9263,N_8116);
nand U11390 (N_11390,N_9711,N_9129);
nand U11391 (N_11391,N_9725,N_8164);
or U11392 (N_11392,N_8201,N_9912);
nor U11393 (N_11393,N_9404,N_8146);
and U11394 (N_11394,N_9162,N_9456);
nand U11395 (N_11395,N_8287,N_9625);
or U11396 (N_11396,N_9160,N_9902);
nand U11397 (N_11397,N_9629,N_9452);
and U11398 (N_11398,N_8875,N_9723);
xor U11399 (N_11399,N_9077,N_8229);
and U11400 (N_11400,N_8202,N_8073);
xor U11401 (N_11401,N_9002,N_9008);
or U11402 (N_11402,N_8969,N_9386);
nand U11403 (N_11403,N_9106,N_8570);
or U11404 (N_11404,N_9829,N_9397);
nand U11405 (N_11405,N_8689,N_9531);
nand U11406 (N_11406,N_9607,N_9623);
and U11407 (N_11407,N_8893,N_8524);
and U11408 (N_11408,N_8110,N_8022);
xnor U11409 (N_11409,N_9274,N_8742);
nand U11410 (N_11410,N_8052,N_8196);
nand U11411 (N_11411,N_9175,N_9123);
and U11412 (N_11412,N_9409,N_9025);
and U11413 (N_11413,N_8056,N_9188);
nor U11414 (N_11414,N_9748,N_8919);
and U11415 (N_11415,N_9231,N_9920);
xnor U11416 (N_11416,N_9871,N_9371);
nand U11417 (N_11417,N_8130,N_8666);
or U11418 (N_11418,N_9561,N_9448);
nor U11419 (N_11419,N_8526,N_8958);
and U11420 (N_11420,N_8672,N_9815);
nand U11421 (N_11421,N_8096,N_9337);
nand U11422 (N_11422,N_8656,N_9142);
nor U11423 (N_11423,N_9174,N_8515);
nor U11424 (N_11424,N_9024,N_8765);
or U11425 (N_11425,N_8281,N_8532);
nand U11426 (N_11426,N_9314,N_9755);
or U11427 (N_11427,N_9923,N_8606);
and U11428 (N_11428,N_8685,N_8457);
or U11429 (N_11429,N_8382,N_8603);
or U11430 (N_11430,N_8586,N_8180);
or U11431 (N_11431,N_9865,N_9782);
nor U11432 (N_11432,N_9427,N_9599);
xnor U11433 (N_11433,N_9549,N_9084);
nor U11434 (N_11434,N_8255,N_8642);
nand U11435 (N_11435,N_9522,N_8774);
nand U11436 (N_11436,N_9417,N_9678);
nor U11437 (N_11437,N_9839,N_9626);
xnor U11438 (N_11438,N_9038,N_9659);
and U11439 (N_11439,N_8009,N_8504);
or U11440 (N_11440,N_8622,N_8468);
nand U11441 (N_11441,N_8232,N_8123);
or U11442 (N_11442,N_9019,N_8846);
nor U11443 (N_11443,N_9315,N_9048);
nand U11444 (N_11444,N_9523,N_8157);
nand U11445 (N_11445,N_9963,N_8772);
and U11446 (N_11446,N_9767,N_8608);
nor U11447 (N_11447,N_8508,N_8400);
nand U11448 (N_11448,N_8625,N_9488);
xnor U11449 (N_11449,N_8542,N_8041);
or U11450 (N_11450,N_8789,N_9455);
nand U11451 (N_11451,N_9010,N_8565);
nand U11452 (N_11452,N_9518,N_8755);
or U11453 (N_11453,N_8730,N_9387);
or U11454 (N_11454,N_9729,N_8948);
nand U11455 (N_11455,N_8978,N_9649);
nand U11456 (N_11456,N_8383,N_8535);
nand U11457 (N_11457,N_9272,N_8051);
and U11458 (N_11458,N_9291,N_9431);
nor U11459 (N_11459,N_8251,N_9016);
and U11460 (N_11460,N_9336,N_9950);
nor U11461 (N_11461,N_9286,N_9898);
or U11462 (N_11462,N_8175,N_9225);
or U11463 (N_11463,N_9241,N_8729);
nor U11464 (N_11464,N_9065,N_9692);
or U11465 (N_11465,N_9149,N_9336);
xnor U11466 (N_11466,N_8225,N_9423);
nand U11467 (N_11467,N_8278,N_8344);
nand U11468 (N_11468,N_8097,N_8499);
and U11469 (N_11469,N_9410,N_9653);
nand U11470 (N_11470,N_8698,N_9119);
xor U11471 (N_11471,N_9426,N_8193);
nand U11472 (N_11472,N_9020,N_9488);
xor U11473 (N_11473,N_8596,N_9853);
xor U11474 (N_11474,N_8131,N_8051);
nand U11475 (N_11475,N_8311,N_9212);
or U11476 (N_11476,N_9304,N_8645);
nand U11477 (N_11477,N_9984,N_8544);
nor U11478 (N_11478,N_8082,N_8484);
nor U11479 (N_11479,N_8598,N_8356);
nor U11480 (N_11480,N_8048,N_8196);
nand U11481 (N_11481,N_9401,N_8344);
nor U11482 (N_11482,N_8157,N_9225);
and U11483 (N_11483,N_8047,N_9749);
and U11484 (N_11484,N_8431,N_8206);
and U11485 (N_11485,N_8370,N_8191);
and U11486 (N_11486,N_8027,N_9326);
nor U11487 (N_11487,N_9954,N_9058);
or U11488 (N_11488,N_8911,N_9567);
nand U11489 (N_11489,N_8271,N_8590);
nand U11490 (N_11490,N_8907,N_9349);
or U11491 (N_11491,N_8682,N_9595);
or U11492 (N_11492,N_9245,N_8918);
nor U11493 (N_11493,N_8435,N_8343);
nand U11494 (N_11494,N_8787,N_9245);
nor U11495 (N_11495,N_8188,N_9186);
or U11496 (N_11496,N_9205,N_9156);
or U11497 (N_11497,N_8116,N_9437);
xor U11498 (N_11498,N_9619,N_9643);
nand U11499 (N_11499,N_9899,N_9242);
xnor U11500 (N_11500,N_9508,N_8280);
nand U11501 (N_11501,N_9223,N_9772);
nor U11502 (N_11502,N_8958,N_8374);
nand U11503 (N_11503,N_9224,N_8756);
or U11504 (N_11504,N_9380,N_9756);
or U11505 (N_11505,N_9707,N_8438);
or U11506 (N_11506,N_9075,N_9147);
nand U11507 (N_11507,N_9584,N_8713);
nor U11508 (N_11508,N_9885,N_9197);
nor U11509 (N_11509,N_8116,N_8114);
nor U11510 (N_11510,N_8916,N_8722);
or U11511 (N_11511,N_8357,N_8251);
xor U11512 (N_11512,N_9797,N_8576);
nand U11513 (N_11513,N_8293,N_9615);
nand U11514 (N_11514,N_9288,N_8044);
or U11515 (N_11515,N_8179,N_8100);
xnor U11516 (N_11516,N_8492,N_8572);
xor U11517 (N_11517,N_8427,N_8667);
and U11518 (N_11518,N_9711,N_9997);
nand U11519 (N_11519,N_9523,N_9682);
and U11520 (N_11520,N_9550,N_9945);
nand U11521 (N_11521,N_9034,N_8911);
nand U11522 (N_11522,N_9507,N_9038);
and U11523 (N_11523,N_9609,N_9592);
nor U11524 (N_11524,N_9185,N_8965);
and U11525 (N_11525,N_8745,N_9135);
nand U11526 (N_11526,N_9353,N_8519);
nor U11527 (N_11527,N_9283,N_8442);
xnor U11528 (N_11528,N_8532,N_9912);
nor U11529 (N_11529,N_8181,N_9999);
or U11530 (N_11530,N_8806,N_8852);
and U11531 (N_11531,N_9590,N_9022);
xor U11532 (N_11532,N_9549,N_9846);
nand U11533 (N_11533,N_8294,N_8991);
or U11534 (N_11534,N_9554,N_8555);
nor U11535 (N_11535,N_8318,N_8886);
nor U11536 (N_11536,N_9218,N_8708);
and U11537 (N_11537,N_8540,N_8508);
nor U11538 (N_11538,N_8897,N_9454);
or U11539 (N_11539,N_8198,N_9932);
nand U11540 (N_11540,N_9036,N_9249);
nor U11541 (N_11541,N_8214,N_8073);
nand U11542 (N_11542,N_8971,N_8880);
or U11543 (N_11543,N_9060,N_9970);
xnor U11544 (N_11544,N_8048,N_8188);
xnor U11545 (N_11545,N_8915,N_9388);
nor U11546 (N_11546,N_8417,N_9864);
and U11547 (N_11547,N_9343,N_8785);
xnor U11548 (N_11548,N_9888,N_9481);
and U11549 (N_11549,N_8354,N_8724);
nor U11550 (N_11550,N_9484,N_9938);
or U11551 (N_11551,N_8550,N_8604);
or U11552 (N_11552,N_8738,N_9601);
nand U11553 (N_11553,N_9805,N_9322);
or U11554 (N_11554,N_9464,N_9649);
nand U11555 (N_11555,N_9143,N_8462);
and U11556 (N_11556,N_8221,N_9560);
or U11557 (N_11557,N_9299,N_8682);
nor U11558 (N_11558,N_9499,N_8618);
or U11559 (N_11559,N_8664,N_8147);
nand U11560 (N_11560,N_9514,N_8712);
or U11561 (N_11561,N_8008,N_9696);
nand U11562 (N_11562,N_8200,N_8001);
nand U11563 (N_11563,N_8940,N_9303);
xnor U11564 (N_11564,N_8897,N_9820);
and U11565 (N_11565,N_8333,N_8825);
nand U11566 (N_11566,N_8332,N_9244);
nor U11567 (N_11567,N_9309,N_9630);
nor U11568 (N_11568,N_9837,N_8956);
or U11569 (N_11569,N_9282,N_8537);
nand U11570 (N_11570,N_9827,N_8752);
and U11571 (N_11571,N_9404,N_9243);
and U11572 (N_11572,N_8739,N_9569);
nor U11573 (N_11573,N_8539,N_9981);
nand U11574 (N_11574,N_8023,N_9552);
or U11575 (N_11575,N_9514,N_9977);
xor U11576 (N_11576,N_8110,N_8958);
or U11577 (N_11577,N_8495,N_9046);
and U11578 (N_11578,N_9190,N_9412);
nor U11579 (N_11579,N_8995,N_9524);
or U11580 (N_11580,N_9536,N_8572);
nand U11581 (N_11581,N_9016,N_9543);
nand U11582 (N_11582,N_8332,N_9698);
xnor U11583 (N_11583,N_9483,N_9407);
or U11584 (N_11584,N_8577,N_8038);
xor U11585 (N_11585,N_8353,N_9893);
nand U11586 (N_11586,N_8498,N_8448);
nand U11587 (N_11587,N_9660,N_9586);
and U11588 (N_11588,N_8018,N_9206);
or U11589 (N_11589,N_8973,N_8959);
nor U11590 (N_11590,N_9049,N_8792);
or U11591 (N_11591,N_9222,N_8318);
and U11592 (N_11592,N_8870,N_9536);
nor U11593 (N_11593,N_9196,N_9271);
or U11594 (N_11594,N_8543,N_9363);
nor U11595 (N_11595,N_8268,N_9793);
and U11596 (N_11596,N_9358,N_9146);
nor U11597 (N_11597,N_8685,N_8282);
xnor U11598 (N_11598,N_8452,N_9871);
nand U11599 (N_11599,N_8707,N_8336);
or U11600 (N_11600,N_8925,N_8244);
or U11601 (N_11601,N_8159,N_9307);
nand U11602 (N_11602,N_8150,N_9181);
xor U11603 (N_11603,N_8051,N_8141);
and U11604 (N_11604,N_9764,N_9271);
or U11605 (N_11605,N_9754,N_9809);
or U11606 (N_11606,N_9671,N_8648);
xnor U11607 (N_11607,N_8688,N_9659);
nand U11608 (N_11608,N_8923,N_9344);
or U11609 (N_11609,N_9164,N_9754);
xor U11610 (N_11610,N_9699,N_8779);
nor U11611 (N_11611,N_9936,N_9010);
nor U11612 (N_11612,N_9488,N_9404);
or U11613 (N_11613,N_9427,N_9865);
and U11614 (N_11614,N_9410,N_8184);
xnor U11615 (N_11615,N_8075,N_9381);
and U11616 (N_11616,N_8991,N_9575);
nand U11617 (N_11617,N_9714,N_8577);
or U11618 (N_11618,N_8125,N_8454);
nand U11619 (N_11619,N_8017,N_8601);
or U11620 (N_11620,N_8273,N_9202);
and U11621 (N_11621,N_9556,N_9722);
nor U11622 (N_11622,N_8017,N_8950);
and U11623 (N_11623,N_8781,N_8941);
or U11624 (N_11624,N_9507,N_8110);
nand U11625 (N_11625,N_9823,N_9478);
and U11626 (N_11626,N_9525,N_8025);
and U11627 (N_11627,N_9329,N_9846);
or U11628 (N_11628,N_8183,N_8641);
nand U11629 (N_11629,N_9237,N_8043);
nand U11630 (N_11630,N_9958,N_9237);
and U11631 (N_11631,N_8610,N_8222);
nand U11632 (N_11632,N_8394,N_9569);
or U11633 (N_11633,N_8356,N_9826);
nand U11634 (N_11634,N_9537,N_9653);
or U11635 (N_11635,N_8830,N_8022);
or U11636 (N_11636,N_9861,N_8946);
and U11637 (N_11637,N_8942,N_8364);
nand U11638 (N_11638,N_8839,N_8873);
nor U11639 (N_11639,N_9632,N_9576);
xnor U11640 (N_11640,N_8031,N_9455);
or U11641 (N_11641,N_8766,N_9355);
nor U11642 (N_11642,N_9750,N_8070);
or U11643 (N_11643,N_9189,N_9734);
nand U11644 (N_11644,N_8174,N_9469);
nor U11645 (N_11645,N_8238,N_9454);
nand U11646 (N_11646,N_9949,N_8738);
nor U11647 (N_11647,N_8166,N_9815);
nand U11648 (N_11648,N_8614,N_9188);
xor U11649 (N_11649,N_9407,N_9089);
and U11650 (N_11650,N_9935,N_9279);
nand U11651 (N_11651,N_9163,N_8223);
or U11652 (N_11652,N_8187,N_8510);
nand U11653 (N_11653,N_8583,N_8994);
or U11654 (N_11654,N_9618,N_8997);
nor U11655 (N_11655,N_8947,N_9428);
or U11656 (N_11656,N_9118,N_8365);
nand U11657 (N_11657,N_9723,N_9003);
nor U11658 (N_11658,N_8887,N_8373);
or U11659 (N_11659,N_8936,N_9471);
xnor U11660 (N_11660,N_9592,N_8677);
or U11661 (N_11661,N_9941,N_8948);
nor U11662 (N_11662,N_8283,N_9730);
and U11663 (N_11663,N_9742,N_9189);
nor U11664 (N_11664,N_9254,N_8357);
or U11665 (N_11665,N_8354,N_8214);
xor U11666 (N_11666,N_9217,N_9097);
nand U11667 (N_11667,N_9009,N_8495);
and U11668 (N_11668,N_8967,N_8636);
and U11669 (N_11669,N_8670,N_9691);
nand U11670 (N_11670,N_9939,N_8800);
and U11671 (N_11671,N_9011,N_8636);
nand U11672 (N_11672,N_9618,N_8639);
nor U11673 (N_11673,N_9066,N_8895);
nand U11674 (N_11674,N_8832,N_9859);
nand U11675 (N_11675,N_8839,N_8753);
and U11676 (N_11676,N_8348,N_8229);
and U11677 (N_11677,N_9767,N_8431);
or U11678 (N_11678,N_9059,N_9024);
and U11679 (N_11679,N_9668,N_9796);
nor U11680 (N_11680,N_9566,N_8331);
nand U11681 (N_11681,N_8060,N_9622);
nor U11682 (N_11682,N_8631,N_9261);
and U11683 (N_11683,N_8275,N_9310);
nor U11684 (N_11684,N_8459,N_8864);
xor U11685 (N_11685,N_9836,N_9093);
nand U11686 (N_11686,N_9080,N_8980);
or U11687 (N_11687,N_8430,N_9257);
and U11688 (N_11688,N_9027,N_8989);
and U11689 (N_11689,N_9421,N_9474);
nor U11690 (N_11690,N_9741,N_8193);
or U11691 (N_11691,N_9608,N_8039);
or U11692 (N_11692,N_9991,N_9360);
and U11693 (N_11693,N_8399,N_8755);
and U11694 (N_11694,N_8275,N_8093);
nand U11695 (N_11695,N_9690,N_9313);
nor U11696 (N_11696,N_9686,N_9947);
nand U11697 (N_11697,N_8624,N_8369);
nor U11698 (N_11698,N_8898,N_9222);
nor U11699 (N_11699,N_8331,N_9596);
nor U11700 (N_11700,N_9202,N_9652);
and U11701 (N_11701,N_9741,N_8758);
or U11702 (N_11702,N_9665,N_8659);
or U11703 (N_11703,N_9726,N_9713);
and U11704 (N_11704,N_9505,N_9279);
nand U11705 (N_11705,N_9641,N_8690);
nor U11706 (N_11706,N_9903,N_9948);
nand U11707 (N_11707,N_9349,N_8846);
or U11708 (N_11708,N_8780,N_9185);
and U11709 (N_11709,N_8072,N_8088);
and U11710 (N_11710,N_9961,N_8010);
or U11711 (N_11711,N_8277,N_8678);
nor U11712 (N_11712,N_9489,N_8805);
xnor U11713 (N_11713,N_9389,N_8752);
nand U11714 (N_11714,N_8409,N_8237);
nor U11715 (N_11715,N_9869,N_9988);
nand U11716 (N_11716,N_9440,N_9307);
nand U11717 (N_11717,N_8092,N_8785);
or U11718 (N_11718,N_8768,N_8569);
nand U11719 (N_11719,N_9583,N_9579);
and U11720 (N_11720,N_8201,N_9173);
nor U11721 (N_11721,N_9987,N_8443);
or U11722 (N_11722,N_8682,N_9091);
xnor U11723 (N_11723,N_8880,N_9007);
nor U11724 (N_11724,N_8812,N_8050);
and U11725 (N_11725,N_9489,N_9571);
or U11726 (N_11726,N_9727,N_8770);
nand U11727 (N_11727,N_9553,N_9820);
nor U11728 (N_11728,N_9004,N_9987);
nand U11729 (N_11729,N_8515,N_9870);
and U11730 (N_11730,N_8691,N_8203);
nor U11731 (N_11731,N_9087,N_8320);
nand U11732 (N_11732,N_9708,N_9023);
nor U11733 (N_11733,N_9629,N_9946);
nand U11734 (N_11734,N_8667,N_8097);
nor U11735 (N_11735,N_8918,N_9526);
or U11736 (N_11736,N_8723,N_8835);
nand U11737 (N_11737,N_9340,N_9409);
nor U11738 (N_11738,N_8500,N_8985);
nand U11739 (N_11739,N_8691,N_9577);
or U11740 (N_11740,N_9549,N_8744);
or U11741 (N_11741,N_9642,N_9494);
nor U11742 (N_11742,N_9658,N_8456);
nor U11743 (N_11743,N_8686,N_9174);
nand U11744 (N_11744,N_9417,N_9379);
nand U11745 (N_11745,N_8549,N_8231);
and U11746 (N_11746,N_9846,N_9938);
xnor U11747 (N_11747,N_8802,N_9132);
nand U11748 (N_11748,N_8345,N_9844);
or U11749 (N_11749,N_9681,N_8165);
xor U11750 (N_11750,N_8452,N_9298);
or U11751 (N_11751,N_9188,N_9385);
nor U11752 (N_11752,N_8561,N_8667);
nand U11753 (N_11753,N_8996,N_8521);
nor U11754 (N_11754,N_9850,N_8979);
and U11755 (N_11755,N_9772,N_9080);
nand U11756 (N_11756,N_8429,N_9990);
nor U11757 (N_11757,N_8843,N_9381);
nor U11758 (N_11758,N_8705,N_8960);
nand U11759 (N_11759,N_9379,N_8234);
or U11760 (N_11760,N_8841,N_8548);
nor U11761 (N_11761,N_9472,N_9900);
and U11762 (N_11762,N_8121,N_9755);
or U11763 (N_11763,N_8166,N_9784);
or U11764 (N_11764,N_9027,N_9533);
nor U11765 (N_11765,N_9350,N_9569);
nor U11766 (N_11766,N_8616,N_9235);
nand U11767 (N_11767,N_8524,N_8067);
nand U11768 (N_11768,N_9800,N_9095);
and U11769 (N_11769,N_9751,N_9257);
nor U11770 (N_11770,N_8257,N_9473);
and U11771 (N_11771,N_8437,N_8171);
and U11772 (N_11772,N_8195,N_9026);
xor U11773 (N_11773,N_9992,N_9190);
nor U11774 (N_11774,N_8970,N_8828);
nor U11775 (N_11775,N_8884,N_8540);
xnor U11776 (N_11776,N_9733,N_8128);
and U11777 (N_11777,N_9821,N_8098);
and U11778 (N_11778,N_9648,N_9001);
nand U11779 (N_11779,N_8798,N_8048);
or U11780 (N_11780,N_8452,N_9332);
and U11781 (N_11781,N_9186,N_8568);
nand U11782 (N_11782,N_9889,N_8339);
or U11783 (N_11783,N_9355,N_8660);
or U11784 (N_11784,N_9960,N_9868);
nor U11785 (N_11785,N_9093,N_9783);
and U11786 (N_11786,N_9578,N_8354);
nand U11787 (N_11787,N_9184,N_9600);
nor U11788 (N_11788,N_8876,N_9948);
and U11789 (N_11789,N_9468,N_9743);
nand U11790 (N_11790,N_8911,N_9400);
or U11791 (N_11791,N_9086,N_8632);
nand U11792 (N_11792,N_8793,N_9170);
and U11793 (N_11793,N_9490,N_9359);
or U11794 (N_11794,N_9131,N_9392);
nand U11795 (N_11795,N_8798,N_9471);
or U11796 (N_11796,N_8568,N_9581);
and U11797 (N_11797,N_8090,N_9613);
or U11798 (N_11798,N_9853,N_9324);
nor U11799 (N_11799,N_9955,N_8996);
xor U11800 (N_11800,N_8264,N_8984);
nand U11801 (N_11801,N_8979,N_8991);
xnor U11802 (N_11802,N_9663,N_8507);
nand U11803 (N_11803,N_8157,N_9496);
nor U11804 (N_11804,N_9702,N_9242);
and U11805 (N_11805,N_8709,N_8088);
and U11806 (N_11806,N_8272,N_8198);
or U11807 (N_11807,N_9497,N_9256);
and U11808 (N_11808,N_9124,N_8768);
and U11809 (N_11809,N_8580,N_9609);
nor U11810 (N_11810,N_8363,N_8314);
and U11811 (N_11811,N_8521,N_9572);
nor U11812 (N_11812,N_8662,N_8446);
and U11813 (N_11813,N_9148,N_8437);
and U11814 (N_11814,N_8341,N_8935);
and U11815 (N_11815,N_9556,N_8349);
nor U11816 (N_11816,N_8255,N_9694);
or U11817 (N_11817,N_8643,N_9798);
and U11818 (N_11818,N_9538,N_8888);
nor U11819 (N_11819,N_8735,N_9430);
nand U11820 (N_11820,N_8758,N_9781);
or U11821 (N_11821,N_8473,N_8608);
xor U11822 (N_11822,N_8668,N_8500);
nor U11823 (N_11823,N_9157,N_8316);
and U11824 (N_11824,N_8351,N_9408);
and U11825 (N_11825,N_9230,N_8065);
nand U11826 (N_11826,N_9985,N_8493);
xor U11827 (N_11827,N_8711,N_9621);
or U11828 (N_11828,N_9378,N_9545);
nand U11829 (N_11829,N_8085,N_9630);
or U11830 (N_11830,N_9718,N_9196);
or U11831 (N_11831,N_8401,N_9506);
and U11832 (N_11832,N_9822,N_8415);
xnor U11833 (N_11833,N_9032,N_8267);
or U11834 (N_11834,N_9825,N_8551);
or U11835 (N_11835,N_9527,N_9148);
or U11836 (N_11836,N_9613,N_8894);
and U11837 (N_11837,N_8324,N_8889);
xor U11838 (N_11838,N_9340,N_8357);
and U11839 (N_11839,N_9887,N_8335);
nor U11840 (N_11840,N_9369,N_8156);
nor U11841 (N_11841,N_8478,N_9356);
xor U11842 (N_11842,N_8068,N_8259);
nor U11843 (N_11843,N_8625,N_9628);
xor U11844 (N_11844,N_8536,N_9214);
nor U11845 (N_11845,N_9477,N_9179);
or U11846 (N_11846,N_8527,N_9620);
xnor U11847 (N_11847,N_8741,N_8023);
and U11848 (N_11848,N_9458,N_8885);
xnor U11849 (N_11849,N_9260,N_8456);
xnor U11850 (N_11850,N_8768,N_8909);
or U11851 (N_11851,N_9785,N_9791);
or U11852 (N_11852,N_8403,N_9165);
nor U11853 (N_11853,N_8533,N_8934);
and U11854 (N_11854,N_8255,N_9000);
or U11855 (N_11855,N_9336,N_8907);
nor U11856 (N_11856,N_8807,N_8107);
and U11857 (N_11857,N_9812,N_8787);
or U11858 (N_11858,N_8647,N_8541);
or U11859 (N_11859,N_9005,N_9250);
and U11860 (N_11860,N_8170,N_9364);
or U11861 (N_11861,N_9555,N_9846);
nor U11862 (N_11862,N_9204,N_9840);
or U11863 (N_11863,N_9862,N_8101);
nand U11864 (N_11864,N_9061,N_8478);
nand U11865 (N_11865,N_8874,N_9901);
xnor U11866 (N_11866,N_8164,N_8728);
and U11867 (N_11867,N_8047,N_9477);
nor U11868 (N_11868,N_8187,N_8432);
nand U11869 (N_11869,N_8579,N_9085);
and U11870 (N_11870,N_8780,N_8261);
xor U11871 (N_11871,N_8432,N_8003);
or U11872 (N_11872,N_9107,N_8815);
nor U11873 (N_11873,N_9552,N_8225);
nand U11874 (N_11874,N_8753,N_8534);
nor U11875 (N_11875,N_9545,N_9736);
and U11876 (N_11876,N_9560,N_9052);
xnor U11877 (N_11877,N_9285,N_9139);
nor U11878 (N_11878,N_9429,N_8740);
nand U11879 (N_11879,N_9061,N_9465);
nand U11880 (N_11880,N_8276,N_9354);
and U11881 (N_11881,N_8716,N_8413);
nand U11882 (N_11882,N_8139,N_8265);
nor U11883 (N_11883,N_8453,N_9319);
and U11884 (N_11884,N_9811,N_8617);
xor U11885 (N_11885,N_9993,N_9314);
nand U11886 (N_11886,N_9889,N_9490);
nor U11887 (N_11887,N_9372,N_8618);
nand U11888 (N_11888,N_8901,N_8981);
or U11889 (N_11889,N_9377,N_9509);
and U11890 (N_11890,N_9807,N_9933);
nor U11891 (N_11891,N_8098,N_8076);
and U11892 (N_11892,N_8299,N_8691);
nor U11893 (N_11893,N_9899,N_9821);
nor U11894 (N_11894,N_9969,N_9911);
nor U11895 (N_11895,N_9871,N_8475);
or U11896 (N_11896,N_9609,N_9437);
and U11897 (N_11897,N_9374,N_9065);
or U11898 (N_11898,N_9032,N_9831);
nor U11899 (N_11899,N_8818,N_8621);
nand U11900 (N_11900,N_8027,N_8065);
and U11901 (N_11901,N_8862,N_8751);
xor U11902 (N_11902,N_9261,N_8978);
and U11903 (N_11903,N_8884,N_9850);
nor U11904 (N_11904,N_8622,N_9704);
nor U11905 (N_11905,N_9070,N_9664);
or U11906 (N_11906,N_9019,N_9732);
nor U11907 (N_11907,N_8678,N_8252);
and U11908 (N_11908,N_8787,N_8743);
or U11909 (N_11909,N_8434,N_8904);
and U11910 (N_11910,N_9917,N_9183);
and U11911 (N_11911,N_8674,N_9568);
or U11912 (N_11912,N_8160,N_9309);
or U11913 (N_11913,N_9651,N_9531);
xor U11914 (N_11914,N_8128,N_9399);
nor U11915 (N_11915,N_9783,N_8425);
nand U11916 (N_11916,N_9394,N_9224);
and U11917 (N_11917,N_9843,N_8326);
nor U11918 (N_11918,N_9656,N_9323);
xor U11919 (N_11919,N_9004,N_8443);
or U11920 (N_11920,N_8661,N_9157);
xnor U11921 (N_11921,N_8180,N_8676);
or U11922 (N_11922,N_9162,N_8792);
or U11923 (N_11923,N_8174,N_8681);
and U11924 (N_11924,N_8914,N_9447);
nand U11925 (N_11925,N_9534,N_8187);
nor U11926 (N_11926,N_8309,N_8613);
nor U11927 (N_11927,N_8652,N_9851);
nor U11928 (N_11928,N_8595,N_9345);
or U11929 (N_11929,N_8696,N_9903);
xnor U11930 (N_11930,N_9213,N_9765);
or U11931 (N_11931,N_9988,N_9255);
nand U11932 (N_11932,N_9467,N_9752);
or U11933 (N_11933,N_8680,N_8101);
and U11934 (N_11934,N_8113,N_9942);
nand U11935 (N_11935,N_9461,N_8719);
nor U11936 (N_11936,N_8151,N_9789);
xor U11937 (N_11937,N_9753,N_8449);
nand U11938 (N_11938,N_9969,N_9968);
xor U11939 (N_11939,N_9991,N_8185);
and U11940 (N_11940,N_8489,N_8477);
nor U11941 (N_11941,N_8040,N_9652);
xor U11942 (N_11942,N_8496,N_9355);
or U11943 (N_11943,N_9452,N_9354);
nand U11944 (N_11944,N_9968,N_9628);
nor U11945 (N_11945,N_8721,N_8969);
nand U11946 (N_11946,N_8114,N_9134);
and U11947 (N_11947,N_9907,N_8613);
nor U11948 (N_11948,N_9368,N_8059);
nor U11949 (N_11949,N_8157,N_9665);
nand U11950 (N_11950,N_9953,N_8195);
or U11951 (N_11951,N_8814,N_8747);
nor U11952 (N_11952,N_8395,N_8982);
xor U11953 (N_11953,N_8010,N_8812);
or U11954 (N_11954,N_9969,N_8635);
nand U11955 (N_11955,N_9895,N_8504);
or U11956 (N_11956,N_8583,N_9848);
nor U11957 (N_11957,N_9514,N_8951);
and U11958 (N_11958,N_9794,N_8483);
and U11959 (N_11959,N_9104,N_8726);
nand U11960 (N_11960,N_8276,N_8261);
nand U11961 (N_11961,N_9671,N_8691);
xor U11962 (N_11962,N_8592,N_8031);
or U11963 (N_11963,N_8234,N_9047);
nor U11964 (N_11964,N_9123,N_8771);
nor U11965 (N_11965,N_8794,N_8575);
or U11966 (N_11966,N_9169,N_8491);
or U11967 (N_11967,N_8874,N_8826);
nand U11968 (N_11968,N_9573,N_8400);
or U11969 (N_11969,N_8453,N_8870);
nand U11970 (N_11970,N_8387,N_9740);
or U11971 (N_11971,N_8818,N_8718);
and U11972 (N_11972,N_9661,N_8859);
and U11973 (N_11973,N_8714,N_8335);
xnor U11974 (N_11974,N_9429,N_8301);
xnor U11975 (N_11975,N_8746,N_9768);
nor U11976 (N_11976,N_9317,N_9204);
and U11977 (N_11977,N_9435,N_8058);
and U11978 (N_11978,N_8677,N_9171);
or U11979 (N_11979,N_8499,N_8892);
or U11980 (N_11980,N_9204,N_8284);
xnor U11981 (N_11981,N_9758,N_9842);
and U11982 (N_11982,N_8571,N_8941);
nand U11983 (N_11983,N_8871,N_9837);
nand U11984 (N_11984,N_9047,N_8709);
nand U11985 (N_11985,N_9255,N_9720);
nor U11986 (N_11986,N_8084,N_9830);
nor U11987 (N_11987,N_9228,N_8952);
and U11988 (N_11988,N_8010,N_8714);
xnor U11989 (N_11989,N_8891,N_8132);
and U11990 (N_11990,N_8054,N_8393);
nand U11991 (N_11991,N_9617,N_9897);
or U11992 (N_11992,N_8020,N_8281);
xnor U11993 (N_11993,N_9066,N_8375);
and U11994 (N_11994,N_8939,N_9186);
nor U11995 (N_11995,N_9647,N_9690);
nor U11996 (N_11996,N_9340,N_9104);
nor U11997 (N_11997,N_8490,N_8530);
and U11998 (N_11998,N_8876,N_8943);
or U11999 (N_11999,N_9030,N_9986);
xor U12000 (N_12000,N_10114,N_11331);
and U12001 (N_12001,N_10013,N_10941);
nand U12002 (N_12002,N_10936,N_11569);
or U12003 (N_12003,N_11734,N_10319);
and U12004 (N_12004,N_11028,N_10543);
xnor U12005 (N_12005,N_11723,N_10824);
nor U12006 (N_12006,N_11253,N_11902);
nand U12007 (N_12007,N_11947,N_10624);
or U12008 (N_12008,N_11285,N_10009);
and U12009 (N_12009,N_11323,N_11779);
and U12010 (N_12010,N_10580,N_10890);
nand U12011 (N_12011,N_11116,N_10460);
nor U12012 (N_12012,N_11373,N_10225);
and U12013 (N_12013,N_11059,N_11393);
and U12014 (N_12014,N_11615,N_10625);
and U12015 (N_12015,N_11362,N_11913);
nor U12016 (N_12016,N_10370,N_11103);
nor U12017 (N_12017,N_10354,N_11578);
nand U12018 (N_12018,N_11279,N_11290);
and U12019 (N_12019,N_11490,N_10305);
nor U12020 (N_12020,N_11056,N_11080);
nand U12021 (N_12021,N_11260,N_10125);
and U12022 (N_12022,N_11875,N_11602);
or U12023 (N_12023,N_11938,N_10002);
or U12024 (N_12024,N_11223,N_11701);
xnor U12025 (N_12025,N_10011,N_11960);
or U12026 (N_12026,N_11273,N_10537);
and U12027 (N_12027,N_10250,N_11882);
nor U12028 (N_12028,N_11504,N_10791);
nor U12029 (N_12029,N_10016,N_10898);
nor U12030 (N_12030,N_10885,N_10939);
and U12031 (N_12031,N_10818,N_10320);
nor U12032 (N_12032,N_11427,N_11349);
nand U12033 (N_12033,N_10949,N_10375);
nor U12034 (N_12034,N_11567,N_11943);
and U12035 (N_12035,N_11963,N_11942);
nand U12036 (N_12036,N_10028,N_11957);
nand U12037 (N_12037,N_11852,N_11999);
and U12038 (N_12038,N_11948,N_10730);
nand U12039 (N_12039,N_10501,N_10602);
or U12040 (N_12040,N_11842,N_11733);
and U12041 (N_12041,N_11495,N_11257);
nor U12042 (N_12042,N_11980,N_10097);
nor U12043 (N_12043,N_11752,N_11741);
nor U12044 (N_12044,N_11995,N_11453);
and U12045 (N_12045,N_10119,N_10261);
and U12046 (N_12046,N_11841,N_11365);
and U12047 (N_12047,N_11093,N_11621);
or U12048 (N_12048,N_10476,N_11936);
nor U12049 (N_12049,N_10378,N_10411);
xnor U12050 (N_12050,N_11356,N_11193);
nand U12051 (N_12051,N_11929,N_11836);
nor U12052 (N_12052,N_10557,N_10118);
nor U12053 (N_12053,N_10166,N_11659);
nand U12054 (N_12054,N_11039,N_11529);
xnor U12055 (N_12055,N_11809,N_10217);
nand U12056 (N_12056,N_11541,N_10406);
and U12057 (N_12057,N_11689,N_11386);
nand U12058 (N_12058,N_10396,N_11525);
nor U12059 (N_12059,N_10671,N_10470);
nand U12060 (N_12060,N_10259,N_10598);
nand U12061 (N_12061,N_10137,N_10763);
xnor U12062 (N_12062,N_11345,N_10260);
and U12063 (N_12063,N_10752,N_10645);
nand U12064 (N_12064,N_10353,N_10201);
nand U12065 (N_12065,N_11114,N_10915);
and U12066 (N_12066,N_10636,N_10242);
nand U12067 (N_12067,N_11821,N_11755);
nand U12068 (N_12068,N_10697,N_11280);
nor U12069 (N_12069,N_11473,N_10386);
and U12070 (N_12070,N_11790,N_11117);
and U12071 (N_12071,N_11204,N_11289);
nor U12072 (N_12072,N_10427,N_11079);
nor U12073 (N_12073,N_11464,N_10734);
and U12074 (N_12074,N_10569,N_11712);
and U12075 (N_12075,N_11085,N_11441);
or U12076 (N_12076,N_11224,N_11787);
nor U12077 (N_12077,N_10776,N_11819);
nand U12078 (N_12078,N_10819,N_11873);
nor U12079 (N_12079,N_10715,N_10672);
nor U12080 (N_12080,N_11477,N_10960);
nor U12081 (N_12081,N_11596,N_10657);
nor U12082 (N_12082,N_11861,N_10572);
and U12083 (N_12083,N_10177,N_11840);
xnor U12084 (N_12084,N_11683,N_10417);
nor U12085 (N_12085,N_11372,N_10942);
nor U12086 (N_12086,N_10500,N_10079);
xnor U12087 (N_12087,N_11795,N_10879);
nand U12088 (N_12088,N_11951,N_10409);
or U12089 (N_12089,N_11579,N_10803);
and U12090 (N_12090,N_10200,N_11670);
xnor U12091 (N_12091,N_10640,N_10480);
and U12092 (N_12092,N_10967,N_11815);
nand U12093 (N_12093,N_11187,N_11926);
nor U12094 (N_12094,N_10271,N_11876);
or U12095 (N_12095,N_11057,N_10509);
nand U12096 (N_12096,N_11435,N_11968);
nor U12097 (N_12097,N_10920,N_11429);
nand U12098 (N_12098,N_10466,N_10094);
nor U12099 (N_12099,N_10756,N_10506);
xor U12100 (N_12100,N_10683,N_10514);
and U12101 (N_12101,N_10443,N_11493);
or U12102 (N_12102,N_11329,N_10704);
and U12103 (N_12103,N_11250,N_11405);
or U12104 (N_12104,N_11912,N_11737);
and U12105 (N_12105,N_11856,N_11857);
xor U12106 (N_12106,N_10037,N_11715);
nor U12107 (N_12107,N_10815,N_10491);
nand U12108 (N_12108,N_10058,N_10027);
or U12109 (N_12109,N_10451,N_10980);
or U12110 (N_12110,N_11886,N_10767);
nor U12111 (N_12111,N_10799,N_11570);
or U12112 (N_12112,N_10010,N_11169);
or U12113 (N_12113,N_10905,N_11027);
nor U12114 (N_12114,N_10232,N_10168);
and U12115 (N_12115,N_11890,N_11012);
and U12116 (N_12116,N_11837,N_10336);
and U12117 (N_12117,N_10782,N_10038);
nand U12118 (N_12118,N_10800,N_11054);
nor U12119 (N_12119,N_10182,N_11887);
and U12120 (N_12120,N_10264,N_11108);
xnor U12121 (N_12121,N_10877,N_11696);
and U12122 (N_12122,N_10066,N_10104);
or U12123 (N_12123,N_11316,N_11711);
or U12124 (N_12124,N_11480,N_10779);
xnor U12125 (N_12125,N_11959,N_11195);
or U12126 (N_12126,N_10255,N_11051);
or U12127 (N_12127,N_11786,N_11909);
or U12128 (N_12128,N_11687,N_11158);
nor U12129 (N_12129,N_10964,N_10132);
and U12130 (N_12130,N_11443,N_10424);
nor U12131 (N_12131,N_10282,N_11774);
and U12132 (N_12132,N_10280,N_11807);
and U12133 (N_12133,N_11391,N_10662);
and U12134 (N_12134,N_11749,N_10064);
xnor U12135 (N_12135,N_10315,N_11969);
nor U12136 (N_12136,N_11694,N_10031);
or U12137 (N_12137,N_11036,N_11258);
xnor U12138 (N_12138,N_10220,N_10361);
or U12139 (N_12139,N_11921,N_10993);
nand U12140 (N_12140,N_10821,N_11645);
nand U12141 (N_12141,N_11277,N_11679);
nand U12142 (N_12142,N_10895,N_10733);
and U12143 (N_12143,N_11061,N_10758);
and U12144 (N_12144,N_11585,N_11352);
and U12145 (N_12145,N_11680,N_11516);
or U12146 (N_12146,N_10067,N_11282);
nor U12147 (N_12147,N_11798,N_11152);
or U12148 (N_12148,N_10873,N_10971);
xor U12149 (N_12149,N_10918,N_10213);
or U12150 (N_12150,N_10210,N_11165);
nor U12151 (N_12151,N_11469,N_10026);
or U12152 (N_12152,N_10073,N_11151);
nand U12153 (N_12153,N_11467,N_10741);
and U12154 (N_12154,N_10281,N_11869);
or U12155 (N_12155,N_11859,N_10328);
or U12156 (N_12156,N_11436,N_11924);
nor U12157 (N_12157,N_10953,N_11744);
nand U12158 (N_12158,N_10212,N_10444);
and U12159 (N_12159,N_10740,N_11501);
nand U12160 (N_12160,N_10442,N_10035);
and U12161 (N_12161,N_11997,N_11914);
xor U12162 (N_12162,N_11183,N_11139);
and U12163 (N_12163,N_10146,N_10738);
and U12164 (N_12164,N_11376,N_10827);
xor U12165 (N_12165,N_10687,N_10797);
or U12166 (N_12166,N_10087,N_10390);
or U12167 (N_12167,N_11720,N_10348);
and U12168 (N_12168,N_10665,N_10228);
nand U12169 (N_12169,N_11291,N_11633);
or U12170 (N_12170,N_10700,N_11024);
and U12171 (N_12171,N_10193,N_11910);
nand U12172 (N_12172,N_10399,N_11398);
xnor U12173 (N_12173,N_11557,N_11883);
nand U12174 (N_12174,N_10292,N_10528);
nor U12175 (N_12175,N_10224,N_10802);
and U12176 (N_12176,N_10948,N_11911);
nand U12177 (N_12177,N_10136,N_11555);
or U12178 (N_12178,N_11827,N_10601);
nor U12179 (N_12179,N_11472,N_10901);
or U12180 (N_12180,N_10078,N_11377);
nand U12181 (N_12181,N_10681,N_11142);
and U12182 (N_12182,N_11474,N_10830);
nor U12183 (N_12183,N_11483,N_10532);
nor U12184 (N_12184,N_10098,N_10963);
nor U12185 (N_12185,N_11603,N_10731);
nor U12186 (N_12186,N_10892,N_10142);
xnor U12187 (N_12187,N_10436,N_10191);
nor U12188 (N_12188,N_10121,N_11197);
xor U12189 (N_12189,N_10042,N_11903);
and U12190 (N_12190,N_11115,N_11485);
xor U12191 (N_12191,N_10127,N_10973);
and U12192 (N_12192,N_10760,N_11242);
or U12193 (N_12193,N_11239,N_11375);
nand U12194 (N_12194,N_10547,N_11979);
nand U12195 (N_12195,N_10065,N_11574);
and U12196 (N_12196,N_11806,N_10339);
or U12197 (N_12197,N_10732,N_10274);
nor U12198 (N_12198,N_10387,N_11799);
or U12199 (N_12199,N_10600,N_10108);
nand U12200 (N_12200,N_10128,N_10458);
or U12201 (N_12201,N_10710,N_10579);
nand U12202 (N_12202,N_10302,N_10654);
nor U12203 (N_12203,N_10587,N_10908);
nor U12204 (N_12204,N_10440,N_11199);
or U12205 (N_12205,N_10996,N_11706);
and U12206 (N_12206,N_10124,N_10183);
xnor U12207 (N_12207,N_10769,N_11157);
or U12208 (N_12208,N_11496,N_10642);
nand U12209 (N_12209,N_10004,N_11104);
and U12210 (N_12210,N_10817,N_10207);
or U12211 (N_12211,N_10946,N_11425);
or U12212 (N_12212,N_11030,N_10568);
and U12213 (N_12213,N_11818,N_10825);
or U12214 (N_12214,N_10888,N_10268);
and U12215 (N_12215,N_11410,N_10607);
or U12216 (N_12216,N_11845,N_11381);
and U12217 (N_12217,N_11571,N_11267);
or U12218 (N_12218,N_11753,N_10321);
nor U12219 (N_12219,N_11003,N_11272);
nor U12220 (N_12220,N_11964,N_11288);
or U12221 (N_12221,N_10017,N_10858);
xor U12222 (N_12222,N_10916,N_11539);
nand U12223 (N_12223,N_11259,N_10432);
or U12224 (N_12224,N_11090,N_11327);
nor U12225 (N_12225,N_10482,N_10337);
nand U12226 (N_12226,N_10428,N_11904);
or U12227 (N_12227,N_10205,N_10103);
nor U12228 (N_12228,N_10754,N_11017);
nor U12229 (N_12229,N_10795,N_10927);
and U12230 (N_12230,N_10332,N_11828);
or U12231 (N_12231,N_10284,N_11967);
and U12232 (N_12232,N_10403,N_11897);
nor U12233 (N_12233,N_11811,N_11756);
or U12234 (N_12234,N_11109,N_11359);
or U12235 (N_12235,N_10473,N_10839);
or U12236 (N_12236,N_10433,N_11072);
nor U12237 (N_12237,N_11233,N_10614);
nor U12238 (N_12238,N_10024,N_10149);
nand U12239 (N_12239,N_10472,N_11933);
or U12240 (N_12240,N_10707,N_11006);
and U12241 (N_12241,N_11830,N_11363);
and U12242 (N_12242,N_10369,N_10603);
or U12243 (N_12243,N_11048,N_11606);
xor U12244 (N_12244,N_11867,N_10402);
or U12245 (N_12245,N_10021,N_10489);
nor U12246 (N_12246,N_11150,N_11216);
nand U12247 (N_12247,N_11013,N_10604);
nand U12248 (N_12248,N_10430,N_10512);
nor U12249 (N_12249,N_10870,N_10486);
nand U12250 (N_12250,N_10831,N_10069);
nand U12251 (N_12251,N_10163,N_10335);
nand U12252 (N_12252,N_10230,N_11684);
or U12253 (N_12253,N_11793,N_11510);
and U12254 (N_12254,N_10780,N_10517);
and U12255 (N_12255,N_10077,N_10140);
nand U12256 (N_12256,N_10222,N_11099);
xnor U12257 (N_12257,N_10739,N_11452);
or U12258 (N_12258,N_11309,N_10570);
xor U12259 (N_12259,N_10747,N_10750);
or U12260 (N_12260,N_11255,N_11731);
or U12261 (N_12261,N_11294,N_11692);
nand U12262 (N_12262,N_11163,N_11556);
nand U12263 (N_12263,N_10120,N_10711);
or U12264 (N_12264,N_10955,N_10931);
or U12265 (N_12265,N_10900,N_11524);
nand U12266 (N_12266,N_10468,N_10434);
and U12267 (N_12267,N_10566,N_11847);
nor U12268 (N_12268,N_10599,N_11025);
or U12269 (N_12269,N_11804,N_10863);
nor U12270 (N_12270,N_11986,N_11045);
or U12271 (N_12271,N_11052,N_11388);
and U12272 (N_12272,N_11205,N_11401);
nand U12273 (N_12273,N_10195,N_10743);
and U12274 (N_12274,N_11854,N_11851);
xnor U12275 (N_12275,N_11447,N_11387);
nor U12276 (N_12276,N_11584,N_11125);
nor U12277 (N_12277,N_11385,N_11306);
nor U12278 (N_12278,N_11087,N_10666);
nand U12279 (N_12279,N_11984,N_10360);
and U12280 (N_12280,N_10699,N_11860);
nor U12281 (N_12281,N_10634,N_11132);
nor U12282 (N_12282,N_10934,N_10415);
nor U12283 (N_12283,N_10656,N_11635);
or U12284 (N_12284,N_11497,N_10806);
nand U12285 (N_12285,N_10952,N_10513);
or U12286 (N_12286,N_10619,N_11534);
nor U12287 (N_12287,N_10391,N_10596);
or U12288 (N_12288,N_10522,N_11412);
and U12289 (N_12289,N_10032,N_11319);
xnor U12290 (N_12290,N_10223,N_10880);
and U12291 (N_12291,N_10413,N_11838);
xor U12292 (N_12292,N_11714,N_10521);
or U12293 (N_12293,N_10385,N_11620);
nand U12294 (N_12294,N_10446,N_11426);
nand U12295 (N_12295,N_10772,N_11608);
and U12296 (N_12296,N_10194,N_11378);
nand U12297 (N_12297,N_10856,N_11595);
or U12298 (N_12298,N_10994,N_11275);
xor U12299 (N_12299,N_11026,N_11403);
or U12300 (N_12300,N_10325,N_10524);
nand U12301 (N_12301,N_10046,N_11332);
or U12302 (N_12302,N_10499,N_10490);
or U12303 (N_12303,N_10074,N_11976);
or U12304 (N_12304,N_11075,N_11461);
and U12305 (N_12305,N_11666,N_10903);
nor U12306 (N_12306,N_11161,N_11989);
or U12307 (N_12307,N_11225,N_11191);
nor U12308 (N_12308,N_10530,N_11862);
nor U12309 (N_12309,N_10309,N_10133);
nand U12310 (N_12310,N_10093,N_11081);
or U12311 (N_12311,N_10560,N_10254);
xnor U12312 (N_12312,N_11318,N_11287);
nor U12313 (N_12313,N_10310,N_10816);
nor U12314 (N_12314,N_10584,N_10567);
nor U12315 (N_12315,N_10467,N_11777);
nor U12316 (N_12316,N_11783,N_11629);
xnor U12317 (N_12317,N_11126,N_10383);
nand U12318 (N_12318,N_11144,N_10643);
nor U12319 (N_12319,N_10940,N_10812);
nand U12320 (N_12320,N_10419,N_11350);
or U12321 (N_12321,N_11727,N_10979);
nand U12322 (N_12322,N_11624,N_10169);
or U12323 (N_12323,N_10729,N_11507);
and U12324 (N_12324,N_11729,N_10048);
or U12325 (N_12325,N_10622,N_10199);
or U12326 (N_12326,N_11586,N_10494);
nor U12327 (N_12327,N_10068,N_11214);
nand U12328 (N_12328,N_10544,N_11992);
nand U12329 (N_12329,N_11747,N_11983);
nor U12330 (N_12330,N_10976,N_10593);
or U12331 (N_12331,N_10631,N_10454);
and U12332 (N_12332,N_11704,N_11589);
and U12333 (N_12333,N_11797,N_10418);
nor U12334 (N_12334,N_11432,N_11422);
nand U12335 (N_12335,N_10678,N_10868);
and U12336 (N_12336,N_11010,N_11424);
or U12337 (N_12337,N_10836,N_10693);
nand U12338 (N_12338,N_10295,N_11702);
and U12339 (N_12339,N_10652,N_10327);
xnor U12340 (N_12340,N_10926,N_10561);
or U12341 (N_12341,N_10753,N_10331);
nand U12342 (N_12342,N_10041,N_10562);
or U12343 (N_12343,N_11966,N_11245);
nor U12344 (N_12344,N_10841,N_10591);
or U12345 (N_12345,N_11708,N_11721);
nor U12346 (N_12346,N_10096,N_10893);
nand U12347 (N_12347,N_10278,N_11005);
and U12348 (N_12348,N_11935,N_10674);
or U12349 (N_12349,N_10357,N_10236);
and U12350 (N_12350,N_11074,N_11750);
nor U12351 (N_12351,N_10653,N_10809);
nor U12352 (N_12352,N_10366,N_11043);
nor U12353 (N_12353,N_10912,N_11899);
and U12354 (N_12354,N_10275,N_11993);
nand U12355 (N_12355,N_11227,N_10371);
nand U12356 (N_12356,N_11462,N_11945);
nand U12357 (N_12357,N_11654,N_11455);
and U12358 (N_12358,N_11757,N_11949);
nand U12359 (N_12359,N_10368,N_10938);
and U12360 (N_12360,N_11858,N_10243);
or U12361 (N_12361,N_11212,N_10983);
nor U12362 (N_12362,N_10526,N_10350);
and U12363 (N_12363,N_11816,N_10574);
nor U12364 (N_12364,N_11397,N_11977);
and U12365 (N_12365,N_11996,N_10173);
nor U12366 (N_12366,N_11143,N_11665);
nor U12367 (N_12367,N_11725,N_10006);
or U12368 (N_12368,N_11732,N_11409);
and U12369 (N_12369,N_10899,N_10082);
and U12370 (N_12370,N_10762,N_10751);
nand U12371 (N_12371,N_10606,N_11137);
and U12372 (N_12372,N_11210,N_10340);
or U12373 (N_12373,N_11448,N_10478);
or U12374 (N_12374,N_10655,N_11208);
nand U12375 (N_12375,N_10755,N_10714);
nand U12376 (N_12376,N_10857,N_10465);
and U12377 (N_12377,N_11370,N_11008);
xnor U12378 (N_12378,N_10745,N_11658);
nor U12379 (N_12379,N_10055,N_11218);
and U12380 (N_12380,N_10712,N_11179);
or U12381 (N_12381,N_11812,N_10450);
nor U12382 (N_12382,N_10285,N_11893);
xnor U12383 (N_12383,N_11740,N_10582);
and U12384 (N_12384,N_11475,N_10209);
nor U12385 (N_12385,N_10904,N_11759);
nand U12386 (N_12386,N_10464,N_10594);
or U12387 (N_12387,N_11905,N_11874);
xnor U12388 (N_12388,N_11609,N_11825);
or U12389 (N_12389,N_10052,N_11826);
and U12390 (N_12390,N_11270,N_11313);
and U12391 (N_12391,N_11268,N_11791);
or U12392 (N_12392,N_10047,N_11789);
nor U12393 (N_12393,N_10053,N_10477);
xor U12394 (N_12394,N_10105,N_11296);
nor U12395 (N_12395,N_11865,N_10299);
nor U12396 (N_12396,N_11023,N_11685);
nor U12397 (N_12397,N_11358,N_11196);
or U12398 (N_12398,N_11533,N_10637);
or U12399 (N_12399,N_10279,N_11411);
xor U12400 (N_12400,N_10578,N_10054);
and U12401 (N_12401,N_10291,N_11408);
and U12402 (N_12402,N_11062,N_11367);
and U12403 (N_12403,N_10377,N_10644);
nand U12404 (N_12404,N_10043,N_11011);
or U12405 (N_12405,N_11674,N_11123);
nand U12406 (N_12406,N_11746,N_11022);
and U12407 (N_12407,N_11406,N_11961);
nand U12408 (N_12408,N_11042,N_11190);
nor U12409 (N_12409,N_10921,N_10367);
nand U12410 (N_12410,N_11738,N_11389);
or U12411 (N_12411,N_10757,N_11065);
nand U12412 (N_12412,N_10785,N_11597);
or U12413 (N_12413,N_10176,N_11632);
or U12414 (N_12414,N_10688,N_11440);
and U12415 (N_12415,N_10313,N_11465);
and U12416 (N_12416,N_10342,N_10110);
nor U12417 (N_12417,N_11780,N_11077);
and U12418 (N_12418,N_11201,N_10449);
nor U12419 (N_12419,N_11168,N_10889);
or U12420 (N_12420,N_11982,N_11407);
and U12421 (N_12421,N_11040,N_10850);
nand U12422 (N_12422,N_10558,N_10551);
and U12423 (N_12423,N_11050,N_11751);
or U12424 (N_12424,N_10535,N_11972);
nand U12425 (N_12425,N_10376,N_10090);
nor U12426 (N_12426,N_10160,N_10860);
or U12427 (N_12427,N_10958,N_10076);
and U12428 (N_12428,N_11069,N_11127);
nand U12429 (N_12429,N_11593,N_10629);
and U12430 (N_12430,N_10559,N_11298);
or U12431 (N_12431,N_11129,N_10961);
and U12432 (N_12432,N_11623,N_10759);
or U12433 (N_12433,N_11086,N_10420);
xnor U12434 (N_12434,N_10798,N_11559);
xor U12435 (N_12435,N_11044,N_11211);
and U12436 (N_12436,N_11021,N_11653);
or U12437 (N_12437,N_11417,N_11922);
nand U12438 (N_12438,N_10853,N_10188);
and U12439 (N_12439,N_10696,N_11987);
and U12440 (N_12440,N_11229,N_10977);
and U12441 (N_12441,N_11519,N_10667);
or U12442 (N_12442,N_11113,N_11369);
nand U12443 (N_12443,N_11944,N_11335);
nand U12444 (N_12444,N_10917,N_10029);
nor U12445 (N_12445,N_10247,N_11112);
nor U12446 (N_12446,N_10650,N_11324);
and U12447 (N_12447,N_10575,N_11293);
or U12448 (N_12448,N_11975,N_11400);
nand U12449 (N_12449,N_11209,N_11540);
nor U12450 (N_12450,N_11667,N_11889);
nor U12451 (N_12451,N_10749,N_11384);
nor U12452 (N_12452,N_11492,N_11119);
nand U12453 (N_12453,N_11107,N_10106);
and U12454 (N_12454,N_11499,N_10138);
nand U12455 (N_12455,N_10887,N_11908);
or U12456 (N_12456,N_10516,N_11906);
and U12457 (N_12457,N_10364,N_10304);
nand U12458 (N_12458,N_11430,N_11418);
nor U12459 (N_12459,N_10453,N_10075);
nand U12460 (N_12460,N_10982,N_10703);
xor U12461 (N_12461,N_11357,N_11479);
and U12462 (N_12462,N_11064,N_10646);
xor U12463 (N_12463,N_11450,N_11284);
nand U12464 (N_12464,N_11466,N_11100);
and U12465 (N_12465,N_11058,N_11468);
or U12466 (N_12466,N_11060,N_11000);
or U12467 (N_12467,N_10635,N_11764);
nor U12468 (N_12468,N_11299,N_10725);
and U12469 (N_12469,N_11866,N_11256);
or U12470 (N_12470,N_11442,N_10192);
nand U12471 (N_12471,N_10358,N_11135);
nor U12472 (N_12472,N_10153,N_11545);
nand U12473 (N_12473,N_11523,N_11509);
or U12474 (N_12474,N_11552,N_10206);
and U12475 (N_12475,N_11067,N_11678);
or U12476 (N_12476,N_11614,N_10170);
nand U12477 (N_12477,N_11071,N_11928);
and U12478 (N_12478,N_11094,N_10648);
or U12479 (N_12479,N_11326,N_11537);
nor U12480 (N_12480,N_11513,N_11891);
and U12481 (N_12481,N_11394,N_11034);
or U12482 (N_12482,N_11953,N_11834);
nand U12483 (N_12483,N_11251,N_11970);
nand U12484 (N_12484,N_10608,N_10867);
nand U12485 (N_12485,N_10229,N_11894);
nand U12486 (N_12486,N_11153,N_10972);
nor U12487 (N_12487,N_10766,N_10422);
or U12488 (N_12488,N_10832,N_11796);
nand U12489 (N_12489,N_10862,N_10611);
or U12490 (N_12490,N_10245,N_11155);
nor U12491 (N_12491,N_10985,N_11149);
or U12492 (N_12492,N_11124,N_11128);
nand U12493 (N_12493,N_11577,N_10384);
or U12494 (N_12494,N_10437,N_10698);
or U12495 (N_12495,N_11334,N_10553);
xor U12496 (N_12496,N_10523,N_10585);
nand U12497 (N_12497,N_10615,N_10826);
nand U12498 (N_12498,N_11498,N_10684);
or U12499 (N_12499,N_10668,N_11771);
or U12500 (N_12500,N_10719,N_10144);
or U12501 (N_12501,N_10589,N_10095);
or U12502 (N_12502,N_10995,N_11049);
nor U12503 (N_12503,N_11348,N_10115);
and U12504 (N_12504,N_10311,N_10240);
or U12505 (N_12505,N_11146,N_11396);
or U12506 (N_12506,N_10796,N_11337);
nor U12507 (N_12507,N_10515,N_10541);
or U12508 (N_12508,N_11662,N_10333);
or U12509 (N_12509,N_11184,N_11248);
nor U12510 (N_12510,N_11171,N_11974);
nand U12511 (N_12511,N_10117,N_11200);
and U12512 (N_12512,N_10198,N_11705);
or U12513 (N_12513,N_10380,N_11222);
and U12514 (N_12514,N_11220,N_10874);
nor U12515 (N_12515,N_10113,N_10974);
nand U12516 (N_12516,N_10861,N_10702);
or U12517 (N_12517,N_10022,N_11286);
and U12518 (N_12518,N_11344,N_10287);
nand U12519 (N_12519,N_11471,N_11766);
xor U12520 (N_12520,N_11754,N_10063);
and U12521 (N_12521,N_11330,N_11916);
or U12522 (N_12522,N_11527,N_10894);
or U12523 (N_12523,N_10793,N_11767);
xnor U12524 (N_12524,N_11033,N_11843);
and U12525 (N_12525,N_10019,N_11338);
xnor U12526 (N_12526,N_11340,N_11591);
nor U12527 (N_12527,N_11382,N_11283);
or U12528 (N_12528,N_11800,N_10999);
and U12529 (N_12529,N_11550,N_10081);
and U12530 (N_12530,N_11600,N_11743);
xnor U12531 (N_12531,N_10546,N_10141);
xnor U12532 (N_12532,N_10249,N_10033);
nand U12533 (N_12533,N_10875,N_10493);
and U12534 (N_12534,N_10801,N_11677);
xnor U12535 (N_12535,N_11675,N_10677);
nor U12536 (N_12536,N_10778,N_10276);
or U12537 (N_12537,N_11133,N_10876);
and U12538 (N_12538,N_10518,N_11962);
nor U12539 (N_12539,N_10709,N_11181);
or U12540 (N_12540,N_10135,N_10161);
nand U12541 (N_12541,N_10346,N_10408);
or U12542 (N_12542,N_11660,N_10592);
nand U12543 (N_12543,N_11402,N_10429);
or U12544 (N_12544,N_10221,N_11955);
and U12545 (N_12545,N_11106,N_10987);
or U12546 (N_12546,N_10435,N_11568);
or U12547 (N_12547,N_11007,N_11937);
and U12548 (N_12548,N_11985,N_11276);
or U12549 (N_12549,N_11768,N_11794);
nor U12550 (N_12550,N_10246,N_11078);
and U12551 (N_12551,N_10781,N_10761);
nor U12552 (N_12552,N_11551,N_11898);
or U12553 (N_12553,N_11881,N_10507);
nand U12554 (N_12554,N_11952,N_11346);
nand U12555 (N_12555,N_11434,N_11230);
xor U12556 (N_12556,N_11742,N_11354);
and U12557 (N_12557,N_11785,N_11646);
xor U12558 (N_12558,N_10267,N_11231);
or U12559 (N_12559,N_11506,N_11451);
nor U12560 (N_12560,N_11548,N_11445);
or U12561 (N_12561,N_11878,N_11037);
or U12562 (N_12562,N_11526,N_11091);
nor U12563 (N_12563,N_10990,N_10823);
nand U12564 (N_12564,N_11252,N_10717);
nor U12565 (N_12565,N_11301,N_10158);
nor U12566 (N_12566,N_10923,N_11254);
or U12567 (N_12567,N_11032,N_10548);
nor U12568 (N_12568,N_11173,N_11940);
xnor U12569 (N_12569,N_10573,N_10581);
or U12570 (N_12570,N_11649,N_11950);
or U12571 (N_12571,N_11990,N_11489);
nand U12572 (N_12572,N_10187,N_10253);
nand U12573 (N_12573,N_10928,N_10639);
and U12574 (N_12574,N_10937,N_10393);
nor U12575 (N_12575,N_11088,N_10777);
and U12576 (N_12576,N_11131,N_11644);
nor U12577 (N_12577,N_10563,N_11531);
nand U12578 (N_12578,N_10381,N_11604);
nor U12579 (N_12579,N_11719,N_10070);
and U12580 (N_12580,N_10978,N_10211);
and U12581 (N_12581,N_10379,N_10349);
and U12582 (N_12582,N_10112,N_11419);
or U12583 (N_12583,N_11215,N_11651);
or U12584 (N_12584,N_11102,N_10056);
nand U12585 (N_12585,N_11488,N_11300);
nand U12586 (N_12586,N_11808,N_10913);
nand U12587 (N_12587,N_11832,N_10626);
nand U12588 (N_12588,N_10590,N_10620);
and U12589 (N_12589,N_10617,N_11046);
or U12590 (N_12590,N_11542,N_11835);
and U12591 (N_12591,N_10503,N_10421);
xor U12592 (N_12592,N_11941,N_11317);
and U12593 (N_12593,N_10156,N_11110);
and U12594 (N_12594,N_10556,N_10632);
xor U12595 (N_12595,N_10479,N_10265);
nor U12596 (N_12596,N_10510,N_11491);
or U12597 (N_12597,N_11176,N_10618);
and U12598 (N_12598,N_10159,N_10447);
nor U12599 (N_12599,N_11175,N_11848);
and U12600 (N_12600,N_10147,N_11784);
nand U12601 (N_12601,N_10459,N_11460);
xor U12602 (N_12602,N_11872,N_10441);
nand U12603 (N_12603,N_11415,N_10914);
and U12604 (N_12604,N_11892,N_10588);
or U12605 (N_12605,N_10988,N_10283);
nor U12606 (N_12606,N_10944,N_10012);
and U12607 (N_12607,N_11709,N_10215);
or U12608 (N_12608,N_11515,N_11379);
nor U12609 (N_12609,N_10545,N_10045);
nor U12610 (N_12610,N_11844,N_10686);
and U12611 (N_12611,N_10804,N_11770);
or U12612 (N_12612,N_10084,N_11014);
and U12613 (N_12613,N_10998,N_11041);
nor U12614 (N_12614,N_10849,N_10404);
nand U12615 (N_12615,N_11638,N_11657);
nand U12616 (N_12616,N_11138,N_11864);
nor U12617 (N_12617,N_10455,N_10181);
nor U12618 (N_12618,N_10872,N_11295);
xnor U12619 (N_12619,N_10787,N_11713);
xor U12620 (N_12620,N_10986,N_11020);
nor U12621 (N_12621,N_10508,N_11605);
nor U12622 (N_12622,N_11304,N_10484);
nand U12623 (N_12623,N_11228,N_11156);
nand U12624 (N_12624,N_10186,N_10388);
nor U12625 (N_12625,N_11502,N_10813);
xor U12626 (N_12626,N_11971,N_10151);
or U12627 (N_12627,N_10294,N_10527);
nor U12628 (N_12628,N_10431,N_10092);
or U12629 (N_12629,N_10577,N_11601);
or U12630 (N_12630,N_10911,N_10296);
nand U12631 (N_12631,N_11627,N_11178);
or U12632 (N_12632,N_11803,N_11339);
nand U12633 (N_12633,N_11001,N_11676);
nand U12634 (N_12634,N_11167,N_10457);
and U12635 (N_12635,N_10469,N_11002);
nand U12636 (N_12636,N_11722,N_11939);
and U12637 (N_12637,N_10951,N_10519);
nand U12638 (N_12638,N_11120,N_10882);
nand U12639 (N_12639,N_10610,N_11626);
and U12640 (N_12640,N_11244,N_11839);
and U12641 (N_12641,N_10475,N_10638);
or U12642 (N_12642,N_11029,N_11444);
nor U12643 (N_12643,N_10235,N_10126);
nand U12644 (N_12644,N_11583,N_11958);
nand U12645 (N_12645,N_11697,N_10790);
or U12646 (N_12646,N_10298,N_10909);
nand U12647 (N_12647,N_11236,N_10670);
nor U12648 (N_12648,N_10162,N_10794);
xnor U12649 (N_12649,N_10189,N_10204);
nor U12650 (N_12650,N_10723,N_11735);
and U12651 (N_12651,N_10290,N_10925);
or U12652 (N_12652,N_11760,N_10185);
nor U12653 (N_12653,N_10727,N_10001);
nand U12654 (N_12654,N_10647,N_11637);
xor U12655 (N_12655,N_11748,N_10748);
and U12656 (N_12656,N_11122,N_10843);
or U12657 (N_12657,N_11226,N_10462);
and U12658 (N_12658,N_11849,N_11084);
and U12659 (N_12659,N_10613,N_10609);
or U12660 (N_12660,N_10910,N_10184);
or U12661 (N_12661,N_11009,N_11154);
nor U12662 (N_12662,N_10051,N_10695);
nand U12663 (N_12663,N_10190,N_11884);
or U12664 (N_12664,N_11850,N_10992);
or U12665 (N_12665,N_11981,N_11642);
nor U12666 (N_12666,N_11562,N_11333);
or U12667 (N_12667,N_11549,N_10689);
or U12668 (N_12668,N_10906,N_10682);
xor U12669 (N_12669,N_10742,N_10145);
nor U12670 (N_12670,N_10989,N_10030);
or U12671 (N_12671,N_10884,N_10564);
or U12672 (N_12672,N_11763,N_11576);
nand U12673 (N_12673,N_10628,N_10829);
and U12674 (N_12674,N_10784,N_11564);
nand U12675 (N_12675,N_10673,N_10716);
nor U12676 (N_12676,N_10497,N_10765);
xor U12677 (N_12677,N_11765,N_11611);
nand U12678 (N_12678,N_10929,N_11607);
or U12679 (N_12679,N_11581,N_11431);
and U12680 (N_12680,N_10771,N_10023);
or U12681 (N_12681,N_11234,N_11863);
or U12682 (N_12682,N_11068,N_10966);
nand U12683 (N_12683,N_11414,N_10044);
nor U12684 (N_12684,N_10134,N_11416);
nor U12685 (N_12685,N_11145,N_11612);
nor U12686 (N_12686,N_10997,N_10805);
and U12687 (N_12687,N_10091,N_11159);
and U12688 (N_12688,N_11587,N_11035);
or U12689 (N_12689,N_10227,N_10485);
nor U12690 (N_12690,N_10401,N_10736);
and U12691 (N_12691,N_11792,N_10616);
and U12692 (N_12692,N_11308,N_10363);
and U12693 (N_12693,N_10343,N_11558);
nand U12694 (N_12694,N_11217,N_11189);
and U12695 (N_12695,N_10721,N_11917);
and U12696 (N_12696,N_11814,N_11476);
or U12697 (N_12697,N_11055,N_11698);
xnor U12698 (N_12698,N_11089,N_11243);
and U12699 (N_12699,N_10970,N_11776);
xor U12700 (N_12700,N_11802,N_11923);
and U12701 (N_12701,N_11631,N_11508);
and U12702 (N_12702,N_11016,N_11769);
or U12703 (N_12703,N_10015,N_10314);
nand U12704 (N_12704,N_10216,N_10612);
nand U12705 (N_12705,N_10663,N_10293);
or U12706 (N_12706,N_10968,N_10775);
or U12707 (N_12707,N_10538,N_10018);
or U12708 (N_12708,N_10203,N_11946);
nand U12709 (N_12709,N_10595,N_10111);
nand U12710 (N_12710,N_11328,N_10897);
xor U12711 (N_12711,N_11082,N_10174);
and U12712 (N_12712,N_11610,N_10945);
or U12713 (N_12713,N_10452,N_11824);
nor U12714 (N_12714,N_10014,N_10323);
or U12715 (N_12715,N_11213,N_10878);
xnor U12716 (N_12716,N_10359,N_11566);
or U12717 (N_12717,N_11805,N_10416);
nand U12718 (N_12718,N_11901,N_11588);
or U12719 (N_12719,N_11221,N_10902);
nand U12720 (N_12720,N_11521,N_10828);
and U12721 (N_12721,N_10308,N_10175);
nor U12722 (N_12722,N_10398,N_10273);
nor U12723 (N_12723,N_11066,N_11505);
nand U12724 (N_12724,N_10851,N_11264);
xnor U12725 (N_12725,N_11546,N_10352);
nand U12726 (N_12726,N_11292,N_10633);
nor U12727 (N_12727,N_11141,N_10820);
and U12728 (N_12728,N_10101,N_11994);
nor U12729 (N_12729,N_10196,N_10786);
or U12730 (N_12730,N_10744,N_11925);
and U12731 (N_12731,N_11281,N_10237);
xor U12732 (N_12732,N_10180,N_10724);
nor U12733 (N_12733,N_11383,N_10481);
and U12734 (N_12734,N_10881,N_11745);
xnor U12735 (N_12735,N_10701,N_10172);
or U12736 (N_12736,N_11261,N_10488);
nor U12737 (N_12737,N_10492,N_10344);
xnor U12738 (N_12738,N_10143,N_11572);
or U12739 (N_12739,N_11919,N_10504);
nor U12740 (N_12740,N_11182,N_10330);
xnor U12741 (N_12741,N_10842,N_10007);
nand U12742 (N_12742,N_10641,N_10036);
and U12743 (N_12743,N_10131,N_11266);
and U12744 (N_12744,N_11661,N_10179);
and U12745 (N_12745,N_10773,N_10373);
nor U12746 (N_12746,N_10407,N_10057);
and U12747 (N_12747,N_11663,N_10288);
nor U12748 (N_12748,N_10838,N_11915);
nand U12749 (N_12749,N_11015,N_11380);
or U12750 (N_12750,N_10252,N_10919);
and U12751 (N_12751,N_11758,N_10855);
or U12752 (N_12752,N_11625,N_10852);
and U12753 (N_12753,N_10891,N_11871);
nor U12754 (N_12754,N_10152,N_11553);
and U12755 (N_12755,N_11822,N_11673);
nand U12756 (N_12756,N_11482,N_11310);
nand U12757 (N_12757,N_10326,N_11174);
nor U12758 (N_12758,N_10329,N_11371);
and U12759 (N_12759,N_11194,N_11314);
nand U12760 (N_12760,N_11263,N_10316);
xor U12761 (N_12761,N_10848,N_10394);
nand U12762 (N_12762,N_11395,N_11031);
nand U12763 (N_12763,N_10341,N_10814);
nand U12764 (N_12764,N_10307,N_11342);
nand U12765 (N_12765,N_11095,N_11716);
and U12766 (N_12766,N_11707,N_10788);
and U12767 (N_12767,N_10129,N_10975);
nor U12768 (N_12768,N_10164,N_10178);
nor U12769 (N_12769,N_11198,N_11366);
or U12770 (N_12770,N_10496,N_10737);
nand U12771 (N_12771,N_11736,N_11192);
and U12772 (N_12772,N_11297,N_10658);
nor U12773 (N_12773,N_10008,N_11690);
and U12774 (N_12774,N_10322,N_10869);
or U12775 (N_12775,N_10060,N_10627);
or U12776 (N_12776,N_10414,N_10157);
or U12777 (N_12777,N_11166,N_10536);
or U12778 (N_12778,N_11249,N_11932);
or U12779 (N_12779,N_10597,N_11278);
and U12780 (N_12780,N_10991,N_11514);
or U12781 (N_12781,N_11896,N_11180);
xor U12782 (N_12782,N_10935,N_11820);
xnor U12783 (N_12783,N_11111,N_10395);
nor U12784 (N_12784,N_10859,N_11647);
or U12785 (N_12785,N_11164,N_11618);
or U12786 (N_12786,N_11761,N_11092);
nand U12787 (N_12787,N_11817,N_10000);
nand U12788 (N_12788,N_10907,N_10382);
nand U12789 (N_12789,N_10025,N_11421);
nand U12790 (N_12790,N_10706,N_11463);
xor U12791 (N_12791,N_10659,N_11535);
nand U12792 (N_12792,N_10456,N_11105);
xor U12793 (N_12793,N_10251,N_10218);
nand U12794 (N_12794,N_10372,N_11628);
and U12795 (N_12795,N_11656,N_11073);
nor U12796 (N_12796,N_10410,N_11710);
and U12797 (N_12797,N_10540,N_10154);
and U12798 (N_12798,N_11669,N_11616);
or U12799 (N_12799,N_10685,N_10630);
and U12800 (N_12800,N_11590,N_10461);
nor U12801 (N_12801,N_10957,N_11511);
or U12802 (N_12802,N_11619,N_10834);
nand U12803 (N_12803,N_11973,N_10233);
and U12804 (N_12804,N_11781,N_11641);
and U12805 (N_12805,N_11547,N_11520);
nand U12806 (N_12806,N_10525,N_10583);
or U12807 (N_12807,N_11888,N_11500);
nand U12808 (N_12808,N_10981,N_11575);
and U12809 (N_12809,N_10947,N_10324);
or U12810 (N_12810,N_10768,N_10533);
and U12811 (N_12811,N_10241,N_11762);
xor U12812 (N_12812,N_11927,N_10351);
and U12813 (N_12813,N_11998,N_10708);
nand U12814 (N_12814,N_10837,N_10347);
or U12815 (N_12815,N_10238,N_10511);
nand U12816 (N_12816,N_11478,N_10984);
nand U12817 (N_12817,N_11920,N_11565);
or U12818 (N_12818,N_10623,N_11262);
and U12819 (N_12819,N_10847,N_11918);
nand U12820 (N_12820,N_10197,N_11147);
and U12821 (N_12821,N_11271,N_11170);
nand U12822 (N_12822,N_10520,N_10059);
nand U12823 (N_12823,N_11718,N_11594);
nand U12824 (N_12824,N_11598,N_11801);
nand U12825 (N_12825,N_10214,N_10713);
and U12826 (N_12826,N_11449,N_10003);
or U12827 (N_12827,N_11773,N_10130);
nand U12828 (N_12828,N_11360,N_10155);
nor U12829 (N_12829,N_11991,N_11560);
nand U12830 (N_12830,N_11691,N_11321);
nor U12831 (N_12831,N_11703,N_11413);
nand U12832 (N_12832,N_11833,N_11517);
nor U12833 (N_12833,N_10020,N_11265);
xnor U12834 (N_12834,N_10792,N_10165);
or U12835 (N_12835,N_11428,N_10554);
and U12836 (N_12836,N_11954,N_11652);
nor U12837 (N_12837,N_10720,N_11188);
and U12838 (N_12838,N_10277,N_10746);
or U12839 (N_12839,N_11681,N_11672);
or U12840 (N_12840,N_10705,N_11724);
nor U12841 (N_12841,N_10664,N_10651);
or U12842 (N_12842,N_11238,N_11655);
and U12843 (N_12843,N_11868,N_10049);
nor U12844 (N_12844,N_10550,N_10896);
and U12845 (N_12845,N_11855,N_11353);
and U12846 (N_12846,N_11355,N_10718);
or U12847 (N_12847,N_11368,N_10808);
nor U12848 (N_12848,N_10694,N_11341);
and U12849 (N_12849,N_10445,N_11235);
nor U12850 (N_12850,N_10552,N_10392);
or U12851 (N_12851,N_11053,N_10061);
xor U12852 (N_12852,N_10100,N_10542);
or U12853 (N_12853,N_10969,N_10080);
xor U12854 (N_12854,N_10692,N_10262);
nor U12855 (N_12855,N_11775,N_11522);
nor U12856 (N_12856,N_11810,N_11446);
xor U12857 (N_12857,N_10085,N_11347);
nand U12858 (N_12858,N_11241,N_10866);
xor U12859 (N_12859,N_10345,N_11311);
or U12860 (N_12860,N_10231,N_11459);
nand U12861 (N_12861,N_11726,N_11247);
nand U12862 (N_12862,N_10423,N_11686);
and U12863 (N_12863,N_11664,N_10529);
or U12864 (N_12864,N_11671,N_11639);
nand U12865 (N_12865,N_11885,N_10950);
xnor U12866 (N_12866,N_11823,N_10844);
or U12867 (N_12867,N_11336,N_11877);
or U12868 (N_12868,N_10483,N_11668);
and U12869 (N_12869,N_10675,N_10807);
nor U12870 (N_12870,N_11978,N_11693);
and U12871 (N_12871,N_10463,N_10965);
or U12872 (N_12872,N_11070,N_11307);
nor U12873 (N_12873,N_11004,N_11518);
nor U12874 (N_12874,N_10930,N_10586);
or U12875 (N_12875,N_10062,N_11134);
nand U12876 (N_12876,N_10289,N_10202);
nor U12877 (N_12877,N_11831,N_11439);
or U12878 (N_12878,N_11934,N_11592);
nand U12879 (N_12879,N_11312,N_10439);
or U12880 (N_12880,N_11543,N_10448);
nand U12881 (N_12881,N_10495,N_10691);
nor U12882 (N_12882,N_10040,N_11148);
and U12883 (N_12883,N_11561,N_11530);
or U12884 (N_12884,N_11390,N_10258);
nand U12885 (N_12885,N_11322,N_11203);
and U12886 (N_12886,N_10148,N_10471);
nand U12887 (N_12887,N_10956,N_11420);
or U12888 (N_12888,N_10039,N_11582);
and U12889 (N_12889,N_11207,N_10770);
or U12890 (N_12890,N_10239,N_11185);
and U12891 (N_12891,N_10726,N_10924);
xnor U12892 (N_12892,N_10263,N_11503);
nand U12893 (N_12893,N_11237,N_11648);
nand U12894 (N_12894,N_11494,N_11470);
nand U12895 (N_12895,N_10679,N_11739);
nand U12896 (N_12896,N_11076,N_11457);
nand U12897 (N_12897,N_11162,N_11870);
nand U12898 (N_12898,N_11121,N_11351);
nand U12899 (N_12899,N_10426,N_11130);
nor U12900 (N_12900,N_10099,N_11486);
and U12901 (N_12901,N_11160,N_10789);
or U12902 (N_12902,N_10811,N_10502);
nor U12903 (N_12903,N_10962,N_10764);
and U12904 (N_12904,N_10425,N_10306);
and U12905 (N_12905,N_10722,N_11636);
and U12906 (N_12906,N_10086,N_11931);
and U12907 (N_12907,N_11240,N_11399);
nor U12908 (N_12908,N_10783,N_10071);
or U12909 (N_12909,N_10959,N_10854);
or U12910 (N_12910,N_10865,N_11219);
or U12911 (N_12911,N_11433,N_11202);
nand U12912 (N_12912,N_11538,N_10438);
or U12913 (N_12913,N_10286,N_10109);
and U12914 (N_12914,N_10660,N_10303);
and U12915 (N_12915,N_10487,N_11512);
nand U12916 (N_12916,N_10389,N_10400);
xor U12917 (N_12917,N_11544,N_10257);
xor U12918 (N_12918,N_10840,N_10102);
nor U12919 (N_12919,N_10397,N_10576);
and U12920 (N_12920,N_10005,N_11038);
nand U12921 (N_12921,N_10534,N_10301);
xnor U12922 (N_12922,N_10122,N_11186);
xor U12923 (N_12923,N_11140,N_10565);
and U12924 (N_12924,N_10833,N_10505);
xnor U12925 (N_12925,N_10680,N_10226);
nor U12926 (N_12926,N_11361,N_11404);
or U12927 (N_12927,N_10571,N_10338);
xnor U12928 (N_12928,N_10539,N_10248);
and U12929 (N_12929,N_10835,N_10822);
and U12930 (N_12930,N_10549,N_11136);
nor U12931 (N_12931,N_11630,N_11047);
and U12932 (N_12932,N_11599,N_11688);
and U12933 (N_12933,N_11206,N_11640);
nor U12934 (N_12934,N_10266,N_10943);
and U12935 (N_12935,N_10244,N_11965);
or U12936 (N_12936,N_11364,N_10365);
and U12937 (N_12937,N_10088,N_10555);
and U12938 (N_12938,N_10072,N_11617);
nand U12939 (N_12939,N_10845,N_10234);
or U12940 (N_12940,N_10300,N_10150);
nor U12941 (N_12941,N_10167,N_11458);
xnor U12942 (N_12942,N_10107,N_11782);
and U12943 (N_12943,N_10272,N_10932);
xnor U12944 (N_12944,N_10356,N_10871);
or U12945 (N_12945,N_11320,N_11788);
or U12946 (N_12946,N_11018,N_11302);
and U12947 (N_12947,N_11895,N_11554);
nand U12948 (N_12948,N_11700,N_10649);
or U12949 (N_12949,N_11269,N_10474);
nor U12950 (N_12950,N_10269,N_10690);
nand U12951 (N_12951,N_11098,N_11573);
and U12952 (N_12952,N_10676,N_11956);
nand U12953 (N_12953,N_11246,N_11563);
nand U12954 (N_12954,N_10531,N_10864);
nand U12955 (N_12955,N_11232,N_10034);
xor U12956 (N_12956,N_10621,N_11019);
or U12957 (N_12957,N_10728,N_10405);
nand U12958 (N_12958,N_10774,N_10270);
and U12959 (N_12959,N_10846,N_11846);
nor U12960 (N_12960,N_10050,N_10922);
and U12961 (N_12961,N_10318,N_11172);
nor U12962 (N_12962,N_10498,N_11438);
and U12963 (N_12963,N_11423,N_11303);
or U12964 (N_12964,N_11325,N_11374);
nor U12965 (N_12965,N_11622,N_11634);
nor U12966 (N_12966,N_11829,N_10317);
nor U12967 (N_12967,N_11083,N_10171);
or U12968 (N_12968,N_10886,N_11118);
and U12969 (N_12969,N_11650,N_10123);
and U12970 (N_12970,N_10208,N_10954);
and U12971 (N_12971,N_11643,N_11484);
and U12972 (N_12972,N_10661,N_11613);
nand U12973 (N_12973,N_11454,N_11528);
and U12974 (N_12974,N_11813,N_11456);
or U12975 (N_12975,N_11682,N_11695);
xor U12976 (N_12976,N_11343,N_11907);
and U12977 (N_12977,N_11988,N_11930);
or U12978 (N_12978,N_10933,N_11177);
and U12979 (N_12979,N_11879,N_10083);
xor U12980 (N_12980,N_11481,N_11392);
or U12981 (N_12981,N_10312,N_10810);
and U12982 (N_12982,N_11880,N_10256);
and U12983 (N_12983,N_10605,N_11536);
and U12984 (N_12984,N_10735,N_11305);
and U12985 (N_12985,N_11772,N_11717);
and U12986 (N_12986,N_10089,N_11580);
or U12987 (N_12987,N_11101,N_10412);
nand U12988 (N_12988,N_10374,N_11274);
and U12989 (N_12989,N_10669,N_11437);
and U12990 (N_12990,N_11097,N_11487);
and U12991 (N_12991,N_10883,N_11853);
or U12992 (N_12992,N_11730,N_11699);
nor U12993 (N_12993,N_10116,N_11900);
and U12994 (N_12994,N_11728,N_10139);
nor U12995 (N_12995,N_10355,N_11063);
and U12996 (N_12996,N_10334,N_10362);
nor U12997 (N_12997,N_11532,N_11315);
and U12998 (N_12998,N_10297,N_11778);
and U12999 (N_12999,N_11096,N_10219);
or U13000 (N_13000,N_11629,N_11683);
and U13001 (N_13001,N_10364,N_10369);
nor U13002 (N_13002,N_10516,N_10640);
nand U13003 (N_13003,N_11748,N_10368);
and U13004 (N_13004,N_10755,N_10352);
nor U13005 (N_13005,N_10680,N_10459);
or U13006 (N_13006,N_11862,N_11758);
nand U13007 (N_13007,N_11622,N_11974);
nand U13008 (N_13008,N_11476,N_10769);
and U13009 (N_13009,N_11163,N_10774);
nor U13010 (N_13010,N_10339,N_10246);
nand U13011 (N_13011,N_10422,N_11696);
nand U13012 (N_13012,N_10856,N_11538);
xor U13013 (N_13013,N_11192,N_10758);
and U13014 (N_13014,N_10811,N_11591);
nor U13015 (N_13015,N_11011,N_11388);
or U13016 (N_13016,N_10438,N_10403);
nand U13017 (N_13017,N_10943,N_11971);
or U13018 (N_13018,N_11429,N_11503);
nand U13019 (N_13019,N_10752,N_11232);
and U13020 (N_13020,N_10406,N_11166);
or U13021 (N_13021,N_10723,N_11358);
nor U13022 (N_13022,N_11346,N_11116);
or U13023 (N_13023,N_11587,N_11856);
nor U13024 (N_13024,N_11445,N_10938);
or U13025 (N_13025,N_11390,N_11860);
or U13026 (N_13026,N_10607,N_10493);
or U13027 (N_13027,N_10132,N_11272);
xor U13028 (N_13028,N_11268,N_10266);
or U13029 (N_13029,N_10627,N_11491);
and U13030 (N_13030,N_11266,N_11984);
and U13031 (N_13031,N_11244,N_11115);
nor U13032 (N_13032,N_10544,N_10428);
or U13033 (N_13033,N_10277,N_10917);
and U13034 (N_13034,N_10711,N_11252);
and U13035 (N_13035,N_11492,N_10159);
nor U13036 (N_13036,N_11190,N_11553);
and U13037 (N_13037,N_10083,N_10403);
nor U13038 (N_13038,N_10530,N_10771);
or U13039 (N_13039,N_11587,N_11520);
nand U13040 (N_13040,N_10444,N_10925);
and U13041 (N_13041,N_10281,N_10148);
or U13042 (N_13042,N_10825,N_11282);
nor U13043 (N_13043,N_10799,N_11414);
nor U13044 (N_13044,N_10832,N_10949);
nor U13045 (N_13045,N_11414,N_11556);
or U13046 (N_13046,N_11525,N_11024);
or U13047 (N_13047,N_10159,N_11159);
nor U13048 (N_13048,N_10523,N_11809);
xnor U13049 (N_13049,N_10957,N_11691);
or U13050 (N_13050,N_11868,N_10710);
and U13051 (N_13051,N_11950,N_11682);
or U13052 (N_13052,N_11189,N_10587);
or U13053 (N_13053,N_10942,N_10563);
nand U13054 (N_13054,N_10319,N_10233);
or U13055 (N_13055,N_11318,N_10496);
nor U13056 (N_13056,N_11476,N_10281);
nor U13057 (N_13057,N_11941,N_10871);
nor U13058 (N_13058,N_10963,N_10704);
or U13059 (N_13059,N_10997,N_11869);
or U13060 (N_13060,N_11182,N_10554);
or U13061 (N_13061,N_10867,N_11201);
nor U13062 (N_13062,N_11104,N_11148);
xnor U13063 (N_13063,N_11422,N_10468);
or U13064 (N_13064,N_11286,N_10335);
nand U13065 (N_13065,N_11399,N_11496);
and U13066 (N_13066,N_11357,N_11302);
xnor U13067 (N_13067,N_11435,N_10326);
or U13068 (N_13068,N_10599,N_11127);
nor U13069 (N_13069,N_11235,N_11465);
xor U13070 (N_13070,N_11898,N_11367);
or U13071 (N_13071,N_11266,N_10209);
and U13072 (N_13072,N_11704,N_10007);
or U13073 (N_13073,N_11451,N_10083);
or U13074 (N_13074,N_11342,N_10723);
and U13075 (N_13075,N_11707,N_11744);
nor U13076 (N_13076,N_11855,N_10848);
nor U13077 (N_13077,N_10296,N_11106);
or U13078 (N_13078,N_11968,N_11502);
nor U13079 (N_13079,N_10712,N_10179);
nand U13080 (N_13080,N_10523,N_11976);
xor U13081 (N_13081,N_10287,N_11385);
nand U13082 (N_13082,N_10081,N_10253);
nor U13083 (N_13083,N_11320,N_10916);
or U13084 (N_13084,N_10277,N_10998);
or U13085 (N_13085,N_10546,N_11057);
or U13086 (N_13086,N_11600,N_10991);
nor U13087 (N_13087,N_11582,N_10473);
nor U13088 (N_13088,N_10744,N_11281);
and U13089 (N_13089,N_11223,N_11917);
nor U13090 (N_13090,N_10962,N_10588);
xor U13091 (N_13091,N_10800,N_11683);
and U13092 (N_13092,N_10088,N_11236);
and U13093 (N_13093,N_11961,N_11103);
xor U13094 (N_13094,N_11093,N_10685);
and U13095 (N_13095,N_11514,N_11449);
nand U13096 (N_13096,N_11541,N_10587);
and U13097 (N_13097,N_10195,N_10505);
or U13098 (N_13098,N_10609,N_11061);
xnor U13099 (N_13099,N_10672,N_11294);
xnor U13100 (N_13100,N_11099,N_11569);
nand U13101 (N_13101,N_10551,N_11910);
and U13102 (N_13102,N_11885,N_10824);
xnor U13103 (N_13103,N_10769,N_10256);
and U13104 (N_13104,N_11740,N_11690);
nand U13105 (N_13105,N_10562,N_11627);
or U13106 (N_13106,N_11826,N_11956);
and U13107 (N_13107,N_10928,N_10942);
or U13108 (N_13108,N_11062,N_10601);
xnor U13109 (N_13109,N_11651,N_10752);
nand U13110 (N_13110,N_10043,N_11429);
nand U13111 (N_13111,N_10004,N_11269);
and U13112 (N_13112,N_11450,N_10996);
or U13113 (N_13113,N_10910,N_10598);
and U13114 (N_13114,N_10726,N_11689);
or U13115 (N_13115,N_11939,N_11525);
xor U13116 (N_13116,N_10641,N_10923);
nor U13117 (N_13117,N_11687,N_10819);
nand U13118 (N_13118,N_10024,N_10442);
nor U13119 (N_13119,N_11525,N_10742);
and U13120 (N_13120,N_11698,N_11012);
nand U13121 (N_13121,N_11456,N_10073);
nor U13122 (N_13122,N_10141,N_10225);
nor U13123 (N_13123,N_10931,N_10124);
nand U13124 (N_13124,N_11391,N_11988);
and U13125 (N_13125,N_11860,N_10333);
nor U13126 (N_13126,N_11736,N_10182);
nand U13127 (N_13127,N_10731,N_10506);
or U13128 (N_13128,N_10800,N_10425);
nor U13129 (N_13129,N_10446,N_11153);
or U13130 (N_13130,N_10205,N_10119);
xnor U13131 (N_13131,N_10074,N_11205);
nand U13132 (N_13132,N_10998,N_10316);
or U13133 (N_13133,N_10597,N_10669);
or U13134 (N_13134,N_11182,N_10083);
or U13135 (N_13135,N_10520,N_11779);
nor U13136 (N_13136,N_10767,N_11556);
and U13137 (N_13137,N_10803,N_11045);
nor U13138 (N_13138,N_11554,N_10931);
nor U13139 (N_13139,N_10857,N_10458);
and U13140 (N_13140,N_10856,N_11561);
nand U13141 (N_13141,N_10166,N_10782);
and U13142 (N_13142,N_11818,N_10356);
or U13143 (N_13143,N_10191,N_10612);
or U13144 (N_13144,N_11353,N_11085);
and U13145 (N_13145,N_10412,N_10614);
or U13146 (N_13146,N_11833,N_11279);
and U13147 (N_13147,N_11691,N_10950);
and U13148 (N_13148,N_10063,N_11549);
nor U13149 (N_13149,N_10699,N_11450);
or U13150 (N_13150,N_10107,N_10907);
nand U13151 (N_13151,N_10532,N_10707);
nor U13152 (N_13152,N_10666,N_11364);
or U13153 (N_13153,N_11060,N_11746);
and U13154 (N_13154,N_11701,N_10966);
nor U13155 (N_13155,N_11420,N_10715);
and U13156 (N_13156,N_11686,N_11191);
nand U13157 (N_13157,N_10055,N_10736);
nand U13158 (N_13158,N_11019,N_11871);
nand U13159 (N_13159,N_10417,N_11477);
nor U13160 (N_13160,N_11278,N_10514);
and U13161 (N_13161,N_10994,N_10008);
nand U13162 (N_13162,N_11244,N_11676);
and U13163 (N_13163,N_11713,N_10800);
and U13164 (N_13164,N_10835,N_10434);
nand U13165 (N_13165,N_10482,N_11489);
or U13166 (N_13166,N_11482,N_10291);
and U13167 (N_13167,N_10298,N_11724);
or U13168 (N_13168,N_10773,N_10670);
xor U13169 (N_13169,N_11105,N_10034);
or U13170 (N_13170,N_10705,N_11463);
nand U13171 (N_13171,N_11282,N_11542);
nor U13172 (N_13172,N_11522,N_10276);
nand U13173 (N_13173,N_10834,N_10349);
and U13174 (N_13174,N_10397,N_11716);
or U13175 (N_13175,N_10868,N_10996);
nand U13176 (N_13176,N_10073,N_11558);
nand U13177 (N_13177,N_11616,N_10715);
or U13178 (N_13178,N_11700,N_10090);
or U13179 (N_13179,N_10350,N_10082);
and U13180 (N_13180,N_10694,N_11189);
nor U13181 (N_13181,N_11313,N_10274);
or U13182 (N_13182,N_10177,N_11570);
and U13183 (N_13183,N_10345,N_10637);
and U13184 (N_13184,N_11379,N_11925);
or U13185 (N_13185,N_10885,N_11883);
xnor U13186 (N_13186,N_11874,N_11367);
or U13187 (N_13187,N_11847,N_10170);
and U13188 (N_13188,N_10911,N_11487);
nand U13189 (N_13189,N_10259,N_10093);
nand U13190 (N_13190,N_11257,N_10346);
nand U13191 (N_13191,N_11005,N_10711);
or U13192 (N_13192,N_10941,N_10483);
or U13193 (N_13193,N_10378,N_10047);
nand U13194 (N_13194,N_11845,N_10004);
nor U13195 (N_13195,N_10935,N_10547);
xor U13196 (N_13196,N_10414,N_11095);
nor U13197 (N_13197,N_10897,N_10355);
or U13198 (N_13198,N_11860,N_10727);
nand U13199 (N_13199,N_10165,N_11576);
or U13200 (N_13200,N_10247,N_11401);
nor U13201 (N_13201,N_11027,N_11418);
nor U13202 (N_13202,N_10440,N_10772);
nor U13203 (N_13203,N_10082,N_10353);
xnor U13204 (N_13204,N_11507,N_11517);
nand U13205 (N_13205,N_11405,N_10588);
xor U13206 (N_13206,N_11992,N_10646);
nand U13207 (N_13207,N_10301,N_10069);
nand U13208 (N_13208,N_11714,N_11579);
nand U13209 (N_13209,N_11556,N_11763);
or U13210 (N_13210,N_11199,N_10788);
nand U13211 (N_13211,N_11154,N_10323);
or U13212 (N_13212,N_10493,N_11409);
or U13213 (N_13213,N_11921,N_11773);
xnor U13214 (N_13214,N_10274,N_11378);
xnor U13215 (N_13215,N_10133,N_11243);
xor U13216 (N_13216,N_10077,N_10551);
or U13217 (N_13217,N_11932,N_11034);
nor U13218 (N_13218,N_11213,N_10762);
nand U13219 (N_13219,N_11717,N_10175);
or U13220 (N_13220,N_11056,N_10151);
nor U13221 (N_13221,N_10498,N_11128);
and U13222 (N_13222,N_10611,N_11526);
nand U13223 (N_13223,N_11171,N_10564);
nor U13224 (N_13224,N_10963,N_11799);
and U13225 (N_13225,N_11220,N_11432);
or U13226 (N_13226,N_11065,N_10415);
and U13227 (N_13227,N_11823,N_11717);
nand U13228 (N_13228,N_11524,N_11820);
nand U13229 (N_13229,N_11714,N_10342);
or U13230 (N_13230,N_10644,N_11149);
nand U13231 (N_13231,N_11402,N_10316);
and U13232 (N_13232,N_11576,N_11500);
xor U13233 (N_13233,N_10895,N_10475);
nor U13234 (N_13234,N_10959,N_11668);
xnor U13235 (N_13235,N_11280,N_11985);
nor U13236 (N_13236,N_11429,N_10205);
nor U13237 (N_13237,N_11605,N_10072);
nor U13238 (N_13238,N_10670,N_10454);
or U13239 (N_13239,N_11414,N_11359);
nor U13240 (N_13240,N_11214,N_11325);
and U13241 (N_13241,N_10132,N_11942);
nor U13242 (N_13242,N_10072,N_10642);
nor U13243 (N_13243,N_11096,N_11285);
or U13244 (N_13244,N_10070,N_10755);
or U13245 (N_13245,N_10175,N_10754);
and U13246 (N_13246,N_11790,N_11605);
nor U13247 (N_13247,N_10616,N_10352);
and U13248 (N_13248,N_11045,N_10205);
and U13249 (N_13249,N_11190,N_10391);
xnor U13250 (N_13250,N_11556,N_10253);
nand U13251 (N_13251,N_10622,N_11887);
nand U13252 (N_13252,N_10708,N_10229);
nand U13253 (N_13253,N_10406,N_11946);
nand U13254 (N_13254,N_10182,N_11665);
or U13255 (N_13255,N_11255,N_10179);
nor U13256 (N_13256,N_10204,N_10979);
and U13257 (N_13257,N_11011,N_11880);
nor U13258 (N_13258,N_11043,N_10624);
or U13259 (N_13259,N_10586,N_11331);
and U13260 (N_13260,N_11259,N_10877);
and U13261 (N_13261,N_11029,N_11175);
xor U13262 (N_13262,N_11366,N_10400);
nor U13263 (N_13263,N_11266,N_11645);
or U13264 (N_13264,N_10827,N_11491);
and U13265 (N_13265,N_11692,N_11543);
xor U13266 (N_13266,N_11711,N_10888);
nor U13267 (N_13267,N_10328,N_10961);
nand U13268 (N_13268,N_10357,N_11847);
nor U13269 (N_13269,N_10324,N_11152);
and U13270 (N_13270,N_10307,N_11850);
nand U13271 (N_13271,N_10582,N_11635);
or U13272 (N_13272,N_11856,N_11133);
nor U13273 (N_13273,N_11961,N_11292);
nand U13274 (N_13274,N_10494,N_10946);
xnor U13275 (N_13275,N_10843,N_11720);
and U13276 (N_13276,N_10182,N_11834);
nor U13277 (N_13277,N_10371,N_11037);
or U13278 (N_13278,N_10952,N_11113);
or U13279 (N_13279,N_11604,N_11865);
nor U13280 (N_13280,N_10415,N_10265);
or U13281 (N_13281,N_11642,N_10981);
and U13282 (N_13282,N_10440,N_10586);
or U13283 (N_13283,N_10648,N_11296);
xor U13284 (N_13284,N_11700,N_10143);
nand U13285 (N_13285,N_10141,N_11288);
nor U13286 (N_13286,N_10581,N_10728);
nand U13287 (N_13287,N_11231,N_10556);
nor U13288 (N_13288,N_10190,N_11317);
nor U13289 (N_13289,N_11255,N_11752);
nand U13290 (N_13290,N_10740,N_11426);
xnor U13291 (N_13291,N_10930,N_10319);
or U13292 (N_13292,N_11108,N_11289);
and U13293 (N_13293,N_10754,N_11851);
or U13294 (N_13294,N_10391,N_11678);
xor U13295 (N_13295,N_11821,N_11053);
and U13296 (N_13296,N_10082,N_10589);
nor U13297 (N_13297,N_11221,N_10770);
xnor U13298 (N_13298,N_10101,N_11426);
and U13299 (N_13299,N_10529,N_10831);
or U13300 (N_13300,N_10002,N_11698);
xor U13301 (N_13301,N_10040,N_10660);
and U13302 (N_13302,N_10763,N_10250);
or U13303 (N_13303,N_10341,N_11949);
xor U13304 (N_13304,N_11262,N_11907);
nand U13305 (N_13305,N_11382,N_10257);
and U13306 (N_13306,N_11855,N_11483);
xnor U13307 (N_13307,N_10586,N_11173);
or U13308 (N_13308,N_11312,N_10582);
or U13309 (N_13309,N_11472,N_10663);
nand U13310 (N_13310,N_10364,N_10102);
or U13311 (N_13311,N_11893,N_10059);
or U13312 (N_13312,N_11384,N_11110);
xnor U13313 (N_13313,N_10234,N_11697);
nand U13314 (N_13314,N_11349,N_10071);
nor U13315 (N_13315,N_11280,N_11752);
and U13316 (N_13316,N_11235,N_10432);
xnor U13317 (N_13317,N_11286,N_10382);
nand U13318 (N_13318,N_11657,N_10140);
nor U13319 (N_13319,N_11391,N_11688);
nor U13320 (N_13320,N_11227,N_10704);
nor U13321 (N_13321,N_11092,N_11006);
or U13322 (N_13322,N_11702,N_10188);
and U13323 (N_13323,N_11991,N_11358);
nor U13324 (N_13324,N_11604,N_10810);
and U13325 (N_13325,N_10181,N_11575);
or U13326 (N_13326,N_11769,N_11007);
and U13327 (N_13327,N_11503,N_11591);
and U13328 (N_13328,N_11435,N_11186);
nor U13329 (N_13329,N_10444,N_10579);
nand U13330 (N_13330,N_10154,N_10998);
or U13331 (N_13331,N_10552,N_10646);
or U13332 (N_13332,N_10089,N_11644);
and U13333 (N_13333,N_11962,N_10119);
nor U13334 (N_13334,N_10866,N_11579);
nor U13335 (N_13335,N_10084,N_10755);
xor U13336 (N_13336,N_11115,N_10758);
or U13337 (N_13337,N_11102,N_10937);
nand U13338 (N_13338,N_11434,N_10873);
nand U13339 (N_13339,N_11661,N_10610);
or U13340 (N_13340,N_11031,N_11062);
or U13341 (N_13341,N_10509,N_10856);
nor U13342 (N_13342,N_11194,N_10729);
or U13343 (N_13343,N_10735,N_11803);
or U13344 (N_13344,N_11901,N_10792);
xor U13345 (N_13345,N_11284,N_10885);
xnor U13346 (N_13346,N_11389,N_11823);
or U13347 (N_13347,N_10148,N_10552);
or U13348 (N_13348,N_10296,N_10511);
or U13349 (N_13349,N_10790,N_11616);
or U13350 (N_13350,N_10664,N_11420);
and U13351 (N_13351,N_10144,N_11359);
nor U13352 (N_13352,N_11660,N_10147);
or U13353 (N_13353,N_11989,N_11663);
nor U13354 (N_13354,N_11665,N_10980);
or U13355 (N_13355,N_11920,N_11134);
and U13356 (N_13356,N_10480,N_10243);
and U13357 (N_13357,N_10330,N_10802);
or U13358 (N_13358,N_10723,N_10651);
nand U13359 (N_13359,N_10423,N_10064);
and U13360 (N_13360,N_10073,N_11394);
or U13361 (N_13361,N_10010,N_10202);
or U13362 (N_13362,N_11049,N_11935);
xnor U13363 (N_13363,N_10744,N_11032);
or U13364 (N_13364,N_10426,N_11502);
and U13365 (N_13365,N_11733,N_10534);
xnor U13366 (N_13366,N_10482,N_10599);
and U13367 (N_13367,N_10879,N_10400);
or U13368 (N_13368,N_10952,N_11979);
or U13369 (N_13369,N_10669,N_11844);
nand U13370 (N_13370,N_10025,N_10143);
or U13371 (N_13371,N_10202,N_10701);
nor U13372 (N_13372,N_11318,N_11090);
or U13373 (N_13373,N_10369,N_11454);
or U13374 (N_13374,N_10413,N_11526);
and U13375 (N_13375,N_10150,N_11755);
and U13376 (N_13376,N_11445,N_11012);
or U13377 (N_13377,N_10458,N_11540);
or U13378 (N_13378,N_11882,N_10800);
or U13379 (N_13379,N_10381,N_11499);
nor U13380 (N_13380,N_10828,N_10682);
or U13381 (N_13381,N_10188,N_10104);
or U13382 (N_13382,N_11452,N_11152);
or U13383 (N_13383,N_10122,N_11813);
nand U13384 (N_13384,N_11331,N_11043);
nand U13385 (N_13385,N_10221,N_10724);
and U13386 (N_13386,N_11032,N_10099);
nor U13387 (N_13387,N_11708,N_11224);
nand U13388 (N_13388,N_10252,N_10439);
or U13389 (N_13389,N_10706,N_10790);
nor U13390 (N_13390,N_11796,N_11843);
and U13391 (N_13391,N_10084,N_10156);
nor U13392 (N_13392,N_10927,N_11680);
or U13393 (N_13393,N_10797,N_11024);
nand U13394 (N_13394,N_10888,N_11384);
nand U13395 (N_13395,N_11938,N_11337);
and U13396 (N_13396,N_10689,N_11083);
nor U13397 (N_13397,N_10050,N_10141);
or U13398 (N_13398,N_11387,N_11631);
nand U13399 (N_13399,N_11461,N_11541);
or U13400 (N_13400,N_11564,N_11845);
nor U13401 (N_13401,N_10284,N_11466);
nand U13402 (N_13402,N_11711,N_10127);
nor U13403 (N_13403,N_11656,N_11945);
xnor U13404 (N_13404,N_10614,N_11859);
xor U13405 (N_13405,N_11359,N_11412);
nor U13406 (N_13406,N_11940,N_10919);
and U13407 (N_13407,N_10335,N_10629);
nand U13408 (N_13408,N_10956,N_11885);
nand U13409 (N_13409,N_11579,N_10147);
or U13410 (N_13410,N_10489,N_10131);
nor U13411 (N_13411,N_10362,N_10380);
or U13412 (N_13412,N_10008,N_10933);
nand U13413 (N_13413,N_11224,N_10760);
xnor U13414 (N_13414,N_11553,N_10298);
or U13415 (N_13415,N_10495,N_11767);
or U13416 (N_13416,N_10809,N_11459);
or U13417 (N_13417,N_10633,N_10430);
or U13418 (N_13418,N_11880,N_11721);
nand U13419 (N_13419,N_11518,N_11420);
or U13420 (N_13420,N_11815,N_11826);
and U13421 (N_13421,N_10831,N_11857);
and U13422 (N_13422,N_11798,N_10412);
and U13423 (N_13423,N_11022,N_11406);
nor U13424 (N_13424,N_11646,N_11706);
nand U13425 (N_13425,N_10615,N_11999);
and U13426 (N_13426,N_11291,N_10455);
nor U13427 (N_13427,N_11319,N_11103);
nand U13428 (N_13428,N_10254,N_11157);
or U13429 (N_13429,N_11634,N_11453);
or U13430 (N_13430,N_10224,N_11413);
and U13431 (N_13431,N_11785,N_10174);
nand U13432 (N_13432,N_11953,N_10131);
nor U13433 (N_13433,N_11333,N_11457);
and U13434 (N_13434,N_11866,N_11914);
nand U13435 (N_13435,N_11368,N_11286);
or U13436 (N_13436,N_11351,N_10249);
nand U13437 (N_13437,N_10618,N_11520);
nor U13438 (N_13438,N_10117,N_11321);
nand U13439 (N_13439,N_11391,N_10666);
or U13440 (N_13440,N_11247,N_10929);
nand U13441 (N_13441,N_11957,N_11196);
nand U13442 (N_13442,N_10730,N_10859);
or U13443 (N_13443,N_11016,N_11826);
nand U13444 (N_13444,N_11648,N_10320);
nand U13445 (N_13445,N_11077,N_11428);
nor U13446 (N_13446,N_10770,N_11325);
nand U13447 (N_13447,N_10782,N_11978);
nor U13448 (N_13448,N_10226,N_11231);
nand U13449 (N_13449,N_10035,N_10437);
or U13450 (N_13450,N_10411,N_10642);
nand U13451 (N_13451,N_10417,N_11693);
and U13452 (N_13452,N_10031,N_10986);
nand U13453 (N_13453,N_11188,N_11844);
nand U13454 (N_13454,N_10558,N_10089);
nand U13455 (N_13455,N_10951,N_11622);
nand U13456 (N_13456,N_10815,N_11989);
and U13457 (N_13457,N_10581,N_10568);
nand U13458 (N_13458,N_10615,N_11564);
or U13459 (N_13459,N_10444,N_10450);
nand U13460 (N_13460,N_10267,N_10075);
nor U13461 (N_13461,N_11355,N_10746);
nor U13462 (N_13462,N_11685,N_10473);
nand U13463 (N_13463,N_11158,N_11624);
or U13464 (N_13464,N_10627,N_10506);
or U13465 (N_13465,N_10835,N_11926);
or U13466 (N_13466,N_11957,N_10672);
and U13467 (N_13467,N_11758,N_10384);
and U13468 (N_13468,N_10207,N_11235);
or U13469 (N_13469,N_10817,N_10355);
xor U13470 (N_13470,N_11279,N_11810);
or U13471 (N_13471,N_11215,N_10343);
xor U13472 (N_13472,N_11155,N_10947);
or U13473 (N_13473,N_10062,N_10151);
nand U13474 (N_13474,N_11458,N_11369);
and U13475 (N_13475,N_10283,N_11850);
and U13476 (N_13476,N_10407,N_11167);
or U13477 (N_13477,N_11680,N_10466);
nor U13478 (N_13478,N_10392,N_11770);
nand U13479 (N_13479,N_10195,N_11022);
nor U13480 (N_13480,N_10172,N_11053);
nor U13481 (N_13481,N_10069,N_10515);
or U13482 (N_13482,N_10586,N_11763);
and U13483 (N_13483,N_11639,N_10546);
and U13484 (N_13484,N_10005,N_11961);
nor U13485 (N_13485,N_10182,N_11020);
or U13486 (N_13486,N_10441,N_11992);
or U13487 (N_13487,N_10029,N_10795);
or U13488 (N_13488,N_10272,N_10789);
or U13489 (N_13489,N_11051,N_10840);
or U13490 (N_13490,N_10942,N_10548);
nand U13491 (N_13491,N_11144,N_10999);
nand U13492 (N_13492,N_11784,N_10324);
and U13493 (N_13493,N_11346,N_10492);
or U13494 (N_13494,N_11145,N_10879);
or U13495 (N_13495,N_10712,N_11013);
nor U13496 (N_13496,N_11433,N_10549);
and U13497 (N_13497,N_11092,N_10338);
or U13498 (N_13498,N_10037,N_11621);
nor U13499 (N_13499,N_10739,N_10650);
nand U13500 (N_13500,N_11642,N_10833);
nor U13501 (N_13501,N_11578,N_11839);
xnor U13502 (N_13502,N_10431,N_10868);
or U13503 (N_13503,N_10342,N_10526);
or U13504 (N_13504,N_11606,N_11439);
nand U13505 (N_13505,N_10299,N_10802);
nand U13506 (N_13506,N_10004,N_11106);
or U13507 (N_13507,N_11804,N_10439);
and U13508 (N_13508,N_10551,N_10207);
and U13509 (N_13509,N_11541,N_11213);
and U13510 (N_13510,N_11364,N_11624);
xnor U13511 (N_13511,N_11740,N_10909);
and U13512 (N_13512,N_10737,N_11926);
or U13513 (N_13513,N_11731,N_11065);
xor U13514 (N_13514,N_10827,N_11839);
nor U13515 (N_13515,N_11971,N_11744);
nor U13516 (N_13516,N_10114,N_10966);
or U13517 (N_13517,N_11918,N_11368);
nand U13518 (N_13518,N_11759,N_10888);
nor U13519 (N_13519,N_10664,N_10033);
nor U13520 (N_13520,N_11116,N_11647);
nand U13521 (N_13521,N_11958,N_11458);
nand U13522 (N_13522,N_10409,N_10675);
nand U13523 (N_13523,N_11159,N_11799);
and U13524 (N_13524,N_10663,N_10027);
nand U13525 (N_13525,N_11361,N_11488);
nand U13526 (N_13526,N_10868,N_11798);
xnor U13527 (N_13527,N_11173,N_11311);
nand U13528 (N_13528,N_10071,N_10805);
and U13529 (N_13529,N_10499,N_10791);
or U13530 (N_13530,N_11088,N_10284);
xor U13531 (N_13531,N_11744,N_10598);
nand U13532 (N_13532,N_11103,N_10361);
and U13533 (N_13533,N_11973,N_11810);
nor U13534 (N_13534,N_11065,N_11348);
or U13535 (N_13535,N_10199,N_10940);
nand U13536 (N_13536,N_10419,N_10846);
nor U13537 (N_13537,N_10336,N_10374);
xor U13538 (N_13538,N_11600,N_10532);
nor U13539 (N_13539,N_11365,N_10866);
and U13540 (N_13540,N_11835,N_11061);
and U13541 (N_13541,N_10570,N_10949);
or U13542 (N_13542,N_11945,N_11610);
or U13543 (N_13543,N_11033,N_10327);
and U13544 (N_13544,N_11531,N_11185);
and U13545 (N_13545,N_11130,N_10135);
nor U13546 (N_13546,N_11589,N_11381);
and U13547 (N_13547,N_11710,N_11852);
or U13548 (N_13548,N_11796,N_10895);
and U13549 (N_13549,N_11013,N_11091);
or U13550 (N_13550,N_11187,N_10395);
or U13551 (N_13551,N_10624,N_11179);
nand U13552 (N_13552,N_11009,N_10113);
nor U13553 (N_13553,N_10762,N_11031);
nand U13554 (N_13554,N_10599,N_10211);
nor U13555 (N_13555,N_10682,N_11811);
nor U13556 (N_13556,N_10162,N_11302);
nor U13557 (N_13557,N_10833,N_11164);
xor U13558 (N_13558,N_11932,N_11656);
or U13559 (N_13559,N_10880,N_11192);
nor U13560 (N_13560,N_10534,N_10744);
nor U13561 (N_13561,N_10155,N_10370);
and U13562 (N_13562,N_10798,N_10643);
or U13563 (N_13563,N_10499,N_11322);
nand U13564 (N_13564,N_10561,N_10644);
nor U13565 (N_13565,N_10964,N_11684);
or U13566 (N_13566,N_11303,N_11197);
nand U13567 (N_13567,N_11936,N_10455);
and U13568 (N_13568,N_10768,N_10277);
or U13569 (N_13569,N_10806,N_11986);
or U13570 (N_13570,N_11943,N_10185);
nand U13571 (N_13571,N_10078,N_11679);
nand U13572 (N_13572,N_11135,N_11741);
nand U13573 (N_13573,N_10861,N_10159);
or U13574 (N_13574,N_11354,N_10984);
xor U13575 (N_13575,N_10637,N_10061);
and U13576 (N_13576,N_11196,N_10669);
nand U13577 (N_13577,N_10008,N_10262);
nor U13578 (N_13578,N_10293,N_11220);
nand U13579 (N_13579,N_11609,N_10258);
and U13580 (N_13580,N_10795,N_10958);
nor U13581 (N_13581,N_11140,N_11543);
or U13582 (N_13582,N_11542,N_11467);
nand U13583 (N_13583,N_11131,N_10709);
nand U13584 (N_13584,N_11467,N_11199);
nor U13585 (N_13585,N_11559,N_10393);
or U13586 (N_13586,N_11399,N_10018);
and U13587 (N_13587,N_10435,N_11561);
or U13588 (N_13588,N_11922,N_11837);
or U13589 (N_13589,N_11932,N_10685);
or U13590 (N_13590,N_10277,N_11481);
nand U13591 (N_13591,N_11918,N_10950);
nand U13592 (N_13592,N_11572,N_10370);
or U13593 (N_13593,N_10191,N_11119);
nor U13594 (N_13594,N_10953,N_10532);
nand U13595 (N_13595,N_11523,N_11869);
nor U13596 (N_13596,N_11542,N_11364);
xnor U13597 (N_13597,N_10712,N_11069);
or U13598 (N_13598,N_10191,N_11642);
nand U13599 (N_13599,N_11577,N_10463);
or U13600 (N_13600,N_10385,N_11555);
or U13601 (N_13601,N_11821,N_11510);
and U13602 (N_13602,N_10162,N_10041);
or U13603 (N_13603,N_10503,N_10559);
xnor U13604 (N_13604,N_11393,N_11483);
xnor U13605 (N_13605,N_11053,N_11626);
nand U13606 (N_13606,N_11140,N_10885);
and U13607 (N_13607,N_11491,N_11114);
or U13608 (N_13608,N_10991,N_10742);
nand U13609 (N_13609,N_11035,N_11495);
nor U13610 (N_13610,N_11115,N_10649);
xor U13611 (N_13611,N_11838,N_10418);
or U13612 (N_13612,N_11090,N_10692);
xnor U13613 (N_13613,N_11529,N_11947);
nand U13614 (N_13614,N_10490,N_11092);
and U13615 (N_13615,N_11178,N_11336);
and U13616 (N_13616,N_10127,N_11436);
and U13617 (N_13617,N_11885,N_11173);
xnor U13618 (N_13618,N_11608,N_11532);
nand U13619 (N_13619,N_11098,N_10146);
nor U13620 (N_13620,N_10619,N_11181);
or U13621 (N_13621,N_11078,N_11761);
and U13622 (N_13622,N_10417,N_10830);
or U13623 (N_13623,N_10657,N_10555);
xnor U13624 (N_13624,N_11587,N_10649);
and U13625 (N_13625,N_10642,N_10638);
nand U13626 (N_13626,N_11211,N_10995);
xor U13627 (N_13627,N_11293,N_11584);
and U13628 (N_13628,N_10337,N_11514);
nand U13629 (N_13629,N_10089,N_11247);
or U13630 (N_13630,N_11015,N_11688);
or U13631 (N_13631,N_11192,N_10777);
xor U13632 (N_13632,N_11310,N_10155);
and U13633 (N_13633,N_11796,N_10674);
and U13634 (N_13634,N_11810,N_11614);
and U13635 (N_13635,N_11194,N_10365);
nand U13636 (N_13636,N_11012,N_11349);
nand U13637 (N_13637,N_10568,N_10637);
nand U13638 (N_13638,N_11834,N_11060);
nor U13639 (N_13639,N_10102,N_11517);
and U13640 (N_13640,N_11131,N_11343);
or U13641 (N_13641,N_11918,N_11756);
or U13642 (N_13642,N_10097,N_11589);
or U13643 (N_13643,N_11670,N_11934);
or U13644 (N_13644,N_10607,N_10152);
xor U13645 (N_13645,N_10874,N_11159);
and U13646 (N_13646,N_11700,N_11413);
nor U13647 (N_13647,N_11597,N_11715);
or U13648 (N_13648,N_11322,N_10338);
and U13649 (N_13649,N_10875,N_11627);
nand U13650 (N_13650,N_10545,N_11613);
nand U13651 (N_13651,N_11876,N_10623);
or U13652 (N_13652,N_10993,N_10877);
and U13653 (N_13653,N_11464,N_10381);
or U13654 (N_13654,N_11348,N_10772);
or U13655 (N_13655,N_10570,N_10343);
xnor U13656 (N_13656,N_10479,N_11182);
or U13657 (N_13657,N_11263,N_10542);
or U13658 (N_13658,N_11395,N_10519);
xnor U13659 (N_13659,N_10096,N_10043);
nor U13660 (N_13660,N_11312,N_11760);
nor U13661 (N_13661,N_10490,N_10889);
or U13662 (N_13662,N_11364,N_11086);
nor U13663 (N_13663,N_11410,N_11694);
nand U13664 (N_13664,N_10344,N_10879);
and U13665 (N_13665,N_10623,N_10284);
and U13666 (N_13666,N_10227,N_10707);
nor U13667 (N_13667,N_11466,N_11652);
nand U13668 (N_13668,N_11214,N_10868);
nor U13669 (N_13669,N_11649,N_11749);
nand U13670 (N_13670,N_10111,N_10374);
nor U13671 (N_13671,N_11521,N_10232);
and U13672 (N_13672,N_11921,N_11216);
nand U13673 (N_13673,N_11809,N_11016);
and U13674 (N_13674,N_11496,N_11021);
and U13675 (N_13675,N_10757,N_11650);
nor U13676 (N_13676,N_11236,N_11997);
nor U13677 (N_13677,N_10385,N_11348);
nor U13678 (N_13678,N_10762,N_10088);
nor U13679 (N_13679,N_10367,N_10317);
xor U13680 (N_13680,N_11864,N_11358);
xnor U13681 (N_13681,N_10481,N_11667);
nand U13682 (N_13682,N_10298,N_10505);
nor U13683 (N_13683,N_10817,N_10526);
or U13684 (N_13684,N_11352,N_11654);
or U13685 (N_13685,N_10764,N_11153);
and U13686 (N_13686,N_11552,N_10589);
and U13687 (N_13687,N_11769,N_10701);
nor U13688 (N_13688,N_10507,N_11622);
nor U13689 (N_13689,N_10238,N_10941);
xnor U13690 (N_13690,N_10918,N_10203);
nand U13691 (N_13691,N_11464,N_11336);
or U13692 (N_13692,N_11633,N_11436);
and U13693 (N_13693,N_11985,N_10645);
nand U13694 (N_13694,N_11059,N_11071);
and U13695 (N_13695,N_10321,N_11985);
nor U13696 (N_13696,N_11564,N_10448);
xnor U13697 (N_13697,N_11103,N_11934);
and U13698 (N_13698,N_11897,N_11530);
xor U13699 (N_13699,N_10892,N_10928);
nor U13700 (N_13700,N_11117,N_10019);
nand U13701 (N_13701,N_10486,N_10287);
and U13702 (N_13702,N_10984,N_11201);
nor U13703 (N_13703,N_11610,N_10981);
and U13704 (N_13704,N_11443,N_10366);
nor U13705 (N_13705,N_11305,N_10596);
nand U13706 (N_13706,N_10823,N_10963);
nor U13707 (N_13707,N_10242,N_11715);
or U13708 (N_13708,N_11012,N_10847);
nand U13709 (N_13709,N_10478,N_10851);
nand U13710 (N_13710,N_10207,N_11591);
and U13711 (N_13711,N_10678,N_11020);
nand U13712 (N_13712,N_11865,N_11633);
and U13713 (N_13713,N_11436,N_11988);
xnor U13714 (N_13714,N_10876,N_11018);
or U13715 (N_13715,N_11882,N_10189);
nand U13716 (N_13716,N_11592,N_11216);
nand U13717 (N_13717,N_11416,N_10231);
xnor U13718 (N_13718,N_10930,N_10403);
nand U13719 (N_13719,N_10963,N_11160);
xor U13720 (N_13720,N_10511,N_10292);
nor U13721 (N_13721,N_11126,N_10096);
nand U13722 (N_13722,N_11940,N_11112);
nor U13723 (N_13723,N_11096,N_10998);
and U13724 (N_13724,N_10598,N_10899);
xnor U13725 (N_13725,N_10812,N_11856);
or U13726 (N_13726,N_10690,N_10483);
and U13727 (N_13727,N_11730,N_11721);
or U13728 (N_13728,N_11993,N_11534);
or U13729 (N_13729,N_10391,N_10854);
nand U13730 (N_13730,N_10012,N_10364);
and U13731 (N_13731,N_11337,N_10031);
or U13732 (N_13732,N_11750,N_11881);
nand U13733 (N_13733,N_10614,N_10492);
or U13734 (N_13734,N_10538,N_10448);
and U13735 (N_13735,N_11793,N_10343);
xnor U13736 (N_13736,N_11101,N_10825);
nand U13737 (N_13737,N_10517,N_11494);
and U13738 (N_13738,N_10564,N_10360);
and U13739 (N_13739,N_11641,N_10505);
nor U13740 (N_13740,N_11392,N_10806);
and U13741 (N_13741,N_11186,N_11541);
and U13742 (N_13742,N_11171,N_11669);
nor U13743 (N_13743,N_11675,N_11330);
and U13744 (N_13744,N_10762,N_10554);
nor U13745 (N_13745,N_10052,N_11553);
nand U13746 (N_13746,N_10105,N_11197);
and U13747 (N_13747,N_11869,N_11410);
nor U13748 (N_13748,N_11171,N_10844);
nor U13749 (N_13749,N_11172,N_10012);
or U13750 (N_13750,N_11860,N_10589);
nand U13751 (N_13751,N_10815,N_11293);
nor U13752 (N_13752,N_10167,N_10866);
nand U13753 (N_13753,N_10419,N_11412);
xnor U13754 (N_13754,N_10169,N_10176);
and U13755 (N_13755,N_11290,N_10464);
and U13756 (N_13756,N_10619,N_11268);
and U13757 (N_13757,N_11889,N_10809);
and U13758 (N_13758,N_11675,N_11565);
or U13759 (N_13759,N_11510,N_10717);
or U13760 (N_13760,N_11478,N_11075);
and U13761 (N_13761,N_11747,N_11728);
nor U13762 (N_13762,N_11240,N_11047);
nand U13763 (N_13763,N_11949,N_10389);
nand U13764 (N_13764,N_11566,N_11616);
and U13765 (N_13765,N_11152,N_11300);
nand U13766 (N_13766,N_11387,N_10268);
and U13767 (N_13767,N_11989,N_11440);
or U13768 (N_13768,N_10428,N_10321);
or U13769 (N_13769,N_11643,N_11833);
or U13770 (N_13770,N_11451,N_10541);
or U13771 (N_13771,N_11021,N_10983);
xor U13772 (N_13772,N_10057,N_10663);
or U13773 (N_13773,N_11036,N_10262);
nand U13774 (N_13774,N_10002,N_11780);
nor U13775 (N_13775,N_11052,N_10356);
and U13776 (N_13776,N_10289,N_11951);
nor U13777 (N_13777,N_11063,N_11932);
nand U13778 (N_13778,N_10715,N_11609);
or U13779 (N_13779,N_10092,N_10764);
xnor U13780 (N_13780,N_10581,N_10912);
and U13781 (N_13781,N_11961,N_10454);
xor U13782 (N_13782,N_10112,N_11104);
and U13783 (N_13783,N_11832,N_11738);
nor U13784 (N_13784,N_10790,N_11710);
nor U13785 (N_13785,N_11991,N_10448);
nand U13786 (N_13786,N_11339,N_10838);
and U13787 (N_13787,N_10820,N_11359);
nor U13788 (N_13788,N_10425,N_10071);
and U13789 (N_13789,N_11522,N_10898);
nor U13790 (N_13790,N_10622,N_10737);
and U13791 (N_13791,N_10147,N_10415);
nor U13792 (N_13792,N_10862,N_10369);
nand U13793 (N_13793,N_11926,N_11043);
nor U13794 (N_13794,N_11434,N_10123);
or U13795 (N_13795,N_11762,N_11658);
nor U13796 (N_13796,N_11562,N_11935);
and U13797 (N_13797,N_11906,N_11759);
nand U13798 (N_13798,N_11364,N_10225);
nand U13799 (N_13799,N_10154,N_10445);
nor U13800 (N_13800,N_10774,N_10538);
xor U13801 (N_13801,N_11201,N_10811);
or U13802 (N_13802,N_10837,N_10433);
and U13803 (N_13803,N_11301,N_11275);
or U13804 (N_13804,N_11711,N_10382);
xnor U13805 (N_13805,N_10593,N_11921);
or U13806 (N_13806,N_11138,N_11438);
or U13807 (N_13807,N_11024,N_10803);
or U13808 (N_13808,N_10373,N_11026);
or U13809 (N_13809,N_10248,N_11313);
and U13810 (N_13810,N_11430,N_10344);
nor U13811 (N_13811,N_11252,N_10745);
nand U13812 (N_13812,N_10730,N_10539);
and U13813 (N_13813,N_11451,N_11538);
nand U13814 (N_13814,N_10589,N_11763);
nand U13815 (N_13815,N_10168,N_11574);
and U13816 (N_13816,N_11051,N_11968);
nor U13817 (N_13817,N_10849,N_11444);
nand U13818 (N_13818,N_11221,N_10321);
nor U13819 (N_13819,N_10895,N_10699);
and U13820 (N_13820,N_11037,N_10437);
nand U13821 (N_13821,N_10603,N_10887);
nor U13822 (N_13822,N_11002,N_10826);
nand U13823 (N_13823,N_11869,N_11717);
nand U13824 (N_13824,N_10435,N_11387);
or U13825 (N_13825,N_11063,N_10497);
xnor U13826 (N_13826,N_11924,N_11296);
nand U13827 (N_13827,N_11840,N_10497);
nand U13828 (N_13828,N_10357,N_11878);
nor U13829 (N_13829,N_11379,N_11650);
and U13830 (N_13830,N_10616,N_11192);
and U13831 (N_13831,N_10652,N_10881);
or U13832 (N_13832,N_11865,N_10146);
xor U13833 (N_13833,N_10808,N_11448);
nand U13834 (N_13834,N_10851,N_11407);
nand U13835 (N_13835,N_10980,N_10237);
and U13836 (N_13836,N_11654,N_10795);
xnor U13837 (N_13837,N_10877,N_10431);
nand U13838 (N_13838,N_10422,N_11022);
and U13839 (N_13839,N_11246,N_10739);
nor U13840 (N_13840,N_10540,N_10508);
nor U13841 (N_13841,N_11145,N_11472);
nand U13842 (N_13842,N_10143,N_11946);
or U13843 (N_13843,N_11310,N_11981);
nor U13844 (N_13844,N_10483,N_10034);
nor U13845 (N_13845,N_10517,N_10116);
and U13846 (N_13846,N_10213,N_11534);
or U13847 (N_13847,N_11532,N_10266);
and U13848 (N_13848,N_10839,N_11503);
or U13849 (N_13849,N_11952,N_11587);
and U13850 (N_13850,N_11964,N_11227);
and U13851 (N_13851,N_10923,N_11773);
nand U13852 (N_13852,N_11774,N_11305);
nand U13853 (N_13853,N_10783,N_10330);
or U13854 (N_13854,N_10080,N_10006);
xnor U13855 (N_13855,N_11849,N_10243);
xor U13856 (N_13856,N_11172,N_11631);
xor U13857 (N_13857,N_11189,N_10482);
or U13858 (N_13858,N_10338,N_11054);
or U13859 (N_13859,N_10891,N_11333);
nand U13860 (N_13860,N_10609,N_11911);
nand U13861 (N_13861,N_11794,N_11909);
nor U13862 (N_13862,N_11082,N_11869);
and U13863 (N_13863,N_10555,N_10378);
and U13864 (N_13864,N_10112,N_11113);
nor U13865 (N_13865,N_10951,N_10655);
xnor U13866 (N_13866,N_10752,N_10385);
nor U13867 (N_13867,N_10705,N_10287);
nor U13868 (N_13868,N_11973,N_11415);
or U13869 (N_13869,N_10762,N_10108);
nor U13870 (N_13870,N_10422,N_11351);
nor U13871 (N_13871,N_10103,N_10773);
nand U13872 (N_13872,N_10919,N_10385);
nor U13873 (N_13873,N_10151,N_10965);
or U13874 (N_13874,N_11463,N_10975);
nand U13875 (N_13875,N_10182,N_11302);
or U13876 (N_13876,N_11821,N_10965);
xnor U13877 (N_13877,N_11910,N_10840);
or U13878 (N_13878,N_10495,N_11776);
xnor U13879 (N_13879,N_11836,N_11569);
nand U13880 (N_13880,N_11299,N_10061);
nand U13881 (N_13881,N_11352,N_11790);
or U13882 (N_13882,N_10819,N_10351);
and U13883 (N_13883,N_11931,N_11471);
nor U13884 (N_13884,N_10879,N_10097);
nor U13885 (N_13885,N_11984,N_11759);
nor U13886 (N_13886,N_10315,N_10032);
nand U13887 (N_13887,N_10490,N_10691);
and U13888 (N_13888,N_11514,N_10150);
nand U13889 (N_13889,N_11511,N_11893);
and U13890 (N_13890,N_10636,N_11617);
or U13891 (N_13891,N_11932,N_10428);
nand U13892 (N_13892,N_10314,N_11164);
nor U13893 (N_13893,N_10639,N_10191);
or U13894 (N_13894,N_10021,N_10955);
nor U13895 (N_13895,N_11415,N_11915);
nand U13896 (N_13896,N_11325,N_10687);
nor U13897 (N_13897,N_11524,N_11476);
xnor U13898 (N_13898,N_10522,N_10573);
or U13899 (N_13899,N_10806,N_11100);
xor U13900 (N_13900,N_10785,N_10228);
or U13901 (N_13901,N_11466,N_11797);
or U13902 (N_13902,N_11820,N_11253);
nand U13903 (N_13903,N_10894,N_11678);
or U13904 (N_13904,N_10982,N_10736);
or U13905 (N_13905,N_10198,N_11840);
or U13906 (N_13906,N_10536,N_11478);
nand U13907 (N_13907,N_10373,N_10125);
nor U13908 (N_13908,N_11634,N_10473);
or U13909 (N_13909,N_11614,N_11313);
nor U13910 (N_13910,N_10391,N_11174);
or U13911 (N_13911,N_11315,N_11250);
and U13912 (N_13912,N_11175,N_11523);
and U13913 (N_13913,N_11370,N_11801);
nand U13914 (N_13914,N_11834,N_10173);
or U13915 (N_13915,N_11409,N_11229);
or U13916 (N_13916,N_10999,N_11186);
nor U13917 (N_13917,N_11723,N_11443);
nand U13918 (N_13918,N_10672,N_11031);
or U13919 (N_13919,N_10905,N_10146);
nand U13920 (N_13920,N_11344,N_11612);
nor U13921 (N_13921,N_10507,N_10891);
nand U13922 (N_13922,N_11054,N_11994);
and U13923 (N_13923,N_11951,N_10852);
nor U13924 (N_13924,N_10448,N_10064);
nor U13925 (N_13925,N_11204,N_11349);
and U13926 (N_13926,N_11753,N_11322);
or U13927 (N_13927,N_11166,N_11639);
or U13928 (N_13928,N_11773,N_11971);
xor U13929 (N_13929,N_11979,N_11096);
and U13930 (N_13930,N_11477,N_10622);
and U13931 (N_13931,N_11005,N_10887);
nand U13932 (N_13932,N_10009,N_10765);
nand U13933 (N_13933,N_10498,N_11951);
or U13934 (N_13934,N_11106,N_10345);
nor U13935 (N_13935,N_10309,N_11910);
and U13936 (N_13936,N_11498,N_10476);
or U13937 (N_13937,N_10296,N_11050);
xor U13938 (N_13938,N_10718,N_10019);
nand U13939 (N_13939,N_11007,N_10004);
nor U13940 (N_13940,N_11532,N_11442);
nor U13941 (N_13941,N_11030,N_11358);
or U13942 (N_13942,N_11303,N_10136);
nand U13943 (N_13943,N_11531,N_11730);
nor U13944 (N_13944,N_11377,N_11863);
nand U13945 (N_13945,N_11719,N_10844);
or U13946 (N_13946,N_11605,N_10888);
or U13947 (N_13947,N_11942,N_10988);
nor U13948 (N_13948,N_10717,N_10123);
xnor U13949 (N_13949,N_11246,N_11127);
nand U13950 (N_13950,N_11572,N_11126);
nand U13951 (N_13951,N_10257,N_11480);
or U13952 (N_13952,N_11590,N_10635);
nor U13953 (N_13953,N_10701,N_11226);
and U13954 (N_13954,N_11303,N_11446);
nand U13955 (N_13955,N_11767,N_10734);
or U13956 (N_13956,N_11542,N_11079);
nor U13957 (N_13957,N_11079,N_11424);
or U13958 (N_13958,N_10265,N_11398);
nor U13959 (N_13959,N_10915,N_11487);
or U13960 (N_13960,N_10116,N_11840);
and U13961 (N_13961,N_10547,N_10608);
nand U13962 (N_13962,N_11030,N_10924);
or U13963 (N_13963,N_10326,N_10316);
and U13964 (N_13964,N_10103,N_11490);
nand U13965 (N_13965,N_10377,N_11181);
and U13966 (N_13966,N_10628,N_11494);
nand U13967 (N_13967,N_11266,N_10260);
nor U13968 (N_13968,N_10080,N_11661);
or U13969 (N_13969,N_10373,N_11989);
or U13970 (N_13970,N_10002,N_10091);
or U13971 (N_13971,N_10352,N_10467);
or U13972 (N_13972,N_11959,N_11774);
or U13973 (N_13973,N_10502,N_10687);
or U13974 (N_13974,N_11580,N_10963);
nand U13975 (N_13975,N_11123,N_10320);
nor U13976 (N_13976,N_10119,N_11423);
or U13977 (N_13977,N_10775,N_11621);
nand U13978 (N_13978,N_10667,N_10958);
nor U13979 (N_13979,N_10193,N_11610);
nand U13980 (N_13980,N_10269,N_10397);
nor U13981 (N_13981,N_10496,N_11140);
or U13982 (N_13982,N_10279,N_10157);
nand U13983 (N_13983,N_10542,N_10504);
nor U13984 (N_13984,N_11413,N_11204);
and U13985 (N_13985,N_11149,N_11013);
nand U13986 (N_13986,N_10059,N_11346);
and U13987 (N_13987,N_11045,N_11613);
or U13988 (N_13988,N_10086,N_10321);
nor U13989 (N_13989,N_11979,N_11502);
or U13990 (N_13990,N_10747,N_11005);
nor U13991 (N_13991,N_10817,N_10100);
xor U13992 (N_13992,N_10465,N_10227);
or U13993 (N_13993,N_10651,N_11607);
nor U13994 (N_13994,N_10394,N_11162);
nand U13995 (N_13995,N_10944,N_11554);
xnor U13996 (N_13996,N_10816,N_10188);
nand U13997 (N_13997,N_10150,N_10325);
or U13998 (N_13998,N_11048,N_10986);
nand U13999 (N_13999,N_11159,N_10620);
or U14000 (N_14000,N_13470,N_13297);
nor U14001 (N_14001,N_13747,N_13525);
nor U14002 (N_14002,N_13983,N_12706);
and U14003 (N_14003,N_12058,N_13932);
nor U14004 (N_14004,N_13440,N_13799);
or U14005 (N_14005,N_12890,N_13516);
nand U14006 (N_14006,N_12402,N_12632);
and U14007 (N_14007,N_12611,N_13284);
and U14008 (N_14008,N_13679,N_13328);
nand U14009 (N_14009,N_12384,N_12283);
or U14010 (N_14010,N_12392,N_12715);
nand U14011 (N_14011,N_12489,N_12593);
and U14012 (N_14012,N_13064,N_13999);
nand U14013 (N_14013,N_12996,N_13864);
nand U14014 (N_14014,N_13500,N_12792);
nor U14015 (N_14015,N_12955,N_12126);
and U14016 (N_14016,N_13019,N_12147);
or U14017 (N_14017,N_13131,N_12563);
nor U14018 (N_14018,N_13826,N_12021);
nand U14019 (N_14019,N_12139,N_12301);
nor U14020 (N_14020,N_13503,N_13234);
nand U14021 (N_14021,N_12666,N_13363);
nand U14022 (N_14022,N_13740,N_13242);
and U14023 (N_14023,N_13785,N_13137);
nor U14024 (N_14024,N_13406,N_12461);
and U14025 (N_14025,N_13955,N_13190);
or U14026 (N_14026,N_12808,N_12032);
nor U14027 (N_14027,N_12754,N_12149);
nand U14028 (N_14028,N_12709,N_13228);
and U14029 (N_14029,N_12441,N_13385);
xnor U14030 (N_14030,N_13578,N_12339);
or U14031 (N_14031,N_12500,N_12958);
nor U14032 (N_14032,N_13038,N_12068);
xor U14033 (N_14033,N_13293,N_13037);
or U14034 (N_14034,N_13984,N_13023);
and U14035 (N_14035,N_13399,N_12663);
and U14036 (N_14036,N_13791,N_12986);
nand U14037 (N_14037,N_13689,N_13353);
nand U14038 (N_14038,N_13295,N_13752);
nand U14039 (N_14039,N_13255,N_12214);
nand U14040 (N_14040,N_12991,N_13236);
nor U14041 (N_14041,N_12901,N_12553);
and U14042 (N_14042,N_13584,N_12687);
nor U14043 (N_14043,N_13445,N_12420);
and U14044 (N_14044,N_13271,N_13910);
and U14045 (N_14045,N_12667,N_13370);
xnor U14046 (N_14046,N_13581,N_13960);
nand U14047 (N_14047,N_12195,N_13104);
nand U14048 (N_14048,N_12286,N_12485);
or U14049 (N_14049,N_12790,N_13311);
nand U14050 (N_14050,N_12970,N_13648);
or U14051 (N_14051,N_13152,N_12132);
or U14052 (N_14052,N_13178,N_12721);
nand U14053 (N_14053,N_12226,N_12730);
xor U14054 (N_14054,N_12848,N_12377);
and U14055 (N_14055,N_12580,N_12004);
nor U14056 (N_14056,N_13382,N_13062);
or U14057 (N_14057,N_13036,N_12560);
and U14058 (N_14058,N_13527,N_12151);
nand U14059 (N_14059,N_13303,N_12934);
or U14060 (N_14060,N_13354,N_13582);
and U14061 (N_14061,N_13246,N_12293);
or U14062 (N_14062,N_12654,N_12192);
nand U14063 (N_14063,N_13260,N_13014);
and U14064 (N_14064,N_13274,N_12840);
or U14065 (N_14065,N_13823,N_12146);
nand U14066 (N_14066,N_13788,N_12207);
or U14067 (N_14067,N_13034,N_12902);
or U14068 (N_14068,N_13216,N_12024);
nand U14069 (N_14069,N_13229,N_12087);
and U14070 (N_14070,N_12354,N_13640);
or U14071 (N_14071,N_13737,N_13951);
nand U14072 (N_14072,N_13085,N_12127);
and U14073 (N_14073,N_12271,N_13974);
and U14074 (N_14074,N_13868,N_13614);
and U14075 (N_14075,N_12287,N_12400);
or U14076 (N_14076,N_13549,N_12622);
and U14077 (N_14077,N_12887,N_12874);
and U14078 (N_14078,N_13817,N_12152);
and U14079 (N_14079,N_13753,N_12397);
or U14080 (N_14080,N_13298,N_13941);
nor U14081 (N_14081,N_13646,N_12007);
nor U14082 (N_14082,N_12182,N_12279);
nor U14083 (N_14083,N_12569,N_13644);
nand U14084 (N_14084,N_13025,N_13774);
and U14085 (N_14085,N_13082,N_12717);
nor U14086 (N_14086,N_13781,N_13600);
and U14087 (N_14087,N_12265,N_12871);
nor U14088 (N_14088,N_12559,N_12819);
xnor U14089 (N_14089,N_13800,N_12741);
nor U14090 (N_14090,N_12575,N_13147);
or U14091 (N_14091,N_13869,N_12909);
or U14092 (N_14092,N_12398,N_13334);
nand U14093 (N_14093,N_12117,N_12690);
or U14094 (N_14094,N_12346,N_13724);
nor U14095 (N_14095,N_12948,N_12777);
or U14096 (N_14096,N_12734,N_12409);
nand U14097 (N_14097,N_12046,N_12325);
and U14098 (N_14098,N_12637,N_12048);
nor U14099 (N_14099,N_12743,N_12401);
nand U14100 (N_14100,N_13453,N_13667);
nand U14101 (N_14101,N_12495,N_12655);
and U14102 (N_14102,N_13562,N_13077);
xor U14103 (N_14103,N_12618,N_12203);
nor U14104 (N_14104,N_12491,N_13009);
or U14105 (N_14105,N_13623,N_12793);
or U14106 (N_14106,N_12482,N_12361);
and U14107 (N_14107,N_13565,N_12037);
and U14108 (N_14108,N_13043,N_12445);
nand U14109 (N_14109,N_13890,N_13498);
nor U14110 (N_14110,N_12988,N_13267);
nor U14111 (N_14111,N_12221,N_13163);
and U14112 (N_14112,N_13276,N_12903);
xor U14113 (N_14113,N_13030,N_13931);
or U14114 (N_14114,N_13074,N_13059);
nand U14115 (N_14115,N_13844,N_12710);
xnor U14116 (N_14116,N_13249,N_12538);
nor U14117 (N_14117,N_13031,N_12699);
nand U14118 (N_14118,N_13764,N_12638);
nand U14119 (N_14119,N_12814,N_13843);
or U14120 (N_14120,N_13994,N_13111);
or U14121 (N_14121,N_12052,N_12012);
nor U14122 (N_14122,N_12408,N_13365);
nor U14123 (N_14123,N_12344,N_13547);
nand U14124 (N_14124,N_13192,N_13292);
nor U14125 (N_14125,N_13911,N_13656);
and U14126 (N_14126,N_12382,N_12574);
xor U14127 (N_14127,N_12025,N_12413);
nand U14128 (N_14128,N_13548,N_12326);
nor U14129 (N_14129,N_12463,N_13758);
nand U14130 (N_14130,N_12103,N_12034);
xnor U14131 (N_14131,N_13005,N_12817);
and U14132 (N_14132,N_13641,N_13786);
nand U14133 (N_14133,N_13891,N_12291);
and U14134 (N_14134,N_13027,N_13842);
nand U14135 (N_14135,N_12171,N_12959);
and U14136 (N_14136,N_12650,N_12543);
and U14137 (N_14137,N_12360,N_12930);
and U14138 (N_14138,N_12086,N_13230);
and U14139 (N_14139,N_12143,N_12381);
and U14140 (N_14140,N_13324,N_13838);
nand U14141 (N_14141,N_12807,N_13596);
and U14142 (N_14142,N_12492,N_12515);
nand U14143 (N_14143,N_13712,N_12614);
and U14144 (N_14144,N_13322,N_12705);
or U14145 (N_14145,N_13150,N_13316);
nor U14146 (N_14146,N_13928,N_12477);
or U14147 (N_14147,N_12315,N_13155);
nor U14148 (N_14148,N_12573,N_12035);
or U14149 (N_14149,N_12349,N_13233);
nor U14150 (N_14150,N_12856,N_12732);
xor U14151 (N_14151,N_12904,N_13706);
and U14152 (N_14152,N_13405,N_12030);
nand U14153 (N_14153,N_13522,N_12765);
nand U14154 (N_14154,N_13134,N_12911);
nor U14155 (N_14155,N_13409,N_13946);
xor U14156 (N_14156,N_12850,N_13750);
nor U14157 (N_14157,N_13687,N_12177);
and U14158 (N_14158,N_12708,N_12141);
nand U14159 (N_14159,N_13921,N_13875);
nand U14160 (N_14160,N_13020,N_13815);
nor U14161 (N_14161,N_13472,N_13671);
and U14162 (N_14162,N_13375,N_13452);
nor U14163 (N_14163,N_13532,N_12334);
xor U14164 (N_14164,N_13502,N_13290);
and U14165 (N_14165,N_12205,N_13389);
xor U14166 (N_14166,N_12063,N_12078);
or U14167 (N_14167,N_12605,N_13579);
and U14168 (N_14168,N_13924,N_13078);
or U14169 (N_14169,N_13696,N_12648);
or U14170 (N_14170,N_13598,N_13165);
or U14171 (N_14171,N_13980,N_12936);
nor U14172 (N_14172,N_13431,N_13259);
or U14173 (N_14173,N_13092,N_12504);
and U14174 (N_14174,N_13917,N_13942);
and U14175 (N_14175,N_12855,N_12827);
nand U14176 (N_14176,N_13220,N_12125);
nand U14177 (N_14177,N_12093,N_13632);
or U14178 (N_14178,N_13203,N_13854);
nor U14179 (N_14179,N_12939,N_12649);
nand U14180 (N_14180,N_12308,N_12977);
nand U14181 (N_14181,N_13210,N_12506);
or U14182 (N_14182,N_13149,N_12832);
or U14183 (N_14183,N_13386,N_13438);
and U14184 (N_14184,N_12665,N_12115);
or U14185 (N_14185,N_13376,N_13849);
nand U14186 (N_14186,N_13506,N_13425);
nand U14187 (N_14187,N_12623,N_13168);
nand U14188 (N_14188,N_13148,N_13618);
and U14189 (N_14189,N_12825,N_13877);
nor U14190 (N_14190,N_13310,N_13110);
xnor U14191 (N_14191,N_13668,N_13746);
nand U14192 (N_14192,N_13585,N_13199);
nor U14193 (N_14193,N_12659,N_12130);
xor U14194 (N_14194,N_13902,N_13349);
nor U14195 (N_14195,N_13624,N_13546);
nand U14196 (N_14196,N_13238,N_13702);
or U14197 (N_14197,N_13021,N_12795);
nor U14198 (N_14198,N_12558,N_13279);
xnor U14199 (N_14199,N_13524,N_12222);
or U14200 (N_14200,N_13132,N_13734);
nand U14201 (N_14201,N_13167,N_13464);
nand U14202 (N_14202,N_12245,N_12042);
or U14203 (N_14203,N_12752,N_13308);
or U14204 (N_14204,N_13957,N_12277);
and U14205 (N_14205,N_13235,N_13559);
xnor U14206 (N_14206,N_12106,N_13639);
nor U14207 (N_14207,N_13839,N_12950);
and U14208 (N_14208,N_12036,N_13424);
and U14209 (N_14209,N_12641,N_12391);
or U14210 (N_14210,N_12739,N_12520);
and U14211 (N_14211,N_13627,N_12867);
nand U14212 (N_14212,N_12471,N_13088);
nand U14213 (N_14213,N_13364,N_13056);
or U14214 (N_14214,N_13756,N_13853);
nor U14215 (N_14215,N_12059,N_13248);
nor U14216 (N_14216,N_12260,N_13900);
and U14217 (N_14217,N_13244,N_12513);
and U14218 (N_14218,N_12439,N_13561);
and U14219 (N_14219,N_13697,N_12875);
nor U14220 (N_14220,N_13985,N_13465);
nor U14221 (N_14221,N_13934,N_12144);
and U14222 (N_14222,N_13554,N_13283);
or U14223 (N_14223,N_13612,N_13218);
or U14224 (N_14224,N_13926,N_12989);
and U14225 (N_14225,N_12418,N_12925);
and U14226 (N_14226,N_13176,N_12259);
xor U14227 (N_14227,N_12588,N_13556);
or U14228 (N_14228,N_13213,N_13987);
nand U14229 (N_14229,N_13492,N_12834);
and U14230 (N_14230,N_13589,N_12027);
or U14231 (N_14231,N_12707,N_12081);
xor U14232 (N_14232,N_13829,N_12133);
nor U14233 (N_14233,N_12180,N_12165);
or U14234 (N_14234,N_13380,N_13243);
nand U14235 (N_14235,N_12051,N_12138);
or U14236 (N_14236,N_12336,N_12497);
xor U14237 (N_14237,N_12862,N_13061);
nand U14238 (N_14238,N_13499,N_13908);
nand U14239 (N_14239,N_13903,N_12800);
and U14240 (N_14240,N_12586,N_12285);
and U14241 (N_14241,N_13675,N_13181);
or U14242 (N_14242,N_12280,N_13620);
and U14243 (N_14243,N_13378,N_12128);
or U14244 (N_14244,N_13509,N_13856);
nor U14245 (N_14245,N_13964,N_13265);
nand U14246 (N_14246,N_12744,N_13997);
nor U14247 (N_14247,N_13913,N_12483);
and U14248 (N_14248,N_12858,N_12072);
or U14249 (N_14249,N_13377,N_12778);
xor U14250 (N_14250,N_12969,N_12047);
nor U14251 (N_14251,N_13511,N_13571);
or U14252 (N_14252,N_13693,N_13227);
xnor U14253 (N_14253,N_12869,N_12829);
nor U14254 (N_14254,N_13266,N_13550);
nor U14255 (N_14255,N_12246,N_13143);
and U14256 (N_14256,N_12430,N_13262);
nand U14257 (N_14257,N_12425,N_13809);
nand U14258 (N_14258,N_12366,N_13277);
xnor U14259 (N_14259,N_12517,N_13806);
and U14260 (N_14260,N_12949,N_13824);
or U14261 (N_14261,N_13454,N_13179);
and U14262 (N_14262,N_12772,N_12374);
or U14263 (N_14263,N_12242,N_12179);
xnor U14264 (N_14264,N_12473,N_12906);
nor U14265 (N_14265,N_12505,N_13976);
nor U14266 (N_14266,N_12303,N_13615);
or U14267 (N_14267,N_13848,N_13374);
xor U14268 (N_14268,N_12818,N_12766);
and U14269 (N_14269,N_13003,N_13935);
xnor U14270 (N_14270,N_12241,N_13046);
or U14271 (N_14271,N_13886,N_13422);
or U14272 (N_14272,N_12444,N_12635);
nor U14273 (N_14273,N_13186,N_12561);
nor U14274 (N_14274,N_12446,N_13223);
or U14275 (N_14275,N_12175,N_12951);
nand U14276 (N_14276,N_13988,N_13760);
and U14277 (N_14277,N_13096,N_12940);
xor U14278 (N_14278,N_12692,N_12050);
nand U14279 (N_14279,N_13588,N_13771);
and U14280 (N_14280,N_12481,N_12161);
nand U14281 (N_14281,N_12597,N_12947);
nor U14282 (N_14282,N_13282,N_12116);
nand U14283 (N_14283,N_13742,N_13820);
or U14284 (N_14284,N_13950,N_13479);
nand U14285 (N_14285,N_12284,N_13075);
and U14286 (N_14286,N_13225,N_12987);
xor U14287 (N_14287,N_13494,N_13850);
nor U14288 (N_14288,N_12000,N_12900);
nand U14289 (N_14289,N_13807,N_13202);
or U14290 (N_14290,N_13072,N_12348);
and U14291 (N_14291,N_13156,N_12319);
nand U14292 (N_14292,N_13307,N_13501);
nand U14293 (N_14293,N_13125,N_13659);
and U14294 (N_14294,N_13810,N_12201);
or U14295 (N_14295,N_13531,N_12797);
or U14296 (N_14296,N_13718,N_13859);
nand U14297 (N_14297,N_13553,N_13677);
nand U14298 (N_14298,N_12095,N_13874);
or U14299 (N_14299,N_12262,N_13087);
and U14300 (N_14300,N_12544,N_13523);
or U14301 (N_14301,N_13154,N_12619);
nor U14302 (N_14302,N_12981,N_13049);
and U14303 (N_14303,N_12438,N_12337);
and U14304 (N_14304,N_12140,N_12256);
nand U14305 (N_14305,N_13631,N_12738);
and U14306 (N_14306,N_12521,N_13595);
nor U14307 (N_14307,N_13507,N_12548);
nor U14308 (N_14308,N_13312,N_12258);
nand U14309 (N_14309,N_13812,N_13684);
nand U14310 (N_14310,N_13183,N_12647);
nor U14311 (N_14311,N_12254,N_13775);
or U14312 (N_14312,N_12695,N_13899);
or U14313 (N_14313,N_12101,N_13306);
nor U14314 (N_14314,N_12314,N_12001);
and U14315 (N_14315,N_12672,N_13457);
or U14316 (N_14316,N_13714,N_12718);
nor U14317 (N_14317,N_13545,N_13885);
and U14318 (N_14318,N_13825,N_13197);
nand U14319 (N_14319,N_12676,N_13336);
nor U14320 (N_14320,N_13570,N_12434);
nor U14321 (N_14321,N_12252,N_13289);
and U14322 (N_14322,N_12514,N_13731);
nand U14323 (N_14323,N_12080,N_12350);
and U14324 (N_14324,N_13819,N_13100);
and U14325 (N_14325,N_13784,N_13726);
and U14326 (N_14326,N_13315,N_12599);
or U14327 (N_14327,N_12837,N_12528);
nor U14328 (N_14328,N_12555,N_12568);
nand U14329 (N_14329,N_12172,N_12610);
or U14330 (N_14330,N_12933,N_13654);
nor U14331 (N_14331,N_12484,N_13576);
nand U14332 (N_14332,N_13184,N_13541);
xor U14333 (N_14333,N_13108,N_13194);
xor U14334 (N_14334,N_12196,N_12762);
and U14335 (N_14335,N_13397,N_12711);
nor U14336 (N_14336,N_13122,N_12703);
nand U14337 (N_14337,N_12853,N_12719);
nor U14338 (N_14338,N_13323,N_13206);
xnor U14339 (N_14339,N_13818,N_12889);
and U14340 (N_14340,N_12104,N_12627);
nor U14341 (N_14341,N_13068,N_13113);
nand U14342 (N_14342,N_12922,N_13369);
xnor U14343 (N_14343,N_12435,N_12253);
nor U14344 (N_14344,N_13160,N_13371);
nor U14345 (N_14345,N_13907,N_12056);
nor U14346 (N_14346,N_12886,N_12764);
nand U14347 (N_14347,N_12552,N_13664);
and U14348 (N_14348,N_12657,N_13604);
xnor U14349 (N_14349,N_12460,N_13929);
nor U14350 (N_14350,N_13655,N_12341);
nor U14351 (N_14351,N_12202,N_12494);
and U14352 (N_14352,N_13580,N_13429);
nor U14353 (N_14353,N_12861,N_13953);
or U14354 (N_14354,N_12096,N_12689);
and U14355 (N_14355,N_12740,N_13822);
or U14356 (N_14356,N_12183,N_13480);
xnor U14357 (N_14357,N_13944,N_13215);
and U14358 (N_14358,N_12530,N_13733);
or U14359 (N_14359,N_12244,N_13381);
or U14360 (N_14360,N_12748,N_12028);
nand U14361 (N_14361,N_12522,N_12062);
nand U14362 (N_14362,N_13728,N_13383);
nor U14363 (N_14363,N_13066,N_12876);
or U14364 (N_14364,N_12071,N_13852);
or U14365 (N_14365,N_13407,N_13945);
and U14366 (N_14366,N_12114,N_13488);
or U14367 (N_14367,N_12219,N_12251);
nor U14368 (N_14368,N_13977,N_12108);
nand U14369 (N_14369,N_12602,N_12269);
nor U14370 (N_14370,N_12255,N_12963);
nand U14371 (N_14371,N_13801,N_12664);
nand U14372 (N_14372,N_12008,N_12982);
and U14373 (N_14373,N_12342,N_13103);
or U14374 (N_14374,N_12804,N_12684);
nor U14375 (N_14375,N_13071,N_12426);
nor U14376 (N_14376,N_12608,N_13504);
or U14377 (N_14377,N_13070,N_13552);
and U14378 (N_14378,N_12170,N_12921);
xnor U14379 (N_14379,N_12228,N_13278);
nor U14380 (N_14380,N_12968,N_12352);
nor U14381 (N_14381,N_13441,N_12920);
and U14382 (N_14382,N_12169,N_12498);
nand U14383 (N_14383,N_12967,N_12019);
or U14384 (N_14384,N_13893,N_12002);
nor U14385 (N_14385,N_13958,N_13463);
nor U14386 (N_14386,N_12020,N_13765);
nor U14387 (N_14387,N_13133,N_13772);
nor U14388 (N_14388,N_12109,N_13432);
xor U14389 (N_14389,N_12784,N_12749);
or U14390 (N_14390,N_12005,N_12961);
or U14391 (N_14391,N_12459,N_12155);
xor U14392 (N_14392,N_12525,N_12200);
and U14393 (N_14393,N_13217,N_13567);
or U14394 (N_14394,N_13270,N_13471);
nand U14395 (N_14395,N_13643,N_12979);
and U14396 (N_14396,N_12164,N_13970);
nor U14397 (N_14397,N_13889,N_13358);
nor U14398 (N_14398,N_13346,N_13073);
or U14399 (N_14399,N_12865,N_12223);
or U14400 (N_14400,N_12576,N_13749);
nand U14401 (N_14401,N_13141,N_12849);
nand U14402 (N_14402,N_13384,N_12429);
or U14403 (N_14403,N_13613,N_12216);
and U14404 (N_14404,N_12176,N_13201);
nand U14405 (N_14405,N_13416,N_13288);
nand U14406 (N_14406,N_13520,N_12779);
nand U14407 (N_14407,N_12124,N_12788);
or U14408 (N_14408,N_12296,N_12330);
or U14409 (N_14409,N_12596,N_12773);
nor U14410 (N_14410,N_13028,N_12229);
and U14411 (N_14411,N_12466,N_12268);
or U14412 (N_14412,N_13300,N_13343);
nor U14413 (N_14413,N_12828,N_12038);
and U14414 (N_14414,N_12533,N_12085);
or U14415 (N_14415,N_13779,N_12549);
or U14416 (N_14416,N_13337,N_13713);
and U14417 (N_14417,N_12810,N_12363);
xor U14418 (N_14418,N_12026,N_13564);
xnor U14419 (N_14419,N_13535,N_13896);
and U14420 (N_14420,N_13254,N_13540);
and U14421 (N_14421,N_12159,N_12224);
nand U14422 (N_14422,N_13808,N_12454);
nor U14423 (N_14423,N_13401,N_13200);
nor U14424 (N_14424,N_12541,N_12225);
xnor U14425 (N_14425,N_13835,N_13840);
xor U14426 (N_14426,N_13493,N_12938);
and U14427 (N_14427,N_13495,N_13123);
and U14428 (N_14428,N_12199,N_13339);
or U14429 (N_14429,N_12298,N_12780);
and U14430 (N_14430,N_13606,N_12057);
or U14431 (N_14431,N_13577,N_12092);
nand U14432 (N_14432,N_12720,N_12617);
nand U14433 (N_14433,N_12209,N_12462);
nor U14434 (N_14434,N_13053,N_13770);
and U14435 (N_14435,N_13166,N_12220);
or U14436 (N_14436,N_12156,N_13139);
nand U14437 (N_14437,N_12111,N_13880);
or U14438 (N_14438,N_13013,N_13098);
nor U14439 (N_14439,N_13973,N_13633);
or U14440 (N_14440,N_13544,N_12831);
nand U14441 (N_14441,N_13418,N_12148);
xor U14442 (N_14442,N_12113,N_13661);
nand U14443 (N_14443,N_12317,N_12864);
nor U14444 (N_14444,N_12450,N_13601);
or U14445 (N_14445,N_12859,N_13219);
nand U14446 (N_14446,N_12501,N_12359);
nor U14447 (N_14447,N_12173,N_12276);
and U14448 (N_14448,N_12395,N_12661);
or U14449 (N_14449,N_13833,N_13239);
and U14450 (N_14450,N_12189,N_13876);
and U14451 (N_14451,N_12524,N_13174);
nor U14452 (N_14452,N_12410,N_12150);
xnor U14453 (N_14453,N_13164,N_13039);
nor U14454 (N_14454,N_13954,N_12662);
and U14455 (N_14455,N_12616,N_13302);
nand U14456 (N_14456,N_13816,N_13140);
nand U14457 (N_14457,N_12585,N_12288);
and U14458 (N_14458,N_13794,N_13831);
nand U14459 (N_14459,N_13171,N_13996);
nor U14460 (N_14460,N_12083,N_13721);
and U14461 (N_14461,N_13790,N_13426);
nor U14462 (N_14462,N_12197,N_13858);
nand U14463 (N_14463,N_13777,N_12935);
nor U14464 (N_14464,N_13975,N_13280);
and U14465 (N_14465,N_12835,N_13635);
nand U14466 (N_14466,N_13528,N_13967);
nor U14467 (N_14467,N_13940,N_13933);
nand U14468 (N_14468,N_13396,N_12868);
nor U14469 (N_14469,N_12074,N_12230);
and U14470 (N_14470,N_13566,N_12365);
nor U14471 (N_14471,N_12275,N_13894);
or U14472 (N_14472,N_13360,N_13617);
nand U14473 (N_14473,N_12943,N_12327);
and U14474 (N_14474,N_13915,N_13237);
nand U14475 (N_14475,N_13883,N_12786);
nor U14476 (N_14476,N_13832,N_13437);
and U14477 (N_14477,N_12476,N_13699);
nand U14478 (N_14478,N_13845,N_13625);
and U14479 (N_14479,N_13252,N_13189);
nand U14480 (N_14480,N_12671,N_12333);
nand U14481 (N_14481,N_13011,N_13359);
xor U14482 (N_14482,N_12973,N_13783);
nor U14483 (N_14483,N_12456,N_12488);
nand U14484 (N_14484,N_12860,N_12419);
nand U14485 (N_14485,N_12039,N_12578);
or U14486 (N_14486,N_12644,N_12053);
or U14487 (N_14487,N_13408,N_12511);
and U14488 (N_14488,N_13345,N_13700);
and U14489 (N_14489,N_12273,N_12424);
nor U14490 (N_14490,N_13415,N_13628);
nor U14491 (N_14491,N_12682,N_12898);
or U14492 (N_14492,N_13256,N_13971);
xor U14493 (N_14493,N_12907,N_13231);
nor U14494 (N_14494,N_13789,N_13146);
nand U14495 (N_14495,N_12335,N_12213);
nand U14496 (N_14496,N_12751,N_12677);
nand U14497 (N_14497,N_13330,N_12670);
nor U14498 (N_14498,N_12210,N_12383);
and U14499 (N_14499,N_12066,N_13253);
nand U14500 (N_14500,N_12746,N_13117);
xnor U14501 (N_14501,N_13695,N_12846);
or U14502 (N_14502,N_12787,N_13390);
nor U14503 (N_14503,N_13079,N_12512);
and U14504 (N_14504,N_13313,N_12964);
nand U14505 (N_14505,N_13272,N_13694);
nor U14506 (N_14506,N_12119,N_13862);
xor U14507 (N_14507,N_13447,N_13102);
nand U14508 (N_14508,N_12099,N_13709);
xor U14509 (N_14509,N_13209,N_13754);
nand U14510 (N_14510,N_12370,N_12107);
or U14511 (N_14511,N_12041,N_13318);
nor U14512 (N_14512,N_13138,N_12502);
nor U14513 (N_14513,N_13673,N_13796);
nand U14514 (N_14514,N_12393,N_12713);
and U14515 (N_14515,N_13670,N_13530);
nand U14516 (N_14516,N_12312,N_13033);
and U14517 (N_14517,N_12023,N_12415);
or U14518 (N_14518,N_13837,N_13678);
nand U14519 (N_14519,N_13109,N_12239);
or U14520 (N_14520,N_13372,N_12351);
and U14521 (N_14521,N_13773,N_13723);
nand U14522 (N_14522,N_13060,N_13466);
and U14523 (N_14523,N_13419,N_13982);
nor U14524 (N_14524,N_12416,N_12974);
xnor U14525 (N_14525,N_13662,N_12154);
or U14526 (N_14526,N_13768,N_13681);
nand U14527 (N_14527,N_12009,N_12168);
or U14528 (N_14528,N_12436,N_13095);
nor U14529 (N_14529,N_13622,N_12945);
or U14530 (N_14530,N_12376,N_12369);
or U14531 (N_14531,N_12013,N_13586);
nand U14532 (N_14532,N_13483,N_13449);
and U14533 (N_14533,N_13484,N_12941);
and U14534 (N_14534,N_12971,N_13912);
and U14535 (N_14535,N_12022,N_13024);
nor U14536 (N_14536,N_13170,N_13392);
nor U14537 (N_14537,N_12112,N_12761);
or U14538 (N_14538,N_13331,N_12680);
and U14539 (N_14539,N_13748,N_12595);
and U14540 (N_14540,N_13497,N_12880);
nand U14541 (N_14541,N_12231,N_13881);
nor U14542 (N_14542,N_13172,N_12537);
or U14543 (N_14543,N_13051,N_13081);
or U14544 (N_14544,N_12639,N_12633);
or U14545 (N_14545,N_13067,N_12763);
nor U14546 (N_14546,N_12879,N_13188);
and U14547 (N_14547,N_13895,N_13605);
or U14548 (N_14548,N_13214,N_12044);
nor U14549 (N_14549,N_12163,N_13680);
nor U14550 (N_14550,N_13510,N_12531);
and U14551 (N_14551,N_13448,N_13226);
nor U14552 (N_14552,N_12733,N_12508);
nor U14553 (N_14553,N_12496,N_12073);
xor U14554 (N_14554,N_13966,N_13686);
and U14555 (N_14555,N_12479,N_12857);
or U14556 (N_14556,N_12307,N_13413);
nor U14557 (N_14557,N_12914,N_12615);
and U14558 (N_14558,N_13787,N_12443);
nand U14559 (N_14559,N_12523,N_12211);
nor U14560 (N_14560,N_12499,N_13803);
and U14561 (N_14561,N_12653,N_13763);
or U14562 (N_14562,N_12668,N_12033);
nand U14563 (N_14563,N_13568,N_13542);
or U14564 (N_14564,N_13676,N_12324);
nand U14565 (N_14565,N_13182,N_12406);
xor U14566 (N_14566,N_12414,N_13222);
xnor U14567 (N_14567,N_12338,N_13663);
nor U14568 (N_14568,N_13846,N_13433);
and U14569 (N_14569,N_12905,N_13482);
nor U14570 (N_14570,N_12031,N_12895);
nand U14571 (N_14571,N_13097,N_13521);
and U14572 (N_14572,N_12571,N_12404);
and U14573 (N_14573,N_12844,N_12329);
and U14574 (N_14574,N_13317,N_12387);
nor U14575 (N_14575,N_12332,N_13391);
or U14576 (N_14576,N_12546,N_13045);
nand U14577 (N_14577,N_13968,N_13979);
xor U14578 (N_14578,N_12120,N_12320);
nor U14579 (N_14579,N_13121,N_13091);
and U14580 (N_14580,N_12625,N_12581);
and U14581 (N_14581,N_12411,N_12423);
nor U14582 (N_14582,N_13356,N_13321);
and U14583 (N_14583,N_13513,N_13333);
nand U14584 (N_14584,N_12321,N_13514);
or U14585 (N_14585,N_12768,N_12257);
nand U14586 (N_14586,N_12620,N_13575);
and U14587 (N_14587,N_12193,N_12704);
and U14588 (N_14588,N_13811,N_12160);
nor U14589 (N_14589,N_12881,N_12248);
nor U14590 (N_14590,N_12727,N_13373);
nor U14591 (N_14591,N_12735,N_12980);
or U14592 (N_14592,N_13674,N_12142);
nand U14593 (N_14593,N_13434,N_12892);
nand U14594 (N_14594,N_12587,N_12966);
nor U14595 (N_14595,N_12305,N_12131);
nand U14596 (N_14596,N_12045,N_13467);
nor U14597 (N_14597,N_12470,N_13338);
nand U14598 (N_14598,N_13720,N_13802);
nor U14599 (N_14599,N_12656,N_13240);
and U14600 (N_14600,N_12328,N_13159);
xnor U14601 (N_14601,N_13047,N_12316);
or U14602 (N_14602,N_12437,N_12917);
nand U14603 (N_14603,N_13963,N_13927);
and U14604 (N_14604,N_12217,N_13518);
nand U14605 (N_14605,N_12493,N_13533);
xnor U14606 (N_14606,N_13065,N_12908);
and U14607 (N_14607,N_13919,N_13821);
or U14608 (N_14608,N_13296,N_13871);
or U14609 (N_14609,N_12490,N_12801);
or U14610 (N_14610,N_12486,N_13637);
nand U14611 (N_14611,N_12206,N_12812);
nand U14612 (N_14612,N_12070,N_13814);
or U14613 (N_14613,N_13018,N_12358);
nand U14614 (N_14614,N_13145,N_12453);
nor U14615 (N_14615,N_13344,N_12636);
nor U14616 (N_14616,N_13735,N_13211);
xor U14617 (N_14617,N_13287,N_13716);
nor U14618 (N_14618,N_12783,N_13127);
or U14619 (N_14619,N_12806,N_13191);
and U14620 (N_14620,N_12888,N_13340);
nand U14621 (N_14621,N_13827,N_13126);
or U14622 (N_14622,N_12915,N_12263);
or U14623 (N_14623,N_12527,N_13379);
and U14624 (N_14624,N_12675,N_12060);
and U14625 (N_14625,N_12345,N_12824);
or U14626 (N_14626,N_13001,N_12535);
and U14627 (N_14627,N_13325,N_12185);
or U14628 (N_14628,N_13157,N_13563);
and U14629 (N_14629,N_13704,N_13793);
nor U14630 (N_14630,N_12882,N_12282);
or U14631 (N_14631,N_13486,N_12278);
nand U14632 (N_14632,N_12166,N_12069);
or U14633 (N_14633,N_12049,N_12306);
nand U14634 (N_14634,N_12310,N_13326);
nand U14635 (N_14635,N_13867,N_12565);
or U14636 (N_14636,N_12469,N_13142);
or U14637 (N_14637,N_13120,N_13715);
nor U14638 (N_14638,N_12157,N_12403);
nand U14639 (N_14639,N_13430,N_13387);
and U14640 (N_14640,N_12584,N_13291);
or U14641 (N_14641,N_12364,N_13922);
nor U14642 (N_14642,N_13634,N_12006);
or U14643 (N_14643,N_12088,N_13795);
nor U14644 (N_14644,N_12681,N_12702);
nor U14645 (N_14645,N_13069,N_12651);
nand U14646 (N_14646,N_12992,N_13690);
and U14647 (N_14647,N_12272,N_13828);
and U14648 (N_14648,N_12728,N_13672);
nor U14649 (N_14649,N_12110,N_13569);
and U14650 (N_14650,N_12630,N_12927);
xor U14651 (N_14651,N_13329,N_12084);
or U14652 (N_14652,N_12998,N_12805);
nand U14653 (N_14653,N_12134,N_12570);
nor U14654 (N_14654,N_12356,N_13042);
or U14655 (N_14655,N_12158,N_12723);
nor U14656 (N_14656,N_12557,N_12842);
nor U14657 (N_14657,N_12724,N_13558);
and U14658 (N_14658,N_13048,N_12640);
nor U14659 (N_14659,N_13861,N_12082);
nor U14660 (N_14660,N_13834,N_13410);
and U14661 (N_14661,N_13857,N_12536);
nand U14662 (N_14662,N_13769,N_13597);
or U14663 (N_14663,N_13208,N_12181);
or U14664 (N_14664,N_12186,N_13017);
nor U14665 (N_14665,N_13981,N_13008);
nand U14666 (N_14666,N_13309,N_12816);
nand U14667 (N_14667,N_13649,N_12270);
or U14668 (N_14668,N_12238,N_12731);
and U14669 (N_14669,N_13089,N_13459);
nand U14670 (N_14670,N_13180,N_13583);
nand U14671 (N_14671,N_13736,N_13055);
or U14672 (N_14672,N_12693,N_13865);
or U14673 (N_14673,N_12843,N_12924);
nand U14674 (N_14674,N_12507,N_13707);
and U14675 (N_14675,N_12755,N_13978);
and U14676 (N_14676,N_12572,N_13135);
nor U14677 (N_14677,N_12067,N_12822);
or U14678 (N_14678,N_13299,N_12609);
and U14679 (N_14679,N_12318,N_13993);
or U14680 (N_14680,N_13412,N_12975);
or U14681 (N_14681,N_13435,N_13755);
nand U14682 (N_14682,N_12598,N_13136);
nor U14683 (N_14683,N_12442,N_13269);
and U14684 (N_14684,N_13076,N_13116);
nor U14685 (N_14685,N_13551,N_13263);
and U14686 (N_14686,N_13574,N_12621);
nand U14687 (N_14687,N_12162,N_12952);
nand U14688 (N_14688,N_13652,N_13196);
nand U14689 (N_14689,N_12838,N_13063);
xor U14690 (N_14690,N_12600,N_12153);
and U14691 (N_14691,N_13878,N_12700);
or U14692 (N_14692,N_13086,N_12794);
nor U14693 (N_14693,N_12378,N_13711);
and U14694 (N_14694,N_12929,N_12055);
and U14695 (N_14695,N_13320,N_12642);
nand U14696 (N_14696,N_13281,N_13557);
xor U14697 (N_14697,N_13404,N_12264);
or U14698 (N_14698,N_12261,N_12089);
or U14699 (N_14699,N_12697,N_13645);
nor U14700 (N_14700,N_12603,N_13327);
nand U14701 (N_14701,N_12355,N_13341);
nor U14702 (N_14702,N_13892,N_13805);
or U14703 (N_14703,N_13939,N_13032);
nand U14704 (N_14704,N_13144,N_12685);
or U14705 (N_14705,N_13537,N_12962);
nand U14706 (N_14706,N_13792,N_12872);
or U14707 (N_14707,N_12926,N_13490);
nor U14708 (N_14708,N_12516,N_13161);
nor U14709 (N_14709,N_12589,N_13860);
nor U14710 (N_14710,N_12372,N_12545);
nor U14711 (N_14711,N_12547,N_12757);
or U14712 (N_14712,N_12455,N_12340);
nor U14713 (N_14713,N_13611,N_12960);
or U14714 (N_14714,N_13478,N_13956);
or U14715 (N_14715,N_12885,N_13348);
or U14716 (N_14716,N_12405,N_13257);
and U14717 (N_14717,N_12643,N_13741);
nand U14718 (N_14718,N_13543,N_13587);
and U14719 (N_14719,N_13169,N_12467);
or U14720 (N_14720,N_12564,N_12129);
and U14721 (N_14721,N_12604,N_13361);
xor U14722 (N_14722,N_13403,N_12919);
or U14723 (N_14723,N_12893,N_13474);
or U14724 (N_14724,N_13995,N_12789);
or U14725 (N_14725,N_13591,N_12396);
or U14726 (N_14726,N_13534,N_13366);
and U14727 (N_14727,N_12607,N_12726);
nor U14728 (N_14728,N_13193,N_12075);
nor U14729 (N_14729,N_13388,N_13705);
or U14730 (N_14730,N_12944,N_13090);
or U14731 (N_14731,N_12910,N_12577);
and U14732 (N_14732,N_13515,N_13275);
nand U14733 (N_14733,N_13106,N_13608);
nor U14734 (N_14734,N_13949,N_13112);
or U14735 (N_14735,N_13732,N_12054);
nand U14736 (N_14736,N_12534,N_12821);
or U14737 (N_14737,N_12631,N_12894);
and U14738 (N_14738,N_12820,N_13347);
xor U14739 (N_14739,N_13529,N_13477);
or U14740 (N_14740,N_13847,N_13642);
and U14741 (N_14741,N_13698,N_12669);
and U14742 (N_14742,N_13717,N_12591);
or U14743 (N_14743,N_13398,N_12208);
nor U14744 (N_14744,N_12448,N_13666);
or U14745 (N_14745,N_12065,N_13335);
nand U14746 (N_14746,N_12781,N_12311);
nor U14747 (N_14747,N_12722,N_13099);
and U14748 (N_14748,N_13936,N_13475);
xor U14749 (N_14749,N_13301,N_13538);
or U14750 (N_14750,N_12999,N_12798);
xor U14751 (N_14751,N_12551,N_13224);
nand U14752 (N_14752,N_13517,N_12540);
and U14753 (N_14753,N_13004,N_12343);
and U14754 (N_14754,N_12347,N_12204);
nor U14755 (N_14755,N_13851,N_12745);
and U14756 (N_14756,N_12464,N_13872);
and U14757 (N_14757,N_12826,N_12691);
and U14758 (N_14758,N_13084,N_13701);
or U14759 (N_14759,N_12729,N_13798);
nor U14760 (N_14760,N_12145,N_12796);
xnor U14761 (N_14761,N_12357,N_13175);
or U14762 (N_14762,N_12916,N_12289);
nand U14763 (N_14763,N_13417,N_13969);
and U14764 (N_14764,N_13052,N_13151);
or U14765 (N_14765,N_13294,N_12725);
or U14766 (N_14766,N_12937,N_12368);
or U14767 (N_14767,N_12747,N_13710);
or U14768 (N_14768,N_13158,N_13395);
nand U14769 (N_14769,N_13657,N_13050);
or U14770 (N_14770,N_12447,N_13187);
nand U14771 (N_14771,N_13450,N_12431);
nor U14772 (N_14772,N_13925,N_12953);
nor U14773 (N_14773,N_12375,N_13508);
and U14774 (N_14774,N_12629,N_12198);
nand U14775 (N_14775,N_12247,N_13739);
or U14776 (N_14776,N_12736,N_12562);
nor U14777 (N_14777,N_13619,N_12017);
nor U14778 (N_14778,N_12567,N_12815);
nand U14779 (N_14779,N_13264,N_12243);
nand U14780 (N_14780,N_12854,N_12123);
and U14781 (N_14781,N_12760,N_12539);
nand U14782 (N_14782,N_13669,N_12122);
and U14783 (N_14783,N_12003,N_12457);
nor U14784 (N_14784,N_12297,N_13469);
and U14785 (N_14785,N_13616,N_12836);
xor U14786 (N_14786,N_13804,N_13992);
and U14787 (N_14787,N_13394,N_13114);
nand U14788 (N_14788,N_13044,N_13512);
or U14789 (N_14789,N_13797,N_12542);
nor U14790 (N_14790,N_12716,N_13990);
nor U14791 (N_14791,N_13920,N_12519);
nand U14792 (N_14792,N_12811,N_12417);
and U14793 (N_14793,N_13650,N_13603);
nand U14794 (N_14794,N_13607,N_12756);
or U14795 (N_14795,N_12532,N_12215);
nor U14796 (N_14796,N_12452,N_13245);
nor U14797 (N_14797,N_13692,N_12769);
and U14798 (N_14798,N_12759,N_13762);
and U14799 (N_14799,N_12174,N_13909);
or U14800 (N_14800,N_12852,N_13572);
nor U14801 (N_14801,N_12299,N_13986);
xnor U14802 (N_14802,N_13342,N_12472);
and U14803 (N_14803,N_13462,N_12839);
or U14804 (N_14804,N_13015,N_12556);
xnor U14805 (N_14805,N_13682,N_13439);
nor U14806 (N_14806,N_13427,N_12863);
nor U14807 (N_14807,N_12097,N_13058);
nor U14808 (N_14808,N_13411,N_13991);
and U14809 (N_14809,N_13357,N_13468);
nor U14810 (N_14810,N_13258,N_12371);
and U14811 (N_14811,N_13665,N_12634);
nand U14812 (N_14812,N_12813,N_12884);
and U14813 (N_14813,N_13767,N_12094);
nand U14814 (N_14814,N_13610,N_13476);
or U14815 (N_14815,N_12712,N_12386);
or U14816 (N_14816,N_12353,N_13250);
nor U14817 (N_14817,N_13629,N_13866);
nand U14818 (N_14818,N_12331,N_12509);
or U14819 (N_14819,N_12976,N_12972);
or U14820 (N_14820,N_13093,N_13352);
and U14821 (N_14821,N_13730,N_12785);
xnor U14822 (N_14822,N_13592,N_12121);
and U14823 (N_14823,N_12782,N_12458);
nand U14824 (N_14824,N_12582,N_13456);
or U14825 (N_14825,N_13423,N_13006);
nor U14826 (N_14826,N_12190,N_12187);
nand U14827 (N_14827,N_13884,N_13083);
or U14828 (N_14828,N_12136,N_12468);
and U14829 (N_14829,N_12188,N_13207);
nand U14830 (N_14830,N_13057,N_13813);
nand U14831 (N_14831,N_13841,N_13487);
and U14832 (N_14832,N_12601,N_12932);
and U14833 (N_14833,N_13938,N_12428);
nor U14834 (N_14834,N_12015,N_12883);
nand U14835 (N_14835,N_13273,N_12809);
and U14836 (N_14836,N_13882,N_12389);
nand U14837 (N_14837,N_13593,N_12678);
or U14838 (N_14838,N_12767,N_13204);
nor U14839 (N_14839,N_12518,N_13251);
xor U14840 (N_14840,N_12694,N_12698);
nor U14841 (N_14841,N_13719,N_12118);
and U14842 (N_14842,N_12841,N_13766);
or U14843 (N_14843,N_12674,N_12701);
nand U14844 (N_14844,N_13609,N_12750);
xnor U14845 (N_14845,N_13153,N_13247);
nand U14846 (N_14846,N_12422,N_12235);
or U14847 (N_14847,N_12946,N_13026);
and U14848 (N_14848,N_12313,N_13961);
or U14849 (N_14849,N_13177,N_13040);
nand U14850 (N_14850,N_13626,N_13703);
nand U14851 (N_14851,N_12249,N_12645);
and U14852 (N_14852,N_13916,N_13232);
or U14853 (N_14853,N_13491,N_12679);
xnor U14854 (N_14854,N_12997,N_13972);
nor U14855 (N_14855,N_13285,N_13905);
and U14856 (N_14856,N_12449,N_13526);
or U14857 (N_14857,N_13002,N_12232);
and U14858 (N_14858,N_12526,N_13455);
and U14859 (N_14859,N_13010,N_13101);
or U14860 (N_14860,N_12737,N_12823);
or U14861 (N_14861,N_12323,N_13162);
and U14862 (N_14862,N_12984,N_13118);
nor U14863 (N_14863,N_12014,N_12079);
nand U14864 (N_14864,N_13481,N_13124);
nand U14865 (N_14865,N_13599,N_12673);
and U14866 (N_14866,N_13261,N_12302);
or U14867 (N_14867,N_12510,N_13745);
nor U14868 (N_14868,N_12029,N_12753);
nor U14869 (N_14869,N_13041,N_13035);
or U14870 (N_14870,N_12385,N_13998);
and U14871 (N_14871,N_12696,N_13054);
or U14872 (N_14872,N_12791,N_12427);
xnor U14873 (N_14873,N_12626,N_12896);
and U14874 (N_14874,N_13446,N_13268);
nand U14875 (N_14875,N_12294,N_13887);
xnor U14876 (N_14876,N_12440,N_13130);
and U14877 (N_14877,N_13355,N_12774);
nor U14878 (N_14878,N_12990,N_12612);
nor U14879 (N_14879,N_13350,N_12833);
or U14880 (N_14880,N_12866,N_12475);
or U14881 (N_14881,N_12407,N_12931);
xnor U14882 (N_14882,N_12891,N_12878);
and U14883 (N_14883,N_13685,N_12592);
nand U14884 (N_14884,N_12993,N_13400);
nor U14885 (N_14885,N_12178,N_12942);
nor U14886 (N_14886,N_13621,N_12281);
nor U14887 (N_14887,N_13519,N_12421);
xor U14888 (N_14888,N_12184,N_12102);
and U14889 (N_14889,N_12290,N_12274);
nand U14890 (N_14890,N_13873,N_12240);
and U14891 (N_14891,N_13658,N_13708);
nor U14892 (N_14892,N_12295,N_13943);
or U14893 (N_14893,N_13594,N_12061);
or U14894 (N_14894,N_13778,N_13947);
and U14895 (N_14895,N_12995,N_12994);
nor U14896 (N_14896,N_12362,N_12899);
and U14897 (N_14897,N_13870,N_12613);
nor U14898 (N_14898,N_12978,N_13780);
nor U14899 (N_14899,N_13012,N_12873);
nor U14900 (N_14900,N_12799,N_13221);
xor U14901 (N_14901,N_13952,N_12090);
nand U14902 (N_14902,N_13729,N_13904);
nor U14903 (N_14903,N_12590,N_13332);
and U14904 (N_14904,N_12227,N_13029);
or U14905 (N_14905,N_13560,N_13367);
or U14906 (N_14906,N_12770,N_13573);
nand U14907 (N_14907,N_12394,N_12250);
nor U14908 (N_14908,N_12594,N_12105);
or U14909 (N_14909,N_13863,N_12040);
nor U14910 (N_14910,N_13351,N_12965);
or U14911 (N_14911,N_13362,N_12474);
or U14912 (N_14912,N_12554,N_13722);
nor U14913 (N_14913,N_13195,N_13725);
nor U14914 (N_14914,N_12771,N_13918);
nand U14915 (N_14915,N_13000,N_12212);
nor U14916 (N_14916,N_12683,N_12529);
nand U14917 (N_14917,N_12167,N_12043);
nor U14918 (N_14918,N_13683,N_13129);
nand U14919 (N_14919,N_12646,N_13744);
nor U14920 (N_14920,N_12016,N_13930);
nand U14921 (N_14921,N_12292,N_13428);
and U14922 (N_14922,N_13776,N_13660);
and U14923 (N_14923,N_12897,N_12432);
or U14924 (N_14924,N_12912,N_13761);
nand U14925 (N_14925,N_13906,N_12758);
nor U14926 (N_14926,N_12309,N_13241);
nor U14927 (N_14927,N_13959,N_13473);
and U14928 (N_14928,N_12660,N_12234);
and U14929 (N_14929,N_12658,N_12550);
or U14930 (N_14930,N_13319,N_12237);
nor U14931 (N_14931,N_12098,N_13128);
nand U14932 (N_14932,N_13314,N_12983);
nor U14933 (N_14933,N_12367,N_12566);
and U14934 (N_14934,N_13937,N_12304);
or U14935 (N_14935,N_13636,N_12011);
and U14936 (N_14936,N_13602,N_13119);
or U14937 (N_14937,N_13414,N_12236);
nor U14938 (N_14938,N_13539,N_13305);
or U14939 (N_14939,N_13647,N_12802);
and U14940 (N_14940,N_13688,N_13016);
nor U14941 (N_14941,N_12233,N_13505);
or U14942 (N_14942,N_13022,N_12923);
nand U14943 (N_14943,N_13751,N_13759);
nor U14944 (N_14944,N_13757,N_12928);
or U14945 (N_14945,N_13555,N_13830);
or U14946 (N_14946,N_13115,N_13451);
or U14947 (N_14947,N_12300,N_12399);
or U14948 (N_14948,N_12322,N_12742);
nor U14949 (N_14949,N_13420,N_13914);
or U14950 (N_14950,N_13205,N_12776);
nand U14951 (N_14951,N_13402,N_13304);
nand U14952 (N_14952,N_13007,N_13080);
xor U14953 (N_14953,N_12803,N_13393);
and U14954 (N_14954,N_12194,N_12077);
and U14955 (N_14955,N_13965,N_12412);
xor U14956 (N_14956,N_12918,N_13094);
or U14957 (N_14957,N_13855,N_12830);
or U14958 (N_14958,N_12465,N_12686);
and U14959 (N_14959,N_12010,N_12487);
and U14960 (N_14960,N_12956,N_13691);
nand U14961 (N_14961,N_12480,N_13897);
nand U14962 (N_14962,N_12100,N_12451);
or U14963 (N_14963,N_12266,N_12877);
nand U14964 (N_14964,N_13898,N_12433);
and U14965 (N_14965,N_13638,N_12076);
or U14966 (N_14966,N_13948,N_12503);
nor U14967 (N_14967,N_12845,N_13496);
and U14968 (N_14968,N_12583,N_12957);
or U14969 (N_14969,N_13105,N_13901);
or U14970 (N_14970,N_13879,N_13782);
nand U14971 (N_14971,N_13962,N_13443);
xor U14972 (N_14972,N_12218,N_13536);
and U14973 (N_14973,N_13198,N_13888);
xor U14974 (N_14974,N_12380,N_12137);
nor U14975 (N_14975,N_13743,N_13460);
or U14976 (N_14976,N_12373,N_13630);
nand U14977 (N_14977,N_12652,N_12579);
xnor U14978 (N_14978,N_12913,N_12954);
or U14979 (N_14979,N_13107,N_13444);
and U14980 (N_14980,N_12688,N_13173);
nand U14981 (N_14981,N_12064,N_13738);
and U14982 (N_14982,N_12624,N_13212);
nand U14983 (N_14983,N_13727,N_12388);
and U14984 (N_14984,N_13836,N_12628);
nand U14985 (N_14985,N_13923,N_12018);
nor U14986 (N_14986,N_12267,N_12851);
and U14987 (N_14987,N_12714,N_13286);
nor U14988 (N_14988,N_13185,N_12390);
or U14989 (N_14989,N_13436,N_12775);
or U14990 (N_14990,N_13989,N_12135);
nand U14991 (N_14991,N_12847,N_12478);
and U14992 (N_14992,N_13461,N_13368);
or U14993 (N_14993,N_13442,N_13590);
and U14994 (N_14994,N_12870,N_13458);
or U14995 (N_14995,N_13653,N_12091);
or U14996 (N_14996,N_12606,N_13651);
nor U14997 (N_14997,N_12985,N_12191);
nand U14998 (N_14998,N_12379,N_13489);
and U14999 (N_14999,N_13421,N_13485);
nand U15000 (N_15000,N_12891,N_12627);
or U15001 (N_15001,N_12808,N_13932);
or U15002 (N_15002,N_13929,N_13890);
or U15003 (N_15003,N_12383,N_13805);
or U15004 (N_15004,N_13769,N_13486);
nor U15005 (N_15005,N_13601,N_12804);
or U15006 (N_15006,N_13068,N_12318);
nand U15007 (N_15007,N_13699,N_12186);
xnor U15008 (N_15008,N_13951,N_12636);
and U15009 (N_15009,N_12341,N_13384);
nor U15010 (N_15010,N_12807,N_13168);
or U15011 (N_15011,N_12711,N_13158);
nand U15012 (N_15012,N_13581,N_13958);
or U15013 (N_15013,N_13599,N_12738);
nor U15014 (N_15014,N_13596,N_13849);
nand U15015 (N_15015,N_13028,N_12178);
or U15016 (N_15016,N_13487,N_12945);
nand U15017 (N_15017,N_12991,N_13750);
and U15018 (N_15018,N_12751,N_12896);
and U15019 (N_15019,N_13772,N_13007);
or U15020 (N_15020,N_13675,N_12184);
or U15021 (N_15021,N_13079,N_13536);
nand U15022 (N_15022,N_12723,N_12671);
and U15023 (N_15023,N_12956,N_13913);
and U15024 (N_15024,N_13950,N_12309);
nor U15025 (N_15025,N_13990,N_12307);
nor U15026 (N_15026,N_12783,N_12450);
xnor U15027 (N_15027,N_12450,N_12988);
or U15028 (N_15028,N_12216,N_12683);
and U15029 (N_15029,N_12025,N_12834);
nor U15030 (N_15030,N_13355,N_13817);
nor U15031 (N_15031,N_13341,N_12708);
nand U15032 (N_15032,N_13354,N_12323);
and U15033 (N_15033,N_12784,N_12657);
and U15034 (N_15034,N_13303,N_13306);
nand U15035 (N_15035,N_13292,N_13088);
or U15036 (N_15036,N_12680,N_12501);
and U15037 (N_15037,N_12004,N_13159);
nor U15038 (N_15038,N_12946,N_13967);
nand U15039 (N_15039,N_12049,N_12017);
nor U15040 (N_15040,N_13713,N_13382);
nand U15041 (N_15041,N_13327,N_13167);
nor U15042 (N_15042,N_12033,N_13212);
or U15043 (N_15043,N_12710,N_12028);
nand U15044 (N_15044,N_13994,N_12329);
or U15045 (N_15045,N_13122,N_13469);
nor U15046 (N_15046,N_12882,N_13917);
nor U15047 (N_15047,N_13006,N_13952);
or U15048 (N_15048,N_12338,N_12679);
nor U15049 (N_15049,N_13339,N_13702);
or U15050 (N_15050,N_13257,N_12403);
or U15051 (N_15051,N_12427,N_13921);
and U15052 (N_15052,N_12767,N_13864);
xor U15053 (N_15053,N_12786,N_12299);
xnor U15054 (N_15054,N_12535,N_13139);
and U15055 (N_15055,N_12704,N_12295);
and U15056 (N_15056,N_13482,N_12676);
nor U15057 (N_15057,N_12793,N_12251);
nor U15058 (N_15058,N_12859,N_12406);
or U15059 (N_15059,N_12124,N_12775);
and U15060 (N_15060,N_12148,N_13089);
and U15061 (N_15061,N_13530,N_12347);
nand U15062 (N_15062,N_12673,N_13753);
and U15063 (N_15063,N_12657,N_13797);
nand U15064 (N_15064,N_12346,N_12451);
xnor U15065 (N_15065,N_13868,N_13117);
or U15066 (N_15066,N_13303,N_13535);
nand U15067 (N_15067,N_12835,N_12954);
nor U15068 (N_15068,N_12593,N_13570);
or U15069 (N_15069,N_13932,N_12731);
nand U15070 (N_15070,N_12726,N_12634);
and U15071 (N_15071,N_12313,N_13484);
nor U15072 (N_15072,N_12851,N_12988);
nand U15073 (N_15073,N_12653,N_12777);
or U15074 (N_15074,N_13362,N_13190);
or U15075 (N_15075,N_13792,N_12129);
and U15076 (N_15076,N_12340,N_13445);
or U15077 (N_15077,N_13772,N_13102);
nor U15078 (N_15078,N_13713,N_12168);
and U15079 (N_15079,N_12077,N_13818);
nand U15080 (N_15080,N_12280,N_13590);
and U15081 (N_15081,N_12744,N_13882);
and U15082 (N_15082,N_13392,N_12467);
and U15083 (N_15083,N_12171,N_13242);
and U15084 (N_15084,N_13004,N_12180);
and U15085 (N_15085,N_12866,N_13070);
and U15086 (N_15086,N_13034,N_13216);
nand U15087 (N_15087,N_12015,N_12035);
nor U15088 (N_15088,N_12552,N_13507);
nand U15089 (N_15089,N_13638,N_12169);
nand U15090 (N_15090,N_13957,N_13828);
xnor U15091 (N_15091,N_12094,N_13977);
nor U15092 (N_15092,N_13418,N_13152);
xor U15093 (N_15093,N_12283,N_13391);
nand U15094 (N_15094,N_13479,N_13646);
nand U15095 (N_15095,N_13451,N_13953);
or U15096 (N_15096,N_12073,N_12269);
or U15097 (N_15097,N_13898,N_12479);
and U15098 (N_15098,N_13564,N_12454);
nand U15099 (N_15099,N_12023,N_12552);
and U15100 (N_15100,N_13820,N_12021);
nor U15101 (N_15101,N_13852,N_13176);
nor U15102 (N_15102,N_12702,N_12574);
or U15103 (N_15103,N_13334,N_12694);
or U15104 (N_15104,N_12710,N_13123);
nand U15105 (N_15105,N_12532,N_13056);
xor U15106 (N_15106,N_13269,N_13003);
nor U15107 (N_15107,N_13355,N_12087);
nor U15108 (N_15108,N_12953,N_12976);
nor U15109 (N_15109,N_13136,N_12482);
and U15110 (N_15110,N_12022,N_12816);
nor U15111 (N_15111,N_12480,N_12384);
or U15112 (N_15112,N_13916,N_13293);
nor U15113 (N_15113,N_12222,N_12593);
or U15114 (N_15114,N_13408,N_13587);
xnor U15115 (N_15115,N_13574,N_13714);
nor U15116 (N_15116,N_12044,N_13238);
and U15117 (N_15117,N_13289,N_12274);
and U15118 (N_15118,N_12189,N_12707);
nor U15119 (N_15119,N_12291,N_12664);
nor U15120 (N_15120,N_13802,N_13233);
nor U15121 (N_15121,N_13165,N_12878);
nand U15122 (N_15122,N_13390,N_13950);
and U15123 (N_15123,N_12680,N_12713);
or U15124 (N_15124,N_12470,N_12511);
nand U15125 (N_15125,N_12086,N_12630);
or U15126 (N_15126,N_12460,N_12492);
nand U15127 (N_15127,N_13380,N_12908);
and U15128 (N_15128,N_12091,N_12064);
and U15129 (N_15129,N_12080,N_13778);
or U15130 (N_15130,N_13932,N_12504);
or U15131 (N_15131,N_12011,N_13301);
or U15132 (N_15132,N_13145,N_13022);
and U15133 (N_15133,N_12576,N_12873);
nand U15134 (N_15134,N_12371,N_13489);
or U15135 (N_15135,N_13035,N_13899);
nor U15136 (N_15136,N_13978,N_12390);
or U15137 (N_15137,N_13799,N_13282);
nand U15138 (N_15138,N_13537,N_12060);
nor U15139 (N_15139,N_12234,N_13509);
xnor U15140 (N_15140,N_13709,N_13720);
nand U15141 (N_15141,N_12320,N_12408);
nor U15142 (N_15142,N_12396,N_13724);
nor U15143 (N_15143,N_13247,N_13213);
nor U15144 (N_15144,N_13910,N_13836);
nand U15145 (N_15145,N_12806,N_13735);
nor U15146 (N_15146,N_12333,N_12517);
or U15147 (N_15147,N_13476,N_12525);
nand U15148 (N_15148,N_13854,N_13783);
and U15149 (N_15149,N_12752,N_13723);
and U15150 (N_15150,N_12774,N_13151);
or U15151 (N_15151,N_12453,N_13184);
nor U15152 (N_15152,N_12992,N_13164);
nor U15153 (N_15153,N_13957,N_12952);
nor U15154 (N_15154,N_13865,N_12705);
nand U15155 (N_15155,N_13172,N_12848);
nand U15156 (N_15156,N_12403,N_12716);
and U15157 (N_15157,N_13573,N_13489);
or U15158 (N_15158,N_12020,N_12459);
nand U15159 (N_15159,N_12153,N_12735);
nand U15160 (N_15160,N_13261,N_13055);
nor U15161 (N_15161,N_12910,N_12572);
nor U15162 (N_15162,N_12102,N_13358);
nand U15163 (N_15163,N_13479,N_13655);
nand U15164 (N_15164,N_12949,N_12434);
and U15165 (N_15165,N_12344,N_12797);
and U15166 (N_15166,N_12859,N_13200);
nand U15167 (N_15167,N_13449,N_12539);
xor U15168 (N_15168,N_13980,N_12191);
nor U15169 (N_15169,N_12839,N_12835);
xor U15170 (N_15170,N_13290,N_13082);
or U15171 (N_15171,N_12617,N_12767);
nand U15172 (N_15172,N_12000,N_12084);
nor U15173 (N_15173,N_12676,N_13890);
or U15174 (N_15174,N_12870,N_12588);
nor U15175 (N_15175,N_12151,N_13397);
or U15176 (N_15176,N_13088,N_13602);
or U15177 (N_15177,N_12013,N_12130);
nand U15178 (N_15178,N_13699,N_13658);
and U15179 (N_15179,N_13715,N_12210);
or U15180 (N_15180,N_12105,N_13920);
nor U15181 (N_15181,N_12476,N_13319);
nor U15182 (N_15182,N_12298,N_12079);
and U15183 (N_15183,N_12431,N_13487);
and U15184 (N_15184,N_13713,N_13817);
or U15185 (N_15185,N_12543,N_12723);
and U15186 (N_15186,N_13649,N_12330);
nand U15187 (N_15187,N_13062,N_13012);
nand U15188 (N_15188,N_13553,N_13546);
nor U15189 (N_15189,N_13157,N_13371);
or U15190 (N_15190,N_13282,N_13908);
and U15191 (N_15191,N_12692,N_13468);
and U15192 (N_15192,N_13308,N_12163);
or U15193 (N_15193,N_12956,N_12297);
or U15194 (N_15194,N_13533,N_13464);
or U15195 (N_15195,N_12896,N_12776);
or U15196 (N_15196,N_12956,N_13167);
and U15197 (N_15197,N_12998,N_12166);
nor U15198 (N_15198,N_12841,N_12750);
nand U15199 (N_15199,N_13432,N_13197);
and U15200 (N_15200,N_12770,N_12060);
and U15201 (N_15201,N_13937,N_13482);
nor U15202 (N_15202,N_12873,N_12925);
nor U15203 (N_15203,N_13810,N_13745);
and U15204 (N_15204,N_12140,N_12139);
and U15205 (N_15205,N_12336,N_13662);
and U15206 (N_15206,N_12495,N_13458);
nand U15207 (N_15207,N_12717,N_13565);
nand U15208 (N_15208,N_13143,N_13280);
nand U15209 (N_15209,N_12285,N_13844);
nor U15210 (N_15210,N_13119,N_13340);
and U15211 (N_15211,N_12078,N_13442);
and U15212 (N_15212,N_12725,N_12576);
nor U15213 (N_15213,N_12719,N_12794);
and U15214 (N_15214,N_13411,N_13962);
xnor U15215 (N_15215,N_13878,N_12482);
nor U15216 (N_15216,N_12758,N_13255);
or U15217 (N_15217,N_12645,N_13548);
nor U15218 (N_15218,N_12688,N_12999);
nand U15219 (N_15219,N_13016,N_13894);
or U15220 (N_15220,N_12269,N_13615);
nor U15221 (N_15221,N_12176,N_13804);
and U15222 (N_15222,N_13640,N_12465);
xnor U15223 (N_15223,N_12471,N_13617);
nand U15224 (N_15224,N_13500,N_13656);
or U15225 (N_15225,N_13964,N_13105);
and U15226 (N_15226,N_12102,N_13346);
and U15227 (N_15227,N_13921,N_12031);
nor U15228 (N_15228,N_13968,N_12463);
or U15229 (N_15229,N_13748,N_13485);
nor U15230 (N_15230,N_13661,N_13046);
or U15231 (N_15231,N_13390,N_12928);
or U15232 (N_15232,N_12684,N_12360);
nand U15233 (N_15233,N_12109,N_13132);
xnor U15234 (N_15234,N_13086,N_13723);
or U15235 (N_15235,N_12008,N_12338);
nand U15236 (N_15236,N_13395,N_13324);
nand U15237 (N_15237,N_13939,N_13295);
or U15238 (N_15238,N_13794,N_13594);
and U15239 (N_15239,N_12685,N_12213);
or U15240 (N_15240,N_12922,N_12056);
nand U15241 (N_15241,N_12896,N_12184);
and U15242 (N_15242,N_12214,N_12314);
nor U15243 (N_15243,N_13072,N_13577);
nand U15244 (N_15244,N_13606,N_13776);
or U15245 (N_15245,N_13923,N_12251);
and U15246 (N_15246,N_12781,N_13305);
nor U15247 (N_15247,N_13588,N_13835);
nor U15248 (N_15248,N_12581,N_13232);
or U15249 (N_15249,N_12717,N_13626);
nand U15250 (N_15250,N_13986,N_13541);
and U15251 (N_15251,N_13692,N_12401);
nand U15252 (N_15252,N_12000,N_12204);
or U15253 (N_15253,N_13399,N_13554);
nand U15254 (N_15254,N_13107,N_13734);
nand U15255 (N_15255,N_12038,N_12806);
or U15256 (N_15256,N_12517,N_12140);
or U15257 (N_15257,N_13905,N_13030);
and U15258 (N_15258,N_13126,N_12661);
and U15259 (N_15259,N_12871,N_12894);
and U15260 (N_15260,N_12839,N_12197);
or U15261 (N_15261,N_13092,N_12233);
xnor U15262 (N_15262,N_12002,N_13351);
and U15263 (N_15263,N_12877,N_12596);
xnor U15264 (N_15264,N_13917,N_12401);
or U15265 (N_15265,N_13908,N_12029);
nand U15266 (N_15266,N_12987,N_13914);
and U15267 (N_15267,N_13546,N_12411);
nand U15268 (N_15268,N_13610,N_13560);
nor U15269 (N_15269,N_13366,N_13369);
xor U15270 (N_15270,N_13852,N_13168);
nand U15271 (N_15271,N_12709,N_13020);
nand U15272 (N_15272,N_13190,N_12410);
or U15273 (N_15273,N_12682,N_13612);
or U15274 (N_15274,N_12696,N_12207);
nor U15275 (N_15275,N_12077,N_12054);
and U15276 (N_15276,N_12617,N_13846);
nand U15277 (N_15277,N_13782,N_12717);
and U15278 (N_15278,N_13597,N_13893);
nor U15279 (N_15279,N_13580,N_12759);
nor U15280 (N_15280,N_12820,N_12459);
nand U15281 (N_15281,N_13261,N_12798);
nand U15282 (N_15282,N_13299,N_13975);
or U15283 (N_15283,N_13971,N_12039);
nor U15284 (N_15284,N_12566,N_13185);
nor U15285 (N_15285,N_13200,N_12483);
nor U15286 (N_15286,N_12323,N_12381);
and U15287 (N_15287,N_13827,N_12070);
nor U15288 (N_15288,N_12763,N_13771);
and U15289 (N_15289,N_13808,N_13228);
nand U15290 (N_15290,N_12671,N_13839);
nand U15291 (N_15291,N_13934,N_13421);
xnor U15292 (N_15292,N_12683,N_12767);
nor U15293 (N_15293,N_12834,N_12400);
nand U15294 (N_15294,N_13183,N_12639);
nor U15295 (N_15295,N_13995,N_12182);
and U15296 (N_15296,N_12464,N_12019);
xor U15297 (N_15297,N_13479,N_12694);
nor U15298 (N_15298,N_12996,N_12224);
or U15299 (N_15299,N_12583,N_13088);
and U15300 (N_15300,N_13349,N_12937);
and U15301 (N_15301,N_12345,N_13963);
nor U15302 (N_15302,N_13398,N_13322);
nor U15303 (N_15303,N_13532,N_13644);
nand U15304 (N_15304,N_13125,N_13869);
nand U15305 (N_15305,N_13870,N_13372);
nor U15306 (N_15306,N_13293,N_12240);
or U15307 (N_15307,N_13668,N_12984);
or U15308 (N_15308,N_13718,N_12117);
xnor U15309 (N_15309,N_13340,N_13221);
and U15310 (N_15310,N_12530,N_13329);
and U15311 (N_15311,N_12306,N_13542);
or U15312 (N_15312,N_13865,N_12954);
or U15313 (N_15313,N_13963,N_12344);
xnor U15314 (N_15314,N_12850,N_13393);
or U15315 (N_15315,N_13091,N_12339);
nor U15316 (N_15316,N_13679,N_12208);
or U15317 (N_15317,N_13969,N_12256);
xor U15318 (N_15318,N_13110,N_13895);
nand U15319 (N_15319,N_12213,N_12795);
and U15320 (N_15320,N_12659,N_13528);
nand U15321 (N_15321,N_13292,N_13716);
xnor U15322 (N_15322,N_13307,N_13821);
xnor U15323 (N_15323,N_12725,N_13991);
nand U15324 (N_15324,N_12087,N_12098);
and U15325 (N_15325,N_13953,N_13471);
xor U15326 (N_15326,N_13835,N_12447);
nand U15327 (N_15327,N_13757,N_13832);
and U15328 (N_15328,N_12673,N_12524);
xnor U15329 (N_15329,N_12173,N_12609);
and U15330 (N_15330,N_12257,N_12965);
or U15331 (N_15331,N_13790,N_12031);
nor U15332 (N_15332,N_13885,N_12073);
nor U15333 (N_15333,N_13114,N_12930);
or U15334 (N_15334,N_13701,N_13129);
nand U15335 (N_15335,N_12380,N_13654);
nor U15336 (N_15336,N_12189,N_12766);
nand U15337 (N_15337,N_12895,N_12654);
nand U15338 (N_15338,N_12206,N_13987);
and U15339 (N_15339,N_12778,N_12749);
xor U15340 (N_15340,N_13762,N_13563);
nor U15341 (N_15341,N_13829,N_12930);
or U15342 (N_15342,N_13289,N_13515);
nor U15343 (N_15343,N_13365,N_12928);
nand U15344 (N_15344,N_13652,N_13747);
xor U15345 (N_15345,N_13915,N_12997);
nor U15346 (N_15346,N_12408,N_12539);
and U15347 (N_15347,N_12775,N_13782);
or U15348 (N_15348,N_13228,N_12302);
nand U15349 (N_15349,N_12636,N_12818);
xor U15350 (N_15350,N_12517,N_13023);
nand U15351 (N_15351,N_12668,N_12286);
xnor U15352 (N_15352,N_12517,N_13896);
or U15353 (N_15353,N_12498,N_12470);
and U15354 (N_15354,N_12244,N_13942);
nor U15355 (N_15355,N_12368,N_13022);
or U15356 (N_15356,N_12890,N_12816);
xnor U15357 (N_15357,N_13336,N_13002);
nand U15358 (N_15358,N_12622,N_13039);
nor U15359 (N_15359,N_12644,N_12432);
nand U15360 (N_15360,N_13699,N_12937);
xor U15361 (N_15361,N_13280,N_12465);
and U15362 (N_15362,N_12313,N_12458);
nand U15363 (N_15363,N_12583,N_12488);
nand U15364 (N_15364,N_12540,N_12237);
nor U15365 (N_15365,N_13567,N_13513);
or U15366 (N_15366,N_12006,N_13105);
or U15367 (N_15367,N_13198,N_12614);
nor U15368 (N_15368,N_12973,N_12633);
or U15369 (N_15369,N_12005,N_13659);
nor U15370 (N_15370,N_13581,N_12543);
nor U15371 (N_15371,N_13361,N_12722);
nor U15372 (N_15372,N_12311,N_13848);
xor U15373 (N_15373,N_13133,N_13034);
xnor U15374 (N_15374,N_13548,N_13884);
nor U15375 (N_15375,N_13515,N_13670);
nand U15376 (N_15376,N_12551,N_13910);
or U15377 (N_15377,N_13409,N_13004);
nor U15378 (N_15378,N_12431,N_12369);
nor U15379 (N_15379,N_13421,N_13231);
nand U15380 (N_15380,N_12151,N_13800);
and U15381 (N_15381,N_12983,N_13712);
nor U15382 (N_15382,N_12673,N_12034);
and U15383 (N_15383,N_12140,N_12144);
and U15384 (N_15384,N_13563,N_12563);
and U15385 (N_15385,N_13592,N_13124);
or U15386 (N_15386,N_13122,N_13112);
and U15387 (N_15387,N_12334,N_13583);
and U15388 (N_15388,N_12959,N_12359);
nor U15389 (N_15389,N_13454,N_13513);
xor U15390 (N_15390,N_12059,N_12727);
or U15391 (N_15391,N_12901,N_12761);
nor U15392 (N_15392,N_12360,N_12608);
or U15393 (N_15393,N_12593,N_13099);
or U15394 (N_15394,N_13770,N_13183);
nand U15395 (N_15395,N_12722,N_13031);
xnor U15396 (N_15396,N_13987,N_12970);
and U15397 (N_15397,N_13250,N_12177);
nor U15398 (N_15398,N_12754,N_12093);
nor U15399 (N_15399,N_12792,N_13241);
nand U15400 (N_15400,N_13043,N_12008);
nand U15401 (N_15401,N_12428,N_12611);
or U15402 (N_15402,N_13814,N_13788);
nor U15403 (N_15403,N_12880,N_12846);
and U15404 (N_15404,N_13638,N_12241);
nand U15405 (N_15405,N_13254,N_13284);
xor U15406 (N_15406,N_13426,N_12447);
and U15407 (N_15407,N_13205,N_13898);
nand U15408 (N_15408,N_12082,N_12477);
or U15409 (N_15409,N_12203,N_13356);
xnor U15410 (N_15410,N_12581,N_13940);
or U15411 (N_15411,N_13633,N_12593);
and U15412 (N_15412,N_12443,N_12238);
nand U15413 (N_15413,N_12503,N_12157);
nor U15414 (N_15414,N_12436,N_12386);
and U15415 (N_15415,N_13419,N_13673);
or U15416 (N_15416,N_12683,N_12453);
or U15417 (N_15417,N_12796,N_12835);
nor U15418 (N_15418,N_13289,N_12064);
or U15419 (N_15419,N_13869,N_12026);
and U15420 (N_15420,N_13493,N_12325);
nor U15421 (N_15421,N_12126,N_13048);
or U15422 (N_15422,N_12159,N_12913);
nand U15423 (N_15423,N_13285,N_13012);
xnor U15424 (N_15424,N_13662,N_12131);
nand U15425 (N_15425,N_13063,N_13894);
and U15426 (N_15426,N_13475,N_13408);
nor U15427 (N_15427,N_13298,N_13777);
or U15428 (N_15428,N_13981,N_13530);
xnor U15429 (N_15429,N_12102,N_13624);
and U15430 (N_15430,N_12438,N_13495);
nor U15431 (N_15431,N_13958,N_13171);
nor U15432 (N_15432,N_12776,N_13281);
nor U15433 (N_15433,N_12818,N_12815);
nand U15434 (N_15434,N_13937,N_12788);
or U15435 (N_15435,N_12868,N_13125);
and U15436 (N_15436,N_12477,N_12590);
and U15437 (N_15437,N_13150,N_13127);
nand U15438 (N_15438,N_13664,N_12031);
nand U15439 (N_15439,N_13285,N_12011);
and U15440 (N_15440,N_12469,N_12019);
nor U15441 (N_15441,N_12257,N_13027);
xnor U15442 (N_15442,N_12188,N_12772);
nor U15443 (N_15443,N_13521,N_12599);
xor U15444 (N_15444,N_12491,N_13277);
nand U15445 (N_15445,N_12412,N_13859);
nor U15446 (N_15446,N_13085,N_12418);
nand U15447 (N_15447,N_12518,N_12848);
nor U15448 (N_15448,N_12764,N_13884);
and U15449 (N_15449,N_13683,N_12535);
or U15450 (N_15450,N_13174,N_12420);
or U15451 (N_15451,N_12351,N_12123);
or U15452 (N_15452,N_13536,N_12735);
or U15453 (N_15453,N_13573,N_13789);
or U15454 (N_15454,N_12654,N_13695);
and U15455 (N_15455,N_12263,N_12120);
xor U15456 (N_15456,N_13004,N_13329);
nand U15457 (N_15457,N_13872,N_12495);
and U15458 (N_15458,N_12106,N_12796);
and U15459 (N_15459,N_13745,N_12426);
and U15460 (N_15460,N_12999,N_12859);
nor U15461 (N_15461,N_13174,N_13285);
or U15462 (N_15462,N_13682,N_12647);
nor U15463 (N_15463,N_13146,N_13082);
or U15464 (N_15464,N_12866,N_12509);
xnor U15465 (N_15465,N_12902,N_13641);
nor U15466 (N_15466,N_12910,N_13897);
nor U15467 (N_15467,N_12994,N_12397);
and U15468 (N_15468,N_12509,N_13546);
xor U15469 (N_15469,N_12012,N_12946);
and U15470 (N_15470,N_13322,N_12982);
xnor U15471 (N_15471,N_13484,N_12664);
or U15472 (N_15472,N_13312,N_12223);
or U15473 (N_15473,N_12420,N_12597);
or U15474 (N_15474,N_12653,N_12778);
and U15475 (N_15475,N_13025,N_12396);
nand U15476 (N_15476,N_13642,N_12333);
nor U15477 (N_15477,N_12886,N_13294);
nand U15478 (N_15478,N_12693,N_13882);
nor U15479 (N_15479,N_13412,N_12191);
or U15480 (N_15480,N_12773,N_12188);
or U15481 (N_15481,N_12093,N_13749);
or U15482 (N_15482,N_12342,N_12677);
xnor U15483 (N_15483,N_13176,N_12881);
nor U15484 (N_15484,N_13490,N_13219);
or U15485 (N_15485,N_12941,N_13068);
nor U15486 (N_15486,N_12621,N_13816);
or U15487 (N_15487,N_13140,N_12422);
and U15488 (N_15488,N_12505,N_13223);
and U15489 (N_15489,N_12661,N_12499);
nor U15490 (N_15490,N_12868,N_12817);
xor U15491 (N_15491,N_13554,N_12340);
and U15492 (N_15492,N_12615,N_12650);
and U15493 (N_15493,N_13454,N_13875);
nor U15494 (N_15494,N_12924,N_13656);
and U15495 (N_15495,N_13736,N_12834);
and U15496 (N_15496,N_12336,N_12487);
and U15497 (N_15497,N_13408,N_12313);
or U15498 (N_15498,N_13780,N_13421);
or U15499 (N_15499,N_13734,N_12253);
or U15500 (N_15500,N_12529,N_12121);
nand U15501 (N_15501,N_13354,N_12617);
or U15502 (N_15502,N_13492,N_13227);
nor U15503 (N_15503,N_13565,N_13758);
nand U15504 (N_15504,N_12048,N_13465);
or U15505 (N_15505,N_12914,N_12531);
or U15506 (N_15506,N_13608,N_12713);
nand U15507 (N_15507,N_13215,N_13704);
or U15508 (N_15508,N_13654,N_13445);
nand U15509 (N_15509,N_13119,N_13140);
or U15510 (N_15510,N_12897,N_12878);
nor U15511 (N_15511,N_12685,N_13984);
or U15512 (N_15512,N_13846,N_13635);
nand U15513 (N_15513,N_12571,N_13375);
or U15514 (N_15514,N_13692,N_13677);
nand U15515 (N_15515,N_12962,N_12983);
and U15516 (N_15516,N_13479,N_12663);
xnor U15517 (N_15517,N_12104,N_12304);
nand U15518 (N_15518,N_13247,N_13776);
xor U15519 (N_15519,N_12604,N_13736);
and U15520 (N_15520,N_13810,N_12587);
or U15521 (N_15521,N_13395,N_13725);
xor U15522 (N_15522,N_12794,N_13342);
nand U15523 (N_15523,N_12104,N_12686);
xor U15524 (N_15524,N_13119,N_12669);
nor U15525 (N_15525,N_12265,N_12435);
and U15526 (N_15526,N_12738,N_12274);
and U15527 (N_15527,N_13391,N_13656);
nand U15528 (N_15528,N_13138,N_12173);
and U15529 (N_15529,N_12151,N_13096);
or U15530 (N_15530,N_13809,N_13572);
xor U15531 (N_15531,N_13011,N_12973);
or U15532 (N_15532,N_13442,N_12494);
nand U15533 (N_15533,N_12806,N_13296);
nor U15534 (N_15534,N_12362,N_13115);
nand U15535 (N_15535,N_13542,N_13633);
and U15536 (N_15536,N_12363,N_12859);
nor U15537 (N_15537,N_12821,N_13030);
nand U15538 (N_15538,N_12888,N_13771);
nand U15539 (N_15539,N_13545,N_12815);
nor U15540 (N_15540,N_12395,N_13047);
and U15541 (N_15541,N_13686,N_12210);
nor U15542 (N_15542,N_12440,N_12010);
nand U15543 (N_15543,N_13914,N_12780);
xor U15544 (N_15544,N_12406,N_13283);
or U15545 (N_15545,N_13433,N_12294);
nand U15546 (N_15546,N_13628,N_12073);
nand U15547 (N_15547,N_12138,N_12807);
or U15548 (N_15548,N_12567,N_12144);
xor U15549 (N_15549,N_12464,N_13287);
nor U15550 (N_15550,N_13819,N_12827);
and U15551 (N_15551,N_12348,N_12057);
nand U15552 (N_15552,N_12468,N_12263);
or U15553 (N_15553,N_12421,N_13156);
nor U15554 (N_15554,N_13428,N_12874);
nand U15555 (N_15555,N_12778,N_12493);
nor U15556 (N_15556,N_13087,N_12642);
and U15557 (N_15557,N_12986,N_12465);
and U15558 (N_15558,N_12184,N_12206);
nor U15559 (N_15559,N_13923,N_12618);
nor U15560 (N_15560,N_12015,N_12390);
nand U15561 (N_15561,N_12753,N_13879);
nand U15562 (N_15562,N_12246,N_13161);
xor U15563 (N_15563,N_12919,N_13411);
and U15564 (N_15564,N_13710,N_12295);
nor U15565 (N_15565,N_13028,N_13879);
nand U15566 (N_15566,N_12910,N_13534);
xnor U15567 (N_15567,N_13517,N_12679);
or U15568 (N_15568,N_13331,N_13479);
nand U15569 (N_15569,N_12884,N_12649);
and U15570 (N_15570,N_12024,N_13359);
nand U15571 (N_15571,N_12284,N_13739);
xnor U15572 (N_15572,N_12489,N_13768);
and U15573 (N_15573,N_13281,N_13667);
nor U15574 (N_15574,N_12499,N_13747);
and U15575 (N_15575,N_12290,N_12276);
and U15576 (N_15576,N_12090,N_13218);
xnor U15577 (N_15577,N_12561,N_12201);
or U15578 (N_15578,N_12863,N_12408);
nand U15579 (N_15579,N_13213,N_12125);
nand U15580 (N_15580,N_12388,N_12798);
or U15581 (N_15581,N_12236,N_12982);
or U15582 (N_15582,N_12426,N_12819);
nor U15583 (N_15583,N_13918,N_13853);
nand U15584 (N_15584,N_13225,N_12330);
or U15585 (N_15585,N_13606,N_12211);
nor U15586 (N_15586,N_13885,N_13443);
nor U15587 (N_15587,N_13614,N_12447);
or U15588 (N_15588,N_12462,N_13494);
or U15589 (N_15589,N_13037,N_13295);
xor U15590 (N_15590,N_12487,N_13564);
or U15591 (N_15591,N_13212,N_13617);
nand U15592 (N_15592,N_13564,N_12323);
and U15593 (N_15593,N_13526,N_13759);
nor U15594 (N_15594,N_12167,N_12284);
or U15595 (N_15595,N_12015,N_13852);
and U15596 (N_15596,N_12250,N_13986);
xnor U15597 (N_15597,N_12449,N_12764);
xor U15598 (N_15598,N_13727,N_12725);
and U15599 (N_15599,N_12384,N_12740);
or U15600 (N_15600,N_12316,N_13483);
nand U15601 (N_15601,N_13972,N_13208);
or U15602 (N_15602,N_13324,N_13616);
nand U15603 (N_15603,N_13055,N_13663);
or U15604 (N_15604,N_12495,N_13736);
xor U15605 (N_15605,N_12176,N_12570);
or U15606 (N_15606,N_12848,N_13269);
nand U15607 (N_15607,N_13905,N_12976);
nor U15608 (N_15608,N_12821,N_12718);
xnor U15609 (N_15609,N_12677,N_12979);
or U15610 (N_15610,N_12909,N_12215);
or U15611 (N_15611,N_12937,N_13832);
nor U15612 (N_15612,N_12809,N_13022);
or U15613 (N_15613,N_13593,N_12829);
nand U15614 (N_15614,N_12960,N_12639);
and U15615 (N_15615,N_13301,N_13738);
nand U15616 (N_15616,N_13375,N_12099);
nor U15617 (N_15617,N_12530,N_12939);
nor U15618 (N_15618,N_13975,N_12667);
xnor U15619 (N_15619,N_13435,N_12313);
nor U15620 (N_15620,N_13526,N_12380);
and U15621 (N_15621,N_12816,N_12959);
xnor U15622 (N_15622,N_13733,N_12306);
nand U15623 (N_15623,N_13140,N_13865);
xnor U15624 (N_15624,N_13984,N_13022);
nand U15625 (N_15625,N_12601,N_12326);
nand U15626 (N_15626,N_12786,N_13261);
or U15627 (N_15627,N_13877,N_13524);
nor U15628 (N_15628,N_12259,N_12268);
nor U15629 (N_15629,N_12597,N_13658);
and U15630 (N_15630,N_12275,N_13480);
and U15631 (N_15631,N_13123,N_12360);
or U15632 (N_15632,N_12975,N_13719);
or U15633 (N_15633,N_12660,N_13744);
nor U15634 (N_15634,N_12047,N_12884);
and U15635 (N_15635,N_13230,N_13226);
nor U15636 (N_15636,N_12917,N_12307);
nand U15637 (N_15637,N_13600,N_13382);
or U15638 (N_15638,N_13598,N_13544);
nand U15639 (N_15639,N_13508,N_12687);
and U15640 (N_15640,N_13154,N_12753);
nor U15641 (N_15641,N_12047,N_12873);
nor U15642 (N_15642,N_12646,N_12852);
or U15643 (N_15643,N_13531,N_13886);
xor U15644 (N_15644,N_13224,N_12557);
nand U15645 (N_15645,N_13880,N_13898);
xor U15646 (N_15646,N_12450,N_13477);
nor U15647 (N_15647,N_12647,N_13561);
nand U15648 (N_15648,N_13842,N_13792);
xnor U15649 (N_15649,N_13845,N_13682);
nor U15650 (N_15650,N_13170,N_12522);
xnor U15651 (N_15651,N_12671,N_13214);
nor U15652 (N_15652,N_13017,N_13414);
xor U15653 (N_15653,N_13521,N_13597);
and U15654 (N_15654,N_12238,N_12958);
and U15655 (N_15655,N_12462,N_13001);
nand U15656 (N_15656,N_13124,N_12178);
nor U15657 (N_15657,N_13702,N_13086);
nand U15658 (N_15658,N_13124,N_13423);
xor U15659 (N_15659,N_12510,N_13163);
xor U15660 (N_15660,N_12688,N_12117);
or U15661 (N_15661,N_13144,N_13320);
or U15662 (N_15662,N_12212,N_13408);
and U15663 (N_15663,N_13067,N_12018);
or U15664 (N_15664,N_13740,N_13939);
nor U15665 (N_15665,N_12157,N_12557);
and U15666 (N_15666,N_12721,N_13337);
nand U15667 (N_15667,N_13034,N_12526);
xnor U15668 (N_15668,N_13209,N_12602);
nor U15669 (N_15669,N_12839,N_12556);
or U15670 (N_15670,N_12359,N_13094);
xnor U15671 (N_15671,N_13994,N_13566);
nand U15672 (N_15672,N_13940,N_12219);
or U15673 (N_15673,N_12037,N_13640);
and U15674 (N_15674,N_13046,N_13613);
and U15675 (N_15675,N_13220,N_12786);
and U15676 (N_15676,N_12205,N_13710);
or U15677 (N_15677,N_13630,N_12361);
nand U15678 (N_15678,N_13251,N_12085);
and U15679 (N_15679,N_13716,N_13311);
or U15680 (N_15680,N_13434,N_12352);
nand U15681 (N_15681,N_13355,N_13113);
or U15682 (N_15682,N_12527,N_13110);
nand U15683 (N_15683,N_12988,N_12759);
and U15684 (N_15684,N_13362,N_12980);
and U15685 (N_15685,N_13534,N_12230);
nor U15686 (N_15686,N_13462,N_13789);
xnor U15687 (N_15687,N_13294,N_12906);
nand U15688 (N_15688,N_12261,N_13088);
nand U15689 (N_15689,N_13589,N_12216);
and U15690 (N_15690,N_13918,N_13931);
nor U15691 (N_15691,N_13654,N_13110);
nor U15692 (N_15692,N_12263,N_12773);
or U15693 (N_15693,N_13353,N_12136);
xnor U15694 (N_15694,N_13452,N_12310);
and U15695 (N_15695,N_13888,N_13668);
nor U15696 (N_15696,N_13541,N_13216);
or U15697 (N_15697,N_12063,N_12869);
nand U15698 (N_15698,N_13686,N_13301);
nor U15699 (N_15699,N_13061,N_13157);
or U15700 (N_15700,N_13076,N_12759);
nor U15701 (N_15701,N_12175,N_13721);
and U15702 (N_15702,N_13117,N_12265);
xor U15703 (N_15703,N_12877,N_12909);
nand U15704 (N_15704,N_12403,N_12314);
nand U15705 (N_15705,N_12508,N_12059);
or U15706 (N_15706,N_12369,N_12713);
and U15707 (N_15707,N_13534,N_13246);
nand U15708 (N_15708,N_13272,N_13542);
and U15709 (N_15709,N_12493,N_13377);
nor U15710 (N_15710,N_13971,N_13951);
nor U15711 (N_15711,N_13065,N_13395);
nor U15712 (N_15712,N_12727,N_12715);
and U15713 (N_15713,N_12841,N_12369);
nor U15714 (N_15714,N_12679,N_13332);
nand U15715 (N_15715,N_13648,N_12475);
or U15716 (N_15716,N_12366,N_13009);
nor U15717 (N_15717,N_12672,N_13474);
nand U15718 (N_15718,N_12790,N_13594);
nor U15719 (N_15719,N_13075,N_13675);
nor U15720 (N_15720,N_12799,N_12769);
nor U15721 (N_15721,N_13638,N_12330);
and U15722 (N_15722,N_13944,N_12248);
or U15723 (N_15723,N_12407,N_13999);
or U15724 (N_15724,N_12436,N_13880);
and U15725 (N_15725,N_12265,N_12692);
nor U15726 (N_15726,N_12329,N_13904);
or U15727 (N_15727,N_13987,N_12897);
and U15728 (N_15728,N_13933,N_12253);
and U15729 (N_15729,N_12500,N_13316);
and U15730 (N_15730,N_13097,N_12420);
and U15731 (N_15731,N_13527,N_13449);
nand U15732 (N_15732,N_13222,N_13883);
and U15733 (N_15733,N_13036,N_12547);
or U15734 (N_15734,N_13534,N_13552);
or U15735 (N_15735,N_13321,N_12628);
nor U15736 (N_15736,N_12761,N_13677);
nand U15737 (N_15737,N_12611,N_13234);
or U15738 (N_15738,N_12110,N_12734);
and U15739 (N_15739,N_12574,N_12975);
or U15740 (N_15740,N_13961,N_13483);
and U15741 (N_15741,N_13596,N_12478);
and U15742 (N_15742,N_12857,N_13171);
nand U15743 (N_15743,N_12105,N_12451);
nand U15744 (N_15744,N_12447,N_12778);
or U15745 (N_15745,N_12101,N_12553);
and U15746 (N_15746,N_12658,N_12309);
and U15747 (N_15747,N_13155,N_12480);
or U15748 (N_15748,N_13970,N_13421);
nand U15749 (N_15749,N_12599,N_12182);
or U15750 (N_15750,N_12585,N_13857);
and U15751 (N_15751,N_13927,N_13445);
nand U15752 (N_15752,N_13955,N_12120);
nor U15753 (N_15753,N_12148,N_12073);
or U15754 (N_15754,N_12467,N_13852);
nand U15755 (N_15755,N_13329,N_12999);
nor U15756 (N_15756,N_12649,N_12858);
and U15757 (N_15757,N_12954,N_12881);
and U15758 (N_15758,N_13972,N_13029);
nor U15759 (N_15759,N_12108,N_12660);
nor U15760 (N_15760,N_13127,N_13562);
or U15761 (N_15761,N_13930,N_13361);
or U15762 (N_15762,N_13451,N_13054);
and U15763 (N_15763,N_12615,N_12997);
or U15764 (N_15764,N_12324,N_13182);
nor U15765 (N_15765,N_13572,N_12075);
nor U15766 (N_15766,N_12257,N_12850);
xnor U15767 (N_15767,N_13246,N_12256);
nor U15768 (N_15768,N_12045,N_13093);
nand U15769 (N_15769,N_13727,N_13774);
xnor U15770 (N_15770,N_12601,N_12849);
or U15771 (N_15771,N_12397,N_12284);
and U15772 (N_15772,N_13980,N_13103);
xor U15773 (N_15773,N_12417,N_13118);
nand U15774 (N_15774,N_13346,N_12439);
or U15775 (N_15775,N_13220,N_13730);
nor U15776 (N_15776,N_13033,N_12869);
or U15777 (N_15777,N_13878,N_12620);
and U15778 (N_15778,N_13593,N_12374);
nand U15779 (N_15779,N_12205,N_13034);
and U15780 (N_15780,N_13094,N_12295);
or U15781 (N_15781,N_12838,N_13041);
nand U15782 (N_15782,N_13583,N_13204);
and U15783 (N_15783,N_12882,N_13540);
xor U15784 (N_15784,N_13555,N_13105);
or U15785 (N_15785,N_12084,N_12274);
or U15786 (N_15786,N_13361,N_13299);
nand U15787 (N_15787,N_13010,N_12386);
and U15788 (N_15788,N_12670,N_13750);
nor U15789 (N_15789,N_12125,N_13562);
or U15790 (N_15790,N_13559,N_13367);
nand U15791 (N_15791,N_12155,N_13501);
nand U15792 (N_15792,N_13144,N_12256);
or U15793 (N_15793,N_13418,N_12812);
nor U15794 (N_15794,N_12618,N_13556);
and U15795 (N_15795,N_13570,N_13080);
nand U15796 (N_15796,N_13884,N_13643);
or U15797 (N_15797,N_13961,N_12646);
nor U15798 (N_15798,N_12746,N_13290);
nand U15799 (N_15799,N_13593,N_12413);
or U15800 (N_15800,N_13161,N_12383);
or U15801 (N_15801,N_12243,N_12060);
and U15802 (N_15802,N_13732,N_13630);
nand U15803 (N_15803,N_13602,N_13531);
nor U15804 (N_15804,N_13503,N_13741);
or U15805 (N_15805,N_12144,N_12166);
and U15806 (N_15806,N_13136,N_13757);
nor U15807 (N_15807,N_12185,N_13762);
nand U15808 (N_15808,N_12049,N_13581);
or U15809 (N_15809,N_13840,N_13426);
nand U15810 (N_15810,N_13395,N_12416);
xor U15811 (N_15811,N_13027,N_12223);
and U15812 (N_15812,N_13491,N_13972);
or U15813 (N_15813,N_12188,N_12611);
or U15814 (N_15814,N_13370,N_13476);
and U15815 (N_15815,N_12107,N_13301);
nand U15816 (N_15816,N_12669,N_13906);
or U15817 (N_15817,N_13901,N_12165);
or U15818 (N_15818,N_12718,N_13665);
or U15819 (N_15819,N_12126,N_13059);
nand U15820 (N_15820,N_13864,N_12155);
or U15821 (N_15821,N_13590,N_13159);
nor U15822 (N_15822,N_13831,N_13897);
or U15823 (N_15823,N_13883,N_12187);
nand U15824 (N_15824,N_12788,N_13384);
or U15825 (N_15825,N_13522,N_13211);
and U15826 (N_15826,N_13806,N_13323);
nand U15827 (N_15827,N_12685,N_12543);
nor U15828 (N_15828,N_13508,N_13064);
or U15829 (N_15829,N_12394,N_13458);
or U15830 (N_15830,N_13823,N_13628);
or U15831 (N_15831,N_13640,N_13167);
nor U15832 (N_15832,N_12375,N_13082);
xor U15833 (N_15833,N_12752,N_13340);
nand U15834 (N_15834,N_12373,N_13289);
xnor U15835 (N_15835,N_12163,N_12753);
nand U15836 (N_15836,N_12273,N_13430);
or U15837 (N_15837,N_13602,N_12915);
nor U15838 (N_15838,N_13550,N_12368);
or U15839 (N_15839,N_13982,N_13402);
xor U15840 (N_15840,N_12984,N_12873);
or U15841 (N_15841,N_12574,N_12458);
or U15842 (N_15842,N_13533,N_12778);
or U15843 (N_15843,N_13107,N_12867);
nand U15844 (N_15844,N_12422,N_12980);
or U15845 (N_15845,N_12268,N_12736);
xor U15846 (N_15846,N_12424,N_13029);
and U15847 (N_15847,N_13454,N_13951);
and U15848 (N_15848,N_13060,N_13355);
and U15849 (N_15849,N_12245,N_12584);
nor U15850 (N_15850,N_12885,N_12781);
nor U15851 (N_15851,N_13458,N_13287);
and U15852 (N_15852,N_13770,N_12499);
or U15853 (N_15853,N_13326,N_13338);
xnor U15854 (N_15854,N_12055,N_13184);
or U15855 (N_15855,N_13747,N_12305);
nand U15856 (N_15856,N_13404,N_12683);
and U15857 (N_15857,N_12015,N_12792);
nor U15858 (N_15858,N_13520,N_12978);
nor U15859 (N_15859,N_12380,N_13847);
nor U15860 (N_15860,N_13930,N_12908);
nor U15861 (N_15861,N_13205,N_12039);
and U15862 (N_15862,N_12180,N_13709);
and U15863 (N_15863,N_13120,N_13425);
nand U15864 (N_15864,N_13029,N_13622);
or U15865 (N_15865,N_13439,N_12004);
nand U15866 (N_15866,N_12268,N_13922);
nand U15867 (N_15867,N_13688,N_13523);
xor U15868 (N_15868,N_13310,N_12373);
nand U15869 (N_15869,N_12485,N_13456);
nor U15870 (N_15870,N_13900,N_12387);
nand U15871 (N_15871,N_12896,N_13318);
nor U15872 (N_15872,N_13578,N_13086);
or U15873 (N_15873,N_13960,N_13981);
or U15874 (N_15874,N_13229,N_12883);
nand U15875 (N_15875,N_12414,N_13853);
xor U15876 (N_15876,N_13951,N_12781);
or U15877 (N_15877,N_13809,N_13337);
xnor U15878 (N_15878,N_12188,N_13155);
xnor U15879 (N_15879,N_12334,N_13082);
nor U15880 (N_15880,N_12648,N_12675);
and U15881 (N_15881,N_13287,N_13678);
nand U15882 (N_15882,N_12947,N_13510);
xor U15883 (N_15883,N_12764,N_12275);
and U15884 (N_15884,N_13813,N_13150);
xor U15885 (N_15885,N_13286,N_13105);
nand U15886 (N_15886,N_12640,N_13413);
or U15887 (N_15887,N_12480,N_12934);
xor U15888 (N_15888,N_13485,N_12961);
nand U15889 (N_15889,N_13074,N_12275);
nor U15890 (N_15890,N_13428,N_12379);
nor U15891 (N_15891,N_12449,N_13115);
xnor U15892 (N_15892,N_13893,N_13028);
xnor U15893 (N_15893,N_13200,N_12991);
nand U15894 (N_15894,N_13818,N_12698);
nand U15895 (N_15895,N_12602,N_13988);
nand U15896 (N_15896,N_13788,N_13602);
xor U15897 (N_15897,N_13533,N_12886);
and U15898 (N_15898,N_13703,N_12694);
nor U15899 (N_15899,N_12064,N_13529);
xor U15900 (N_15900,N_12098,N_12023);
or U15901 (N_15901,N_12960,N_13550);
and U15902 (N_15902,N_13216,N_12407);
and U15903 (N_15903,N_13413,N_13954);
nand U15904 (N_15904,N_13347,N_12684);
nor U15905 (N_15905,N_13497,N_12944);
and U15906 (N_15906,N_12716,N_12255);
nand U15907 (N_15907,N_12538,N_12629);
nor U15908 (N_15908,N_13641,N_13155);
nand U15909 (N_15909,N_13236,N_12555);
nand U15910 (N_15910,N_13744,N_13434);
nand U15911 (N_15911,N_13002,N_13464);
or U15912 (N_15912,N_12896,N_13158);
nand U15913 (N_15913,N_13457,N_13969);
and U15914 (N_15914,N_13534,N_12499);
or U15915 (N_15915,N_13639,N_13138);
or U15916 (N_15916,N_12102,N_12680);
and U15917 (N_15917,N_12130,N_12856);
and U15918 (N_15918,N_13964,N_12489);
and U15919 (N_15919,N_13224,N_12353);
nand U15920 (N_15920,N_12683,N_13198);
nand U15921 (N_15921,N_12984,N_13068);
nor U15922 (N_15922,N_13144,N_13266);
nand U15923 (N_15923,N_12563,N_13179);
or U15924 (N_15924,N_12631,N_13395);
nor U15925 (N_15925,N_12723,N_12891);
or U15926 (N_15926,N_13094,N_12379);
xor U15927 (N_15927,N_12313,N_12675);
or U15928 (N_15928,N_12112,N_13355);
xnor U15929 (N_15929,N_13032,N_12109);
or U15930 (N_15930,N_13215,N_13516);
nand U15931 (N_15931,N_12212,N_13973);
nand U15932 (N_15932,N_13005,N_13519);
and U15933 (N_15933,N_12756,N_13158);
nor U15934 (N_15934,N_12745,N_13505);
nand U15935 (N_15935,N_12593,N_12834);
or U15936 (N_15936,N_12346,N_13528);
and U15937 (N_15937,N_12408,N_13549);
xnor U15938 (N_15938,N_12194,N_13559);
xnor U15939 (N_15939,N_13053,N_13069);
and U15940 (N_15940,N_12275,N_13905);
nand U15941 (N_15941,N_13173,N_12019);
and U15942 (N_15942,N_12050,N_12358);
nand U15943 (N_15943,N_13270,N_13103);
and U15944 (N_15944,N_12881,N_12800);
and U15945 (N_15945,N_13665,N_12104);
or U15946 (N_15946,N_13949,N_12545);
or U15947 (N_15947,N_13879,N_13983);
and U15948 (N_15948,N_13689,N_12417);
xor U15949 (N_15949,N_12288,N_13093);
and U15950 (N_15950,N_13286,N_13929);
nor U15951 (N_15951,N_12047,N_13998);
nand U15952 (N_15952,N_13052,N_13406);
nor U15953 (N_15953,N_13243,N_12286);
and U15954 (N_15954,N_13909,N_13719);
xnor U15955 (N_15955,N_13472,N_12210);
or U15956 (N_15956,N_13300,N_12228);
nand U15957 (N_15957,N_13161,N_13542);
or U15958 (N_15958,N_12910,N_12017);
or U15959 (N_15959,N_12828,N_13661);
xor U15960 (N_15960,N_13691,N_13250);
nor U15961 (N_15961,N_13825,N_12081);
or U15962 (N_15962,N_12677,N_12411);
and U15963 (N_15963,N_12038,N_13060);
nand U15964 (N_15964,N_13308,N_12019);
nor U15965 (N_15965,N_13351,N_12558);
or U15966 (N_15966,N_12566,N_12926);
and U15967 (N_15967,N_13327,N_12833);
or U15968 (N_15968,N_13642,N_13536);
and U15969 (N_15969,N_12381,N_13290);
nand U15970 (N_15970,N_13086,N_12614);
and U15971 (N_15971,N_12009,N_12302);
and U15972 (N_15972,N_12404,N_13204);
and U15973 (N_15973,N_13801,N_12938);
nand U15974 (N_15974,N_12864,N_13877);
nand U15975 (N_15975,N_12708,N_12852);
or U15976 (N_15976,N_12633,N_12780);
or U15977 (N_15977,N_13555,N_13840);
nand U15978 (N_15978,N_12840,N_13056);
or U15979 (N_15979,N_13121,N_13015);
and U15980 (N_15980,N_13660,N_13808);
or U15981 (N_15981,N_13642,N_12854);
nand U15982 (N_15982,N_13400,N_12999);
or U15983 (N_15983,N_13715,N_13113);
nor U15984 (N_15984,N_13158,N_12565);
or U15985 (N_15985,N_13676,N_13293);
nand U15986 (N_15986,N_12081,N_12693);
or U15987 (N_15987,N_13095,N_12035);
nand U15988 (N_15988,N_12451,N_12545);
or U15989 (N_15989,N_12783,N_13805);
or U15990 (N_15990,N_12493,N_13805);
and U15991 (N_15991,N_13533,N_12984);
nand U15992 (N_15992,N_13405,N_12496);
xor U15993 (N_15993,N_13798,N_12806);
or U15994 (N_15994,N_12040,N_12263);
xnor U15995 (N_15995,N_12199,N_12873);
nor U15996 (N_15996,N_13986,N_13005);
nor U15997 (N_15997,N_12369,N_13783);
nor U15998 (N_15998,N_12740,N_13628);
or U15999 (N_15999,N_12026,N_13798);
nor U16000 (N_16000,N_14525,N_14519);
or U16001 (N_16001,N_15465,N_14791);
nor U16002 (N_16002,N_14285,N_14298);
or U16003 (N_16003,N_14774,N_15925);
or U16004 (N_16004,N_14685,N_15919);
nor U16005 (N_16005,N_15365,N_14984);
nor U16006 (N_16006,N_15179,N_15795);
nand U16007 (N_16007,N_14709,N_14428);
or U16008 (N_16008,N_15697,N_14863);
and U16009 (N_16009,N_14434,N_14312);
or U16010 (N_16010,N_15609,N_15630);
nor U16011 (N_16011,N_14197,N_14206);
and U16012 (N_16012,N_15954,N_15330);
or U16013 (N_16013,N_14419,N_14003);
and U16014 (N_16014,N_15092,N_14891);
or U16015 (N_16015,N_15978,N_15643);
nand U16016 (N_16016,N_14758,N_14126);
nand U16017 (N_16017,N_14114,N_15757);
nand U16018 (N_16018,N_14269,N_14476);
nor U16019 (N_16019,N_14388,N_15865);
nand U16020 (N_16020,N_14590,N_15773);
or U16021 (N_16021,N_15046,N_15903);
or U16022 (N_16022,N_14760,N_14091);
nor U16023 (N_16023,N_15811,N_14949);
nand U16024 (N_16024,N_15584,N_14461);
or U16025 (N_16025,N_14327,N_14673);
nand U16026 (N_16026,N_14310,N_15950);
nor U16027 (N_16027,N_15771,N_14786);
nand U16028 (N_16028,N_15891,N_15900);
or U16029 (N_16029,N_14264,N_15449);
nand U16030 (N_16030,N_14575,N_14082);
nor U16031 (N_16031,N_14391,N_14515);
or U16032 (N_16032,N_14379,N_15955);
and U16033 (N_16033,N_15794,N_15393);
and U16034 (N_16034,N_15830,N_15062);
and U16035 (N_16035,N_14740,N_15076);
nor U16036 (N_16036,N_14293,N_14372);
and U16037 (N_16037,N_15091,N_14314);
xor U16038 (N_16038,N_15959,N_15305);
nor U16039 (N_16039,N_15364,N_14968);
nand U16040 (N_16040,N_14290,N_14976);
nor U16041 (N_16041,N_15575,N_14313);
or U16042 (N_16042,N_14231,N_14061);
nor U16043 (N_16043,N_14973,N_15034);
xnor U16044 (N_16044,N_14803,N_14636);
nand U16045 (N_16045,N_14606,N_14223);
xor U16046 (N_16046,N_15392,N_15132);
or U16047 (N_16047,N_15505,N_14492);
and U16048 (N_16048,N_14352,N_15486);
nor U16049 (N_16049,N_15413,N_15787);
and U16050 (N_16050,N_14805,N_15473);
or U16051 (N_16051,N_15633,N_14701);
or U16052 (N_16052,N_15451,N_15147);
or U16053 (N_16053,N_14794,N_14437);
nand U16054 (N_16054,N_15809,N_15253);
nor U16055 (N_16055,N_15241,N_14455);
nor U16056 (N_16056,N_15359,N_14315);
nor U16057 (N_16057,N_14363,N_14203);
xor U16058 (N_16058,N_15075,N_15420);
nor U16059 (N_16059,N_15382,N_14488);
nor U16060 (N_16060,N_15112,N_14523);
nor U16061 (N_16061,N_15597,N_15129);
nand U16062 (N_16062,N_14975,N_15769);
nand U16063 (N_16063,N_15541,N_15661);
or U16064 (N_16064,N_14602,N_14044);
nor U16065 (N_16065,N_14864,N_15144);
nand U16066 (N_16066,N_14167,N_15206);
nor U16067 (N_16067,N_14565,N_14398);
or U16068 (N_16068,N_15628,N_14268);
or U16069 (N_16069,N_15426,N_15437);
and U16070 (N_16070,N_14212,N_14539);
nand U16071 (N_16071,N_15434,N_15414);
nor U16072 (N_16072,N_15855,N_14107);
nand U16073 (N_16073,N_15588,N_14109);
and U16074 (N_16074,N_14422,N_14882);
and U16075 (N_16075,N_14302,N_14651);
nor U16076 (N_16076,N_14104,N_14219);
and U16077 (N_16077,N_14746,N_15782);
and U16078 (N_16078,N_14354,N_14335);
nand U16079 (N_16079,N_15512,N_14035);
or U16080 (N_16080,N_14272,N_14262);
nor U16081 (N_16081,N_14271,N_14042);
or U16082 (N_16082,N_15470,N_14407);
and U16083 (N_16083,N_15174,N_15133);
or U16084 (N_16084,N_15587,N_15495);
or U16085 (N_16085,N_14823,N_14039);
nand U16086 (N_16086,N_15840,N_15694);
or U16087 (N_16087,N_15126,N_14904);
nand U16088 (N_16088,N_14304,N_15515);
or U16089 (N_16089,N_14678,N_15490);
and U16090 (N_16090,N_14639,N_15309);
nand U16091 (N_16091,N_15337,N_14119);
or U16092 (N_16092,N_15931,N_14291);
nor U16093 (N_16093,N_14917,N_14466);
or U16094 (N_16094,N_14650,N_15537);
or U16095 (N_16095,N_14001,N_15806);
nand U16096 (N_16096,N_15025,N_15064);
or U16097 (N_16097,N_15984,N_14587);
nand U16098 (N_16098,N_14225,N_15156);
or U16099 (N_16099,N_14654,N_14100);
and U16100 (N_16100,N_15883,N_14883);
and U16101 (N_16101,N_15405,N_14374);
nor U16102 (N_16102,N_15496,N_14604);
nor U16103 (N_16103,N_14273,N_15790);
nor U16104 (N_16104,N_15606,N_15032);
xor U16105 (N_16105,N_14266,N_14308);
and U16106 (N_16106,N_14911,N_14614);
and U16107 (N_16107,N_15378,N_14189);
nand U16108 (N_16108,N_14198,N_14284);
and U16109 (N_16109,N_14669,N_14161);
xor U16110 (N_16110,N_14748,N_14265);
nand U16111 (N_16111,N_15605,N_15745);
nor U16112 (N_16112,N_14887,N_14494);
xor U16113 (N_16113,N_15325,N_14759);
or U16114 (N_16114,N_14845,N_14021);
and U16115 (N_16115,N_15298,N_14593);
nand U16116 (N_16116,N_14369,N_14784);
nand U16117 (N_16117,N_15059,N_15729);
nand U16118 (N_16118,N_15121,N_15868);
nor U16119 (N_16119,N_14873,N_15700);
or U16120 (N_16120,N_15508,N_14665);
nor U16121 (N_16121,N_15219,N_15583);
or U16122 (N_16122,N_15637,N_15109);
nor U16123 (N_16123,N_15224,N_14950);
nor U16124 (N_16124,N_15912,N_15755);
nand U16125 (N_16125,N_15957,N_15388);
or U16126 (N_16126,N_15577,N_14453);
or U16127 (N_16127,N_15923,N_14815);
or U16128 (N_16128,N_15525,N_14139);
nor U16129 (N_16129,N_14421,N_14509);
nand U16130 (N_16130,N_15417,N_15114);
nand U16131 (N_16131,N_14910,N_14877);
nor U16132 (N_16132,N_14839,N_14698);
nor U16133 (N_16133,N_15598,N_14329);
and U16134 (N_16134,N_15935,N_15138);
or U16135 (N_16135,N_14844,N_14380);
nor U16136 (N_16136,N_15350,N_15613);
nand U16137 (N_16137,N_14981,N_15024);
nor U16138 (N_16138,N_15140,N_14277);
nand U16139 (N_16139,N_14624,N_15313);
and U16140 (N_16140,N_15137,N_15906);
nor U16141 (N_16141,N_15646,N_15674);
or U16142 (N_16142,N_15779,N_14827);
and U16143 (N_16143,N_14344,N_15012);
or U16144 (N_16144,N_15679,N_14516);
nand U16145 (N_16145,N_15115,N_15676);
or U16146 (N_16146,N_14690,N_14037);
nand U16147 (N_16147,N_14214,N_14501);
nand U16148 (N_16148,N_14713,N_14148);
nand U16149 (N_16149,N_14207,N_14829);
nand U16150 (N_16150,N_14720,N_14643);
xnor U16151 (N_16151,N_15274,N_15998);
and U16152 (N_16152,N_15848,N_14259);
or U16153 (N_16153,N_14584,N_14945);
xnor U16154 (N_16154,N_15705,N_14529);
nand U16155 (N_16155,N_14051,N_15345);
nand U16156 (N_16156,N_15460,N_15347);
or U16157 (N_16157,N_15220,N_14648);
xor U16158 (N_16158,N_14856,N_14835);
and U16159 (N_16159,N_14158,N_14837);
or U16160 (N_16160,N_15479,N_15462);
or U16161 (N_16161,N_15673,N_15463);
nand U16162 (N_16162,N_15439,N_14510);
nor U16163 (N_16163,N_15469,N_14169);
and U16164 (N_16164,N_15030,N_14806);
nor U16165 (N_16165,N_15159,N_15722);
and U16166 (N_16166,N_14804,N_14424);
or U16167 (N_16167,N_15400,N_14581);
and U16168 (N_16168,N_15847,N_15027);
nand U16169 (N_16169,N_15678,N_14482);
or U16170 (N_16170,N_15639,N_14394);
or U16171 (N_16171,N_15358,N_14280);
xnor U16172 (N_16172,N_14731,N_14495);
nor U16173 (N_16173,N_15956,N_14792);
or U16174 (N_16174,N_15975,N_15073);
or U16175 (N_16175,N_14449,N_14465);
and U16176 (N_16176,N_14807,N_15792);
or U16177 (N_16177,N_15620,N_14719);
nand U16178 (N_16178,N_14591,N_14386);
nor U16179 (N_16179,N_14777,N_14186);
or U16180 (N_16180,N_15546,N_14228);
xnor U16181 (N_16181,N_15250,N_14348);
nand U16182 (N_16182,N_15349,N_14742);
nor U16183 (N_16183,N_15742,N_15893);
nor U16184 (N_16184,N_15670,N_14103);
nand U16185 (N_16185,N_15681,N_15895);
nand U16186 (N_16186,N_14825,N_15461);
or U16187 (N_16187,N_15653,N_14957);
or U16188 (N_16188,N_14063,N_14121);
or U16189 (N_16189,N_14953,N_14297);
or U16190 (N_16190,N_15228,N_15016);
nand U16191 (N_16191,N_14582,N_15863);
xor U16192 (N_16192,N_14566,N_14649);
or U16193 (N_16193,N_14847,N_14326);
nand U16194 (N_16194,N_14729,N_15264);
and U16195 (N_16195,N_15827,N_14890);
nor U16196 (N_16196,N_15858,N_15177);
nand U16197 (N_16197,N_14595,N_14652);
nand U16198 (N_16198,N_15524,N_15611);
nand U16199 (N_16199,N_15019,N_15712);
or U16200 (N_16200,N_14099,N_14535);
nand U16201 (N_16201,N_14281,N_15727);
xor U16202 (N_16202,N_14420,N_15738);
or U16203 (N_16203,N_14937,N_15514);
nor U16204 (N_16204,N_14627,N_15821);
nor U16205 (N_16205,N_15938,N_15867);
nand U16206 (N_16206,N_15979,N_15006);
and U16207 (N_16207,N_15185,N_15176);
or U16208 (N_16208,N_15520,N_14337);
nand U16209 (N_16209,N_14641,N_15339);
nor U16210 (N_16210,N_15615,N_14242);
or U16211 (N_16211,N_14403,N_15162);
nor U16212 (N_16212,N_14903,N_15856);
or U16213 (N_16213,N_15737,N_14834);
nand U16214 (N_16214,N_14022,N_14520);
xor U16215 (N_16215,N_14571,N_15892);
nand U16216 (N_16216,N_15235,N_14232);
xnor U16217 (N_16217,N_14245,N_14353);
or U16218 (N_16218,N_14017,N_14014);
and U16219 (N_16219,N_14468,N_15355);
nor U16220 (N_16220,N_15041,N_14160);
xnor U16221 (N_16221,N_14876,N_15381);
nor U16222 (N_16222,N_14721,N_15318);
or U16223 (N_16223,N_14728,N_15194);
and U16224 (N_16224,N_14090,N_15455);
nor U16225 (N_16225,N_14514,N_14123);
xor U16226 (N_16226,N_14412,N_14828);
nand U16227 (N_16227,N_15949,N_14912);
nand U16228 (N_16228,N_15864,N_14447);
nor U16229 (N_16229,N_14763,N_14059);
nand U16230 (N_16230,N_14630,N_14768);
and U16231 (N_16231,N_15994,N_15932);
or U16232 (N_16232,N_14282,N_15277);
nor U16233 (N_16233,N_15839,N_15168);
nand U16234 (N_16234,N_15270,N_14870);
or U16235 (N_16235,N_15053,N_15433);
nand U16236 (N_16236,N_15367,N_14801);
xor U16237 (N_16237,N_14754,N_14441);
and U16238 (N_16238,N_15902,N_14795);
nand U16239 (N_16239,N_14283,N_15214);
or U16240 (N_16240,N_14301,N_15435);
or U16241 (N_16241,N_15578,N_15532);
nand U16242 (N_16242,N_15299,N_15846);
nor U16243 (N_16243,N_15280,N_14317);
nand U16244 (N_16244,N_15651,N_14410);
and U16245 (N_16245,N_15262,N_14397);
xnor U16246 (N_16246,N_15748,N_14577);
nand U16247 (N_16247,N_14350,N_15838);
or U16248 (N_16248,N_15982,N_14629);
or U16249 (N_16249,N_15011,N_14248);
and U16250 (N_16250,N_15842,N_15884);
or U16251 (N_16251,N_14880,N_15338);
or U16252 (N_16252,N_15936,N_14444);
nor U16253 (N_16253,N_15110,N_14857);
nor U16254 (N_16254,N_15832,N_14311);
nor U16255 (N_16255,N_14075,N_15389);
and U16256 (N_16256,N_14462,N_14176);
and U16257 (N_16257,N_14905,N_14128);
nor U16258 (N_16258,N_15669,N_15829);
and U16259 (N_16259,N_14249,N_14540);
nand U16260 (N_16260,N_15283,N_14377);
or U16261 (N_16261,N_15560,N_14963);
xor U16262 (N_16262,N_15047,N_14137);
nor U16263 (N_16263,N_15209,N_15725);
xnor U16264 (N_16264,N_14522,N_15079);
xor U16265 (N_16265,N_15622,N_15428);
xnor U16266 (N_16266,N_15887,N_14031);
nor U16267 (N_16267,N_14151,N_14722);
nor U16268 (N_16268,N_15852,N_15986);
and U16269 (N_16269,N_14508,N_14771);
nand U16270 (N_16270,N_14147,N_14555);
or U16271 (N_16271,N_14362,N_14276);
and U16272 (N_16272,N_14788,N_14846);
and U16273 (N_16273,N_15111,N_14443);
xor U16274 (N_16274,N_14251,N_14964);
xor U16275 (N_16275,N_14108,N_15728);
and U16276 (N_16276,N_15559,N_15551);
nand U16277 (N_16277,N_14469,N_15482);
and U16278 (N_16278,N_14755,N_14113);
or U16279 (N_16279,N_14024,N_14002);
nand U16280 (N_16280,N_15203,N_15487);
or U16281 (N_16281,N_14382,N_14097);
nor U16282 (N_16282,N_14977,N_15749);
and U16283 (N_16283,N_15962,N_15198);
and U16284 (N_16284,N_15552,N_15410);
and U16285 (N_16285,N_14322,N_14433);
nand U16286 (N_16286,N_14843,N_15644);
nor U16287 (N_16287,N_14320,N_14533);
nor U16288 (N_16288,N_15934,N_15005);
and U16289 (N_16289,N_15010,N_14413);
nand U16290 (N_16290,N_14637,N_15844);
and U16291 (N_16291,N_15056,N_14171);
and U16292 (N_16292,N_14078,N_15103);
nor U16293 (N_16293,N_14416,N_15610);
and U16294 (N_16294,N_15668,N_14400);
or U16295 (N_16295,N_14838,N_15545);
and U16296 (N_16296,N_15672,N_14941);
nor U16297 (N_16297,N_15627,N_14138);
or U16298 (N_16298,N_14146,N_15450);
or U16299 (N_16299,N_15961,N_14193);
and U16300 (N_16300,N_15859,N_14733);
or U16301 (N_16301,N_14765,N_14702);
nor U16302 (N_16302,N_14734,N_14725);
and U16303 (N_16303,N_15617,N_14745);
or U16304 (N_16304,N_14338,N_14454);
nand U16305 (N_16305,N_14048,N_15511);
and U16306 (N_16306,N_15974,N_14275);
or U16307 (N_16307,N_15314,N_15108);
or U16308 (N_16308,N_14478,N_15503);
nand U16309 (N_16309,N_15734,N_14756);
and U16310 (N_16310,N_15399,N_15322);
or U16311 (N_16311,N_15044,N_15295);
xnor U16312 (N_16312,N_14684,N_15993);
nor U16313 (N_16313,N_15150,N_15265);
nand U16314 (N_16314,N_15008,N_15783);
or U16315 (N_16315,N_15599,N_15256);
nor U16316 (N_16316,N_14347,N_15101);
nor U16317 (N_16317,N_14036,N_15402);
or U16318 (N_16318,N_14484,N_15762);
and U16319 (N_16319,N_15180,N_14157);
nor U16320 (N_16320,N_14967,N_15777);
nor U16321 (N_16321,N_15078,N_14694);
nand U16322 (N_16322,N_15823,N_14747);
nand U16323 (N_16323,N_15564,N_14946);
or U16324 (N_16324,N_14389,N_14503);
nand U16325 (N_16325,N_15098,N_15491);
nand U16326 (N_16326,N_15039,N_15683);
nor U16327 (N_16327,N_14767,N_14655);
nor U16328 (N_16328,N_15415,N_14802);
xnor U16329 (N_16329,N_15269,N_14600);
nand U16330 (N_16330,N_15862,N_15908);
and U16331 (N_16331,N_15703,N_14188);
or U16332 (N_16332,N_14782,N_15123);
and U16333 (N_16333,N_15094,N_15650);
nor U16334 (N_16334,N_15544,N_15145);
xor U16335 (N_16335,N_15087,N_15621);
nor U16336 (N_16336,N_14739,N_14371);
or U16337 (N_16337,N_14030,N_15286);
or U16338 (N_16338,N_15197,N_15326);
and U16339 (N_16339,N_14130,N_14339);
nand U16340 (N_16340,N_15464,N_15813);
nor U16341 (N_16341,N_14050,N_15040);
or U16342 (N_16342,N_15441,N_14136);
nor U16343 (N_16343,N_15243,N_14247);
and U16344 (N_16344,N_15352,N_15539);
or U16345 (N_16345,N_15261,N_15763);
or U16346 (N_16346,N_14589,N_14274);
and U16347 (N_16347,N_14717,N_14598);
xnor U16348 (N_16348,N_14451,N_14106);
xor U16349 (N_16349,N_15589,N_14491);
nand U16350 (N_16350,N_15648,N_14653);
or U16351 (N_16351,N_15636,N_14092);
nand U16352 (N_16352,N_14253,N_14922);
nand U16353 (N_16353,N_15721,N_15665);
and U16354 (N_16354,N_14987,N_15788);
nor U16355 (N_16355,N_15408,N_14303);
or U16356 (N_16356,N_15289,N_15558);
and U16357 (N_16357,N_14543,N_14230);
xnor U16358 (N_16358,N_15770,N_14355);
nand U16359 (N_16359,N_14766,N_14808);
nand U16360 (N_16360,N_14735,N_14028);
and U16361 (N_16361,N_14683,N_14578);
nor U16362 (N_16362,N_14162,N_14526);
xnor U16363 (N_16363,N_14871,N_15474);
xor U16364 (N_16364,N_14789,N_15193);
and U16365 (N_16365,N_15234,N_15869);
or U16366 (N_16366,N_15785,N_15212);
and U16367 (N_16367,N_14635,N_15945);
or U16368 (N_16368,N_15088,N_15102);
or U16369 (N_16369,N_14738,N_14278);
nand U16370 (N_16370,N_15328,N_15805);
or U16371 (N_16371,N_15675,N_14330);
nor U16372 (N_16372,N_15845,N_15944);
and U16373 (N_16373,N_15375,N_14496);
and U16374 (N_16374,N_14961,N_14243);
or U16375 (N_16375,N_15063,N_15376);
nor U16376 (N_16376,N_15018,N_15985);
nor U16377 (N_16377,N_15816,N_15001);
nor U16378 (N_16378,N_15036,N_14418);
nor U16379 (N_16379,N_14594,N_15761);
and U16380 (N_16380,N_14633,N_15374);
nor U16381 (N_16381,N_15756,N_15686);
nor U16382 (N_16382,N_15124,N_14580);
xor U16383 (N_16383,N_15894,N_14296);
and U16384 (N_16384,N_14027,N_15475);
nor U16385 (N_16385,N_14551,N_14170);
xnor U16386 (N_16386,N_14087,N_15638);
and U16387 (N_16387,N_14813,N_15361);
and U16388 (N_16388,N_14568,N_14375);
and U16389 (N_16389,N_15710,N_15764);
or U16390 (N_16390,N_15017,N_15576);
or U16391 (N_16391,N_14885,N_15684);
and U16392 (N_16392,N_14955,N_14192);
nor U16393 (N_16393,N_15566,N_14164);
or U16394 (N_16394,N_15336,N_15320);
nand U16395 (N_16395,N_14153,N_15819);
or U16396 (N_16396,N_15850,N_14920);
nand U16397 (N_16397,N_15310,N_14707);
nor U16398 (N_16398,N_15281,N_14548);
and U16399 (N_16399,N_15983,N_15999);
nor U16400 (N_16400,N_14246,N_14178);
nor U16401 (N_16401,N_15579,N_14145);
nand U16402 (N_16402,N_15929,N_15752);
and U16403 (N_16403,N_15548,N_15372);
and U16404 (N_16404,N_15107,N_14133);
xor U16405 (N_16405,N_15574,N_15074);
and U16406 (N_16406,N_15726,N_15951);
and U16407 (N_16407,N_14493,N_14120);
and U16408 (N_16408,N_14438,N_15724);
or U16409 (N_16409,N_14716,N_14902);
or U16410 (N_16410,N_15000,N_15942);
or U16411 (N_16411,N_15937,N_14626);
nor U16412 (N_16412,N_14261,N_14215);
nand U16413 (N_16413,N_15458,N_14617);
or U16414 (N_16414,N_15227,N_15632);
xor U16415 (N_16415,N_14088,N_14235);
nor U16416 (N_16416,N_15704,N_15204);
nand U16417 (N_16417,N_14205,N_14840);
or U16418 (N_16418,N_15086,N_15713);
nand U16419 (N_16419,N_15746,N_14750);
or U16420 (N_16420,N_14965,N_15516);
nand U16421 (N_16421,N_15290,N_14122);
or U16422 (N_16422,N_14899,N_14393);
nor U16423 (N_16423,N_15872,N_14209);
nor U16424 (N_16424,N_15125,N_14116);
nor U16425 (N_16425,N_14677,N_15416);
or U16426 (N_16426,N_14986,N_15618);
nor U16427 (N_16427,N_14611,N_15128);
and U16428 (N_16428,N_15561,N_14854);
nand U16429 (N_16429,N_15278,N_14471);
and U16430 (N_16430,N_14569,N_15153);
or U16431 (N_16431,N_14111,N_15254);
nor U16432 (N_16432,N_15766,N_14681);
nor U16433 (N_16433,N_15205,N_15424);
and U16434 (N_16434,N_15456,N_14559);
nand U16435 (N_16435,N_15438,N_15952);
nor U16436 (N_16436,N_15554,N_15861);
and U16437 (N_16437,N_14150,N_15067);
nor U16438 (N_16438,N_15500,N_14980);
nor U16439 (N_16439,N_14570,N_15498);
or U16440 (N_16440,N_14066,N_15387);
nor U16441 (N_16441,N_14159,N_14019);
xnor U16442 (N_16442,N_15489,N_15750);
and U16443 (N_16443,N_15051,N_14190);
or U16444 (N_16444,N_14409,N_15760);
nand U16445 (N_16445,N_15948,N_15828);
nor U16446 (N_16446,N_15077,N_14221);
nand U16447 (N_16447,N_14213,N_15165);
nor U16448 (N_16448,N_15476,N_14898);
nor U16449 (N_16449,N_15781,N_14865);
or U16450 (N_16450,N_14043,N_15292);
nor U16451 (N_16451,N_15175,N_15022);
nor U16452 (N_16452,N_15042,N_15876);
and U16453 (N_16453,N_14435,N_15089);
or U16454 (N_16454,N_14279,N_15021);
or U16455 (N_16455,N_14489,N_15664);
nor U16456 (N_16456,N_15789,N_14200);
and U16457 (N_16457,N_15407,N_14737);
or U16458 (N_16458,N_15901,N_14609);
nand U16459 (N_16459,N_15989,N_14874);
and U16460 (N_16460,N_14426,N_15642);
nor U16461 (N_16461,N_14105,N_14757);
nor U16462 (N_16462,N_14006,N_15068);
nor U16463 (N_16463,N_15173,N_15351);
nand U16464 (N_16464,N_15333,N_14647);
nor U16465 (N_16465,N_14459,N_14692);
and U16466 (N_16466,N_14552,N_14554);
or U16467 (N_16467,N_15874,N_15249);
nor U16468 (N_16468,N_14381,N_14185);
nand U16469 (N_16469,N_15709,N_14060);
nor U16470 (N_16470,N_14993,N_15425);
xor U16471 (N_16471,N_14990,N_15826);
and U16472 (N_16472,N_15033,N_15189);
and U16473 (N_16473,N_15659,N_14054);
xor U16474 (N_16474,N_15431,N_14612);
nand U16475 (N_16475,N_15368,N_15273);
and U16476 (N_16476,N_14892,N_15690);
nor U16477 (N_16477,N_15301,N_14816);
and U16478 (N_16478,N_14970,N_14487);
nand U16479 (N_16479,N_15526,N_15453);
nor U16480 (N_16480,N_15802,N_14373);
xnor U16481 (N_16481,N_14546,N_15521);
xnor U16482 (N_16482,N_15196,N_14255);
and U16483 (N_16483,N_15055,N_15607);
or U16484 (N_16484,N_14849,N_14076);
nand U16485 (N_16485,N_15191,N_15649);
or U16486 (N_16486,N_15166,N_15481);
xnor U16487 (N_16487,N_15065,N_14370);
nand U16488 (N_16488,N_14007,N_15799);
nor U16489 (N_16489,N_15857,N_15446);
or U16490 (N_16490,N_14172,N_15641);
or U16491 (N_16491,N_15880,N_14041);
nor U16492 (N_16492,N_14718,N_15246);
nor U16493 (N_16493,N_15323,N_15720);
and U16494 (N_16494,N_15677,N_14842);
nand U16495 (N_16495,N_15404,N_15953);
nand U16496 (N_16496,N_15711,N_14972);
nor U16497 (N_16497,N_14557,N_14244);
nor U16498 (N_16498,N_15139,N_15626);
nand U16499 (N_16499,N_14483,N_14708);
nand U16500 (N_16500,N_15398,N_14693);
and U16501 (N_16501,N_14321,N_14399);
nand U16502 (N_16502,N_15570,N_14787);
and U16503 (N_16503,N_15383,N_15656);
nor U16504 (N_16504,N_14878,N_14086);
or U16505 (N_16505,N_15097,N_14697);
or U16506 (N_16506,N_14081,N_14342);
and U16507 (N_16507,N_15164,N_15366);
nand U16508 (N_16508,N_14714,N_15430);
or U16509 (N_16509,N_14799,N_15775);
and U16510 (N_16510,N_15815,N_15595);
nand U16511 (N_16511,N_15625,N_14962);
xnor U16512 (N_16512,N_15841,N_15997);
nor U16513 (N_16513,N_15335,N_14679);
nor U16514 (N_16514,N_14621,N_14236);
nand U16515 (N_16515,N_15152,N_14779);
nand U16516 (N_16516,N_15810,N_14895);
nand U16517 (N_16517,N_15634,N_15751);
or U16518 (N_16518,N_15488,N_15553);
nor U16519 (N_16519,N_15267,N_14016);
nor U16520 (N_16520,N_15232,N_15692);
and U16521 (N_16521,N_15995,N_15853);
or U16522 (N_16522,N_15804,N_14065);
nand U16523 (N_16523,N_14009,N_15909);
nand U16524 (N_16524,N_15377,N_14727);
or U16525 (N_16525,N_14642,N_15406);
and U16526 (N_16526,N_15612,N_15066);
nand U16527 (N_16527,N_15971,N_15167);
nor U16528 (N_16528,N_15028,N_14850);
xor U16529 (N_16529,N_14936,N_14112);
or U16530 (N_16530,N_15026,N_15327);
nor U16531 (N_16531,N_14810,N_15218);
nand U16532 (N_16532,N_14919,N_14346);
xnor U16533 (N_16533,N_15940,N_14458);
and U16534 (N_16534,N_14928,N_14095);
or U16535 (N_16535,N_15141,N_14931);
or U16536 (N_16536,N_14442,N_15049);
nor U16537 (N_16537,N_15183,N_15118);
nor U16538 (N_16538,N_14680,N_15237);
nor U16539 (N_16539,N_14603,N_14723);
xor U16540 (N_16540,N_15741,N_14025);
or U16541 (N_16541,N_14183,N_14517);
nand U16542 (N_16542,N_14913,N_15100);
nand U16543 (N_16543,N_14676,N_15136);
nor U16544 (N_16544,N_15084,N_14940);
nor U16545 (N_16545,N_14574,N_15342);
xnor U16546 (N_16546,N_14662,N_15562);
and U16547 (N_16547,N_14744,N_14456);
and U16548 (N_16548,N_14541,N_15403);
and U16549 (N_16549,N_15427,N_14477);
and U16550 (N_16550,N_15468,N_14040);
and U16551 (N_16551,N_14942,N_14997);
nand U16552 (N_16552,N_15767,N_14199);
nand U16553 (N_16553,N_15740,N_14411);
nor U16554 (N_16554,N_14820,N_14549);
nand U16555 (N_16555,N_15851,N_14547);
nand U16556 (N_16556,N_15968,N_15373);
nand U16557 (N_16557,N_14974,N_14288);
xor U16558 (N_16558,N_15660,N_15718);
or U16559 (N_16559,N_15356,N_15835);
nand U16560 (N_16560,N_15023,N_14324);
xor U16561 (N_16561,N_14307,N_14991);
nand U16562 (N_16562,N_14888,N_15216);
or U16563 (N_16563,N_15691,N_15494);
nand U16564 (N_16564,N_15836,N_14306);
xnor U16565 (N_16565,N_15987,N_15260);
nand U16566 (N_16566,N_15303,N_14405);
nand U16567 (N_16567,N_15824,N_15890);
or U16568 (N_16568,N_15568,N_14859);
nor U16569 (N_16569,N_15739,N_15523);
nand U16570 (N_16570,N_14700,N_15914);
xor U16571 (N_16571,N_14084,N_14797);
nand U16572 (N_16572,N_15172,N_15332);
nand U16573 (N_16573,N_14867,N_14638);
or U16574 (N_16574,N_15753,N_14906);
or U16575 (N_16575,N_14140,N_15095);
or U16576 (N_16576,N_15031,N_14256);
nor U16577 (N_16577,N_14406,N_14915);
nor U16578 (N_16578,N_15918,N_15324);
nand U16579 (N_16579,N_14367,N_15747);
nand U16580 (N_16580,N_15702,N_14179);
xnor U16581 (N_16581,N_15723,N_14926);
xnor U16582 (N_16582,N_15946,N_15831);
nand U16583 (N_16583,N_14340,N_14196);
and U16584 (N_16584,N_14538,N_15257);
or U16585 (N_16585,N_14969,N_15538);
and U16586 (N_16586,N_15758,N_15226);
nand U16587 (N_16587,N_14318,N_14174);
and U16588 (N_16588,N_14896,N_15395);
nand U16589 (N_16589,N_14333,N_15231);
and U16590 (N_16590,N_14573,N_14029);
nand U16591 (N_16591,N_14047,N_15540);
nand U16592 (N_16592,N_14222,N_14077);
nand U16593 (N_16593,N_14132,N_14884);
or U16594 (N_16594,N_15543,N_15184);
and U16595 (N_16595,N_14596,N_14250);
nor U16596 (N_16596,N_14989,N_14672);
nor U16597 (N_16597,N_15104,N_15276);
and U16598 (N_16598,N_14094,N_15719);
or U16599 (N_16599,N_14811,N_14187);
nor U16600 (N_16600,N_14234,N_15663);
nor U16601 (N_16601,N_14010,N_15910);
or U16602 (N_16602,N_14916,N_14415);
nor U16603 (N_16603,N_15331,N_15300);
xor U16604 (N_16604,N_14659,N_14216);
nand U16605 (N_16605,N_15421,N_15759);
nor U16606 (N_16606,N_14227,N_15357);
nor U16607 (N_16607,N_14085,N_15223);
or U16608 (N_16608,N_15680,N_15090);
or U16609 (N_16609,N_14079,N_15412);
nand U16610 (N_16610,N_15926,N_15947);
and U16611 (N_16611,N_15009,N_14294);
xnor U16612 (N_16612,N_14592,N_14536);
and U16613 (N_16613,N_15014,N_15860);
nand U16614 (N_16614,N_15966,N_14474);
and U16615 (N_16615,N_15207,N_15291);
nor U16616 (N_16616,N_15791,N_15043);
and U16617 (N_16617,N_14328,N_14824);
and U16618 (N_16618,N_14252,N_14323);
or U16619 (N_16619,N_14505,N_15963);
nand U16620 (N_16620,N_15113,N_15477);
nand U16621 (N_16621,N_15754,N_15127);
and U16622 (N_16622,N_15870,N_15471);
nor U16623 (N_16623,N_15151,N_14992);
nor U16624 (N_16624,N_14118,N_14613);
nand U16625 (N_16625,N_14045,N_14448);
or U16626 (N_16626,N_15348,N_14732);
or U16627 (N_16627,N_14663,N_15981);
nor U16628 (N_16628,N_14518,N_14008);
nor U16629 (N_16629,N_14956,N_14524);
or U16630 (N_16630,N_15671,N_14770);
nor U16631 (N_16631,N_14220,N_15507);
and U16632 (N_16632,N_15635,N_14907);
or U16633 (N_16633,N_14781,N_15082);
and U16634 (N_16634,N_15837,N_14368);
nand U16635 (N_16635,N_15822,N_14218);
or U16636 (N_16636,N_15143,N_14545);
xnor U16637 (N_16637,N_15154,N_14332);
nor U16638 (N_16638,N_14263,N_14623);
nor U16639 (N_16639,N_14954,N_15600);
or U16640 (N_16640,N_14861,N_14848);
nand U16641 (N_16641,N_15131,N_14131);
and U16642 (N_16642,N_14532,N_15513);
or U16643 (N_16643,N_14034,N_14064);
xor U16644 (N_16644,N_15288,N_14068);
nand U16645 (N_16645,N_14927,N_14463);
or U16646 (N_16646,N_14237,N_15797);
and U16647 (N_16647,N_15969,N_15499);
or U16648 (N_16648,N_14319,N_15155);
nand U16649 (N_16649,N_15970,N_15602);
xor U16650 (N_16650,N_15509,N_15555);
and U16651 (N_16651,N_15778,N_15608);
nor U16652 (N_16652,N_14819,N_15334);
nand U16653 (N_16653,N_14616,N_14013);
nand U16654 (N_16654,N_14923,N_14909);
or U16655 (N_16655,N_15459,N_15849);
nor U16656 (N_16656,N_14818,N_14822);
and U16657 (N_16657,N_15549,N_14417);
or U16658 (N_16658,N_15230,N_15875);
xor U16659 (N_16659,N_14165,N_15519);
nor U16660 (N_16660,N_15666,N_15881);
nand U16661 (N_16661,N_15187,N_15765);
nor U16662 (N_16662,N_15585,N_15236);
nand U16663 (N_16663,N_14258,N_15447);
and U16664 (N_16664,N_15531,N_15038);
nand U16665 (N_16665,N_15442,N_14831);
or U16666 (N_16666,N_14632,N_15213);
and U16667 (N_16667,N_15279,N_15130);
and U16668 (N_16668,N_14481,N_14599);
and U16669 (N_16669,N_15980,N_15255);
and U16670 (N_16670,N_14155,N_14486);
or U16671 (N_16671,N_15603,N_14879);
or U16672 (N_16672,N_14944,N_14897);
nor U16673 (N_16673,N_15647,N_15083);
or U16674 (N_16674,N_14129,N_14240);
nor U16675 (N_16675,N_15582,N_14073);
nor U16676 (N_16676,N_14142,N_15263);
nor U16677 (N_16677,N_14141,N_14101);
or U16678 (N_16678,N_15529,N_15522);
nand U16679 (N_16679,N_15157,N_14295);
or U16680 (N_16680,N_14334,N_14836);
or U16681 (N_16681,N_14996,N_14661);
nand U16682 (N_16682,N_14705,N_14349);
or U16683 (N_16683,N_14656,N_14556);
nor U16684 (N_16684,N_15244,N_15182);
nor U16685 (N_16685,N_14893,N_14585);
nand U16686 (N_16686,N_15135,N_15854);
or U16687 (N_16687,N_14168,N_14550);
and U16688 (N_16688,N_14404,N_15394);
and U16689 (N_16689,N_15380,N_14135);
and U16690 (N_16690,N_14376,N_14724);
or U16691 (N_16691,N_14408,N_15594);
nand U16692 (N_16692,N_14175,N_14619);
or U16693 (N_16693,N_14387,N_14149);
nand U16694 (N_16694,N_15866,N_15933);
nor U16695 (N_16695,N_15071,N_15550);
nand U16696 (N_16696,N_15069,N_14640);
nand U16697 (N_16697,N_15343,N_15258);
nor U16698 (N_16698,N_15798,N_15793);
nand U16699 (N_16699,N_15052,N_15907);
nand U16700 (N_16700,N_14300,N_14675);
or U16701 (N_16701,N_15467,N_14497);
or U16702 (N_16702,N_14812,N_14862);
nor U16703 (N_16703,N_14056,N_14886);
and U16704 (N_16704,N_15445,N_15877);
nor U16705 (N_16705,N_15708,N_14790);
and U16706 (N_16706,N_14507,N_14383);
and U16707 (N_16707,N_15271,N_15629);
nand U16708 (N_16708,N_14358,N_14872);
nand U16709 (N_16709,N_15735,N_15662);
or U16710 (N_16710,N_15386,N_15563);
nor U16711 (N_16711,N_14500,N_15454);
xnor U16712 (N_16712,N_14152,N_14226);
and U16713 (N_16713,N_15385,N_15252);
xor U16714 (N_16714,N_15506,N_15820);
nand U16715 (N_16715,N_14645,N_14439);
nand U16716 (N_16716,N_14696,N_14071);
xnor U16717 (N_16717,N_14325,N_15807);
and U16718 (N_16718,N_14670,N_15714);
nor U16719 (N_16719,N_15924,N_15004);
nor U16720 (N_16720,N_15492,N_15282);
nand U16721 (N_16721,N_14096,N_14004);
and U16722 (N_16722,N_14351,N_14826);
or U16723 (N_16723,N_14628,N_14080);
and U16724 (N_16724,N_15478,N_15340);
nor U16725 (N_16725,N_14772,N_14666);
nor U16726 (N_16726,N_15285,N_14634);
nor U16727 (N_16727,N_15928,N_14553);
or U16728 (N_16728,N_15731,N_15436);
nand U16729 (N_16729,N_14423,N_15889);
nand U16730 (N_16730,N_15743,N_14115);
and U16731 (N_16731,N_14378,N_14445);
nand U16732 (N_16732,N_15353,N_14689);
xor U16733 (N_16733,N_15315,N_14682);
and U16734 (N_16734,N_14703,N_15080);
and U16735 (N_16735,N_15211,N_15354);
nor U16736 (N_16736,N_15796,N_15485);
or U16737 (N_16737,N_15534,N_15484);
or U16738 (N_16738,N_14588,N_14914);
or U16739 (N_16739,N_14032,N_15768);
nand U16740 (N_16740,N_14579,N_15652);
nand U16741 (N_16741,N_15106,N_14537);
nand U16742 (N_16742,N_14357,N_15913);
and U16743 (N_16743,N_15483,N_14430);
nand U16744 (N_16744,N_15287,N_14506);
and U16745 (N_16745,N_14583,N_15547);
or U16746 (N_16746,N_14706,N_15530);
or U16747 (N_16747,N_14401,N_14033);
and U16748 (N_16748,N_15586,N_14286);
or U16749 (N_16749,N_15645,N_15814);
nand U16750 (N_16750,N_15429,N_14070);
or U16751 (N_16751,N_14000,N_15808);
or U16752 (N_16752,N_15229,N_15916);
and U16753 (N_16753,N_15921,N_15440);
or U16754 (N_16754,N_15341,N_15581);
nand U16755 (N_16755,N_14971,N_14935);
nor U16756 (N_16756,N_15251,N_15780);
or U16757 (N_16757,N_15452,N_15888);
or U16758 (N_16758,N_14182,N_15116);
nor U16759 (N_16759,N_14467,N_14270);
nor U16760 (N_16760,N_15007,N_15225);
nand U16761 (N_16761,N_14875,N_15202);
nor U16762 (N_16762,N_15142,N_15943);
nor U16763 (N_16763,N_15899,N_14900);
nor U16764 (N_16764,N_15054,N_15533);
nor U16765 (N_16765,N_15319,N_14058);
xor U16766 (N_16766,N_15148,N_15119);
or U16767 (N_16767,N_14202,N_14124);
nand U16768 (N_16768,N_14191,N_14156);
nand U16769 (N_16769,N_15293,N_14646);
or U16770 (N_16770,N_15122,N_14241);
nor U16771 (N_16771,N_14163,N_15401);
or U16772 (N_16772,N_14894,N_15886);
or U16773 (N_16773,N_14254,N_14932);
nand U16774 (N_16774,N_15593,N_15569);
nor U16775 (N_16775,N_14939,N_14201);
and U16776 (N_16776,N_14814,N_14918);
xor U16777 (N_16777,N_15170,N_14809);
or U16778 (N_16778,N_15911,N_14597);
or U16779 (N_16779,N_15698,N_14395);
nand U16780 (N_16780,N_14083,N_14195);
or U16781 (N_16781,N_15596,N_15658);
or U16782 (N_16782,N_15699,N_14299);
nor U16783 (N_16783,N_15825,N_14607);
and U16784 (N_16784,N_15927,N_15619);
and U16785 (N_16785,N_14359,N_14074);
or U16786 (N_16786,N_14753,N_14688);
and U16787 (N_16787,N_15873,N_15432);
or U16788 (N_16788,N_15571,N_15715);
or U16789 (N_16789,N_15178,N_14472);
or U16790 (N_16790,N_15744,N_15991);
nand U16791 (N_16791,N_14921,N_14457);
nand U16792 (N_16792,N_15896,N_15247);
and U16793 (N_16793,N_14947,N_14562);
or U16794 (N_16794,N_14951,N_15517);
or U16795 (N_16795,N_14336,N_14396);
and U16796 (N_16796,N_15904,N_14671);
nand U16797 (N_16797,N_14154,N_15307);
nor U16798 (N_16798,N_15411,N_14994);
or U16799 (N_16799,N_15706,N_14289);
and U16800 (N_16800,N_15567,N_14015);
nor U16801 (N_16801,N_14062,N_14392);
nand U16802 (N_16802,N_14667,N_14983);
nor U16803 (N_16803,N_14504,N_15466);
nor U16804 (N_16804,N_14361,N_14239);
and U16805 (N_16805,N_15363,N_14356);
or U16806 (N_16806,N_15390,N_14958);
nand U16807 (N_16807,N_14925,N_15208);
and U16808 (N_16808,N_14026,N_15072);
or U16809 (N_16809,N_15013,N_14217);
xor U16810 (N_16810,N_14144,N_15784);
nand U16811 (N_16811,N_14544,N_15171);
or U16812 (N_16812,N_15266,N_14177);
and U16813 (N_16813,N_14622,N_15992);
nand U16814 (N_16814,N_15573,N_15316);
nor U16815 (N_16815,N_14513,N_14889);
and U16816 (N_16816,N_15210,N_14194);
xnor U16817 (N_16817,N_14817,N_14558);
nand U16818 (N_16818,N_14563,N_15201);
nand U16819 (N_16819,N_15693,N_14012);
nor U16820 (N_16820,N_14260,N_14117);
and U16821 (N_16821,N_14440,N_15685);
xnor U16822 (N_16822,N_14869,N_14134);
nand U16823 (N_16823,N_15624,N_14712);
nand U16824 (N_16824,N_14674,N_14365);
nand U16825 (N_16825,N_15572,N_14102);
nand U16826 (N_16826,N_15614,N_14366);
or U16827 (N_16827,N_15370,N_15591);
nor U16828 (N_16828,N_14615,N_14473);
and U16829 (N_16829,N_15379,N_15423);
nand U16830 (N_16830,N_14948,N_15818);
and U16831 (N_16831,N_15772,N_15015);
nor U16832 (N_16832,N_15730,N_15557);
and U16833 (N_16833,N_14210,N_14752);
and U16834 (N_16834,N_15616,N_15812);
nor U16835 (N_16835,N_14561,N_15965);
xor U16836 (N_16836,N_14143,N_15536);
nand U16837 (N_16837,N_14470,N_14173);
and U16838 (N_16838,N_14309,N_15190);
nor U16839 (N_16839,N_15542,N_14644);
nor U16840 (N_16840,N_15239,N_15221);
or U16841 (N_16841,N_15590,N_14052);
or U16842 (N_16842,N_15105,N_15419);
and U16843 (N_16843,N_14292,N_15146);
nor U16844 (N_16844,N_15081,N_14999);
or U16845 (N_16845,N_14726,N_15655);
nor U16846 (N_16846,N_15060,N_15149);
and U16847 (N_16847,N_15960,N_15048);
or U16848 (N_16848,N_15117,N_14778);
nor U16849 (N_16849,N_14345,N_15493);
or U16850 (N_16850,N_14046,N_14866);
or U16851 (N_16851,N_14127,N_14995);
or U16852 (N_16852,N_15871,N_15134);
nand U16853 (N_16853,N_15321,N_14528);
nor U16854 (N_16854,N_14018,N_15973);
and U16855 (N_16855,N_15510,N_14934);
nand U16856 (N_16856,N_14427,N_15941);
or U16857 (N_16857,N_15346,N_14446);
nand U16858 (N_16858,N_14761,N_15057);
xnor U16859 (N_16859,N_15682,N_15657);
and U16860 (N_16860,N_15275,N_15397);
and U16861 (N_16861,N_14360,N_14452);
or U16862 (N_16862,N_14125,N_14608);
nand U16863 (N_16863,N_15035,N_15242);
nor U16864 (N_16864,N_14780,N_14432);
nand U16865 (N_16865,N_14711,N_14180);
nand U16866 (N_16866,N_15002,N_14572);
or U16867 (N_16867,N_15369,N_14038);
and U16868 (N_16868,N_15188,N_14110);
and U16869 (N_16869,N_15786,N_14564);
and U16870 (N_16870,N_14901,N_14499);
nor U16871 (N_16871,N_15186,N_15045);
and U16872 (N_16872,N_14979,N_14414);
nand U16873 (N_16873,N_14933,N_15716);
nand U16874 (N_16874,N_15834,N_14741);
nor U16875 (N_16875,N_14710,N_15215);
and U16876 (N_16876,N_14860,N_14257);
and U16877 (N_16877,N_14343,N_14610);
nor U16878 (N_16878,N_15701,N_14620);
nor U16879 (N_16879,N_14699,N_15915);
nand U16880 (N_16880,N_15418,N_15443);
nand U16881 (N_16881,N_15689,N_15200);
and U16882 (N_16882,N_14093,N_15003);
nand U16883 (N_16883,N_14089,N_15604);
nor U16884 (N_16884,N_15360,N_15817);
and U16885 (N_16885,N_14316,N_15391);
nor U16886 (N_16886,N_14841,N_15885);
nand U16887 (N_16887,N_14211,N_15317);
nor U16888 (N_16888,N_15199,N_14464);
or U16889 (N_16889,N_15163,N_14485);
nand U16890 (N_16890,N_14966,N_14502);
or U16891 (N_16891,N_15245,N_14985);
and U16892 (N_16892,N_14511,N_15776);
nand U16893 (N_16893,N_15878,N_14851);
or U16894 (N_16894,N_15058,N_14475);
or U16895 (N_16895,N_15688,N_14924);
or U16896 (N_16896,N_14053,N_15384);
nor U16897 (N_16897,N_15917,N_14166);
or U16898 (N_16898,N_14479,N_15535);
nand U16899 (N_16899,N_14704,N_15311);
nand U16900 (N_16900,N_14833,N_15905);
and U16901 (N_16901,N_15037,N_14776);
nor U16902 (N_16902,N_15707,N_14450);
and U16903 (N_16903,N_14881,N_15181);
nor U16904 (N_16904,N_15939,N_14023);
nand U16905 (N_16905,N_14049,N_15696);
or U16906 (N_16906,N_15501,N_14521);
nor U16907 (N_16907,N_15988,N_14530);
nand U16908 (N_16908,N_15020,N_14567);
nor U16909 (N_16909,N_15296,N_14005);
nor U16910 (N_16910,N_14385,N_15272);
nand U16911 (N_16911,N_14943,N_14527);
and U16912 (N_16912,N_15996,N_14715);
nand U16913 (N_16913,N_15480,N_15527);
xnor U16914 (N_16914,N_14783,N_14793);
nand U16915 (N_16915,N_14658,N_15920);
nand U16916 (N_16916,N_14938,N_15195);
xor U16917 (N_16917,N_15158,N_15695);
and U16918 (N_16918,N_15556,N_15580);
and U16919 (N_16919,N_15667,N_15472);
nand U16920 (N_16920,N_15396,N_14798);
and U16921 (N_16921,N_14020,N_15502);
or U16922 (N_16922,N_15099,N_15736);
nand U16923 (N_16923,N_15990,N_14631);
nor U16924 (N_16924,N_15843,N_15050);
and U16925 (N_16925,N_14762,N_15096);
or U16926 (N_16926,N_15240,N_15733);
and U16927 (N_16927,N_15192,N_14695);
and U16928 (N_16928,N_15259,N_14601);
or U16929 (N_16929,N_14305,N_14431);
and U16930 (N_16930,N_14436,N_14691);
nor U16931 (N_16931,N_15631,N_14764);
and U16932 (N_16932,N_15623,N_14429);
and U16933 (N_16933,N_15774,N_15967);
nand U16934 (N_16934,N_15308,N_15654);
xnor U16935 (N_16935,N_15120,N_15977);
and U16936 (N_16936,N_14908,N_14238);
xnor U16937 (N_16937,N_14402,N_14208);
nand U16938 (N_16938,N_14287,N_15371);
nand U16939 (N_16939,N_14560,N_15294);
nand U16940 (N_16940,N_15457,N_15070);
xnor U16941 (N_16941,N_14224,N_14341);
xor U16942 (N_16942,N_14660,N_14773);
and U16943 (N_16943,N_14930,N_14055);
or U16944 (N_16944,N_15687,N_15800);
and U16945 (N_16945,N_14785,N_15964);
nor U16946 (N_16946,N_14982,N_14730);
xor U16947 (N_16947,N_14960,N_14229);
nand U16948 (N_16948,N_14498,N_15029);
or U16949 (N_16949,N_14858,N_15565);
nor U16950 (N_16950,N_15233,N_14605);
and U16951 (N_16951,N_14586,N_14204);
and U16952 (N_16952,N_15306,N_15422);
or U16953 (N_16953,N_14390,N_14057);
and U16954 (N_16954,N_15592,N_15312);
or U16955 (N_16955,N_15833,N_14384);
nand U16956 (N_16956,N_14576,N_15302);
nand U16957 (N_16957,N_14978,N_14542);
or U16958 (N_16958,N_14069,N_14686);
and U16959 (N_16959,N_15930,N_15497);
nor U16960 (N_16960,N_14331,N_15160);
nor U16961 (N_16961,N_15448,N_15329);
or U16962 (N_16962,N_14233,N_14868);
or U16963 (N_16963,N_14618,N_14929);
or U16964 (N_16964,N_15222,N_15518);
nand U16965 (N_16965,N_15801,N_15284);
xor U16966 (N_16966,N_15717,N_15444);
or U16967 (N_16967,N_14687,N_14534);
or U16968 (N_16968,N_14664,N_14959);
and U16969 (N_16969,N_15732,N_14743);
nand U16970 (N_16970,N_14067,N_15504);
and U16971 (N_16971,N_14072,N_14832);
and U16972 (N_16972,N_15897,N_15268);
xnor U16973 (N_16973,N_15161,N_15882);
and U16974 (N_16974,N_15362,N_14769);
xnor U16975 (N_16975,N_15898,N_15169);
and U16976 (N_16976,N_15304,N_14775);
and U16977 (N_16977,N_14952,N_14821);
or U16978 (N_16978,N_14800,N_15879);
or U16979 (N_16979,N_15248,N_15803);
and U16980 (N_16980,N_14830,N_14184);
or U16981 (N_16981,N_14668,N_14751);
and U16982 (N_16982,N_14512,N_15601);
and U16983 (N_16983,N_15972,N_14796);
xor U16984 (N_16984,N_14011,N_14657);
and U16985 (N_16985,N_14855,N_14267);
or U16986 (N_16986,N_14098,N_14181);
or U16987 (N_16987,N_15409,N_14853);
xor U16988 (N_16988,N_15085,N_14490);
and U16989 (N_16989,N_15217,N_14998);
and U16990 (N_16990,N_14480,N_15238);
nor U16991 (N_16991,N_15344,N_15922);
and U16992 (N_16992,N_14749,N_15093);
nand U16993 (N_16993,N_14460,N_14988);
nand U16994 (N_16994,N_14531,N_14425);
or U16995 (N_16995,N_15976,N_15958);
or U16996 (N_16996,N_14852,N_14625);
and U16997 (N_16997,N_14364,N_15297);
nor U16998 (N_16998,N_14736,N_15528);
or U16999 (N_16999,N_15640,N_15061);
or U17000 (N_17000,N_15625,N_15312);
or U17001 (N_17001,N_15328,N_15873);
nand U17002 (N_17002,N_14760,N_14466);
nor U17003 (N_17003,N_14224,N_15217);
nor U17004 (N_17004,N_15815,N_14979);
and U17005 (N_17005,N_14717,N_14216);
or U17006 (N_17006,N_14647,N_15398);
nor U17007 (N_17007,N_15498,N_14846);
nor U17008 (N_17008,N_14072,N_15587);
and U17009 (N_17009,N_14968,N_14954);
nand U17010 (N_17010,N_15755,N_14491);
nor U17011 (N_17011,N_15673,N_15838);
nor U17012 (N_17012,N_15009,N_14111);
nand U17013 (N_17013,N_15769,N_14239);
nand U17014 (N_17014,N_14237,N_15893);
xor U17015 (N_17015,N_15354,N_14095);
and U17016 (N_17016,N_14609,N_15659);
or U17017 (N_17017,N_14626,N_14265);
nor U17018 (N_17018,N_15764,N_15312);
nor U17019 (N_17019,N_15287,N_15118);
nor U17020 (N_17020,N_15442,N_14625);
xor U17021 (N_17021,N_15062,N_14536);
and U17022 (N_17022,N_14733,N_14284);
or U17023 (N_17023,N_14579,N_14367);
nand U17024 (N_17024,N_14599,N_14983);
and U17025 (N_17025,N_14884,N_15061);
nand U17026 (N_17026,N_14700,N_15151);
nand U17027 (N_17027,N_15663,N_14209);
nand U17028 (N_17028,N_15280,N_15106);
or U17029 (N_17029,N_14552,N_14165);
nor U17030 (N_17030,N_14050,N_15520);
nor U17031 (N_17031,N_15065,N_14905);
nand U17032 (N_17032,N_14934,N_14845);
nor U17033 (N_17033,N_14162,N_15853);
or U17034 (N_17034,N_15036,N_14365);
xnor U17035 (N_17035,N_14014,N_14053);
nor U17036 (N_17036,N_15769,N_14275);
or U17037 (N_17037,N_15427,N_14652);
or U17038 (N_17038,N_15216,N_14015);
nand U17039 (N_17039,N_15068,N_15368);
nor U17040 (N_17040,N_15957,N_14704);
and U17041 (N_17041,N_15668,N_14794);
and U17042 (N_17042,N_15862,N_15636);
nand U17043 (N_17043,N_15633,N_14707);
nor U17044 (N_17044,N_14976,N_14398);
and U17045 (N_17045,N_14219,N_15309);
nand U17046 (N_17046,N_15789,N_14145);
xor U17047 (N_17047,N_15828,N_14304);
or U17048 (N_17048,N_14928,N_15680);
nand U17049 (N_17049,N_15790,N_15288);
or U17050 (N_17050,N_14417,N_15723);
or U17051 (N_17051,N_15469,N_15375);
or U17052 (N_17052,N_14098,N_14871);
nor U17053 (N_17053,N_15970,N_14954);
nand U17054 (N_17054,N_15623,N_15719);
nand U17055 (N_17055,N_15262,N_14205);
or U17056 (N_17056,N_15374,N_15409);
nand U17057 (N_17057,N_15890,N_15010);
nand U17058 (N_17058,N_15490,N_15892);
nand U17059 (N_17059,N_14866,N_15030);
nor U17060 (N_17060,N_15686,N_14600);
nor U17061 (N_17061,N_14275,N_15601);
and U17062 (N_17062,N_15343,N_14134);
or U17063 (N_17063,N_15743,N_14729);
nor U17064 (N_17064,N_15610,N_15275);
nand U17065 (N_17065,N_14495,N_14339);
or U17066 (N_17066,N_14901,N_14913);
xnor U17067 (N_17067,N_14842,N_14235);
nand U17068 (N_17068,N_14779,N_14077);
and U17069 (N_17069,N_14478,N_14774);
nor U17070 (N_17070,N_15660,N_14036);
and U17071 (N_17071,N_15026,N_14012);
or U17072 (N_17072,N_14068,N_14208);
and U17073 (N_17073,N_14725,N_14356);
and U17074 (N_17074,N_14610,N_14883);
nor U17075 (N_17075,N_14700,N_14056);
and U17076 (N_17076,N_14694,N_14512);
nand U17077 (N_17077,N_15500,N_15462);
nor U17078 (N_17078,N_14316,N_15304);
nand U17079 (N_17079,N_15106,N_14930);
and U17080 (N_17080,N_14794,N_15949);
nor U17081 (N_17081,N_15977,N_14989);
nor U17082 (N_17082,N_14878,N_15154);
nor U17083 (N_17083,N_15842,N_15650);
or U17084 (N_17084,N_15761,N_14124);
or U17085 (N_17085,N_15557,N_14361);
or U17086 (N_17086,N_15113,N_14583);
and U17087 (N_17087,N_15502,N_14429);
nand U17088 (N_17088,N_15972,N_14213);
or U17089 (N_17089,N_15917,N_15576);
nor U17090 (N_17090,N_15985,N_15884);
xnor U17091 (N_17091,N_15082,N_15514);
and U17092 (N_17092,N_15139,N_15222);
nand U17093 (N_17093,N_15511,N_14169);
or U17094 (N_17094,N_14980,N_15116);
and U17095 (N_17095,N_14851,N_15072);
nor U17096 (N_17096,N_15426,N_15258);
nand U17097 (N_17097,N_14894,N_15251);
or U17098 (N_17098,N_14365,N_14997);
nor U17099 (N_17099,N_14322,N_14513);
or U17100 (N_17100,N_14911,N_14165);
nor U17101 (N_17101,N_14689,N_14040);
nand U17102 (N_17102,N_14742,N_14907);
and U17103 (N_17103,N_15570,N_14123);
xnor U17104 (N_17104,N_14808,N_14443);
nor U17105 (N_17105,N_15214,N_15838);
nand U17106 (N_17106,N_14490,N_14749);
nand U17107 (N_17107,N_14096,N_14386);
and U17108 (N_17108,N_15133,N_15100);
nand U17109 (N_17109,N_14265,N_15742);
and U17110 (N_17110,N_15458,N_14200);
nor U17111 (N_17111,N_15925,N_15731);
and U17112 (N_17112,N_15350,N_14349);
nand U17113 (N_17113,N_14012,N_14335);
xor U17114 (N_17114,N_15929,N_15830);
nor U17115 (N_17115,N_15803,N_14851);
and U17116 (N_17116,N_15214,N_14132);
or U17117 (N_17117,N_14307,N_14472);
nor U17118 (N_17118,N_15604,N_15869);
nor U17119 (N_17119,N_14324,N_14669);
or U17120 (N_17120,N_15014,N_14104);
and U17121 (N_17121,N_14132,N_14445);
or U17122 (N_17122,N_15644,N_14826);
nand U17123 (N_17123,N_15578,N_15134);
xor U17124 (N_17124,N_14911,N_14356);
and U17125 (N_17125,N_15764,N_14588);
xnor U17126 (N_17126,N_14622,N_15820);
or U17127 (N_17127,N_15315,N_14982);
nor U17128 (N_17128,N_14843,N_15016);
and U17129 (N_17129,N_15408,N_14753);
or U17130 (N_17130,N_15030,N_14781);
nor U17131 (N_17131,N_14092,N_15808);
nand U17132 (N_17132,N_14185,N_15185);
or U17133 (N_17133,N_15358,N_14461);
nor U17134 (N_17134,N_14741,N_15143);
nand U17135 (N_17135,N_14863,N_14865);
or U17136 (N_17136,N_14690,N_15989);
nand U17137 (N_17137,N_14529,N_15002);
nor U17138 (N_17138,N_15756,N_14857);
and U17139 (N_17139,N_14121,N_15001);
or U17140 (N_17140,N_15301,N_15981);
nor U17141 (N_17141,N_14561,N_14778);
xnor U17142 (N_17142,N_14984,N_14284);
or U17143 (N_17143,N_15807,N_14286);
nand U17144 (N_17144,N_14256,N_14112);
nor U17145 (N_17145,N_14203,N_15632);
or U17146 (N_17146,N_15393,N_14541);
nand U17147 (N_17147,N_14793,N_15936);
nand U17148 (N_17148,N_14769,N_15929);
or U17149 (N_17149,N_14802,N_14749);
nor U17150 (N_17150,N_14155,N_15512);
or U17151 (N_17151,N_15985,N_15925);
and U17152 (N_17152,N_14620,N_15351);
or U17153 (N_17153,N_15766,N_15155);
and U17154 (N_17154,N_15520,N_14997);
or U17155 (N_17155,N_15107,N_14526);
nor U17156 (N_17156,N_14342,N_15922);
nor U17157 (N_17157,N_14708,N_14080);
and U17158 (N_17158,N_14036,N_15074);
or U17159 (N_17159,N_15646,N_15123);
nand U17160 (N_17160,N_14608,N_15424);
nor U17161 (N_17161,N_15100,N_14482);
nor U17162 (N_17162,N_14708,N_15150);
nand U17163 (N_17163,N_14864,N_15363);
and U17164 (N_17164,N_14100,N_14067);
or U17165 (N_17165,N_14084,N_15640);
or U17166 (N_17166,N_15665,N_15391);
xor U17167 (N_17167,N_14514,N_15972);
nor U17168 (N_17168,N_15715,N_14690);
and U17169 (N_17169,N_14758,N_14646);
or U17170 (N_17170,N_15466,N_14501);
or U17171 (N_17171,N_14992,N_14975);
nor U17172 (N_17172,N_14807,N_14854);
nand U17173 (N_17173,N_14022,N_14711);
or U17174 (N_17174,N_15231,N_14567);
and U17175 (N_17175,N_15845,N_15684);
xor U17176 (N_17176,N_15095,N_15317);
and U17177 (N_17177,N_14010,N_15442);
nand U17178 (N_17178,N_14112,N_14500);
nand U17179 (N_17179,N_14718,N_14416);
nand U17180 (N_17180,N_15668,N_14778);
nand U17181 (N_17181,N_15915,N_14289);
nand U17182 (N_17182,N_14518,N_14886);
xor U17183 (N_17183,N_14459,N_15069);
xor U17184 (N_17184,N_14930,N_15041);
xnor U17185 (N_17185,N_15085,N_14928);
nor U17186 (N_17186,N_15528,N_14879);
nor U17187 (N_17187,N_14415,N_14983);
xor U17188 (N_17188,N_15263,N_14823);
nor U17189 (N_17189,N_15280,N_15387);
and U17190 (N_17190,N_15215,N_15497);
nor U17191 (N_17191,N_14553,N_14819);
and U17192 (N_17192,N_14840,N_14499);
or U17193 (N_17193,N_14704,N_15689);
nand U17194 (N_17194,N_14557,N_14848);
or U17195 (N_17195,N_15348,N_14730);
nand U17196 (N_17196,N_15060,N_14881);
nor U17197 (N_17197,N_14743,N_15745);
or U17198 (N_17198,N_15204,N_14033);
nor U17199 (N_17199,N_15373,N_14764);
and U17200 (N_17200,N_15682,N_14838);
nor U17201 (N_17201,N_15360,N_14215);
nand U17202 (N_17202,N_14875,N_14192);
and U17203 (N_17203,N_15158,N_14486);
xor U17204 (N_17204,N_15650,N_14976);
nand U17205 (N_17205,N_14468,N_15919);
and U17206 (N_17206,N_14665,N_14173);
nand U17207 (N_17207,N_14084,N_15148);
and U17208 (N_17208,N_14301,N_14989);
xor U17209 (N_17209,N_14891,N_14707);
nand U17210 (N_17210,N_14385,N_14780);
nor U17211 (N_17211,N_14032,N_15451);
or U17212 (N_17212,N_14441,N_15654);
nor U17213 (N_17213,N_14452,N_15393);
and U17214 (N_17214,N_15146,N_15406);
nor U17215 (N_17215,N_14179,N_15438);
nor U17216 (N_17216,N_14267,N_14613);
nand U17217 (N_17217,N_14300,N_14713);
nand U17218 (N_17218,N_15292,N_14098);
nor U17219 (N_17219,N_14876,N_15870);
and U17220 (N_17220,N_15339,N_14453);
and U17221 (N_17221,N_14143,N_14437);
and U17222 (N_17222,N_14466,N_14449);
nand U17223 (N_17223,N_14046,N_15981);
nand U17224 (N_17224,N_15357,N_15302);
nand U17225 (N_17225,N_15172,N_15013);
xor U17226 (N_17226,N_15710,N_14408);
nor U17227 (N_17227,N_14132,N_14863);
and U17228 (N_17228,N_15783,N_15071);
and U17229 (N_17229,N_14631,N_14015);
nor U17230 (N_17230,N_15351,N_15389);
or U17231 (N_17231,N_14245,N_15414);
nor U17232 (N_17232,N_14900,N_14713);
nor U17233 (N_17233,N_15384,N_15707);
nor U17234 (N_17234,N_14891,N_15571);
nor U17235 (N_17235,N_15354,N_14862);
xor U17236 (N_17236,N_14424,N_15295);
and U17237 (N_17237,N_14221,N_15481);
or U17238 (N_17238,N_15484,N_15827);
and U17239 (N_17239,N_15784,N_14375);
nand U17240 (N_17240,N_14156,N_14099);
nor U17241 (N_17241,N_15400,N_14324);
or U17242 (N_17242,N_15182,N_15835);
xnor U17243 (N_17243,N_14285,N_15615);
or U17244 (N_17244,N_15648,N_14923);
or U17245 (N_17245,N_15453,N_14742);
xor U17246 (N_17246,N_15826,N_15669);
and U17247 (N_17247,N_14213,N_15904);
or U17248 (N_17248,N_15257,N_15858);
nand U17249 (N_17249,N_15874,N_14741);
and U17250 (N_17250,N_14312,N_14886);
nor U17251 (N_17251,N_15939,N_14227);
nor U17252 (N_17252,N_14013,N_14108);
xnor U17253 (N_17253,N_15211,N_15067);
or U17254 (N_17254,N_14979,N_15843);
or U17255 (N_17255,N_15763,N_15203);
nand U17256 (N_17256,N_14632,N_15240);
nand U17257 (N_17257,N_15148,N_14137);
nand U17258 (N_17258,N_15225,N_15985);
and U17259 (N_17259,N_14054,N_14536);
and U17260 (N_17260,N_15659,N_14289);
and U17261 (N_17261,N_15729,N_14486);
or U17262 (N_17262,N_14332,N_15994);
nor U17263 (N_17263,N_14086,N_14323);
and U17264 (N_17264,N_14242,N_15369);
nand U17265 (N_17265,N_15237,N_14199);
nand U17266 (N_17266,N_15264,N_15091);
or U17267 (N_17267,N_15758,N_14438);
or U17268 (N_17268,N_15424,N_15529);
and U17269 (N_17269,N_15779,N_14914);
or U17270 (N_17270,N_15317,N_14794);
xnor U17271 (N_17271,N_15065,N_15320);
nand U17272 (N_17272,N_15706,N_15539);
and U17273 (N_17273,N_14412,N_14611);
nor U17274 (N_17274,N_14026,N_15265);
nand U17275 (N_17275,N_15607,N_14559);
or U17276 (N_17276,N_14527,N_14571);
nand U17277 (N_17277,N_15871,N_14685);
and U17278 (N_17278,N_15846,N_14336);
or U17279 (N_17279,N_14263,N_14124);
and U17280 (N_17280,N_14672,N_15164);
nand U17281 (N_17281,N_14475,N_14867);
nor U17282 (N_17282,N_14594,N_15645);
nand U17283 (N_17283,N_15548,N_14005);
nand U17284 (N_17284,N_15991,N_14582);
and U17285 (N_17285,N_14831,N_14817);
and U17286 (N_17286,N_15845,N_14047);
xor U17287 (N_17287,N_14600,N_14425);
nor U17288 (N_17288,N_14027,N_15368);
and U17289 (N_17289,N_14849,N_15717);
and U17290 (N_17290,N_14656,N_15804);
nand U17291 (N_17291,N_15626,N_14929);
and U17292 (N_17292,N_15230,N_15927);
nand U17293 (N_17293,N_15566,N_14910);
or U17294 (N_17294,N_15331,N_15371);
nor U17295 (N_17295,N_15396,N_15011);
nand U17296 (N_17296,N_14541,N_15104);
or U17297 (N_17297,N_15028,N_15571);
or U17298 (N_17298,N_14069,N_14457);
nand U17299 (N_17299,N_15211,N_15560);
or U17300 (N_17300,N_15235,N_14521);
and U17301 (N_17301,N_15273,N_14238);
xnor U17302 (N_17302,N_15729,N_15299);
xor U17303 (N_17303,N_15076,N_14162);
nor U17304 (N_17304,N_14664,N_15007);
xnor U17305 (N_17305,N_14944,N_14548);
and U17306 (N_17306,N_14667,N_14467);
or U17307 (N_17307,N_15400,N_15583);
and U17308 (N_17308,N_14598,N_15888);
nand U17309 (N_17309,N_15007,N_15050);
nor U17310 (N_17310,N_15768,N_15670);
nor U17311 (N_17311,N_15544,N_15152);
nand U17312 (N_17312,N_15858,N_14094);
or U17313 (N_17313,N_14841,N_15043);
and U17314 (N_17314,N_14874,N_15033);
or U17315 (N_17315,N_14836,N_15545);
xor U17316 (N_17316,N_15359,N_15530);
or U17317 (N_17317,N_15217,N_15524);
and U17318 (N_17318,N_15322,N_15088);
xnor U17319 (N_17319,N_14417,N_15491);
and U17320 (N_17320,N_15115,N_15673);
nor U17321 (N_17321,N_14570,N_15399);
nor U17322 (N_17322,N_14860,N_15372);
or U17323 (N_17323,N_14714,N_14020);
nand U17324 (N_17324,N_15508,N_14453);
nand U17325 (N_17325,N_14217,N_15705);
nor U17326 (N_17326,N_15656,N_15821);
and U17327 (N_17327,N_14304,N_14917);
nor U17328 (N_17328,N_15666,N_14622);
nor U17329 (N_17329,N_14703,N_15905);
and U17330 (N_17330,N_14108,N_15967);
nand U17331 (N_17331,N_15478,N_15809);
nor U17332 (N_17332,N_14092,N_15208);
nor U17333 (N_17333,N_15666,N_14787);
and U17334 (N_17334,N_15683,N_14543);
nor U17335 (N_17335,N_14610,N_15817);
and U17336 (N_17336,N_15656,N_15265);
and U17337 (N_17337,N_15917,N_14207);
or U17338 (N_17338,N_14459,N_15337);
and U17339 (N_17339,N_15760,N_15344);
and U17340 (N_17340,N_15034,N_15470);
or U17341 (N_17341,N_14567,N_14786);
or U17342 (N_17342,N_15198,N_15153);
nor U17343 (N_17343,N_15063,N_14142);
or U17344 (N_17344,N_15824,N_15502);
and U17345 (N_17345,N_15504,N_15068);
or U17346 (N_17346,N_14107,N_14715);
nor U17347 (N_17347,N_15094,N_14490);
and U17348 (N_17348,N_14275,N_14564);
nor U17349 (N_17349,N_14630,N_15130);
nand U17350 (N_17350,N_14922,N_14155);
or U17351 (N_17351,N_15655,N_14933);
nor U17352 (N_17352,N_15002,N_14802);
nand U17353 (N_17353,N_15964,N_15021);
xor U17354 (N_17354,N_14503,N_15877);
nor U17355 (N_17355,N_15740,N_15814);
nor U17356 (N_17356,N_15298,N_14085);
or U17357 (N_17357,N_15785,N_15599);
nand U17358 (N_17358,N_14622,N_15971);
or U17359 (N_17359,N_14748,N_14302);
or U17360 (N_17360,N_15759,N_15669);
nor U17361 (N_17361,N_15818,N_15149);
xnor U17362 (N_17362,N_15134,N_14167);
nor U17363 (N_17363,N_14517,N_14722);
nand U17364 (N_17364,N_15580,N_15280);
or U17365 (N_17365,N_15682,N_15081);
xnor U17366 (N_17366,N_15043,N_14572);
nand U17367 (N_17367,N_14592,N_14319);
or U17368 (N_17368,N_14713,N_14279);
and U17369 (N_17369,N_14496,N_14807);
nand U17370 (N_17370,N_14068,N_14203);
nor U17371 (N_17371,N_15454,N_15915);
or U17372 (N_17372,N_15456,N_15532);
nand U17373 (N_17373,N_15002,N_15168);
xnor U17374 (N_17374,N_15357,N_14432);
nor U17375 (N_17375,N_14840,N_14433);
nor U17376 (N_17376,N_14648,N_14027);
or U17377 (N_17377,N_15508,N_14520);
and U17378 (N_17378,N_14937,N_15098);
nor U17379 (N_17379,N_15770,N_15366);
and U17380 (N_17380,N_14276,N_15164);
and U17381 (N_17381,N_14186,N_15695);
nor U17382 (N_17382,N_15991,N_15977);
nand U17383 (N_17383,N_14887,N_15840);
nand U17384 (N_17384,N_14521,N_14686);
and U17385 (N_17385,N_15535,N_15720);
and U17386 (N_17386,N_15446,N_14850);
xnor U17387 (N_17387,N_15895,N_14319);
or U17388 (N_17388,N_15221,N_14558);
and U17389 (N_17389,N_14178,N_15181);
or U17390 (N_17390,N_15073,N_15313);
or U17391 (N_17391,N_15971,N_14895);
nand U17392 (N_17392,N_15766,N_15271);
or U17393 (N_17393,N_14732,N_15978);
nor U17394 (N_17394,N_15611,N_15325);
or U17395 (N_17395,N_14557,N_14432);
xnor U17396 (N_17396,N_15712,N_15217);
or U17397 (N_17397,N_15347,N_15543);
nand U17398 (N_17398,N_14854,N_15696);
nor U17399 (N_17399,N_15389,N_14731);
nor U17400 (N_17400,N_14968,N_15179);
nor U17401 (N_17401,N_14152,N_15692);
xnor U17402 (N_17402,N_15613,N_14296);
nor U17403 (N_17403,N_15472,N_15389);
or U17404 (N_17404,N_15250,N_14681);
or U17405 (N_17405,N_14572,N_15906);
nand U17406 (N_17406,N_15209,N_15473);
or U17407 (N_17407,N_15067,N_15501);
nand U17408 (N_17408,N_14267,N_14629);
or U17409 (N_17409,N_14360,N_14070);
and U17410 (N_17410,N_14273,N_15924);
nor U17411 (N_17411,N_14943,N_15501);
nor U17412 (N_17412,N_15626,N_15123);
and U17413 (N_17413,N_14260,N_14253);
and U17414 (N_17414,N_14477,N_14866);
nand U17415 (N_17415,N_15300,N_15479);
nand U17416 (N_17416,N_14275,N_15453);
nor U17417 (N_17417,N_14950,N_15371);
nand U17418 (N_17418,N_14033,N_15978);
and U17419 (N_17419,N_14000,N_14937);
nor U17420 (N_17420,N_14623,N_14586);
nor U17421 (N_17421,N_14848,N_15932);
or U17422 (N_17422,N_15231,N_15257);
and U17423 (N_17423,N_15300,N_14229);
and U17424 (N_17424,N_14325,N_14793);
nand U17425 (N_17425,N_15839,N_14370);
nor U17426 (N_17426,N_14736,N_14478);
and U17427 (N_17427,N_14449,N_14730);
xor U17428 (N_17428,N_15933,N_14573);
xor U17429 (N_17429,N_14554,N_14483);
nand U17430 (N_17430,N_15424,N_14136);
or U17431 (N_17431,N_14025,N_14755);
xor U17432 (N_17432,N_14042,N_15705);
and U17433 (N_17433,N_14246,N_15214);
nand U17434 (N_17434,N_14142,N_14298);
nor U17435 (N_17435,N_15050,N_14287);
or U17436 (N_17436,N_14596,N_15233);
nand U17437 (N_17437,N_15240,N_14481);
xnor U17438 (N_17438,N_15354,N_14108);
nand U17439 (N_17439,N_14749,N_15583);
or U17440 (N_17440,N_14842,N_15859);
or U17441 (N_17441,N_15531,N_15070);
and U17442 (N_17442,N_14489,N_15548);
or U17443 (N_17443,N_14437,N_15501);
nor U17444 (N_17444,N_14901,N_15137);
nand U17445 (N_17445,N_15041,N_14758);
and U17446 (N_17446,N_14329,N_14500);
and U17447 (N_17447,N_14946,N_14025);
nand U17448 (N_17448,N_14166,N_15997);
and U17449 (N_17449,N_15180,N_14659);
and U17450 (N_17450,N_14126,N_14661);
nand U17451 (N_17451,N_14941,N_15754);
and U17452 (N_17452,N_14413,N_15692);
and U17453 (N_17453,N_15627,N_14033);
and U17454 (N_17454,N_15539,N_15026);
nor U17455 (N_17455,N_14901,N_15371);
and U17456 (N_17456,N_15196,N_15124);
and U17457 (N_17457,N_15503,N_14187);
and U17458 (N_17458,N_15087,N_14924);
xor U17459 (N_17459,N_15384,N_14370);
or U17460 (N_17460,N_15293,N_14844);
or U17461 (N_17461,N_15336,N_14663);
and U17462 (N_17462,N_15447,N_14002);
nor U17463 (N_17463,N_15525,N_15613);
or U17464 (N_17464,N_15494,N_14084);
and U17465 (N_17465,N_14985,N_14100);
or U17466 (N_17466,N_14988,N_15902);
or U17467 (N_17467,N_14142,N_15100);
nor U17468 (N_17468,N_14881,N_15737);
and U17469 (N_17469,N_15844,N_15721);
or U17470 (N_17470,N_14030,N_14092);
xor U17471 (N_17471,N_15135,N_15430);
or U17472 (N_17472,N_14261,N_15262);
or U17473 (N_17473,N_15458,N_14492);
nand U17474 (N_17474,N_15433,N_14299);
or U17475 (N_17475,N_14102,N_15271);
nor U17476 (N_17476,N_14407,N_15265);
or U17477 (N_17477,N_15202,N_15402);
or U17478 (N_17478,N_14289,N_15316);
and U17479 (N_17479,N_14815,N_14450);
or U17480 (N_17480,N_14004,N_14190);
nor U17481 (N_17481,N_14682,N_14654);
and U17482 (N_17482,N_15871,N_14560);
or U17483 (N_17483,N_14939,N_15197);
nor U17484 (N_17484,N_15754,N_14272);
nor U17485 (N_17485,N_14901,N_15828);
xnor U17486 (N_17486,N_15452,N_14119);
nand U17487 (N_17487,N_15556,N_14819);
nor U17488 (N_17488,N_14802,N_14553);
nor U17489 (N_17489,N_14624,N_15521);
xor U17490 (N_17490,N_15694,N_15199);
nor U17491 (N_17491,N_14518,N_14965);
nor U17492 (N_17492,N_14067,N_14160);
nand U17493 (N_17493,N_14848,N_15266);
nand U17494 (N_17494,N_15984,N_14189);
and U17495 (N_17495,N_15573,N_15040);
or U17496 (N_17496,N_15250,N_14670);
nand U17497 (N_17497,N_15161,N_14978);
and U17498 (N_17498,N_14649,N_14539);
nand U17499 (N_17499,N_15304,N_14978);
nor U17500 (N_17500,N_15068,N_14571);
nor U17501 (N_17501,N_14814,N_15681);
and U17502 (N_17502,N_14720,N_15015);
and U17503 (N_17503,N_14720,N_14677);
nand U17504 (N_17504,N_15958,N_14058);
or U17505 (N_17505,N_15848,N_14566);
nand U17506 (N_17506,N_14208,N_14661);
nor U17507 (N_17507,N_14358,N_14566);
or U17508 (N_17508,N_15053,N_15987);
or U17509 (N_17509,N_14109,N_15756);
and U17510 (N_17510,N_15680,N_15724);
nand U17511 (N_17511,N_14348,N_15346);
nor U17512 (N_17512,N_14031,N_14823);
and U17513 (N_17513,N_15392,N_14233);
nor U17514 (N_17514,N_15908,N_15519);
nand U17515 (N_17515,N_14316,N_15513);
and U17516 (N_17516,N_15725,N_14350);
nor U17517 (N_17517,N_15933,N_14251);
or U17518 (N_17518,N_15457,N_15723);
nor U17519 (N_17519,N_14443,N_14155);
or U17520 (N_17520,N_14594,N_14242);
nor U17521 (N_17521,N_15870,N_15477);
nor U17522 (N_17522,N_15666,N_14702);
nand U17523 (N_17523,N_14144,N_14422);
or U17524 (N_17524,N_15092,N_15205);
nor U17525 (N_17525,N_14390,N_15139);
or U17526 (N_17526,N_15263,N_15619);
nor U17527 (N_17527,N_14619,N_14859);
or U17528 (N_17528,N_15168,N_15470);
nand U17529 (N_17529,N_15403,N_14516);
xnor U17530 (N_17530,N_14206,N_15508);
nor U17531 (N_17531,N_14958,N_15470);
nand U17532 (N_17532,N_14754,N_14845);
and U17533 (N_17533,N_15295,N_14283);
nand U17534 (N_17534,N_14301,N_14749);
or U17535 (N_17535,N_15027,N_14470);
and U17536 (N_17536,N_14723,N_15888);
xor U17537 (N_17537,N_15154,N_15582);
and U17538 (N_17538,N_14137,N_15222);
xor U17539 (N_17539,N_15744,N_15613);
or U17540 (N_17540,N_15004,N_14155);
or U17541 (N_17541,N_15400,N_15628);
xnor U17542 (N_17542,N_14007,N_14412);
nand U17543 (N_17543,N_14323,N_15845);
nand U17544 (N_17544,N_14349,N_15022);
and U17545 (N_17545,N_14258,N_15311);
or U17546 (N_17546,N_14097,N_15646);
and U17547 (N_17547,N_15448,N_15874);
or U17548 (N_17548,N_14186,N_15133);
or U17549 (N_17549,N_14759,N_15136);
nor U17550 (N_17550,N_14637,N_14398);
nand U17551 (N_17551,N_15994,N_15870);
nor U17552 (N_17552,N_14535,N_14902);
and U17553 (N_17553,N_14548,N_15216);
and U17554 (N_17554,N_14340,N_15816);
nor U17555 (N_17555,N_15048,N_14742);
and U17556 (N_17556,N_15394,N_14113);
nand U17557 (N_17557,N_15285,N_15221);
or U17558 (N_17558,N_14266,N_14700);
nor U17559 (N_17559,N_14056,N_15979);
and U17560 (N_17560,N_15163,N_15386);
and U17561 (N_17561,N_15686,N_15905);
nor U17562 (N_17562,N_14219,N_14217);
xnor U17563 (N_17563,N_15551,N_15111);
and U17564 (N_17564,N_14063,N_15192);
or U17565 (N_17565,N_14247,N_14215);
and U17566 (N_17566,N_14437,N_14466);
xor U17567 (N_17567,N_15865,N_15903);
and U17568 (N_17568,N_14379,N_15200);
nand U17569 (N_17569,N_15372,N_15963);
nor U17570 (N_17570,N_14360,N_15797);
and U17571 (N_17571,N_14760,N_15407);
and U17572 (N_17572,N_14518,N_14157);
or U17573 (N_17573,N_15713,N_14534);
nand U17574 (N_17574,N_14394,N_14866);
and U17575 (N_17575,N_15159,N_15587);
nand U17576 (N_17576,N_15715,N_15036);
and U17577 (N_17577,N_15965,N_15300);
nor U17578 (N_17578,N_14856,N_15062);
nand U17579 (N_17579,N_15491,N_14806);
or U17580 (N_17580,N_15981,N_14656);
and U17581 (N_17581,N_15955,N_15197);
nand U17582 (N_17582,N_14471,N_15601);
nand U17583 (N_17583,N_14770,N_15696);
and U17584 (N_17584,N_14777,N_15472);
nand U17585 (N_17585,N_15426,N_14322);
nor U17586 (N_17586,N_15606,N_14024);
nand U17587 (N_17587,N_15936,N_15937);
nor U17588 (N_17588,N_14743,N_14321);
and U17589 (N_17589,N_14312,N_14917);
nand U17590 (N_17590,N_14601,N_15621);
or U17591 (N_17591,N_15313,N_14977);
or U17592 (N_17592,N_15134,N_15111);
and U17593 (N_17593,N_15815,N_15603);
nand U17594 (N_17594,N_14013,N_15612);
or U17595 (N_17595,N_15186,N_15980);
nand U17596 (N_17596,N_15213,N_15247);
or U17597 (N_17597,N_15620,N_15667);
nand U17598 (N_17598,N_14544,N_14003);
nand U17599 (N_17599,N_15479,N_15122);
or U17600 (N_17600,N_15128,N_15526);
nor U17601 (N_17601,N_14246,N_15720);
nand U17602 (N_17602,N_14559,N_14998);
nor U17603 (N_17603,N_14436,N_15631);
or U17604 (N_17604,N_14797,N_15345);
nand U17605 (N_17605,N_15471,N_14692);
and U17606 (N_17606,N_14598,N_14909);
nand U17607 (N_17607,N_15525,N_15023);
nor U17608 (N_17608,N_14981,N_15943);
nand U17609 (N_17609,N_15961,N_14040);
and U17610 (N_17610,N_15977,N_14492);
nand U17611 (N_17611,N_14523,N_15751);
and U17612 (N_17612,N_14123,N_15608);
nor U17613 (N_17613,N_14499,N_15593);
or U17614 (N_17614,N_14522,N_15679);
or U17615 (N_17615,N_14651,N_14693);
and U17616 (N_17616,N_14237,N_14216);
and U17617 (N_17617,N_14177,N_15468);
xnor U17618 (N_17618,N_14628,N_14845);
xor U17619 (N_17619,N_15482,N_15942);
and U17620 (N_17620,N_15264,N_15895);
nor U17621 (N_17621,N_15319,N_15563);
nand U17622 (N_17622,N_15092,N_15447);
nor U17623 (N_17623,N_15569,N_15952);
and U17624 (N_17624,N_14620,N_14303);
or U17625 (N_17625,N_15902,N_14730);
nor U17626 (N_17626,N_15488,N_15343);
and U17627 (N_17627,N_15327,N_14491);
nor U17628 (N_17628,N_14769,N_14000);
and U17629 (N_17629,N_14417,N_15385);
nand U17630 (N_17630,N_14653,N_14222);
nand U17631 (N_17631,N_15638,N_14199);
or U17632 (N_17632,N_15238,N_15554);
nor U17633 (N_17633,N_15392,N_14053);
xnor U17634 (N_17634,N_14150,N_15054);
and U17635 (N_17635,N_15725,N_14265);
or U17636 (N_17636,N_15108,N_15234);
and U17637 (N_17637,N_14540,N_14547);
nor U17638 (N_17638,N_14211,N_14839);
nor U17639 (N_17639,N_14645,N_15679);
or U17640 (N_17640,N_15833,N_15671);
nand U17641 (N_17641,N_15834,N_14721);
or U17642 (N_17642,N_14637,N_15350);
xor U17643 (N_17643,N_14956,N_15808);
or U17644 (N_17644,N_14248,N_14043);
nor U17645 (N_17645,N_15738,N_14392);
nand U17646 (N_17646,N_15371,N_14358);
or U17647 (N_17647,N_14664,N_14476);
nand U17648 (N_17648,N_14486,N_15899);
nand U17649 (N_17649,N_14793,N_15064);
nand U17650 (N_17650,N_15571,N_15594);
or U17651 (N_17651,N_15445,N_15621);
and U17652 (N_17652,N_14974,N_15607);
xor U17653 (N_17653,N_15573,N_15847);
or U17654 (N_17654,N_14275,N_15057);
nor U17655 (N_17655,N_14127,N_15566);
nand U17656 (N_17656,N_15572,N_15468);
nor U17657 (N_17657,N_15396,N_15119);
or U17658 (N_17658,N_14702,N_15766);
or U17659 (N_17659,N_15062,N_14483);
nand U17660 (N_17660,N_15275,N_15970);
nor U17661 (N_17661,N_14813,N_15590);
xor U17662 (N_17662,N_14842,N_15465);
or U17663 (N_17663,N_15031,N_14836);
xor U17664 (N_17664,N_14421,N_15128);
and U17665 (N_17665,N_15775,N_15741);
nor U17666 (N_17666,N_14959,N_15703);
nor U17667 (N_17667,N_14472,N_15413);
nor U17668 (N_17668,N_15628,N_15073);
nor U17669 (N_17669,N_14261,N_14606);
nor U17670 (N_17670,N_14105,N_15817);
or U17671 (N_17671,N_15831,N_14774);
and U17672 (N_17672,N_14192,N_14098);
nand U17673 (N_17673,N_14744,N_14006);
xnor U17674 (N_17674,N_15281,N_14496);
nand U17675 (N_17675,N_14960,N_15188);
and U17676 (N_17676,N_15668,N_14750);
nor U17677 (N_17677,N_15787,N_14085);
nor U17678 (N_17678,N_15757,N_14164);
nand U17679 (N_17679,N_14916,N_14238);
nand U17680 (N_17680,N_14482,N_15210);
nor U17681 (N_17681,N_15677,N_14632);
nand U17682 (N_17682,N_15024,N_15052);
nor U17683 (N_17683,N_15006,N_14550);
or U17684 (N_17684,N_15110,N_15152);
or U17685 (N_17685,N_14681,N_15479);
nand U17686 (N_17686,N_15538,N_14097);
and U17687 (N_17687,N_15559,N_15289);
and U17688 (N_17688,N_14951,N_15546);
and U17689 (N_17689,N_14450,N_14941);
or U17690 (N_17690,N_15377,N_15891);
or U17691 (N_17691,N_14856,N_14834);
or U17692 (N_17692,N_15220,N_14531);
and U17693 (N_17693,N_15847,N_15649);
nor U17694 (N_17694,N_14971,N_14933);
nand U17695 (N_17695,N_15541,N_15587);
and U17696 (N_17696,N_14963,N_15518);
xnor U17697 (N_17697,N_14915,N_15754);
nand U17698 (N_17698,N_15255,N_15055);
and U17699 (N_17699,N_15284,N_15030);
or U17700 (N_17700,N_15544,N_15214);
or U17701 (N_17701,N_15176,N_15435);
and U17702 (N_17702,N_14266,N_15023);
nor U17703 (N_17703,N_15715,N_14201);
nor U17704 (N_17704,N_15255,N_14480);
xnor U17705 (N_17705,N_15920,N_15020);
nor U17706 (N_17706,N_14280,N_14187);
nand U17707 (N_17707,N_14989,N_14704);
nor U17708 (N_17708,N_15025,N_15113);
nor U17709 (N_17709,N_14019,N_14358);
and U17710 (N_17710,N_15734,N_15707);
or U17711 (N_17711,N_15130,N_15001);
nor U17712 (N_17712,N_15310,N_15453);
xnor U17713 (N_17713,N_15975,N_14209);
nor U17714 (N_17714,N_15275,N_14521);
nand U17715 (N_17715,N_15697,N_15653);
nor U17716 (N_17716,N_15987,N_14312);
or U17717 (N_17717,N_15378,N_15387);
nor U17718 (N_17718,N_14845,N_15633);
nor U17719 (N_17719,N_15603,N_15897);
or U17720 (N_17720,N_14794,N_14027);
or U17721 (N_17721,N_14396,N_14495);
nor U17722 (N_17722,N_15079,N_15228);
nand U17723 (N_17723,N_15631,N_14297);
nand U17724 (N_17724,N_14729,N_14856);
or U17725 (N_17725,N_14865,N_14717);
or U17726 (N_17726,N_14362,N_15303);
and U17727 (N_17727,N_14296,N_15229);
xor U17728 (N_17728,N_15552,N_14964);
and U17729 (N_17729,N_15812,N_14209);
and U17730 (N_17730,N_14198,N_14638);
nor U17731 (N_17731,N_14837,N_15572);
and U17732 (N_17732,N_15465,N_15214);
nor U17733 (N_17733,N_15707,N_15990);
or U17734 (N_17734,N_14928,N_15870);
and U17735 (N_17735,N_14427,N_14792);
nor U17736 (N_17736,N_14006,N_15063);
and U17737 (N_17737,N_14074,N_14680);
and U17738 (N_17738,N_15427,N_15079);
nand U17739 (N_17739,N_15008,N_15947);
and U17740 (N_17740,N_14562,N_14970);
and U17741 (N_17741,N_14760,N_15524);
or U17742 (N_17742,N_14386,N_14341);
nand U17743 (N_17743,N_15925,N_14965);
and U17744 (N_17744,N_15488,N_15417);
or U17745 (N_17745,N_15554,N_15305);
xor U17746 (N_17746,N_15004,N_14027);
nand U17747 (N_17747,N_14032,N_14310);
or U17748 (N_17748,N_14044,N_14299);
or U17749 (N_17749,N_15186,N_15624);
or U17750 (N_17750,N_15059,N_14368);
nand U17751 (N_17751,N_14177,N_14471);
nand U17752 (N_17752,N_15166,N_15325);
and U17753 (N_17753,N_15375,N_15233);
xor U17754 (N_17754,N_14880,N_14031);
xnor U17755 (N_17755,N_14637,N_14891);
nand U17756 (N_17756,N_15200,N_14601);
and U17757 (N_17757,N_14802,N_15981);
or U17758 (N_17758,N_14973,N_15022);
nand U17759 (N_17759,N_14594,N_14225);
nand U17760 (N_17760,N_15712,N_14290);
nor U17761 (N_17761,N_15095,N_15108);
nand U17762 (N_17762,N_14508,N_14398);
xor U17763 (N_17763,N_14597,N_14118);
or U17764 (N_17764,N_14229,N_14936);
or U17765 (N_17765,N_14033,N_15253);
and U17766 (N_17766,N_14103,N_14838);
or U17767 (N_17767,N_14973,N_15907);
and U17768 (N_17768,N_14761,N_15578);
and U17769 (N_17769,N_15774,N_15795);
nand U17770 (N_17770,N_14461,N_14276);
and U17771 (N_17771,N_15737,N_14965);
and U17772 (N_17772,N_15480,N_14074);
and U17773 (N_17773,N_14484,N_15407);
and U17774 (N_17774,N_14574,N_15487);
nor U17775 (N_17775,N_15366,N_15882);
or U17776 (N_17776,N_15261,N_15456);
xnor U17777 (N_17777,N_14944,N_15470);
and U17778 (N_17778,N_15248,N_14546);
xnor U17779 (N_17779,N_14944,N_15752);
nor U17780 (N_17780,N_15618,N_15836);
nand U17781 (N_17781,N_14546,N_14816);
nor U17782 (N_17782,N_14870,N_14793);
nor U17783 (N_17783,N_14986,N_15625);
or U17784 (N_17784,N_15484,N_15547);
or U17785 (N_17785,N_15762,N_15764);
nor U17786 (N_17786,N_15104,N_14433);
nor U17787 (N_17787,N_14610,N_14528);
and U17788 (N_17788,N_15135,N_15764);
nor U17789 (N_17789,N_15970,N_15483);
or U17790 (N_17790,N_15183,N_14817);
nor U17791 (N_17791,N_14448,N_15350);
or U17792 (N_17792,N_14882,N_15484);
nor U17793 (N_17793,N_15703,N_15579);
nor U17794 (N_17794,N_15278,N_14229);
nor U17795 (N_17795,N_14246,N_15275);
nor U17796 (N_17796,N_14641,N_15647);
and U17797 (N_17797,N_15887,N_15830);
nor U17798 (N_17798,N_15565,N_15994);
and U17799 (N_17799,N_15730,N_15440);
nor U17800 (N_17800,N_15957,N_14988);
and U17801 (N_17801,N_15456,N_15957);
and U17802 (N_17802,N_15683,N_15850);
or U17803 (N_17803,N_15504,N_15138);
and U17804 (N_17804,N_14651,N_14527);
or U17805 (N_17805,N_15533,N_15663);
nand U17806 (N_17806,N_14788,N_14593);
nand U17807 (N_17807,N_15524,N_15233);
or U17808 (N_17808,N_15549,N_15030);
nor U17809 (N_17809,N_15458,N_15374);
nor U17810 (N_17810,N_14577,N_14286);
and U17811 (N_17811,N_14515,N_15343);
nor U17812 (N_17812,N_15025,N_14580);
or U17813 (N_17813,N_15327,N_14473);
or U17814 (N_17814,N_14088,N_14127);
nand U17815 (N_17815,N_14550,N_14595);
nor U17816 (N_17816,N_15901,N_14840);
nand U17817 (N_17817,N_15854,N_15463);
nor U17818 (N_17818,N_14049,N_15467);
or U17819 (N_17819,N_14555,N_15660);
xor U17820 (N_17820,N_14920,N_15628);
nand U17821 (N_17821,N_14748,N_15460);
nor U17822 (N_17822,N_15111,N_15044);
nand U17823 (N_17823,N_15367,N_15916);
nand U17824 (N_17824,N_14157,N_14387);
xnor U17825 (N_17825,N_15956,N_14312);
nor U17826 (N_17826,N_15373,N_15991);
or U17827 (N_17827,N_15273,N_15138);
nand U17828 (N_17828,N_15168,N_14550);
and U17829 (N_17829,N_14065,N_14705);
and U17830 (N_17830,N_15289,N_14083);
nor U17831 (N_17831,N_14786,N_14976);
or U17832 (N_17832,N_14312,N_14818);
nor U17833 (N_17833,N_14995,N_15489);
and U17834 (N_17834,N_15703,N_15528);
nor U17835 (N_17835,N_14974,N_14549);
or U17836 (N_17836,N_15366,N_15472);
or U17837 (N_17837,N_15656,N_14907);
or U17838 (N_17838,N_14723,N_15591);
or U17839 (N_17839,N_14778,N_15666);
nor U17840 (N_17840,N_15496,N_14758);
nand U17841 (N_17841,N_14804,N_14649);
and U17842 (N_17842,N_15034,N_15403);
and U17843 (N_17843,N_14125,N_14615);
or U17844 (N_17844,N_15812,N_15033);
or U17845 (N_17845,N_15746,N_14042);
xnor U17846 (N_17846,N_14393,N_15430);
or U17847 (N_17847,N_15799,N_14830);
xor U17848 (N_17848,N_15394,N_14573);
or U17849 (N_17849,N_15026,N_15955);
and U17850 (N_17850,N_14484,N_14004);
or U17851 (N_17851,N_14354,N_14071);
and U17852 (N_17852,N_14883,N_15877);
nor U17853 (N_17853,N_14389,N_15426);
nor U17854 (N_17854,N_15603,N_14279);
or U17855 (N_17855,N_15632,N_15890);
or U17856 (N_17856,N_14589,N_15870);
nand U17857 (N_17857,N_14639,N_15344);
nand U17858 (N_17858,N_14396,N_15671);
and U17859 (N_17859,N_14383,N_15471);
nand U17860 (N_17860,N_14589,N_14361);
or U17861 (N_17861,N_14665,N_14700);
nor U17862 (N_17862,N_15769,N_15868);
or U17863 (N_17863,N_14771,N_14192);
nor U17864 (N_17864,N_14592,N_14670);
or U17865 (N_17865,N_15055,N_15169);
and U17866 (N_17866,N_14681,N_14950);
or U17867 (N_17867,N_15638,N_15407);
nand U17868 (N_17868,N_15904,N_14423);
xor U17869 (N_17869,N_14072,N_14342);
and U17870 (N_17870,N_15614,N_15225);
and U17871 (N_17871,N_14700,N_15521);
nor U17872 (N_17872,N_14960,N_15337);
or U17873 (N_17873,N_14576,N_14102);
nand U17874 (N_17874,N_15545,N_14035);
xnor U17875 (N_17875,N_15165,N_15418);
and U17876 (N_17876,N_15437,N_14939);
nand U17877 (N_17877,N_14535,N_15839);
nand U17878 (N_17878,N_14665,N_15501);
nor U17879 (N_17879,N_15719,N_15414);
xnor U17880 (N_17880,N_15873,N_14218);
or U17881 (N_17881,N_14406,N_14971);
nand U17882 (N_17882,N_15135,N_14465);
and U17883 (N_17883,N_14402,N_14258);
and U17884 (N_17884,N_15696,N_15485);
nand U17885 (N_17885,N_15437,N_14965);
nor U17886 (N_17886,N_14790,N_14860);
or U17887 (N_17887,N_15117,N_14319);
and U17888 (N_17888,N_15958,N_15906);
nor U17889 (N_17889,N_15375,N_14203);
or U17890 (N_17890,N_14979,N_15823);
or U17891 (N_17891,N_14529,N_14771);
nor U17892 (N_17892,N_14323,N_15208);
and U17893 (N_17893,N_15036,N_14027);
nand U17894 (N_17894,N_14164,N_14613);
and U17895 (N_17895,N_15289,N_14498);
or U17896 (N_17896,N_15502,N_14224);
nor U17897 (N_17897,N_15444,N_14148);
nor U17898 (N_17898,N_14196,N_14660);
nor U17899 (N_17899,N_15478,N_14117);
and U17900 (N_17900,N_15293,N_14277);
nand U17901 (N_17901,N_14394,N_15219);
nor U17902 (N_17902,N_14880,N_14025);
or U17903 (N_17903,N_14185,N_14257);
nand U17904 (N_17904,N_15408,N_15155);
or U17905 (N_17905,N_15539,N_14987);
and U17906 (N_17906,N_15202,N_15797);
and U17907 (N_17907,N_14794,N_15904);
or U17908 (N_17908,N_15485,N_15204);
nand U17909 (N_17909,N_15294,N_15848);
xnor U17910 (N_17910,N_14727,N_15403);
and U17911 (N_17911,N_14585,N_14210);
xnor U17912 (N_17912,N_15050,N_15371);
nor U17913 (N_17913,N_14825,N_15470);
or U17914 (N_17914,N_15832,N_14587);
and U17915 (N_17915,N_14898,N_15964);
and U17916 (N_17916,N_15398,N_15336);
or U17917 (N_17917,N_15069,N_15647);
xor U17918 (N_17918,N_14574,N_15509);
nand U17919 (N_17919,N_14498,N_15682);
nor U17920 (N_17920,N_15596,N_15578);
nand U17921 (N_17921,N_15245,N_15439);
xor U17922 (N_17922,N_15265,N_14738);
nor U17923 (N_17923,N_15013,N_15471);
xnor U17924 (N_17924,N_14470,N_15015);
nor U17925 (N_17925,N_15197,N_14901);
or U17926 (N_17926,N_14045,N_14303);
or U17927 (N_17927,N_15163,N_14664);
or U17928 (N_17928,N_15860,N_15339);
xnor U17929 (N_17929,N_14878,N_14908);
and U17930 (N_17930,N_14703,N_14878);
and U17931 (N_17931,N_15568,N_14992);
or U17932 (N_17932,N_15034,N_14331);
nand U17933 (N_17933,N_15046,N_15849);
or U17934 (N_17934,N_15498,N_14416);
nor U17935 (N_17935,N_14059,N_14075);
and U17936 (N_17936,N_14749,N_15809);
nand U17937 (N_17937,N_14315,N_14267);
or U17938 (N_17938,N_15642,N_14783);
and U17939 (N_17939,N_14978,N_14253);
and U17940 (N_17940,N_15851,N_15425);
or U17941 (N_17941,N_14321,N_15259);
or U17942 (N_17942,N_15336,N_15180);
or U17943 (N_17943,N_15322,N_14388);
and U17944 (N_17944,N_15725,N_14523);
nor U17945 (N_17945,N_15779,N_15579);
nor U17946 (N_17946,N_14156,N_15879);
or U17947 (N_17947,N_14507,N_15485);
nor U17948 (N_17948,N_14772,N_14310);
or U17949 (N_17949,N_15188,N_14228);
nand U17950 (N_17950,N_15427,N_15476);
or U17951 (N_17951,N_14178,N_14700);
xor U17952 (N_17952,N_14422,N_15145);
nor U17953 (N_17953,N_14188,N_15988);
or U17954 (N_17954,N_15874,N_15502);
xnor U17955 (N_17955,N_14448,N_14006);
nor U17956 (N_17956,N_15387,N_15011);
and U17957 (N_17957,N_14884,N_15475);
nor U17958 (N_17958,N_15275,N_14594);
nor U17959 (N_17959,N_14921,N_15132);
and U17960 (N_17960,N_15104,N_15897);
or U17961 (N_17961,N_15752,N_15602);
and U17962 (N_17962,N_14008,N_15216);
or U17963 (N_17963,N_15665,N_14542);
xor U17964 (N_17964,N_15078,N_15224);
and U17965 (N_17965,N_14624,N_14495);
nand U17966 (N_17966,N_14432,N_14775);
nand U17967 (N_17967,N_15182,N_15099);
nand U17968 (N_17968,N_14556,N_14242);
nand U17969 (N_17969,N_14119,N_15842);
nor U17970 (N_17970,N_14108,N_15388);
nand U17971 (N_17971,N_14667,N_14697);
nand U17972 (N_17972,N_14717,N_15080);
nor U17973 (N_17973,N_14352,N_15711);
and U17974 (N_17974,N_14420,N_14717);
xor U17975 (N_17975,N_14841,N_15465);
and U17976 (N_17976,N_15823,N_15288);
or U17977 (N_17977,N_14122,N_15687);
and U17978 (N_17978,N_14016,N_15280);
nor U17979 (N_17979,N_15730,N_14426);
and U17980 (N_17980,N_15631,N_14074);
or U17981 (N_17981,N_14273,N_15579);
xor U17982 (N_17982,N_15730,N_14043);
or U17983 (N_17983,N_15747,N_14533);
xor U17984 (N_17984,N_15221,N_14333);
and U17985 (N_17985,N_14377,N_14900);
nor U17986 (N_17986,N_15958,N_14411);
nand U17987 (N_17987,N_15123,N_14495);
and U17988 (N_17988,N_15019,N_15874);
nor U17989 (N_17989,N_14008,N_14652);
nor U17990 (N_17990,N_15725,N_15286);
xnor U17991 (N_17991,N_14587,N_15224);
and U17992 (N_17992,N_15250,N_14823);
or U17993 (N_17993,N_15798,N_15328);
nand U17994 (N_17994,N_15385,N_15533);
and U17995 (N_17995,N_15818,N_15387);
nor U17996 (N_17996,N_15479,N_15118);
and U17997 (N_17997,N_14881,N_14147);
nand U17998 (N_17998,N_14415,N_14530);
xor U17999 (N_17999,N_14063,N_14203);
and U18000 (N_18000,N_16230,N_17938);
nor U18001 (N_18001,N_17769,N_17946);
nor U18002 (N_18002,N_17614,N_17015);
and U18003 (N_18003,N_16142,N_17825);
nor U18004 (N_18004,N_16840,N_16351);
or U18005 (N_18005,N_16410,N_17048);
nand U18006 (N_18006,N_16323,N_17371);
and U18007 (N_18007,N_17680,N_16588);
nor U18008 (N_18008,N_16949,N_16032);
and U18009 (N_18009,N_16655,N_17995);
nand U18010 (N_18010,N_16468,N_17489);
or U18011 (N_18011,N_16113,N_16549);
nand U18012 (N_18012,N_16589,N_16563);
or U18013 (N_18013,N_16418,N_16141);
nor U18014 (N_18014,N_17333,N_16612);
nor U18015 (N_18015,N_16764,N_17844);
nor U18016 (N_18016,N_17984,N_16704);
or U18017 (N_18017,N_16930,N_16147);
nor U18018 (N_18018,N_16438,N_17171);
nand U18019 (N_18019,N_16648,N_16683);
or U18020 (N_18020,N_17024,N_16297);
nand U18021 (N_18021,N_16682,N_17109);
nand U18022 (N_18022,N_17519,N_16278);
or U18023 (N_18023,N_16865,N_17941);
and U18024 (N_18024,N_16693,N_16432);
nor U18025 (N_18025,N_17804,N_17552);
or U18026 (N_18026,N_17923,N_16999);
or U18027 (N_18027,N_17916,N_16611);
nand U18028 (N_18028,N_16659,N_16478);
and U18029 (N_18029,N_17172,N_17367);
nand U18030 (N_18030,N_17113,N_17554);
nand U18031 (N_18031,N_17343,N_16644);
nand U18032 (N_18032,N_16606,N_17594);
nand U18033 (N_18033,N_17885,N_16863);
nand U18034 (N_18034,N_16150,N_17880);
nor U18035 (N_18035,N_17381,N_16448);
or U18036 (N_18036,N_17985,N_16143);
nor U18037 (N_18037,N_16969,N_17467);
and U18038 (N_18038,N_17005,N_16347);
or U18039 (N_18039,N_16381,N_16285);
xor U18040 (N_18040,N_16100,N_16484);
nand U18041 (N_18041,N_16650,N_17702);
nor U18042 (N_18042,N_16262,N_17002);
or U18043 (N_18043,N_17642,N_16112);
and U18044 (N_18044,N_16900,N_17476);
xnor U18045 (N_18045,N_16867,N_17562);
and U18046 (N_18046,N_16377,N_16986);
xnor U18047 (N_18047,N_16958,N_17021);
nor U18048 (N_18048,N_17484,N_16575);
nor U18049 (N_18049,N_17589,N_16360);
nor U18050 (N_18050,N_16171,N_17396);
nand U18051 (N_18051,N_17060,N_17188);
and U18052 (N_18052,N_16767,N_16678);
and U18053 (N_18053,N_17560,N_17913);
and U18054 (N_18054,N_16831,N_16107);
or U18055 (N_18055,N_16873,N_16316);
nor U18056 (N_18056,N_17225,N_16102);
nand U18057 (N_18057,N_17276,N_17287);
xor U18058 (N_18058,N_17696,N_16241);
or U18059 (N_18059,N_17265,N_16376);
or U18060 (N_18060,N_16572,N_16551);
and U18061 (N_18061,N_17622,N_17167);
nand U18062 (N_18062,N_17295,N_17737);
nor U18063 (N_18063,N_17008,N_16668);
nand U18064 (N_18064,N_17848,N_16548);
nand U18065 (N_18065,N_16200,N_16138);
or U18066 (N_18066,N_17464,N_17253);
and U18067 (N_18067,N_17184,N_17471);
nand U18068 (N_18068,N_16750,N_16491);
nor U18069 (N_18069,N_17847,N_16148);
nor U18070 (N_18070,N_17711,N_16294);
and U18071 (N_18071,N_16779,N_17776);
nand U18072 (N_18072,N_16918,N_17255);
and U18073 (N_18073,N_16281,N_16803);
xnor U18074 (N_18074,N_16737,N_16028);
or U18075 (N_18075,N_17348,N_16591);
xnor U18076 (N_18076,N_16385,N_16215);
nor U18077 (N_18077,N_17293,N_17139);
nand U18078 (N_18078,N_16774,N_16666);
or U18079 (N_18079,N_17423,N_16717);
nor U18080 (N_18080,N_16079,N_16495);
or U18081 (N_18081,N_17877,N_16783);
nand U18082 (N_18082,N_16406,N_17685);
nand U18083 (N_18083,N_17821,N_17179);
and U18084 (N_18084,N_16229,N_16136);
nand U18085 (N_18085,N_16832,N_17756);
and U18086 (N_18086,N_16736,N_17676);
nor U18087 (N_18087,N_17585,N_16159);
and U18088 (N_18088,N_17195,N_16508);
nand U18089 (N_18089,N_17173,N_16125);
nor U18090 (N_18090,N_16466,N_17502);
or U18091 (N_18091,N_17736,N_17338);
nand U18092 (N_18092,N_16210,N_16293);
nand U18093 (N_18093,N_16341,N_17105);
nand U18094 (N_18094,N_17742,N_17237);
and U18095 (N_18095,N_16637,N_17727);
nand U18096 (N_18096,N_17836,N_17949);
nor U18097 (N_18097,N_17865,N_17812);
or U18098 (N_18098,N_17539,N_17340);
or U18099 (N_18099,N_16092,N_17695);
and U18100 (N_18100,N_16409,N_17615);
xor U18101 (N_18101,N_16415,N_16841);
and U18102 (N_18102,N_16676,N_16905);
nand U18103 (N_18103,N_17267,N_16393);
nor U18104 (N_18104,N_17486,N_16835);
or U18105 (N_18105,N_16787,N_16025);
or U18106 (N_18106,N_16480,N_16698);
or U18107 (N_18107,N_16095,N_16621);
or U18108 (N_18108,N_16272,N_16234);
nand U18109 (N_18109,N_16027,N_17244);
nand U18110 (N_18110,N_16423,N_17904);
nand U18111 (N_18111,N_17196,N_17601);
or U18112 (N_18112,N_17254,N_17639);
nand U18113 (N_18113,N_17439,N_17477);
or U18114 (N_18114,N_17407,N_16592);
nor U18115 (N_18115,N_17270,N_16008);
nand U18116 (N_18116,N_17433,N_17337);
and U18117 (N_18117,N_17915,N_17029);
nor U18118 (N_18118,N_16651,N_16614);
and U18119 (N_18119,N_17741,N_17643);
xor U18120 (N_18120,N_16332,N_17954);
xor U18121 (N_18121,N_16538,N_17217);
or U18122 (N_18122,N_17548,N_16753);
nand U18123 (N_18123,N_16732,N_17799);
nand U18124 (N_18124,N_17198,N_16653);
or U18125 (N_18125,N_16977,N_17768);
nor U18126 (N_18126,N_17305,N_17070);
nor U18127 (N_18127,N_16400,N_17550);
and U18128 (N_18128,N_17996,N_17505);
or U18129 (N_18129,N_17272,N_16174);
or U18130 (N_18130,N_16980,N_17587);
or U18131 (N_18131,N_16191,N_16635);
nor U18132 (N_18132,N_17186,N_16935);
or U18133 (N_18133,N_16435,N_16688);
nor U18134 (N_18134,N_17876,N_17118);
nor U18135 (N_18135,N_16439,N_16273);
nor U18136 (N_18136,N_17025,N_17677);
or U18137 (N_18137,N_17827,N_17809);
nor U18138 (N_18138,N_16477,N_16228);
nand U18139 (N_18139,N_16392,N_16288);
nand U18140 (N_18140,N_17636,N_16103);
and U18141 (N_18141,N_16859,N_16854);
or U18142 (N_18142,N_17302,N_16946);
and U18143 (N_18143,N_16602,N_16601);
or U18144 (N_18144,N_17782,N_17602);
and U18145 (N_18145,N_16349,N_17992);
nand U18146 (N_18146,N_16872,N_17250);
nor U18147 (N_18147,N_17240,N_17482);
nor U18148 (N_18148,N_17811,N_17845);
xnor U18149 (N_18149,N_17864,N_16511);
xor U18150 (N_18150,N_16098,N_16353);
and U18151 (N_18151,N_17752,N_16401);
or U18152 (N_18152,N_16154,N_16494);
and U18153 (N_18153,N_16785,N_17950);
or U18154 (N_18154,N_16308,N_16450);
xnor U18155 (N_18155,N_17387,N_17147);
nand U18156 (N_18156,N_16836,N_16296);
or U18157 (N_18157,N_16616,N_17064);
nand U18158 (N_18158,N_16099,N_16012);
nor U18159 (N_18159,N_16673,N_17824);
and U18160 (N_18160,N_16366,N_17556);
xnor U18161 (N_18161,N_16885,N_17584);
and U18162 (N_18162,N_16679,N_17717);
or U18163 (N_18163,N_16249,N_16336);
or U18164 (N_18164,N_17249,N_17599);
nor U18165 (N_18165,N_16137,N_16071);
nand U18166 (N_18166,N_17134,N_16500);
and U18167 (N_18167,N_17124,N_17054);
and U18168 (N_18168,N_17859,N_16800);
xor U18169 (N_18169,N_17221,N_16735);
nor U18170 (N_18170,N_17947,N_17291);
and U18171 (N_18171,N_17185,N_17573);
nand U18172 (N_18172,N_17716,N_16761);
nor U18173 (N_18173,N_17391,N_17405);
xnor U18174 (N_18174,N_16738,N_17873);
nor U18175 (N_18175,N_17942,N_17389);
or U18176 (N_18176,N_17878,N_17434);
or U18177 (N_18177,N_16037,N_17213);
or U18178 (N_18178,N_16157,N_17088);
and U18179 (N_18179,N_16583,N_17849);
or U18180 (N_18180,N_17369,N_16305);
nand U18181 (N_18181,N_16260,N_16994);
and U18182 (N_18182,N_17259,N_17735);
nand U18183 (N_18183,N_17000,N_16163);
nor U18184 (N_18184,N_17819,N_16340);
nor U18185 (N_18185,N_17416,N_16839);
and U18186 (N_18186,N_17504,N_16057);
or U18187 (N_18187,N_17038,N_17073);
and U18188 (N_18188,N_16674,N_17428);
or U18189 (N_18189,N_16654,N_16536);
nand U18190 (N_18190,N_16164,N_16266);
or U18191 (N_18191,N_16675,N_16680);
nand U18192 (N_18192,N_16198,N_16667);
and U18193 (N_18193,N_16901,N_17500);
nand U18194 (N_18194,N_16145,N_17511);
and U18195 (N_18195,N_17801,N_16554);
and U18196 (N_18196,N_16017,N_17398);
nand U18197 (N_18197,N_17401,N_16408);
and U18198 (N_18198,N_16453,N_17781);
and U18199 (N_18199,N_17778,N_17708);
or U18200 (N_18200,N_16819,N_17612);
nand U18201 (N_18201,N_16757,N_17662);
nand U18202 (N_18202,N_17275,N_16561);
and U18203 (N_18203,N_17055,N_17532);
nor U18204 (N_18204,N_17432,N_16302);
nor U18205 (N_18205,N_16727,N_16007);
xor U18206 (N_18206,N_16492,N_17062);
or U18207 (N_18207,N_17830,N_16250);
or U18208 (N_18208,N_17582,N_17775);
nor U18209 (N_18209,N_17030,N_16503);
or U18210 (N_18210,N_17903,N_17951);
or U18211 (N_18211,N_16166,N_17354);
nand U18212 (N_18212,N_17637,N_16715);
or U18213 (N_18213,N_17375,N_16402);
nor U18214 (N_18214,N_16733,N_16327);
nor U18215 (N_18215,N_16627,N_17318);
nor U18216 (N_18216,N_16827,N_16289);
or U18217 (N_18217,N_16066,N_17980);
and U18218 (N_18218,N_17262,N_16259);
nand U18219 (N_18219,N_17478,N_17579);
xnor U18220 (N_18220,N_16421,N_16747);
nor U18221 (N_18221,N_17663,N_17260);
nand U18222 (N_18222,N_16797,N_17613);
nand U18223 (N_18223,N_17450,N_17943);
or U18224 (N_18224,N_16760,N_16178);
nor U18225 (N_18225,N_16989,N_16501);
or U18226 (N_18226,N_16093,N_17926);
nor U18227 (N_18227,N_17378,N_17852);
or U18228 (N_18228,N_17598,N_16237);
nand U18229 (N_18229,N_17521,N_16261);
nor U18230 (N_18230,N_16852,N_16874);
nor U18231 (N_18231,N_17967,N_17501);
and U18232 (N_18232,N_16485,N_17816);
xor U18233 (N_18233,N_17085,N_17133);
or U18234 (N_18234,N_17854,N_16313);
and U18235 (N_18235,N_17264,N_17686);
or U18236 (N_18236,N_17688,N_16721);
and U18237 (N_18237,N_17412,N_16463);
or U18238 (N_18238,N_17571,N_16245);
nor U18239 (N_18239,N_17493,N_16580);
xnor U18240 (N_18240,N_16033,N_17309);
nand U18241 (N_18241,N_17789,N_16844);
and U18242 (N_18242,N_17136,N_16906);
and U18243 (N_18243,N_16587,N_16371);
or U18244 (N_18244,N_17870,N_17409);
xnor U18245 (N_18245,N_16746,N_16405);
nand U18246 (N_18246,N_17491,N_17116);
or U18247 (N_18247,N_16603,N_16222);
and U18248 (N_18248,N_17581,N_17959);
nor U18249 (N_18249,N_17067,N_17568);
or U18250 (N_18250,N_16233,N_17119);
or U18251 (N_18251,N_17110,N_16047);
xor U18252 (N_18252,N_16074,N_16253);
or U18253 (N_18253,N_16447,N_17017);
and U18254 (N_18254,N_17473,N_17525);
nand U18255 (N_18255,N_16236,N_17235);
nor U18256 (N_18256,N_16975,N_17207);
nand U18257 (N_18257,N_17933,N_16365);
nor U18258 (N_18258,N_16443,N_16576);
and U18259 (N_18259,N_16306,N_16342);
nor U18260 (N_18260,N_17080,N_16567);
nand U18261 (N_18261,N_16355,N_17430);
nand U18262 (N_18262,N_16181,N_16828);
nand U18263 (N_18263,N_16629,N_17211);
and U18264 (N_18264,N_17961,N_16584);
and U18265 (N_18265,N_16581,N_17499);
and U18266 (N_18266,N_17414,N_16502);
nor U18267 (N_18267,N_17796,N_17014);
and U18268 (N_18268,N_17475,N_16891);
nor U18269 (N_18269,N_16525,N_16451);
or U18270 (N_18270,N_16642,N_17011);
nor U18271 (N_18271,N_16345,N_17436);
and U18272 (N_18272,N_17956,N_17049);
nor U18273 (N_18273,N_16346,N_17290);
nor U18274 (N_18274,N_16833,N_17991);
nor U18275 (N_18275,N_17284,N_17580);
nand U18276 (N_18276,N_17128,N_16045);
nor U18277 (N_18277,N_16597,N_17965);
or U18278 (N_18278,N_16252,N_17152);
xor U18279 (N_18279,N_16445,N_17953);
or U18280 (N_18280,N_16383,N_17181);
nor U18281 (N_18281,N_16813,N_16686);
or U18282 (N_18282,N_17150,N_17127);
and U18283 (N_18283,N_16195,N_17679);
nor U18284 (N_18284,N_17624,N_16647);
nor U18285 (N_18285,N_17729,N_16378);
nand U18286 (N_18286,N_17114,N_16938);
nor U18287 (N_18287,N_16015,N_16156);
or U18288 (N_18288,N_16035,N_16023);
xor U18289 (N_18289,N_17009,N_16943);
and U18290 (N_18290,N_16334,N_17115);
or U18291 (N_18291,N_17681,N_16789);
nand U18292 (N_18292,N_16490,N_16911);
nand U18293 (N_18293,N_17656,N_16209);
nand U18294 (N_18294,N_17631,N_16177);
or U18295 (N_18295,N_16806,N_16457);
nor U18296 (N_18296,N_16304,N_16907);
or U18297 (N_18297,N_17962,N_16090);
or U18298 (N_18298,N_16036,N_17772);
nand U18299 (N_18299,N_17555,N_16188);
and U18300 (N_18300,N_16579,N_16462);
nand U18301 (N_18301,N_17419,N_16546);
nor U18302 (N_18302,N_17061,N_17872);
nor U18303 (N_18303,N_17321,N_16981);
or U18304 (N_18304,N_16424,N_16689);
xnor U18305 (N_18305,N_16419,N_16772);
and U18306 (N_18306,N_17100,N_17749);
and U18307 (N_18307,N_16056,N_16104);
or U18308 (N_18308,N_17862,N_17590);
xnor U18309 (N_18309,N_16712,N_17395);
or U18310 (N_18310,N_16613,N_16399);
nor U18311 (N_18311,N_16170,N_16773);
xnor U18312 (N_18312,N_17047,N_16719);
and U18313 (N_18313,N_16184,N_16054);
and U18314 (N_18314,N_17835,N_17514);
or U18315 (N_18315,N_16769,N_16542);
nor U18316 (N_18316,N_16582,N_17480);
or U18317 (N_18317,N_16433,N_17528);
nand U18318 (N_18318,N_16126,N_16691);
nor U18319 (N_18319,N_17721,N_16111);
or U18320 (N_18320,N_16734,N_17111);
nor U18321 (N_18321,N_16444,N_17045);
and U18322 (N_18322,N_16837,N_16251);
or U18323 (N_18323,N_17292,N_17328);
nand U18324 (N_18324,N_16880,N_16173);
nand U18325 (N_18325,N_17059,N_17683);
nand U18326 (N_18326,N_16596,N_17924);
and U18327 (N_18327,N_17345,N_17699);
and U18328 (N_18328,N_17065,N_16489);
xnor U18329 (N_18329,N_16223,N_16776);
nor U18330 (N_18330,N_16566,N_17393);
and U18331 (N_18331,N_16373,N_17744);
nand U18332 (N_18332,N_16268,N_16775);
and U18333 (N_18333,N_16220,N_17731);
and U18334 (N_18334,N_17842,N_17588);
and U18335 (N_18335,N_16106,N_16310);
nor U18336 (N_18336,N_17754,N_16179);
nor U18337 (N_18337,N_16124,N_16531);
nand U18338 (N_18338,N_16553,N_16461);
or U18339 (N_18339,N_16050,N_17191);
and U18340 (N_18340,N_16205,N_17958);
nor U18341 (N_18341,N_16456,N_17549);
and U18342 (N_18342,N_16522,N_16625);
xnor U18343 (N_18343,N_17162,N_17868);
nor U18344 (N_18344,N_16506,N_17041);
and U18345 (N_18345,N_16329,N_16845);
and U18346 (N_18346,N_16314,N_17356);
or U18347 (N_18347,N_17529,N_17839);
nor U18348 (N_18348,N_17906,N_16758);
nor U18349 (N_18349,N_16826,N_16780);
and U18350 (N_18350,N_16458,N_17881);
nand U18351 (N_18351,N_17705,N_17875);
and U18352 (N_18352,N_17036,N_16876);
nand U18353 (N_18353,N_17765,N_17141);
or U18354 (N_18354,N_16232,N_16607);
or U18355 (N_18355,N_16105,N_17183);
and U18356 (N_18356,N_16076,N_17052);
nor U18357 (N_18357,N_16088,N_16893);
and U18358 (N_18358,N_17397,N_16487);
and U18359 (N_18359,N_16847,N_17204);
nor U18360 (N_18360,N_17784,N_17547);
nand U18361 (N_18361,N_16545,N_16641);
and U18362 (N_18362,N_16794,N_17763);
nor U18363 (N_18363,N_16869,N_16834);
and U18364 (N_18364,N_16799,N_16067);
nor U18365 (N_18365,N_16743,N_17077);
or U18366 (N_18366,N_16357,N_16632);
and U18367 (N_18367,N_17905,N_16527);
nor U18368 (N_18368,N_17296,N_17056);
and U18369 (N_18369,N_16442,N_16540);
nor U18370 (N_18370,N_17545,N_17071);
and U18371 (N_18371,N_17583,N_16896);
nand U18372 (N_18372,N_16291,N_16254);
or U18373 (N_18373,N_17972,N_16328);
xnor U18374 (N_18374,N_17818,N_16778);
nand U18375 (N_18375,N_16877,N_16537);
nand U18376 (N_18376,N_16481,N_17530);
nand U18377 (N_18377,N_17593,N_16963);
nor U18378 (N_18378,N_16870,N_17326);
nor U18379 (N_18379,N_16765,N_17233);
nor U18380 (N_18380,N_17146,N_16805);
nand U18381 (N_18381,N_16344,N_17750);
and U18382 (N_18382,N_16923,N_16019);
and U18383 (N_18383,N_16211,N_17299);
nor U18384 (N_18384,N_16031,N_16060);
and U18385 (N_18385,N_16941,N_16550);
nand U18386 (N_18386,N_17462,N_17066);
and U18387 (N_18387,N_16182,N_17570);
and U18388 (N_18388,N_16335,N_16729);
and U18389 (N_18389,N_17666,N_16269);
xor U18390 (N_18390,N_16745,N_16243);
or U18391 (N_18391,N_16802,N_16897);
nand U18392 (N_18392,N_17723,N_17828);
nand U18393 (N_18393,N_17882,N_17334);
nor U18394 (N_18394,N_17586,N_17997);
nor U18395 (N_18395,N_16922,N_17003);
nor U18396 (N_18396,N_16043,N_16333);
xor U18397 (N_18397,N_16299,N_17994);
and U18398 (N_18398,N_17851,N_16942);
and U18399 (N_18399,N_17447,N_17856);
nor U18400 (N_18400,N_16749,N_16437);
or U18401 (N_18401,N_17352,N_17960);
nand U18402 (N_18402,N_16082,N_16725);
or U18403 (N_18403,N_17704,N_17018);
nand U18404 (N_18404,N_16115,N_16343);
xor U18405 (N_18405,N_16473,N_17630);
or U18406 (N_18406,N_16264,N_17086);
or U18407 (N_18407,N_17617,N_16982);
or U18408 (N_18408,N_17918,N_17155);
and U18409 (N_18409,N_17046,N_17470);
nor U18410 (N_18410,N_17385,N_16726);
or U18411 (N_18411,N_17945,N_16798);
or U18412 (N_18412,N_16882,N_17382);
xor U18413 (N_18413,N_17129,N_17667);
or U18414 (N_18414,N_16878,N_17982);
nand U18415 (N_18415,N_17700,N_17939);
nor U18416 (N_18416,N_16338,N_17983);
xnor U18417 (N_18417,N_16752,N_16889);
or U18418 (N_18418,N_17928,N_17001);
nand U18419 (N_18419,N_16920,N_17031);
nor U18420 (N_18420,N_16227,N_17888);
and U18421 (N_18421,N_16059,N_17883);
and U18422 (N_18422,N_17420,N_17379);
nor U18423 (N_18423,N_17725,N_16731);
xnor U18424 (N_18424,N_16646,N_16562);
or U18425 (N_18425,N_16441,N_17764);
nand U18426 (N_18426,N_17898,N_17900);
nand U18427 (N_18427,N_16777,N_17513);
or U18428 (N_18428,N_16853,N_17576);
or U18429 (N_18429,N_17930,N_16356);
nor U18430 (N_18430,N_16690,N_17037);
nand U18431 (N_18431,N_17357,N_17206);
nor U18432 (N_18432,N_16397,N_17438);
and U18433 (N_18433,N_16792,N_17542);
nor U18434 (N_18434,N_16620,N_16068);
or U18435 (N_18435,N_17595,N_16394);
nand U18436 (N_18436,N_16003,N_17411);
nand U18437 (N_18437,N_17329,N_17652);
xor U18438 (N_18438,N_17222,N_16534);
or U18439 (N_18439,N_16464,N_16883);
nand U18440 (N_18440,N_17189,N_17361);
and U18441 (N_18441,N_17874,N_16149);
nand U18442 (N_18442,N_17494,N_16011);
nand U18443 (N_18443,N_17834,N_16022);
and U18444 (N_18444,N_16710,N_17279);
or U18445 (N_18445,N_17914,N_17449);
or U18446 (N_18446,N_17618,N_16671);
xor U18447 (N_18447,N_17032,N_16959);
nand U18448 (N_18448,N_17330,N_17761);
or U18449 (N_18449,N_17665,N_17553);
nand U18450 (N_18450,N_16702,N_16073);
nor U18451 (N_18451,N_16657,N_17692);
nand U18452 (N_18452,N_16324,N_17429);
nor U18453 (N_18453,N_16153,N_17368);
and U18454 (N_18454,N_16339,N_16699);
or U18455 (N_18455,N_16816,N_16425);
nand U18456 (N_18456,N_16626,N_17831);
and U18457 (N_18457,N_17336,N_17485);
and U18458 (N_18458,N_16380,N_17090);
nor U18459 (N_18459,N_17694,N_16311);
nor U18460 (N_18460,N_17795,N_16244);
nand U18461 (N_18461,N_17650,N_17390);
or U18462 (N_18462,N_17981,N_17460);
and U18463 (N_18463,N_17523,N_17912);
nor U18464 (N_18464,N_17896,N_16984);
nor U18465 (N_18465,N_16993,N_16168);
or U18466 (N_18466,N_16005,N_17843);
and U18467 (N_18467,N_16312,N_16390);
xnor U18468 (N_18468,N_16034,N_16782);
nand U18469 (N_18469,N_16814,N_16129);
or U18470 (N_18470,N_16716,N_16565);
nand U18471 (N_18471,N_17280,N_16135);
xor U18472 (N_18472,N_17151,N_17413);
nand U18473 (N_18473,N_16564,N_16714);
nand U18474 (N_18474,N_16224,N_17869);
nor U18475 (N_18475,N_17281,N_16978);
nand U18476 (N_18476,N_17771,N_17163);
nand U18477 (N_18477,N_16422,N_17948);
and U18478 (N_18478,N_17793,N_17016);
and U18479 (N_18479,N_16917,N_16430);
or U18480 (N_18480,N_17807,N_17963);
nand U18481 (N_18481,N_17194,N_17245);
nand U18482 (N_18482,N_17861,N_16483);
or U18483 (N_18483,N_17452,N_17803);
or U18484 (N_18484,N_17312,N_16768);
and U18485 (N_18485,N_16957,N_17786);
and U18486 (N_18486,N_17040,N_16002);
nor U18487 (N_18487,N_16072,N_17712);
nor U18488 (N_18488,N_17425,N_16670);
nor U18489 (N_18489,N_16242,N_16434);
and U18490 (N_18490,N_16204,N_17023);
nor U18491 (N_18491,N_16751,N_16910);
and U18492 (N_18492,N_17574,N_16979);
and U18493 (N_18493,N_17437,N_17376);
xor U18494 (N_18494,N_16513,N_16722);
nand U18495 (N_18495,N_16295,N_17012);
nor U18496 (N_18496,N_17575,N_16578);
and U18497 (N_18497,N_17838,N_17664);
or U18498 (N_18498,N_17748,N_17937);
or U18499 (N_18499,N_16026,N_17657);
or U18500 (N_18500,N_16207,N_16953);
nand U18501 (N_18501,N_17977,N_17687);
xor U18502 (N_18502,N_17899,N_16014);
or U18503 (N_18503,N_17158,N_16991);
xnor U18504 (N_18504,N_16412,N_16146);
nand U18505 (N_18505,N_17603,N_16039);
nor U18506 (N_18506,N_16042,N_16524);
nand U18507 (N_18507,N_16199,N_17506);
nand U18508 (N_18508,N_17286,N_16172);
and U18509 (N_18509,N_16348,N_17964);
nor U18510 (N_18510,N_16130,N_17408);
nor U18511 (N_18511,N_16382,N_16284);
and U18512 (N_18512,N_16208,N_17201);
or U18513 (N_18513,N_16809,N_17509);
nor U18514 (N_18514,N_16552,N_16465);
or U18515 (N_18515,N_16692,N_17282);
and U18516 (N_18516,N_16155,N_17440);
and U18517 (N_18517,N_16730,N_17907);
or U18518 (N_18518,N_17344,N_17074);
nand U18519 (N_18519,N_16604,N_16414);
nand U18520 (N_18520,N_17693,N_17658);
nor U18521 (N_18521,N_16420,N_16619);
or U18522 (N_18522,N_16871,N_17374);
nor U18523 (N_18523,N_17808,N_17126);
or U18524 (N_18524,N_17920,N_17193);
or U18525 (N_18525,N_17004,N_16781);
nand U18526 (N_18526,N_17653,N_16934);
or U18527 (N_18527,N_16862,N_17682);
and U18528 (N_18528,N_16598,N_17911);
and U18529 (N_18529,N_16431,N_16370);
or U18530 (N_18530,N_16820,N_16608);
nand U18531 (N_18531,N_17468,N_17145);
nor U18532 (N_18532,N_17832,N_17459);
or U18533 (N_18533,N_17271,N_16411);
nor U18534 (N_18534,N_16857,N_17301);
nand U18535 (N_18535,N_16379,N_17463);
xor U18536 (N_18536,N_17335,N_17866);
or U18537 (N_18537,N_16203,N_16040);
nand U18538 (N_18538,N_17323,N_17453);
nand U18539 (N_18539,N_16196,N_17079);
xnor U18540 (N_18540,N_16618,N_16571);
and U18541 (N_18541,N_16915,N_16988);
or U18542 (N_18542,N_17488,N_16937);
xnor U18543 (N_18543,N_17841,N_17597);
or U18544 (N_18544,N_17675,N_17076);
xor U18545 (N_18545,N_16771,N_17616);
and U18546 (N_18546,N_17927,N_16998);
and U18547 (N_18547,N_16913,N_16996);
nor U18548 (N_18548,N_16556,N_17410);
and U18549 (N_18549,N_17169,N_16038);
or U18550 (N_18550,N_16560,N_16856);
and U18551 (N_18551,N_16908,N_17230);
and U18552 (N_18552,N_17239,N_17691);
and U18553 (N_18553,N_17435,N_16939);
nand U18554 (N_18554,N_16940,N_16677);
xor U18555 (N_18555,N_16713,N_17377);
and U18556 (N_18556,N_16077,N_16881);
and U18557 (N_18557,N_17709,N_16369);
and U18558 (N_18558,N_17557,N_17890);
nand U18559 (N_18559,N_16116,N_17989);
nand U18560 (N_18560,N_16009,N_17891);
xnor U18561 (N_18561,N_16640,N_17892);
nand U18562 (N_18562,N_17922,N_17739);
nor U18563 (N_18563,N_17515,N_16695);
xnor U18564 (N_18564,N_17117,N_17707);
or U18565 (N_18565,N_17633,N_17728);
nand U18566 (N_18566,N_17098,N_16089);
nor U18567 (N_18567,N_16892,N_16240);
nor U18568 (N_18568,N_17112,N_17517);
or U18569 (N_18569,N_16162,N_16449);
or U18570 (N_18570,N_17274,N_16928);
and U18571 (N_18571,N_16221,N_16529);
nand U18572 (N_18572,N_17518,N_17406);
nand U18573 (N_18573,N_17082,N_17178);
and U18574 (N_18574,N_16337,N_16265);
nand U18575 (N_18575,N_16740,N_17512);
nor U18576 (N_18576,N_17713,N_16194);
xnor U18577 (N_18577,N_17577,N_16824);
and U18578 (N_18578,N_16945,N_17770);
xnor U18579 (N_18579,N_16387,N_17738);
and U18580 (N_18580,N_16049,N_16914);
or U18581 (N_18581,N_17626,N_16652);
xnor U18582 (N_18582,N_17578,N_16318);
or U18583 (N_18583,N_17747,N_17627);
and U18584 (N_18584,N_17710,N_16788);
nor U18585 (N_18585,N_16663,N_16701);
nor U18586 (N_18586,N_16610,N_16004);
nor U18587 (N_18587,N_17533,N_16763);
nand U18588 (N_18588,N_16358,N_16094);
nand U18589 (N_18589,N_17932,N_16290);
nor U18590 (N_18590,N_16898,N_16951);
nand U18591 (N_18591,N_16139,N_16669);
xnor U18592 (N_18592,N_17457,N_17733);
or U18593 (N_18593,N_17083,N_16724);
nand U18594 (N_18594,N_17889,N_17231);
nor U18595 (N_18595,N_16656,N_16926);
nor U18596 (N_18596,N_16118,N_16454);
nand U18597 (N_18597,N_17655,N_16064);
nor U18598 (N_18598,N_17199,N_17561);
or U18599 (N_18599,N_16955,N_16594);
or U18600 (N_18600,N_17089,N_16427);
or U18601 (N_18601,N_16643,N_17660);
or U18602 (N_18602,N_16665,N_16255);
nand U18603 (N_18603,N_17600,N_16687);
nor U18604 (N_18604,N_16516,N_17149);
xor U18605 (N_18605,N_16275,N_16965);
or U18606 (N_18606,N_16486,N_17901);
nand U18607 (N_18607,N_16428,N_16916);
nand U18608 (N_18608,N_16759,N_16041);
and U18609 (N_18609,N_17672,N_17566);
nor U18610 (N_18610,N_16995,N_16950);
nand U18611 (N_18611,N_16658,N_17507);
xnor U18612 (N_18612,N_16661,N_17125);
or U18613 (N_18613,N_16006,N_16851);
nor U18614 (N_18614,N_16160,N_16615);
xor U18615 (N_18615,N_16664,N_17315);
and U18616 (N_18616,N_17443,N_16407);
or U18617 (N_18617,N_17659,N_16052);
xor U18618 (N_18618,N_16144,N_17640);
nor U18619 (N_18619,N_17591,N_17252);
nand U18620 (N_18620,N_16849,N_16352);
nor U18621 (N_18621,N_16708,N_17160);
nand U18622 (N_18622,N_17197,N_17974);
nand U18623 (N_18623,N_17777,N_16622);
and U18624 (N_18624,N_16887,N_16151);
and U18625 (N_18625,N_16509,N_16389);
nand U18626 (N_18626,N_17107,N_16467);
and U18627 (N_18627,N_16706,N_17404);
nor U18628 (N_18628,N_17148,N_17909);
and U18629 (N_18629,N_17122,N_16754);
nor U18630 (N_18630,N_16842,N_16201);
nor U18631 (N_18631,N_17242,N_17730);
nor U18632 (N_18632,N_17860,N_16320);
and U18633 (N_18633,N_17289,N_16808);
or U18634 (N_18634,N_17753,N_17810);
and U18635 (N_18635,N_17645,N_16815);
nand U18636 (N_18636,N_17081,N_17092);
nand U18637 (N_18637,N_17732,N_16013);
nand U18638 (N_18638,N_17386,N_17641);
nand U18639 (N_18639,N_16544,N_16990);
nor U18640 (N_18640,N_16681,N_17164);
and U18641 (N_18641,N_17322,N_17646);
nor U18642 (N_18642,N_17919,N_16152);
or U18643 (N_18643,N_17448,N_17910);
nand U18644 (N_18644,N_17611,N_16605);
and U18645 (N_18645,N_17936,N_17867);
xnor U18646 (N_18646,N_16120,N_17605);
and U18647 (N_18647,N_17543,N_17341);
nand U18648 (N_18648,N_17531,N_17058);
nor U18649 (N_18649,N_16055,N_16925);
nor U18650 (N_18650,N_17853,N_17142);
xor U18651 (N_18651,N_17300,N_16384);
nand U18652 (N_18652,N_17138,N_16791);
and U18653 (N_18653,N_17102,N_16577);
xor U18654 (N_18654,N_17203,N_17033);
and U18655 (N_18655,N_17269,N_17427);
nor U18656 (N_18656,N_16956,N_16286);
nor U18657 (N_18657,N_17773,N_17628);
nand U18658 (N_18658,N_17075,N_17902);
and U18659 (N_18659,N_16121,N_16711);
xnor U18660 (N_18660,N_16624,N_16966);
and U18661 (N_18661,N_17714,N_16183);
or U18662 (N_18662,N_17153,N_16547);
and U18663 (N_18663,N_16087,N_16117);
nor U18664 (N_18664,N_17893,N_17288);
nand U18665 (N_18665,N_17261,N_16645);
or U18666 (N_18666,N_17418,N_16075);
and U18667 (N_18667,N_17487,N_16766);
and U18668 (N_18668,N_16091,N_16696);
xnor U18669 (N_18669,N_16097,N_16123);
nand U18670 (N_18670,N_16631,N_16301);
or U18671 (N_18671,N_17212,N_17156);
nand U18672 (N_18672,N_17342,N_17346);
and U18673 (N_18673,N_16630,N_17241);
nand U18674 (N_18674,N_17106,N_17952);
nor U18675 (N_18675,N_16169,N_17724);
or U18676 (N_18676,N_17451,N_16848);
nand U18677 (N_18677,N_17415,N_17043);
and U18678 (N_18678,N_17791,N_17373);
nand U18679 (N_18679,N_16961,N_17726);
nand U18680 (N_18680,N_16235,N_16256);
or U18681 (N_18681,N_16267,N_17010);
nand U18682 (N_18682,N_17522,N_16127);
nor U18683 (N_18683,N_17303,N_17099);
or U18684 (N_18684,N_16292,N_17564);
nand U18685 (N_18685,N_17258,N_16276);
or U18686 (N_18686,N_16519,N_16623);
or U18687 (N_18687,N_16884,N_17224);
nand U18688 (N_18688,N_16515,N_16363);
xnor U18689 (N_18689,N_16460,N_16756);
nand U18690 (N_18690,N_17743,N_17349);
and U18691 (N_18691,N_17715,N_16000);
nor U18692 (N_18692,N_17256,N_16590);
nor U18693 (N_18693,N_16470,N_17520);
and U18694 (N_18694,N_16784,N_16762);
nor U18695 (N_18695,N_16231,N_16855);
nor U18696 (N_18696,N_16530,N_17446);
nand U18697 (N_18697,N_16279,N_17084);
and U18698 (N_18698,N_17537,N_16559);
nor U18699 (N_18699,N_16404,N_16921);
or U18700 (N_18700,N_16599,N_17546);
xnor U18701 (N_18701,N_17779,N_17285);
and U18702 (N_18702,N_16469,N_17607);
and U18703 (N_18703,N_17734,N_17159);
or U18704 (N_18704,N_17608,N_16903);
nand U18705 (N_18705,N_17347,N_17251);
or U18706 (N_18706,N_17671,N_17455);
and U18707 (N_18707,N_17331,N_16497);
or U18708 (N_18708,N_17697,N_17895);
nor U18709 (N_18709,N_17226,N_17223);
nor U18710 (N_18710,N_16636,N_17722);
nand U18711 (N_18711,N_17720,N_16331);
xnor U18712 (N_18712,N_17698,N_16029);
nor U18713 (N_18713,N_17277,N_16309);
nand U18714 (N_18714,N_17654,N_16350);
or U18715 (N_18715,N_16197,N_16948);
nor U18716 (N_18716,N_17516,N_16983);
and U18717 (N_18717,N_16225,N_16185);
and U18718 (N_18718,N_17766,N_16660);
and U18719 (N_18719,N_17706,N_16860);
nand U18720 (N_18720,N_17210,N_16080);
and U18721 (N_18721,N_17497,N_16974);
nor U18722 (N_18722,N_16226,N_17297);
nand U18723 (N_18723,N_17332,N_17986);
xor U18724 (N_18724,N_17897,N_17673);
nand U18725 (N_18725,N_17311,N_16257);
and U18726 (N_18726,N_16971,N_17325);
or U18727 (N_18727,N_16175,N_16398);
nand U18728 (N_18728,N_16628,N_16728);
nor U18729 (N_18729,N_16812,N_17674);
nor U18730 (N_18730,N_16807,N_17802);
or U18731 (N_18731,N_16046,N_16694);
nor U18732 (N_18732,N_16101,N_17934);
or U18733 (N_18733,N_16684,N_17372);
nor U18734 (N_18734,N_17007,N_16452);
and U18735 (N_18735,N_17886,N_16528);
and U18736 (N_18736,N_17317,N_16330);
nand U18737 (N_18737,N_17751,N_17044);
and U18738 (N_18738,N_16214,N_16507);
or U18739 (N_18739,N_16440,N_17180);
xor U18740 (N_18740,N_17175,N_17209);
or U18741 (N_18741,N_16846,N_17805);
or U18742 (N_18742,N_16518,N_16672);
nor U18743 (N_18743,N_17057,N_17774);
and U18744 (N_18744,N_17304,N_16471);
nor U18745 (N_18745,N_17474,N_16317);
nor U18746 (N_18746,N_16403,N_16247);
nor U18747 (N_18747,N_17108,N_17563);
nor U18748 (N_18748,N_17165,N_16744);
and U18749 (N_18749,N_17422,N_16741);
nand U18750 (N_18750,N_17817,N_17174);
nand U18751 (N_18751,N_16187,N_17632);
xor U18752 (N_18752,N_17218,N_16703);
and U18753 (N_18753,N_16326,N_17190);
and U18754 (N_18754,N_17823,N_16367);
and U18755 (N_18755,N_16748,N_17123);
xnor U18756 (N_18756,N_16569,N_16997);
or U18757 (N_18757,N_16858,N_16078);
nand U18758 (N_18758,N_17701,N_17944);
and U18759 (N_18759,N_17978,N_17510);
nor U18760 (N_18760,N_17740,N_17324);
and U18761 (N_18761,N_17976,N_16709);
and U18762 (N_18762,N_17365,N_17762);
xor U18763 (N_18763,N_17176,N_16218);
nor U18764 (N_18764,N_17026,N_17822);
or U18765 (N_18765,N_16823,N_17759);
nor U18766 (N_18766,N_17019,N_17042);
nor U18767 (N_18767,N_16051,N_17894);
nand U18768 (N_18768,N_16895,N_16526);
xnor U18769 (N_18769,N_17306,N_16931);
nor U18770 (N_18770,N_17940,N_17465);
nor U18771 (N_18771,N_16217,N_16319);
nand U18772 (N_18772,N_17846,N_16161);
and U18773 (N_18773,N_16739,N_17202);
nand U18774 (N_18774,N_16639,N_17458);
or U18775 (N_18775,N_16960,N_16083);
and U18776 (N_18776,N_16416,N_17998);
or U18777 (N_18777,N_16964,N_17606);
nand U18778 (N_18778,N_17268,N_16165);
and U18779 (N_18779,N_16246,N_16976);
nand U18780 (N_18780,N_16742,N_17154);
nor U18781 (N_18781,N_16322,N_16843);
and U18782 (N_18782,N_17388,N_17403);
or U18783 (N_18783,N_17469,N_17551);
nand U18784 (N_18784,N_17970,N_17931);
nand U18785 (N_18785,N_17957,N_17215);
and U18786 (N_18786,N_17973,N_17028);
and U18787 (N_18787,N_16810,N_17187);
and U18788 (N_18788,N_16417,N_17999);
nor U18789 (N_18789,N_17620,N_17758);
xor U18790 (N_18790,N_16239,N_16557);
nor U18791 (N_18791,N_17104,N_17400);
nand U18792 (N_18792,N_17339,N_16167);
nor U18793 (N_18793,N_16018,N_16817);
nor U18794 (N_18794,N_17320,N_16804);
nor U18795 (N_18795,N_16396,N_16298);
or U18796 (N_18796,N_16541,N_17227);
nand U18797 (N_18797,N_17572,N_17442);
xor U18798 (N_18798,N_16568,N_16426);
nand U18799 (N_18799,N_16593,N_16944);
and U18800 (N_18800,N_16069,N_17535);
nor U18801 (N_18801,N_16570,N_16888);
or U18802 (N_18802,N_17454,N_17649);
nand U18803 (N_18803,N_16109,N_16962);
nand U18804 (N_18804,N_16368,N_17219);
or U18805 (N_18805,N_16793,N_16476);
or U18806 (N_18806,N_17490,N_16520);
nand U18807 (N_18807,N_17035,N_17840);
or U18808 (N_18808,N_16132,N_17091);
nor U18809 (N_18809,N_16952,N_17767);
nor U18810 (N_18810,N_16886,N_16119);
nand U18811 (N_18811,N_16718,N_17140);
nor U18812 (N_18812,N_17216,N_17635);
xor U18813 (N_18813,N_16001,N_17200);
and U18814 (N_18814,N_17596,N_17355);
xor U18815 (N_18815,N_17013,N_16030);
nand U18816 (N_18816,N_17135,N_17383);
nor U18817 (N_18817,N_17745,N_16555);
nor U18818 (N_18818,N_16307,N_16573);
xor U18819 (N_18819,N_16133,N_17170);
or U18820 (N_18820,N_17558,N_16372);
nand U18821 (N_18821,N_16248,N_16216);
or U18822 (N_18822,N_17316,N_17785);
or U18823 (N_18823,N_16685,N_16300);
or U18824 (N_18824,N_16638,N_16044);
or U18825 (N_18825,N_17157,N_16053);
or U18826 (N_18826,N_17313,N_16446);
and U18827 (N_18827,N_17871,N_16609);
or U18828 (N_18828,N_16662,N_16933);
and U18829 (N_18829,N_17629,N_16700);
nand U18830 (N_18830,N_17621,N_17243);
or U18831 (N_18831,N_17863,N_16021);
nand U18832 (N_18832,N_17668,N_16361);
nand U18833 (N_18833,N_17887,N_17783);
or U18834 (N_18834,N_17718,N_16386);
nor U18835 (N_18835,N_17604,N_17792);
and U18836 (N_18836,N_17638,N_16202);
nor U18837 (N_18837,N_17993,N_16649);
or U18838 (N_18838,N_17689,N_17908);
or U18839 (N_18839,N_16063,N_16514);
nor U18840 (N_18840,N_16496,N_16321);
nor U18841 (N_18841,N_17120,N_17351);
nor U18842 (N_18842,N_17283,N_17298);
nor U18843 (N_18843,N_16482,N_16801);
and U18844 (N_18844,N_17039,N_17634);
and U18845 (N_18845,N_16062,N_17794);
nor U18846 (N_18846,N_16912,N_16128);
nor U18847 (N_18847,N_17498,N_16212);
and U18848 (N_18848,N_16475,N_16586);
xnor U18849 (N_18849,N_17544,N_17310);
and U18850 (N_18850,N_17399,N_17094);
xnor U18851 (N_18851,N_16967,N_16270);
nand U18852 (N_18852,N_16790,N_17760);
nor U18853 (N_18853,N_16024,N_16081);
nand U18854 (N_18854,N_17370,N_16829);
nand U18855 (N_18855,N_17678,N_17559);
nand U18856 (N_18856,N_17472,N_17362);
and U18857 (N_18857,N_17684,N_17806);
and U18858 (N_18858,N_16535,N_16822);
or U18859 (N_18859,N_16436,N_16488);
or U18860 (N_18860,N_17358,N_16413);
nand U18861 (N_18861,N_16325,N_16830);
nand U18862 (N_18862,N_16504,N_16795);
nor U18863 (N_18863,N_16864,N_17884);
nor U18864 (N_18864,N_17266,N_16375);
nor U18865 (N_18865,N_17492,N_17101);
or U18866 (N_18866,N_17757,N_17719);
nor U18867 (N_18867,N_17095,N_16122);
and U18868 (N_18868,N_17850,N_17935);
or U18869 (N_18869,N_16258,N_16512);
and U18870 (N_18870,N_17855,N_16850);
and U18871 (N_18871,N_16354,N_16890);
nor U18872 (N_18872,N_17503,N_17565);
and U18873 (N_18873,N_16374,N_17979);
nand U18874 (N_18874,N_16193,N_17619);
and U18875 (N_18875,N_17096,N_16283);
nand U18876 (N_18876,N_17670,N_16770);
and U18877 (N_18877,N_16523,N_17798);
xnor U18878 (N_18878,N_17364,N_17925);
or U18879 (N_18879,N_17787,N_16280);
or U18880 (N_18880,N_17121,N_17988);
and U18881 (N_18881,N_17208,N_17248);
nor U18882 (N_18882,N_16617,N_16992);
and U18883 (N_18883,N_16010,N_16282);
nor U18884 (N_18884,N_16479,N_17294);
nor U18885 (N_18885,N_16595,N_16020);
and U18886 (N_18886,N_16786,N_17220);
or U18887 (N_18887,N_17247,N_17444);
or U18888 (N_18888,N_17837,N_17353);
xor U18889 (N_18889,N_17508,N_17538);
nand U18890 (N_18890,N_16821,N_16875);
nor U18891 (N_18891,N_16972,N_16932);
nor U18892 (N_18892,N_17567,N_16899);
and U18893 (N_18893,N_17879,N_17257);
or U18894 (N_18894,N_17966,N_16521);
and U18895 (N_18895,N_17380,N_17540);
xnor U18896 (N_18896,N_17534,N_16505);
and U18897 (N_18897,N_17063,N_16909);
and U18898 (N_18898,N_16927,N_17987);
and U18899 (N_18899,N_17093,N_17971);
nor U18900 (N_18900,N_17921,N_16016);
and U18901 (N_18901,N_16947,N_17228);
nand U18902 (N_18902,N_17205,N_17651);
and U18903 (N_18903,N_17072,N_16904);
nor U18904 (N_18904,N_16498,N_17214);
nand U18905 (N_18905,N_16134,N_17661);
xor U18906 (N_18906,N_17813,N_16510);
and U18907 (N_18907,N_17669,N_17968);
nand U18908 (N_18908,N_16929,N_16263);
nor U18909 (N_18909,N_16818,N_16287);
xnor U18910 (N_18910,N_16455,N_17755);
and U18911 (N_18911,N_16395,N_17392);
and U18912 (N_18912,N_17168,N_17833);
xnor U18913 (N_18913,N_16954,N_16902);
or U18914 (N_18914,N_17319,N_17609);
nor U18915 (N_18915,N_17246,N_17273);
nor U18916 (N_18916,N_17417,N_16924);
and U18917 (N_18917,N_16058,N_16140);
or U18918 (N_18918,N_17780,N_16585);
and U18919 (N_18919,N_17969,N_17166);
and U18920 (N_18920,N_17569,N_17161);
or U18921 (N_18921,N_17541,N_16277);
nor U18922 (N_18922,N_17182,N_16868);
or U18923 (N_18923,N_17130,N_17456);
and U18924 (N_18924,N_16359,N_17481);
and U18925 (N_18925,N_16987,N_16084);
nor U18926 (N_18926,N_17053,N_17278);
xnor U18927 (N_18927,N_17078,N_16936);
nor U18928 (N_18928,N_17087,N_17479);
nor U18929 (N_18929,N_16388,N_17858);
and U18930 (N_18930,N_17097,N_17366);
xor U18931 (N_18931,N_17526,N_17236);
and U18932 (N_18932,N_17020,N_16158);
nor U18933 (N_18933,N_16633,N_17384);
or U18934 (N_18934,N_17441,N_17648);
or U18935 (N_18935,N_17929,N_17050);
xor U18936 (N_18936,N_17027,N_16085);
nand U18937 (N_18937,N_16315,N_16811);
xor U18938 (N_18938,N_17797,N_16189);
and U18939 (N_18939,N_16391,N_17690);
and U18940 (N_18940,N_17466,N_17402);
and U18941 (N_18941,N_16131,N_16474);
xor U18942 (N_18942,N_17527,N_16755);
or U18943 (N_18943,N_17815,N_17788);
nor U18944 (N_18944,N_17069,N_16238);
nor U18945 (N_18945,N_16539,N_17975);
and U18946 (N_18946,N_16110,N_17445);
nor U18947 (N_18947,N_17232,N_16213);
or U18948 (N_18948,N_17431,N_16970);
and U18949 (N_18949,N_17461,N_16517);
nand U18950 (N_18950,N_16499,N_16861);
or U18951 (N_18951,N_17610,N_17746);
or U18952 (N_18952,N_17137,N_17814);
and U18953 (N_18953,N_17143,N_16493);
nand U18954 (N_18954,N_17820,N_17238);
nand U18955 (N_18955,N_17426,N_17308);
and U18956 (N_18956,N_17790,N_17359);
nor U18957 (N_18957,N_17536,N_16362);
and U18958 (N_18958,N_17592,N_16364);
and U18959 (N_18959,N_16086,N_16180);
and U18960 (N_18960,N_17022,N_17192);
nor U18961 (N_18961,N_17421,N_17177);
nor U18962 (N_18962,N_17826,N_16879);
xor U18963 (N_18963,N_16206,N_16574);
and U18964 (N_18964,N_17524,N_16176);
or U18965 (N_18965,N_16707,N_16190);
or U18966 (N_18966,N_17857,N_16558);
xnor U18967 (N_18967,N_17068,N_16825);
and U18968 (N_18968,N_16838,N_17307);
and U18969 (N_18969,N_16985,N_17263);
and U18970 (N_18970,N_17829,N_17955);
nor U18971 (N_18971,N_17644,N_16429);
or U18972 (N_18972,N_17034,N_16866);
or U18973 (N_18973,N_17132,N_16274);
and U18974 (N_18974,N_17350,N_17647);
or U18975 (N_18975,N_16271,N_17314);
nand U18976 (N_18976,N_17800,N_17144);
nand U18977 (N_18977,N_16723,N_17495);
or U18978 (N_18978,N_16968,N_16472);
nor U18979 (N_18979,N_17623,N_16600);
nand U18980 (N_18980,N_17703,N_17006);
nor U18981 (N_18981,N_17360,N_16108);
nand U18982 (N_18982,N_16634,N_16303);
nand U18983 (N_18983,N_16186,N_17424);
nor U18984 (N_18984,N_16096,N_16543);
and U18985 (N_18985,N_16973,N_17483);
nor U18986 (N_18986,N_17496,N_16048);
and U18987 (N_18987,N_17103,N_16919);
nor U18988 (N_18988,N_16697,N_17229);
nand U18989 (N_18989,N_17234,N_16219);
nand U18990 (N_18990,N_16070,N_16533);
or U18991 (N_18991,N_17051,N_17363);
nand U18992 (N_18992,N_16532,N_16459);
or U18993 (N_18993,N_16705,N_17990);
nand U18994 (N_18994,N_16192,N_16114);
or U18995 (N_18995,N_16720,N_16796);
nand U18996 (N_18996,N_17394,N_16065);
nand U18997 (N_18997,N_17327,N_17131);
or U18998 (N_18998,N_17625,N_17917);
and U18999 (N_18999,N_16894,N_16061);
nor U19000 (N_19000,N_16188,N_17283);
nand U19001 (N_19001,N_16665,N_16269);
and U19002 (N_19002,N_17888,N_16628);
nand U19003 (N_19003,N_16413,N_16162);
or U19004 (N_19004,N_17993,N_17724);
or U19005 (N_19005,N_17228,N_17547);
or U19006 (N_19006,N_17809,N_17112);
nand U19007 (N_19007,N_17502,N_17132);
and U19008 (N_19008,N_16765,N_16923);
nand U19009 (N_19009,N_17702,N_17560);
and U19010 (N_19010,N_17075,N_17680);
and U19011 (N_19011,N_17652,N_16255);
or U19012 (N_19012,N_17836,N_17387);
nor U19013 (N_19013,N_17029,N_17255);
nand U19014 (N_19014,N_16156,N_17456);
nand U19015 (N_19015,N_17886,N_17299);
or U19016 (N_19016,N_17575,N_16855);
and U19017 (N_19017,N_16876,N_16745);
and U19018 (N_19018,N_16685,N_17047);
nor U19019 (N_19019,N_17760,N_16688);
nor U19020 (N_19020,N_16630,N_16996);
or U19021 (N_19021,N_16106,N_16657);
and U19022 (N_19022,N_16934,N_17841);
and U19023 (N_19023,N_16522,N_17067);
and U19024 (N_19024,N_17336,N_17079);
nand U19025 (N_19025,N_16154,N_16801);
nand U19026 (N_19026,N_17609,N_16334);
xor U19027 (N_19027,N_17226,N_16705);
and U19028 (N_19028,N_17699,N_16495);
or U19029 (N_19029,N_17872,N_16713);
or U19030 (N_19030,N_16295,N_16391);
nor U19031 (N_19031,N_17306,N_16342);
and U19032 (N_19032,N_17721,N_17304);
nor U19033 (N_19033,N_16856,N_16236);
or U19034 (N_19034,N_16932,N_17824);
and U19035 (N_19035,N_16691,N_17606);
nand U19036 (N_19036,N_16187,N_16789);
and U19037 (N_19037,N_17106,N_17982);
xnor U19038 (N_19038,N_16552,N_16753);
or U19039 (N_19039,N_16407,N_17598);
nor U19040 (N_19040,N_17962,N_17630);
nor U19041 (N_19041,N_17578,N_17170);
nand U19042 (N_19042,N_17785,N_17158);
and U19043 (N_19043,N_16548,N_17097);
nand U19044 (N_19044,N_17215,N_16138);
nor U19045 (N_19045,N_17316,N_16470);
and U19046 (N_19046,N_16016,N_17740);
xor U19047 (N_19047,N_16577,N_17836);
xor U19048 (N_19048,N_16716,N_17440);
and U19049 (N_19049,N_16711,N_16268);
nand U19050 (N_19050,N_17754,N_17050);
nand U19051 (N_19051,N_16518,N_17688);
nand U19052 (N_19052,N_17875,N_17295);
nor U19053 (N_19053,N_17199,N_16095);
or U19054 (N_19054,N_16964,N_17234);
or U19055 (N_19055,N_17775,N_16507);
and U19056 (N_19056,N_16972,N_16061);
nor U19057 (N_19057,N_16470,N_17990);
nor U19058 (N_19058,N_17601,N_16889);
and U19059 (N_19059,N_17937,N_17593);
or U19060 (N_19060,N_16138,N_17473);
nand U19061 (N_19061,N_17638,N_16428);
nand U19062 (N_19062,N_17661,N_16224);
and U19063 (N_19063,N_16800,N_16421);
nand U19064 (N_19064,N_17478,N_17913);
nand U19065 (N_19065,N_16758,N_16131);
nand U19066 (N_19066,N_17161,N_16031);
and U19067 (N_19067,N_17200,N_16039);
and U19068 (N_19068,N_17278,N_17689);
or U19069 (N_19069,N_17557,N_17112);
nand U19070 (N_19070,N_16105,N_17585);
or U19071 (N_19071,N_16401,N_16595);
nand U19072 (N_19072,N_16811,N_16386);
and U19073 (N_19073,N_16466,N_16648);
nand U19074 (N_19074,N_17066,N_17284);
or U19075 (N_19075,N_16001,N_17692);
xnor U19076 (N_19076,N_17191,N_16009);
nand U19077 (N_19077,N_16245,N_16806);
xnor U19078 (N_19078,N_17216,N_16401);
xnor U19079 (N_19079,N_16674,N_17069);
nor U19080 (N_19080,N_16938,N_17685);
or U19081 (N_19081,N_16836,N_16151);
and U19082 (N_19082,N_17480,N_16892);
nor U19083 (N_19083,N_17593,N_17694);
or U19084 (N_19084,N_16606,N_17870);
nor U19085 (N_19085,N_16095,N_16191);
and U19086 (N_19086,N_17048,N_17021);
nor U19087 (N_19087,N_17013,N_17522);
nand U19088 (N_19088,N_16655,N_17811);
xor U19089 (N_19089,N_16968,N_17655);
or U19090 (N_19090,N_17112,N_17800);
xor U19091 (N_19091,N_17222,N_16444);
nor U19092 (N_19092,N_16652,N_17492);
or U19093 (N_19093,N_17788,N_16988);
and U19094 (N_19094,N_16732,N_16256);
and U19095 (N_19095,N_17013,N_17921);
and U19096 (N_19096,N_16165,N_16315);
nand U19097 (N_19097,N_16960,N_16112);
or U19098 (N_19098,N_17556,N_17105);
or U19099 (N_19099,N_16329,N_17692);
xnor U19100 (N_19100,N_16499,N_16911);
nand U19101 (N_19101,N_16654,N_16730);
or U19102 (N_19102,N_17868,N_16978);
and U19103 (N_19103,N_17873,N_17904);
nand U19104 (N_19104,N_17553,N_17918);
nand U19105 (N_19105,N_17289,N_16890);
xnor U19106 (N_19106,N_16632,N_16892);
or U19107 (N_19107,N_16740,N_16043);
nor U19108 (N_19108,N_16427,N_16330);
nand U19109 (N_19109,N_17547,N_17502);
nor U19110 (N_19110,N_17329,N_16689);
nand U19111 (N_19111,N_16081,N_16616);
nor U19112 (N_19112,N_16461,N_17881);
or U19113 (N_19113,N_16589,N_17512);
nor U19114 (N_19114,N_16386,N_16085);
xor U19115 (N_19115,N_17641,N_16563);
or U19116 (N_19116,N_16313,N_17358);
and U19117 (N_19117,N_17759,N_17067);
nor U19118 (N_19118,N_16560,N_17553);
and U19119 (N_19119,N_16021,N_17721);
and U19120 (N_19120,N_16673,N_17093);
nor U19121 (N_19121,N_17487,N_16546);
xor U19122 (N_19122,N_16300,N_17165);
nand U19123 (N_19123,N_16611,N_17568);
nand U19124 (N_19124,N_16567,N_16214);
xor U19125 (N_19125,N_17571,N_16225);
nand U19126 (N_19126,N_17491,N_16964);
nand U19127 (N_19127,N_16622,N_16204);
xor U19128 (N_19128,N_16978,N_17943);
nor U19129 (N_19129,N_17860,N_16638);
nor U19130 (N_19130,N_17077,N_16689);
or U19131 (N_19131,N_16858,N_16087);
and U19132 (N_19132,N_17191,N_17604);
nand U19133 (N_19133,N_17621,N_16554);
xor U19134 (N_19134,N_16205,N_17657);
nand U19135 (N_19135,N_16895,N_17814);
nor U19136 (N_19136,N_17147,N_17955);
or U19137 (N_19137,N_17882,N_17496);
nand U19138 (N_19138,N_17761,N_17094);
and U19139 (N_19139,N_17931,N_16430);
nor U19140 (N_19140,N_17348,N_16403);
nand U19141 (N_19141,N_16422,N_17634);
or U19142 (N_19142,N_17558,N_17244);
nor U19143 (N_19143,N_17829,N_16213);
nor U19144 (N_19144,N_16874,N_16772);
nand U19145 (N_19145,N_17632,N_16915);
nor U19146 (N_19146,N_16349,N_17414);
nor U19147 (N_19147,N_17449,N_16197);
or U19148 (N_19148,N_17716,N_16111);
or U19149 (N_19149,N_17826,N_16478);
or U19150 (N_19150,N_17677,N_16800);
nor U19151 (N_19151,N_16762,N_16288);
nand U19152 (N_19152,N_17295,N_17008);
or U19153 (N_19153,N_17060,N_16353);
or U19154 (N_19154,N_16547,N_17348);
and U19155 (N_19155,N_16153,N_16388);
nor U19156 (N_19156,N_17408,N_17261);
nor U19157 (N_19157,N_17938,N_17702);
nor U19158 (N_19158,N_16042,N_17462);
nand U19159 (N_19159,N_17277,N_16824);
nand U19160 (N_19160,N_17221,N_16469);
nand U19161 (N_19161,N_16119,N_16647);
and U19162 (N_19162,N_17256,N_16041);
or U19163 (N_19163,N_17133,N_17624);
xor U19164 (N_19164,N_17349,N_17961);
xor U19165 (N_19165,N_17749,N_17225);
nand U19166 (N_19166,N_17308,N_16477);
or U19167 (N_19167,N_16978,N_16883);
or U19168 (N_19168,N_16487,N_16372);
nor U19169 (N_19169,N_16587,N_17005);
or U19170 (N_19170,N_17448,N_17418);
and U19171 (N_19171,N_16662,N_16400);
nor U19172 (N_19172,N_16352,N_16852);
nand U19173 (N_19173,N_17124,N_17175);
nor U19174 (N_19174,N_16448,N_17368);
and U19175 (N_19175,N_17513,N_16221);
or U19176 (N_19176,N_16711,N_16421);
or U19177 (N_19177,N_16909,N_16207);
and U19178 (N_19178,N_17181,N_17318);
nand U19179 (N_19179,N_16249,N_17121);
nand U19180 (N_19180,N_16745,N_17259);
xor U19181 (N_19181,N_17011,N_17682);
and U19182 (N_19182,N_16053,N_16106);
or U19183 (N_19183,N_16068,N_16661);
nand U19184 (N_19184,N_17304,N_17454);
or U19185 (N_19185,N_16514,N_17034);
nor U19186 (N_19186,N_17309,N_17560);
nand U19187 (N_19187,N_17209,N_17446);
or U19188 (N_19188,N_16074,N_16416);
and U19189 (N_19189,N_16527,N_17479);
and U19190 (N_19190,N_16385,N_17754);
and U19191 (N_19191,N_17812,N_16190);
or U19192 (N_19192,N_16992,N_17737);
nand U19193 (N_19193,N_17771,N_16224);
nand U19194 (N_19194,N_17717,N_16046);
and U19195 (N_19195,N_17118,N_17952);
nor U19196 (N_19196,N_16402,N_16692);
nor U19197 (N_19197,N_17797,N_17580);
xnor U19198 (N_19198,N_17197,N_17738);
nand U19199 (N_19199,N_16852,N_16502);
nand U19200 (N_19200,N_16215,N_16083);
xor U19201 (N_19201,N_17682,N_17065);
nand U19202 (N_19202,N_17140,N_16014);
nand U19203 (N_19203,N_17173,N_17192);
and U19204 (N_19204,N_16733,N_16306);
nand U19205 (N_19205,N_16714,N_17987);
or U19206 (N_19206,N_16857,N_17505);
nor U19207 (N_19207,N_17818,N_17415);
xnor U19208 (N_19208,N_16071,N_16485);
xor U19209 (N_19209,N_17982,N_17042);
nand U19210 (N_19210,N_16304,N_17604);
and U19211 (N_19211,N_17626,N_17035);
nand U19212 (N_19212,N_17162,N_16774);
nand U19213 (N_19213,N_17802,N_17031);
or U19214 (N_19214,N_16502,N_17788);
and U19215 (N_19215,N_16354,N_17713);
nor U19216 (N_19216,N_16418,N_17965);
xnor U19217 (N_19217,N_16455,N_17410);
xnor U19218 (N_19218,N_16540,N_16220);
nor U19219 (N_19219,N_16144,N_16492);
xnor U19220 (N_19220,N_16680,N_17791);
nor U19221 (N_19221,N_16029,N_17494);
or U19222 (N_19222,N_16058,N_17587);
or U19223 (N_19223,N_17434,N_16146);
nand U19224 (N_19224,N_17499,N_16373);
xnor U19225 (N_19225,N_16520,N_17600);
nor U19226 (N_19226,N_17976,N_16192);
nand U19227 (N_19227,N_17568,N_16048);
nor U19228 (N_19228,N_16445,N_16909);
or U19229 (N_19229,N_16275,N_16439);
and U19230 (N_19230,N_17638,N_16279);
xor U19231 (N_19231,N_16187,N_17405);
nor U19232 (N_19232,N_17456,N_16777);
nor U19233 (N_19233,N_17819,N_17482);
xor U19234 (N_19234,N_17221,N_16677);
xor U19235 (N_19235,N_16373,N_16975);
or U19236 (N_19236,N_16984,N_17684);
and U19237 (N_19237,N_16749,N_17702);
nor U19238 (N_19238,N_17710,N_17739);
and U19239 (N_19239,N_16242,N_17177);
or U19240 (N_19240,N_16523,N_16517);
nand U19241 (N_19241,N_17012,N_17718);
or U19242 (N_19242,N_17045,N_16084);
or U19243 (N_19243,N_16408,N_16247);
or U19244 (N_19244,N_17604,N_17617);
nand U19245 (N_19245,N_17799,N_16221);
and U19246 (N_19246,N_16344,N_16894);
nor U19247 (N_19247,N_17640,N_16079);
and U19248 (N_19248,N_16323,N_17366);
nand U19249 (N_19249,N_16112,N_16386);
and U19250 (N_19250,N_17106,N_17996);
and U19251 (N_19251,N_16053,N_17716);
and U19252 (N_19252,N_16969,N_17127);
and U19253 (N_19253,N_16513,N_17343);
or U19254 (N_19254,N_16783,N_16742);
or U19255 (N_19255,N_16537,N_17346);
nor U19256 (N_19256,N_16899,N_17588);
and U19257 (N_19257,N_16304,N_16116);
nand U19258 (N_19258,N_16479,N_16958);
or U19259 (N_19259,N_16169,N_17045);
or U19260 (N_19260,N_16067,N_17358);
nor U19261 (N_19261,N_17090,N_16345);
and U19262 (N_19262,N_17155,N_17380);
nor U19263 (N_19263,N_17531,N_17823);
nor U19264 (N_19264,N_17996,N_16868);
and U19265 (N_19265,N_17983,N_17531);
nand U19266 (N_19266,N_17333,N_17606);
nand U19267 (N_19267,N_16333,N_16912);
nand U19268 (N_19268,N_16842,N_17476);
nor U19269 (N_19269,N_16755,N_17689);
or U19270 (N_19270,N_16068,N_17412);
xor U19271 (N_19271,N_17541,N_17177);
xnor U19272 (N_19272,N_16740,N_16147);
and U19273 (N_19273,N_16698,N_17523);
nand U19274 (N_19274,N_16944,N_17343);
or U19275 (N_19275,N_16586,N_16240);
xnor U19276 (N_19276,N_16221,N_16848);
or U19277 (N_19277,N_16649,N_17341);
nand U19278 (N_19278,N_16462,N_16950);
nand U19279 (N_19279,N_17762,N_17904);
nand U19280 (N_19280,N_16623,N_17430);
and U19281 (N_19281,N_16526,N_17063);
nand U19282 (N_19282,N_16877,N_16850);
nor U19283 (N_19283,N_16634,N_17594);
or U19284 (N_19284,N_17476,N_17704);
and U19285 (N_19285,N_17873,N_16208);
or U19286 (N_19286,N_16710,N_17535);
nand U19287 (N_19287,N_16320,N_16887);
nand U19288 (N_19288,N_16209,N_16388);
and U19289 (N_19289,N_17352,N_17687);
nor U19290 (N_19290,N_17435,N_16188);
or U19291 (N_19291,N_16820,N_17469);
xor U19292 (N_19292,N_17443,N_17175);
nand U19293 (N_19293,N_16722,N_16350);
and U19294 (N_19294,N_16084,N_17146);
xor U19295 (N_19295,N_17865,N_17027);
or U19296 (N_19296,N_16117,N_16297);
and U19297 (N_19297,N_17984,N_16505);
nand U19298 (N_19298,N_17863,N_17205);
nand U19299 (N_19299,N_17068,N_16799);
or U19300 (N_19300,N_17787,N_17268);
nor U19301 (N_19301,N_17811,N_17553);
nand U19302 (N_19302,N_16069,N_17192);
or U19303 (N_19303,N_16449,N_16690);
nor U19304 (N_19304,N_17495,N_17552);
nor U19305 (N_19305,N_16431,N_16783);
and U19306 (N_19306,N_16894,N_16435);
and U19307 (N_19307,N_16487,N_17597);
and U19308 (N_19308,N_16699,N_16463);
nor U19309 (N_19309,N_16238,N_16474);
nand U19310 (N_19310,N_16752,N_16995);
or U19311 (N_19311,N_17946,N_16749);
or U19312 (N_19312,N_17660,N_17202);
and U19313 (N_19313,N_17466,N_17954);
and U19314 (N_19314,N_17342,N_16625);
nor U19315 (N_19315,N_17574,N_17657);
nor U19316 (N_19316,N_16344,N_16419);
nand U19317 (N_19317,N_16278,N_16821);
or U19318 (N_19318,N_17234,N_17068);
nor U19319 (N_19319,N_17707,N_17501);
nor U19320 (N_19320,N_16934,N_16940);
or U19321 (N_19321,N_17699,N_17748);
and U19322 (N_19322,N_16915,N_16568);
or U19323 (N_19323,N_16175,N_16375);
nand U19324 (N_19324,N_17598,N_16976);
nor U19325 (N_19325,N_16189,N_16787);
or U19326 (N_19326,N_16558,N_17035);
nand U19327 (N_19327,N_16417,N_16418);
and U19328 (N_19328,N_16383,N_16355);
and U19329 (N_19329,N_17678,N_17198);
nor U19330 (N_19330,N_17628,N_16903);
nand U19331 (N_19331,N_17279,N_17160);
and U19332 (N_19332,N_16141,N_16912);
xnor U19333 (N_19333,N_17444,N_16342);
nor U19334 (N_19334,N_16097,N_17607);
xor U19335 (N_19335,N_17176,N_17963);
xnor U19336 (N_19336,N_16056,N_16179);
or U19337 (N_19337,N_16014,N_16779);
nand U19338 (N_19338,N_17473,N_17102);
and U19339 (N_19339,N_16161,N_17514);
xor U19340 (N_19340,N_16660,N_16373);
and U19341 (N_19341,N_17260,N_16512);
nor U19342 (N_19342,N_16441,N_17200);
nand U19343 (N_19343,N_16942,N_16076);
and U19344 (N_19344,N_16274,N_17270);
xnor U19345 (N_19345,N_16047,N_16989);
and U19346 (N_19346,N_17582,N_16198);
and U19347 (N_19347,N_16044,N_17985);
nor U19348 (N_19348,N_16258,N_16911);
nand U19349 (N_19349,N_16312,N_17596);
and U19350 (N_19350,N_17082,N_17210);
or U19351 (N_19351,N_16276,N_17986);
xor U19352 (N_19352,N_17152,N_16554);
nand U19353 (N_19353,N_17980,N_16464);
nor U19354 (N_19354,N_17211,N_17384);
or U19355 (N_19355,N_17995,N_17630);
nor U19356 (N_19356,N_17992,N_16231);
and U19357 (N_19357,N_16904,N_17843);
nand U19358 (N_19358,N_17193,N_16880);
nor U19359 (N_19359,N_17819,N_16064);
or U19360 (N_19360,N_16512,N_17684);
or U19361 (N_19361,N_16877,N_16673);
nand U19362 (N_19362,N_16804,N_17893);
nor U19363 (N_19363,N_17459,N_17610);
nor U19364 (N_19364,N_17288,N_16343);
nand U19365 (N_19365,N_17890,N_16530);
nor U19366 (N_19366,N_17345,N_16345);
or U19367 (N_19367,N_16013,N_17843);
or U19368 (N_19368,N_17834,N_17169);
and U19369 (N_19369,N_17631,N_17528);
or U19370 (N_19370,N_16340,N_17689);
or U19371 (N_19371,N_17136,N_16066);
and U19372 (N_19372,N_16813,N_16788);
nand U19373 (N_19373,N_17305,N_16780);
or U19374 (N_19374,N_17941,N_17637);
nor U19375 (N_19375,N_17677,N_17866);
or U19376 (N_19376,N_17217,N_16480);
or U19377 (N_19377,N_17582,N_17885);
and U19378 (N_19378,N_16736,N_16416);
nor U19379 (N_19379,N_17105,N_17203);
or U19380 (N_19380,N_17026,N_17222);
xnor U19381 (N_19381,N_16850,N_17869);
or U19382 (N_19382,N_17469,N_16534);
and U19383 (N_19383,N_16247,N_16007);
nor U19384 (N_19384,N_16650,N_17024);
or U19385 (N_19385,N_16075,N_16608);
nor U19386 (N_19386,N_17677,N_16820);
nor U19387 (N_19387,N_17657,N_17150);
nor U19388 (N_19388,N_16268,N_16013);
or U19389 (N_19389,N_16198,N_16297);
xor U19390 (N_19390,N_16590,N_16298);
and U19391 (N_19391,N_16718,N_16414);
nor U19392 (N_19392,N_16093,N_16170);
nor U19393 (N_19393,N_16615,N_17963);
and U19394 (N_19394,N_17116,N_17731);
and U19395 (N_19395,N_16762,N_16272);
nor U19396 (N_19396,N_17316,N_17827);
nand U19397 (N_19397,N_17703,N_17154);
and U19398 (N_19398,N_16138,N_16064);
and U19399 (N_19399,N_17388,N_16784);
nor U19400 (N_19400,N_17981,N_16563);
nor U19401 (N_19401,N_16901,N_16342);
and U19402 (N_19402,N_16436,N_17685);
or U19403 (N_19403,N_17287,N_17180);
xnor U19404 (N_19404,N_16026,N_16998);
and U19405 (N_19405,N_16199,N_17228);
nand U19406 (N_19406,N_17583,N_17936);
xor U19407 (N_19407,N_16397,N_17434);
nand U19408 (N_19408,N_16814,N_16480);
nor U19409 (N_19409,N_17565,N_17220);
nor U19410 (N_19410,N_17458,N_16822);
or U19411 (N_19411,N_17621,N_16084);
and U19412 (N_19412,N_17792,N_16588);
nor U19413 (N_19413,N_17254,N_17383);
nor U19414 (N_19414,N_17647,N_17680);
xor U19415 (N_19415,N_17534,N_16787);
nand U19416 (N_19416,N_17694,N_16264);
nand U19417 (N_19417,N_16098,N_16212);
nor U19418 (N_19418,N_16968,N_17890);
nor U19419 (N_19419,N_17890,N_16080);
nand U19420 (N_19420,N_17282,N_17601);
nand U19421 (N_19421,N_16634,N_17431);
nand U19422 (N_19422,N_17740,N_17554);
or U19423 (N_19423,N_17717,N_17714);
and U19424 (N_19424,N_17004,N_16488);
nor U19425 (N_19425,N_17822,N_17767);
nand U19426 (N_19426,N_17145,N_16676);
nor U19427 (N_19427,N_17961,N_17635);
nand U19428 (N_19428,N_17779,N_17955);
nor U19429 (N_19429,N_16689,N_16358);
or U19430 (N_19430,N_16115,N_17629);
or U19431 (N_19431,N_16872,N_16438);
xnor U19432 (N_19432,N_17922,N_17277);
nand U19433 (N_19433,N_16952,N_16132);
and U19434 (N_19434,N_16364,N_16725);
nand U19435 (N_19435,N_17251,N_17088);
or U19436 (N_19436,N_17950,N_17164);
or U19437 (N_19437,N_17188,N_17391);
and U19438 (N_19438,N_17352,N_16812);
nor U19439 (N_19439,N_16407,N_16486);
and U19440 (N_19440,N_16060,N_17805);
or U19441 (N_19441,N_16775,N_16334);
or U19442 (N_19442,N_17817,N_17820);
and U19443 (N_19443,N_16442,N_17449);
xor U19444 (N_19444,N_17139,N_17382);
and U19445 (N_19445,N_16832,N_17802);
or U19446 (N_19446,N_17182,N_16653);
and U19447 (N_19447,N_16529,N_16939);
xnor U19448 (N_19448,N_17514,N_16781);
or U19449 (N_19449,N_16272,N_16642);
nand U19450 (N_19450,N_17354,N_16736);
nor U19451 (N_19451,N_16854,N_16235);
or U19452 (N_19452,N_16864,N_16574);
nor U19453 (N_19453,N_16514,N_16384);
nor U19454 (N_19454,N_17200,N_16162);
nand U19455 (N_19455,N_16327,N_16090);
or U19456 (N_19456,N_17930,N_16751);
or U19457 (N_19457,N_17247,N_16097);
nand U19458 (N_19458,N_16735,N_16099);
and U19459 (N_19459,N_16254,N_16390);
or U19460 (N_19460,N_17610,N_16218);
nand U19461 (N_19461,N_16622,N_17370);
nand U19462 (N_19462,N_16083,N_16904);
nand U19463 (N_19463,N_16887,N_16029);
nand U19464 (N_19464,N_17502,N_17906);
and U19465 (N_19465,N_16065,N_16001);
or U19466 (N_19466,N_17280,N_17074);
and U19467 (N_19467,N_17302,N_16675);
nand U19468 (N_19468,N_17972,N_16180);
and U19469 (N_19469,N_17544,N_16980);
nor U19470 (N_19470,N_16832,N_16479);
or U19471 (N_19471,N_17561,N_16801);
and U19472 (N_19472,N_16767,N_16492);
or U19473 (N_19473,N_17637,N_16617);
nor U19474 (N_19474,N_17672,N_17112);
nand U19475 (N_19475,N_17824,N_16016);
nor U19476 (N_19476,N_16540,N_17641);
nand U19477 (N_19477,N_16432,N_16089);
and U19478 (N_19478,N_17567,N_17533);
or U19479 (N_19479,N_16463,N_16889);
nor U19480 (N_19480,N_17155,N_16758);
or U19481 (N_19481,N_16736,N_17633);
and U19482 (N_19482,N_16207,N_17364);
and U19483 (N_19483,N_17684,N_16722);
nor U19484 (N_19484,N_17685,N_17331);
or U19485 (N_19485,N_17259,N_17302);
and U19486 (N_19486,N_17892,N_17895);
and U19487 (N_19487,N_16953,N_17540);
and U19488 (N_19488,N_17849,N_16027);
xor U19489 (N_19489,N_16960,N_16911);
nor U19490 (N_19490,N_17733,N_16961);
nand U19491 (N_19491,N_16861,N_16768);
nand U19492 (N_19492,N_17441,N_17183);
nor U19493 (N_19493,N_17856,N_17237);
nand U19494 (N_19494,N_17874,N_17906);
nor U19495 (N_19495,N_17071,N_17099);
and U19496 (N_19496,N_17546,N_17550);
or U19497 (N_19497,N_17620,N_16932);
and U19498 (N_19498,N_17792,N_16394);
nand U19499 (N_19499,N_16819,N_16673);
nand U19500 (N_19500,N_17236,N_17813);
nor U19501 (N_19501,N_16360,N_16249);
and U19502 (N_19502,N_16096,N_17807);
or U19503 (N_19503,N_16699,N_17301);
and U19504 (N_19504,N_16209,N_17882);
nand U19505 (N_19505,N_17730,N_16055);
and U19506 (N_19506,N_16105,N_17771);
and U19507 (N_19507,N_17263,N_17368);
and U19508 (N_19508,N_16741,N_16282);
and U19509 (N_19509,N_16676,N_16024);
and U19510 (N_19510,N_17546,N_16141);
and U19511 (N_19511,N_17539,N_17570);
and U19512 (N_19512,N_17105,N_16867);
and U19513 (N_19513,N_16742,N_17636);
nor U19514 (N_19514,N_16432,N_16078);
xnor U19515 (N_19515,N_17214,N_17532);
and U19516 (N_19516,N_16989,N_17211);
nor U19517 (N_19517,N_16914,N_17792);
nor U19518 (N_19518,N_16718,N_16562);
nor U19519 (N_19519,N_17923,N_17702);
or U19520 (N_19520,N_16346,N_16947);
and U19521 (N_19521,N_16342,N_16280);
or U19522 (N_19522,N_17561,N_17264);
nand U19523 (N_19523,N_17173,N_16768);
and U19524 (N_19524,N_17143,N_16589);
and U19525 (N_19525,N_16759,N_16096);
nand U19526 (N_19526,N_17564,N_16825);
and U19527 (N_19527,N_16140,N_16253);
nand U19528 (N_19528,N_16656,N_17483);
or U19529 (N_19529,N_16864,N_16368);
and U19530 (N_19530,N_16365,N_16361);
nand U19531 (N_19531,N_17339,N_17195);
nor U19532 (N_19532,N_17878,N_17609);
xnor U19533 (N_19533,N_17857,N_17272);
or U19534 (N_19534,N_16218,N_16029);
nor U19535 (N_19535,N_16813,N_17206);
nor U19536 (N_19536,N_17658,N_16324);
or U19537 (N_19537,N_16961,N_16316);
xor U19538 (N_19538,N_17456,N_17689);
or U19539 (N_19539,N_16432,N_16806);
and U19540 (N_19540,N_16609,N_17105);
nor U19541 (N_19541,N_16771,N_16067);
nor U19542 (N_19542,N_17915,N_17783);
and U19543 (N_19543,N_16972,N_17876);
and U19544 (N_19544,N_16277,N_16516);
and U19545 (N_19545,N_16116,N_17585);
or U19546 (N_19546,N_16650,N_17522);
nor U19547 (N_19547,N_16611,N_16484);
nand U19548 (N_19548,N_16665,N_17061);
nand U19549 (N_19549,N_17058,N_17932);
or U19550 (N_19550,N_16460,N_16365);
xnor U19551 (N_19551,N_17957,N_17150);
nand U19552 (N_19552,N_16770,N_16761);
nand U19553 (N_19553,N_17708,N_17207);
nor U19554 (N_19554,N_17464,N_17722);
nor U19555 (N_19555,N_16158,N_16387);
nor U19556 (N_19556,N_16024,N_17782);
nor U19557 (N_19557,N_16023,N_17606);
and U19558 (N_19558,N_16192,N_16555);
or U19559 (N_19559,N_16317,N_16669);
or U19560 (N_19560,N_16198,N_17979);
or U19561 (N_19561,N_16216,N_17573);
and U19562 (N_19562,N_17313,N_16523);
and U19563 (N_19563,N_17652,N_16028);
or U19564 (N_19564,N_17897,N_17291);
and U19565 (N_19565,N_17439,N_16703);
nor U19566 (N_19566,N_17888,N_17181);
and U19567 (N_19567,N_16252,N_17845);
nor U19568 (N_19568,N_17862,N_17293);
or U19569 (N_19569,N_16338,N_17964);
xor U19570 (N_19570,N_17326,N_17318);
nor U19571 (N_19571,N_16495,N_17622);
xnor U19572 (N_19572,N_17071,N_17470);
and U19573 (N_19573,N_16633,N_16266);
nand U19574 (N_19574,N_16486,N_17656);
nand U19575 (N_19575,N_16355,N_16310);
nand U19576 (N_19576,N_16422,N_17613);
nand U19577 (N_19577,N_16815,N_16693);
nand U19578 (N_19578,N_17949,N_16929);
nor U19579 (N_19579,N_16558,N_17588);
and U19580 (N_19580,N_17929,N_16821);
nand U19581 (N_19581,N_16003,N_16311);
and U19582 (N_19582,N_16604,N_17957);
nor U19583 (N_19583,N_17150,N_17037);
or U19584 (N_19584,N_16345,N_17866);
xnor U19585 (N_19585,N_17696,N_17353);
nor U19586 (N_19586,N_16066,N_17988);
nand U19587 (N_19587,N_16384,N_16346);
nand U19588 (N_19588,N_16526,N_16428);
nor U19589 (N_19589,N_16516,N_17567);
nand U19590 (N_19590,N_16755,N_16465);
or U19591 (N_19591,N_16205,N_16273);
xnor U19592 (N_19592,N_16755,N_16470);
nor U19593 (N_19593,N_16977,N_17568);
nor U19594 (N_19594,N_16732,N_16906);
or U19595 (N_19595,N_17067,N_17945);
or U19596 (N_19596,N_16710,N_16302);
xnor U19597 (N_19597,N_16721,N_17172);
and U19598 (N_19598,N_17995,N_16941);
or U19599 (N_19599,N_16795,N_17171);
or U19600 (N_19600,N_16501,N_16095);
or U19601 (N_19601,N_16626,N_17326);
or U19602 (N_19602,N_17516,N_17860);
nor U19603 (N_19603,N_17221,N_17812);
and U19604 (N_19604,N_16023,N_16490);
or U19605 (N_19605,N_17686,N_17648);
and U19606 (N_19606,N_16419,N_17203);
and U19607 (N_19607,N_17615,N_16150);
or U19608 (N_19608,N_17760,N_17214);
nor U19609 (N_19609,N_17288,N_16976);
and U19610 (N_19610,N_17984,N_17660);
nor U19611 (N_19611,N_17713,N_16091);
nand U19612 (N_19612,N_16596,N_17969);
and U19613 (N_19613,N_16879,N_17073);
and U19614 (N_19614,N_16779,N_16073);
or U19615 (N_19615,N_16114,N_17745);
and U19616 (N_19616,N_16622,N_16706);
or U19617 (N_19617,N_16680,N_16768);
and U19618 (N_19618,N_17371,N_17576);
or U19619 (N_19619,N_16826,N_17101);
or U19620 (N_19620,N_16201,N_16916);
or U19621 (N_19621,N_17650,N_16583);
and U19622 (N_19622,N_16904,N_17640);
nand U19623 (N_19623,N_17686,N_17861);
or U19624 (N_19624,N_16269,N_16277);
and U19625 (N_19625,N_17868,N_17963);
or U19626 (N_19626,N_17269,N_17801);
or U19627 (N_19627,N_17107,N_17637);
or U19628 (N_19628,N_17881,N_17972);
or U19629 (N_19629,N_17980,N_17757);
xor U19630 (N_19630,N_17444,N_16571);
nand U19631 (N_19631,N_16831,N_17672);
nor U19632 (N_19632,N_16501,N_16938);
nand U19633 (N_19633,N_16370,N_17259);
and U19634 (N_19634,N_17011,N_16852);
nor U19635 (N_19635,N_17247,N_16088);
and U19636 (N_19636,N_16160,N_17706);
or U19637 (N_19637,N_17553,N_17902);
or U19638 (N_19638,N_17284,N_16550);
and U19639 (N_19639,N_17070,N_16874);
or U19640 (N_19640,N_16381,N_17667);
nor U19641 (N_19641,N_16160,N_16563);
nand U19642 (N_19642,N_17879,N_17697);
nor U19643 (N_19643,N_16184,N_17736);
xnor U19644 (N_19644,N_17302,N_17047);
xor U19645 (N_19645,N_17878,N_17646);
nand U19646 (N_19646,N_16478,N_16864);
and U19647 (N_19647,N_16205,N_17867);
or U19648 (N_19648,N_17339,N_17413);
or U19649 (N_19649,N_16638,N_16102);
nor U19650 (N_19650,N_16476,N_16834);
nor U19651 (N_19651,N_16806,N_17459);
nor U19652 (N_19652,N_16740,N_16910);
nor U19653 (N_19653,N_16887,N_16924);
nor U19654 (N_19654,N_16134,N_16178);
and U19655 (N_19655,N_16061,N_17697);
nor U19656 (N_19656,N_16786,N_16430);
nor U19657 (N_19657,N_16481,N_16772);
and U19658 (N_19658,N_16363,N_17476);
and U19659 (N_19659,N_16375,N_16228);
nor U19660 (N_19660,N_16040,N_16668);
nand U19661 (N_19661,N_16267,N_17904);
nand U19662 (N_19662,N_16822,N_16761);
and U19663 (N_19663,N_17140,N_16914);
nor U19664 (N_19664,N_17425,N_16328);
nand U19665 (N_19665,N_16601,N_16396);
nand U19666 (N_19666,N_16075,N_17583);
or U19667 (N_19667,N_17373,N_16798);
or U19668 (N_19668,N_16723,N_17003);
or U19669 (N_19669,N_16202,N_17066);
xor U19670 (N_19670,N_16070,N_17310);
or U19671 (N_19671,N_16973,N_16639);
or U19672 (N_19672,N_16015,N_16298);
nand U19673 (N_19673,N_17438,N_17281);
nand U19674 (N_19674,N_16344,N_16740);
nand U19675 (N_19675,N_16338,N_16353);
nand U19676 (N_19676,N_16114,N_16087);
xnor U19677 (N_19677,N_16485,N_17544);
and U19678 (N_19678,N_16085,N_16272);
or U19679 (N_19679,N_16931,N_16234);
nor U19680 (N_19680,N_16727,N_17467);
nand U19681 (N_19681,N_16599,N_17278);
nand U19682 (N_19682,N_17917,N_16444);
or U19683 (N_19683,N_17724,N_16202);
nand U19684 (N_19684,N_16946,N_16898);
or U19685 (N_19685,N_17317,N_16022);
nor U19686 (N_19686,N_16574,N_16196);
and U19687 (N_19687,N_17793,N_17183);
or U19688 (N_19688,N_17303,N_16882);
and U19689 (N_19689,N_16576,N_16469);
nand U19690 (N_19690,N_16511,N_17801);
nand U19691 (N_19691,N_16953,N_16059);
and U19692 (N_19692,N_17358,N_17128);
nand U19693 (N_19693,N_17709,N_16710);
or U19694 (N_19694,N_16616,N_16087);
nor U19695 (N_19695,N_16487,N_17918);
xor U19696 (N_19696,N_16801,N_16643);
nor U19697 (N_19697,N_16082,N_16636);
and U19698 (N_19698,N_17210,N_17002);
or U19699 (N_19699,N_17021,N_16884);
or U19700 (N_19700,N_17590,N_16546);
nand U19701 (N_19701,N_17033,N_16288);
xor U19702 (N_19702,N_17886,N_16654);
and U19703 (N_19703,N_17879,N_16845);
and U19704 (N_19704,N_17787,N_16877);
nor U19705 (N_19705,N_16526,N_17719);
nand U19706 (N_19706,N_17971,N_17458);
nand U19707 (N_19707,N_17135,N_16905);
nand U19708 (N_19708,N_16938,N_16283);
and U19709 (N_19709,N_16741,N_17007);
nand U19710 (N_19710,N_16511,N_17700);
and U19711 (N_19711,N_16504,N_17169);
nand U19712 (N_19712,N_17876,N_17497);
and U19713 (N_19713,N_17054,N_17679);
nor U19714 (N_19714,N_17653,N_17739);
xor U19715 (N_19715,N_16950,N_16290);
nor U19716 (N_19716,N_17596,N_17917);
nand U19717 (N_19717,N_16259,N_17043);
or U19718 (N_19718,N_16831,N_16133);
nand U19719 (N_19719,N_16286,N_17167);
nor U19720 (N_19720,N_17326,N_17598);
nor U19721 (N_19721,N_16616,N_17395);
nand U19722 (N_19722,N_16033,N_17554);
nor U19723 (N_19723,N_17590,N_17865);
nand U19724 (N_19724,N_17448,N_17780);
nor U19725 (N_19725,N_17010,N_17452);
nor U19726 (N_19726,N_17429,N_16677);
nor U19727 (N_19727,N_16141,N_17926);
xnor U19728 (N_19728,N_17943,N_17376);
and U19729 (N_19729,N_17077,N_16178);
or U19730 (N_19730,N_17889,N_16683);
nor U19731 (N_19731,N_17729,N_17946);
and U19732 (N_19732,N_16326,N_17610);
or U19733 (N_19733,N_17628,N_16464);
nand U19734 (N_19734,N_17731,N_16350);
or U19735 (N_19735,N_17604,N_16145);
and U19736 (N_19736,N_16342,N_16552);
and U19737 (N_19737,N_16165,N_17183);
nand U19738 (N_19738,N_16524,N_17109);
xnor U19739 (N_19739,N_17532,N_16624);
xor U19740 (N_19740,N_17029,N_17291);
nand U19741 (N_19741,N_17675,N_16093);
xor U19742 (N_19742,N_16288,N_17655);
or U19743 (N_19743,N_17348,N_17307);
or U19744 (N_19744,N_16081,N_16041);
nor U19745 (N_19745,N_17805,N_17355);
nand U19746 (N_19746,N_17355,N_17667);
or U19747 (N_19747,N_16425,N_16822);
and U19748 (N_19748,N_17177,N_17246);
or U19749 (N_19749,N_17099,N_17156);
nand U19750 (N_19750,N_16664,N_17861);
nor U19751 (N_19751,N_16376,N_16352);
or U19752 (N_19752,N_17611,N_16170);
nor U19753 (N_19753,N_16719,N_16154);
nor U19754 (N_19754,N_16692,N_16548);
or U19755 (N_19755,N_16421,N_16414);
nand U19756 (N_19756,N_16810,N_17785);
and U19757 (N_19757,N_16967,N_17361);
nand U19758 (N_19758,N_16834,N_16786);
nand U19759 (N_19759,N_17754,N_16296);
nor U19760 (N_19760,N_16825,N_16532);
and U19761 (N_19761,N_17006,N_16870);
or U19762 (N_19762,N_16505,N_17226);
or U19763 (N_19763,N_17778,N_16214);
or U19764 (N_19764,N_17734,N_16265);
nor U19765 (N_19765,N_17535,N_17452);
or U19766 (N_19766,N_17722,N_17443);
and U19767 (N_19767,N_17410,N_17843);
nor U19768 (N_19768,N_16419,N_16314);
nand U19769 (N_19769,N_17541,N_16274);
nand U19770 (N_19770,N_16442,N_17117);
nor U19771 (N_19771,N_16058,N_17204);
nand U19772 (N_19772,N_16020,N_17794);
nor U19773 (N_19773,N_16910,N_17314);
and U19774 (N_19774,N_17879,N_17430);
nor U19775 (N_19775,N_17704,N_16168);
nor U19776 (N_19776,N_17371,N_16092);
and U19777 (N_19777,N_17111,N_16551);
nor U19778 (N_19778,N_17433,N_16760);
and U19779 (N_19779,N_17615,N_17165);
xnor U19780 (N_19780,N_16468,N_16974);
or U19781 (N_19781,N_16365,N_16139);
or U19782 (N_19782,N_17250,N_16461);
or U19783 (N_19783,N_17389,N_17097);
nand U19784 (N_19784,N_17528,N_16563);
xnor U19785 (N_19785,N_17192,N_17597);
and U19786 (N_19786,N_17416,N_16305);
nor U19787 (N_19787,N_16588,N_16495);
or U19788 (N_19788,N_17058,N_16850);
nor U19789 (N_19789,N_16693,N_16153);
nor U19790 (N_19790,N_17462,N_17354);
nand U19791 (N_19791,N_16289,N_17142);
or U19792 (N_19792,N_16612,N_16349);
nand U19793 (N_19793,N_16807,N_16086);
and U19794 (N_19794,N_16456,N_16399);
nor U19795 (N_19795,N_17352,N_17005);
nor U19796 (N_19796,N_16541,N_17933);
nor U19797 (N_19797,N_16837,N_17661);
nor U19798 (N_19798,N_17412,N_17066);
nand U19799 (N_19799,N_16849,N_16821);
and U19800 (N_19800,N_16453,N_17323);
nand U19801 (N_19801,N_17539,N_16433);
nand U19802 (N_19802,N_17969,N_16669);
xor U19803 (N_19803,N_17548,N_16764);
nand U19804 (N_19804,N_17881,N_17527);
nor U19805 (N_19805,N_16385,N_17621);
nand U19806 (N_19806,N_16505,N_16921);
or U19807 (N_19807,N_17381,N_17017);
nand U19808 (N_19808,N_16380,N_16310);
nor U19809 (N_19809,N_17150,N_16599);
and U19810 (N_19810,N_17244,N_16970);
nor U19811 (N_19811,N_16697,N_17370);
nor U19812 (N_19812,N_16071,N_16984);
xnor U19813 (N_19813,N_16621,N_16393);
and U19814 (N_19814,N_16257,N_17744);
nand U19815 (N_19815,N_17233,N_16372);
nor U19816 (N_19816,N_17196,N_17298);
and U19817 (N_19817,N_17391,N_17215);
or U19818 (N_19818,N_16590,N_16676);
or U19819 (N_19819,N_17796,N_17874);
or U19820 (N_19820,N_17140,N_17176);
or U19821 (N_19821,N_17614,N_16354);
nor U19822 (N_19822,N_16030,N_16471);
nor U19823 (N_19823,N_17523,N_17965);
nand U19824 (N_19824,N_17660,N_17941);
xnor U19825 (N_19825,N_16382,N_17532);
or U19826 (N_19826,N_17458,N_16601);
nor U19827 (N_19827,N_17527,N_17496);
or U19828 (N_19828,N_17591,N_16142);
nand U19829 (N_19829,N_16614,N_16094);
nor U19830 (N_19830,N_16316,N_17336);
nor U19831 (N_19831,N_16240,N_17285);
xor U19832 (N_19832,N_16550,N_16964);
or U19833 (N_19833,N_16247,N_16731);
nand U19834 (N_19834,N_16702,N_16075);
nand U19835 (N_19835,N_16173,N_16446);
xnor U19836 (N_19836,N_17051,N_17269);
and U19837 (N_19837,N_17726,N_17435);
and U19838 (N_19838,N_16587,N_16881);
nor U19839 (N_19839,N_17043,N_16113);
nor U19840 (N_19840,N_16879,N_17417);
nor U19841 (N_19841,N_16139,N_17712);
and U19842 (N_19842,N_16534,N_17628);
or U19843 (N_19843,N_16180,N_17790);
or U19844 (N_19844,N_17928,N_16044);
nor U19845 (N_19845,N_17995,N_16866);
nor U19846 (N_19846,N_16600,N_17690);
nand U19847 (N_19847,N_17568,N_16809);
nor U19848 (N_19848,N_17461,N_17844);
xnor U19849 (N_19849,N_16287,N_16973);
and U19850 (N_19850,N_17100,N_16324);
nor U19851 (N_19851,N_16112,N_16862);
and U19852 (N_19852,N_17566,N_17666);
and U19853 (N_19853,N_16943,N_17089);
xnor U19854 (N_19854,N_17425,N_16972);
nand U19855 (N_19855,N_17623,N_16118);
and U19856 (N_19856,N_17812,N_17526);
nor U19857 (N_19857,N_17460,N_17713);
nor U19858 (N_19858,N_17417,N_17030);
nand U19859 (N_19859,N_17011,N_16674);
and U19860 (N_19860,N_16314,N_17962);
nor U19861 (N_19861,N_17930,N_16925);
nand U19862 (N_19862,N_16457,N_17172);
or U19863 (N_19863,N_17771,N_17756);
and U19864 (N_19864,N_17243,N_17285);
xnor U19865 (N_19865,N_17949,N_16958);
and U19866 (N_19866,N_17878,N_17268);
nand U19867 (N_19867,N_17881,N_17570);
and U19868 (N_19868,N_17032,N_17981);
or U19869 (N_19869,N_16576,N_16892);
xor U19870 (N_19870,N_16020,N_16265);
and U19871 (N_19871,N_17483,N_16086);
and U19872 (N_19872,N_16673,N_16490);
and U19873 (N_19873,N_16243,N_17228);
nor U19874 (N_19874,N_16285,N_17820);
nand U19875 (N_19875,N_17996,N_16901);
xnor U19876 (N_19876,N_16554,N_17386);
and U19877 (N_19877,N_17840,N_16979);
or U19878 (N_19878,N_17771,N_16545);
nor U19879 (N_19879,N_16381,N_16138);
nor U19880 (N_19880,N_17691,N_16156);
nand U19881 (N_19881,N_17756,N_17538);
nor U19882 (N_19882,N_17212,N_16794);
and U19883 (N_19883,N_16117,N_17353);
xnor U19884 (N_19884,N_16162,N_16819);
nand U19885 (N_19885,N_16679,N_16640);
nand U19886 (N_19886,N_17704,N_17660);
nand U19887 (N_19887,N_16441,N_16210);
nand U19888 (N_19888,N_17930,N_17297);
nor U19889 (N_19889,N_17066,N_16195);
or U19890 (N_19890,N_16729,N_17639);
or U19891 (N_19891,N_16346,N_16032);
or U19892 (N_19892,N_17935,N_16007);
nor U19893 (N_19893,N_17616,N_16353);
or U19894 (N_19894,N_16780,N_16829);
nor U19895 (N_19895,N_17828,N_17883);
or U19896 (N_19896,N_16119,N_16939);
and U19897 (N_19897,N_16876,N_17217);
nand U19898 (N_19898,N_16923,N_17305);
nor U19899 (N_19899,N_17866,N_16201);
nand U19900 (N_19900,N_16516,N_17880);
and U19901 (N_19901,N_16304,N_16425);
nand U19902 (N_19902,N_16962,N_17877);
nor U19903 (N_19903,N_17067,N_16548);
nand U19904 (N_19904,N_16109,N_17546);
and U19905 (N_19905,N_16626,N_17542);
nand U19906 (N_19906,N_17069,N_16637);
nand U19907 (N_19907,N_17121,N_17873);
nand U19908 (N_19908,N_16030,N_17867);
and U19909 (N_19909,N_16174,N_17140);
nand U19910 (N_19910,N_17328,N_16540);
nand U19911 (N_19911,N_17383,N_17734);
nor U19912 (N_19912,N_16644,N_16502);
nor U19913 (N_19913,N_16630,N_16171);
nand U19914 (N_19914,N_17603,N_17066);
or U19915 (N_19915,N_16836,N_16359);
or U19916 (N_19916,N_16319,N_16980);
or U19917 (N_19917,N_16841,N_17145);
nor U19918 (N_19918,N_17989,N_17520);
nor U19919 (N_19919,N_17750,N_17297);
nand U19920 (N_19920,N_16834,N_16317);
nand U19921 (N_19921,N_17711,N_16902);
and U19922 (N_19922,N_17734,N_16716);
and U19923 (N_19923,N_17732,N_16720);
nor U19924 (N_19924,N_17090,N_16739);
xnor U19925 (N_19925,N_16206,N_16377);
nand U19926 (N_19926,N_16023,N_17951);
nor U19927 (N_19927,N_17633,N_17298);
nand U19928 (N_19928,N_17913,N_17698);
nor U19929 (N_19929,N_16110,N_16076);
nand U19930 (N_19930,N_17517,N_16688);
nand U19931 (N_19931,N_16011,N_16170);
nand U19932 (N_19932,N_16396,N_17029);
and U19933 (N_19933,N_17489,N_17101);
nor U19934 (N_19934,N_17061,N_17969);
xor U19935 (N_19935,N_17392,N_16699);
xnor U19936 (N_19936,N_17984,N_16586);
or U19937 (N_19937,N_17714,N_16502);
xnor U19938 (N_19938,N_17884,N_16971);
nand U19939 (N_19939,N_17133,N_16105);
or U19940 (N_19940,N_16593,N_17567);
xnor U19941 (N_19941,N_17211,N_16639);
or U19942 (N_19942,N_17212,N_16763);
nor U19943 (N_19943,N_17094,N_17605);
nor U19944 (N_19944,N_17065,N_17668);
or U19945 (N_19945,N_16186,N_16902);
or U19946 (N_19946,N_16593,N_16548);
and U19947 (N_19947,N_17612,N_17715);
xnor U19948 (N_19948,N_16963,N_16891);
and U19949 (N_19949,N_17030,N_16883);
xor U19950 (N_19950,N_16718,N_16015);
and U19951 (N_19951,N_17806,N_16497);
or U19952 (N_19952,N_16398,N_16368);
nand U19953 (N_19953,N_17699,N_16533);
nor U19954 (N_19954,N_17089,N_16041);
and U19955 (N_19955,N_16018,N_16645);
nor U19956 (N_19956,N_16581,N_17363);
nor U19957 (N_19957,N_16414,N_17417);
or U19958 (N_19958,N_16156,N_17202);
nand U19959 (N_19959,N_17245,N_16123);
nor U19960 (N_19960,N_17189,N_17392);
or U19961 (N_19961,N_16219,N_16132);
nand U19962 (N_19962,N_16218,N_16589);
nor U19963 (N_19963,N_16167,N_16590);
and U19964 (N_19964,N_16561,N_17397);
nor U19965 (N_19965,N_16704,N_17673);
nand U19966 (N_19966,N_17127,N_16399);
xor U19967 (N_19967,N_17956,N_17180);
or U19968 (N_19968,N_16425,N_17039);
nor U19969 (N_19969,N_17231,N_17546);
or U19970 (N_19970,N_16271,N_16883);
or U19971 (N_19971,N_16141,N_17894);
or U19972 (N_19972,N_16815,N_16275);
nor U19973 (N_19973,N_17843,N_16213);
and U19974 (N_19974,N_17840,N_16036);
or U19975 (N_19975,N_17996,N_16774);
nor U19976 (N_19976,N_16503,N_16434);
nand U19977 (N_19977,N_17657,N_16512);
nand U19978 (N_19978,N_17553,N_16543);
and U19979 (N_19979,N_16650,N_17879);
or U19980 (N_19980,N_17333,N_17588);
nand U19981 (N_19981,N_17131,N_16948);
or U19982 (N_19982,N_16502,N_17396);
and U19983 (N_19983,N_16189,N_17910);
nand U19984 (N_19984,N_17934,N_17869);
xor U19985 (N_19985,N_16962,N_17613);
nand U19986 (N_19986,N_16510,N_16581);
or U19987 (N_19987,N_17262,N_16712);
nand U19988 (N_19988,N_17042,N_16607);
and U19989 (N_19989,N_17869,N_16601);
or U19990 (N_19990,N_17364,N_16040);
and U19991 (N_19991,N_16911,N_17131);
or U19992 (N_19992,N_17497,N_17227);
or U19993 (N_19993,N_16398,N_16921);
or U19994 (N_19994,N_16770,N_16483);
xnor U19995 (N_19995,N_17124,N_16167);
or U19996 (N_19996,N_17323,N_16194);
nor U19997 (N_19997,N_16170,N_16405);
and U19998 (N_19998,N_16545,N_17616);
nor U19999 (N_19999,N_16801,N_17982);
nand UO_0 (O_0,N_18990,N_18534);
nand UO_1 (O_1,N_19620,N_19907);
or UO_2 (O_2,N_19989,N_18513);
xnor UO_3 (O_3,N_18321,N_18351);
and UO_4 (O_4,N_18674,N_19468);
and UO_5 (O_5,N_18000,N_19806);
xor UO_6 (O_6,N_18655,N_18396);
nor UO_7 (O_7,N_18066,N_19978);
and UO_8 (O_8,N_19729,N_19628);
nand UO_9 (O_9,N_19476,N_18353);
nor UO_10 (O_10,N_19138,N_18656);
or UO_11 (O_11,N_18085,N_19260);
or UO_12 (O_12,N_18070,N_19642);
or UO_13 (O_13,N_19245,N_19947);
nor UO_14 (O_14,N_18912,N_18336);
and UO_15 (O_15,N_18958,N_18339);
or UO_16 (O_16,N_18617,N_18436);
nor UO_17 (O_17,N_18419,N_18376);
or UO_18 (O_18,N_18448,N_19125);
nor UO_19 (O_19,N_18140,N_18638);
nand UO_20 (O_20,N_19095,N_19536);
and UO_21 (O_21,N_18544,N_19890);
and UO_22 (O_22,N_19933,N_18897);
nand UO_23 (O_23,N_19054,N_18112);
xor UO_24 (O_24,N_18155,N_19117);
and UO_25 (O_25,N_18610,N_18464);
or UO_26 (O_26,N_19851,N_19188);
and UO_27 (O_27,N_18168,N_18802);
xor UO_28 (O_28,N_19588,N_19661);
and UO_29 (O_29,N_19964,N_19398);
nor UO_30 (O_30,N_18987,N_19387);
nor UO_31 (O_31,N_19747,N_19562);
nor UO_32 (O_32,N_18695,N_19896);
nand UO_33 (O_33,N_18154,N_18174);
and UO_34 (O_34,N_18394,N_18426);
and UO_35 (O_35,N_18265,N_18182);
or UO_36 (O_36,N_19845,N_19945);
and UO_37 (O_37,N_19208,N_18184);
nor UO_38 (O_38,N_18312,N_19505);
and UO_39 (O_39,N_18226,N_18496);
nand UO_40 (O_40,N_19233,N_19999);
nor UO_41 (O_41,N_19785,N_19883);
or UO_42 (O_42,N_19289,N_19370);
and UO_43 (O_43,N_19241,N_19464);
or UO_44 (O_44,N_19650,N_18243);
and UO_45 (O_45,N_18531,N_19832);
nand UO_46 (O_46,N_18960,N_18091);
and UO_47 (O_47,N_19328,N_18849);
and UO_48 (O_48,N_19744,N_19919);
nor UO_49 (O_49,N_19728,N_18388);
nand UO_50 (O_50,N_18803,N_18716);
or UO_51 (O_51,N_19962,N_18625);
xor UO_52 (O_52,N_18221,N_18129);
and UO_53 (O_53,N_18751,N_19878);
nand UO_54 (O_54,N_18056,N_19093);
or UO_55 (O_55,N_19110,N_19101);
nand UO_56 (O_56,N_19762,N_18955);
nand UO_57 (O_57,N_18765,N_19655);
or UO_58 (O_58,N_18600,N_19251);
xnor UO_59 (O_59,N_18220,N_18555);
or UO_60 (O_60,N_19614,N_19686);
or UO_61 (O_61,N_18564,N_19580);
nand UO_62 (O_62,N_18694,N_18477);
xor UO_63 (O_63,N_18144,N_19960);
and UO_64 (O_64,N_19705,N_19771);
and UO_65 (O_65,N_18314,N_18398);
and UO_66 (O_66,N_19910,N_19394);
nor UO_67 (O_67,N_18292,N_19106);
or UO_68 (O_68,N_19200,N_18186);
or UO_69 (O_69,N_19731,N_19234);
nor UO_70 (O_70,N_19203,N_19593);
nand UO_71 (O_71,N_18627,N_18896);
and UO_72 (O_72,N_19629,N_19915);
nand UO_73 (O_73,N_18532,N_19291);
and UO_74 (O_74,N_18787,N_19697);
nor UO_75 (O_75,N_19146,N_19649);
xnor UO_76 (O_76,N_18658,N_19176);
nor UO_77 (O_77,N_19267,N_19918);
or UO_78 (O_78,N_19459,N_19209);
or UO_79 (O_79,N_19455,N_18171);
nor UO_80 (O_80,N_18246,N_19175);
or UO_81 (O_81,N_19134,N_18445);
xor UO_82 (O_82,N_18961,N_19560);
and UO_83 (O_83,N_18365,N_19607);
or UO_84 (O_84,N_19952,N_18846);
xor UO_85 (O_85,N_19699,N_18263);
and UO_86 (O_86,N_18789,N_19058);
nor UO_87 (O_87,N_18392,N_18071);
and UO_88 (O_88,N_18428,N_18300);
xnor UO_89 (O_89,N_19740,N_19040);
or UO_90 (O_90,N_19339,N_19774);
nor UO_91 (O_91,N_19271,N_18516);
or UO_92 (O_92,N_19862,N_18784);
and UO_93 (O_93,N_19107,N_18796);
and UO_94 (O_94,N_19128,N_19715);
nand UO_95 (O_95,N_19645,N_18476);
nor UO_96 (O_96,N_19198,N_18950);
nor UO_97 (O_97,N_19658,N_18211);
nor UO_98 (O_98,N_19957,N_19470);
xnor UO_99 (O_99,N_19707,N_19244);
and UO_100 (O_100,N_19948,N_19124);
and UO_101 (O_101,N_19524,N_19376);
nand UO_102 (O_102,N_19502,N_19078);
and UO_103 (O_103,N_18239,N_19207);
nor UO_104 (O_104,N_19534,N_18889);
nand UO_105 (O_105,N_19154,N_19369);
and UO_106 (O_106,N_19453,N_18382);
or UO_107 (O_107,N_19055,N_19503);
nand UO_108 (O_108,N_18947,N_18838);
nand UO_109 (O_109,N_19222,N_18370);
or UO_110 (O_110,N_19804,N_18812);
xor UO_111 (O_111,N_19392,N_18387);
or UO_112 (O_112,N_19386,N_18390);
and UO_113 (O_113,N_19533,N_18008);
nand UO_114 (O_114,N_18311,N_19908);
and UO_115 (O_115,N_18984,N_18668);
nand UO_116 (O_116,N_18180,N_19229);
nand UO_117 (O_117,N_18165,N_19623);
nand UO_118 (O_118,N_19640,N_19263);
or UO_119 (O_119,N_18736,N_19850);
xor UO_120 (O_120,N_18420,N_18946);
or UO_121 (O_121,N_19954,N_18639);
nor UO_122 (O_122,N_18726,N_19827);
nor UO_123 (O_123,N_18910,N_18703);
nor UO_124 (O_124,N_19600,N_18842);
nor UO_125 (O_125,N_19252,N_18623);
or UO_126 (O_126,N_18994,N_19424);
nand UO_127 (O_127,N_19433,N_19777);
nor UO_128 (O_128,N_18528,N_18741);
nand UO_129 (O_129,N_19706,N_18356);
nand UO_130 (O_130,N_18636,N_18414);
xnor UO_131 (O_131,N_19246,N_19282);
nand UO_132 (O_132,N_18179,N_18911);
nand UO_133 (O_133,N_18457,N_18223);
or UO_134 (O_134,N_19020,N_18233);
or UO_135 (O_135,N_19683,N_19480);
and UO_136 (O_136,N_19381,N_18641);
nand UO_137 (O_137,N_18764,N_18041);
nand UO_138 (O_138,N_18898,N_19326);
and UO_139 (O_139,N_18925,N_18815);
nand UO_140 (O_140,N_18722,N_18199);
or UO_141 (O_141,N_18702,N_18409);
or UO_142 (O_142,N_19063,N_19323);
and UO_143 (O_143,N_19135,N_18735);
and UO_144 (O_144,N_19047,N_19546);
nor UO_145 (O_145,N_19216,N_19321);
and UO_146 (O_146,N_18498,N_18432);
and UO_147 (O_147,N_19105,N_19288);
xnor UO_148 (O_148,N_19692,N_18196);
and UO_149 (O_149,N_19936,N_18685);
or UO_150 (O_150,N_19928,N_19319);
and UO_151 (O_151,N_18714,N_18197);
and UO_152 (O_152,N_19094,N_19912);
or UO_153 (O_153,N_19894,N_18433);
and UO_154 (O_154,N_19859,N_18093);
nor UO_155 (O_155,N_18575,N_19284);
nand UO_156 (O_156,N_18616,N_18704);
or UO_157 (O_157,N_19172,N_18101);
nor UO_158 (O_158,N_18999,N_18319);
or UO_159 (O_159,N_18021,N_18074);
nor UO_160 (O_160,N_18135,N_18385);
and UO_161 (O_161,N_19494,N_18378);
and UO_162 (O_162,N_18176,N_19287);
xnor UO_163 (O_163,N_19577,N_18201);
xnor UO_164 (O_164,N_18829,N_19713);
nor UO_165 (O_165,N_18595,N_19190);
nor UO_166 (O_166,N_19052,N_19021);
or UO_167 (O_167,N_18153,N_19364);
and UO_168 (O_168,N_18208,N_19102);
nor UO_169 (O_169,N_18111,N_18285);
nand UO_170 (O_170,N_19196,N_19192);
and UO_171 (O_171,N_18443,N_19709);
nand UO_172 (O_172,N_19872,N_18416);
or UO_173 (O_173,N_19255,N_19738);
nor UO_174 (O_174,N_19438,N_19512);
or UO_175 (O_175,N_18523,N_18017);
nand UO_176 (O_176,N_19286,N_19174);
nand UO_177 (O_177,N_18137,N_19171);
nor UO_178 (O_178,N_19905,N_18866);
and UO_179 (O_179,N_18650,N_18767);
or UO_180 (O_180,N_19025,N_18497);
nor UO_181 (O_181,N_19653,N_19368);
and UO_182 (O_182,N_18412,N_18522);
nor UO_183 (O_183,N_19545,N_18280);
nand UO_184 (O_184,N_18320,N_19404);
and UO_185 (O_185,N_18380,N_18649);
or UO_186 (O_186,N_19811,N_18247);
or UO_187 (O_187,N_18423,N_19017);
nor UO_188 (O_188,N_19210,N_18257);
xnor UO_189 (O_189,N_18537,N_19903);
xor UO_190 (O_190,N_19922,N_19079);
nand UO_191 (O_191,N_19719,N_18482);
nand UO_192 (O_192,N_19589,N_19002);
and UO_193 (O_193,N_19920,N_18205);
and UO_194 (O_194,N_19767,N_19247);
xor UO_195 (O_195,N_18928,N_18559);
nand UO_196 (O_196,N_18922,N_18556);
and UO_197 (O_197,N_18222,N_19576);
or UO_198 (O_198,N_19344,N_18809);
nand UO_199 (O_199,N_19264,N_19089);
nand UO_200 (O_200,N_19179,N_19592);
and UO_201 (O_201,N_19735,N_19197);
nor UO_202 (O_202,N_19914,N_19349);
or UO_203 (O_203,N_19882,N_19754);
and UO_204 (O_204,N_18132,N_18774);
or UO_205 (O_205,N_18373,N_18269);
or UO_206 (O_206,N_19467,N_18102);
xor UO_207 (O_207,N_18980,N_19566);
nand UO_208 (O_208,N_18206,N_19250);
nand UO_209 (O_209,N_18647,N_18402);
or UO_210 (O_210,N_18957,N_19460);
nor UO_211 (O_211,N_19547,N_18012);
nand UO_212 (O_212,N_18274,N_18484);
or UO_213 (O_213,N_19803,N_19334);
nand UO_214 (O_214,N_18622,N_19924);
xnor UO_215 (O_215,N_18368,N_19969);
nor UO_216 (O_216,N_18614,N_18675);
nand UO_217 (O_217,N_19848,N_19057);
and UO_218 (O_218,N_18948,N_19902);
xor UO_219 (O_219,N_18040,N_18251);
nand UO_220 (O_220,N_19342,N_19985);
nor UO_221 (O_221,N_19432,N_18806);
or UO_222 (O_222,N_19929,N_18976);
nand UO_223 (O_223,N_19029,N_19232);
and UO_224 (O_224,N_19316,N_19236);
nand UO_225 (O_225,N_19722,N_19988);
nand UO_226 (O_226,N_19443,N_18400);
or UO_227 (O_227,N_19998,N_19330);
nor UO_228 (O_228,N_19013,N_18893);
or UO_229 (O_229,N_18903,N_19130);
nor UO_230 (O_230,N_19516,N_18565);
and UO_231 (O_231,N_19809,N_19582);
or UO_232 (O_232,N_18539,N_18217);
and UO_233 (O_233,N_18177,N_19164);
or UO_234 (O_234,N_19431,N_18367);
xor UO_235 (O_235,N_19761,N_19698);
nand UO_236 (O_236,N_18830,N_18969);
or UO_237 (O_237,N_19290,N_19519);
and UO_238 (O_238,N_18526,N_19955);
or UO_239 (O_239,N_19590,N_19075);
xor UO_240 (O_240,N_19652,N_18277);
xor UO_241 (O_241,N_19363,N_19294);
nor UO_242 (O_242,N_18700,N_19568);
nand UO_243 (O_243,N_18613,N_19412);
and UO_244 (O_244,N_19836,N_19755);
nand UO_245 (O_245,N_18250,N_18527);
and UO_246 (O_246,N_19940,N_18634);
nand UO_247 (O_247,N_18086,N_19726);
xnor UO_248 (O_248,N_19753,N_19569);
nand UO_249 (O_249,N_19454,N_19579);
nand UO_250 (O_250,N_19508,N_18372);
or UO_251 (O_251,N_19926,N_19925);
xor UO_252 (O_252,N_18779,N_18082);
or UO_253 (O_253,N_18921,N_18363);
nand UO_254 (O_254,N_19700,N_19001);
and UO_255 (O_255,N_18288,N_18282);
and UO_256 (O_256,N_18752,N_19157);
and UO_257 (O_257,N_18275,N_18072);
and UO_258 (O_258,N_18002,N_18146);
nand UO_259 (O_259,N_19621,N_19169);
and UO_260 (O_260,N_19227,N_19921);
nand UO_261 (O_261,N_19975,N_19701);
xnor UO_262 (O_262,N_19854,N_19829);
or UO_263 (O_263,N_19830,N_19420);
and UO_264 (O_264,N_18192,N_18869);
nand UO_265 (O_265,N_19504,N_19356);
nand UO_266 (O_266,N_18972,N_18608);
and UO_267 (O_267,N_19156,N_18490);
xor UO_268 (O_268,N_19279,N_18589);
xnor UO_269 (O_269,N_18261,N_18081);
nand UO_270 (O_270,N_19606,N_19783);
xnor UO_271 (O_271,N_19009,N_19423);
xnor UO_272 (O_272,N_19441,N_18709);
nand UO_273 (O_273,N_19211,N_18032);
nor UO_274 (O_274,N_18511,N_18507);
and UO_275 (O_275,N_19817,N_19496);
or UO_276 (O_276,N_19951,N_18895);
and UO_277 (O_277,N_18771,N_18410);
and UO_278 (O_278,N_18548,N_18749);
nand UO_279 (O_279,N_18579,N_18064);
or UO_280 (O_280,N_19177,N_18856);
nand UO_281 (O_281,N_19765,N_19053);
and UO_282 (O_282,N_18262,N_18268);
nor UO_283 (O_283,N_19307,N_19627);
nand UO_284 (O_284,N_18149,N_18831);
nor UO_285 (O_285,N_18106,N_19388);
nor UO_286 (O_286,N_19067,N_19973);
and UO_287 (O_287,N_19361,N_19449);
nand UO_288 (O_288,N_19535,N_18238);
nand UO_289 (O_289,N_19796,N_19165);
nand UO_290 (O_290,N_18393,N_18533);
and UO_291 (O_291,N_19343,N_18989);
or UO_292 (O_292,N_19314,N_19204);
or UO_293 (O_293,N_18494,N_19133);
nand UO_294 (O_294,N_19421,N_18127);
nor UO_295 (O_295,N_19126,N_19108);
xor UO_296 (O_296,N_19630,N_19776);
or UO_297 (O_297,N_18746,N_18814);
and UO_298 (O_298,N_18940,N_19272);
xnor UO_299 (O_299,N_18346,N_19888);
or UO_300 (O_300,N_18791,N_18003);
nor UO_301 (O_301,N_18159,N_18847);
nor UO_302 (O_302,N_18121,N_19695);
nor UO_303 (O_303,N_18648,N_18857);
or UO_304 (O_304,N_19594,N_18954);
xor UO_305 (O_305,N_19734,N_18185);
or UO_306 (O_306,N_19139,N_19268);
or UO_307 (O_307,N_19028,N_18078);
and UO_308 (O_308,N_19514,N_18670);
and UO_309 (O_309,N_18991,N_18444);
or UO_310 (O_310,N_18978,N_18286);
nor UO_311 (O_311,N_18871,N_19375);
nor UO_312 (O_312,N_18745,N_19743);
or UO_313 (O_313,N_19173,N_18643);
nand UO_314 (O_314,N_18953,N_19643);
xor UO_315 (O_315,N_19218,N_18384);
and UO_316 (O_316,N_18328,N_19819);
and UO_317 (O_317,N_18937,N_18418);
or UO_318 (O_318,N_18793,N_18541);
or UO_319 (O_319,N_18979,N_18660);
nand UO_320 (O_320,N_19930,N_18050);
nor UO_321 (O_321,N_18248,N_19355);
nand UO_322 (O_322,N_18504,N_18447);
nand UO_323 (O_323,N_18562,N_19983);
nand UO_324 (O_324,N_19730,N_19875);
xor UO_325 (O_325,N_19010,N_19669);
nand UO_326 (O_326,N_19059,N_19301);
or UO_327 (O_327,N_19217,N_19618);
nand UO_328 (O_328,N_18203,N_19037);
nor UO_329 (O_329,N_18296,N_18308);
nand UO_330 (O_330,N_19893,N_18437);
nand UO_331 (O_331,N_18932,N_19061);
xor UO_332 (O_332,N_19942,N_19261);
xnor UO_333 (O_333,N_19320,N_19240);
nor UO_334 (O_334,N_19635,N_19664);
or UO_335 (O_335,N_18891,N_19115);
nor UO_336 (O_336,N_18337,N_19971);
or UO_337 (O_337,N_18792,N_18267);
nor UO_338 (O_338,N_19153,N_19889);
nor UO_339 (O_339,N_19313,N_18941);
and UO_340 (O_340,N_18923,N_19539);
nor UO_341 (O_341,N_18480,N_19549);
nor UO_342 (O_342,N_18453,N_18729);
nand UO_343 (O_343,N_18687,N_19790);
or UO_344 (O_344,N_19688,N_19651);
or UO_345 (O_345,N_18501,N_18717);
or UO_346 (O_346,N_18048,N_18043);
or UO_347 (O_347,N_18234,N_19159);
nor UO_348 (O_348,N_19880,N_18738);
nor UO_349 (O_349,N_18963,N_19308);
and UO_350 (O_350,N_18152,N_19167);
and UO_351 (O_351,N_19555,N_19745);
nor UO_352 (O_352,N_18175,N_19481);
and UO_353 (O_353,N_18119,N_19140);
and UO_354 (O_354,N_18599,N_19026);
nor UO_355 (O_355,N_18229,N_19711);
xor UO_356 (O_356,N_18241,N_18334);
or UO_357 (O_357,N_19853,N_19961);
nand UO_358 (O_358,N_19400,N_18033);
nand UO_359 (O_359,N_18543,N_18934);
nor UO_360 (O_360,N_18381,N_18573);
or UO_361 (O_361,N_19795,N_18742);
nand UO_362 (O_362,N_19870,N_18983);
or UO_363 (O_363,N_18586,N_18907);
nand UO_364 (O_364,N_18971,N_18473);
and UO_365 (O_365,N_18966,N_18109);
and UO_366 (O_366,N_18026,N_18888);
or UO_367 (O_367,N_18905,N_19895);
nand UO_368 (O_368,N_19221,N_18389);
xnor UO_369 (O_369,N_18868,N_18689);
and UO_370 (O_370,N_19488,N_18609);
nand UO_371 (O_371,N_19082,N_18567);
nor UO_372 (O_372,N_18434,N_19044);
and UO_373 (O_373,N_19529,N_18631);
nor UO_374 (O_374,N_19136,N_19518);
and UO_375 (O_375,N_19414,N_18122);
nand UO_376 (O_376,N_19193,N_19565);
nor UO_377 (O_377,N_18283,N_18521);
nand UO_378 (O_378,N_19742,N_19366);
xnor UO_379 (O_379,N_18065,N_19039);
or UO_380 (O_380,N_19527,N_18785);
nor UO_381 (O_381,N_18369,N_19521);
and UO_382 (O_382,N_19770,N_19679);
and UO_383 (O_383,N_19358,N_19958);
and UO_384 (O_384,N_18343,N_18640);
or UO_385 (O_385,N_19265,N_18667);
or UO_386 (O_386,N_19150,N_19036);
and UO_387 (O_387,N_19407,N_19837);
or UO_388 (O_388,N_19030,N_19479);
and UO_389 (O_389,N_18917,N_19501);
xnor UO_390 (O_390,N_18455,N_18313);
and UO_391 (O_391,N_19763,N_19548);
nand UO_392 (O_392,N_18190,N_19758);
and UO_393 (O_393,N_18699,N_19716);
and UO_394 (O_394,N_19725,N_18161);
or UO_395 (O_395,N_18029,N_18141);
nor UO_396 (O_396,N_18446,N_18881);
nor UO_397 (O_397,N_19909,N_19143);
nor UO_398 (O_398,N_19354,N_18143);
and UO_399 (O_399,N_19202,N_18691);
and UO_400 (O_400,N_18988,N_18724);
or UO_401 (O_401,N_18929,N_18676);
xnor UO_402 (O_402,N_19487,N_19877);
or UO_403 (O_403,N_18302,N_18580);
or UO_404 (O_404,N_18266,N_19016);
nor UO_405 (O_405,N_19223,N_18025);
xnor UO_406 (O_406,N_19199,N_18510);
or UO_407 (O_407,N_18572,N_18323);
nand UO_408 (O_408,N_18350,N_19826);
xnor UO_409 (O_409,N_19045,N_19794);
nor UO_410 (O_410,N_18273,N_18100);
and UO_411 (O_411,N_19617,N_18128);
and UO_412 (O_412,N_18331,N_18031);
and UO_413 (O_413,N_19303,N_18466);
nor UO_414 (O_414,N_18974,N_18158);
nand UO_415 (O_415,N_18028,N_18770);
nor UO_416 (O_416,N_19469,N_18139);
nor UO_417 (O_417,N_18560,N_18569);
or UO_418 (O_418,N_19074,N_18620);
or UO_419 (O_419,N_18827,N_19219);
xor UO_420 (O_420,N_19641,N_19923);
nand UO_421 (O_421,N_18181,N_18468);
or UO_422 (O_422,N_19112,N_18212);
or UO_423 (O_423,N_19557,N_19511);
and UO_424 (O_424,N_18347,N_18290);
or UO_425 (O_425,N_18680,N_19011);
nand UO_426 (O_426,N_19867,N_18295);
or UO_427 (O_427,N_19163,N_18693);
nand UO_428 (O_428,N_19257,N_18879);
or UO_429 (O_429,N_18918,N_18582);
or UO_430 (O_430,N_19773,N_18354);
nand UO_431 (O_431,N_18679,N_18970);
nor UO_432 (O_432,N_19406,N_18299);
and UO_433 (O_433,N_19022,N_18520);
or UO_434 (O_434,N_18104,N_19943);
or UO_435 (O_435,N_19605,N_19673);
xor UO_436 (O_436,N_19799,N_18678);
xor UO_437 (O_437,N_19357,N_18098);
xnor UO_438 (O_438,N_19946,N_18492);
or UO_439 (O_439,N_18659,N_18189);
nand UO_440 (O_440,N_19064,N_19517);
nand UO_441 (O_441,N_18187,N_19178);
nor UO_442 (O_442,N_18366,N_18927);
or UO_443 (O_443,N_18820,N_19004);
and UO_444 (O_444,N_18499,N_18877);
nand UO_445 (O_445,N_19426,N_18645);
nor UO_446 (O_446,N_18194,N_19083);
xor UO_447 (O_447,N_18982,N_18027);
nand UO_448 (O_448,N_18046,N_18483);
nand UO_449 (O_449,N_19906,N_18942);
or UO_450 (O_450,N_19823,N_18768);
and UO_451 (O_451,N_18215,N_18756);
or UO_452 (O_452,N_18935,N_19189);
nand UO_453 (O_453,N_18281,N_18481);
nor UO_454 (O_454,N_19005,N_18757);
xor UO_455 (O_455,N_18506,N_18166);
or UO_456 (O_456,N_18084,N_19863);
and UO_457 (O_457,N_19530,N_18530);
or UO_458 (O_458,N_18873,N_19458);
nor UO_459 (O_459,N_19325,N_19226);
xnor UO_460 (O_460,N_19992,N_18327);
nand UO_461 (O_461,N_19937,N_18408);
and UO_462 (O_462,N_19152,N_18549);
nor UO_463 (O_463,N_19253,N_19374);
and UO_464 (O_464,N_19865,N_19499);
nand UO_465 (O_465,N_19601,N_19417);
xor UO_466 (O_466,N_19493,N_19141);
nand UO_467 (O_467,N_18782,N_19060);
nand UO_468 (O_468,N_19559,N_18606);
or UO_469 (O_469,N_19348,N_18469);
or UO_470 (O_470,N_19484,N_18886);
xor UO_471 (O_471,N_18023,N_19411);
or UO_472 (O_472,N_19185,N_19702);
nand UO_473 (O_473,N_18800,N_18349);
and UO_474 (O_474,N_18228,N_19636);
or UO_475 (O_475,N_18242,N_18405);
nand UO_476 (O_476,N_19007,N_18962);
and UO_477 (O_477,N_18315,N_18474);
or UO_478 (O_478,N_18841,N_18264);
nand UO_479 (O_479,N_18256,N_18630);
xnor UO_480 (O_480,N_19531,N_19876);
nand UO_481 (O_481,N_19231,N_18244);
nand UO_482 (O_482,N_18591,N_18202);
nor UO_483 (O_483,N_19254,N_19416);
nor UO_484 (O_484,N_18125,N_18355);
xor UO_485 (O_485,N_18906,N_19119);
or UO_486 (O_486,N_19810,N_18798);
nand UO_487 (O_487,N_18590,N_18061);
nor UO_488 (O_488,N_18865,N_19564);
or UO_489 (O_489,N_19148,N_19329);
and UO_490 (O_490,N_18692,N_18092);
and UO_491 (O_491,N_19122,N_19023);
nor UO_492 (O_492,N_18581,N_18051);
nor UO_493 (O_493,N_18107,N_18303);
or UO_494 (O_494,N_19570,N_19733);
nor UO_495 (O_495,N_19098,N_19506);
xnor UO_496 (O_496,N_18424,N_18688);
nor UO_497 (O_497,N_18517,N_19238);
and UO_498 (O_498,N_18379,N_19038);
or UO_499 (O_499,N_18096,N_18117);
and UO_500 (O_500,N_18493,N_18431);
nor UO_501 (O_501,N_19677,N_18227);
and UO_502 (O_502,N_19587,N_18330);
xnor UO_503 (O_503,N_18475,N_18844);
or UO_504 (O_504,N_18594,N_18169);
and UO_505 (O_505,N_19583,N_19898);
xnor UO_506 (O_506,N_19447,N_18981);
nand UO_507 (O_507,N_18778,N_19638);
or UO_508 (O_508,N_18718,N_18006);
nand UO_509 (O_509,N_18628,N_18750);
nor UO_510 (O_510,N_19622,N_18095);
and UO_511 (O_511,N_19379,N_19155);
or UO_512 (O_512,N_18547,N_18605);
or UO_513 (O_513,N_19684,N_19276);
or UO_514 (O_514,N_19080,N_18421);
or UO_515 (O_515,N_19739,N_19120);
xnor UO_516 (O_516,N_18305,N_18157);
xnor UO_517 (O_517,N_19278,N_18998);
nor UO_518 (O_518,N_19789,N_18884);
and UO_519 (O_519,N_18053,N_19456);
and UO_520 (O_520,N_19674,N_19913);
or UO_521 (O_521,N_18583,N_19385);
or UO_522 (O_522,N_19402,N_19938);
and UO_523 (O_523,N_19389,N_18259);
nand UO_524 (O_524,N_19435,N_18099);
or UO_525 (O_525,N_18759,N_18134);
and UO_526 (O_526,N_19613,N_19212);
nor UO_527 (O_527,N_18890,N_18876);
or UO_528 (O_528,N_19225,N_18338);
or UO_529 (O_529,N_18772,N_19097);
or UO_530 (O_530,N_18835,N_18375);
xor UO_531 (O_531,N_19522,N_19784);
nand UO_532 (O_532,N_18352,N_18094);
or UO_533 (O_533,N_18325,N_18007);
nor UO_534 (O_534,N_19297,N_18672);
or UO_535 (O_535,N_19220,N_18823);
nor UO_536 (O_536,N_19031,N_19243);
or UO_537 (O_537,N_18123,N_18601);
or UO_538 (O_538,N_19269,N_19248);
and UO_539 (O_539,N_19422,N_18404);
or UO_540 (O_540,N_18845,N_19213);
nor UO_541 (O_541,N_18304,N_19553);
nor UO_542 (O_542,N_19970,N_19507);
or UO_543 (O_543,N_18723,N_18058);
nand UO_544 (O_544,N_19681,N_18374);
nor UO_545 (O_545,N_18677,N_19873);
and UO_546 (O_546,N_19485,N_19831);
xor UO_547 (O_547,N_19772,N_19446);
or UO_548 (O_548,N_19835,N_19675);
nand UO_549 (O_549,N_18832,N_19885);
or UO_550 (O_550,N_18529,N_18036);
and UO_551 (O_551,N_18860,N_19390);
nor UO_552 (O_552,N_18880,N_18807);
nor UO_553 (O_553,N_19822,N_19256);
nand UO_554 (O_554,N_18824,N_19884);
and UO_555 (O_555,N_18992,N_19891);
and UO_556 (O_556,N_19086,N_18160);
nand UO_557 (O_557,N_18758,N_18450);
nand UO_558 (O_558,N_18114,N_18883);
nor UO_559 (O_559,N_18088,N_19365);
and UO_560 (O_560,N_19224,N_18413);
nor UO_561 (O_561,N_18875,N_19048);
xnor UO_562 (O_562,N_18933,N_19551);
nor UO_563 (O_563,N_18825,N_18062);
or UO_564 (O_564,N_18120,N_18826);
or UO_565 (O_565,N_18566,N_18801);
nand UO_566 (O_566,N_19371,N_18452);
nand UO_567 (O_567,N_18495,N_19425);
and UO_568 (O_568,N_18850,N_18422);
or UO_569 (O_569,N_19085,N_18542);
or UO_570 (O_570,N_18427,N_19346);
nand UO_571 (O_571,N_18042,N_18967);
nor UO_572 (O_572,N_19682,N_18710);
xor UO_573 (O_573,N_18430,N_19554);
or UO_574 (O_574,N_19662,N_18682);
or UO_575 (O_575,N_19678,N_19586);
and UO_576 (O_576,N_19825,N_18551);
nand UO_577 (O_577,N_19249,N_19746);
nand UO_578 (O_578,N_19160,N_18348);
xor UO_579 (O_579,N_19008,N_19899);
and UO_580 (O_580,N_19984,N_18706);
or UO_581 (O_581,N_18236,N_19195);
nand UO_582 (O_582,N_19595,N_18822);
or UO_583 (O_583,N_18395,N_18044);
and UO_584 (O_584,N_19779,N_18287);
and UO_585 (O_585,N_18009,N_18901);
nand UO_586 (O_586,N_19616,N_18219);
nor UO_587 (O_587,N_18054,N_18781);
and UO_588 (O_588,N_19520,N_18993);
or UO_589 (O_589,N_18681,N_18103);
nand UO_590 (O_590,N_19186,N_18615);
or UO_591 (O_591,N_18001,N_18843);
nor UO_592 (O_592,N_18401,N_19897);
or UO_593 (O_593,N_18545,N_18553);
and UO_594 (O_594,N_18069,N_19604);
or UO_595 (O_595,N_19081,N_18938);
nor UO_596 (O_596,N_18230,N_18775);
and UO_597 (O_597,N_19935,N_18237);
and UO_598 (O_598,N_18949,N_18010);
nor UO_599 (O_599,N_18894,N_18755);
and UO_600 (O_600,N_19096,N_18588);
nand UO_601 (O_601,N_19123,N_18425);
or UO_602 (O_602,N_18293,N_19861);
nor UO_603 (O_603,N_18018,N_19332);
xor UO_604 (O_604,N_19187,N_19561);
and UO_605 (O_605,N_19027,N_19121);
nand UO_606 (O_606,N_18509,N_18612);
and UO_607 (O_607,N_18249,N_19091);
nand UO_608 (O_608,N_18819,N_18253);
nor UO_609 (O_609,N_19637,N_19856);
and UO_610 (O_610,N_18839,N_18810);
nand UO_611 (O_611,N_19603,N_18836);
nand UO_612 (O_612,N_18766,N_18454);
and UO_613 (O_613,N_19457,N_19841);
and UO_614 (O_614,N_18731,N_19273);
xnor UO_615 (O_615,N_18654,N_19104);
nand UO_616 (O_616,N_18943,N_18646);
nand UO_617 (O_617,N_19166,N_19667);
or UO_618 (O_618,N_19317,N_18231);
and UO_619 (O_619,N_18361,N_19088);
nor UO_620 (O_620,N_19927,N_19544);
and UO_621 (O_621,N_19968,N_19858);
or UO_622 (O_622,N_19959,N_18113);
nand UO_623 (O_623,N_19384,N_19465);
nor UO_624 (O_624,N_18357,N_18733);
xnor UO_625 (O_625,N_19668,N_18584);
and UO_626 (O_626,N_19990,N_18944);
nand UO_627 (O_627,N_18952,N_18435);
xor UO_628 (O_628,N_19280,N_18326);
or UO_629 (O_629,N_19812,N_19687);
and UO_630 (O_630,N_19721,N_19656);
and UO_631 (O_631,N_19428,N_19076);
nor UO_632 (O_632,N_18852,N_19298);
xnor UO_633 (O_633,N_19483,N_18945);
and UO_634 (O_634,N_19963,N_19111);
nand UO_635 (O_635,N_18224,N_18173);
nand UO_636 (O_636,N_18204,N_19610);
nand UO_637 (O_637,N_19228,N_18959);
or UO_638 (O_638,N_18585,N_18142);
or UO_639 (O_639,N_19181,N_19000);
or UO_640 (O_640,N_18429,N_18116);
nor UO_641 (O_641,N_19168,N_19050);
or UO_642 (O_642,N_19500,N_19950);
nand UO_643 (O_643,N_19981,N_18817);
or UO_644 (O_644,N_18799,N_18397);
and UO_645 (O_645,N_19676,N_19144);
or UO_646 (O_646,N_18035,N_19538);
nand UO_647 (O_647,N_19396,N_19413);
and UO_648 (O_648,N_19846,N_18924);
nand UO_649 (O_649,N_19552,N_18618);
nor UO_650 (O_650,N_18167,N_19035);
nor UO_651 (O_651,N_18811,N_19840);
xnor UO_652 (O_652,N_18318,N_19737);
or UO_653 (O_653,N_19575,N_18951);
or UO_654 (O_654,N_18730,N_19275);
nor UO_655 (O_655,N_19597,N_18671);
nand UO_656 (O_656,N_19452,N_18459);
or UO_657 (O_657,N_18725,N_19051);
or UO_658 (O_658,N_18821,N_19347);
nor UO_659 (O_659,N_18406,N_18684);
nor UO_660 (O_660,N_19310,N_19418);
and UO_661 (O_661,N_19997,N_18195);
or UO_662 (O_662,N_18118,N_18360);
or UO_663 (O_663,N_19787,N_18727);
and UO_664 (O_664,N_19340,N_19170);
xnor UO_665 (O_665,N_18045,N_19995);
or UO_666 (O_666,N_19285,N_18763);
nand UO_667 (O_667,N_19006,N_18828);
nor UO_668 (O_668,N_18156,N_19359);
xor UO_669 (O_669,N_18130,N_19602);
and UO_670 (O_670,N_19274,N_18973);
or UO_671 (O_671,N_18872,N_19373);
nor UO_672 (O_672,N_19537,N_18005);
nand UO_673 (O_673,N_18743,N_19077);
and UO_674 (O_674,N_18683,N_19598);
nor UO_675 (O_675,N_18345,N_18097);
nor UO_676 (O_676,N_18626,N_19046);
and UO_677 (O_677,N_18721,N_19147);
or UO_678 (O_678,N_19482,N_18637);
and UO_679 (O_679,N_18279,N_18131);
xnor UO_680 (O_680,N_18577,N_18769);
xnor UO_681 (O_681,N_18022,N_18449);
nor UO_682 (O_682,N_18364,N_19377);
nor UO_683 (O_683,N_19277,N_18711);
xor UO_684 (O_684,N_19573,N_19864);
xor UO_685 (O_685,N_18052,N_18015);
and UO_686 (O_686,N_18278,N_18624);
xnor UO_687 (O_687,N_18518,N_18762);
or UO_688 (O_688,N_19574,N_18439);
or UO_689 (O_689,N_19855,N_19691);
nand UO_690 (O_690,N_19292,N_18783);
or UO_691 (O_691,N_19869,N_18887);
nor UO_692 (O_692,N_19703,N_18471);
nand UO_693 (O_693,N_18914,N_19309);
and UO_694 (O_694,N_18170,N_19849);
nor UO_695 (O_695,N_19931,N_18407);
and UO_696 (O_696,N_18773,N_18861);
nand UO_697 (O_697,N_19515,N_19191);
xnor UO_698 (O_698,N_18508,N_18892);
nor UO_699 (O_699,N_18908,N_19657);
nor UO_700 (O_700,N_19351,N_19162);
nor UO_701 (O_701,N_19510,N_19723);
nor UO_702 (O_702,N_19033,N_19736);
and UO_703 (O_703,N_18383,N_18193);
and UO_704 (O_704,N_19151,N_18411);
nand UO_705 (O_705,N_18163,N_18621);
and UO_706 (O_706,N_19615,N_19917);
nor UO_707 (O_707,N_18108,N_18593);
nor UO_708 (O_708,N_18188,N_19932);
nand UO_709 (O_709,N_18525,N_19397);
nand UO_710 (O_710,N_19475,N_18997);
nand UO_711 (O_711,N_18172,N_19724);
nand UO_712 (O_712,N_18276,N_19572);
nor UO_713 (O_713,N_19788,N_19833);
nand UO_714 (O_714,N_19710,N_18298);
or UO_715 (O_715,N_18309,N_19092);
nand UO_716 (O_716,N_18067,N_19235);
and UO_717 (O_717,N_19237,N_18147);
nand UO_718 (O_718,N_18329,N_19965);
and UO_719 (O_719,N_18138,N_18747);
nand UO_720 (O_720,N_18863,N_19214);
nand UO_721 (O_721,N_19584,N_18524);
or UO_722 (O_722,N_18576,N_19430);
nor UO_723 (O_723,N_19769,N_18975);
or UO_724 (O_724,N_18460,N_19403);
nor UO_725 (O_725,N_18665,N_19383);
xnor UO_726 (O_726,N_19436,N_19802);
and UO_727 (O_727,N_19820,N_19042);
and UO_728 (O_728,N_18059,N_19798);
and UO_729 (O_729,N_18148,N_18899);
nor UO_730 (O_730,N_18546,N_19599);
or UO_731 (O_731,N_18011,N_18777);
xor UO_732 (O_732,N_19070,N_19879);
nand UO_733 (O_733,N_18240,N_19672);
nand UO_734 (O_734,N_19956,N_19100);
or UO_735 (O_735,N_18207,N_19834);
and UO_736 (O_736,N_19689,N_19184);
and UO_737 (O_737,N_18030,N_18603);
or UO_738 (O_738,N_18359,N_19944);
or UO_739 (O_739,N_18075,N_19194);
or UO_740 (O_740,N_18090,N_19986);
nor UO_741 (O_741,N_18324,N_18232);
and UO_742 (O_742,N_19338,N_18644);
or UO_743 (O_743,N_18760,N_19129);
nand UO_744 (O_744,N_19782,N_19149);
nand UO_745 (O_745,N_19018,N_19327);
xor UO_746 (O_746,N_19205,N_18690);
nand UO_747 (O_747,N_19382,N_19791);
and UO_748 (O_748,N_19072,N_18882);
and UO_749 (O_749,N_19732,N_18417);
nor UO_750 (O_750,N_18834,N_19633);
nor UO_751 (O_751,N_18456,N_18462);
nor UO_752 (O_752,N_19118,N_19881);
nand UO_753 (O_753,N_18344,N_19720);
nand UO_754 (O_754,N_19295,N_19526);
xnor UO_755 (O_755,N_19816,N_18403);
nor UO_756 (O_756,N_18294,N_18060);
or UO_757 (O_757,N_18016,N_19807);
nand UO_758 (O_758,N_19230,N_18079);
or UO_759 (O_759,N_18761,N_18024);
nand UO_760 (O_760,N_18728,N_19490);
and UO_761 (O_761,N_19611,N_18635);
nor UO_762 (O_762,N_19322,N_18391);
xnor UO_763 (O_763,N_19631,N_19781);
nor UO_764 (O_764,N_19473,N_18235);
nor UO_765 (O_765,N_18748,N_19974);
or UO_766 (O_766,N_19887,N_19367);
nor UO_767 (O_767,N_19182,N_19852);
and UO_768 (O_768,N_19934,N_18858);
and UO_769 (O_769,N_18124,N_18463);
nand UO_770 (O_770,N_19312,N_18840);
and UO_771 (O_771,N_18657,N_19399);
nor UO_772 (O_772,N_18568,N_19069);
nor UO_773 (O_773,N_18465,N_19857);
or UO_774 (O_774,N_19437,N_19337);
xor UO_775 (O_775,N_19012,N_18673);
and UO_776 (O_776,N_18479,N_18486);
and UO_777 (O_777,N_18505,N_18333);
nand UO_778 (O_778,N_19463,N_18965);
nor UO_779 (O_779,N_19283,N_19786);
and UO_780 (O_780,N_18055,N_19813);
and UO_781 (O_781,N_18080,N_18191);
nor UO_782 (O_782,N_19953,N_18900);
xnor UO_783 (O_783,N_19874,N_19281);
xor UO_784 (O_784,N_18587,N_18057);
nand UO_785 (O_785,N_19071,N_19663);
and UO_786 (O_786,N_18804,N_18519);
or UO_787 (O_787,N_19461,N_19302);
and UO_788 (O_788,N_19821,N_18133);
and UO_789 (O_789,N_19318,N_19612);
nand UO_790 (O_790,N_19450,N_19492);
or UO_791 (O_791,N_19472,N_19670);
nand UO_792 (O_792,N_19760,N_18904);
and UO_793 (O_793,N_19632,N_18776);
or UO_794 (O_794,N_19299,N_18340);
or UO_795 (O_795,N_19625,N_19408);
xor UO_796 (O_796,N_19415,N_19991);
or UO_797 (O_797,N_19647,N_18358);
nand UO_798 (O_798,N_19180,N_18734);
nand UO_799 (O_799,N_18162,N_19814);
xnor UO_800 (O_800,N_18753,N_19259);
nor UO_801 (O_801,N_19145,N_19360);
and UO_802 (O_802,N_19941,N_18919);
nand UO_803 (O_803,N_19032,N_19239);
xnor UO_804 (O_804,N_18260,N_18862);
xnor UO_805 (O_805,N_19486,N_18578);
or UO_806 (O_806,N_18322,N_18478);
nand UO_807 (O_807,N_19306,N_18037);
and UO_808 (O_808,N_19759,N_19350);
or UO_809 (O_809,N_18213,N_18105);
or UO_810 (O_810,N_19513,N_19034);
nor UO_811 (O_811,N_19847,N_19563);
nor UO_812 (O_812,N_19336,N_18859);
nand UO_813 (O_813,N_19778,N_19451);
and UO_814 (O_814,N_19987,N_19066);
nor UO_815 (O_815,N_18451,N_18697);
nand UO_816 (O_816,N_18739,N_18653);
nor UO_817 (O_817,N_18651,N_19440);
nand UO_818 (O_818,N_18377,N_18795);
and UO_819 (O_819,N_19489,N_19293);
nor UO_820 (O_820,N_18855,N_18301);
nor UO_821 (O_821,N_19694,N_18666);
nand UO_822 (O_822,N_18837,N_19142);
or UO_823 (O_823,N_19871,N_19498);
and UO_824 (O_824,N_19003,N_18136);
or UO_825 (O_825,N_19304,N_19979);
nand UO_826 (O_826,N_18744,N_18604);
and UO_827 (O_827,N_18977,N_18126);
nand UO_828 (O_828,N_19591,N_19532);
nor UO_829 (O_829,N_18867,N_18472);
nand UO_830 (O_830,N_18306,N_18909);
and UO_831 (O_831,N_18790,N_18720);
nor UO_832 (O_832,N_19646,N_18502);
nand UO_833 (O_833,N_18254,N_18964);
nand UO_834 (O_834,N_19523,N_19015);
or UO_835 (O_835,N_19866,N_18642);
xor UO_836 (O_836,N_19976,N_19775);
nand UO_837 (O_837,N_19904,N_18632);
nor UO_838 (O_838,N_19362,N_19993);
nor UO_839 (O_839,N_18740,N_19099);
and UO_840 (O_840,N_18874,N_19393);
nor UO_841 (O_841,N_18574,N_19900);
or UO_842 (O_842,N_18557,N_19838);
or UO_843 (O_843,N_19542,N_18307);
and UO_844 (O_844,N_19886,N_18485);
or UO_845 (O_845,N_18145,N_18371);
and UO_846 (O_846,N_18317,N_18916);
xnor UO_847 (O_847,N_19797,N_19793);
xor UO_848 (O_848,N_19911,N_18619);
nand UO_849 (O_849,N_19444,N_18818);
nand UO_850 (O_850,N_18512,N_19049);
and UO_851 (O_851,N_18561,N_19391);
nor UO_852 (O_852,N_18607,N_19315);
and UO_853 (O_853,N_19748,N_19462);
or UO_854 (O_854,N_19751,N_19410);
nand UO_855 (O_855,N_19266,N_19660);
nand UO_856 (O_856,N_18014,N_18284);
nor UO_857 (O_857,N_19405,N_19901);
or UO_858 (O_858,N_18034,N_18939);
or UO_859 (O_859,N_19495,N_19624);
nor UO_860 (O_860,N_19608,N_18077);
nand UO_861 (O_861,N_18209,N_19491);
or UO_862 (O_862,N_18049,N_18297);
nor UO_863 (O_863,N_19509,N_18491);
or UO_864 (O_864,N_19116,N_19550);
or UO_865 (O_865,N_18754,N_19980);
nor UO_866 (O_866,N_18039,N_18885);
or UO_867 (O_867,N_18020,N_18833);
nor UO_868 (O_868,N_18805,N_19714);
nor UO_869 (O_869,N_18255,N_18289);
or UO_870 (O_870,N_18854,N_19671);
nor UO_871 (O_871,N_18995,N_19567);
or UO_872 (O_872,N_18013,N_19427);
and UO_873 (O_873,N_18598,N_18878);
nand UO_874 (O_874,N_19062,N_19805);
xor UO_875 (O_875,N_18200,N_19844);
or UO_876 (O_876,N_18272,N_19558);
or UO_877 (O_877,N_19448,N_18629);
nand UO_878 (O_878,N_18652,N_19619);
and UO_879 (O_879,N_19818,N_19585);
and UO_880 (O_880,N_19949,N_19659);
nor UO_881 (O_881,N_19131,N_18662);
xor UO_882 (O_882,N_19114,N_19839);
xnor UO_883 (O_883,N_18083,N_18930);
nor UO_884 (O_884,N_18488,N_19718);
nand UO_885 (O_885,N_19708,N_19756);
or UO_886 (O_886,N_18386,N_19073);
nor UO_887 (O_887,N_18737,N_18538);
nand UO_888 (O_888,N_19068,N_18151);
xor UO_889 (O_889,N_19996,N_18902);
xnor UO_890 (O_890,N_19127,N_19648);
and UO_891 (O_891,N_19024,N_18708);
nor UO_892 (O_892,N_18985,N_19132);
nor UO_893 (O_893,N_19768,N_19801);
and UO_894 (O_894,N_19445,N_18780);
and UO_895 (O_895,N_19466,N_19966);
or UO_896 (O_896,N_19380,N_18225);
or UO_897 (O_897,N_19808,N_19262);
nand UO_898 (O_898,N_19824,N_19639);
nor UO_899 (O_899,N_19258,N_19161);
or UO_900 (O_900,N_18956,N_18438);
nand UO_901 (O_901,N_18535,N_18503);
nor UO_902 (O_902,N_18470,N_18110);
and UO_903 (O_903,N_19815,N_18698);
and UO_904 (O_904,N_19084,N_18252);
and UO_905 (O_905,N_19158,N_18936);
and UO_906 (O_906,N_19065,N_18732);
nand UO_907 (O_907,N_18713,N_19696);
xnor UO_908 (O_908,N_18864,N_19041);
nand UO_909 (O_909,N_19352,N_18788);
and UO_910 (O_910,N_19741,N_19967);
nand UO_911 (O_911,N_19977,N_18461);
nor UO_912 (O_912,N_18596,N_18214);
and UO_913 (O_913,N_18986,N_18571);
nor UO_914 (O_914,N_18602,N_19401);
nor UO_915 (O_915,N_18915,N_18686);
and UO_916 (O_916,N_18558,N_19982);
xnor UO_917 (O_917,N_19113,N_18210);
nor UO_918 (O_918,N_18063,N_19665);
nand UO_919 (O_919,N_18310,N_19766);
nor UO_920 (O_920,N_18087,N_18467);
or UO_921 (O_921,N_18515,N_18198);
or UO_922 (O_922,N_19478,N_19474);
nor UO_923 (O_923,N_19043,N_19727);
xor UO_924 (O_924,N_19442,N_19596);
and UO_925 (O_925,N_18550,N_19860);
nor UO_926 (O_926,N_18178,N_19780);
and UO_927 (O_927,N_19409,N_18570);
or UO_928 (O_928,N_19183,N_18245);
and UO_929 (O_929,N_18813,N_19215);
or UO_930 (O_930,N_19842,N_19916);
and UO_931 (O_931,N_18489,N_19556);
and UO_932 (O_932,N_19331,N_19439);
nand UO_933 (O_933,N_18664,N_19311);
nor UO_934 (O_934,N_19206,N_18661);
nor UO_935 (O_935,N_18920,N_19690);
nand UO_936 (O_936,N_19581,N_18316);
nand UO_937 (O_937,N_18808,N_19333);
nor UO_938 (O_938,N_19471,N_18633);
nor UO_939 (O_939,N_19541,N_18563);
nor UO_940 (O_940,N_18441,N_18332);
or UO_941 (O_941,N_18931,N_19353);
nor UO_942 (O_942,N_19750,N_18554);
and UO_943 (O_943,N_19324,N_18335);
nand UO_944 (O_944,N_18597,N_19543);
and UO_945 (O_945,N_18270,N_19201);
or UO_946 (O_946,N_19395,N_18705);
and UO_947 (O_947,N_19335,N_19378);
xor UO_948 (O_948,N_18848,N_19609);
or UO_949 (O_949,N_19540,N_19305);
nand UO_950 (O_950,N_18218,N_18258);
and UO_951 (O_951,N_18913,N_18794);
nor UO_952 (O_952,N_19090,N_18715);
xnor UO_953 (O_953,N_18816,N_18341);
nand UO_954 (O_954,N_18968,N_19712);
and UO_955 (O_955,N_19419,N_19994);
nand UO_956 (O_956,N_18536,N_18853);
nor UO_957 (O_957,N_18164,N_18926);
nand UO_958 (O_958,N_18500,N_18870);
nor UO_959 (O_959,N_19939,N_19109);
xnor UO_960 (O_960,N_18719,N_19868);
or UO_961 (O_961,N_18073,N_19571);
nand UO_962 (O_962,N_18150,N_18399);
nand UO_963 (O_963,N_18996,N_19843);
nand UO_964 (O_964,N_19693,N_18797);
or UO_965 (O_965,N_19792,N_19704);
or UO_966 (O_966,N_19372,N_19634);
nand UO_967 (O_967,N_19137,N_19434);
or UO_968 (O_968,N_19749,N_19497);
nor UO_969 (O_969,N_18458,N_19014);
and UO_970 (O_970,N_19828,N_18415);
and UO_971 (O_971,N_19345,N_19685);
nand UO_972 (O_972,N_18851,N_19103);
or UO_973 (O_973,N_19717,N_19019);
and UO_974 (O_974,N_19429,N_18115);
and UO_975 (O_975,N_19242,N_18540);
and UO_976 (O_976,N_19296,N_19528);
nand UO_977 (O_977,N_19644,N_18076);
or UO_978 (O_978,N_19525,N_18786);
nor UO_979 (O_979,N_19477,N_18004);
xnor UO_980 (O_980,N_19764,N_18089);
nor UO_981 (O_981,N_18701,N_19757);
nor UO_982 (O_982,N_18514,N_19680);
or UO_983 (O_983,N_18068,N_18183);
nand UO_984 (O_984,N_18216,N_18019);
and UO_985 (O_985,N_18047,N_18707);
or UO_986 (O_986,N_19752,N_19626);
nor UO_987 (O_987,N_19056,N_18552);
nand UO_988 (O_988,N_19300,N_18669);
or UO_989 (O_989,N_18440,N_18038);
nand UO_990 (O_990,N_18611,N_19800);
xor UO_991 (O_991,N_18696,N_19666);
and UO_992 (O_992,N_19341,N_19892);
xnor UO_993 (O_993,N_19972,N_19270);
nor UO_994 (O_994,N_18271,N_18442);
or UO_995 (O_995,N_18487,N_18291);
or UO_996 (O_996,N_18663,N_19578);
nor UO_997 (O_997,N_19087,N_18712);
nor UO_998 (O_998,N_19654,N_18592);
nor UO_999 (O_999,N_18362,N_18342);
nand UO_1000 (O_1000,N_19737,N_19807);
and UO_1001 (O_1001,N_19011,N_18924);
nand UO_1002 (O_1002,N_18407,N_18257);
nand UO_1003 (O_1003,N_18185,N_18328);
and UO_1004 (O_1004,N_19190,N_19964);
or UO_1005 (O_1005,N_18938,N_18530);
or UO_1006 (O_1006,N_19733,N_19481);
nand UO_1007 (O_1007,N_19078,N_18131);
and UO_1008 (O_1008,N_19887,N_18750);
nand UO_1009 (O_1009,N_18057,N_18868);
xnor UO_1010 (O_1010,N_19860,N_19150);
or UO_1011 (O_1011,N_19742,N_18969);
and UO_1012 (O_1012,N_19872,N_19003);
or UO_1013 (O_1013,N_19557,N_19370);
nand UO_1014 (O_1014,N_18982,N_18177);
or UO_1015 (O_1015,N_18290,N_18764);
nand UO_1016 (O_1016,N_18441,N_19121);
nand UO_1017 (O_1017,N_18048,N_19473);
xnor UO_1018 (O_1018,N_19369,N_19965);
nand UO_1019 (O_1019,N_18256,N_18904);
nor UO_1020 (O_1020,N_19344,N_18673);
and UO_1021 (O_1021,N_19394,N_18384);
nor UO_1022 (O_1022,N_18596,N_19235);
nor UO_1023 (O_1023,N_19564,N_19971);
nor UO_1024 (O_1024,N_19342,N_18982);
or UO_1025 (O_1025,N_18970,N_19571);
and UO_1026 (O_1026,N_18535,N_19854);
nor UO_1027 (O_1027,N_18428,N_18282);
or UO_1028 (O_1028,N_18015,N_18345);
or UO_1029 (O_1029,N_18089,N_19076);
nor UO_1030 (O_1030,N_19496,N_18808);
nand UO_1031 (O_1031,N_18489,N_18968);
nand UO_1032 (O_1032,N_19970,N_18705);
nor UO_1033 (O_1033,N_19456,N_18584);
or UO_1034 (O_1034,N_18213,N_18151);
xor UO_1035 (O_1035,N_19033,N_18891);
or UO_1036 (O_1036,N_19279,N_18727);
and UO_1037 (O_1037,N_19062,N_19103);
nand UO_1038 (O_1038,N_19630,N_18770);
and UO_1039 (O_1039,N_19506,N_18098);
xor UO_1040 (O_1040,N_18696,N_18103);
or UO_1041 (O_1041,N_19344,N_18614);
nand UO_1042 (O_1042,N_18952,N_19046);
xor UO_1043 (O_1043,N_18739,N_18474);
or UO_1044 (O_1044,N_19830,N_19311);
nor UO_1045 (O_1045,N_19467,N_18828);
or UO_1046 (O_1046,N_18102,N_18291);
nand UO_1047 (O_1047,N_19384,N_19611);
or UO_1048 (O_1048,N_19161,N_18452);
and UO_1049 (O_1049,N_19492,N_18800);
or UO_1050 (O_1050,N_19811,N_18206);
or UO_1051 (O_1051,N_19473,N_18222);
or UO_1052 (O_1052,N_18790,N_18454);
nor UO_1053 (O_1053,N_19542,N_19553);
or UO_1054 (O_1054,N_19162,N_18810);
nor UO_1055 (O_1055,N_19746,N_19809);
or UO_1056 (O_1056,N_19316,N_18407);
or UO_1057 (O_1057,N_19889,N_18909);
and UO_1058 (O_1058,N_18992,N_18877);
nor UO_1059 (O_1059,N_19086,N_19899);
and UO_1060 (O_1060,N_18849,N_18607);
or UO_1061 (O_1061,N_18612,N_18949);
and UO_1062 (O_1062,N_19997,N_18665);
and UO_1063 (O_1063,N_18630,N_18791);
and UO_1064 (O_1064,N_18319,N_18524);
xnor UO_1065 (O_1065,N_19846,N_18874);
or UO_1066 (O_1066,N_19373,N_19298);
xnor UO_1067 (O_1067,N_19718,N_19277);
nand UO_1068 (O_1068,N_19969,N_19722);
nand UO_1069 (O_1069,N_18279,N_18847);
or UO_1070 (O_1070,N_18939,N_18102);
nor UO_1071 (O_1071,N_18675,N_19317);
or UO_1072 (O_1072,N_19348,N_18223);
nand UO_1073 (O_1073,N_18871,N_19726);
and UO_1074 (O_1074,N_19120,N_18128);
xor UO_1075 (O_1075,N_18777,N_18888);
xnor UO_1076 (O_1076,N_19606,N_19823);
xnor UO_1077 (O_1077,N_19370,N_19873);
nor UO_1078 (O_1078,N_18646,N_19018);
or UO_1079 (O_1079,N_18321,N_18069);
nor UO_1080 (O_1080,N_19180,N_19248);
nor UO_1081 (O_1081,N_18889,N_18545);
nand UO_1082 (O_1082,N_18048,N_18372);
and UO_1083 (O_1083,N_19814,N_19395);
nor UO_1084 (O_1084,N_18907,N_19885);
and UO_1085 (O_1085,N_19759,N_18025);
nand UO_1086 (O_1086,N_18800,N_18516);
or UO_1087 (O_1087,N_18290,N_19245);
nand UO_1088 (O_1088,N_19283,N_19575);
and UO_1089 (O_1089,N_18316,N_19194);
and UO_1090 (O_1090,N_18627,N_19801);
nand UO_1091 (O_1091,N_18393,N_19013);
and UO_1092 (O_1092,N_18044,N_18348);
and UO_1093 (O_1093,N_18799,N_19103);
and UO_1094 (O_1094,N_19778,N_18697);
and UO_1095 (O_1095,N_19878,N_18957);
and UO_1096 (O_1096,N_19892,N_18974);
nand UO_1097 (O_1097,N_19263,N_18328);
nor UO_1098 (O_1098,N_18374,N_19178);
or UO_1099 (O_1099,N_18685,N_19540);
nor UO_1100 (O_1100,N_19702,N_18268);
xnor UO_1101 (O_1101,N_19208,N_18420);
nand UO_1102 (O_1102,N_18465,N_19217);
or UO_1103 (O_1103,N_18374,N_19156);
and UO_1104 (O_1104,N_19097,N_19831);
nand UO_1105 (O_1105,N_18113,N_18680);
and UO_1106 (O_1106,N_18195,N_18701);
and UO_1107 (O_1107,N_19215,N_19661);
or UO_1108 (O_1108,N_18038,N_18004);
nand UO_1109 (O_1109,N_19578,N_19572);
nand UO_1110 (O_1110,N_18593,N_18061);
nand UO_1111 (O_1111,N_19679,N_19651);
and UO_1112 (O_1112,N_18578,N_18181);
nand UO_1113 (O_1113,N_18290,N_19605);
and UO_1114 (O_1114,N_19519,N_19239);
xnor UO_1115 (O_1115,N_19649,N_18100);
nand UO_1116 (O_1116,N_18810,N_19095);
or UO_1117 (O_1117,N_19765,N_18223);
and UO_1118 (O_1118,N_18630,N_19376);
nor UO_1119 (O_1119,N_19185,N_19748);
nand UO_1120 (O_1120,N_19515,N_19622);
nand UO_1121 (O_1121,N_18032,N_18972);
or UO_1122 (O_1122,N_19353,N_19273);
nand UO_1123 (O_1123,N_18056,N_18546);
and UO_1124 (O_1124,N_19853,N_19904);
nand UO_1125 (O_1125,N_19778,N_18137);
nor UO_1126 (O_1126,N_19412,N_18727);
and UO_1127 (O_1127,N_19086,N_19672);
nand UO_1128 (O_1128,N_19691,N_18310);
or UO_1129 (O_1129,N_19785,N_18537);
or UO_1130 (O_1130,N_18420,N_19344);
nand UO_1131 (O_1131,N_18556,N_19921);
or UO_1132 (O_1132,N_19354,N_19591);
nand UO_1133 (O_1133,N_18789,N_18195);
and UO_1134 (O_1134,N_18203,N_19983);
or UO_1135 (O_1135,N_19253,N_19356);
nor UO_1136 (O_1136,N_19601,N_18172);
nand UO_1137 (O_1137,N_18024,N_18642);
nor UO_1138 (O_1138,N_18931,N_18301);
nand UO_1139 (O_1139,N_18002,N_18086);
or UO_1140 (O_1140,N_19386,N_18759);
nor UO_1141 (O_1141,N_18285,N_18965);
or UO_1142 (O_1142,N_18594,N_19291);
nand UO_1143 (O_1143,N_18911,N_19355);
nand UO_1144 (O_1144,N_19023,N_18073);
and UO_1145 (O_1145,N_19423,N_18190);
or UO_1146 (O_1146,N_18137,N_19270);
and UO_1147 (O_1147,N_18245,N_18439);
nand UO_1148 (O_1148,N_19820,N_19981);
and UO_1149 (O_1149,N_19588,N_19540);
xnor UO_1150 (O_1150,N_18535,N_18221);
nor UO_1151 (O_1151,N_19420,N_19784);
or UO_1152 (O_1152,N_19687,N_18939);
or UO_1153 (O_1153,N_19687,N_18334);
xnor UO_1154 (O_1154,N_18219,N_18071);
nand UO_1155 (O_1155,N_18177,N_18989);
or UO_1156 (O_1156,N_19141,N_18732);
or UO_1157 (O_1157,N_18850,N_18551);
nor UO_1158 (O_1158,N_19529,N_19448);
or UO_1159 (O_1159,N_19186,N_19083);
or UO_1160 (O_1160,N_18780,N_19686);
and UO_1161 (O_1161,N_19199,N_19523);
or UO_1162 (O_1162,N_18016,N_19442);
or UO_1163 (O_1163,N_18325,N_19918);
and UO_1164 (O_1164,N_18980,N_18131);
nor UO_1165 (O_1165,N_18228,N_18261);
nor UO_1166 (O_1166,N_19556,N_19648);
nor UO_1167 (O_1167,N_19592,N_19765);
nor UO_1168 (O_1168,N_19959,N_19459);
xor UO_1169 (O_1169,N_18094,N_19614);
nor UO_1170 (O_1170,N_18708,N_18637);
and UO_1171 (O_1171,N_19470,N_18863);
nor UO_1172 (O_1172,N_18691,N_19888);
nor UO_1173 (O_1173,N_19825,N_18567);
nand UO_1174 (O_1174,N_18599,N_19282);
and UO_1175 (O_1175,N_18320,N_18346);
and UO_1176 (O_1176,N_18561,N_19461);
nand UO_1177 (O_1177,N_18613,N_18692);
nand UO_1178 (O_1178,N_18875,N_18728);
and UO_1179 (O_1179,N_18057,N_18920);
nand UO_1180 (O_1180,N_19969,N_18666);
nor UO_1181 (O_1181,N_19902,N_19419);
and UO_1182 (O_1182,N_18428,N_18873);
or UO_1183 (O_1183,N_19776,N_18929);
nand UO_1184 (O_1184,N_18593,N_19009);
nand UO_1185 (O_1185,N_19178,N_18916);
xnor UO_1186 (O_1186,N_18140,N_18416);
nand UO_1187 (O_1187,N_18840,N_18905);
and UO_1188 (O_1188,N_19889,N_19049);
and UO_1189 (O_1189,N_19450,N_18570);
and UO_1190 (O_1190,N_19682,N_18364);
or UO_1191 (O_1191,N_19810,N_18947);
xnor UO_1192 (O_1192,N_18759,N_18735);
nand UO_1193 (O_1193,N_19784,N_19648);
or UO_1194 (O_1194,N_19243,N_18282);
or UO_1195 (O_1195,N_18404,N_19125);
and UO_1196 (O_1196,N_18624,N_19112);
nor UO_1197 (O_1197,N_18868,N_18753);
and UO_1198 (O_1198,N_19831,N_19588);
and UO_1199 (O_1199,N_18595,N_18439);
nor UO_1200 (O_1200,N_18407,N_19247);
nor UO_1201 (O_1201,N_19982,N_18799);
and UO_1202 (O_1202,N_19984,N_18064);
nand UO_1203 (O_1203,N_19018,N_18760);
or UO_1204 (O_1204,N_18154,N_19752);
nor UO_1205 (O_1205,N_18076,N_18277);
xor UO_1206 (O_1206,N_18027,N_19982);
or UO_1207 (O_1207,N_19142,N_18289);
xnor UO_1208 (O_1208,N_19450,N_18214);
nor UO_1209 (O_1209,N_19417,N_19808);
nand UO_1210 (O_1210,N_19149,N_19592);
or UO_1211 (O_1211,N_18024,N_18690);
nor UO_1212 (O_1212,N_18789,N_19226);
or UO_1213 (O_1213,N_18267,N_19892);
or UO_1214 (O_1214,N_19088,N_18337);
and UO_1215 (O_1215,N_19622,N_18560);
nand UO_1216 (O_1216,N_19962,N_18776);
and UO_1217 (O_1217,N_19121,N_19536);
or UO_1218 (O_1218,N_19904,N_18291);
and UO_1219 (O_1219,N_19087,N_18746);
and UO_1220 (O_1220,N_19182,N_18230);
nand UO_1221 (O_1221,N_19014,N_18761);
nor UO_1222 (O_1222,N_19050,N_19962);
or UO_1223 (O_1223,N_18241,N_18481);
nand UO_1224 (O_1224,N_19471,N_19798);
nor UO_1225 (O_1225,N_18324,N_18921);
nor UO_1226 (O_1226,N_19980,N_18274);
and UO_1227 (O_1227,N_18670,N_19421);
and UO_1228 (O_1228,N_19030,N_19531);
and UO_1229 (O_1229,N_18795,N_18578);
nor UO_1230 (O_1230,N_19290,N_18022);
and UO_1231 (O_1231,N_19314,N_19384);
or UO_1232 (O_1232,N_18479,N_19478);
or UO_1233 (O_1233,N_18654,N_18057);
nor UO_1234 (O_1234,N_19695,N_18449);
xnor UO_1235 (O_1235,N_19709,N_18264);
or UO_1236 (O_1236,N_18047,N_19324);
xor UO_1237 (O_1237,N_19990,N_19564);
nand UO_1238 (O_1238,N_19260,N_18917);
nor UO_1239 (O_1239,N_18863,N_18651);
nand UO_1240 (O_1240,N_18144,N_18677);
nor UO_1241 (O_1241,N_19609,N_19164);
and UO_1242 (O_1242,N_19401,N_18447);
nor UO_1243 (O_1243,N_18400,N_19952);
nor UO_1244 (O_1244,N_18790,N_18424);
nor UO_1245 (O_1245,N_19225,N_19661);
and UO_1246 (O_1246,N_18786,N_18344);
nand UO_1247 (O_1247,N_18525,N_18503);
nor UO_1248 (O_1248,N_19866,N_19198);
nor UO_1249 (O_1249,N_19415,N_19514);
or UO_1250 (O_1250,N_18423,N_19571);
or UO_1251 (O_1251,N_19535,N_18119);
nor UO_1252 (O_1252,N_19228,N_19518);
and UO_1253 (O_1253,N_18630,N_18567);
xnor UO_1254 (O_1254,N_18780,N_18535);
xnor UO_1255 (O_1255,N_19063,N_19214);
and UO_1256 (O_1256,N_18806,N_18616);
nor UO_1257 (O_1257,N_18479,N_19261);
or UO_1258 (O_1258,N_19338,N_18102);
or UO_1259 (O_1259,N_18390,N_18704);
nor UO_1260 (O_1260,N_18676,N_19437);
nor UO_1261 (O_1261,N_18414,N_19795);
nand UO_1262 (O_1262,N_19052,N_19663);
and UO_1263 (O_1263,N_18735,N_18395);
nand UO_1264 (O_1264,N_19492,N_19385);
xnor UO_1265 (O_1265,N_19571,N_18465);
nor UO_1266 (O_1266,N_19911,N_19179);
and UO_1267 (O_1267,N_18398,N_19602);
nand UO_1268 (O_1268,N_19401,N_19825);
or UO_1269 (O_1269,N_18066,N_19973);
nand UO_1270 (O_1270,N_18593,N_19192);
nand UO_1271 (O_1271,N_19633,N_18841);
or UO_1272 (O_1272,N_19236,N_18421);
and UO_1273 (O_1273,N_18974,N_18614);
or UO_1274 (O_1274,N_18781,N_19687);
and UO_1275 (O_1275,N_19878,N_19102);
nor UO_1276 (O_1276,N_18946,N_19431);
nand UO_1277 (O_1277,N_18932,N_18547);
nor UO_1278 (O_1278,N_19816,N_18707);
or UO_1279 (O_1279,N_18714,N_18362);
and UO_1280 (O_1280,N_19450,N_18452);
and UO_1281 (O_1281,N_19841,N_19809);
xor UO_1282 (O_1282,N_18196,N_19670);
xnor UO_1283 (O_1283,N_19244,N_19140);
or UO_1284 (O_1284,N_18330,N_19683);
or UO_1285 (O_1285,N_19680,N_18418);
xnor UO_1286 (O_1286,N_18083,N_19847);
and UO_1287 (O_1287,N_18769,N_19243);
nand UO_1288 (O_1288,N_19551,N_19678);
or UO_1289 (O_1289,N_19402,N_18258);
nor UO_1290 (O_1290,N_19352,N_19779);
nor UO_1291 (O_1291,N_19577,N_19641);
xor UO_1292 (O_1292,N_18526,N_18641);
and UO_1293 (O_1293,N_18882,N_18570);
or UO_1294 (O_1294,N_18531,N_19293);
or UO_1295 (O_1295,N_18503,N_19002);
nand UO_1296 (O_1296,N_18191,N_18476);
nor UO_1297 (O_1297,N_18756,N_19703);
or UO_1298 (O_1298,N_18544,N_18642);
nand UO_1299 (O_1299,N_19968,N_19982);
nand UO_1300 (O_1300,N_19352,N_18982);
and UO_1301 (O_1301,N_19393,N_18848);
or UO_1302 (O_1302,N_18655,N_18088);
nand UO_1303 (O_1303,N_18739,N_19337);
or UO_1304 (O_1304,N_18369,N_18829);
nand UO_1305 (O_1305,N_19267,N_18242);
and UO_1306 (O_1306,N_19059,N_19830);
and UO_1307 (O_1307,N_19233,N_19228);
or UO_1308 (O_1308,N_19320,N_19959);
xnor UO_1309 (O_1309,N_19099,N_18590);
nand UO_1310 (O_1310,N_19894,N_18124);
and UO_1311 (O_1311,N_19335,N_18506);
nor UO_1312 (O_1312,N_18000,N_19425);
nor UO_1313 (O_1313,N_18312,N_18932);
nor UO_1314 (O_1314,N_18964,N_19977);
or UO_1315 (O_1315,N_18404,N_18402);
nand UO_1316 (O_1316,N_18621,N_19771);
nand UO_1317 (O_1317,N_18394,N_19401);
xor UO_1318 (O_1318,N_19668,N_19231);
nor UO_1319 (O_1319,N_18190,N_19976);
nor UO_1320 (O_1320,N_18752,N_18974);
nand UO_1321 (O_1321,N_19233,N_18422);
nor UO_1322 (O_1322,N_18160,N_18013);
nor UO_1323 (O_1323,N_19422,N_18361);
and UO_1324 (O_1324,N_18702,N_18297);
or UO_1325 (O_1325,N_18705,N_18416);
nor UO_1326 (O_1326,N_18632,N_18824);
nor UO_1327 (O_1327,N_18174,N_18298);
and UO_1328 (O_1328,N_18441,N_18072);
nand UO_1329 (O_1329,N_18869,N_19055);
nor UO_1330 (O_1330,N_18156,N_19139);
or UO_1331 (O_1331,N_18452,N_19485);
or UO_1332 (O_1332,N_18893,N_19082);
nand UO_1333 (O_1333,N_19409,N_18320);
xnor UO_1334 (O_1334,N_18900,N_18087);
nor UO_1335 (O_1335,N_19200,N_18355);
and UO_1336 (O_1336,N_18589,N_19941);
nand UO_1337 (O_1337,N_18223,N_19137);
nand UO_1338 (O_1338,N_19308,N_19859);
nand UO_1339 (O_1339,N_18971,N_19475);
and UO_1340 (O_1340,N_18781,N_19085);
nor UO_1341 (O_1341,N_19141,N_18250);
nor UO_1342 (O_1342,N_18157,N_18617);
or UO_1343 (O_1343,N_19483,N_19969);
nor UO_1344 (O_1344,N_18074,N_19672);
or UO_1345 (O_1345,N_18851,N_19624);
or UO_1346 (O_1346,N_18698,N_19948);
nand UO_1347 (O_1347,N_19679,N_19875);
nand UO_1348 (O_1348,N_18420,N_19689);
and UO_1349 (O_1349,N_18517,N_18669);
nor UO_1350 (O_1350,N_18221,N_19443);
nand UO_1351 (O_1351,N_18758,N_18262);
or UO_1352 (O_1352,N_18636,N_19369);
and UO_1353 (O_1353,N_19828,N_18144);
nor UO_1354 (O_1354,N_18674,N_18787);
nor UO_1355 (O_1355,N_18252,N_19874);
nor UO_1356 (O_1356,N_18210,N_18280);
or UO_1357 (O_1357,N_18546,N_18951);
nand UO_1358 (O_1358,N_19949,N_18611);
nor UO_1359 (O_1359,N_19957,N_19093);
xnor UO_1360 (O_1360,N_19489,N_18387);
nor UO_1361 (O_1361,N_19153,N_19804);
nor UO_1362 (O_1362,N_19812,N_19793);
or UO_1363 (O_1363,N_19759,N_19495);
nor UO_1364 (O_1364,N_18447,N_19902);
and UO_1365 (O_1365,N_18098,N_19292);
and UO_1366 (O_1366,N_18417,N_18571);
or UO_1367 (O_1367,N_19416,N_19658);
nand UO_1368 (O_1368,N_19867,N_19520);
or UO_1369 (O_1369,N_18417,N_19433);
and UO_1370 (O_1370,N_18500,N_18177);
nor UO_1371 (O_1371,N_18777,N_18780);
nor UO_1372 (O_1372,N_19239,N_19950);
or UO_1373 (O_1373,N_18129,N_18941);
or UO_1374 (O_1374,N_18417,N_19248);
nand UO_1375 (O_1375,N_19152,N_18673);
xor UO_1376 (O_1376,N_19469,N_18789);
nor UO_1377 (O_1377,N_19813,N_19517);
and UO_1378 (O_1378,N_18505,N_19492);
nor UO_1379 (O_1379,N_18398,N_18409);
nand UO_1380 (O_1380,N_18932,N_19059);
and UO_1381 (O_1381,N_19494,N_18748);
nor UO_1382 (O_1382,N_19737,N_18112);
or UO_1383 (O_1383,N_19566,N_18291);
and UO_1384 (O_1384,N_19109,N_19267);
nand UO_1385 (O_1385,N_19502,N_18839);
nand UO_1386 (O_1386,N_19716,N_18479);
and UO_1387 (O_1387,N_18788,N_18919);
nand UO_1388 (O_1388,N_18367,N_19222);
or UO_1389 (O_1389,N_18009,N_18144);
nor UO_1390 (O_1390,N_19185,N_19814);
or UO_1391 (O_1391,N_19995,N_18380);
nand UO_1392 (O_1392,N_19407,N_19032);
nor UO_1393 (O_1393,N_18757,N_18632);
nor UO_1394 (O_1394,N_19735,N_19396);
nand UO_1395 (O_1395,N_19378,N_18152);
or UO_1396 (O_1396,N_19030,N_19755);
xnor UO_1397 (O_1397,N_18847,N_18474);
nand UO_1398 (O_1398,N_19205,N_18993);
or UO_1399 (O_1399,N_19755,N_19728);
or UO_1400 (O_1400,N_18680,N_18085);
or UO_1401 (O_1401,N_19286,N_18437);
xor UO_1402 (O_1402,N_19121,N_19512);
nand UO_1403 (O_1403,N_18266,N_19443);
nor UO_1404 (O_1404,N_19457,N_19381);
nand UO_1405 (O_1405,N_19293,N_19434);
nand UO_1406 (O_1406,N_19048,N_19126);
and UO_1407 (O_1407,N_19155,N_19552);
xnor UO_1408 (O_1408,N_19787,N_19402);
or UO_1409 (O_1409,N_18576,N_18963);
and UO_1410 (O_1410,N_19942,N_19710);
or UO_1411 (O_1411,N_18435,N_19189);
xor UO_1412 (O_1412,N_19256,N_19381);
and UO_1413 (O_1413,N_18286,N_19881);
nand UO_1414 (O_1414,N_19624,N_18169);
nor UO_1415 (O_1415,N_19649,N_19581);
or UO_1416 (O_1416,N_19470,N_19789);
and UO_1417 (O_1417,N_19456,N_18955);
or UO_1418 (O_1418,N_18452,N_19742);
or UO_1419 (O_1419,N_18823,N_18802);
nor UO_1420 (O_1420,N_19439,N_18261);
or UO_1421 (O_1421,N_18388,N_19417);
nand UO_1422 (O_1422,N_18844,N_19648);
nand UO_1423 (O_1423,N_19348,N_18339);
xnor UO_1424 (O_1424,N_19822,N_19295);
and UO_1425 (O_1425,N_18217,N_18408);
or UO_1426 (O_1426,N_19832,N_18155);
nor UO_1427 (O_1427,N_18069,N_19889);
and UO_1428 (O_1428,N_19742,N_19712);
or UO_1429 (O_1429,N_19731,N_19399);
nor UO_1430 (O_1430,N_19542,N_18255);
or UO_1431 (O_1431,N_18982,N_19153);
nand UO_1432 (O_1432,N_18334,N_19060);
and UO_1433 (O_1433,N_18165,N_18332);
nor UO_1434 (O_1434,N_18450,N_19517);
nor UO_1435 (O_1435,N_18540,N_19815);
and UO_1436 (O_1436,N_18360,N_18981);
xnor UO_1437 (O_1437,N_18968,N_18791);
and UO_1438 (O_1438,N_18917,N_18435);
and UO_1439 (O_1439,N_19586,N_18375);
nor UO_1440 (O_1440,N_18225,N_18900);
and UO_1441 (O_1441,N_18615,N_19081);
or UO_1442 (O_1442,N_18049,N_19493);
nor UO_1443 (O_1443,N_18851,N_19484);
nand UO_1444 (O_1444,N_19525,N_19750);
nor UO_1445 (O_1445,N_18771,N_19373);
nor UO_1446 (O_1446,N_18909,N_18379);
or UO_1447 (O_1447,N_19477,N_19191);
or UO_1448 (O_1448,N_19676,N_19719);
and UO_1449 (O_1449,N_19289,N_19611);
nor UO_1450 (O_1450,N_19682,N_18418);
xor UO_1451 (O_1451,N_18592,N_19788);
nand UO_1452 (O_1452,N_19653,N_18031);
or UO_1453 (O_1453,N_18214,N_18061);
nand UO_1454 (O_1454,N_18326,N_19048);
nand UO_1455 (O_1455,N_19294,N_18773);
nor UO_1456 (O_1456,N_19540,N_19789);
nor UO_1457 (O_1457,N_19905,N_18031);
nand UO_1458 (O_1458,N_19645,N_18792);
and UO_1459 (O_1459,N_18032,N_18989);
and UO_1460 (O_1460,N_18337,N_19089);
or UO_1461 (O_1461,N_18794,N_19314);
nand UO_1462 (O_1462,N_19107,N_19851);
nand UO_1463 (O_1463,N_19315,N_19798);
or UO_1464 (O_1464,N_19900,N_18246);
xnor UO_1465 (O_1465,N_19543,N_18202);
nand UO_1466 (O_1466,N_19222,N_19113);
and UO_1467 (O_1467,N_19726,N_18801);
nand UO_1468 (O_1468,N_18400,N_18342);
nor UO_1469 (O_1469,N_18785,N_18685);
or UO_1470 (O_1470,N_19386,N_19596);
nand UO_1471 (O_1471,N_19284,N_19567);
and UO_1472 (O_1472,N_18866,N_18622);
nor UO_1473 (O_1473,N_19762,N_19441);
and UO_1474 (O_1474,N_18507,N_18006);
nand UO_1475 (O_1475,N_19217,N_19330);
and UO_1476 (O_1476,N_18861,N_19752);
nor UO_1477 (O_1477,N_18926,N_19296);
or UO_1478 (O_1478,N_19190,N_19752);
nand UO_1479 (O_1479,N_19287,N_18709);
or UO_1480 (O_1480,N_18640,N_19431);
nor UO_1481 (O_1481,N_19642,N_18185);
nand UO_1482 (O_1482,N_18279,N_19256);
nor UO_1483 (O_1483,N_19075,N_18853);
nor UO_1484 (O_1484,N_18750,N_19097);
nand UO_1485 (O_1485,N_19221,N_19241);
nand UO_1486 (O_1486,N_19424,N_18903);
nor UO_1487 (O_1487,N_19795,N_19023);
nand UO_1488 (O_1488,N_18888,N_18502);
nand UO_1489 (O_1489,N_19487,N_19646);
xor UO_1490 (O_1490,N_18714,N_19848);
or UO_1491 (O_1491,N_19990,N_19121);
nor UO_1492 (O_1492,N_18839,N_18783);
and UO_1493 (O_1493,N_18418,N_19136);
and UO_1494 (O_1494,N_19043,N_18086);
or UO_1495 (O_1495,N_18433,N_19969);
xnor UO_1496 (O_1496,N_18975,N_18793);
nor UO_1497 (O_1497,N_18125,N_18241);
nand UO_1498 (O_1498,N_19808,N_18842);
nand UO_1499 (O_1499,N_18869,N_19918);
nor UO_1500 (O_1500,N_19551,N_18798);
or UO_1501 (O_1501,N_18452,N_18454);
and UO_1502 (O_1502,N_18311,N_19515);
nand UO_1503 (O_1503,N_19965,N_18932);
or UO_1504 (O_1504,N_19045,N_19303);
and UO_1505 (O_1505,N_19883,N_18589);
nand UO_1506 (O_1506,N_18582,N_19294);
nor UO_1507 (O_1507,N_18019,N_19614);
nand UO_1508 (O_1508,N_19189,N_19941);
and UO_1509 (O_1509,N_19206,N_19574);
nand UO_1510 (O_1510,N_19199,N_18982);
or UO_1511 (O_1511,N_19157,N_18181);
or UO_1512 (O_1512,N_18541,N_18719);
nand UO_1513 (O_1513,N_19658,N_18600);
or UO_1514 (O_1514,N_18218,N_19871);
nand UO_1515 (O_1515,N_19539,N_19532);
or UO_1516 (O_1516,N_18493,N_18527);
nor UO_1517 (O_1517,N_18370,N_19877);
xor UO_1518 (O_1518,N_19880,N_18994);
and UO_1519 (O_1519,N_18095,N_19356);
nor UO_1520 (O_1520,N_18149,N_19792);
nor UO_1521 (O_1521,N_18761,N_18691);
and UO_1522 (O_1522,N_18403,N_18502);
nor UO_1523 (O_1523,N_19693,N_18765);
or UO_1524 (O_1524,N_19126,N_18526);
nand UO_1525 (O_1525,N_18536,N_19610);
nor UO_1526 (O_1526,N_19192,N_19489);
or UO_1527 (O_1527,N_19801,N_19811);
or UO_1528 (O_1528,N_19230,N_19949);
nor UO_1529 (O_1529,N_18282,N_19123);
and UO_1530 (O_1530,N_19425,N_18895);
nand UO_1531 (O_1531,N_18290,N_19243);
nor UO_1532 (O_1532,N_19220,N_19016);
nand UO_1533 (O_1533,N_19313,N_19281);
xor UO_1534 (O_1534,N_19885,N_18831);
or UO_1535 (O_1535,N_18152,N_18510);
and UO_1536 (O_1536,N_18939,N_19047);
nor UO_1537 (O_1537,N_19319,N_19775);
or UO_1538 (O_1538,N_19773,N_19810);
nor UO_1539 (O_1539,N_19227,N_18861);
and UO_1540 (O_1540,N_19778,N_18589);
nor UO_1541 (O_1541,N_18633,N_18093);
xnor UO_1542 (O_1542,N_19231,N_18708);
or UO_1543 (O_1543,N_19736,N_18317);
xor UO_1544 (O_1544,N_18235,N_19581);
and UO_1545 (O_1545,N_18066,N_18334);
and UO_1546 (O_1546,N_18751,N_18694);
nor UO_1547 (O_1547,N_19397,N_18875);
nand UO_1548 (O_1548,N_18492,N_19028);
and UO_1549 (O_1549,N_19655,N_19878);
or UO_1550 (O_1550,N_19265,N_19843);
and UO_1551 (O_1551,N_18395,N_19482);
nor UO_1552 (O_1552,N_19052,N_18991);
nand UO_1553 (O_1553,N_18413,N_18123);
nor UO_1554 (O_1554,N_19369,N_18727);
and UO_1555 (O_1555,N_19435,N_19071);
nand UO_1556 (O_1556,N_19854,N_18837);
and UO_1557 (O_1557,N_19313,N_19896);
xor UO_1558 (O_1558,N_18087,N_18536);
xor UO_1559 (O_1559,N_18397,N_18817);
or UO_1560 (O_1560,N_19104,N_19703);
and UO_1561 (O_1561,N_19614,N_19497);
nand UO_1562 (O_1562,N_19359,N_19945);
and UO_1563 (O_1563,N_18086,N_19837);
nor UO_1564 (O_1564,N_19346,N_19153);
nor UO_1565 (O_1565,N_19766,N_18104);
or UO_1566 (O_1566,N_19956,N_18211);
or UO_1567 (O_1567,N_19306,N_18086);
or UO_1568 (O_1568,N_18802,N_19619);
and UO_1569 (O_1569,N_19576,N_18152);
nor UO_1570 (O_1570,N_18485,N_18593);
or UO_1571 (O_1571,N_18539,N_18232);
and UO_1572 (O_1572,N_19947,N_19917);
nor UO_1573 (O_1573,N_19597,N_19869);
nor UO_1574 (O_1574,N_19271,N_19540);
nand UO_1575 (O_1575,N_19518,N_18999);
and UO_1576 (O_1576,N_18768,N_18355);
or UO_1577 (O_1577,N_19542,N_18788);
nor UO_1578 (O_1578,N_18570,N_18108);
nand UO_1579 (O_1579,N_18969,N_18707);
and UO_1580 (O_1580,N_19593,N_18113);
nand UO_1581 (O_1581,N_19490,N_19226);
nand UO_1582 (O_1582,N_18620,N_18848);
nand UO_1583 (O_1583,N_18364,N_18325);
or UO_1584 (O_1584,N_19402,N_19206);
nor UO_1585 (O_1585,N_18988,N_19167);
nand UO_1586 (O_1586,N_18463,N_19797);
nor UO_1587 (O_1587,N_18124,N_18338);
or UO_1588 (O_1588,N_18584,N_18678);
nand UO_1589 (O_1589,N_18313,N_18211);
and UO_1590 (O_1590,N_19721,N_18627);
or UO_1591 (O_1591,N_18790,N_18703);
and UO_1592 (O_1592,N_18962,N_19908);
and UO_1593 (O_1593,N_19276,N_19070);
or UO_1594 (O_1594,N_18664,N_18216);
or UO_1595 (O_1595,N_18908,N_18971);
and UO_1596 (O_1596,N_19486,N_19306);
and UO_1597 (O_1597,N_18508,N_19534);
nand UO_1598 (O_1598,N_18274,N_19677);
or UO_1599 (O_1599,N_19122,N_18510);
nand UO_1600 (O_1600,N_19191,N_19189);
and UO_1601 (O_1601,N_18506,N_18809);
and UO_1602 (O_1602,N_18518,N_19124);
nor UO_1603 (O_1603,N_19284,N_19089);
xor UO_1604 (O_1604,N_18753,N_19979);
nor UO_1605 (O_1605,N_18553,N_19626);
nor UO_1606 (O_1606,N_18812,N_19024);
xnor UO_1607 (O_1607,N_18391,N_19296);
nor UO_1608 (O_1608,N_18873,N_19694);
and UO_1609 (O_1609,N_18537,N_18257);
xor UO_1610 (O_1610,N_19175,N_18217);
or UO_1611 (O_1611,N_18454,N_18112);
xor UO_1612 (O_1612,N_18022,N_19577);
nand UO_1613 (O_1613,N_18399,N_18454);
nand UO_1614 (O_1614,N_18668,N_18605);
and UO_1615 (O_1615,N_19595,N_19457);
and UO_1616 (O_1616,N_18706,N_19185);
nor UO_1617 (O_1617,N_18807,N_18157);
nand UO_1618 (O_1618,N_18558,N_18483);
and UO_1619 (O_1619,N_19474,N_18966);
xor UO_1620 (O_1620,N_19187,N_18326);
and UO_1621 (O_1621,N_18043,N_19205);
nor UO_1622 (O_1622,N_18459,N_19253);
nand UO_1623 (O_1623,N_19521,N_18890);
or UO_1624 (O_1624,N_18835,N_18671);
nor UO_1625 (O_1625,N_18103,N_18959);
or UO_1626 (O_1626,N_19931,N_18270);
nor UO_1627 (O_1627,N_18327,N_19633);
nor UO_1628 (O_1628,N_19930,N_18084);
nand UO_1629 (O_1629,N_19830,N_18824);
or UO_1630 (O_1630,N_19804,N_19397);
nand UO_1631 (O_1631,N_19565,N_18655);
xnor UO_1632 (O_1632,N_19865,N_19074);
nand UO_1633 (O_1633,N_18973,N_19149);
and UO_1634 (O_1634,N_18486,N_18498);
or UO_1635 (O_1635,N_19566,N_18805);
or UO_1636 (O_1636,N_19126,N_19294);
and UO_1637 (O_1637,N_18433,N_19298);
or UO_1638 (O_1638,N_18491,N_19714);
nor UO_1639 (O_1639,N_19700,N_19909);
xnor UO_1640 (O_1640,N_19250,N_18680);
or UO_1641 (O_1641,N_18170,N_19591);
nand UO_1642 (O_1642,N_18932,N_19295);
and UO_1643 (O_1643,N_18450,N_18715);
nor UO_1644 (O_1644,N_19066,N_19216);
xnor UO_1645 (O_1645,N_19458,N_18386);
nand UO_1646 (O_1646,N_19561,N_18671);
nand UO_1647 (O_1647,N_18970,N_19892);
xnor UO_1648 (O_1648,N_18501,N_19851);
nor UO_1649 (O_1649,N_19237,N_18642);
or UO_1650 (O_1650,N_19558,N_18625);
nand UO_1651 (O_1651,N_19177,N_19014);
nor UO_1652 (O_1652,N_19470,N_19075);
xor UO_1653 (O_1653,N_19916,N_18120);
nor UO_1654 (O_1654,N_19816,N_18784);
or UO_1655 (O_1655,N_18383,N_19544);
and UO_1656 (O_1656,N_19904,N_18143);
or UO_1657 (O_1657,N_18349,N_18573);
xnor UO_1658 (O_1658,N_19572,N_19225);
xor UO_1659 (O_1659,N_18681,N_18748);
or UO_1660 (O_1660,N_19344,N_19858);
and UO_1661 (O_1661,N_19903,N_18113);
nor UO_1662 (O_1662,N_19484,N_19672);
nor UO_1663 (O_1663,N_19118,N_19809);
and UO_1664 (O_1664,N_19127,N_18990);
nor UO_1665 (O_1665,N_18646,N_19882);
nor UO_1666 (O_1666,N_19687,N_19698);
nand UO_1667 (O_1667,N_19137,N_18837);
nor UO_1668 (O_1668,N_19482,N_18662);
or UO_1669 (O_1669,N_19293,N_18212);
nor UO_1670 (O_1670,N_19166,N_19609);
or UO_1671 (O_1671,N_18499,N_19394);
and UO_1672 (O_1672,N_18905,N_19170);
and UO_1673 (O_1673,N_19072,N_18362);
nand UO_1674 (O_1674,N_18609,N_19117);
or UO_1675 (O_1675,N_18712,N_19689);
nand UO_1676 (O_1676,N_18875,N_19336);
nor UO_1677 (O_1677,N_18909,N_19764);
or UO_1678 (O_1678,N_19370,N_18109);
and UO_1679 (O_1679,N_18643,N_19893);
or UO_1680 (O_1680,N_18558,N_19826);
and UO_1681 (O_1681,N_19760,N_18273);
nor UO_1682 (O_1682,N_19866,N_18687);
or UO_1683 (O_1683,N_18906,N_18769);
and UO_1684 (O_1684,N_19556,N_18131);
and UO_1685 (O_1685,N_18883,N_19952);
or UO_1686 (O_1686,N_19969,N_19821);
and UO_1687 (O_1687,N_18419,N_18155);
xnor UO_1688 (O_1688,N_18438,N_18820);
and UO_1689 (O_1689,N_18904,N_19670);
nor UO_1690 (O_1690,N_18364,N_18241);
and UO_1691 (O_1691,N_19496,N_19470);
nand UO_1692 (O_1692,N_18717,N_18357);
nor UO_1693 (O_1693,N_18774,N_18030);
or UO_1694 (O_1694,N_19505,N_18396);
nand UO_1695 (O_1695,N_18065,N_18671);
or UO_1696 (O_1696,N_18534,N_19141);
nand UO_1697 (O_1697,N_19149,N_18125);
nor UO_1698 (O_1698,N_19718,N_19173);
and UO_1699 (O_1699,N_19652,N_18983);
nand UO_1700 (O_1700,N_18008,N_18732);
or UO_1701 (O_1701,N_19905,N_18841);
and UO_1702 (O_1702,N_19397,N_19251);
nand UO_1703 (O_1703,N_19666,N_19471);
nand UO_1704 (O_1704,N_18599,N_18896);
nand UO_1705 (O_1705,N_18379,N_19853);
and UO_1706 (O_1706,N_19662,N_18437);
nand UO_1707 (O_1707,N_19356,N_18691);
nor UO_1708 (O_1708,N_18592,N_18910);
and UO_1709 (O_1709,N_18126,N_18256);
nand UO_1710 (O_1710,N_18228,N_19011);
nor UO_1711 (O_1711,N_19882,N_19080);
xor UO_1712 (O_1712,N_18514,N_18893);
and UO_1713 (O_1713,N_18116,N_18046);
nor UO_1714 (O_1714,N_19501,N_18881);
nand UO_1715 (O_1715,N_19237,N_19663);
and UO_1716 (O_1716,N_18390,N_19998);
and UO_1717 (O_1717,N_19997,N_19738);
nor UO_1718 (O_1718,N_18009,N_18115);
nand UO_1719 (O_1719,N_18495,N_19107);
or UO_1720 (O_1720,N_19687,N_19571);
nor UO_1721 (O_1721,N_19587,N_19548);
or UO_1722 (O_1722,N_18454,N_18062);
nand UO_1723 (O_1723,N_18493,N_19246);
nand UO_1724 (O_1724,N_18760,N_19692);
or UO_1725 (O_1725,N_18640,N_19466);
xor UO_1726 (O_1726,N_18112,N_19586);
or UO_1727 (O_1727,N_19538,N_19303);
nor UO_1728 (O_1728,N_18359,N_18774);
or UO_1729 (O_1729,N_18079,N_19129);
and UO_1730 (O_1730,N_19986,N_18458);
nor UO_1731 (O_1731,N_19619,N_19616);
nor UO_1732 (O_1732,N_19174,N_18718);
and UO_1733 (O_1733,N_19583,N_18680);
nand UO_1734 (O_1734,N_19852,N_19243);
nor UO_1735 (O_1735,N_18757,N_18930);
xor UO_1736 (O_1736,N_19984,N_18433);
nand UO_1737 (O_1737,N_18288,N_19464);
nor UO_1738 (O_1738,N_18397,N_19188);
and UO_1739 (O_1739,N_19225,N_19037);
nor UO_1740 (O_1740,N_18569,N_19673);
nand UO_1741 (O_1741,N_19742,N_18773);
and UO_1742 (O_1742,N_19743,N_18913);
nand UO_1743 (O_1743,N_19358,N_19693);
nor UO_1744 (O_1744,N_19716,N_18116);
nand UO_1745 (O_1745,N_18756,N_18343);
or UO_1746 (O_1746,N_18775,N_18591);
or UO_1747 (O_1747,N_19589,N_18655);
nand UO_1748 (O_1748,N_18529,N_19566);
nor UO_1749 (O_1749,N_18058,N_18492);
or UO_1750 (O_1750,N_18582,N_19653);
nand UO_1751 (O_1751,N_19878,N_19854);
and UO_1752 (O_1752,N_18787,N_18640);
nand UO_1753 (O_1753,N_19088,N_19745);
nand UO_1754 (O_1754,N_18289,N_18132);
and UO_1755 (O_1755,N_19139,N_19862);
or UO_1756 (O_1756,N_19442,N_19837);
nand UO_1757 (O_1757,N_19577,N_18128);
nor UO_1758 (O_1758,N_18312,N_19288);
nand UO_1759 (O_1759,N_18734,N_19893);
nor UO_1760 (O_1760,N_19358,N_18938);
xor UO_1761 (O_1761,N_19147,N_19159);
nor UO_1762 (O_1762,N_18439,N_19280);
and UO_1763 (O_1763,N_19257,N_18459);
nand UO_1764 (O_1764,N_19194,N_18893);
nand UO_1765 (O_1765,N_19584,N_18193);
nand UO_1766 (O_1766,N_19306,N_19174);
nor UO_1767 (O_1767,N_18883,N_19355);
and UO_1768 (O_1768,N_18698,N_18328);
or UO_1769 (O_1769,N_19902,N_19692);
nand UO_1770 (O_1770,N_18924,N_18416);
nand UO_1771 (O_1771,N_19077,N_19715);
nand UO_1772 (O_1772,N_18416,N_18564);
nor UO_1773 (O_1773,N_19332,N_19442);
nand UO_1774 (O_1774,N_19181,N_18804);
and UO_1775 (O_1775,N_19238,N_18354);
and UO_1776 (O_1776,N_18283,N_19490);
nand UO_1777 (O_1777,N_19949,N_19405);
nand UO_1778 (O_1778,N_19653,N_18283);
nor UO_1779 (O_1779,N_19695,N_19955);
or UO_1780 (O_1780,N_18032,N_18073);
and UO_1781 (O_1781,N_18096,N_18305);
and UO_1782 (O_1782,N_19111,N_18643);
and UO_1783 (O_1783,N_19535,N_19170);
or UO_1784 (O_1784,N_19833,N_18795);
or UO_1785 (O_1785,N_19014,N_19755);
or UO_1786 (O_1786,N_18359,N_19545);
nand UO_1787 (O_1787,N_18775,N_19060);
nor UO_1788 (O_1788,N_19339,N_18821);
or UO_1789 (O_1789,N_19034,N_19508);
nor UO_1790 (O_1790,N_19735,N_19462);
nand UO_1791 (O_1791,N_19911,N_19383);
and UO_1792 (O_1792,N_19244,N_18996);
nand UO_1793 (O_1793,N_18639,N_19513);
or UO_1794 (O_1794,N_18304,N_19623);
xnor UO_1795 (O_1795,N_18656,N_18235);
nor UO_1796 (O_1796,N_19186,N_19723);
xnor UO_1797 (O_1797,N_19557,N_19162);
and UO_1798 (O_1798,N_19233,N_18802);
and UO_1799 (O_1799,N_19742,N_18328);
or UO_1800 (O_1800,N_18203,N_18915);
and UO_1801 (O_1801,N_18658,N_18202);
nand UO_1802 (O_1802,N_19324,N_18169);
and UO_1803 (O_1803,N_18483,N_19657);
nand UO_1804 (O_1804,N_19780,N_18685);
or UO_1805 (O_1805,N_19954,N_18876);
and UO_1806 (O_1806,N_19194,N_18612);
nand UO_1807 (O_1807,N_19811,N_19835);
or UO_1808 (O_1808,N_18274,N_18634);
and UO_1809 (O_1809,N_19214,N_18043);
or UO_1810 (O_1810,N_18675,N_18967);
or UO_1811 (O_1811,N_18663,N_18191);
and UO_1812 (O_1812,N_18972,N_19061);
or UO_1813 (O_1813,N_19754,N_19505);
and UO_1814 (O_1814,N_18819,N_19432);
or UO_1815 (O_1815,N_18310,N_18027);
nand UO_1816 (O_1816,N_18870,N_19823);
and UO_1817 (O_1817,N_19537,N_18103);
and UO_1818 (O_1818,N_19904,N_18140);
or UO_1819 (O_1819,N_18674,N_18214);
nand UO_1820 (O_1820,N_18549,N_18494);
or UO_1821 (O_1821,N_18446,N_19874);
or UO_1822 (O_1822,N_18650,N_19740);
and UO_1823 (O_1823,N_18716,N_19269);
and UO_1824 (O_1824,N_19066,N_19105);
or UO_1825 (O_1825,N_19588,N_19213);
or UO_1826 (O_1826,N_18954,N_19413);
nor UO_1827 (O_1827,N_18164,N_19362);
xnor UO_1828 (O_1828,N_19118,N_19666);
or UO_1829 (O_1829,N_18053,N_18932);
or UO_1830 (O_1830,N_18528,N_18423);
nor UO_1831 (O_1831,N_19149,N_18557);
xor UO_1832 (O_1832,N_18740,N_19744);
xnor UO_1833 (O_1833,N_19737,N_19378);
and UO_1834 (O_1834,N_18735,N_19100);
and UO_1835 (O_1835,N_19812,N_18814);
xnor UO_1836 (O_1836,N_18706,N_19417);
xnor UO_1837 (O_1837,N_19374,N_19085);
nand UO_1838 (O_1838,N_19300,N_18180);
or UO_1839 (O_1839,N_19105,N_18037);
or UO_1840 (O_1840,N_19793,N_18423);
and UO_1841 (O_1841,N_18106,N_18595);
and UO_1842 (O_1842,N_19482,N_18218);
xnor UO_1843 (O_1843,N_18776,N_18492);
nand UO_1844 (O_1844,N_18633,N_19583);
nor UO_1845 (O_1845,N_18784,N_18055);
nand UO_1846 (O_1846,N_19686,N_18848);
and UO_1847 (O_1847,N_18623,N_18669);
and UO_1848 (O_1848,N_18931,N_19739);
or UO_1849 (O_1849,N_19434,N_19974);
nand UO_1850 (O_1850,N_19088,N_19618);
nand UO_1851 (O_1851,N_18667,N_19348);
nand UO_1852 (O_1852,N_19111,N_19509);
and UO_1853 (O_1853,N_19248,N_19644);
xnor UO_1854 (O_1854,N_19207,N_19258);
and UO_1855 (O_1855,N_19400,N_18827);
nand UO_1856 (O_1856,N_19018,N_18122);
nand UO_1857 (O_1857,N_18667,N_18278);
nor UO_1858 (O_1858,N_19228,N_19018);
xnor UO_1859 (O_1859,N_19669,N_19355);
nand UO_1860 (O_1860,N_18334,N_19070);
nor UO_1861 (O_1861,N_18629,N_19901);
and UO_1862 (O_1862,N_19613,N_18946);
or UO_1863 (O_1863,N_19552,N_19281);
and UO_1864 (O_1864,N_19629,N_18015);
nand UO_1865 (O_1865,N_18969,N_18718);
xnor UO_1866 (O_1866,N_19879,N_18945);
nor UO_1867 (O_1867,N_19730,N_19162);
nand UO_1868 (O_1868,N_18697,N_18516);
xnor UO_1869 (O_1869,N_18800,N_19581);
xnor UO_1870 (O_1870,N_18495,N_18395);
nor UO_1871 (O_1871,N_18941,N_19512);
nor UO_1872 (O_1872,N_18582,N_18068);
and UO_1873 (O_1873,N_18157,N_19322);
and UO_1874 (O_1874,N_19145,N_18935);
or UO_1875 (O_1875,N_19667,N_19875);
nand UO_1876 (O_1876,N_18170,N_19558);
nor UO_1877 (O_1877,N_18543,N_18010);
xnor UO_1878 (O_1878,N_18025,N_18827);
and UO_1879 (O_1879,N_19417,N_18951);
nand UO_1880 (O_1880,N_18570,N_19479);
and UO_1881 (O_1881,N_18926,N_18454);
nand UO_1882 (O_1882,N_18477,N_18475);
nor UO_1883 (O_1883,N_19357,N_18189);
or UO_1884 (O_1884,N_18359,N_19441);
and UO_1885 (O_1885,N_18543,N_18782);
and UO_1886 (O_1886,N_19935,N_18439);
nor UO_1887 (O_1887,N_19047,N_18599);
nor UO_1888 (O_1888,N_19852,N_18267);
nor UO_1889 (O_1889,N_19315,N_18640);
nand UO_1890 (O_1890,N_18336,N_18445);
or UO_1891 (O_1891,N_18500,N_19936);
or UO_1892 (O_1892,N_18613,N_18660);
and UO_1893 (O_1893,N_18713,N_18718);
or UO_1894 (O_1894,N_18310,N_18450);
or UO_1895 (O_1895,N_18412,N_18456);
xnor UO_1896 (O_1896,N_18486,N_18055);
or UO_1897 (O_1897,N_18135,N_19545);
nand UO_1898 (O_1898,N_18831,N_18939);
xnor UO_1899 (O_1899,N_18485,N_18934);
nor UO_1900 (O_1900,N_18164,N_19774);
nor UO_1901 (O_1901,N_18314,N_18218);
and UO_1902 (O_1902,N_19879,N_18482);
xnor UO_1903 (O_1903,N_18004,N_18641);
nor UO_1904 (O_1904,N_18761,N_18499);
and UO_1905 (O_1905,N_18396,N_18134);
nor UO_1906 (O_1906,N_18975,N_19733);
or UO_1907 (O_1907,N_18363,N_18511);
or UO_1908 (O_1908,N_18545,N_18639);
xnor UO_1909 (O_1909,N_19223,N_18861);
and UO_1910 (O_1910,N_19482,N_19921);
nand UO_1911 (O_1911,N_19695,N_18582);
or UO_1912 (O_1912,N_19973,N_18316);
and UO_1913 (O_1913,N_19451,N_18877);
and UO_1914 (O_1914,N_18873,N_19689);
and UO_1915 (O_1915,N_18977,N_19703);
nand UO_1916 (O_1916,N_19266,N_19231);
or UO_1917 (O_1917,N_18133,N_19823);
nor UO_1918 (O_1918,N_19544,N_19012);
nand UO_1919 (O_1919,N_19410,N_19397);
nor UO_1920 (O_1920,N_18245,N_19643);
and UO_1921 (O_1921,N_18732,N_19201);
or UO_1922 (O_1922,N_19596,N_18142);
and UO_1923 (O_1923,N_18600,N_19748);
nor UO_1924 (O_1924,N_19659,N_18067);
or UO_1925 (O_1925,N_19562,N_18130);
nand UO_1926 (O_1926,N_18319,N_18629);
or UO_1927 (O_1927,N_18769,N_19013);
or UO_1928 (O_1928,N_19026,N_19084);
nor UO_1929 (O_1929,N_19675,N_19867);
and UO_1930 (O_1930,N_18773,N_19855);
nor UO_1931 (O_1931,N_19179,N_18732);
nand UO_1932 (O_1932,N_19728,N_18394);
and UO_1933 (O_1933,N_19967,N_18858);
and UO_1934 (O_1934,N_19881,N_19707);
and UO_1935 (O_1935,N_19275,N_18553);
nand UO_1936 (O_1936,N_18159,N_19165);
nor UO_1937 (O_1937,N_18920,N_19864);
and UO_1938 (O_1938,N_18492,N_18898);
nor UO_1939 (O_1939,N_19390,N_18340);
nor UO_1940 (O_1940,N_18033,N_19488);
and UO_1941 (O_1941,N_19390,N_18077);
or UO_1942 (O_1942,N_18555,N_19511);
and UO_1943 (O_1943,N_18136,N_18690);
xnor UO_1944 (O_1944,N_18906,N_18960);
or UO_1945 (O_1945,N_18526,N_18805);
or UO_1946 (O_1946,N_19499,N_19114);
xor UO_1947 (O_1947,N_18907,N_19995);
nand UO_1948 (O_1948,N_19534,N_19072);
or UO_1949 (O_1949,N_19688,N_18585);
nor UO_1950 (O_1950,N_18272,N_18888);
and UO_1951 (O_1951,N_19013,N_18647);
nor UO_1952 (O_1952,N_19157,N_18925);
or UO_1953 (O_1953,N_18206,N_18801);
nand UO_1954 (O_1954,N_18127,N_19483);
nor UO_1955 (O_1955,N_18410,N_19661);
or UO_1956 (O_1956,N_18580,N_19617);
nor UO_1957 (O_1957,N_19092,N_18096);
nand UO_1958 (O_1958,N_18558,N_18011);
or UO_1959 (O_1959,N_19425,N_19600);
nor UO_1960 (O_1960,N_19084,N_18654);
and UO_1961 (O_1961,N_19195,N_18098);
nor UO_1962 (O_1962,N_18628,N_19200);
nor UO_1963 (O_1963,N_19730,N_19621);
or UO_1964 (O_1964,N_18663,N_18002);
xnor UO_1965 (O_1965,N_18453,N_18439);
xnor UO_1966 (O_1966,N_18370,N_19609);
nor UO_1967 (O_1967,N_19594,N_18721);
nand UO_1968 (O_1968,N_19222,N_18954);
nor UO_1969 (O_1969,N_19920,N_19333);
and UO_1970 (O_1970,N_19275,N_18564);
or UO_1971 (O_1971,N_19298,N_19321);
nor UO_1972 (O_1972,N_19914,N_18435);
nor UO_1973 (O_1973,N_19784,N_19550);
or UO_1974 (O_1974,N_18834,N_19668);
and UO_1975 (O_1975,N_19692,N_18175);
or UO_1976 (O_1976,N_19175,N_18160);
nor UO_1977 (O_1977,N_19771,N_19122);
nor UO_1978 (O_1978,N_19096,N_19374);
nand UO_1979 (O_1979,N_19933,N_18564);
nor UO_1980 (O_1980,N_19182,N_18149);
or UO_1981 (O_1981,N_19635,N_18059);
nor UO_1982 (O_1982,N_19412,N_18336);
nor UO_1983 (O_1983,N_18063,N_18242);
nor UO_1984 (O_1984,N_18215,N_19719);
or UO_1985 (O_1985,N_18288,N_19984);
nand UO_1986 (O_1986,N_18010,N_18854);
nand UO_1987 (O_1987,N_18212,N_19976);
nor UO_1988 (O_1988,N_18782,N_18298);
nor UO_1989 (O_1989,N_18070,N_18898);
or UO_1990 (O_1990,N_18694,N_18829);
nor UO_1991 (O_1991,N_19883,N_19791);
nand UO_1992 (O_1992,N_19432,N_18230);
nand UO_1993 (O_1993,N_18901,N_19851);
nand UO_1994 (O_1994,N_19981,N_18453);
and UO_1995 (O_1995,N_18837,N_19307);
xnor UO_1996 (O_1996,N_18161,N_19599);
nand UO_1997 (O_1997,N_19242,N_18837);
nand UO_1998 (O_1998,N_19528,N_19135);
nor UO_1999 (O_1999,N_19891,N_19646);
nand UO_2000 (O_2000,N_18281,N_18664);
nand UO_2001 (O_2001,N_19886,N_19152);
and UO_2002 (O_2002,N_18471,N_18114);
nor UO_2003 (O_2003,N_19943,N_18258);
and UO_2004 (O_2004,N_19296,N_18852);
nand UO_2005 (O_2005,N_18930,N_19641);
and UO_2006 (O_2006,N_19494,N_19437);
or UO_2007 (O_2007,N_19644,N_19304);
nand UO_2008 (O_2008,N_19491,N_19218);
nand UO_2009 (O_2009,N_18454,N_19273);
nor UO_2010 (O_2010,N_18497,N_19666);
nor UO_2011 (O_2011,N_18492,N_19352);
or UO_2012 (O_2012,N_18382,N_18414);
nor UO_2013 (O_2013,N_18456,N_18979);
and UO_2014 (O_2014,N_18294,N_18950);
or UO_2015 (O_2015,N_18848,N_19672);
and UO_2016 (O_2016,N_18392,N_19091);
nor UO_2017 (O_2017,N_18921,N_19240);
xor UO_2018 (O_2018,N_19026,N_19926);
nand UO_2019 (O_2019,N_18786,N_19078);
and UO_2020 (O_2020,N_18125,N_19342);
or UO_2021 (O_2021,N_18531,N_19409);
nand UO_2022 (O_2022,N_19696,N_18083);
and UO_2023 (O_2023,N_18612,N_18507);
and UO_2024 (O_2024,N_18446,N_19880);
xnor UO_2025 (O_2025,N_19766,N_18334);
xnor UO_2026 (O_2026,N_19597,N_19732);
nor UO_2027 (O_2027,N_18544,N_19213);
xnor UO_2028 (O_2028,N_19329,N_18863);
or UO_2029 (O_2029,N_18259,N_18873);
and UO_2030 (O_2030,N_18526,N_19314);
nor UO_2031 (O_2031,N_18229,N_19453);
and UO_2032 (O_2032,N_19652,N_18697);
nor UO_2033 (O_2033,N_19299,N_18520);
and UO_2034 (O_2034,N_18074,N_18038);
or UO_2035 (O_2035,N_18649,N_18587);
and UO_2036 (O_2036,N_18817,N_18796);
xor UO_2037 (O_2037,N_18565,N_18197);
nor UO_2038 (O_2038,N_19292,N_19825);
and UO_2039 (O_2039,N_18641,N_18914);
or UO_2040 (O_2040,N_18049,N_19865);
or UO_2041 (O_2041,N_18470,N_19586);
or UO_2042 (O_2042,N_19323,N_19139);
nand UO_2043 (O_2043,N_19540,N_18350);
and UO_2044 (O_2044,N_18540,N_19691);
nor UO_2045 (O_2045,N_18820,N_19166);
nor UO_2046 (O_2046,N_18823,N_19166);
nor UO_2047 (O_2047,N_18378,N_19849);
nand UO_2048 (O_2048,N_19975,N_19959);
nand UO_2049 (O_2049,N_19008,N_18319);
or UO_2050 (O_2050,N_18626,N_18748);
or UO_2051 (O_2051,N_18439,N_19621);
nor UO_2052 (O_2052,N_19062,N_19351);
or UO_2053 (O_2053,N_19236,N_19444);
or UO_2054 (O_2054,N_18952,N_19357);
nor UO_2055 (O_2055,N_18473,N_18601);
or UO_2056 (O_2056,N_18523,N_18368);
and UO_2057 (O_2057,N_19300,N_18865);
nor UO_2058 (O_2058,N_19074,N_19161);
and UO_2059 (O_2059,N_18815,N_19308);
and UO_2060 (O_2060,N_18354,N_18552);
and UO_2061 (O_2061,N_18822,N_18515);
nor UO_2062 (O_2062,N_19607,N_18455);
and UO_2063 (O_2063,N_18745,N_18999);
and UO_2064 (O_2064,N_19311,N_18371);
xor UO_2065 (O_2065,N_19514,N_19944);
nor UO_2066 (O_2066,N_19414,N_18397);
nand UO_2067 (O_2067,N_18462,N_18429);
or UO_2068 (O_2068,N_18646,N_18257);
or UO_2069 (O_2069,N_19950,N_18064);
nor UO_2070 (O_2070,N_19547,N_19522);
and UO_2071 (O_2071,N_19783,N_19350);
nor UO_2072 (O_2072,N_19002,N_18923);
or UO_2073 (O_2073,N_18015,N_19081);
and UO_2074 (O_2074,N_19351,N_19096);
nor UO_2075 (O_2075,N_18868,N_18324);
or UO_2076 (O_2076,N_18812,N_19398);
or UO_2077 (O_2077,N_18964,N_19081);
nand UO_2078 (O_2078,N_19563,N_18170);
and UO_2079 (O_2079,N_19111,N_19913);
and UO_2080 (O_2080,N_18326,N_18884);
or UO_2081 (O_2081,N_19320,N_19747);
nor UO_2082 (O_2082,N_19462,N_19810);
nand UO_2083 (O_2083,N_18850,N_18055);
or UO_2084 (O_2084,N_18973,N_19210);
nor UO_2085 (O_2085,N_19057,N_18875);
and UO_2086 (O_2086,N_18208,N_18767);
or UO_2087 (O_2087,N_19317,N_19493);
nor UO_2088 (O_2088,N_19784,N_19247);
or UO_2089 (O_2089,N_19824,N_19882);
xor UO_2090 (O_2090,N_18474,N_18816);
nand UO_2091 (O_2091,N_19290,N_19142);
nand UO_2092 (O_2092,N_19078,N_18530);
xnor UO_2093 (O_2093,N_19948,N_19113);
or UO_2094 (O_2094,N_18291,N_19006);
and UO_2095 (O_2095,N_19050,N_18436);
or UO_2096 (O_2096,N_19813,N_18743);
xnor UO_2097 (O_2097,N_18518,N_19836);
and UO_2098 (O_2098,N_19252,N_19798);
nor UO_2099 (O_2099,N_18819,N_18376);
or UO_2100 (O_2100,N_18595,N_19725);
xor UO_2101 (O_2101,N_18100,N_18294);
nand UO_2102 (O_2102,N_19233,N_18780);
nand UO_2103 (O_2103,N_19574,N_18859);
nand UO_2104 (O_2104,N_19518,N_19123);
nand UO_2105 (O_2105,N_19117,N_18553);
and UO_2106 (O_2106,N_18553,N_18694);
and UO_2107 (O_2107,N_19777,N_18179);
nor UO_2108 (O_2108,N_18347,N_19056);
and UO_2109 (O_2109,N_19642,N_18056);
nor UO_2110 (O_2110,N_18643,N_18031);
nand UO_2111 (O_2111,N_18705,N_19630);
or UO_2112 (O_2112,N_18392,N_18408);
nor UO_2113 (O_2113,N_18121,N_19204);
and UO_2114 (O_2114,N_18176,N_19466);
or UO_2115 (O_2115,N_19332,N_19247);
nor UO_2116 (O_2116,N_18764,N_18424);
nor UO_2117 (O_2117,N_19040,N_19602);
xor UO_2118 (O_2118,N_18149,N_19049);
or UO_2119 (O_2119,N_18086,N_18546);
and UO_2120 (O_2120,N_19944,N_18141);
and UO_2121 (O_2121,N_19741,N_18774);
or UO_2122 (O_2122,N_19606,N_19927);
and UO_2123 (O_2123,N_19947,N_19335);
nand UO_2124 (O_2124,N_18921,N_19050);
and UO_2125 (O_2125,N_19841,N_18197);
nor UO_2126 (O_2126,N_19797,N_18392);
xor UO_2127 (O_2127,N_18118,N_19163);
or UO_2128 (O_2128,N_19050,N_19730);
and UO_2129 (O_2129,N_18364,N_19303);
and UO_2130 (O_2130,N_19737,N_18735);
and UO_2131 (O_2131,N_19312,N_19522);
nand UO_2132 (O_2132,N_18254,N_19009);
nand UO_2133 (O_2133,N_19512,N_18388);
and UO_2134 (O_2134,N_19463,N_18415);
nor UO_2135 (O_2135,N_18397,N_19811);
and UO_2136 (O_2136,N_19870,N_19667);
nor UO_2137 (O_2137,N_19152,N_19663);
nand UO_2138 (O_2138,N_18972,N_18273);
and UO_2139 (O_2139,N_18196,N_19101);
or UO_2140 (O_2140,N_18908,N_18220);
nor UO_2141 (O_2141,N_19820,N_19906);
or UO_2142 (O_2142,N_18867,N_19641);
nor UO_2143 (O_2143,N_19172,N_18080);
nor UO_2144 (O_2144,N_18451,N_19262);
nand UO_2145 (O_2145,N_19042,N_19688);
xor UO_2146 (O_2146,N_18900,N_18847);
nor UO_2147 (O_2147,N_18955,N_19506);
and UO_2148 (O_2148,N_19684,N_18324);
or UO_2149 (O_2149,N_18219,N_18839);
and UO_2150 (O_2150,N_18881,N_18270);
or UO_2151 (O_2151,N_19306,N_19059);
nand UO_2152 (O_2152,N_18259,N_19317);
or UO_2153 (O_2153,N_19343,N_18315);
or UO_2154 (O_2154,N_18674,N_19309);
or UO_2155 (O_2155,N_19045,N_19132);
and UO_2156 (O_2156,N_18929,N_18362);
nand UO_2157 (O_2157,N_18242,N_18812);
nand UO_2158 (O_2158,N_18611,N_18370);
nand UO_2159 (O_2159,N_18863,N_18512);
or UO_2160 (O_2160,N_18009,N_18789);
nor UO_2161 (O_2161,N_18819,N_19173);
or UO_2162 (O_2162,N_18179,N_19554);
or UO_2163 (O_2163,N_19369,N_19815);
and UO_2164 (O_2164,N_19557,N_19765);
nor UO_2165 (O_2165,N_18729,N_18337);
or UO_2166 (O_2166,N_18731,N_19861);
and UO_2167 (O_2167,N_19764,N_19580);
or UO_2168 (O_2168,N_18474,N_19690);
nor UO_2169 (O_2169,N_18596,N_18425);
or UO_2170 (O_2170,N_18495,N_18117);
nor UO_2171 (O_2171,N_18649,N_19623);
nand UO_2172 (O_2172,N_19829,N_18295);
or UO_2173 (O_2173,N_19614,N_19095);
and UO_2174 (O_2174,N_18350,N_18634);
and UO_2175 (O_2175,N_19983,N_19848);
or UO_2176 (O_2176,N_19554,N_19502);
and UO_2177 (O_2177,N_19589,N_18817);
nor UO_2178 (O_2178,N_18024,N_19934);
nand UO_2179 (O_2179,N_19441,N_19764);
xnor UO_2180 (O_2180,N_19161,N_18180);
xor UO_2181 (O_2181,N_19203,N_19042);
nand UO_2182 (O_2182,N_18673,N_19076);
and UO_2183 (O_2183,N_19553,N_18097);
and UO_2184 (O_2184,N_18962,N_19501);
nor UO_2185 (O_2185,N_18539,N_18629);
nand UO_2186 (O_2186,N_19135,N_18670);
nand UO_2187 (O_2187,N_18350,N_18495);
or UO_2188 (O_2188,N_18952,N_19744);
xnor UO_2189 (O_2189,N_18063,N_18689);
and UO_2190 (O_2190,N_19372,N_18142);
nor UO_2191 (O_2191,N_19573,N_18404);
nand UO_2192 (O_2192,N_19885,N_18240);
and UO_2193 (O_2193,N_18472,N_18124);
and UO_2194 (O_2194,N_19148,N_19737);
nand UO_2195 (O_2195,N_18559,N_19002);
nor UO_2196 (O_2196,N_19908,N_19772);
or UO_2197 (O_2197,N_18093,N_19916);
nor UO_2198 (O_2198,N_18312,N_19341);
xor UO_2199 (O_2199,N_19119,N_18498);
nor UO_2200 (O_2200,N_19024,N_19364);
nand UO_2201 (O_2201,N_19448,N_18969);
and UO_2202 (O_2202,N_19272,N_18404);
or UO_2203 (O_2203,N_18046,N_19190);
or UO_2204 (O_2204,N_19844,N_19661);
nor UO_2205 (O_2205,N_18859,N_19021);
or UO_2206 (O_2206,N_18883,N_18100);
or UO_2207 (O_2207,N_18446,N_19665);
nor UO_2208 (O_2208,N_19013,N_18350);
or UO_2209 (O_2209,N_18084,N_18022);
nand UO_2210 (O_2210,N_18906,N_19481);
or UO_2211 (O_2211,N_18697,N_19883);
nand UO_2212 (O_2212,N_19575,N_19089);
nor UO_2213 (O_2213,N_18218,N_19522);
nor UO_2214 (O_2214,N_18986,N_19978);
nor UO_2215 (O_2215,N_18298,N_19665);
or UO_2216 (O_2216,N_18353,N_18905);
nand UO_2217 (O_2217,N_18800,N_19182);
nand UO_2218 (O_2218,N_18164,N_19653);
xnor UO_2219 (O_2219,N_18744,N_19319);
and UO_2220 (O_2220,N_18425,N_19187);
and UO_2221 (O_2221,N_19745,N_18630);
or UO_2222 (O_2222,N_18405,N_18406);
or UO_2223 (O_2223,N_19062,N_19750);
or UO_2224 (O_2224,N_18084,N_19646);
nor UO_2225 (O_2225,N_19313,N_18858);
nor UO_2226 (O_2226,N_19964,N_18672);
xnor UO_2227 (O_2227,N_19102,N_18393);
and UO_2228 (O_2228,N_18721,N_19687);
and UO_2229 (O_2229,N_19958,N_19272);
nand UO_2230 (O_2230,N_18752,N_19819);
nand UO_2231 (O_2231,N_18679,N_18644);
xor UO_2232 (O_2232,N_18671,N_19846);
nor UO_2233 (O_2233,N_19115,N_18790);
nor UO_2234 (O_2234,N_18969,N_19037);
or UO_2235 (O_2235,N_19631,N_18331);
nor UO_2236 (O_2236,N_19625,N_18713);
nand UO_2237 (O_2237,N_19195,N_18397);
xor UO_2238 (O_2238,N_19080,N_18385);
nand UO_2239 (O_2239,N_19075,N_19167);
nand UO_2240 (O_2240,N_18238,N_19691);
nor UO_2241 (O_2241,N_18125,N_18128);
nor UO_2242 (O_2242,N_18332,N_19379);
xor UO_2243 (O_2243,N_19567,N_18940);
nand UO_2244 (O_2244,N_18762,N_18403);
or UO_2245 (O_2245,N_18792,N_18419);
or UO_2246 (O_2246,N_18857,N_19597);
nand UO_2247 (O_2247,N_19503,N_18362);
or UO_2248 (O_2248,N_18535,N_19875);
or UO_2249 (O_2249,N_18145,N_19350);
nand UO_2250 (O_2250,N_18228,N_19614);
xor UO_2251 (O_2251,N_19960,N_19301);
and UO_2252 (O_2252,N_19151,N_18529);
nor UO_2253 (O_2253,N_19555,N_18073);
or UO_2254 (O_2254,N_19774,N_18572);
or UO_2255 (O_2255,N_19674,N_19639);
xor UO_2256 (O_2256,N_19099,N_19638);
xnor UO_2257 (O_2257,N_18793,N_18585);
nand UO_2258 (O_2258,N_18953,N_19814);
nor UO_2259 (O_2259,N_19390,N_19180);
nand UO_2260 (O_2260,N_18507,N_18501);
and UO_2261 (O_2261,N_19622,N_18433);
or UO_2262 (O_2262,N_19081,N_18511);
and UO_2263 (O_2263,N_18844,N_19460);
or UO_2264 (O_2264,N_18877,N_19127);
or UO_2265 (O_2265,N_18907,N_18645);
nor UO_2266 (O_2266,N_18059,N_18467);
nor UO_2267 (O_2267,N_18187,N_18188);
nor UO_2268 (O_2268,N_19217,N_19427);
or UO_2269 (O_2269,N_18625,N_19185);
or UO_2270 (O_2270,N_19627,N_18045);
nand UO_2271 (O_2271,N_19102,N_19897);
or UO_2272 (O_2272,N_18645,N_18592);
and UO_2273 (O_2273,N_19439,N_18280);
or UO_2274 (O_2274,N_19106,N_18972);
xor UO_2275 (O_2275,N_19717,N_18899);
or UO_2276 (O_2276,N_19678,N_19563);
or UO_2277 (O_2277,N_18145,N_18100);
nor UO_2278 (O_2278,N_19837,N_18374);
xor UO_2279 (O_2279,N_18743,N_19024);
nand UO_2280 (O_2280,N_18644,N_18394);
nand UO_2281 (O_2281,N_18161,N_18459);
nand UO_2282 (O_2282,N_19994,N_18874);
nand UO_2283 (O_2283,N_18370,N_19284);
nand UO_2284 (O_2284,N_18584,N_19241);
and UO_2285 (O_2285,N_19958,N_18794);
or UO_2286 (O_2286,N_19766,N_19010);
and UO_2287 (O_2287,N_19705,N_19560);
nor UO_2288 (O_2288,N_18142,N_18242);
nand UO_2289 (O_2289,N_18398,N_19860);
or UO_2290 (O_2290,N_18154,N_19881);
nor UO_2291 (O_2291,N_18759,N_18987);
and UO_2292 (O_2292,N_19595,N_19010);
and UO_2293 (O_2293,N_19168,N_18677);
xnor UO_2294 (O_2294,N_18968,N_19238);
or UO_2295 (O_2295,N_18659,N_18129);
nand UO_2296 (O_2296,N_18436,N_18991);
and UO_2297 (O_2297,N_18326,N_18375);
and UO_2298 (O_2298,N_19041,N_18243);
nand UO_2299 (O_2299,N_18284,N_19806);
nor UO_2300 (O_2300,N_18097,N_18374);
or UO_2301 (O_2301,N_19864,N_19781);
nand UO_2302 (O_2302,N_19009,N_19963);
nand UO_2303 (O_2303,N_19321,N_19761);
or UO_2304 (O_2304,N_19814,N_19641);
or UO_2305 (O_2305,N_18882,N_19683);
and UO_2306 (O_2306,N_19571,N_18598);
nor UO_2307 (O_2307,N_18810,N_19864);
xnor UO_2308 (O_2308,N_19959,N_19981);
and UO_2309 (O_2309,N_18738,N_19125);
nand UO_2310 (O_2310,N_19132,N_18053);
nand UO_2311 (O_2311,N_18123,N_18332);
xor UO_2312 (O_2312,N_18528,N_19016);
nand UO_2313 (O_2313,N_18077,N_18737);
nand UO_2314 (O_2314,N_18898,N_19906);
or UO_2315 (O_2315,N_19859,N_19314);
and UO_2316 (O_2316,N_19340,N_18736);
or UO_2317 (O_2317,N_18489,N_18572);
nor UO_2318 (O_2318,N_19726,N_18907);
nor UO_2319 (O_2319,N_18986,N_18799);
xnor UO_2320 (O_2320,N_18497,N_18872);
and UO_2321 (O_2321,N_19779,N_19030);
nand UO_2322 (O_2322,N_19500,N_19315);
nor UO_2323 (O_2323,N_19929,N_18763);
and UO_2324 (O_2324,N_19572,N_19210);
nor UO_2325 (O_2325,N_18377,N_18950);
nand UO_2326 (O_2326,N_19097,N_19347);
or UO_2327 (O_2327,N_18059,N_18304);
nand UO_2328 (O_2328,N_18674,N_19426);
and UO_2329 (O_2329,N_18723,N_18019);
and UO_2330 (O_2330,N_19373,N_18009);
xnor UO_2331 (O_2331,N_18080,N_19901);
nand UO_2332 (O_2332,N_18525,N_18686);
nor UO_2333 (O_2333,N_18927,N_19577);
nand UO_2334 (O_2334,N_18451,N_18974);
or UO_2335 (O_2335,N_19561,N_19507);
nand UO_2336 (O_2336,N_19567,N_19660);
or UO_2337 (O_2337,N_18792,N_19062);
and UO_2338 (O_2338,N_18089,N_18221);
and UO_2339 (O_2339,N_18399,N_19706);
nand UO_2340 (O_2340,N_19122,N_19406);
and UO_2341 (O_2341,N_19160,N_18658);
or UO_2342 (O_2342,N_18138,N_18045);
and UO_2343 (O_2343,N_18351,N_19853);
nand UO_2344 (O_2344,N_19298,N_19833);
nor UO_2345 (O_2345,N_19486,N_18804);
nand UO_2346 (O_2346,N_19634,N_19179);
nand UO_2347 (O_2347,N_18094,N_18381);
or UO_2348 (O_2348,N_18890,N_18341);
nor UO_2349 (O_2349,N_18328,N_19733);
and UO_2350 (O_2350,N_19257,N_19553);
and UO_2351 (O_2351,N_18875,N_18893);
nor UO_2352 (O_2352,N_18664,N_18071);
and UO_2353 (O_2353,N_18654,N_19420);
and UO_2354 (O_2354,N_18164,N_18295);
or UO_2355 (O_2355,N_19490,N_18607);
or UO_2356 (O_2356,N_18695,N_19636);
nand UO_2357 (O_2357,N_19381,N_19071);
or UO_2358 (O_2358,N_18461,N_19166);
nand UO_2359 (O_2359,N_19651,N_18655);
nor UO_2360 (O_2360,N_18328,N_18581);
or UO_2361 (O_2361,N_18537,N_18376);
nand UO_2362 (O_2362,N_19400,N_19702);
xnor UO_2363 (O_2363,N_18841,N_18956);
and UO_2364 (O_2364,N_19275,N_18882);
or UO_2365 (O_2365,N_19323,N_18366);
or UO_2366 (O_2366,N_19000,N_18587);
nand UO_2367 (O_2367,N_18966,N_19525);
xor UO_2368 (O_2368,N_19874,N_18143);
nor UO_2369 (O_2369,N_18938,N_19392);
or UO_2370 (O_2370,N_19804,N_18011);
or UO_2371 (O_2371,N_19187,N_19263);
or UO_2372 (O_2372,N_18298,N_18365);
nand UO_2373 (O_2373,N_18886,N_18787);
nand UO_2374 (O_2374,N_18202,N_19677);
or UO_2375 (O_2375,N_19607,N_18549);
nand UO_2376 (O_2376,N_19974,N_19089);
or UO_2377 (O_2377,N_19211,N_18733);
and UO_2378 (O_2378,N_19888,N_19158);
and UO_2379 (O_2379,N_19642,N_19713);
nand UO_2380 (O_2380,N_18003,N_19780);
nor UO_2381 (O_2381,N_19234,N_18094);
nor UO_2382 (O_2382,N_19561,N_19048);
nand UO_2383 (O_2383,N_18184,N_18483);
xor UO_2384 (O_2384,N_19809,N_18661);
and UO_2385 (O_2385,N_19376,N_19507);
and UO_2386 (O_2386,N_18113,N_19286);
nand UO_2387 (O_2387,N_18816,N_18306);
and UO_2388 (O_2388,N_19963,N_18004);
nor UO_2389 (O_2389,N_19605,N_19190);
and UO_2390 (O_2390,N_18265,N_19582);
nor UO_2391 (O_2391,N_18167,N_18280);
nand UO_2392 (O_2392,N_19271,N_18670);
nand UO_2393 (O_2393,N_18747,N_19220);
nor UO_2394 (O_2394,N_18865,N_18627);
nor UO_2395 (O_2395,N_19544,N_19911);
or UO_2396 (O_2396,N_19042,N_19015);
nand UO_2397 (O_2397,N_19782,N_18674);
or UO_2398 (O_2398,N_18689,N_18488);
nand UO_2399 (O_2399,N_19400,N_18543);
nand UO_2400 (O_2400,N_18100,N_18415);
or UO_2401 (O_2401,N_18074,N_19235);
nand UO_2402 (O_2402,N_18368,N_18250);
nand UO_2403 (O_2403,N_18786,N_19487);
nor UO_2404 (O_2404,N_18025,N_19520);
and UO_2405 (O_2405,N_18767,N_18976);
and UO_2406 (O_2406,N_19671,N_18642);
and UO_2407 (O_2407,N_18257,N_18909);
or UO_2408 (O_2408,N_19281,N_18054);
or UO_2409 (O_2409,N_18771,N_18463);
or UO_2410 (O_2410,N_18739,N_19809);
and UO_2411 (O_2411,N_19140,N_19241);
nand UO_2412 (O_2412,N_18380,N_19152);
nor UO_2413 (O_2413,N_19590,N_18106);
and UO_2414 (O_2414,N_19113,N_18277);
nand UO_2415 (O_2415,N_18435,N_18744);
nand UO_2416 (O_2416,N_18268,N_18189);
nand UO_2417 (O_2417,N_18953,N_18520);
nor UO_2418 (O_2418,N_19850,N_18880);
or UO_2419 (O_2419,N_19888,N_18437);
or UO_2420 (O_2420,N_18924,N_18762);
nor UO_2421 (O_2421,N_19537,N_19087);
and UO_2422 (O_2422,N_18461,N_19291);
or UO_2423 (O_2423,N_18819,N_19384);
nand UO_2424 (O_2424,N_18562,N_19398);
nand UO_2425 (O_2425,N_18681,N_18182);
nand UO_2426 (O_2426,N_19885,N_19976);
or UO_2427 (O_2427,N_19199,N_18946);
or UO_2428 (O_2428,N_19223,N_18591);
nor UO_2429 (O_2429,N_18591,N_18230);
or UO_2430 (O_2430,N_18581,N_19797);
xor UO_2431 (O_2431,N_19897,N_19217);
nor UO_2432 (O_2432,N_18389,N_18037);
nor UO_2433 (O_2433,N_18517,N_18288);
or UO_2434 (O_2434,N_19864,N_19568);
and UO_2435 (O_2435,N_19146,N_19743);
nand UO_2436 (O_2436,N_18799,N_18098);
or UO_2437 (O_2437,N_19462,N_19319);
xnor UO_2438 (O_2438,N_19932,N_18928);
nand UO_2439 (O_2439,N_18433,N_19944);
and UO_2440 (O_2440,N_19256,N_18113);
and UO_2441 (O_2441,N_18152,N_19876);
nor UO_2442 (O_2442,N_19082,N_19309);
nand UO_2443 (O_2443,N_19397,N_19868);
nand UO_2444 (O_2444,N_19681,N_19932);
and UO_2445 (O_2445,N_18590,N_19746);
nand UO_2446 (O_2446,N_19196,N_18341);
xor UO_2447 (O_2447,N_18524,N_19910);
and UO_2448 (O_2448,N_19474,N_18903);
nand UO_2449 (O_2449,N_18111,N_19472);
nand UO_2450 (O_2450,N_19037,N_19738);
nand UO_2451 (O_2451,N_18033,N_18968);
nand UO_2452 (O_2452,N_18839,N_19534);
or UO_2453 (O_2453,N_19274,N_19098);
nand UO_2454 (O_2454,N_19624,N_18104);
or UO_2455 (O_2455,N_18042,N_19353);
nand UO_2456 (O_2456,N_19962,N_19191);
xnor UO_2457 (O_2457,N_18948,N_18555);
or UO_2458 (O_2458,N_18374,N_18726);
xnor UO_2459 (O_2459,N_18020,N_18037);
or UO_2460 (O_2460,N_19842,N_19930);
nor UO_2461 (O_2461,N_19949,N_19699);
or UO_2462 (O_2462,N_19877,N_18773);
nor UO_2463 (O_2463,N_18390,N_19045);
nand UO_2464 (O_2464,N_19988,N_18058);
nor UO_2465 (O_2465,N_18269,N_18969);
or UO_2466 (O_2466,N_18826,N_19794);
nor UO_2467 (O_2467,N_19180,N_19864);
and UO_2468 (O_2468,N_19335,N_18130);
nor UO_2469 (O_2469,N_18707,N_19244);
and UO_2470 (O_2470,N_19876,N_19921);
nor UO_2471 (O_2471,N_18220,N_19263);
xnor UO_2472 (O_2472,N_19801,N_19750);
nor UO_2473 (O_2473,N_18421,N_19174);
and UO_2474 (O_2474,N_18820,N_19144);
xor UO_2475 (O_2475,N_18517,N_18632);
xor UO_2476 (O_2476,N_19161,N_19007);
or UO_2477 (O_2477,N_18670,N_18442);
nor UO_2478 (O_2478,N_19347,N_18705);
xor UO_2479 (O_2479,N_19574,N_18782);
and UO_2480 (O_2480,N_18324,N_19918);
and UO_2481 (O_2481,N_19870,N_18753);
nand UO_2482 (O_2482,N_18622,N_18224);
nand UO_2483 (O_2483,N_18366,N_18330);
nand UO_2484 (O_2484,N_19469,N_18676);
xor UO_2485 (O_2485,N_18877,N_19909);
and UO_2486 (O_2486,N_18530,N_18762);
nand UO_2487 (O_2487,N_19266,N_18825);
or UO_2488 (O_2488,N_19428,N_18410);
nor UO_2489 (O_2489,N_18920,N_19563);
and UO_2490 (O_2490,N_19714,N_19666);
and UO_2491 (O_2491,N_18227,N_18852);
nand UO_2492 (O_2492,N_18301,N_19251);
or UO_2493 (O_2493,N_18884,N_18925);
nor UO_2494 (O_2494,N_19578,N_18322);
or UO_2495 (O_2495,N_18551,N_19664);
or UO_2496 (O_2496,N_18791,N_18007);
nor UO_2497 (O_2497,N_19995,N_19184);
and UO_2498 (O_2498,N_19129,N_18579);
or UO_2499 (O_2499,N_19955,N_19038);
endmodule