module basic_1500_15000_2000_10_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xor U0 (N_0,In_1441,In_479);
and U1 (N_1,In_968,In_42);
and U2 (N_2,In_736,In_466);
and U3 (N_3,In_553,In_1263);
nor U4 (N_4,In_876,In_778);
xor U5 (N_5,In_510,In_561);
nor U6 (N_6,In_344,In_1354);
xor U7 (N_7,In_258,In_725);
or U8 (N_8,In_250,In_1119);
xor U9 (N_9,In_224,In_418);
xor U10 (N_10,In_757,In_1126);
xnor U11 (N_11,In_305,In_822);
xnor U12 (N_12,In_808,In_57);
xnor U13 (N_13,In_162,In_1059);
xnor U14 (N_14,In_97,In_313);
xor U15 (N_15,In_319,In_1295);
xor U16 (N_16,In_217,In_1363);
nand U17 (N_17,In_973,In_159);
nor U18 (N_18,In_1129,In_491);
and U19 (N_19,In_1134,In_1194);
or U20 (N_20,In_113,In_790);
nand U21 (N_21,In_55,In_147);
or U22 (N_22,In_1311,In_14);
nand U23 (N_23,In_403,In_35);
and U24 (N_24,In_1147,In_1451);
nand U25 (N_25,In_744,In_525);
xor U26 (N_26,In_285,In_15);
xor U27 (N_27,In_229,In_680);
and U28 (N_28,In_1381,In_1056);
nand U29 (N_29,In_289,In_396);
or U30 (N_30,In_27,In_407);
and U31 (N_31,In_1327,In_509);
and U32 (N_32,In_1031,In_464);
xnor U33 (N_33,In_1471,In_656);
nand U34 (N_34,In_648,In_26);
and U35 (N_35,In_1048,In_2);
or U36 (N_36,In_671,In_1369);
and U37 (N_37,In_228,In_722);
nand U38 (N_38,In_379,In_1483);
or U39 (N_39,In_1087,In_1411);
nor U40 (N_40,In_1230,In_904);
nand U41 (N_41,In_153,In_307);
and U42 (N_42,In_293,In_1051);
xor U43 (N_43,In_607,In_552);
xnor U44 (N_44,In_1320,In_686);
nand U45 (N_45,In_538,In_1495);
nand U46 (N_46,In_169,In_706);
xnor U47 (N_47,In_1359,In_1341);
nand U48 (N_48,In_1337,In_184);
and U49 (N_49,In_1437,In_43);
nand U50 (N_50,In_928,In_1460);
nand U51 (N_51,In_991,In_1185);
and U52 (N_52,In_1271,In_683);
nand U53 (N_53,In_892,In_354);
or U54 (N_54,In_1035,In_554);
xnor U55 (N_55,In_106,In_65);
xnor U56 (N_56,In_1082,In_131);
nor U57 (N_57,In_267,In_1218);
and U58 (N_58,In_916,In_74);
and U59 (N_59,In_103,In_748);
nor U60 (N_60,In_277,In_30);
nor U61 (N_61,In_494,In_961);
xor U62 (N_62,In_801,In_815);
nand U63 (N_63,In_109,In_1440);
or U64 (N_64,In_426,In_85);
nor U65 (N_65,In_337,In_1006);
and U66 (N_66,In_1278,In_545);
nand U67 (N_67,In_1050,In_579);
nor U68 (N_68,In_523,In_318);
nand U69 (N_69,In_1165,In_397);
or U70 (N_70,In_457,In_36);
nand U71 (N_71,In_168,In_256);
or U72 (N_72,In_597,In_328);
nand U73 (N_73,In_259,In_828);
nor U74 (N_74,In_998,In_1153);
xor U75 (N_75,In_1308,In_1306);
nor U76 (N_76,In_942,In_1488);
nand U77 (N_77,In_239,In_1497);
nand U78 (N_78,In_681,In_729);
and U79 (N_79,In_284,In_1044);
and U80 (N_80,In_534,In_436);
and U81 (N_81,In_831,In_88);
or U82 (N_82,In_992,In_754);
nand U83 (N_83,In_115,In_616);
nor U84 (N_84,In_170,In_1128);
nor U85 (N_85,In_528,In_1052);
xor U86 (N_86,In_689,In_410);
and U87 (N_87,In_101,In_614);
or U88 (N_88,In_927,In_516);
nor U89 (N_89,In_1221,In_1178);
nand U90 (N_90,In_1074,In_402);
or U91 (N_91,In_272,In_895);
or U92 (N_92,In_1344,In_690);
nor U93 (N_93,In_618,In_434);
nor U94 (N_94,In_529,In_1003);
nor U95 (N_95,In_1092,In_260);
nand U96 (N_96,In_1105,In_1156);
xor U97 (N_97,In_1253,In_165);
nand U98 (N_98,In_726,In_513);
and U99 (N_99,In_1388,In_1386);
nand U100 (N_100,In_732,In_1070);
nor U101 (N_101,In_79,In_160);
xor U102 (N_102,In_66,In_329);
xor U103 (N_103,In_1420,In_1109);
nor U104 (N_104,In_1468,In_455);
xnor U105 (N_105,In_915,In_1205);
nor U106 (N_106,In_874,In_932);
nor U107 (N_107,In_734,In_214);
or U108 (N_108,In_629,In_1414);
or U109 (N_109,In_1115,In_363);
nor U110 (N_110,In_1290,In_1045);
or U111 (N_111,In_143,In_136);
nor U112 (N_112,In_201,In_745);
or U113 (N_113,In_501,In_1355);
or U114 (N_114,In_1004,In_727);
or U115 (N_115,In_39,In_785);
xnor U116 (N_116,In_708,In_1453);
or U117 (N_117,In_70,In_743);
nor U118 (N_118,In_41,In_1088);
nor U119 (N_119,In_1304,In_419);
and U120 (N_120,In_565,In_636);
and U121 (N_121,In_1060,In_580);
nor U122 (N_122,In_204,In_1328);
nand U123 (N_123,In_1356,In_202);
xor U124 (N_124,In_530,In_522);
nor U125 (N_125,In_247,In_1100);
or U126 (N_126,In_886,In_560);
or U127 (N_127,In_1462,In_1346);
nor U128 (N_128,In_1323,In_659);
nand U129 (N_129,In_124,In_837);
or U130 (N_130,In_302,In_769);
nor U131 (N_131,In_638,In_943);
or U132 (N_132,In_612,In_28);
nand U133 (N_133,In_430,In_1436);
nor U134 (N_134,In_888,In_639);
and U135 (N_135,In_46,In_1001);
nand U136 (N_136,In_1431,In_414);
nor U137 (N_137,In_644,In_650);
and U138 (N_138,In_226,In_863);
and U139 (N_139,In_427,In_1423);
and U140 (N_140,In_613,In_849);
or U141 (N_141,In_898,In_38);
or U142 (N_142,In_1293,In_1492);
xnor U143 (N_143,In_733,In_1174);
or U144 (N_144,In_1039,In_399);
or U145 (N_145,In_753,In_723);
nor U146 (N_146,In_702,In_796);
nand U147 (N_147,In_811,In_810);
and U148 (N_148,In_1254,In_1379);
or U149 (N_149,In_975,In_1152);
and U150 (N_150,In_905,In_541);
or U151 (N_151,In_454,In_804);
nand U152 (N_152,In_1400,In_1457);
and U153 (N_153,In_1118,In_87);
xor U154 (N_154,In_884,In_310);
and U155 (N_155,In_728,In_645);
and U156 (N_156,In_295,In_634);
nor U157 (N_157,In_1485,In_472);
xor U158 (N_158,In_1244,In_1260);
nor U159 (N_159,In_1315,In_1104);
nand U160 (N_160,In_969,In_248);
xnor U161 (N_161,In_1120,In_635);
and U162 (N_162,In_1268,In_1009);
or U163 (N_163,In_1287,In_550);
and U164 (N_164,In_1324,In_548);
xor U165 (N_165,In_666,In_742);
nor U166 (N_166,In_1089,In_766);
and U167 (N_167,In_1191,In_405);
and U168 (N_168,In_1421,In_518);
nand U169 (N_169,In_1302,In_1404);
nor U170 (N_170,In_460,In_1209);
nand U171 (N_171,In_1061,In_16);
xnor U172 (N_172,In_314,In_192);
or U173 (N_173,In_1223,In_951);
nand U174 (N_174,In_620,In_1279);
nand U175 (N_175,In_846,In_383);
xnor U176 (N_176,In_21,In_1188);
nor U177 (N_177,In_227,In_1464);
xor U178 (N_178,In_1055,In_572);
nand U179 (N_179,In_151,In_566);
or U180 (N_180,In_6,In_133);
nand U181 (N_181,In_242,In_33);
nand U182 (N_182,In_965,In_1390);
nor U183 (N_183,In_61,In_1330);
and U184 (N_184,In_956,In_206);
and U185 (N_185,In_440,In_263);
xnor U186 (N_186,In_1124,In_406);
nand U187 (N_187,In_118,In_1175);
xor U188 (N_188,In_506,In_531);
nor U189 (N_189,In_1406,In_347);
and U190 (N_190,In_569,In_409);
and U191 (N_191,In_326,In_1317);
nand U192 (N_192,In_1452,In_489);
and U193 (N_193,In_428,In_76);
nand U194 (N_194,In_979,In_1450);
or U195 (N_195,In_843,In_237);
xor U196 (N_196,In_899,In_970);
or U197 (N_197,In_717,In_292);
nor U198 (N_198,In_558,In_497);
xnor U199 (N_199,In_477,In_154);
nor U200 (N_200,In_338,In_661);
xor U201 (N_201,In_448,In_611);
xnor U202 (N_202,In_922,In_1480);
and U203 (N_203,In_606,In_1106);
and U204 (N_204,In_1395,In_1215);
or U205 (N_205,In_1357,In_1176);
or U206 (N_206,In_929,In_17);
or U207 (N_207,In_487,In_142);
xnor U208 (N_208,In_335,In_731);
and U209 (N_209,In_871,In_852);
nand U210 (N_210,In_1241,In_198);
and U211 (N_211,In_1058,In_8);
or U212 (N_212,In_1099,In_191);
nand U213 (N_213,In_1075,In_841);
xnor U214 (N_214,In_1213,In_148);
nor U215 (N_215,In_210,In_171);
nor U216 (N_216,In_178,In_1387);
nor U217 (N_217,In_301,In_1342);
xor U218 (N_218,In_809,In_350);
and U219 (N_219,In_47,In_213);
nor U220 (N_220,In_1367,In_1490);
and U221 (N_221,In_93,In_1292);
nand U222 (N_222,In_1493,In_741);
nor U223 (N_223,In_903,In_37);
xnor U224 (N_224,In_786,In_799);
or U225 (N_225,In_450,In_940);
xnor U226 (N_226,In_834,In_1322);
xor U227 (N_227,In_926,In_972);
or U228 (N_228,In_1073,In_909);
and U229 (N_229,In_880,In_675);
xor U230 (N_230,In_490,In_707);
or U231 (N_231,In_887,In_1439);
and U232 (N_232,In_127,In_271);
nand U233 (N_233,In_574,In_900);
or U234 (N_234,In_23,In_977);
nor U235 (N_235,In_1442,In_135);
xor U236 (N_236,In_1430,In_1011);
and U237 (N_237,In_166,In_80);
xnor U238 (N_238,In_95,In_715);
nor U239 (N_239,In_670,In_334);
nand U240 (N_240,In_444,In_1362);
or U241 (N_241,In_879,In_392);
nand U242 (N_242,In_243,In_1038);
nor U243 (N_243,In_1478,In_1285);
nand U244 (N_244,In_617,In_411);
or U245 (N_245,In_819,In_327);
or U246 (N_246,In_546,In_642);
or U247 (N_247,In_625,In_788);
xnor U248 (N_248,In_539,In_1247);
xor U249 (N_249,In_286,In_628);
nor U250 (N_250,In_1489,In_1094);
nand U251 (N_251,In_760,In_98);
nand U252 (N_252,In_762,In_1310);
nor U253 (N_253,In_573,In_1000);
and U254 (N_254,In_687,In_1085);
nor U255 (N_255,In_798,In_936);
or U256 (N_256,In_300,In_508);
and U257 (N_257,In_980,In_1427);
nor U258 (N_258,In_592,In_861);
or U259 (N_259,In_483,In_1228);
nand U260 (N_260,In_278,In_370);
nor U261 (N_261,In_1277,In_255);
xnor U262 (N_262,In_1412,In_981);
and U263 (N_263,In_603,In_963);
xnor U264 (N_264,In_694,In_114);
nand U265 (N_265,In_835,In_1158);
nor U266 (N_266,In_864,In_69);
and U267 (N_267,In_1198,In_367);
nand U268 (N_268,In_1361,In_1186);
nor U269 (N_269,In_505,In_262);
nand U270 (N_270,In_205,In_1443);
xnor U271 (N_271,In_782,In_682);
xor U272 (N_272,In_657,In_1032);
or U273 (N_273,In_104,In_691);
nand U274 (N_274,In_346,In_1149);
xor U275 (N_275,In_125,In_390);
or U276 (N_276,In_1280,In_873);
or U277 (N_277,In_352,In_461);
nor U278 (N_278,In_976,In_1382);
nor U279 (N_279,In_578,In_287);
and U280 (N_280,In_1066,In_913);
nor U281 (N_281,In_955,In_492);
nor U282 (N_282,In_947,In_498);
nand U283 (N_283,In_854,In_821);
nand U284 (N_284,In_1020,In_817);
nor U285 (N_285,In_152,In_1234);
and U286 (N_286,In_149,In_375);
nor U287 (N_287,In_1047,In_1413);
nand U288 (N_288,In_374,In_230);
or U289 (N_289,In_608,In_1353);
or U290 (N_290,In_218,In_221);
xnor U291 (N_291,In_1481,In_596);
and U292 (N_292,In_1352,In_986);
nand U293 (N_293,In_1063,In_1180);
or U294 (N_294,In_333,In_1130);
and U295 (N_295,In_1496,In_540);
or U296 (N_296,In_339,In_31);
nand U297 (N_297,In_331,In_233);
or U298 (N_298,In_1296,In_366);
or U299 (N_299,In_679,In_476);
xor U300 (N_300,In_829,In_63);
and U301 (N_301,In_1482,In_1166);
nand U302 (N_302,In_1014,In_1057);
and U303 (N_303,In_997,In_34);
or U304 (N_304,In_1107,In_772);
and U305 (N_305,In_438,In_290);
nor U306 (N_306,In_532,In_1091);
xor U307 (N_307,In_459,In_602);
nand U308 (N_308,In_896,In_1373);
nand U309 (N_309,In_1238,In_298);
xnor U310 (N_310,In_1135,In_562);
nand U311 (N_311,In_860,In_132);
or U312 (N_312,In_1143,In_1172);
xor U313 (N_313,In_1385,In_978);
xor U314 (N_314,In_1142,In_1262);
nand U315 (N_315,In_632,In_294);
or U316 (N_316,In_939,In_77);
and U317 (N_317,In_660,In_249);
nor U318 (N_318,In_86,In_1434);
and U319 (N_319,In_674,In_1329);
or U320 (N_320,In_704,In_1173);
nand U321 (N_321,In_373,In_1257);
nor U322 (N_322,In_600,In_1265);
and U323 (N_323,In_412,In_215);
or U324 (N_324,In_996,In_1312);
nand U325 (N_325,In_989,In_1371);
and U326 (N_326,In_515,In_297);
xnor U327 (N_327,In_853,In_779);
and U328 (N_328,In_130,In_1182);
xor U329 (N_329,In_999,In_699);
or U330 (N_330,In_1083,In_1463);
or U331 (N_331,In_1002,In_839);
and U332 (N_332,In_1125,In_914);
nand U333 (N_333,In_212,In_502);
or U334 (N_334,In_1160,In_433);
nor U335 (N_335,In_1336,In_718);
xor U336 (N_336,In_91,In_110);
nand U337 (N_337,In_842,In_594);
and U338 (N_338,In_850,In_1389);
or U339 (N_339,In_1484,In_244);
or U340 (N_340,In_1169,In_164);
and U341 (N_341,In_1475,In_514);
xnor U342 (N_342,In_567,In_838);
nand U343 (N_343,In_868,In_1110);
nor U344 (N_344,In_468,In_1243);
xnor U345 (N_345,In_179,In_1005);
xor U346 (N_346,In_1077,In_685);
nand U347 (N_347,In_107,In_1095);
nand U348 (N_348,In_1467,In_1409);
xor U349 (N_349,In_643,In_441);
or U350 (N_350,In_667,In_1283);
xnor U351 (N_351,In_398,In_931);
xor U352 (N_352,In_568,In_1137);
nand U353 (N_353,In_68,In_1319);
nand U354 (N_354,In_584,In_950);
nor U355 (N_355,In_480,In_341);
nor U356 (N_356,In_739,In_197);
nand U357 (N_357,In_537,In_13);
or U358 (N_358,In_1347,In_245);
nand U359 (N_359,In_496,In_751);
nor U360 (N_360,In_797,In_1183);
nor U361 (N_361,In_885,In_1065);
nor U362 (N_362,In_234,In_121);
xor U363 (N_363,In_40,In_747);
xnor U364 (N_364,In_776,In_145);
and U365 (N_365,In_527,In_581);
and U366 (N_366,In_544,In_408);
and U367 (N_367,In_1240,In_1398);
nor U368 (N_368,In_1393,In_1249);
xnor U369 (N_369,In_1017,In_1372);
nor U370 (N_370,In_1334,In_937);
xnor U371 (N_371,In_281,In_919);
nand U372 (N_372,In_1473,In_1010);
xnor U373 (N_373,In_1447,In_1401);
and U374 (N_374,In_343,In_1054);
nor U375 (N_375,In_655,In_117);
or U376 (N_376,In_238,In_588);
or U377 (N_377,In_813,In_44);
and U378 (N_378,In_173,In_833);
nand U379 (N_379,In_1008,In_425);
nor U380 (N_380,In_1376,In_369);
xnor U381 (N_381,In_355,In_610);
and U382 (N_382,In_1171,In_53);
nor U383 (N_383,In_869,In_1079);
nand U384 (N_384,In_958,In_1053);
nor U385 (N_385,In_296,In_1019);
and U386 (N_386,In_62,In_1);
and U387 (N_387,In_400,In_1219);
or U388 (N_388,In_669,In_823);
xnor U389 (N_389,In_1380,In_1102);
xor U390 (N_390,In_500,In_672);
and U391 (N_391,In_735,In_1466);
and U392 (N_392,In_1159,In_812);
or U393 (N_393,In_1121,In_1141);
nor U394 (N_394,In_911,In_349);
and U395 (N_395,In_1284,In_1225);
and U396 (N_396,In_32,In_158);
xor U397 (N_397,In_356,In_912);
or U398 (N_398,In_604,In_1399);
nor U399 (N_399,In_647,In_771);
nand U400 (N_400,In_83,In_570);
nor U401 (N_401,In_759,In_1132);
or U402 (N_402,In_1227,In_859);
or U403 (N_403,In_814,In_282);
nor U404 (N_404,In_1392,In_1418);
nand U405 (N_405,In_382,In_67);
and U406 (N_406,In_542,In_551);
nor U407 (N_407,In_587,In_1378);
xor U408 (N_408,In_126,In_595);
xnor U409 (N_409,In_624,In_807);
nand U410 (N_410,In_324,In_816);
or U411 (N_411,In_631,In_1199);
or U412 (N_412,In_740,In_189);
xnor U413 (N_413,In_359,In_60);
nor U414 (N_414,In_697,In_340);
xor U415 (N_415,In_139,In_1368);
nand U416 (N_416,In_493,In_1360);
or U417 (N_417,In_1122,In_1021);
and U418 (N_418,In_1248,In_1235);
xnor U419 (N_419,In_45,In_10);
and U420 (N_420,In_721,In_654);
nor U421 (N_421,In_1184,In_1123);
or U422 (N_422,In_897,In_512);
and U423 (N_423,In_1177,In_49);
and U424 (N_424,In_623,In_1154);
xnor U425 (N_425,In_3,In_621);
xor U426 (N_426,In_29,In_288);
xnor U427 (N_427,In_1348,In_474);
or U428 (N_428,In_478,In_1081);
and U429 (N_429,In_1067,In_724);
xnor U430 (N_430,In_330,In_315);
nand U431 (N_431,In_161,In_615);
and U432 (N_432,In_371,In_985);
nor U433 (N_433,In_1449,In_1375);
nand U434 (N_434,In_1338,In_713);
or U435 (N_435,In_445,In_269);
or U436 (N_436,In_609,In_1432);
nand U437 (N_437,In_555,In_1456);
nand U438 (N_438,In_1316,In_1458);
and U439 (N_439,In_653,In_176);
nor U440 (N_440,In_1161,In_712);
xnor U441 (N_441,In_1397,In_378);
nand U442 (N_442,In_1407,In_750);
or U443 (N_443,In_488,In_458);
nor U444 (N_444,In_100,In_856);
nor U445 (N_445,In_589,In_818);
and U446 (N_446,In_1041,In_71);
and U447 (N_447,In_535,In_141);
xor U448 (N_448,In_138,In_1197);
xor U449 (N_449,In_511,In_1196);
and U450 (N_450,In_872,In_695);
nor U451 (N_451,In_203,In_593);
nand U452 (N_452,In_116,In_705);
xor U453 (N_453,In_484,In_181);
or U454 (N_454,In_280,In_1018);
nand U455 (N_455,In_902,In_1261);
nand U456 (N_456,In_982,In_571);
or U457 (N_457,In_676,In_1448);
nand U458 (N_458,In_1417,In_443);
or U459 (N_459,In_768,In_190);
xor U460 (N_460,In_380,In_1428);
nor U461 (N_461,In_391,In_194);
xor U462 (N_462,In_974,In_1402);
nand U463 (N_463,In_948,In_336);
or U464 (N_464,In_200,In_451);
or U465 (N_465,In_720,In_921);
nand U466 (N_466,In_361,In_820);
nor U467 (N_467,In_1189,In_765);
or U468 (N_468,In_485,In_219);
nand U469 (N_469,In_995,In_223);
xnor U470 (N_470,In_946,In_784);
nor U471 (N_471,In_851,In_368);
or U472 (N_472,In_236,In_719);
and U473 (N_473,In_81,In_1012);
nand U474 (N_474,In_640,In_627);
nand U475 (N_475,In_917,In_1433);
nand U476 (N_476,In_1470,In_783);
or U477 (N_477,In_990,In_439);
or U478 (N_478,In_1289,In_0);
nand U479 (N_479,In_257,In_306);
or U480 (N_480,In_1220,In_1291);
or U481 (N_481,In_598,In_429);
nand U482 (N_482,In_456,In_780);
nor U483 (N_483,In_549,In_1049);
and U484 (N_484,In_51,In_1131);
nor U485 (N_485,In_700,In_1117);
nand U486 (N_486,In_193,In_1140);
nor U487 (N_487,In_901,In_1345);
or U488 (N_488,In_345,In_1144);
and U489 (N_489,In_471,In_1046);
nor U490 (N_490,In_1216,In_1181);
and U491 (N_491,In_1259,In_605);
nor U492 (N_492,In_1207,In_415);
and U493 (N_493,In_1139,In_1093);
nor U494 (N_494,In_1258,In_1445);
or U495 (N_495,In_216,In_82);
nand U496 (N_496,In_1394,In_585);
and U497 (N_497,In_266,In_789);
or U498 (N_498,In_830,In_163);
nor U499 (N_499,In_649,In_945);
and U500 (N_500,In_321,In_449);
or U501 (N_501,In_906,In_54);
nand U502 (N_502,In_1101,In_422);
xor U503 (N_503,In_826,In_1276);
nand U504 (N_504,In_1080,In_325);
or U505 (N_505,In_1343,In_1016);
xor U506 (N_506,In_92,In_377);
nor U507 (N_507,In_883,In_180);
nor U508 (N_508,In_1351,In_692);
xnor U509 (N_509,In_1266,In_935);
nand U510 (N_510,In_312,In_241);
nand U511 (N_511,In_1237,In_1071);
and U512 (N_512,In_1435,In_174);
nor U513 (N_513,In_1274,In_1446);
or U514 (N_514,In_1340,In_5);
and U515 (N_515,In_1007,In_1233);
xnor U516 (N_516,In_953,In_420);
nand U517 (N_517,In_1226,In_222);
nor U518 (N_518,In_90,In_252);
nor U519 (N_519,In_738,In_316);
nand U520 (N_520,In_1146,In_1281);
nor U521 (N_521,In_1255,In_1426);
nand U522 (N_522,In_78,In_1335);
and U523 (N_523,In_401,In_1444);
and U524 (N_524,In_12,In_167);
and U525 (N_525,In_50,In_774);
and U526 (N_526,In_320,In_964);
and U527 (N_527,In_908,In_543);
and U528 (N_528,In_1486,In_526);
and U529 (N_529,In_1068,In_1429);
xnor U530 (N_530,In_129,In_150);
nor U531 (N_531,In_413,In_1229);
nand U532 (N_532,In_453,In_791);
nor U533 (N_533,In_847,In_1364);
xnor U534 (N_534,In_867,In_431);
or U535 (N_535,In_209,In_1096);
nand U536 (N_536,In_240,In_806);
nand U537 (N_537,In_1150,In_64);
xnor U538 (N_538,In_469,In_519);
nand U539 (N_539,In_387,In_1210);
and U540 (N_540,In_467,In_793);
or U541 (N_541,In_767,In_1112);
nand U542 (N_542,In_1242,In_1069);
nor U543 (N_543,In_231,In_1422);
and U544 (N_544,In_22,In_1455);
nand U545 (N_545,In_1349,In_533);
xnor U546 (N_546,In_1299,In_72);
and U547 (N_547,In_432,In_524);
and U548 (N_548,In_1162,In_678);
xor U549 (N_549,In_1275,In_365);
nor U550 (N_550,In_24,In_824);
xor U551 (N_551,In_1403,In_73);
nor U552 (N_552,In_388,In_304);
xnor U553 (N_553,In_591,In_144);
or U554 (N_554,In_954,In_664);
xnor U555 (N_555,In_1015,In_463);
nor U556 (N_556,In_737,In_1391);
and U557 (N_557,In_111,In_993);
or U558 (N_558,In_1300,In_389);
and U559 (N_559,In_1499,In_99);
or U560 (N_560,In_1190,In_875);
nand U561 (N_561,In_652,In_437);
or U562 (N_562,In_577,In_372);
and U563 (N_563,In_499,In_186);
or U564 (N_564,In_1269,In_1148);
or U565 (N_565,In_187,In_332);
and U566 (N_566,In_1333,In_1113);
or U567 (N_567,In_677,In_1301);
or U568 (N_568,In_770,In_547);
xnor U569 (N_569,In_9,In_1203);
nor U570 (N_570,In_848,In_1084);
and U571 (N_571,In_795,In_1232);
nand U572 (N_572,In_1114,In_1286);
and U573 (N_573,In_1078,In_857);
nor U574 (N_574,In_711,In_393);
or U575 (N_575,In_128,In_1250);
xor U576 (N_576,In_1042,In_1025);
nand U577 (N_577,In_1157,In_421);
xnor U578 (N_578,In_557,In_251);
nor U579 (N_579,In_1036,In_599);
nand U580 (N_580,In_482,In_264);
xnor U581 (N_581,In_781,In_196);
and U582 (N_582,In_1192,In_761);
and U583 (N_583,In_185,In_11);
or U584 (N_584,In_794,In_1425);
and U585 (N_585,In_619,In_276);
xnor U586 (N_586,In_394,In_1024);
nor U587 (N_587,In_923,In_755);
or U588 (N_588,In_424,In_983);
nor U589 (N_589,In_658,In_1168);
nand U590 (N_590,In_920,In_1111);
or U591 (N_591,In_357,In_265);
or U592 (N_592,In_381,In_1410);
xor U593 (N_593,In_517,In_1370);
or U594 (N_594,In_1321,In_960);
xnor U595 (N_595,In_1365,In_1288);
or U596 (N_596,In_89,In_253);
and U597 (N_597,In_311,In_1033);
xor U598 (N_598,In_586,In_894);
nor U599 (N_599,In_386,In_1222);
nor U600 (N_600,In_417,In_626);
xnor U601 (N_601,In_58,In_637);
or U602 (N_602,In_416,In_1136);
or U603 (N_603,In_246,In_48);
xnor U604 (N_604,In_362,In_108);
nand U605 (N_605,In_1208,In_971);
nand U606 (N_606,In_1187,In_75);
nand U607 (N_607,In_775,In_1029);
or U608 (N_608,In_1090,In_470);
or U609 (N_609,In_1023,In_758);
xnor U610 (N_610,In_1491,In_1098);
nor U611 (N_611,In_423,In_447);
nand U612 (N_612,In_714,In_836);
xnor U613 (N_613,In_1252,In_465);
nor U614 (N_614,In_452,In_1043);
xnor U615 (N_615,In_1477,In_1193);
nand U616 (N_616,In_709,In_890);
xor U617 (N_617,In_188,In_1116);
or U618 (N_618,In_696,In_376);
nor U619 (N_619,In_1313,In_122);
and U620 (N_620,In_1366,In_752);
nand U621 (N_621,In_274,In_1331);
xnor U622 (N_622,In_384,In_475);
or U623 (N_623,In_1027,In_25);
nand U624 (N_624,In_556,In_716);
nand U625 (N_625,In_119,In_1256);
nor U626 (N_626,In_764,In_1272);
nor U627 (N_627,In_925,In_582);
nand U628 (N_628,In_763,In_877);
and U629 (N_629,In_805,In_773);
nand U630 (N_630,In_1170,In_1163);
nor U631 (N_631,In_1474,In_1064);
nand U632 (N_632,In_827,In_275);
xor U633 (N_633,In_504,In_182);
nand U634 (N_634,In_1405,In_1195);
and U635 (N_635,In_1479,In_907);
and U636 (N_636,In_1408,In_1459);
nor U637 (N_637,In_1013,In_123);
xnor U638 (N_638,In_435,In_665);
and U639 (N_639,In_1383,In_299);
nand U640 (N_640,In_521,In_1204);
xor U641 (N_641,In_507,In_1332);
nor U642 (N_642,In_1037,In_930);
or U643 (N_643,In_646,In_941);
nand U644 (N_644,In_1384,In_1498);
or U645 (N_645,In_195,In_1318);
xor U646 (N_646,In_924,In_220);
and U647 (N_647,In_563,In_749);
and U648 (N_648,In_495,In_1179);
or U649 (N_649,In_536,In_1155);
nor U650 (N_650,In_303,In_232);
nor U651 (N_651,In_1246,In_322);
and U652 (N_652,In_268,In_688);
nand U653 (N_653,In_1103,In_1026);
and U654 (N_654,In_1305,In_1145);
nor U655 (N_655,In_967,In_1151);
or U656 (N_656,In_1138,In_146);
and U657 (N_657,In_261,In_1350);
and U658 (N_658,In_641,In_486);
or U659 (N_659,In_446,In_112);
and U660 (N_660,In_1231,In_279);
and U661 (N_661,In_1419,In_137);
xor U662 (N_662,In_962,In_1108);
xnor U663 (N_663,In_1469,In_1325);
or U664 (N_664,In_1040,In_693);
or U665 (N_665,In_1022,In_442);
nor U666 (N_666,In_891,In_473);
nor U667 (N_667,In_1396,In_211);
xor U668 (N_668,In_878,In_787);
nand U669 (N_669,In_1465,In_283);
or U670 (N_670,In_1267,In_730);
nor U671 (N_671,In_701,In_800);
and U672 (N_672,In_358,In_1297);
nand U673 (N_673,In_317,In_1294);
nor U674 (N_674,In_777,In_673);
nand U675 (N_675,In_1264,In_96);
xor U676 (N_676,In_910,In_270);
nand U677 (N_677,In_481,In_1358);
or U678 (N_678,In_952,In_175);
and U679 (N_679,In_870,In_1438);
xnor U680 (N_680,In_235,In_862);
or U681 (N_681,In_1212,In_1236);
nor U682 (N_682,In_1377,In_601);
xor U683 (N_683,In_918,In_1298);
xnor U684 (N_684,In_684,In_208);
xnor U685 (N_685,In_1326,In_7);
nor U686 (N_686,In_622,In_1097);
nor U687 (N_687,In_583,In_1494);
or U688 (N_688,In_756,In_18);
and U689 (N_689,In_858,In_710);
and U690 (N_690,In_559,In_94);
nor U691 (N_691,In_351,In_845);
or U692 (N_692,In_1224,In_1167);
nor U693 (N_693,In_564,In_934);
xor U694 (N_694,In_698,In_966);
nand U695 (N_695,In_1416,In_1309);
nor U696 (N_696,In_662,In_364);
and U697 (N_697,In_1303,In_881);
xnor U698 (N_698,In_105,In_172);
or U699 (N_699,In_893,In_1086);
nand U700 (N_700,In_933,In_19);
nand U701 (N_701,In_348,In_291);
nor U702 (N_702,In_1239,In_140);
and U703 (N_703,In_938,In_1217);
xnor U704 (N_704,In_889,In_52);
and U705 (N_705,In_803,In_882);
nand U706 (N_706,In_957,In_802);
xor U707 (N_707,In_1424,In_590);
nor U708 (N_708,In_840,In_651);
and U709 (N_709,In_395,In_865);
xnor U710 (N_710,In_156,In_199);
nor U711 (N_711,In_959,In_575);
or U712 (N_712,In_825,In_360);
xor U713 (N_713,In_1472,In_703);
xnor U714 (N_714,In_1030,In_832);
or U715 (N_715,In_1206,In_1270);
and U716 (N_716,In_134,In_59);
xor U717 (N_717,In_84,In_1415);
or U718 (N_718,In_309,In_1461);
xnor U719 (N_719,In_1127,In_1282);
or U720 (N_720,In_1072,In_866);
nor U721 (N_721,In_1076,In_1211);
and U722 (N_722,In_120,In_385);
and U723 (N_723,In_1339,In_342);
xor U724 (N_724,In_462,In_1164);
and U725 (N_725,In_949,In_404);
or U726 (N_726,In_1314,In_844);
and U727 (N_727,In_1374,In_1201);
xnor U728 (N_728,In_254,In_663);
nor U729 (N_729,In_994,In_987);
xor U730 (N_730,In_177,In_1487);
and U731 (N_731,In_273,In_56);
and U732 (N_732,In_20,In_308);
or U733 (N_733,In_668,In_4);
and U734 (N_734,In_1028,In_633);
xnor U735 (N_735,In_576,In_1062);
nor U736 (N_736,In_1273,In_323);
or U737 (N_737,In_102,In_1454);
or U738 (N_738,In_1245,In_1034);
nor U739 (N_739,In_1200,In_746);
and U740 (N_740,In_988,In_855);
nor U741 (N_741,In_520,In_984);
and U742 (N_742,In_157,In_353);
xnor U743 (N_743,In_503,In_225);
nor U744 (N_744,In_1202,In_944);
nand U745 (N_745,In_1251,In_207);
xnor U746 (N_746,In_792,In_1133);
and U747 (N_747,In_155,In_630);
and U748 (N_748,In_1476,In_1214);
and U749 (N_749,In_183,In_1307);
and U750 (N_750,In_159,In_715);
or U751 (N_751,In_252,In_796);
nand U752 (N_752,In_326,In_1343);
or U753 (N_753,In_833,In_179);
nand U754 (N_754,In_704,In_1244);
or U755 (N_755,In_438,In_458);
or U756 (N_756,In_1238,In_717);
xnor U757 (N_757,In_1291,In_165);
xnor U758 (N_758,In_771,In_1400);
and U759 (N_759,In_939,In_1270);
nand U760 (N_760,In_1473,In_1051);
and U761 (N_761,In_1400,In_878);
xnor U762 (N_762,In_1496,In_362);
nand U763 (N_763,In_991,In_1375);
or U764 (N_764,In_539,In_1393);
nor U765 (N_765,In_98,In_924);
and U766 (N_766,In_470,In_1483);
and U767 (N_767,In_1496,In_536);
xor U768 (N_768,In_987,In_1224);
nor U769 (N_769,In_992,In_1245);
and U770 (N_770,In_1477,In_799);
nand U771 (N_771,In_211,In_1271);
and U772 (N_772,In_1341,In_1261);
or U773 (N_773,In_1387,In_1451);
nor U774 (N_774,In_1449,In_1041);
xnor U775 (N_775,In_1027,In_317);
nor U776 (N_776,In_50,In_797);
and U777 (N_777,In_699,In_652);
and U778 (N_778,In_1448,In_857);
nand U779 (N_779,In_1303,In_1351);
and U780 (N_780,In_1381,In_90);
nand U781 (N_781,In_1468,In_1076);
nand U782 (N_782,In_829,In_815);
nand U783 (N_783,In_113,In_1352);
and U784 (N_784,In_1096,In_1494);
nor U785 (N_785,In_734,In_923);
nand U786 (N_786,In_1390,In_234);
nand U787 (N_787,In_902,In_741);
nand U788 (N_788,In_740,In_64);
nand U789 (N_789,In_856,In_728);
nor U790 (N_790,In_967,In_345);
nand U791 (N_791,In_969,In_463);
xor U792 (N_792,In_585,In_396);
and U793 (N_793,In_659,In_792);
or U794 (N_794,In_20,In_103);
or U795 (N_795,In_882,In_1136);
nand U796 (N_796,In_917,In_1152);
and U797 (N_797,In_322,In_405);
xnor U798 (N_798,In_762,In_112);
xnor U799 (N_799,In_957,In_1028);
nor U800 (N_800,In_593,In_908);
nand U801 (N_801,In_1013,In_278);
and U802 (N_802,In_165,In_516);
or U803 (N_803,In_727,In_57);
nand U804 (N_804,In_257,In_1193);
and U805 (N_805,In_510,In_1180);
xnor U806 (N_806,In_316,In_137);
nand U807 (N_807,In_1091,In_34);
nor U808 (N_808,In_573,In_319);
nor U809 (N_809,In_1484,In_424);
and U810 (N_810,In_1221,In_312);
and U811 (N_811,In_1305,In_625);
xnor U812 (N_812,In_1384,In_537);
and U813 (N_813,In_1339,In_1028);
nor U814 (N_814,In_794,In_1197);
and U815 (N_815,In_1183,In_145);
nor U816 (N_816,In_569,In_775);
nand U817 (N_817,In_566,In_225);
xnor U818 (N_818,In_608,In_919);
nand U819 (N_819,In_889,In_1130);
nor U820 (N_820,In_1271,In_562);
or U821 (N_821,In_253,In_712);
nand U822 (N_822,In_448,In_189);
xor U823 (N_823,In_326,In_1401);
and U824 (N_824,In_867,In_1317);
xnor U825 (N_825,In_1355,In_122);
xnor U826 (N_826,In_1408,In_202);
xor U827 (N_827,In_688,In_484);
nand U828 (N_828,In_1479,In_906);
or U829 (N_829,In_317,In_1498);
or U830 (N_830,In_613,In_993);
nor U831 (N_831,In_1095,In_680);
xor U832 (N_832,In_1264,In_827);
and U833 (N_833,In_873,In_1031);
xnor U834 (N_834,In_1121,In_325);
or U835 (N_835,In_1495,In_54);
nor U836 (N_836,In_244,In_25);
and U837 (N_837,In_942,In_651);
nor U838 (N_838,In_373,In_695);
nand U839 (N_839,In_279,In_1258);
xor U840 (N_840,In_1398,In_330);
and U841 (N_841,In_874,In_754);
nor U842 (N_842,In_1054,In_766);
nand U843 (N_843,In_1088,In_158);
xor U844 (N_844,In_886,In_450);
and U845 (N_845,In_805,In_574);
or U846 (N_846,In_833,In_484);
xor U847 (N_847,In_824,In_1409);
and U848 (N_848,In_147,In_1308);
nor U849 (N_849,In_19,In_185);
nand U850 (N_850,In_64,In_713);
or U851 (N_851,In_628,In_1184);
xor U852 (N_852,In_1190,In_1135);
nand U853 (N_853,In_809,In_574);
nand U854 (N_854,In_347,In_278);
nor U855 (N_855,In_710,In_299);
and U856 (N_856,In_210,In_687);
nand U857 (N_857,In_508,In_409);
xnor U858 (N_858,In_906,In_899);
nor U859 (N_859,In_880,In_1220);
nand U860 (N_860,In_702,In_1296);
nor U861 (N_861,In_1047,In_160);
xor U862 (N_862,In_1460,In_1105);
or U863 (N_863,In_346,In_956);
nand U864 (N_864,In_418,In_1492);
and U865 (N_865,In_320,In_881);
xor U866 (N_866,In_1081,In_537);
nor U867 (N_867,In_980,In_897);
xnor U868 (N_868,In_1125,In_814);
nand U869 (N_869,In_619,In_696);
xnor U870 (N_870,In_614,In_758);
and U871 (N_871,In_1323,In_415);
or U872 (N_872,In_141,In_1074);
or U873 (N_873,In_1179,In_533);
nand U874 (N_874,In_875,In_999);
and U875 (N_875,In_1343,In_1246);
or U876 (N_876,In_1446,In_1291);
or U877 (N_877,In_153,In_836);
and U878 (N_878,In_1136,In_1489);
nand U879 (N_879,In_107,In_129);
xnor U880 (N_880,In_64,In_1303);
or U881 (N_881,In_922,In_1331);
or U882 (N_882,In_1434,In_588);
nand U883 (N_883,In_1489,In_459);
nand U884 (N_884,In_1068,In_581);
or U885 (N_885,In_382,In_412);
and U886 (N_886,In_277,In_1071);
nand U887 (N_887,In_1373,In_701);
xor U888 (N_888,In_893,In_845);
nor U889 (N_889,In_1272,In_1476);
and U890 (N_890,In_782,In_83);
or U891 (N_891,In_1351,In_1430);
nand U892 (N_892,In_1263,In_1000);
and U893 (N_893,In_1193,In_1244);
or U894 (N_894,In_554,In_779);
and U895 (N_895,In_215,In_886);
or U896 (N_896,In_847,In_843);
nor U897 (N_897,In_827,In_716);
nor U898 (N_898,In_417,In_2);
nand U899 (N_899,In_1161,In_1372);
or U900 (N_900,In_394,In_1034);
or U901 (N_901,In_746,In_962);
nor U902 (N_902,In_173,In_835);
xor U903 (N_903,In_683,In_690);
nand U904 (N_904,In_493,In_901);
or U905 (N_905,In_1394,In_73);
nor U906 (N_906,In_688,In_671);
xnor U907 (N_907,In_713,In_565);
or U908 (N_908,In_629,In_931);
nand U909 (N_909,In_194,In_538);
xor U910 (N_910,In_1224,In_720);
or U911 (N_911,In_731,In_1009);
nor U912 (N_912,In_998,In_1375);
nand U913 (N_913,In_1006,In_228);
nor U914 (N_914,In_428,In_872);
xor U915 (N_915,In_321,In_1137);
xor U916 (N_916,In_761,In_385);
nand U917 (N_917,In_663,In_360);
or U918 (N_918,In_458,In_480);
xnor U919 (N_919,In_486,In_36);
nand U920 (N_920,In_318,In_1070);
xor U921 (N_921,In_888,In_323);
and U922 (N_922,In_188,In_722);
nor U923 (N_923,In_379,In_609);
or U924 (N_924,In_58,In_508);
nand U925 (N_925,In_4,In_453);
xnor U926 (N_926,In_282,In_1175);
nor U927 (N_927,In_1238,In_109);
nor U928 (N_928,In_585,In_317);
or U929 (N_929,In_101,In_799);
nor U930 (N_930,In_1364,In_221);
nand U931 (N_931,In_458,In_710);
and U932 (N_932,In_1082,In_662);
nand U933 (N_933,In_801,In_1180);
and U934 (N_934,In_1114,In_865);
nand U935 (N_935,In_1030,In_356);
nand U936 (N_936,In_1498,In_720);
and U937 (N_937,In_217,In_328);
nor U938 (N_938,In_39,In_622);
xnor U939 (N_939,In_418,In_765);
xor U940 (N_940,In_629,In_1049);
and U941 (N_941,In_108,In_1271);
and U942 (N_942,In_831,In_130);
and U943 (N_943,In_1023,In_910);
nand U944 (N_944,In_175,In_340);
nor U945 (N_945,In_1406,In_693);
nand U946 (N_946,In_518,In_1112);
nor U947 (N_947,In_927,In_10);
xnor U948 (N_948,In_86,In_159);
nand U949 (N_949,In_667,In_795);
and U950 (N_950,In_731,In_1297);
and U951 (N_951,In_396,In_1258);
nor U952 (N_952,In_364,In_1273);
xnor U953 (N_953,In_936,In_1193);
xnor U954 (N_954,In_1351,In_372);
and U955 (N_955,In_1114,In_1266);
nand U956 (N_956,In_195,In_1422);
nand U957 (N_957,In_65,In_120);
xnor U958 (N_958,In_1295,In_960);
nor U959 (N_959,In_1179,In_1499);
xnor U960 (N_960,In_207,In_449);
nand U961 (N_961,In_938,In_1231);
xnor U962 (N_962,In_233,In_445);
and U963 (N_963,In_1305,In_1245);
nand U964 (N_964,In_1309,In_1178);
nand U965 (N_965,In_75,In_1241);
xor U966 (N_966,In_1000,In_56);
nand U967 (N_967,In_1244,In_618);
nor U968 (N_968,In_1027,In_86);
and U969 (N_969,In_1324,In_960);
nand U970 (N_970,In_113,In_151);
xnor U971 (N_971,In_1338,In_794);
xnor U972 (N_972,In_1153,In_259);
or U973 (N_973,In_1091,In_1356);
xnor U974 (N_974,In_395,In_1246);
xor U975 (N_975,In_550,In_1457);
nor U976 (N_976,In_1110,In_797);
and U977 (N_977,In_925,In_802);
or U978 (N_978,In_737,In_693);
or U979 (N_979,In_1329,In_1134);
and U980 (N_980,In_597,In_146);
xnor U981 (N_981,In_430,In_1324);
xor U982 (N_982,In_1433,In_131);
nor U983 (N_983,In_482,In_36);
or U984 (N_984,In_1399,In_628);
xor U985 (N_985,In_320,In_1222);
nor U986 (N_986,In_152,In_508);
nand U987 (N_987,In_934,In_269);
nand U988 (N_988,In_1163,In_1361);
or U989 (N_989,In_412,In_525);
xor U990 (N_990,In_580,In_120);
nor U991 (N_991,In_1241,In_1482);
nor U992 (N_992,In_38,In_19);
nand U993 (N_993,In_1408,In_807);
or U994 (N_994,In_1372,In_913);
xor U995 (N_995,In_164,In_627);
xor U996 (N_996,In_623,In_814);
nor U997 (N_997,In_397,In_770);
nor U998 (N_998,In_1019,In_723);
nand U999 (N_999,In_917,In_1268);
nand U1000 (N_1000,In_725,In_74);
nor U1001 (N_1001,In_1118,In_353);
nor U1002 (N_1002,In_875,In_565);
or U1003 (N_1003,In_1290,In_528);
nand U1004 (N_1004,In_1153,In_865);
and U1005 (N_1005,In_233,In_1214);
nand U1006 (N_1006,In_1049,In_823);
and U1007 (N_1007,In_1138,In_108);
nand U1008 (N_1008,In_800,In_417);
nand U1009 (N_1009,In_714,In_991);
xor U1010 (N_1010,In_1123,In_510);
nor U1011 (N_1011,In_1410,In_643);
nor U1012 (N_1012,In_276,In_271);
nand U1013 (N_1013,In_322,In_10);
xor U1014 (N_1014,In_577,In_867);
xnor U1015 (N_1015,In_92,In_803);
or U1016 (N_1016,In_887,In_309);
and U1017 (N_1017,In_571,In_1414);
nor U1018 (N_1018,In_1296,In_564);
xnor U1019 (N_1019,In_1079,In_1485);
xor U1020 (N_1020,In_1292,In_198);
and U1021 (N_1021,In_967,In_538);
xor U1022 (N_1022,In_607,In_820);
xnor U1023 (N_1023,In_84,In_9);
and U1024 (N_1024,In_1183,In_876);
or U1025 (N_1025,In_482,In_507);
xnor U1026 (N_1026,In_726,In_89);
and U1027 (N_1027,In_957,In_84);
or U1028 (N_1028,In_70,In_1221);
xor U1029 (N_1029,In_126,In_1431);
nand U1030 (N_1030,In_149,In_349);
nand U1031 (N_1031,In_373,In_455);
xor U1032 (N_1032,In_869,In_736);
nor U1033 (N_1033,In_943,In_731);
nor U1034 (N_1034,In_538,In_643);
xor U1035 (N_1035,In_1317,In_48);
and U1036 (N_1036,In_467,In_1207);
nor U1037 (N_1037,In_1338,In_1400);
or U1038 (N_1038,In_984,In_893);
or U1039 (N_1039,In_881,In_751);
nand U1040 (N_1040,In_1115,In_1429);
nand U1041 (N_1041,In_1341,In_123);
nor U1042 (N_1042,In_510,In_1394);
xnor U1043 (N_1043,In_632,In_641);
nor U1044 (N_1044,In_1162,In_1393);
nand U1045 (N_1045,In_932,In_962);
nor U1046 (N_1046,In_1050,In_841);
nand U1047 (N_1047,In_145,In_845);
and U1048 (N_1048,In_459,In_1282);
nand U1049 (N_1049,In_647,In_82);
xor U1050 (N_1050,In_221,In_322);
nand U1051 (N_1051,In_553,In_912);
nor U1052 (N_1052,In_112,In_1458);
or U1053 (N_1053,In_437,In_1262);
nor U1054 (N_1054,In_847,In_291);
xor U1055 (N_1055,In_97,In_62);
and U1056 (N_1056,In_1086,In_36);
xnor U1057 (N_1057,In_487,In_414);
xor U1058 (N_1058,In_840,In_1208);
xor U1059 (N_1059,In_196,In_685);
xnor U1060 (N_1060,In_746,In_523);
nand U1061 (N_1061,In_1248,In_838);
and U1062 (N_1062,In_966,In_263);
and U1063 (N_1063,In_856,In_589);
nor U1064 (N_1064,In_461,In_189);
or U1065 (N_1065,In_580,In_28);
nor U1066 (N_1066,In_275,In_34);
and U1067 (N_1067,In_1069,In_995);
and U1068 (N_1068,In_513,In_975);
xor U1069 (N_1069,In_648,In_326);
or U1070 (N_1070,In_466,In_153);
xor U1071 (N_1071,In_945,In_324);
or U1072 (N_1072,In_545,In_411);
xor U1073 (N_1073,In_729,In_695);
or U1074 (N_1074,In_1413,In_1006);
xor U1075 (N_1075,In_588,In_433);
and U1076 (N_1076,In_169,In_135);
or U1077 (N_1077,In_779,In_516);
nand U1078 (N_1078,In_1260,In_1268);
nor U1079 (N_1079,In_688,In_1265);
and U1080 (N_1080,In_1087,In_1112);
nand U1081 (N_1081,In_266,In_1435);
nor U1082 (N_1082,In_1331,In_1048);
xor U1083 (N_1083,In_307,In_409);
nor U1084 (N_1084,In_1095,In_331);
or U1085 (N_1085,In_1020,In_754);
or U1086 (N_1086,In_376,In_845);
or U1087 (N_1087,In_1174,In_1344);
nor U1088 (N_1088,In_189,In_801);
and U1089 (N_1089,In_856,In_1189);
xor U1090 (N_1090,In_1326,In_1222);
nand U1091 (N_1091,In_29,In_1327);
nor U1092 (N_1092,In_1456,In_1251);
xnor U1093 (N_1093,In_851,In_1029);
xnor U1094 (N_1094,In_537,In_1342);
xnor U1095 (N_1095,In_328,In_157);
or U1096 (N_1096,In_0,In_653);
nor U1097 (N_1097,In_732,In_317);
or U1098 (N_1098,In_965,In_1258);
xnor U1099 (N_1099,In_15,In_1186);
xnor U1100 (N_1100,In_974,In_712);
nor U1101 (N_1101,In_1282,In_812);
and U1102 (N_1102,In_510,In_1153);
nand U1103 (N_1103,In_939,In_1487);
or U1104 (N_1104,In_1402,In_1475);
xor U1105 (N_1105,In_455,In_1498);
nand U1106 (N_1106,In_1461,In_1356);
nand U1107 (N_1107,In_75,In_733);
nor U1108 (N_1108,In_773,In_911);
nand U1109 (N_1109,In_846,In_1340);
nor U1110 (N_1110,In_677,In_310);
xor U1111 (N_1111,In_47,In_529);
and U1112 (N_1112,In_984,In_586);
nand U1113 (N_1113,In_835,In_685);
nor U1114 (N_1114,In_673,In_377);
nand U1115 (N_1115,In_779,In_366);
or U1116 (N_1116,In_1005,In_1191);
and U1117 (N_1117,In_1098,In_1166);
or U1118 (N_1118,In_869,In_516);
and U1119 (N_1119,In_1080,In_1142);
or U1120 (N_1120,In_690,In_527);
or U1121 (N_1121,In_1188,In_427);
or U1122 (N_1122,In_531,In_1169);
nand U1123 (N_1123,In_398,In_523);
or U1124 (N_1124,In_5,In_1294);
or U1125 (N_1125,In_1230,In_1100);
and U1126 (N_1126,In_1132,In_931);
xor U1127 (N_1127,In_1290,In_1158);
nand U1128 (N_1128,In_561,In_425);
xnor U1129 (N_1129,In_1095,In_436);
nand U1130 (N_1130,In_814,In_157);
nor U1131 (N_1131,In_1206,In_1031);
nand U1132 (N_1132,In_108,In_788);
nand U1133 (N_1133,In_1400,In_1193);
xnor U1134 (N_1134,In_87,In_898);
or U1135 (N_1135,In_1411,In_3);
and U1136 (N_1136,In_966,In_709);
and U1137 (N_1137,In_508,In_187);
nand U1138 (N_1138,In_621,In_305);
nor U1139 (N_1139,In_1003,In_1374);
and U1140 (N_1140,In_107,In_1126);
xnor U1141 (N_1141,In_427,In_337);
xnor U1142 (N_1142,In_367,In_989);
or U1143 (N_1143,In_382,In_217);
or U1144 (N_1144,In_475,In_126);
and U1145 (N_1145,In_329,In_94);
nand U1146 (N_1146,In_62,In_882);
or U1147 (N_1147,In_451,In_1180);
and U1148 (N_1148,In_21,In_133);
nor U1149 (N_1149,In_1328,In_1134);
xor U1150 (N_1150,In_1450,In_164);
or U1151 (N_1151,In_1174,In_1076);
xnor U1152 (N_1152,In_1398,In_858);
xor U1153 (N_1153,In_1455,In_1398);
xor U1154 (N_1154,In_344,In_324);
nor U1155 (N_1155,In_1417,In_1085);
or U1156 (N_1156,In_18,In_1010);
xnor U1157 (N_1157,In_1158,In_48);
nor U1158 (N_1158,In_728,In_756);
and U1159 (N_1159,In_402,In_182);
nand U1160 (N_1160,In_450,In_1409);
nor U1161 (N_1161,In_606,In_1244);
nor U1162 (N_1162,In_432,In_703);
nand U1163 (N_1163,In_271,In_273);
or U1164 (N_1164,In_302,In_923);
or U1165 (N_1165,In_942,In_1340);
and U1166 (N_1166,In_924,In_528);
nand U1167 (N_1167,In_483,In_79);
xor U1168 (N_1168,In_172,In_295);
and U1169 (N_1169,In_191,In_1045);
xnor U1170 (N_1170,In_950,In_916);
or U1171 (N_1171,In_405,In_1163);
nor U1172 (N_1172,In_276,In_352);
and U1173 (N_1173,In_991,In_1087);
nand U1174 (N_1174,In_220,In_1337);
and U1175 (N_1175,In_1056,In_231);
or U1176 (N_1176,In_1236,In_469);
xnor U1177 (N_1177,In_52,In_646);
or U1178 (N_1178,In_456,In_60);
and U1179 (N_1179,In_1217,In_6);
or U1180 (N_1180,In_785,In_207);
nor U1181 (N_1181,In_946,In_1042);
or U1182 (N_1182,In_245,In_1459);
xnor U1183 (N_1183,In_1494,In_513);
xor U1184 (N_1184,In_292,In_1099);
or U1185 (N_1185,In_1166,In_319);
and U1186 (N_1186,In_947,In_1218);
and U1187 (N_1187,In_845,In_1049);
or U1188 (N_1188,In_498,In_1271);
xnor U1189 (N_1189,In_522,In_1177);
xor U1190 (N_1190,In_888,In_528);
xnor U1191 (N_1191,In_243,In_1227);
and U1192 (N_1192,In_1354,In_25);
nor U1193 (N_1193,In_705,In_410);
or U1194 (N_1194,In_683,In_771);
or U1195 (N_1195,In_1032,In_1444);
nand U1196 (N_1196,In_1212,In_1250);
nand U1197 (N_1197,In_1237,In_191);
xor U1198 (N_1198,In_1351,In_146);
or U1199 (N_1199,In_1058,In_844);
nor U1200 (N_1200,In_192,In_961);
nor U1201 (N_1201,In_589,In_382);
nand U1202 (N_1202,In_1114,In_407);
nor U1203 (N_1203,In_546,In_889);
or U1204 (N_1204,In_145,In_832);
or U1205 (N_1205,In_426,In_944);
nor U1206 (N_1206,In_454,In_1118);
nand U1207 (N_1207,In_728,In_1166);
nand U1208 (N_1208,In_63,In_207);
nand U1209 (N_1209,In_1172,In_171);
or U1210 (N_1210,In_569,In_1192);
nor U1211 (N_1211,In_872,In_849);
xnor U1212 (N_1212,In_175,In_1424);
and U1213 (N_1213,In_126,In_827);
nor U1214 (N_1214,In_692,In_962);
nand U1215 (N_1215,In_787,In_322);
xor U1216 (N_1216,In_1413,In_660);
or U1217 (N_1217,In_393,In_67);
nor U1218 (N_1218,In_871,In_47);
xnor U1219 (N_1219,In_1449,In_224);
or U1220 (N_1220,In_880,In_558);
and U1221 (N_1221,In_630,In_792);
nor U1222 (N_1222,In_1440,In_895);
nand U1223 (N_1223,In_1226,In_1065);
and U1224 (N_1224,In_524,In_1384);
nor U1225 (N_1225,In_1055,In_366);
or U1226 (N_1226,In_103,In_1473);
nand U1227 (N_1227,In_80,In_976);
and U1228 (N_1228,In_895,In_1367);
or U1229 (N_1229,In_489,In_1139);
nor U1230 (N_1230,In_1075,In_1045);
nor U1231 (N_1231,In_450,In_522);
nor U1232 (N_1232,In_37,In_1347);
or U1233 (N_1233,In_1354,In_688);
nand U1234 (N_1234,In_427,In_567);
nor U1235 (N_1235,In_0,In_655);
and U1236 (N_1236,In_935,In_198);
and U1237 (N_1237,In_820,In_1054);
nor U1238 (N_1238,In_1458,In_453);
xnor U1239 (N_1239,In_483,In_729);
xnor U1240 (N_1240,In_108,In_130);
or U1241 (N_1241,In_1166,In_1084);
nand U1242 (N_1242,In_1310,In_1149);
xnor U1243 (N_1243,In_610,In_682);
nand U1244 (N_1244,In_711,In_1406);
and U1245 (N_1245,In_130,In_246);
or U1246 (N_1246,In_1003,In_879);
xnor U1247 (N_1247,In_171,In_849);
and U1248 (N_1248,In_214,In_657);
and U1249 (N_1249,In_1435,In_1082);
nor U1250 (N_1250,In_1127,In_703);
and U1251 (N_1251,In_525,In_438);
or U1252 (N_1252,In_559,In_278);
and U1253 (N_1253,In_639,In_1443);
nor U1254 (N_1254,In_806,In_823);
and U1255 (N_1255,In_835,In_751);
xor U1256 (N_1256,In_1393,In_1365);
and U1257 (N_1257,In_763,In_1041);
xor U1258 (N_1258,In_1017,In_925);
or U1259 (N_1259,In_921,In_37);
or U1260 (N_1260,In_1310,In_33);
nor U1261 (N_1261,In_1205,In_208);
or U1262 (N_1262,In_675,In_39);
nand U1263 (N_1263,In_1007,In_692);
nand U1264 (N_1264,In_1213,In_604);
nor U1265 (N_1265,In_1360,In_1424);
nand U1266 (N_1266,In_1370,In_180);
and U1267 (N_1267,In_1472,In_353);
and U1268 (N_1268,In_67,In_99);
or U1269 (N_1269,In_187,In_254);
nor U1270 (N_1270,In_1076,In_1173);
or U1271 (N_1271,In_1361,In_1434);
xor U1272 (N_1272,In_787,In_1120);
xor U1273 (N_1273,In_664,In_1142);
or U1274 (N_1274,In_778,In_590);
and U1275 (N_1275,In_383,In_532);
nor U1276 (N_1276,In_684,In_1098);
nand U1277 (N_1277,In_1017,In_389);
nor U1278 (N_1278,In_39,In_939);
and U1279 (N_1279,In_222,In_81);
or U1280 (N_1280,In_131,In_122);
nand U1281 (N_1281,In_157,In_620);
or U1282 (N_1282,In_1488,In_946);
nor U1283 (N_1283,In_493,In_419);
and U1284 (N_1284,In_1143,In_24);
and U1285 (N_1285,In_373,In_959);
or U1286 (N_1286,In_815,In_590);
nand U1287 (N_1287,In_767,In_1383);
or U1288 (N_1288,In_1223,In_410);
nor U1289 (N_1289,In_454,In_1042);
nor U1290 (N_1290,In_571,In_1350);
xnor U1291 (N_1291,In_822,In_965);
and U1292 (N_1292,In_636,In_921);
nor U1293 (N_1293,In_1257,In_1084);
nand U1294 (N_1294,In_255,In_1025);
xnor U1295 (N_1295,In_1226,In_303);
nand U1296 (N_1296,In_1268,In_491);
and U1297 (N_1297,In_978,In_1081);
and U1298 (N_1298,In_1470,In_983);
and U1299 (N_1299,In_627,In_44);
or U1300 (N_1300,In_0,In_489);
and U1301 (N_1301,In_1086,In_1123);
nand U1302 (N_1302,In_166,In_688);
xor U1303 (N_1303,In_47,In_1018);
and U1304 (N_1304,In_1463,In_985);
nand U1305 (N_1305,In_426,In_499);
or U1306 (N_1306,In_1156,In_1432);
nor U1307 (N_1307,In_988,In_195);
or U1308 (N_1308,In_707,In_1064);
nand U1309 (N_1309,In_926,In_242);
nor U1310 (N_1310,In_138,In_146);
and U1311 (N_1311,In_551,In_1426);
or U1312 (N_1312,In_444,In_395);
xor U1313 (N_1313,In_1080,In_436);
and U1314 (N_1314,In_796,In_754);
or U1315 (N_1315,In_44,In_1475);
and U1316 (N_1316,In_1271,In_576);
and U1317 (N_1317,In_580,In_211);
nor U1318 (N_1318,In_204,In_249);
or U1319 (N_1319,In_156,In_411);
nor U1320 (N_1320,In_991,In_924);
nand U1321 (N_1321,In_605,In_407);
and U1322 (N_1322,In_1377,In_1180);
nand U1323 (N_1323,In_1040,In_1354);
or U1324 (N_1324,In_1238,In_75);
nand U1325 (N_1325,In_1243,In_1314);
nor U1326 (N_1326,In_1173,In_676);
nor U1327 (N_1327,In_921,In_592);
and U1328 (N_1328,In_1211,In_1266);
or U1329 (N_1329,In_1384,In_143);
and U1330 (N_1330,In_13,In_288);
nand U1331 (N_1331,In_497,In_233);
or U1332 (N_1332,In_482,In_450);
nor U1333 (N_1333,In_1241,In_565);
nor U1334 (N_1334,In_1426,In_1053);
and U1335 (N_1335,In_1293,In_796);
nor U1336 (N_1336,In_716,In_1334);
nand U1337 (N_1337,In_1282,In_1025);
or U1338 (N_1338,In_577,In_647);
xnor U1339 (N_1339,In_1251,In_284);
nand U1340 (N_1340,In_809,In_589);
xor U1341 (N_1341,In_207,In_512);
nor U1342 (N_1342,In_1027,In_996);
xor U1343 (N_1343,In_994,In_357);
or U1344 (N_1344,In_1232,In_373);
xnor U1345 (N_1345,In_1114,In_476);
and U1346 (N_1346,In_1217,In_1148);
nand U1347 (N_1347,In_1136,In_95);
nor U1348 (N_1348,In_984,In_504);
and U1349 (N_1349,In_1110,In_1103);
xor U1350 (N_1350,In_820,In_293);
nand U1351 (N_1351,In_1038,In_113);
xnor U1352 (N_1352,In_73,In_1018);
nand U1353 (N_1353,In_1173,In_104);
nand U1354 (N_1354,In_1415,In_1303);
or U1355 (N_1355,In_563,In_700);
xor U1356 (N_1356,In_1272,In_979);
nand U1357 (N_1357,In_1275,In_537);
and U1358 (N_1358,In_1155,In_1055);
nand U1359 (N_1359,In_922,In_1174);
nor U1360 (N_1360,In_281,In_188);
nor U1361 (N_1361,In_357,In_733);
nor U1362 (N_1362,In_1187,In_700);
and U1363 (N_1363,In_1421,In_1068);
and U1364 (N_1364,In_815,In_1435);
nor U1365 (N_1365,In_537,In_254);
or U1366 (N_1366,In_613,In_670);
or U1367 (N_1367,In_296,In_1219);
nor U1368 (N_1368,In_359,In_487);
or U1369 (N_1369,In_772,In_1427);
and U1370 (N_1370,In_466,In_1450);
or U1371 (N_1371,In_358,In_724);
or U1372 (N_1372,In_1488,In_64);
or U1373 (N_1373,In_1464,In_310);
nor U1374 (N_1374,In_869,In_194);
and U1375 (N_1375,In_1072,In_1467);
and U1376 (N_1376,In_703,In_150);
or U1377 (N_1377,In_852,In_1062);
or U1378 (N_1378,In_614,In_769);
and U1379 (N_1379,In_1405,In_922);
nand U1380 (N_1380,In_83,In_1102);
nand U1381 (N_1381,In_92,In_1463);
and U1382 (N_1382,In_328,In_949);
nor U1383 (N_1383,In_644,In_38);
or U1384 (N_1384,In_583,In_974);
or U1385 (N_1385,In_759,In_279);
and U1386 (N_1386,In_605,In_666);
xnor U1387 (N_1387,In_15,In_1430);
nand U1388 (N_1388,In_724,In_651);
and U1389 (N_1389,In_264,In_1270);
nand U1390 (N_1390,In_922,In_506);
and U1391 (N_1391,In_871,In_1235);
or U1392 (N_1392,In_580,In_439);
nand U1393 (N_1393,In_500,In_1463);
nor U1394 (N_1394,In_406,In_121);
xor U1395 (N_1395,In_1323,In_520);
and U1396 (N_1396,In_40,In_1252);
nand U1397 (N_1397,In_1014,In_1354);
nor U1398 (N_1398,In_359,In_1078);
nor U1399 (N_1399,In_431,In_796);
or U1400 (N_1400,In_908,In_873);
nor U1401 (N_1401,In_1056,In_137);
or U1402 (N_1402,In_466,In_824);
or U1403 (N_1403,In_1193,In_753);
nand U1404 (N_1404,In_1284,In_1164);
nand U1405 (N_1405,In_492,In_8);
xnor U1406 (N_1406,In_852,In_920);
and U1407 (N_1407,In_702,In_200);
xor U1408 (N_1408,In_857,In_1084);
nor U1409 (N_1409,In_659,In_503);
or U1410 (N_1410,In_1439,In_73);
nand U1411 (N_1411,In_317,In_304);
nor U1412 (N_1412,In_412,In_26);
xor U1413 (N_1413,In_1001,In_971);
xor U1414 (N_1414,In_756,In_578);
xor U1415 (N_1415,In_909,In_590);
xnor U1416 (N_1416,In_220,In_810);
xor U1417 (N_1417,In_618,In_1058);
and U1418 (N_1418,In_404,In_29);
xnor U1419 (N_1419,In_69,In_793);
or U1420 (N_1420,In_1085,In_129);
and U1421 (N_1421,In_768,In_355);
or U1422 (N_1422,In_1363,In_1393);
and U1423 (N_1423,In_1351,In_421);
nor U1424 (N_1424,In_972,In_997);
or U1425 (N_1425,In_229,In_785);
nor U1426 (N_1426,In_802,In_646);
or U1427 (N_1427,In_1387,In_294);
nor U1428 (N_1428,In_1466,In_1109);
or U1429 (N_1429,In_431,In_1375);
nand U1430 (N_1430,In_709,In_293);
xnor U1431 (N_1431,In_929,In_773);
nand U1432 (N_1432,In_568,In_137);
xor U1433 (N_1433,In_1327,In_1013);
xor U1434 (N_1434,In_656,In_1295);
xnor U1435 (N_1435,In_839,In_232);
and U1436 (N_1436,In_475,In_1409);
nor U1437 (N_1437,In_414,In_842);
xor U1438 (N_1438,In_797,In_453);
xnor U1439 (N_1439,In_665,In_268);
or U1440 (N_1440,In_1130,In_603);
nand U1441 (N_1441,In_189,In_555);
xor U1442 (N_1442,In_769,In_188);
or U1443 (N_1443,In_208,In_1416);
xnor U1444 (N_1444,In_1365,In_94);
or U1445 (N_1445,In_1171,In_360);
and U1446 (N_1446,In_52,In_398);
nand U1447 (N_1447,In_1006,In_184);
nand U1448 (N_1448,In_841,In_1498);
or U1449 (N_1449,In_347,In_132);
nor U1450 (N_1450,In_793,In_341);
and U1451 (N_1451,In_624,In_1346);
or U1452 (N_1452,In_1116,In_1144);
nor U1453 (N_1453,In_749,In_475);
nor U1454 (N_1454,In_936,In_289);
or U1455 (N_1455,In_1184,In_982);
and U1456 (N_1456,In_741,In_1214);
or U1457 (N_1457,In_313,In_990);
or U1458 (N_1458,In_755,In_1303);
nor U1459 (N_1459,In_591,In_551);
xnor U1460 (N_1460,In_488,In_146);
and U1461 (N_1461,In_384,In_24);
xor U1462 (N_1462,In_1248,In_1252);
xor U1463 (N_1463,In_881,In_230);
nor U1464 (N_1464,In_1194,In_320);
nor U1465 (N_1465,In_1256,In_631);
nand U1466 (N_1466,In_578,In_274);
nand U1467 (N_1467,In_1366,In_657);
or U1468 (N_1468,In_1438,In_1102);
and U1469 (N_1469,In_485,In_1194);
or U1470 (N_1470,In_1428,In_38);
and U1471 (N_1471,In_141,In_1256);
nand U1472 (N_1472,In_1171,In_1080);
or U1473 (N_1473,In_976,In_151);
xnor U1474 (N_1474,In_907,In_754);
and U1475 (N_1475,In_363,In_1366);
nand U1476 (N_1476,In_697,In_463);
xnor U1477 (N_1477,In_1311,In_301);
xnor U1478 (N_1478,In_204,In_1121);
xnor U1479 (N_1479,In_626,In_1363);
and U1480 (N_1480,In_920,In_289);
xnor U1481 (N_1481,In_520,In_1401);
nand U1482 (N_1482,In_331,In_859);
nor U1483 (N_1483,In_868,In_727);
nand U1484 (N_1484,In_296,In_1158);
nor U1485 (N_1485,In_958,In_72);
nor U1486 (N_1486,In_370,In_1146);
nand U1487 (N_1487,In_1045,In_819);
xnor U1488 (N_1488,In_699,In_1360);
and U1489 (N_1489,In_805,In_1090);
and U1490 (N_1490,In_1336,In_1268);
nor U1491 (N_1491,In_250,In_267);
nand U1492 (N_1492,In_173,In_83);
xnor U1493 (N_1493,In_879,In_713);
nand U1494 (N_1494,In_416,In_336);
xnor U1495 (N_1495,In_1222,In_1228);
or U1496 (N_1496,In_665,In_1087);
or U1497 (N_1497,In_763,In_709);
nor U1498 (N_1498,In_930,In_1479);
nor U1499 (N_1499,In_1068,In_504);
nor U1500 (N_1500,N_607,N_440);
nor U1501 (N_1501,N_617,N_1357);
xor U1502 (N_1502,N_1481,N_411);
nor U1503 (N_1503,N_1423,N_809);
nor U1504 (N_1504,N_1338,N_693);
and U1505 (N_1505,N_1383,N_1415);
and U1506 (N_1506,N_793,N_293);
or U1507 (N_1507,N_787,N_894);
and U1508 (N_1508,N_109,N_111);
and U1509 (N_1509,N_1056,N_1018);
xnor U1510 (N_1510,N_123,N_19);
and U1511 (N_1511,N_813,N_26);
nand U1512 (N_1512,N_1323,N_1327);
nor U1513 (N_1513,N_657,N_1216);
nor U1514 (N_1514,N_135,N_196);
nand U1515 (N_1515,N_997,N_772);
xnor U1516 (N_1516,N_41,N_225);
and U1517 (N_1517,N_1090,N_1226);
or U1518 (N_1518,N_419,N_927);
and U1519 (N_1519,N_391,N_1259);
xor U1520 (N_1520,N_1012,N_403);
and U1521 (N_1521,N_78,N_471);
or U1522 (N_1522,N_1159,N_1104);
xor U1523 (N_1523,N_1266,N_25);
xor U1524 (N_1524,N_1322,N_550);
or U1525 (N_1525,N_500,N_1485);
and U1526 (N_1526,N_838,N_1275);
nor U1527 (N_1527,N_697,N_567);
nand U1528 (N_1528,N_1167,N_475);
and U1529 (N_1529,N_1034,N_1010);
or U1530 (N_1530,N_522,N_1047);
nand U1531 (N_1531,N_844,N_138);
or U1532 (N_1532,N_1042,N_81);
xnor U1533 (N_1533,N_990,N_794);
nand U1534 (N_1534,N_1094,N_1249);
or U1535 (N_1535,N_769,N_387);
or U1536 (N_1536,N_959,N_253);
and U1537 (N_1537,N_18,N_728);
xnor U1538 (N_1538,N_145,N_1314);
nand U1539 (N_1539,N_9,N_1483);
nand U1540 (N_1540,N_1494,N_47);
nand U1541 (N_1541,N_513,N_712);
nor U1542 (N_1542,N_117,N_296);
and U1543 (N_1543,N_1247,N_540);
nand U1544 (N_1544,N_854,N_1022);
nand U1545 (N_1545,N_238,N_953);
nand U1546 (N_1546,N_1472,N_662);
and U1547 (N_1547,N_666,N_1121);
xnor U1548 (N_1548,N_863,N_300);
nand U1549 (N_1549,N_1442,N_1148);
xor U1550 (N_1550,N_966,N_823);
and U1551 (N_1551,N_1214,N_636);
nand U1552 (N_1552,N_1025,N_1120);
xor U1553 (N_1553,N_1113,N_731);
and U1554 (N_1554,N_1039,N_64);
nand U1555 (N_1555,N_1342,N_786);
nor U1556 (N_1556,N_620,N_531);
or U1557 (N_1557,N_1172,N_97);
nor U1558 (N_1558,N_327,N_1096);
xnor U1559 (N_1559,N_398,N_874);
nand U1560 (N_1560,N_736,N_1246);
nor U1561 (N_1561,N_907,N_777);
nor U1562 (N_1562,N_237,N_981);
xnor U1563 (N_1563,N_124,N_158);
xor U1564 (N_1564,N_750,N_1245);
nand U1565 (N_1565,N_416,N_1397);
xor U1566 (N_1566,N_1013,N_877);
or U1567 (N_1567,N_675,N_687);
nor U1568 (N_1568,N_606,N_886);
nand U1569 (N_1569,N_190,N_744);
nor U1570 (N_1570,N_1287,N_696);
xnor U1571 (N_1571,N_1065,N_553);
xnor U1572 (N_1572,N_1142,N_388);
nor U1573 (N_1573,N_951,N_182);
or U1574 (N_1574,N_1345,N_956);
nor U1575 (N_1575,N_1452,N_827);
xor U1576 (N_1576,N_773,N_1054);
xor U1577 (N_1577,N_1382,N_417);
nor U1578 (N_1578,N_458,N_312);
or U1579 (N_1579,N_477,N_702);
xor U1580 (N_1580,N_1294,N_1241);
nor U1581 (N_1581,N_77,N_33);
and U1582 (N_1582,N_895,N_1036);
nand U1583 (N_1583,N_1264,N_861);
or U1584 (N_1584,N_1321,N_1146);
xnor U1585 (N_1585,N_1340,N_940);
and U1586 (N_1586,N_1370,N_992);
nand U1587 (N_1587,N_1369,N_737);
nand U1588 (N_1588,N_1453,N_1414);
nor U1589 (N_1589,N_942,N_1169);
xor U1590 (N_1590,N_324,N_795);
and U1591 (N_1591,N_911,N_1476);
and U1592 (N_1592,N_1011,N_229);
nor U1593 (N_1593,N_441,N_654);
or U1594 (N_1594,N_1209,N_244);
xor U1595 (N_1595,N_1285,N_1400);
or U1596 (N_1596,N_235,N_472);
nor U1597 (N_1597,N_367,N_316);
xnor U1598 (N_1598,N_92,N_671);
or U1599 (N_1599,N_539,N_1071);
or U1600 (N_1600,N_264,N_674);
xnor U1601 (N_1601,N_516,N_122);
or U1602 (N_1602,N_1231,N_962);
or U1603 (N_1603,N_605,N_514);
xor U1604 (N_1604,N_105,N_684);
nor U1605 (N_1605,N_964,N_1250);
nand U1606 (N_1606,N_984,N_554);
nor U1607 (N_1607,N_202,N_217);
xor U1608 (N_1608,N_1390,N_711);
or U1609 (N_1609,N_670,N_851);
or U1610 (N_1610,N_1398,N_385);
nand U1611 (N_1611,N_564,N_914);
xor U1612 (N_1612,N_859,N_631);
xor U1613 (N_1613,N_30,N_192);
and U1614 (N_1614,N_1229,N_379);
xnor U1615 (N_1615,N_855,N_1161);
nand U1616 (N_1616,N_457,N_360);
nand U1617 (N_1617,N_1269,N_936);
nand U1618 (N_1618,N_1286,N_286);
nand U1619 (N_1619,N_35,N_1057);
nor U1620 (N_1620,N_783,N_1242);
nand U1621 (N_1621,N_396,N_447);
and U1622 (N_1622,N_302,N_604);
nor U1623 (N_1623,N_1032,N_893);
nand U1624 (N_1624,N_969,N_1461);
nor U1625 (N_1625,N_985,N_224);
nor U1626 (N_1626,N_162,N_1131);
nand U1627 (N_1627,N_600,N_1111);
and U1628 (N_1628,N_107,N_252);
xnor U1629 (N_1629,N_128,N_856);
nand U1630 (N_1630,N_902,N_713);
and U1631 (N_1631,N_1473,N_198);
nor U1632 (N_1632,N_478,N_717);
and U1633 (N_1633,N_31,N_796);
or U1634 (N_1634,N_944,N_623);
nand U1635 (N_1635,N_1134,N_1464);
nand U1636 (N_1636,N_1387,N_336);
nor U1637 (N_1637,N_347,N_1435);
and U1638 (N_1638,N_114,N_1225);
or U1639 (N_1639,N_493,N_341);
and U1640 (N_1640,N_80,N_928);
nand U1641 (N_1641,N_578,N_1312);
nand U1642 (N_1642,N_807,N_402);
xnor U1643 (N_1643,N_1459,N_200);
nand U1644 (N_1644,N_950,N_948);
and U1645 (N_1645,N_1067,N_1425);
xnor U1646 (N_1646,N_1355,N_1081);
xnor U1647 (N_1647,N_1206,N_38);
nor U1648 (N_1648,N_113,N_186);
and U1649 (N_1649,N_209,N_1135);
xnor U1650 (N_1650,N_259,N_1046);
xor U1651 (N_1651,N_1300,N_467);
nor U1652 (N_1652,N_588,N_837);
xor U1653 (N_1653,N_742,N_1353);
and U1654 (N_1654,N_414,N_1221);
or U1655 (N_1655,N_570,N_504);
nand U1656 (N_1656,N_183,N_497);
and U1657 (N_1657,N_401,N_487);
nand U1658 (N_1658,N_1208,N_133);
nor U1659 (N_1659,N_1122,N_329);
nand U1660 (N_1660,N_939,N_1190);
or U1661 (N_1661,N_210,N_883);
xor U1662 (N_1662,N_543,N_1044);
xnor U1663 (N_1663,N_1298,N_257);
or U1664 (N_1664,N_1176,N_1180);
or U1665 (N_1665,N_1027,N_1449);
or U1666 (N_1666,N_1160,N_484);
and U1667 (N_1667,N_1021,N_1309);
or U1668 (N_1668,N_1063,N_723);
nand U1669 (N_1669,N_1498,N_1106);
or U1670 (N_1670,N_62,N_1162);
and U1671 (N_1671,N_1188,N_880);
or U1672 (N_1672,N_802,N_1381);
nand U1673 (N_1673,N_598,N_1186);
or U1674 (N_1674,N_323,N_1352);
or U1675 (N_1675,N_297,N_634);
xor U1676 (N_1676,N_1201,N_160);
nand U1677 (N_1677,N_551,N_326);
and U1678 (N_1678,N_1361,N_810);
or U1679 (N_1679,N_669,N_1040);
nor U1680 (N_1680,N_625,N_639);
nor U1681 (N_1681,N_1187,N_602);
and U1682 (N_1682,N_1359,N_248);
xor U1683 (N_1683,N_1306,N_292);
nor U1684 (N_1684,N_503,N_1087);
and U1685 (N_1685,N_1307,N_222);
nor U1686 (N_1686,N_592,N_55);
xor U1687 (N_1687,N_685,N_881);
nand U1688 (N_1688,N_1430,N_301);
or U1689 (N_1689,N_265,N_1238);
and U1690 (N_1690,N_740,N_148);
or U1691 (N_1691,N_356,N_947);
nor U1692 (N_1692,N_868,N_197);
or U1693 (N_1693,N_50,N_1458);
nand U1694 (N_1694,N_1165,N_619);
nor U1695 (N_1695,N_1235,N_332);
nand U1696 (N_1696,N_935,N_189);
nor U1697 (N_1697,N_44,N_1137);
and U1698 (N_1698,N_1248,N_1434);
nand U1699 (N_1699,N_5,N_1061);
or U1700 (N_1700,N_1317,N_679);
nor U1701 (N_1701,N_83,N_1474);
or U1702 (N_1702,N_512,N_378);
and U1703 (N_1703,N_1051,N_682);
nor U1704 (N_1704,N_291,N_866);
and U1705 (N_1705,N_1243,N_788);
nand U1706 (N_1706,N_595,N_839);
and U1707 (N_1707,N_89,N_1066);
xnor U1708 (N_1708,N_218,N_11);
nor U1709 (N_1709,N_121,N_1411);
or U1710 (N_1710,N_1107,N_1178);
nor U1711 (N_1711,N_566,N_369);
xor U1712 (N_1712,N_820,N_701);
nor U1713 (N_1713,N_580,N_905);
xnor U1714 (N_1714,N_1199,N_932);
or U1715 (N_1715,N_590,N_1455);
nand U1716 (N_1716,N_216,N_819);
and U1717 (N_1717,N_427,N_315);
or U1718 (N_1718,N_150,N_413);
or U1719 (N_1719,N_1197,N_1110);
or U1720 (N_1720,N_754,N_473);
or U1721 (N_1721,N_331,N_727);
nor U1722 (N_1722,N_609,N_8);
nor U1723 (N_1723,N_1256,N_848);
and U1724 (N_1724,N_364,N_1315);
nand U1725 (N_1725,N_660,N_1484);
nor U1726 (N_1726,N_958,N_1020);
nor U1727 (N_1727,N_1015,N_154);
and U1728 (N_1728,N_699,N_594);
nor U1729 (N_1729,N_873,N_1446);
nor U1730 (N_1730,N_688,N_203);
and U1731 (N_1731,N_562,N_1183);
or U1732 (N_1732,N_184,N_45);
nand U1733 (N_1733,N_370,N_406);
and U1734 (N_1734,N_649,N_1447);
xnor U1735 (N_1735,N_1299,N_1017);
xor U1736 (N_1736,N_1496,N_613);
nand U1737 (N_1737,N_1468,N_785);
nand U1738 (N_1738,N_1076,N_833);
and U1739 (N_1739,N_1212,N_596);
nand U1740 (N_1740,N_1099,N_1093);
nor U1741 (N_1741,N_690,N_890);
nor U1742 (N_1742,N_344,N_1265);
xor U1743 (N_1743,N_1128,N_597);
nand U1744 (N_1744,N_912,N_1410);
xor U1745 (N_1745,N_896,N_394);
nor U1746 (N_1746,N_1333,N_768);
nand U1747 (N_1747,N_1204,N_1329);
nor U1748 (N_1748,N_242,N_1109);
xnor U1749 (N_1749,N_587,N_799);
and U1750 (N_1750,N_151,N_56);
or U1751 (N_1751,N_172,N_1421);
nand U1752 (N_1752,N_395,N_1346);
nor U1753 (N_1753,N_1177,N_954);
nor U1754 (N_1754,N_1336,N_1143);
nor U1755 (N_1755,N_1431,N_285);
or U1756 (N_1756,N_1237,N_1151);
nand U1757 (N_1757,N_668,N_1192);
or U1758 (N_1758,N_987,N_1085);
and U1759 (N_1759,N_689,N_328);
nor U1760 (N_1760,N_1100,N_761);
nor U1761 (N_1761,N_131,N_996);
and U1762 (N_1762,N_271,N_611);
xor U1763 (N_1763,N_599,N_1438);
nor U1764 (N_1764,N_1002,N_745);
and U1765 (N_1765,N_1478,N_865);
and U1766 (N_1766,N_1184,N_412);
nand U1767 (N_1767,N_174,N_349);
xnor U1768 (N_1768,N_1281,N_282);
nand U1769 (N_1769,N_1016,N_1182);
xnor U1770 (N_1770,N_1089,N_194);
or U1771 (N_1771,N_479,N_1296);
and U1772 (N_1772,N_485,N_714);
nand U1773 (N_1773,N_579,N_650);
or U1774 (N_1774,N_977,N_269);
and U1775 (N_1775,N_900,N_1443);
xor U1776 (N_1776,N_14,N_826);
or U1777 (N_1777,N_389,N_1371);
nor U1778 (N_1778,N_1078,N_537);
nand U1779 (N_1779,N_268,N_357);
xor U1780 (N_1780,N_1139,N_1419);
xnor U1781 (N_1781,N_10,N_147);
nand U1782 (N_1782,N_82,N_535);
and U1783 (N_1783,N_716,N_653);
and U1784 (N_1784,N_632,N_638);
and U1785 (N_1785,N_643,N_1083);
nor U1786 (N_1786,N_79,N_1193);
xnor U1787 (N_1787,N_624,N_509);
nand U1788 (N_1788,N_486,N_1215);
nand U1789 (N_1789,N_464,N_492);
nor U1790 (N_1790,N_1429,N_1292);
and U1791 (N_1791,N_399,N_899);
nand U1792 (N_1792,N_618,N_226);
nand U1793 (N_1793,N_1072,N_1460);
nand U1794 (N_1794,N_845,N_988);
nand U1795 (N_1795,N_29,N_307);
nor U1796 (N_1796,N_532,N_303);
or U1797 (N_1797,N_1487,N_1210);
nand U1798 (N_1798,N_305,N_1175);
xnor U1799 (N_1799,N_556,N_559);
xnor U1800 (N_1800,N_1239,N_1005);
or U1801 (N_1801,N_818,N_1466);
xnor U1802 (N_1802,N_904,N_1145);
and U1803 (N_1803,N_589,N_1316);
nand U1804 (N_1804,N_1043,N_835);
or U1805 (N_1805,N_1038,N_1441);
and U1806 (N_1806,N_629,N_284);
xnor U1807 (N_1807,N_1097,N_872);
nor U1808 (N_1808,N_1037,N_1497);
nor U1809 (N_1809,N_1234,N_1077);
and U1810 (N_1810,N_408,N_1075);
xor U1811 (N_1811,N_95,N_152);
xor U1812 (N_1812,N_909,N_937);
nor U1813 (N_1813,N_340,N_755);
and U1814 (N_1814,N_421,N_1117);
xnor U1815 (N_1815,N_630,N_1283);
and U1816 (N_1816,N_180,N_199);
nand U1817 (N_1817,N_63,N_125);
nor U1818 (N_1818,N_847,N_734);
or U1819 (N_1819,N_110,N_656);
nand U1820 (N_1820,N_973,N_922);
nand U1821 (N_1821,N_520,N_474);
nor U1822 (N_1822,N_612,N_781);
xnor U1823 (N_1823,N_967,N_1354);
xor U1824 (N_1824,N_463,N_75);
or U1825 (N_1825,N_166,N_782);
and U1826 (N_1826,N_568,N_1191);
nand U1827 (N_1827,N_976,N_279);
nand U1828 (N_1828,N_1291,N_952);
xnor U1829 (N_1829,N_141,N_1362);
and U1830 (N_1830,N_453,N_765);
and U1831 (N_1831,N_24,N_806);
or U1832 (N_1832,N_1376,N_1262);
xnor U1833 (N_1833,N_508,N_1456);
nor U1834 (N_1834,N_1463,N_862);
nor U1835 (N_1835,N_250,N_343);
nand U1836 (N_1836,N_239,N_885);
nand U1837 (N_1837,N_771,N_706);
nor U1838 (N_1838,N_665,N_748);
xor U1839 (N_1839,N_829,N_1395);
or U1840 (N_1840,N_876,N_3);
xor U1841 (N_1841,N_127,N_214);
xnor U1842 (N_1842,N_94,N_1217);
nor U1843 (N_1843,N_943,N_1490);
nor U1844 (N_1844,N_1045,N_963);
and U1845 (N_1845,N_1372,N_456);
and U1846 (N_1846,N_533,N_1493);
nor U1847 (N_1847,N_735,N_891);
xnor U1848 (N_1848,N_879,N_1006);
and U1849 (N_1849,N_1130,N_1433);
xor U1850 (N_1850,N_1179,N_805);
or U1851 (N_1851,N_283,N_1115);
xor U1852 (N_1852,N_52,N_698);
nor U1853 (N_1853,N_1278,N_433);
xnor U1854 (N_1854,N_930,N_490);
xnor U1855 (N_1855,N_139,N_1138);
or U1856 (N_1856,N_751,N_1150);
nand U1857 (N_1857,N_824,N_730);
nand U1858 (N_1858,N_767,N_635);
or U1859 (N_1859,N_789,N_762);
nor U1860 (N_1860,N_99,N_968);
or U1861 (N_1861,N_319,N_1049);
nor U1862 (N_1862,N_1196,N_651);
and U1863 (N_1863,N_1437,N_933);
xnor U1864 (N_1864,N_569,N_1331);
nor U1865 (N_1865,N_784,N_1272);
nor U1866 (N_1866,N_1213,N_273);
nor U1867 (N_1867,N_119,N_1088);
nor U1868 (N_1868,N_495,N_49);
nand U1869 (N_1869,N_571,N_1198);
nor U1870 (N_1870,N_386,N_832);
nand U1871 (N_1871,N_1279,N_919);
or U1872 (N_1872,N_352,N_374);
nand U1873 (N_1873,N_261,N_418);
xnor U1874 (N_1874,N_800,N_362);
or U1875 (N_1875,N_1310,N_59);
nand U1876 (N_1876,N_1403,N_377);
nor U1877 (N_1877,N_156,N_975);
and U1878 (N_1878,N_234,N_459);
or U1879 (N_1879,N_640,N_330);
nand U1880 (N_1880,N_102,N_310);
or U1881 (N_1881,N_747,N_274);
or U1882 (N_1882,N_206,N_405);
or U1883 (N_1883,N_1062,N_308);
nand U1884 (N_1884,N_167,N_1407);
nor U1885 (N_1885,N_27,N_376);
nand U1886 (N_1886,N_170,N_1350);
nor U1887 (N_1887,N_204,N_628);
xor U1888 (N_1888,N_1203,N_557);
nor U1889 (N_1889,N_814,N_1082);
xor U1890 (N_1890,N_455,N_1399);
nand U1891 (N_1891,N_1079,N_978);
and U1892 (N_1892,N_294,N_1181);
xnor U1893 (N_1893,N_410,N_614);
xnor U1894 (N_1894,N_1147,N_1377);
nand U1895 (N_1895,N_1289,N_211);
nor U1896 (N_1896,N_1149,N_991);
nor U1897 (N_1897,N_529,N_451);
xor U1898 (N_1898,N_758,N_1118);
or U1899 (N_1899,N_354,N_43);
nand U1900 (N_1900,N_449,N_358);
nor U1901 (N_1901,N_1375,N_1488);
and U1902 (N_1902,N_28,N_48);
nor U1903 (N_1903,N_1277,N_1302);
nor U1904 (N_1904,N_1260,N_715);
nor U1905 (N_1905,N_1258,N_98);
nand U1906 (N_1906,N_34,N_1480);
nor U1907 (N_1907,N_429,N_424);
and U1908 (N_1908,N_722,N_830);
nand U1909 (N_1909,N_572,N_677);
or U1910 (N_1910,N_267,N_443);
or U1911 (N_1911,N_171,N_752);
and U1912 (N_1912,N_1450,N_1436);
or U1913 (N_1913,N_317,N_1048);
and U1914 (N_1914,N_36,N_169);
or U1915 (N_1915,N_1301,N_366);
nand U1916 (N_1916,N_1274,N_205);
xnor U1917 (N_1917,N_663,N_1295);
nor U1918 (N_1918,N_1055,N_322);
and U1919 (N_1919,N_915,N_1428);
nor U1920 (N_1920,N_90,N_917);
nand U1921 (N_1921,N_247,N_739);
xnor U1922 (N_1922,N_1084,N_1422);
nor U1923 (N_1923,N_836,N_276);
xnor U1924 (N_1924,N_380,N_920);
or U1925 (N_1925,N_346,N_130);
nor U1926 (N_1926,N_729,N_661);
nor U1927 (N_1927,N_1068,N_393);
nor U1928 (N_1928,N_372,N_334);
nor U1929 (N_1929,N_1347,N_309);
and U1930 (N_1930,N_867,N_995);
nand U1931 (N_1931,N_938,N_149);
and U1932 (N_1932,N_637,N_1127);
xor U1933 (N_1933,N_1267,N_910);
nand U1934 (N_1934,N_1427,N_908);
xnor U1935 (N_1935,N_155,N_586);
and U1936 (N_1936,N_581,N_465);
nand U1937 (N_1937,N_1152,N_0);
nor U1938 (N_1938,N_365,N_1171);
or U1939 (N_1939,N_1348,N_721);
or U1940 (N_1940,N_831,N_648);
nand U1941 (N_1941,N_1330,N_1311);
nor U1942 (N_1942,N_1358,N_207);
nand U1943 (N_1943,N_1409,N_21);
xnor U1944 (N_1944,N_1349,N_955);
nor U1945 (N_1945,N_957,N_1026);
or U1946 (N_1946,N_187,N_195);
nor U1947 (N_1947,N_858,N_469);
xnor U1948 (N_1948,N_295,N_1001);
nor U1949 (N_1949,N_582,N_1380);
nor U1950 (N_1950,N_897,N_1060);
xnor U1951 (N_1951,N_1251,N_161);
nor U1952 (N_1952,N_929,N_1031);
xnor U1953 (N_1953,N_468,N_480);
nand U1954 (N_1954,N_219,N_560);
nand U1955 (N_1955,N_345,N_350);
xor U1956 (N_1956,N_753,N_1366);
or U1957 (N_1957,N_790,N_1332);
or U1958 (N_1958,N_157,N_849);
xor U1959 (N_1959,N_1297,N_763);
xor U1960 (N_1960,N_1489,N_1244);
and U1961 (N_1961,N_1444,N_591);
nor U1962 (N_1962,N_1360,N_888);
nor U1963 (N_1963,N_1392,N_73);
nor U1964 (N_1964,N_710,N_466);
or U1965 (N_1965,N_46,N_719);
nand U1966 (N_1966,N_23,N_61);
and U1967 (N_1967,N_547,N_986);
xnor U1968 (N_1968,N_652,N_1158);
nand U1969 (N_1969,N_1477,N_641);
nor U1970 (N_1970,N_1194,N_889);
nand U1971 (N_1971,N_1365,N_373);
nor U1972 (N_1972,N_57,N_1050);
or U1973 (N_1973,N_980,N_989);
or U1974 (N_1974,N_511,N_452);
nor U1975 (N_1975,N_892,N_1041);
nand U1976 (N_1976,N_444,N_791);
and U1977 (N_1977,N_318,N_103);
or U1978 (N_1978,N_1308,N_339);
and U1979 (N_1979,N_381,N_1499);
nor U1980 (N_1980,N_115,N_519);
or U1981 (N_1981,N_1282,N_488);
nand U1982 (N_1982,N_1378,N_536);
nand U1983 (N_1983,N_12,N_442);
and U1984 (N_1984,N_972,N_703);
xnor U1985 (N_1985,N_1140,N_4);
nor U1986 (N_1986,N_1413,N_870);
or U1987 (N_1987,N_1033,N_801);
nor U1988 (N_1988,N_118,N_143);
or U1989 (N_1989,N_778,N_1418);
and U1990 (N_1990,N_137,N_223);
and U1991 (N_1991,N_1014,N_776);
nor U1992 (N_1992,N_16,N_1024);
nor U1993 (N_1993,N_1386,N_925);
xor U1994 (N_1994,N_407,N_528);
or U1995 (N_1995,N_450,N_1030);
or U1996 (N_1996,N_821,N_1337);
xor U1997 (N_1997,N_246,N_53);
nand U1998 (N_1998,N_439,N_575);
nor U1999 (N_1999,N_1102,N_263);
nand U2000 (N_2000,N_645,N_430);
or U2001 (N_2001,N_1467,N_1163);
xnor U2002 (N_2002,N_1236,N_1114);
and U2003 (N_2003,N_1313,N_659);
and U2004 (N_2004,N_40,N_1335);
xor U2005 (N_2005,N_803,N_853);
and U2006 (N_2006,N_526,N_538);
and U2007 (N_2007,N_1133,N_146);
or U2008 (N_2008,N_351,N_676);
or U2009 (N_2009,N_725,N_924);
nand U2010 (N_2010,N_181,N_277);
or U2011 (N_2011,N_593,N_1154);
nor U2012 (N_2012,N_527,N_1263);
nand U2013 (N_2013,N_320,N_289);
and U2014 (N_2014,N_913,N_1470);
and U2015 (N_2015,N_258,N_811);
and U2016 (N_2016,N_1426,N_979);
nor U2017 (N_2017,N_383,N_1270);
nor U2018 (N_2018,N_1019,N_949);
and U2019 (N_2019,N_236,N_233);
nor U2020 (N_2020,N_521,N_185);
nand U2021 (N_2021,N_523,N_1424);
and U2022 (N_2022,N_941,N_112);
nor U2023 (N_2023,N_1351,N_1164);
xor U2024 (N_2024,N_434,N_871);
xnor U2025 (N_2025,N_615,N_1095);
or U2026 (N_2026,N_266,N_686);
nor U2027 (N_2027,N_1255,N_1166);
nor U2028 (N_2028,N_502,N_290);
nor U2029 (N_2029,N_546,N_42);
and U2030 (N_2030,N_1457,N_573);
or U2031 (N_2031,N_770,N_228);
xor U2032 (N_2032,N_136,N_101);
xnor U2033 (N_2033,N_1482,N_1073);
xnor U2034 (N_2034,N_1339,N_491);
nor U2035 (N_2035,N_58,N_1326);
and U2036 (N_2036,N_1432,N_1029);
nand U2037 (N_2037,N_39,N_60);
nor U2038 (N_2038,N_1394,N_13);
nand U2039 (N_2039,N_1374,N_1440);
and U2040 (N_2040,N_153,N_335);
xnor U2041 (N_2041,N_1373,N_1284);
nor U2042 (N_2042,N_1170,N_1439);
xor U2043 (N_2043,N_1119,N_221);
or U2044 (N_2044,N_1103,N_1125);
and U2045 (N_2045,N_1207,N_1367);
or U2046 (N_2046,N_1227,N_561);
nor U2047 (N_2047,N_2,N_278);
and U2048 (N_2048,N_1086,N_1471);
nand U2049 (N_2049,N_76,N_1268);
nor U2050 (N_2050,N_1124,N_446);
nand U2051 (N_2051,N_545,N_1363);
nand U2052 (N_2052,N_232,N_544);
or U2053 (N_2053,N_193,N_70);
and U2054 (N_2054,N_983,N_709);
or U2055 (N_2055,N_1092,N_1173);
nand U2056 (N_2056,N_840,N_1035);
nand U2057 (N_2057,N_462,N_1053);
nand U2058 (N_2058,N_1064,N_817);
and U2059 (N_2059,N_804,N_1123);
or U2060 (N_2060,N_982,N_1153);
xor U2061 (N_2061,N_1416,N_774);
xor U2062 (N_2062,N_168,N_432);
xor U2063 (N_2063,N_1384,N_517);
or U2064 (N_2064,N_426,N_1156);
nand U2065 (N_2065,N_506,N_392);
and U2066 (N_2066,N_1069,N_348);
and U2067 (N_2067,N_1003,N_321);
nor U2068 (N_2068,N_994,N_87);
and U2069 (N_2069,N_287,N_245);
xor U2070 (N_2070,N_583,N_176);
or U2071 (N_2071,N_22,N_1218);
nand U2072 (N_2072,N_7,N_368);
xnor U2073 (N_2073,N_603,N_1058);
and U2074 (N_2074,N_518,N_1304);
nand U2075 (N_2075,N_681,N_1144);
xor U2076 (N_2076,N_1475,N_220);
or U2077 (N_2077,N_672,N_841);
and U2078 (N_2078,N_1028,N_960);
and U2079 (N_2079,N_1112,N_647);
or U2080 (N_2080,N_549,N_438);
and U2081 (N_2081,N_173,N_240);
or U2082 (N_2082,N_1328,N_177);
and U2083 (N_2083,N_1325,N_1157);
and U2084 (N_2084,N_93,N_163);
or U2085 (N_2085,N_1141,N_355);
or U2086 (N_2086,N_1293,N_792);
and U2087 (N_2087,N_69,N_1007);
nand U2088 (N_2088,N_425,N_1454);
and U2089 (N_2089,N_808,N_1341);
nor U2090 (N_2090,N_116,N_903);
xnor U2091 (N_2091,N_1189,N_132);
or U2092 (N_2092,N_1257,N_1356);
nand U2093 (N_2093,N_626,N_243);
or U2094 (N_2094,N_743,N_333);
xor U2095 (N_2095,N_961,N_724);
and U2096 (N_2096,N_188,N_304);
xor U2097 (N_2097,N_496,N_726);
and U2098 (N_2098,N_882,N_860);
nor U2099 (N_2099,N_610,N_507);
nor U2100 (N_2100,N_633,N_178);
nand U2101 (N_2101,N_371,N_72);
nor U2102 (N_2102,N_104,N_563);
nor U2103 (N_2103,N_534,N_1408);
nand U2104 (N_2104,N_164,N_68);
and U2105 (N_2105,N_934,N_165);
xor U2106 (N_2106,N_1000,N_1129);
nor U2107 (N_2107,N_481,N_1448);
xor U2108 (N_2108,N_552,N_409);
and U2109 (N_2109,N_705,N_1465);
nand U2110 (N_2110,N_227,N_201);
nor U2111 (N_2111,N_15,N_337);
or U2112 (N_2112,N_1200,N_878);
xnor U2113 (N_2113,N_476,N_1228);
nand U2114 (N_2114,N_694,N_1486);
or U2115 (N_2115,N_704,N_733);
nor U2116 (N_2116,N_1385,N_1303);
xor U2117 (N_2117,N_1401,N_828);
nor U2118 (N_2118,N_85,N_524);
nand U2119 (N_2119,N_926,N_1195);
nand U2120 (N_2120,N_1334,N_20);
nand U2121 (N_2121,N_342,N_436);
or U2122 (N_2122,N_86,N_299);
nand U2123 (N_2123,N_760,N_846);
nor U2124 (N_2124,N_191,N_708);
nand U2125 (N_2125,N_483,N_281);
nand U2126 (N_2126,N_812,N_100);
or U2127 (N_2127,N_875,N_489);
or U2128 (N_2128,N_707,N_542);
and U2129 (N_2129,N_1491,N_499);
and U2130 (N_2130,N_363,N_741);
nor U2131 (N_2131,N_732,N_260);
nand U2132 (N_2132,N_691,N_1230);
nand U2133 (N_2133,N_1116,N_655);
xor U2134 (N_2134,N_1253,N_585);
nor U2135 (N_2135,N_96,N_431);
or U2136 (N_2136,N_843,N_437);
nor U2137 (N_2137,N_577,N_361);
nand U2138 (N_2138,N_850,N_1008);
and U2139 (N_2139,N_695,N_66);
nand U2140 (N_2140,N_530,N_400);
or U2141 (N_2141,N_54,N_764);
and U2142 (N_2142,N_1202,N_1222);
and U2143 (N_2143,N_555,N_460);
xor U2144 (N_2144,N_822,N_1174);
or U2145 (N_2145,N_965,N_1126);
xnor U2146 (N_2146,N_683,N_230);
or U2147 (N_2147,N_280,N_1305);
nand U2148 (N_2148,N_1280,N_1168);
nand U2149 (N_2149,N_718,N_325);
or U2150 (N_2150,N_998,N_921);
xor U2151 (N_2151,N_884,N_88);
xor U2152 (N_2152,N_501,N_584);
xnor U2153 (N_2153,N_241,N_1080);
or U2154 (N_2154,N_1495,N_916);
nor U2155 (N_2155,N_1404,N_84);
xor U2156 (N_2156,N_1009,N_1417);
xnor U2157 (N_2157,N_1070,N_775);
nor U2158 (N_2158,N_179,N_1389);
xor U2159 (N_2159,N_797,N_700);
nand U2160 (N_2160,N_1445,N_852);
or U2161 (N_2161,N_1469,N_646);
xnor U2162 (N_2162,N_298,N_215);
and U2163 (N_2163,N_262,N_1132);
xor U2164 (N_2164,N_1391,N_1368);
or U2165 (N_2165,N_1101,N_898);
or U2166 (N_2166,N_313,N_435);
nand U2167 (N_2167,N_720,N_565);
nor U2168 (N_2168,N_470,N_1318);
or U2169 (N_2169,N_667,N_627);
nor U2170 (N_2170,N_1479,N_494);
nor U2171 (N_2171,N_106,N_256);
nor U2172 (N_2172,N_993,N_422);
xor U2173 (N_2173,N_288,N_382);
or U2174 (N_2174,N_749,N_1211);
xor U2175 (N_2175,N_1405,N_375);
nor U2176 (N_2176,N_454,N_1136);
nand U2177 (N_2177,N_1224,N_931);
xnor U2178 (N_2178,N_175,N_275);
nor U2179 (N_2179,N_738,N_397);
and U2180 (N_2180,N_1451,N_815);
and U2181 (N_2181,N_1004,N_1059);
nand U2182 (N_2182,N_857,N_746);
xor U2183 (N_2183,N_1290,N_779);
nand U2184 (N_2184,N_404,N_1155);
nor U2185 (N_2185,N_254,N_1343);
or U2186 (N_2186,N_642,N_510);
and U2187 (N_2187,N_159,N_1254);
xor U2188 (N_2188,N_1205,N_272);
xnor U2189 (N_2189,N_970,N_644);
nand U2190 (N_2190,N_1185,N_658);
nor U2191 (N_2191,N_1074,N_1324);
and U2192 (N_2192,N_461,N_1252);
and U2193 (N_2193,N_1052,N_945);
or U2194 (N_2194,N_1,N_445);
nand U2195 (N_2195,N_270,N_901);
nor U2196 (N_2196,N_306,N_601);
nand U2197 (N_2197,N_1108,N_1364);
or U2198 (N_2198,N_338,N_255);
or U2199 (N_2199,N_608,N_142);
nand U2200 (N_2200,N_1220,N_249);
or U2201 (N_2201,N_32,N_842);
or U2202 (N_2202,N_756,N_1412);
and U2203 (N_2203,N_91,N_1219);
or U2204 (N_2204,N_448,N_1098);
xnor U2205 (N_2205,N_757,N_74);
nand U2206 (N_2206,N_1320,N_1406);
nand U2207 (N_2207,N_231,N_420);
nand U2208 (N_2208,N_1319,N_126);
nand U2209 (N_2209,N_17,N_576);
or U2210 (N_2210,N_482,N_999);
xor U2211 (N_2211,N_1223,N_780);
and U2212 (N_2212,N_208,N_541);
or U2213 (N_2213,N_664,N_1379);
nand U2214 (N_2214,N_498,N_971);
nor U2215 (N_2215,N_1393,N_423);
and U2216 (N_2216,N_1232,N_1023);
xnor U2217 (N_2217,N_1462,N_525);
nand U2218 (N_2218,N_353,N_574);
xor U2219 (N_2219,N_1388,N_622);
nor U2220 (N_2220,N_616,N_1273);
or U2221 (N_2221,N_390,N_384);
and U2222 (N_2222,N_415,N_1420);
and U2223 (N_2223,N_311,N_359);
and U2224 (N_2224,N_1105,N_1396);
or U2225 (N_2225,N_428,N_108);
or U2226 (N_2226,N_51,N_548);
nor U2227 (N_2227,N_1288,N_680);
xnor U2228 (N_2228,N_918,N_923);
or U2229 (N_2229,N_1091,N_798);
xor U2230 (N_2230,N_558,N_120);
or U2231 (N_2231,N_887,N_825);
and U2232 (N_2232,N_1492,N_140);
nor U2233 (N_2233,N_71,N_515);
or U2234 (N_2234,N_1240,N_144);
xor U2235 (N_2235,N_946,N_869);
nand U2236 (N_2236,N_212,N_673);
and U2237 (N_2237,N_1261,N_621);
nor U2238 (N_2238,N_906,N_1276);
nor U2239 (N_2239,N_314,N_678);
nand U2240 (N_2240,N_1402,N_834);
nor U2241 (N_2241,N_251,N_1271);
xor U2242 (N_2242,N_67,N_759);
or U2243 (N_2243,N_692,N_1344);
and U2244 (N_2244,N_1233,N_505);
xor U2245 (N_2245,N_129,N_213);
or U2246 (N_2246,N_134,N_6);
or U2247 (N_2247,N_974,N_864);
and U2248 (N_2248,N_816,N_37);
and U2249 (N_2249,N_65,N_766);
and U2250 (N_2250,N_1011,N_452);
xor U2251 (N_2251,N_33,N_777);
nand U2252 (N_2252,N_542,N_639);
and U2253 (N_2253,N_699,N_497);
or U2254 (N_2254,N_608,N_1118);
xor U2255 (N_2255,N_1119,N_854);
or U2256 (N_2256,N_550,N_1214);
nor U2257 (N_2257,N_1215,N_444);
nand U2258 (N_2258,N_327,N_856);
or U2259 (N_2259,N_894,N_1435);
and U2260 (N_2260,N_1471,N_1144);
nor U2261 (N_2261,N_923,N_1433);
xor U2262 (N_2262,N_228,N_104);
or U2263 (N_2263,N_683,N_407);
nor U2264 (N_2264,N_1484,N_282);
or U2265 (N_2265,N_936,N_987);
and U2266 (N_2266,N_391,N_1104);
and U2267 (N_2267,N_45,N_1114);
xor U2268 (N_2268,N_76,N_178);
xor U2269 (N_2269,N_1464,N_1262);
xnor U2270 (N_2270,N_1409,N_34);
or U2271 (N_2271,N_1011,N_221);
nand U2272 (N_2272,N_1137,N_1469);
nand U2273 (N_2273,N_1239,N_311);
xnor U2274 (N_2274,N_204,N_1008);
or U2275 (N_2275,N_739,N_1095);
or U2276 (N_2276,N_1349,N_26);
and U2277 (N_2277,N_266,N_1199);
nor U2278 (N_2278,N_691,N_279);
nor U2279 (N_2279,N_739,N_841);
and U2280 (N_2280,N_82,N_201);
and U2281 (N_2281,N_227,N_319);
xnor U2282 (N_2282,N_1409,N_1371);
or U2283 (N_2283,N_218,N_308);
or U2284 (N_2284,N_40,N_1079);
and U2285 (N_2285,N_733,N_0);
or U2286 (N_2286,N_814,N_1087);
nor U2287 (N_2287,N_530,N_202);
and U2288 (N_2288,N_1422,N_161);
xor U2289 (N_2289,N_1417,N_1271);
nor U2290 (N_2290,N_1068,N_558);
xor U2291 (N_2291,N_253,N_645);
or U2292 (N_2292,N_1049,N_63);
or U2293 (N_2293,N_919,N_428);
and U2294 (N_2294,N_1378,N_560);
xnor U2295 (N_2295,N_506,N_1273);
or U2296 (N_2296,N_220,N_145);
xnor U2297 (N_2297,N_219,N_399);
nand U2298 (N_2298,N_523,N_1);
and U2299 (N_2299,N_565,N_898);
nor U2300 (N_2300,N_529,N_904);
or U2301 (N_2301,N_288,N_752);
and U2302 (N_2302,N_323,N_1003);
and U2303 (N_2303,N_937,N_1034);
and U2304 (N_2304,N_994,N_1041);
or U2305 (N_2305,N_890,N_1108);
xnor U2306 (N_2306,N_232,N_438);
nand U2307 (N_2307,N_1038,N_877);
nand U2308 (N_2308,N_760,N_1173);
nor U2309 (N_2309,N_339,N_723);
xnor U2310 (N_2310,N_1079,N_1292);
or U2311 (N_2311,N_517,N_107);
or U2312 (N_2312,N_893,N_614);
nor U2313 (N_2313,N_972,N_682);
or U2314 (N_2314,N_1121,N_1225);
xor U2315 (N_2315,N_311,N_804);
or U2316 (N_2316,N_973,N_564);
nand U2317 (N_2317,N_28,N_1115);
nand U2318 (N_2318,N_1155,N_1408);
and U2319 (N_2319,N_1203,N_272);
xnor U2320 (N_2320,N_1011,N_947);
xor U2321 (N_2321,N_1213,N_160);
nand U2322 (N_2322,N_7,N_1074);
nor U2323 (N_2323,N_1013,N_559);
nor U2324 (N_2324,N_745,N_729);
and U2325 (N_2325,N_73,N_964);
xnor U2326 (N_2326,N_736,N_421);
xor U2327 (N_2327,N_447,N_1099);
and U2328 (N_2328,N_742,N_424);
or U2329 (N_2329,N_618,N_283);
or U2330 (N_2330,N_1251,N_236);
or U2331 (N_2331,N_80,N_1138);
and U2332 (N_2332,N_43,N_421);
nand U2333 (N_2333,N_725,N_329);
nor U2334 (N_2334,N_679,N_866);
or U2335 (N_2335,N_502,N_814);
and U2336 (N_2336,N_1182,N_239);
xor U2337 (N_2337,N_143,N_773);
and U2338 (N_2338,N_299,N_1486);
and U2339 (N_2339,N_547,N_1380);
xor U2340 (N_2340,N_733,N_66);
and U2341 (N_2341,N_1228,N_976);
xnor U2342 (N_2342,N_1405,N_82);
and U2343 (N_2343,N_107,N_114);
or U2344 (N_2344,N_927,N_1489);
or U2345 (N_2345,N_977,N_1409);
or U2346 (N_2346,N_561,N_1373);
xor U2347 (N_2347,N_1079,N_381);
nand U2348 (N_2348,N_148,N_58);
and U2349 (N_2349,N_1182,N_370);
nor U2350 (N_2350,N_292,N_294);
nor U2351 (N_2351,N_542,N_1299);
nor U2352 (N_2352,N_748,N_863);
xor U2353 (N_2353,N_400,N_68);
or U2354 (N_2354,N_417,N_1340);
nand U2355 (N_2355,N_578,N_598);
and U2356 (N_2356,N_230,N_722);
and U2357 (N_2357,N_968,N_418);
nor U2358 (N_2358,N_280,N_348);
nor U2359 (N_2359,N_1408,N_1097);
nor U2360 (N_2360,N_43,N_905);
and U2361 (N_2361,N_943,N_475);
xnor U2362 (N_2362,N_106,N_1217);
nor U2363 (N_2363,N_237,N_961);
nand U2364 (N_2364,N_1298,N_858);
xor U2365 (N_2365,N_722,N_550);
and U2366 (N_2366,N_794,N_592);
nand U2367 (N_2367,N_1047,N_1359);
and U2368 (N_2368,N_1408,N_1152);
and U2369 (N_2369,N_1009,N_1353);
and U2370 (N_2370,N_551,N_913);
and U2371 (N_2371,N_1122,N_385);
xor U2372 (N_2372,N_739,N_499);
xnor U2373 (N_2373,N_830,N_597);
and U2374 (N_2374,N_903,N_281);
and U2375 (N_2375,N_345,N_1239);
nor U2376 (N_2376,N_565,N_735);
and U2377 (N_2377,N_701,N_139);
and U2378 (N_2378,N_927,N_670);
or U2379 (N_2379,N_768,N_414);
nor U2380 (N_2380,N_1358,N_664);
nand U2381 (N_2381,N_88,N_534);
or U2382 (N_2382,N_173,N_312);
xnor U2383 (N_2383,N_1403,N_247);
and U2384 (N_2384,N_1269,N_994);
nand U2385 (N_2385,N_358,N_105);
nand U2386 (N_2386,N_1365,N_937);
xnor U2387 (N_2387,N_250,N_430);
nand U2388 (N_2388,N_75,N_668);
or U2389 (N_2389,N_1088,N_1389);
nand U2390 (N_2390,N_1397,N_12);
nand U2391 (N_2391,N_212,N_857);
or U2392 (N_2392,N_845,N_1024);
nor U2393 (N_2393,N_979,N_1427);
or U2394 (N_2394,N_1033,N_497);
and U2395 (N_2395,N_136,N_1402);
nand U2396 (N_2396,N_76,N_1058);
and U2397 (N_2397,N_1230,N_393);
nor U2398 (N_2398,N_896,N_493);
nand U2399 (N_2399,N_179,N_827);
nand U2400 (N_2400,N_904,N_443);
xor U2401 (N_2401,N_1321,N_769);
xor U2402 (N_2402,N_1379,N_722);
xnor U2403 (N_2403,N_594,N_898);
or U2404 (N_2404,N_599,N_839);
nor U2405 (N_2405,N_776,N_579);
nand U2406 (N_2406,N_98,N_723);
and U2407 (N_2407,N_1438,N_425);
nor U2408 (N_2408,N_1425,N_1135);
xor U2409 (N_2409,N_27,N_1374);
nor U2410 (N_2410,N_839,N_1203);
or U2411 (N_2411,N_1136,N_146);
nor U2412 (N_2412,N_310,N_1218);
xnor U2413 (N_2413,N_494,N_575);
nor U2414 (N_2414,N_1433,N_492);
nor U2415 (N_2415,N_107,N_995);
xnor U2416 (N_2416,N_1088,N_220);
xnor U2417 (N_2417,N_1277,N_305);
xnor U2418 (N_2418,N_419,N_543);
nand U2419 (N_2419,N_1359,N_747);
nor U2420 (N_2420,N_407,N_12);
and U2421 (N_2421,N_336,N_1494);
and U2422 (N_2422,N_1296,N_5);
and U2423 (N_2423,N_1328,N_132);
nand U2424 (N_2424,N_1362,N_980);
nor U2425 (N_2425,N_650,N_255);
or U2426 (N_2426,N_414,N_984);
and U2427 (N_2427,N_234,N_404);
or U2428 (N_2428,N_1463,N_301);
xnor U2429 (N_2429,N_1387,N_1264);
or U2430 (N_2430,N_309,N_0);
nand U2431 (N_2431,N_878,N_36);
xor U2432 (N_2432,N_1032,N_94);
nand U2433 (N_2433,N_1395,N_361);
xor U2434 (N_2434,N_659,N_119);
and U2435 (N_2435,N_1225,N_713);
nor U2436 (N_2436,N_332,N_571);
nor U2437 (N_2437,N_459,N_392);
and U2438 (N_2438,N_247,N_991);
nand U2439 (N_2439,N_294,N_1242);
and U2440 (N_2440,N_1295,N_968);
nor U2441 (N_2441,N_611,N_177);
xor U2442 (N_2442,N_660,N_208);
and U2443 (N_2443,N_1121,N_1174);
and U2444 (N_2444,N_1100,N_251);
nor U2445 (N_2445,N_1144,N_197);
and U2446 (N_2446,N_482,N_1219);
nand U2447 (N_2447,N_361,N_53);
or U2448 (N_2448,N_935,N_153);
xor U2449 (N_2449,N_612,N_1167);
nand U2450 (N_2450,N_1220,N_224);
nand U2451 (N_2451,N_134,N_435);
or U2452 (N_2452,N_1216,N_1315);
nor U2453 (N_2453,N_60,N_746);
or U2454 (N_2454,N_651,N_1415);
xnor U2455 (N_2455,N_783,N_1386);
nand U2456 (N_2456,N_91,N_973);
or U2457 (N_2457,N_96,N_389);
and U2458 (N_2458,N_1407,N_159);
nor U2459 (N_2459,N_1165,N_1016);
or U2460 (N_2460,N_111,N_581);
xor U2461 (N_2461,N_105,N_1397);
xnor U2462 (N_2462,N_286,N_6);
nor U2463 (N_2463,N_855,N_747);
nand U2464 (N_2464,N_277,N_982);
and U2465 (N_2465,N_1222,N_337);
and U2466 (N_2466,N_1320,N_287);
nand U2467 (N_2467,N_1304,N_476);
and U2468 (N_2468,N_115,N_1480);
or U2469 (N_2469,N_393,N_520);
nor U2470 (N_2470,N_1360,N_324);
nand U2471 (N_2471,N_1118,N_1026);
xor U2472 (N_2472,N_1487,N_114);
xnor U2473 (N_2473,N_1220,N_424);
nor U2474 (N_2474,N_1394,N_423);
nand U2475 (N_2475,N_127,N_1197);
nand U2476 (N_2476,N_721,N_639);
nand U2477 (N_2477,N_284,N_995);
xnor U2478 (N_2478,N_903,N_663);
or U2479 (N_2479,N_395,N_735);
or U2480 (N_2480,N_1381,N_861);
nand U2481 (N_2481,N_397,N_744);
nor U2482 (N_2482,N_103,N_737);
or U2483 (N_2483,N_1042,N_795);
and U2484 (N_2484,N_836,N_121);
or U2485 (N_2485,N_160,N_100);
nor U2486 (N_2486,N_745,N_433);
and U2487 (N_2487,N_1466,N_592);
nand U2488 (N_2488,N_428,N_1171);
and U2489 (N_2489,N_605,N_62);
and U2490 (N_2490,N_1399,N_1196);
or U2491 (N_2491,N_791,N_522);
xor U2492 (N_2492,N_1076,N_519);
and U2493 (N_2493,N_14,N_1);
nand U2494 (N_2494,N_654,N_919);
nand U2495 (N_2495,N_1148,N_915);
or U2496 (N_2496,N_1298,N_1439);
xnor U2497 (N_2497,N_105,N_1394);
or U2498 (N_2498,N_946,N_546);
or U2499 (N_2499,N_278,N_339);
nand U2500 (N_2500,N_1047,N_1068);
nand U2501 (N_2501,N_694,N_478);
nand U2502 (N_2502,N_1064,N_177);
nor U2503 (N_2503,N_1281,N_1330);
and U2504 (N_2504,N_817,N_1068);
nor U2505 (N_2505,N_464,N_396);
xnor U2506 (N_2506,N_560,N_13);
nor U2507 (N_2507,N_274,N_527);
and U2508 (N_2508,N_1279,N_366);
and U2509 (N_2509,N_279,N_655);
nor U2510 (N_2510,N_814,N_923);
and U2511 (N_2511,N_883,N_667);
xor U2512 (N_2512,N_858,N_503);
xnor U2513 (N_2513,N_177,N_78);
or U2514 (N_2514,N_742,N_1347);
nor U2515 (N_2515,N_249,N_794);
or U2516 (N_2516,N_1394,N_1031);
xor U2517 (N_2517,N_539,N_243);
nor U2518 (N_2518,N_995,N_568);
nor U2519 (N_2519,N_1201,N_1210);
xor U2520 (N_2520,N_363,N_1130);
nand U2521 (N_2521,N_278,N_1048);
nand U2522 (N_2522,N_744,N_1110);
nor U2523 (N_2523,N_176,N_1267);
nor U2524 (N_2524,N_30,N_719);
xnor U2525 (N_2525,N_717,N_246);
nor U2526 (N_2526,N_950,N_937);
or U2527 (N_2527,N_599,N_751);
and U2528 (N_2528,N_1138,N_1098);
or U2529 (N_2529,N_399,N_208);
nand U2530 (N_2530,N_1201,N_1144);
xor U2531 (N_2531,N_1334,N_1138);
or U2532 (N_2532,N_1102,N_3);
nand U2533 (N_2533,N_1312,N_1268);
nor U2534 (N_2534,N_1051,N_62);
xnor U2535 (N_2535,N_76,N_262);
and U2536 (N_2536,N_1005,N_669);
nor U2537 (N_2537,N_1331,N_379);
nor U2538 (N_2538,N_872,N_514);
or U2539 (N_2539,N_809,N_297);
xnor U2540 (N_2540,N_515,N_1497);
xor U2541 (N_2541,N_1001,N_418);
nor U2542 (N_2542,N_546,N_821);
and U2543 (N_2543,N_412,N_804);
nand U2544 (N_2544,N_1257,N_1111);
or U2545 (N_2545,N_675,N_1321);
and U2546 (N_2546,N_1364,N_1442);
or U2547 (N_2547,N_1057,N_316);
and U2548 (N_2548,N_1297,N_320);
nand U2549 (N_2549,N_509,N_1295);
or U2550 (N_2550,N_653,N_1153);
nor U2551 (N_2551,N_1392,N_1038);
nor U2552 (N_2552,N_900,N_779);
and U2553 (N_2553,N_440,N_444);
xor U2554 (N_2554,N_1149,N_1375);
nor U2555 (N_2555,N_1312,N_475);
or U2556 (N_2556,N_911,N_1033);
nand U2557 (N_2557,N_1478,N_1464);
nor U2558 (N_2558,N_660,N_474);
nor U2559 (N_2559,N_1124,N_660);
or U2560 (N_2560,N_575,N_875);
nand U2561 (N_2561,N_287,N_963);
nor U2562 (N_2562,N_1058,N_1032);
nand U2563 (N_2563,N_73,N_574);
or U2564 (N_2564,N_497,N_86);
and U2565 (N_2565,N_1444,N_57);
and U2566 (N_2566,N_383,N_894);
and U2567 (N_2567,N_125,N_1450);
nor U2568 (N_2568,N_1443,N_579);
or U2569 (N_2569,N_454,N_1430);
nand U2570 (N_2570,N_610,N_1144);
xnor U2571 (N_2571,N_612,N_619);
nand U2572 (N_2572,N_83,N_1242);
nand U2573 (N_2573,N_1380,N_1045);
or U2574 (N_2574,N_401,N_1338);
xnor U2575 (N_2575,N_659,N_210);
xnor U2576 (N_2576,N_1408,N_1374);
or U2577 (N_2577,N_174,N_337);
or U2578 (N_2578,N_988,N_749);
or U2579 (N_2579,N_1153,N_473);
nor U2580 (N_2580,N_39,N_616);
xor U2581 (N_2581,N_1089,N_1435);
nor U2582 (N_2582,N_971,N_825);
xor U2583 (N_2583,N_1469,N_1460);
nand U2584 (N_2584,N_657,N_416);
nand U2585 (N_2585,N_115,N_808);
nand U2586 (N_2586,N_141,N_310);
or U2587 (N_2587,N_144,N_71);
and U2588 (N_2588,N_1009,N_689);
or U2589 (N_2589,N_700,N_1480);
nor U2590 (N_2590,N_980,N_1090);
nor U2591 (N_2591,N_1183,N_601);
xor U2592 (N_2592,N_1261,N_702);
xnor U2593 (N_2593,N_250,N_764);
or U2594 (N_2594,N_395,N_24);
xor U2595 (N_2595,N_934,N_1181);
nand U2596 (N_2596,N_576,N_516);
nand U2597 (N_2597,N_1283,N_1008);
or U2598 (N_2598,N_937,N_151);
xor U2599 (N_2599,N_1091,N_1136);
or U2600 (N_2600,N_638,N_1109);
and U2601 (N_2601,N_805,N_1427);
nor U2602 (N_2602,N_554,N_1354);
nor U2603 (N_2603,N_1435,N_738);
or U2604 (N_2604,N_853,N_1135);
nor U2605 (N_2605,N_957,N_1008);
and U2606 (N_2606,N_303,N_203);
nand U2607 (N_2607,N_825,N_54);
and U2608 (N_2608,N_161,N_1107);
or U2609 (N_2609,N_1213,N_392);
and U2610 (N_2610,N_76,N_578);
nor U2611 (N_2611,N_1121,N_104);
nand U2612 (N_2612,N_121,N_1346);
and U2613 (N_2613,N_1053,N_243);
and U2614 (N_2614,N_473,N_96);
nand U2615 (N_2615,N_919,N_703);
and U2616 (N_2616,N_995,N_106);
or U2617 (N_2617,N_1126,N_395);
and U2618 (N_2618,N_972,N_969);
and U2619 (N_2619,N_342,N_1132);
nor U2620 (N_2620,N_528,N_1084);
and U2621 (N_2621,N_928,N_537);
or U2622 (N_2622,N_939,N_1350);
or U2623 (N_2623,N_1316,N_358);
xor U2624 (N_2624,N_433,N_617);
nor U2625 (N_2625,N_1463,N_567);
nor U2626 (N_2626,N_991,N_1471);
xor U2627 (N_2627,N_311,N_481);
and U2628 (N_2628,N_1164,N_401);
nand U2629 (N_2629,N_847,N_195);
and U2630 (N_2630,N_274,N_273);
and U2631 (N_2631,N_870,N_809);
xnor U2632 (N_2632,N_343,N_1374);
nor U2633 (N_2633,N_607,N_306);
and U2634 (N_2634,N_1119,N_663);
or U2635 (N_2635,N_842,N_803);
nand U2636 (N_2636,N_837,N_209);
xor U2637 (N_2637,N_1442,N_1340);
nand U2638 (N_2638,N_763,N_1048);
xor U2639 (N_2639,N_651,N_919);
nand U2640 (N_2640,N_846,N_1113);
nand U2641 (N_2641,N_1100,N_335);
or U2642 (N_2642,N_1041,N_210);
xor U2643 (N_2643,N_584,N_1035);
xnor U2644 (N_2644,N_568,N_1280);
nor U2645 (N_2645,N_1427,N_400);
xor U2646 (N_2646,N_620,N_929);
and U2647 (N_2647,N_466,N_665);
nor U2648 (N_2648,N_234,N_1422);
xnor U2649 (N_2649,N_1186,N_1083);
xor U2650 (N_2650,N_1032,N_524);
xor U2651 (N_2651,N_1028,N_858);
and U2652 (N_2652,N_627,N_307);
nor U2653 (N_2653,N_1462,N_1032);
and U2654 (N_2654,N_1445,N_1489);
nand U2655 (N_2655,N_262,N_1435);
nand U2656 (N_2656,N_796,N_1313);
xor U2657 (N_2657,N_195,N_1098);
and U2658 (N_2658,N_551,N_1065);
xnor U2659 (N_2659,N_76,N_1422);
nand U2660 (N_2660,N_920,N_255);
nand U2661 (N_2661,N_451,N_754);
nand U2662 (N_2662,N_967,N_1190);
nor U2663 (N_2663,N_1340,N_1316);
nor U2664 (N_2664,N_1350,N_196);
xor U2665 (N_2665,N_1258,N_573);
nor U2666 (N_2666,N_193,N_673);
and U2667 (N_2667,N_292,N_185);
nand U2668 (N_2668,N_1009,N_1179);
nand U2669 (N_2669,N_403,N_347);
xor U2670 (N_2670,N_1350,N_1206);
xor U2671 (N_2671,N_968,N_337);
and U2672 (N_2672,N_38,N_745);
xor U2673 (N_2673,N_532,N_1462);
and U2674 (N_2674,N_392,N_763);
nor U2675 (N_2675,N_1127,N_1081);
nand U2676 (N_2676,N_675,N_930);
or U2677 (N_2677,N_1161,N_1347);
or U2678 (N_2678,N_1188,N_354);
and U2679 (N_2679,N_937,N_471);
xnor U2680 (N_2680,N_735,N_1448);
or U2681 (N_2681,N_417,N_429);
and U2682 (N_2682,N_358,N_93);
nor U2683 (N_2683,N_996,N_368);
and U2684 (N_2684,N_1055,N_709);
nand U2685 (N_2685,N_1022,N_926);
xnor U2686 (N_2686,N_974,N_1038);
xor U2687 (N_2687,N_246,N_306);
nand U2688 (N_2688,N_1486,N_759);
nor U2689 (N_2689,N_1324,N_548);
xor U2690 (N_2690,N_467,N_1434);
and U2691 (N_2691,N_201,N_433);
xor U2692 (N_2692,N_69,N_35);
nand U2693 (N_2693,N_702,N_826);
nor U2694 (N_2694,N_904,N_194);
and U2695 (N_2695,N_300,N_935);
and U2696 (N_2696,N_1186,N_1151);
nor U2697 (N_2697,N_1310,N_318);
or U2698 (N_2698,N_19,N_640);
nand U2699 (N_2699,N_1445,N_1108);
nand U2700 (N_2700,N_599,N_931);
xnor U2701 (N_2701,N_1251,N_1235);
nand U2702 (N_2702,N_315,N_1032);
nor U2703 (N_2703,N_388,N_358);
and U2704 (N_2704,N_946,N_1467);
xor U2705 (N_2705,N_1009,N_389);
nor U2706 (N_2706,N_1039,N_84);
nor U2707 (N_2707,N_907,N_483);
and U2708 (N_2708,N_1430,N_256);
nor U2709 (N_2709,N_51,N_703);
xor U2710 (N_2710,N_526,N_1282);
xor U2711 (N_2711,N_63,N_1483);
nand U2712 (N_2712,N_1208,N_121);
nor U2713 (N_2713,N_1402,N_218);
and U2714 (N_2714,N_699,N_1273);
nand U2715 (N_2715,N_66,N_1465);
nand U2716 (N_2716,N_384,N_560);
and U2717 (N_2717,N_1338,N_984);
or U2718 (N_2718,N_293,N_1248);
or U2719 (N_2719,N_93,N_201);
nand U2720 (N_2720,N_46,N_173);
xor U2721 (N_2721,N_1159,N_710);
xor U2722 (N_2722,N_345,N_872);
and U2723 (N_2723,N_916,N_991);
xor U2724 (N_2724,N_308,N_765);
nor U2725 (N_2725,N_6,N_551);
and U2726 (N_2726,N_590,N_1312);
nand U2727 (N_2727,N_694,N_523);
xnor U2728 (N_2728,N_682,N_172);
nand U2729 (N_2729,N_317,N_866);
nand U2730 (N_2730,N_466,N_1210);
or U2731 (N_2731,N_101,N_886);
or U2732 (N_2732,N_383,N_208);
nand U2733 (N_2733,N_201,N_551);
nand U2734 (N_2734,N_168,N_343);
nor U2735 (N_2735,N_762,N_65);
or U2736 (N_2736,N_700,N_513);
nor U2737 (N_2737,N_922,N_341);
xor U2738 (N_2738,N_509,N_1189);
and U2739 (N_2739,N_600,N_80);
or U2740 (N_2740,N_562,N_1339);
and U2741 (N_2741,N_1171,N_431);
nor U2742 (N_2742,N_760,N_1014);
and U2743 (N_2743,N_364,N_510);
xnor U2744 (N_2744,N_1028,N_406);
or U2745 (N_2745,N_1420,N_80);
nor U2746 (N_2746,N_1352,N_1214);
nor U2747 (N_2747,N_126,N_1218);
xor U2748 (N_2748,N_444,N_1180);
nor U2749 (N_2749,N_68,N_794);
nand U2750 (N_2750,N_1208,N_730);
nand U2751 (N_2751,N_137,N_658);
xnor U2752 (N_2752,N_94,N_148);
xor U2753 (N_2753,N_859,N_1036);
or U2754 (N_2754,N_838,N_1105);
or U2755 (N_2755,N_1471,N_314);
nand U2756 (N_2756,N_1452,N_752);
and U2757 (N_2757,N_1278,N_1143);
and U2758 (N_2758,N_1258,N_1044);
nor U2759 (N_2759,N_788,N_1112);
nor U2760 (N_2760,N_902,N_622);
and U2761 (N_2761,N_256,N_504);
and U2762 (N_2762,N_1181,N_8);
nand U2763 (N_2763,N_299,N_933);
or U2764 (N_2764,N_50,N_1422);
and U2765 (N_2765,N_690,N_1189);
and U2766 (N_2766,N_345,N_129);
nand U2767 (N_2767,N_42,N_1067);
nand U2768 (N_2768,N_169,N_94);
nor U2769 (N_2769,N_1498,N_1126);
or U2770 (N_2770,N_274,N_811);
and U2771 (N_2771,N_1141,N_1083);
nand U2772 (N_2772,N_727,N_1180);
xor U2773 (N_2773,N_1288,N_159);
or U2774 (N_2774,N_1425,N_578);
xor U2775 (N_2775,N_724,N_932);
and U2776 (N_2776,N_555,N_497);
xor U2777 (N_2777,N_350,N_844);
nor U2778 (N_2778,N_756,N_1396);
nor U2779 (N_2779,N_501,N_875);
nor U2780 (N_2780,N_128,N_660);
and U2781 (N_2781,N_115,N_375);
and U2782 (N_2782,N_765,N_442);
or U2783 (N_2783,N_940,N_705);
xnor U2784 (N_2784,N_1314,N_481);
nand U2785 (N_2785,N_1043,N_14);
or U2786 (N_2786,N_117,N_61);
xor U2787 (N_2787,N_1370,N_1339);
or U2788 (N_2788,N_487,N_1);
and U2789 (N_2789,N_986,N_502);
or U2790 (N_2790,N_1007,N_194);
xor U2791 (N_2791,N_534,N_859);
and U2792 (N_2792,N_589,N_870);
xor U2793 (N_2793,N_674,N_1223);
nand U2794 (N_2794,N_294,N_1076);
or U2795 (N_2795,N_440,N_822);
and U2796 (N_2796,N_1253,N_1310);
xnor U2797 (N_2797,N_354,N_170);
nor U2798 (N_2798,N_306,N_236);
and U2799 (N_2799,N_1154,N_1250);
nand U2800 (N_2800,N_1383,N_216);
xnor U2801 (N_2801,N_1019,N_123);
nor U2802 (N_2802,N_1236,N_1242);
nand U2803 (N_2803,N_1350,N_319);
xnor U2804 (N_2804,N_1381,N_416);
nand U2805 (N_2805,N_856,N_1374);
xor U2806 (N_2806,N_805,N_801);
or U2807 (N_2807,N_381,N_345);
and U2808 (N_2808,N_268,N_606);
and U2809 (N_2809,N_1293,N_1029);
or U2810 (N_2810,N_762,N_1109);
nor U2811 (N_2811,N_695,N_846);
xor U2812 (N_2812,N_628,N_733);
nand U2813 (N_2813,N_842,N_1490);
or U2814 (N_2814,N_1104,N_1119);
nor U2815 (N_2815,N_568,N_498);
nor U2816 (N_2816,N_262,N_505);
nor U2817 (N_2817,N_1276,N_802);
xor U2818 (N_2818,N_1116,N_116);
nand U2819 (N_2819,N_315,N_735);
and U2820 (N_2820,N_732,N_1442);
nand U2821 (N_2821,N_237,N_139);
nor U2822 (N_2822,N_612,N_1366);
or U2823 (N_2823,N_140,N_334);
nand U2824 (N_2824,N_1145,N_528);
xnor U2825 (N_2825,N_1165,N_1192);
or U2826 (N_2826,N_815,N_585);
xnor U2827 (N_2827,N_317,N_995);
nor U2828 (N_2828,N_1053,N_1050);
xor U2829 (N_2829,N_1277,N_1209);
xnor U2830 (N_2830,N_875,N_901);
or U2831 (N_2831,N_282,N_1231);
xnor U2832 (N_2832,N_377,N_168);
or U2833 (N_2833,N_1314,N_1275);
and U2834 (N_2834,N_719,N_470);
nor U2835 (N_2835,N_1376,N_866);
nor U2836 (N_2836,N_847,N_743);
and U2837 (N_2837,N_230,N_894);
xor U2838 (N_2838,N_340,N_1130);
and U2839 (N_2839,N_1479,N_623);
nand U2840 (N_2840,N_647,N_941);
and U2841 (N_2841,N_1357,N_1347);
nand U2842 (N_2842,N_70,N_1467);
and U2843 (N_2843,N_1019,N_618);
nand U2844 (N_2844,N_1084,N_1236);
xor U2845 (N_2845,N_591,N_498);
or U2846 (N_2846,N_412,N_1352);
xor U2847 (N_2847,N_1009,N_1379);
nor U2848 (N_2848,N_775,N_472);
or U2849 (N_2849,N_387,N_869);
nor U2850 (N_2850,N_1105,N_658);
and U2851 (N_2851,N_681,N_503);
and U2852 (N_2852,N_131,N_603);
or U2853 (N_2853,N_1107,N_1223);
xor U2854 (N_2854,N_740,N_933);
and U2855 (N_2855,N_1184,N_597);
or U2856 (N_2856,N_965,N_486);
nand U2857 (N_2857,N_1211,N_1114);
nand U2858 (N_2858,N_376,N_71);
and U2859 (N_2859,N_138,N_738);
and U2860 (N_2860,N_826,N_1205);
xnor U2861 (N_2861,N_1146,N_893);
nor U2862 (N_2862,N_1401,N_108);
nand U2863 (N_2863,N_1048,N_965);
nor U2864 (N_2864,N_1278,N_33);
or U2865 (N_2865,N_662,N_885);
nand U2866 (N_2866,N_648,N_647);
or U2867 (N_2867,N_83,N_1416);
nor U2868 (N_2868,N_1479,N_424);
xnor U2869 (N_2869,N_512,N_436);
nor U2870 (N_2870,N_470,N_0);
or U2871 (N_2871,N_725,N_1371);
nor U2872 (N_2872,N_451,N_161);
nor U2873 (N_2873,N_1213,N_1107);
or U2874 (N_2874,N_963,N_807);
xnor U2875 (N_2875,N_1437,N_72);
nor U2876 (N_2876,N_719,N_523);
xor U2877 (N_2877,N_655,N_60);
or U2878 (N_2878,N_561,N_223);
and U2879 (N_2879,N_815,N_147);
nand U2880 (N_2880,N_1278,N_959);
and U2881 (N_2881,N_1223,N_836);
or U2882 (N_2882,N_1244,N_1142);
xor U2883 (N_2883,N_670,N_791);
or U2884 (N_2884,N_1375,N_1324);
nand U2885 (N_2885,N_880,N_974);
nand U2886 (N_2886,N_1387,N_115);
and U2887 (N_2887,N_1469,N_1248);
or U2888 (N_2888,N_588,N_1367);
or U2889 (N_2889,N_854,N_1257);
nor U2890 (N_2890,N_225,N_833);
or U2891 (N_2891,N_737,N_266);
or U2892 (N_2892,N_186,N_909);
nand U2893 (N_2893,N_120,N_1149);
xnor U2894 (N_2894,N_220,N_252);
nor U2895 (N_2895,N_834,N_1336);
nor U2896 (N_2896,N_698,N_1486);
nor U2897 (N_2897,N_679,N_410);
and U2898 (N_2898,N_1434,N_1010);
xor U2899 (N_2899,N_1429,N_564);
and U2900 (N_2900,N_78,N_1295);
nor U2901 (N_2901,N_1090,N_505);
and U2902 (N_2902,N_375,N_40);
or U2903 (N_2903,N_1323,N_887);
and U2904 (N_2904,N_877,N_964);
xor U2905 (N_2905,N_1221,N_754);
nor U2906 (N_2906,N_358,N_269);
and U2907 (N_2907,N_504,N_523);
xnor U2908 (N_2908,N_972,N_921);
and U2909 (N_2909,N_155,N_1089);
or U2910 (N_2910,N_1174,N_1427);
and U2911 (N_2911,N_1380,N_588);
xor U2912 (N_2912,N_1389,N_376);
nor U2913 (N_2913,N_654,N_541);
nor U2914 (N_2914,N_350,N_1112);
nand U2915 (N_2915,N_1395,N_1301);
and U2916 (N_2916,N_664,N_808);
xor U2917 (N_2917,N_346,N_409);
xor U2918 (N_2918,N_174,N_82);
xnor U2919 (N_2919,N_932,N_722);
and U2920 (N_2920,N_1160,N_251);
and U2921 (N_2921,N_1092,N_864);
and U2922 (N_2922,N_989,N_1406);
nor U2923 (N_2923,N_818,N_474);
xnor U2924 (N_2924,N_1064,N_875);
nor U2925 (N_2925,N_718,N_686);
nor U2926 (N_2926,N_1243,N_474);
nor U2927 (N_2927,N_436,N_917);
and U2928 (N_2928,N_1174,N_257);
nand U2929 (N_2929,N_887,N_1026);
xnor U2930 (N_2930,N_1401,N_1274);
and U2931 (N_2931,N_607,N_654);
nor U2932 (N_2932,N_1340,N_1407);
xnor U2933 (N_2933,N_290,N_65);
xor U2934 (N_2934,N_1239,N_1257);
or U2935 (N_2935,N_210,N_304);
xnor U2936 (N_2936,N_1310,N_590);
nand U2937 (N_2937,N_1305,N_730);
nand U2938 (N_2938,N_161,N_1090);
xor U2939 (N_2939,N_1399,N_1055);
xor U2940 (N_2940,N_802,N_839);
nor U2941 (N_2941,N_1286,N_590);
nand U2942 (N_2942,N_824,N_1313);
and U2943 (N_2943,N_843,N_139);
and U2944 (N_2944,N_611,N_408);
and U2945 (N_2945,N_445,N_1252);
nand U2946 (N_2946,N_651,N_1137);
or U2947 (N_2947,N_566,N_27);
nor U2948 (N_2948,N_961,N_1278);
nand U2949 (N_2949,N_1434,N_789);
or U2950 (N_2950,N_1063,N_153);
and U2951 (N_2951,N_192,N_114);
nor U2952 (N_2952,N_263,N_248);
nor U2953 (N_2953,N_664,N_30);
xor U2954 (N_2954,N_687,N_1270);
nand U2955 (N_2955,N_803,N_148);
xnor U2956 (N_2956,N_1267,N_486);
nand U2957 (N_2957,N_1371,N_1320);
xnor U2958 (N_2958,N_765,N_334);
and U2959 (N_2959,N_1056,N_1262);
nand U2960 (N_2960,N_874,N_672);
or U2961 (N_2961,N_606,N_970);
or U2962 (N_2962,N_971,N_454);
and U2963 (N_2963,N_359,N_1082);
nor U2964 (N_2964,N_1208,N_157);
or U2965 (N_2965,N_62,N_1362);
nor U2966 (N_2966,N_966,N_542);
or U2967 (N_2967,N_530,N_94);
nor U2968 (N_2968,N_897,N_119);
or U2969 (N_2969,N_1226,N_421);
and U2970 (N_2970,N_507,N_231);
nor U2971 (N_2971,N_779,N_509);
or U2972 (N_2972,N_113,N_590);
and U2973 (N_2973,N_559,N_533);
xnor U2974 (N_2974,N_546,N_1344);
nor U2975 (N_2975,N_576,N_1417);
nor U2976 (N_2976,N_697,N_719);
nor U2977 (N_2977,N_561,N_178);
nand U2978 (N_2978,N_267,N_1164);
or U2979 (N_2979,N_809,N_840);
nor U2980 (N_2980,N_311,N_1324);
nand U2981 (N_2981,N_204,N_789);
and U2982 (N_2982,N_197,N_1233);
nand U2983 (N_2983,N_964,N_451);
nor U2984 (N_2984,N_80,N_1221);
or U2985 (N_2985,N_1417,N_802);
nor U2986 (N_2986,N_823,N_46);
nor U2987 (N_2987,N_101,N_434);
nor U2988 (N_2988,N_1248,N_252);
or U2989 (N_2989,N_626,N_1084);
or U2990 (N_2990,N_346,N_304);
nor U2991 (N_2991,N_947,N_281);
or U2992 (N_2992,N_263,N_284);
xnor U2993 (N_2993,N_1191,N_61);
and U2994 (N_2994,N_1488,N_823);
nand U2995 (N_2995,N_614,N_322);
or U2996 (N_2996,N_998,N_1486);
nor U2997 (N_2997,N_1112,N_74);
xor U2998 (N_2998,N_1290,N_206);
nand U2999 (N_2999,N_679,N_1049);
nand U3000 (N_3000,N_2598,N_2939);
nor U3001 (N_3001,N_2134,N_2098);
nand U3002 (N_3002,N_1891,N_2482);
or U3003 (N_3003,N_2761,N_1819);
nand U3004 (N_3004,N_2656,N_2928);
xnor U3005 (N_3005,N_1999,N_2980);
xor U3006 (N_3006,N_1720,N_1586);
nor U3007 (N_3007,N_1803,N_2399);
or U3008 (N_3008,N_2786,N_1686);
nor U3009 (N_3009,N_1664,N_2231);
nand U3010 (N_3010,N_1680,N_2057);
and U3011 (N_3011,N_1647,N_2702);
nor U3012 (N_3012,N_2618,N_2236);
nor U3013 (N_3013,N_2448,N_2974);
nor U3014 (N_3014,N_1637,N_1911);
or U3015 (N_3015,N_2267,N_2903);
and U3016 (N_3016,N_1544,N_2263);
nand U3017 (N_3017,N_2931,N_2204);
or U3018 (N_3018,N_2216,N_1825);
or U3019 (N_3019,N_2308,N_1745);
and U3020 (N_3020,N_2147,N_2438);
and U3021 (N_3021,N_2678,N_1955);
or U3022 (N_3022,N_1638,N_1603);
nand U3023 (N_3023,N_1748,N_2418);
and U3024 (N_3024,N_1564,N_2342);
xor U3025 (N_3025,N_2392,N_2299);
xnor U3026 (N_3026,N_2082,N_2574);
or U3027 (N_3027,N_2461,N_1714);
nor U3028 (N_3028,N_1979,N_2652);
xor U3029 (N_3029,N_2401,N_2967);
nor U3030 (N_3030,N_2156,N_2773);
or U3031 (N_3031,N_2840,N_2377);
and U3032 (N_3032,N_2422,N_2816);
and U3033 (N_3033,N_1857,N_1532);
and U3034 (N_3034,N_2064,N_1867);
or U3035 (N_3035,N_1796,N_1856);
nor U3036 (N_3036,N_2273,N_1770);
nand U3037 (N_3037,N_1579,N_2164);
xnor U3038 (N_3038,N_2076,N_1562);
nand U3039 (N_3039,N_1820,N_1624);
nor U3040 (N_3040,N_2865,N_2311);
xor U3041 (N_3041,N_2805,N_1845);
or U3042 (N_3042,N_2275,N_2628);
or U3043 (N_3043,N_2845,N_2855);
nor U3044 (N_3044,N_1740,N_2352);
or U3045 (N_3045,N_2955,N_1862);
or U3046 (N_3046,N_1518,N_2527);
and U3047 (N_3047,N_1504,N_2649);
or U3048 (N_3048,N_2543,N_2370);
and U3049 (N_3049,N_2991,N_2480);
xnor U3050 (N_3050,N_2243,N_1906);
nand U3051 (N_3051,N_2639,N_1700);
xnor U3052 (N_3052,N_1998,N_2396);
and U3053 (N_3053,N_2703,N_1724);
nand U3054 (N_3054,N_2798,N_2676);
or U3055 (N_3055,N_1789,N_2810);
nand U3056 (N_3056,N_2672,N_2010);
nand U3057 (N_3057,N_1600,N_1951);
nand U3058 (N_3058,N_2320,N_2075);
nor U3059 (N_3059,N_2822,N_2759);
or U3060 (N_3060,N_1635,N_2358);
xor U3061 (N_3061,N_1786,N_2911);
xor U3062 (N_3062,N_2929,N_2686);
or U3063 (N_3063,N_2409,N_2405);
xor U3064 (N_3064,N_2919,N_1697);
or U3065 (N_3065,N_2525,N_1595);
or U3066 (N_3066,N_2030,N_1732);
nor U3067 (N_3067,N_2593,N_1530);
xnor U3068 (N_3068,N_2671,N_1995);
nand U3069 (N_3069,N_2610,N_2096);
nand U3070 (N_3070,N_2270,N_1869);
and U3071 (N_3071,N_2186,N_2682);
xor U3072 (N_3072,N_2580,N_1520);
xor U3073 (N_3073,N_2766,N_2994);
or U3074 (N_3074,N_1588,N_2454);
nor U3075 (N_3075,N_1811,N_2747);
or U3076 (N_3076,N_1914,N_1500);
nand U3077 (N_3077,N_2103,N_2184);
and U3078 (N_3078,N_1773,N_2723);
or U3079 (N_3079,N_2220,N_2424);
or U3080 (N_3080,N_2572,N_2343);
and U3081 (N_3081,N_1528,N_1986);
or U3082 (N_3082,N_1723,N_2657);
nor U3083 (N_3083,N_2149,N_2157);
nand U3084 (N_3084,N_1958,N_2599);
nand U3085 (N_3085,N_2832,N_1941);
nand U3086 (N_3086,N_1960,N_2895);
nor U3087 (N_3087,N_2188,N_2715);
or U3088 (N_3088,N_1980,N_2627);
xnor U3089 (N_3089,N_1580,N_2779);
or U3090 (N_3090,N_1949,N_2592);
and U3091 (N_3091,N_2026,N_2203);
or U3092 (N_3092,N_1590,N_2468);
or U3093 (N_3093,N_1981,N_1717);
xnor U3094 (N_3094,N_1760,N_2675);
xnor U3095 (N_3095,N_1656,N_2576);
xor U3096 (N_3096,N_2927,N_2340);
xnor U3097 (N_3097,N_2882,N_1541);
xor U3098 (N_3098,N_1808,N_2178);
nor U3099 (N_3099,N_2612,N_2518);
or U3100 (N_3100,N_2160,N_1709);
and U3101 (N_3101,N_1550,N_2004);
xor U3102 (N_3102,N_1666,N_2780);
nand U3103 (N_3103,N_2881,N_2017);
nor U3104 (N_3104,N_2522,N_2775);
and U3105 (N_3105,N_2492,N_2710);
and U3106 (N_3106,N_2361,N_2179);
nand U3107 (N_3107,N_1679,N_2506);
and U3108 (N_3108,N_2722,N_2327);
nor U3109 (N_3109,N_2745,N_1944);
and U3110 (N_3110,N_2106,N_2648);
or U3111 (N_3111,N_2207,N_1910);
and U3112 (N_3112,N_2720,N_1633);
nand U3113 (N_3113,N_1552,N_2472);
xor U3114 (N_3114,N_2641,N_2550);
nor U3115 (N_3115,N_1622,N_2037);
nor U3116 (N_3116,N_2508,N_2502);
nor U3117 (N_3117,N_2287,N_1731);
nor U3118 (N_3118,N_2819,N_2651);
nand U3119 (N_3119,N_1946,N_1954);
nor U3120 (N_3120,N_2283,N_1988);
nand U3121 (N_3121,N_2762,N_2079);
or U3122 (N_3122,N_1851,N_1866);
or U3123 (N_3123,N_2210,N_2754);
or U3124 (N_3124,N_1822,N_1618);
xnor U3125 (N_3125,N_2517,N_2215);
nand U3126 (N_3126,N_2459,N_2326);
xor U3127 (N_3127,N_2796,N_2661);
nor U3128 (N_3128,N_2069,N_2013);
and U3129 (N_3129,N_2042,N_2562);
nand U3130 (N_3130,N_2307,N_1883);
or U3131 (N_3131,N_1991,N_2884);
nand U3132 (N_3132,N_2317,N_2238);
xor U3133 (N_3133,N_2379,N_2202);
nand U3134 (N_3134,N_2772,N_2444);
or U3135 (N_3135,N_2137,N_1719);
or U3136 (N_3136,N_2003,N_2801);
nor U3137 (N_3137,N_2229,N_2705);
and U3138 (N_3138,N_1826,N_1792);
xor U3139 (N_3139,N_1940,N_2054);
nor U3140 (N_3140,N_1976,N_1549);
nor U3141 (N_3141,N_1610,N_2680);
nand U3142 (N_3142,N_2826,N_2494);
or U3143 (N_3143,N_2262,N_1928);
xnor U3144 (N_3144,N_2921,N_2029);
and U3145 (N_3145,N_1535,N_2968);
nand U3146 (N_3146,N_2569,N_1896);
or U3147 (N_3147,N_2012,N_2752);
nand U3148 (N_3148,N_1907,N_2892);
nor U3149 (N_3149,N_2503,N_2567);
xor U3150 (N_3150,N_1568,N_2471);
xnor U3151 (N_3151,N_2337,N_2721);
nor U3152 (N_3152,N_1868,N_1750);
xnor U3153 (N_3153,N_2368,N_2066);
nand U3154 (N_3154,N_2746,N_1961);
and U3155 (N_3155,N_2858,N_1702);
or U3156 (N_3156,N_2078,N_2406);
or U3157 (N_3157,N_2445,N_2331);
or U3158 (N_3158,N_2789,N_1699);
and U3159 (N_3159,N_1764,N_2217);
nor U3160 (N_3160,N_1774,N_2616);
xor U3161 (N_3161,N_2212,N_2191);
xor U3162 (N_3162,N_1917,N_2484);
or U3163 (N_3163,N_2047,N_1627);
nand U3164 (N_3164,N_1524,N_2420);
xor U3165 (N_3165,N_1957,N_2554);
and U3166 (N_3166,N_2211,N_1919);
nor U3167 (N_3167,N_2937,N_2450);
xnor U3168 (N_3168,N_1933,N_1519);
xnor U3169 (N_3169,N_2934,N_2032);
nor U3170 (N_3170,N_1834,N_1583);
or U3171 (N_3171,N_2071,N_2831);
xnor U3172 (N_3172,N_1577,N_2105);
xor U3173 (N_3173,N_2828,N_2899);
nand U3174 (N_3174,N_2850,N_2196);
or U3175 (N_3175,N_2001,N_2834);
or U3176 (N_3176,N_2724,N_1754);
nand U3177 (N_3177,N_2027,N_2585);
nand U3178 (N_3178,N_2116,N_2626);
nand U3179 (N_3179,N_2565,N_2898);
xor U3180 (N_3180,N_2988,N_2334);
nor U3181 (N_3181,N_2132,N_1598);
xor U3182 (N_3182,N_2434,N_2741);
or U3183 (N_3183,N_2481,N_2504);
nor U3184 (N_3184,N_1918,N_2976);
nand U3185 (N_3185,N_1643,N_2848);
nand U3186 (N_3186,N_1926,N_2304);
nor U3187 (N_3187,N_2268,N_2925);
xnor U3188 (N_3188,N_1658,N_2764);
xnor U3189 (N_3189,N_2956,N_1685);
or U3190 (N_3190,N_2624,N_1529);
nor U3191 (N_3191,N_2279,N_2523);
or U3192 (N_3192,N_2346,N_2440);
nor U3193 (N_3193,N_2877,N_2049);
xnor U3194 (N_3194,N_2292,N_1776);
nand U3195 (N_3195,N_2168,N_2587);
and U3196 (N_3196,N_2284,N_2175);
or U3197 (N_3197,N_2663,N_2045);
nor U3198 (N_3198,N_2859,N_1641);
or U3199 (N_3199,N_2473,N_2583);
xnor U3200 (N_3200,N_1945,N_2385);
and U3201 (N_3201,N_2095,N_1874);
nand U3202 (N_3202,N_1526,N_1756);
nand U3203 (N_3203,N_2306,N_2535);
nand U3204 (N_3204,N_2594,N_2600);
and U3205 (N_3205,N_2708,N_2851);
nand U3206 (N_3206,N_2922,N_1547);
and U3207 (N_3207,N_2545,N_2208);
and U3208 (N_3208,N_2341,N_2654);
or U3209 (N_3209,N_2142,N_1971);
nand U3210 (N_3210,N_1950,N_2077);
nand U3211 (N_3211,N_2126,N_2665);
nand U3212 (N_3212,N_1782,N_1892);
or U3213 (N_3213,N_2871,N_2059);
or U3214 (N_3214,N_2835,N_1790);
or U3215 (N_3215,N_2662,N_1501);
nand U3216 (N_3216,N_2920,N_1895);
or U3217 (N_3217,N_2139,N_2799);
nand U3218 (N_3218,N_2735,N_2328);
nand U3219 (N_3219,N_1597,N_1670);
or U3220 (N_3220,N_2866,N_2189);
and U3221 (N_3221,N_1585,N_1565);
or U3222 (N_3222,N_2428,N_2932);
nand U3223 (N_3223,N_1694,N_2415);
or U3224 (N_3224,N_2602,N_1841);
xor U3225 (N_3225,N_2246,N_1592);
and U3226 (N_3226,N_1513,N_2297);
and U3227 (N_3227,N_1576,N_2426);
xnor U3228 (N_3228,N_2023,N_2194);
nand U3229 (N_3229,N_2785,N_1713);
nand U3230 (N_3230,N_2908,N_2818);
xor U3231 (N_3231,N_1571,N_2971);
and U3232 (N_3232,N_1959,N_1992);
or U3233 (N_3233,N_2540,N_2345);
nand U3234 (N_3234,N_1924,N_1842);
nor U3235 (N_3235,N_2951,N_2760);
xor U3236 (N_3236,N_2613,N_1932);
nor U3237 (N_3237,N_2528,N_2259);
nand U3238 (N_3238,N_2041,N_2716);
nand U3239 (N_3239,N_1934,N_1650);
nand U3240 (N_3240,N_2916,N_1506);
or U3241 (N_3241,N_2018,N_1757);
nor U3242 (N_3242,N_2734,N_2282);
nor U3243 (N_3243,N_2684,N_2172);
and U3244 (N_3244,N_2040,N_2193);
nand U3245 (N_3245,N_2872,N_2809);
nor U3246 (N_3246,N_1987,N_2803);
nor U3247 (N_3247,N_2114,N_1574);
nand U3248 (N_3248,N_1768,N_2655);
nor U3249 (N_3249,N_1509,N_1561);
or U3250 (N_3250,N_2725,N_1829);
nor U3251 (N_3251,N_1795,N_2784);
nor U3252 (N_3252,N_2751,N_2441);
or U3253 (N_3253,N_2581,N_2640);
xnor U3254 (N_3254,N_1642,N_2659);
xor U3255 (N_3255,N_2356,N_2309);
or U3256 (N_3256,N_1882,N_1688);
nand U3257 (N_3257,N_2996,N_2841);
xnor U3258 (N_3258,N_1502,N_1880);
nand U3259 (N_3259,N_2591,N_2605);
nand U3260 (N_3260,N_2673,N_2091);
and U3261 (N_3261,N_1948,N_1726);
xnor U3262 (N_3262,N_1693,N_1801);
xnor U3263 (N_3263,N_2897,N_1810);
nand U3264 (N_3264,N_1840,N_2470);
xnor U3265 (N_3265,N_2814,N_2589);
nand U3266 (N_3266,N_1831,N_2237);
and U3267 (N_3267,N_1769,N_2874);
nor U3268 (N_3268,N_1742,N_1990);
nand U3269 (N_3269,N_2883,N_2286);
nand U3270 (N_3270,N_2763,N_1712);
and U3271 (N_3271,N_1860,N_2793);
or U3272 (N_3272,N_2008,N_2509);
nand U3273 (N_3273,N_2487,N_2218);
nand U3274 (N_3274,N_1674,N_2395);
nand U3275 (N_3275,N_2363,N_1863);
or U3276 (N_3276,N_1659,N_1969);
nand U3277 (N_3277,N_1781,N_2107);
or U3278 (N_3278,N_1591,N_1983);
and U3279 (N_3279,N_2915,N_1828);
and U3280 (N_3280,N_2669,N_2936);
nand U3281 (N_3281,N_2644,N_2192);
nand U3282 (N_3282,N_2146,N_2436);
and U3283 (N_3283,N_2889,N_2590);
xor U3284 (N_3284,N_2757,N_1607);
xor U3285 (N_3285,N_1937,N_2141);
xnor U3286 (N_3286,N_2120,N_2620);
nand U3287 (N_3287,N_2083,N_2742);
and U3288 (N_3288,N_1739,N_1871);
nor U3289 (N_3289,N_1661,N_2902);
xnor U3290 (N_3290,N_2281,N_1827);
xnor U3291 (N_3291,N_2711,N_2365);
nand U3292 (N_3292,N_1531,N_2529);
nand U3293 (N_3293,N_2240,N_2310);
nand U3294 (N_3294,N_1551,N_1936);
or U3295 (N_3295,N_2435,N_1935);
and U3296 (N_3296,N_2623,N_2694);
or U3297 (N_3297,N_2174,N_1706);
xnor U3298 (N_3298,N_2695,N_2970);
nor U3299 (N_3299,N_1964,N_1692);
or U3300 (N_3300,N_1623,N_1952);
and U3301 (N_3301,N_1545,N_2097);
nand U3302 (N_3302,N_1735,N_2369);
nor U3303 (N_3303,N_2115,N_2578);
xnor U3304 (N_3304,N_2288,N_1909);
nor U3305 (N_3305,N_2312,N_1730);
xor U3306 (N_3306,N_1836,N_2244);
nor U3307 (N_3307,N_2727,N_2778);
or U3308 (N_3308,N_2548,N_2313);
or U3309 (N_3309,N_1695,N_2315);
nand U3310 (N_3310,N_1974,N_2815);
or U3311 (N_3311,N_1558,N_2539);
and U3312 (N_3312,N_2019,N_2333);
nand U3313 (N_3313,N_1852,N_1663);
xor U3314 (N_3314,N_2873,N_2713);
nor U3315 (N_3315,N_1621,N_1744);
xnor U3316 (N_3316,N_1703,N_1596);
and U3317 (N_3317,N_2296,N_2534);
nor U3318 (N_3318,N_2486,N_2726);
and U3319 (N_3319,N_2755,N_2544);
or U3320 (N_3320,N_2489,N_1722);
xnor U3321 (N_3321,N_2689,N_2087);
nand U3322 (N_3322,N_2635,N_1648);
xor U3323 (N_3323,N_2560,N_2693);
or U3324 (N_3324,N_2802,N_1848);
nor U3325 (N_3325,N_1890,N_2941);
nor U3326 (N_3326,N_2960,N_2190);
xor U3327 (N_3327,N_1727,N_2575);
and U3328 (N_3328,N_2719,N_2986);
and U3329 (N_3329,N_1625,N_1927);
nand U3330 (N_3330,N_1689,N_2009);
xor U3331 (N_3331,N_2099,N_2375);
and U3332 (N_3332,N_1913,N_2953);
or U3333 (N_3333,N_2443,N_2280);
nor U3334 (N_3334,N_2777,N_1861);
nor U3335 (N_3335,N_2151,N_2324);
nor U3336 (N_3336,N_2997,N_1900);
or U3337 (N_3337,N_1609,N_1962);
or U3338 (N_3338,N_2596,N_2864);
and U3339 (N_3339,N_1525,N_2788);
or U3340 (N_3340,N_1865,N_2242);
nor U3341 (N_3341,N_2812,N_2603);
nor U3342 (N_3342,N_2571,N_2500);
and U3343 (N_3343,N_2170,N_2769);
or U3344 (N_3344,N_2442,N_2336);
nand U3345 (N_3345,N_2022,N_1678);
and U3346 (N_3346,N_1575,N_1787);
and U3347 (N_3347,N_1807,N_2414);
or U3348 (N_3348,N_1602,N_1839);
nor U3349 (N_3349,N_2736,N_1718);
nand U3350 (N_3350,N_1902,N_1984);
xnor U3351 (N_3351,N_2371,N_2579);
and U3352 (N_3352,N_2800,N_2373);
nor U3353 (N_3353,N_2039,N_1997);
and U3354 (N_3354,N_2985,N_2833);
and U3355 (N_3355,N_1676,N_2425);
and U3356 (N_3356,N_1746,N_2072);
or U3357 (N_3357,N_1503,N_1557);
and U3358 (N_3358,N_2901,N_1904);
and U3359 (N_3359,N_1707,N_1893);
nor U3360 (N_3360,N_1527,N_1855);
xnor U3361 (N_3361,N_2278,N_2080);
xnor U3362 (N_3362,N_2381,N_1830);
and U3363 (N_3363,N_2260,N_2948);
and U3364 (N_3364,N_2199,N_1687);
nor U3365 (N_3365,N_1738,N_2364);
nand U3366 (N_3366,N_1601,N_2225);
nand U3367 (N_3367,N_1850,N_2094);
or U3368 (N_3368,N_1805,N_2180);
xor U3369 (N_3369,N_1884,N_1751);
or U3370 (N_3370,N_1996,N_2732);
nand U3371 (N_3371,N_2163,N_1705);
nand U3372 (N_3372,N_1716,N_2475);
nor U3373 (N_3373,N_2885,N_2838);
xor U3374 (N_3374,N_2496,N_2771);
and U3375 (N_3375,N_1881,N_1762);
or U3376 (N_3376,N_2677,N_2634);
nor U3377 (N_3377,N_2891,N_2226);
and U3378 (N_3378,N_2923,N_2791);
xor U3379 (N_3379,N_2144,N_1912);
or U3380 (N_3380,N_2704,N_2547);
nor U3381 (N_3381,N_1546,N_1794);
xnor U3382 (N_3382,N_1652,N_1899);
nor U3383 (N_3383,N_1734,N_2538);
nor U3384 (N_3384,N_1741,N_2376);
and U3385 (N_3385,N_2431,N_2501);
nand U3386 (N_3386,N_1885,N_1684);
nand U3387 (N_3387,N_2362,N_2387);
nand U3388 (N_3388,N_1505,N_2338);
nand U3389 (N_3389,N_2255,N_1626);
nor U3390 (N_3390,N_2650,N_2185);
or U3391 (N_3391,N_2491,N_1543);
nor U3392 (N_3392,N_2118,N_2860);
nor U3393 (N_3393,N_2601,N_2797);
and U3394 (N_3394,N_2335,N_2021);
xor U3395 (N_3395,N_2514,N_2645);
xnor U3396 (N_3396,N_1886,N_2697);
xor U3397 (N_3397,N_2016,N_2391);
nor U3398 (N_3398,N_2969,N_2637);
and U3399 (N_3399,N_2944,N_2161);
nand U3400 (N_3400,N_2493,N_1875);
xor U3401 (N_3401,N_2926,N_2987);
nand U3402 (N_3402,N_2169,N_2382);
nand U3403 (N_3403,N_1672,N_2767);
xor U3404 (N_3404,N_1548,N_1930);
nor U3405 (N_3405,N_2148,N_2388);
nand U3406 (N_3406,N_1517,N_2349);
or U3407 (N_3407,N_2323,N_2692);
nand U3408 (N_3408,N_2584,N_2488);
and U3409 (N_3409,N_1662,N_2679);
nor U3410 (N_3410,N_1521,N_2606);
xnor U3411 (N_3411,N_1943,N_1922);
nor U3412 (N_3412,N_2905,N_2269);
xor U3413 (N_3413,N_2261,N_2563);
nand U3414 (N_3414,N_1847,N_1755);
nand U3415 (N_3415,N_2293,N_2930);
xnor U3416 (N_3416,N_2537,N_1814);
nor U3417 (N_3417,N_1898,N_2516);
or U3418 (N_3418,N_1512,N_2294);
nand U3419 (N_3419,N_2564,N_2530);
nand U3420 (N_3420,N_2412,N_2419);
nand U3421 (N_3421,N_1654,N_2521);
xor U3422 (N_3422,N_1977,N_2681);
nor U3423 (N_3423,N_1690,N_2121);
nand U3424 (N_3424,N_2028,N_2133);
xnor U3425 (N_3425,N_2875,N_1594);
or U3426 (N_3426,N_2366,N_2397);
and U3427 (N_3427,N_2894,N_2089);
and U3428 (N_3428,N_2515,N_2140);
xor U3429 (N_3429,N_2453,N_2914);
nor U3430 (N_3430,N_2355,N_2876);
nand U3431 (N_3431,N_2947,N_2108);
or U3432 (N_3432,N_2531,N_2479);
xnor U3433 (N_3433,N_1823,N_2224);
or U3434 (N_3434,N_1715,N_2737);
nand U3435 (N_3435,N_2992,N_2394);
or U3436 (N_3436,N_1667,N_1864);
nand U3437 (N_3437,N_1728,N_1966);
or U3438 (N_3438,N_1779,N_1806);
nor U3439 (N_3439,N_2981,N_2432);
xor U3440 (N_3440,N_2330,N_2466);
and U3441 (N_3441,N_2256,N_2643);
nand U3442 (N_3442,N_2890,N_2808);
nor U3443 (N_3443,N_2497,N_1683);
nor U3444 (N_3444,N_2000,N_1780);
nor U3445 (N_3445,N_2474,N_2556);
xnor U3446 (N_3446,N_2794,N_2664);
nand U3447 (N_3447,N_2232,N_2817);
or U3448 (N_3448,N_2582,N_1587);
or U3449 (N_3449,N_2209,N_2264);
xnor U3450 (N_3450,N_1605,N_2621);
nand U3451 (N_3451,N_2555,N_2429);
xor U3452 (N_3452,N_2081,N_1573);
and U3453 (N_3453,N_2646,N_2520);
nand U3454 (N_3454,N_2253,N_1763);
and U3455 (N_3455,N_1675,N_2943);
xnor U3456 (N_3456,N_2933,N_2350);
nand U3457 (N_3457,N_2744,N_1572);
and U3458 (N_3458,N_2086,N_2046);
or U3459 (N_3459,N_2322,N_2050);
or U3460 (N_3460,N_1761,N_2984);
nand U3461 (N_3461,N_1838,N_2542);
nand U3462 (N_3462,N_2455,N_1634);
xnor U3463 (N_3463,N_2378,N_2549);
xnor U3464 (N_3464,N_2245,N_2187);
or U3465 (N_3465,N_2034,N_2511);
nor U3466 (N_3466,N_2909,N_2325);
and U3467 (N_3467,N_2577,N_1818);
nor U3468 (N_3468,N_2295,N_2913);
and U3469 (N_3469,N_2614,N_2403);
or U3470 (N_3470,N_2007,N_2155);
and U3471 (N_3471,N_2573,N_2490);
xor U3472 (N_3472,N_1593,N_2696);
nor U3473 (N_3473,N_1870,N_2439);
nor U3474 (N_3474,N_2728,N_2667);
nand U3475 (N_3475,N_2965,N_2526);
xor U3476 (N_3476,N_1514,N_2546);
nor U3477 (N_3477,N_2276,N_1733);
xor U3478 (N_3478,N_2888,N_2036);
nor U3479 (N_3479,N_1704,N_2688);
and U3480 (N_3480,N_2867,N_1965);
or U3481 (N_3481,N_2206,N_1536);
and U3482 (N_3482,N_1931,N_2781);
xnor U3483 (N_3483,N_1853,N_2712);
nand U3484 (N_3484,N_2005,N_2125);
xnor U3485 (N_3485,N_2052,N_1534);
or U3486 (N_3486,N_1671,N_1677);
nor U3487 (N_3487,N_2512,N_2128);
nand U3488 (N_3488,N_2999,N_1872);
nor U3489 (N_3489,N_1515,N_2910);
or U3490 (N_3490,N_2239,N_2658);
xnor U3491 (N_3491,N_2853,N_2499);
or U3492 (N_3492,N_2557,N_2464);
xor U3493 (N_3493,N_2837,N_1752);
xor U3494 (N_3494,N_2854,N_2266);
nor U3495 (N_3495,N_1766,N_1632);
and U3496 (N_3496,N_2451,N_1846);
nor U3497 (N_3497,N_2233,N_2699);
and U3498 (N_3498,N_1813,N_2924);
or U3499 (N_3499,N_2998,N_2880);
nor U3500 (N_3500,N_2668,N_2374);
xor U3501 (N_3501,N_1533,N_1584);
nand U3502 (N_3502,N_2958,N_2604);
or U3503 (N_3503,N_1783,N_2433);
or U3504 (N_3504,N_1556,N_2957);
nor U3505 (N_3505,N_2068,N_2961);
and U3506 (N_3506,N_2683,N_2061);
or U3507 (N_3507,N_1655,N_2271);
and U3508 (N_3508,N_2177,N_1832);
or U3509 (N_3509,N_2687,N_1644);
or U3510 (N_3510,N_2990,N_2249);
nor U3511 (N_3511,N_1973,N_1710);
nor U3512 (N_3512,N_1878,N_2561);
or U3513 (N_3513,N_1815,N_2570);
or U3514 (N_3514,N_2247,N_2862);
and U3515 (N_3515,N_1538,N_2863);
and U3516 (N_3516,N_2123,N_2015);
nand U3517 (N_3517,N_2129,N_2975);
or U3518 (N_3518,N_2413,N_2507);
xor U3519 (N_3519,N_2265,N_2241);
nor U3520 (N_3520,N_2896,N_1982);
nand U3521 (N_3521,N_2360,N_2254);
or U3522 (N_3522,N_2055,N_2353);
nand U3523 (N_3523,N_2607,N_2993);
and U3524 (N_3524,N_2774,N_2390);
and U3525 (N_3525,N_2790,N_2093);
xor U3526 (N_3526,N_2989,N_1619);
and U3527 (N_3527,N_1660,N_2830);
xor U3528 (N_3528,N_2014,N_2868);
nand U3529 (N_3529,N_2033,N_2408);
nand U3530 (N_3530,N_2213,N_2964);
nand U3531 (N_3531,N_2973,N_2940);
xnor U3532 (N_3532,N_2740,N_1743);
nor U3533 (N_3533,N_1873,N_2171);
nor U3534 (N_3534,N_2617,N_1978);
or U3535 (N_3535,N_2044,N_2824);
and U3536 (N_3536,N_1802,N_1698);
nor U3537 (N_3537,N_2285,N_1809);
xnor U3538 (N_3538,N_2768,N_1889);
nand U3539 (N_3539,N_2787,N_2938);
nor U3540 (N_3540,N_1629,N_2205);
nor U3541 (N_3541,N_1725,N_2329);
nand U3542 (N_3542,N_2197,N_1901);
xnor U3543 (N_3543,N_2359,N_1975);
nor U3544 (N_3544,N_2417,N_2056);
xnor U3545 (N_3545,N_1589,N_2465);
and U3546 (N_3546,N_1553,N_1877);
nor U3547 (N_3547,N_1833,N_2101);
nor U3548 (N_3548,N_2136,N_2104);
and U3549 (N_3549,N_1791,N_1908);
nand U3550 (N_3550,N_2060,N_2950);
nand U3551 (N_3551,N_2138,N_2608);
nor U3552 (N_3552,N_2402,N_2456);
xnor U3553 (N_3553,N_1523,N_2063);
xnor U3554 (N_3554,N_2222,N_2298);
nand U3555 (N_3555,N_1785,N_2462);
or U3556 (N_3556,N_1804,N_2536);
nor U3557 (N_3557,N_2478,N_2303);
nand U3558 (N_3558,N_1620,N_2458);
or U3559 (N_3559,N_2006,N_1611);
nand U3560 (N_3560,N_2631,N_2053);
xor U3561 (N_3561,N_2935,N_2219);
xnor U3562 (N_3562,N_2348,N_1888);
and U3563 (N_3563,N_1915,N_2959);
nand U3564 (N_3564,N_1793,N_2861);
or U3565 (N_3565,N_2558,N_2452);
nand U3566 (N_3566,N_2670,N_2846);
nor U3567 (N_3567,N_1905,N_1612);
xor U3568 (N_3568,N_2559,N_2700);
xnor U3569 (N_3569,N_2393,N_1972);
xor U3570 (N_3570,N_2130,N_2782);
nand U3571 (N_3571,N_2386,N_1985);
and U3572 (N_3572,N_1649,N_2449);
or U3573 (N_3573,N_1797,N_2918);
or U3574 (N_3574,N_2302,N_2423);
nand U3575 (N_3575,N_2446,N_2532);
or U3576 (N_3576,N_2900,N_2383);
xnor U3577 (N_3577,N_2167,N_2886);
nand U3578 (N_3578,N_2709,N_1925);
and U3579 (N_3579,N_1858,N_2945);
and U3580 (N_3580,N_2380,N_1758);
xor U3581 (N_3581,N_1708,N_2251);
or U3582 (N_3582,N_1854,N_2483);
or U3583 (N_3583,N_2852,N_2421);
and U3584 (N_3584,N_2201,N_2113);
or U3585 (N_3585,N_2660,N_2733);
xnor U3586 (N_3586,N_2743,N_1897);
nor U3587 (N_3587,N_2729,N_2917);
and U3588 (N_3588,N_1691,N_2159);
nor U3589 (N_3589,N_2806,N_2291);
nor U3590 (N_3590,N_2776,N_1508);
and U3591 (N_3591,N_2002,N_2811);
nor U3592 (N_3592,N_2551,N_1887);
nand U3593 (N_3593,N_2165,N_2351);
nor U3594 (N_3594,N_1879,N_2274);
or U3595 (N_3595,N_2666,N_1923);
nor U3596 (N_3596,N_2907,N_1696);
nor U3597 (N_3597,N_2117,N_2622);
xor U3598 (N_3598,N_2820,N_2879);
nand U3599 (N_3599,N_2318,N_2731);
or U3600 (N_3600,N_2485,N_2813);
and U3601 (N_3601,N_2354,N_1507);
xnor U3602 (N_3602,N_2062,N_2691);
or U3603 (N_3603,N_1682,N_2150);
and U3604 (N_3604,N_2597,N_1765);
and U3605 (N_3605,N_2717,N_2463);
and U3606 (N_3606,N_1614,N_1929);
and U3607 (N_3607,N_1665,N_2690);
xnor U3608 (N_3608,N_1968,N_1798);
and U3609 (N_3609,N_2615,N_2427);
xnor U3610 (N_3610,N_2758,N_1615);
or U3611 (N_3611,N_2519,N_2119);
nand U3612 (N_3612,N_1560,N_2065);
nor U3613 (N_3613,N_2102,N_2416);
and U3614 (N_3614,N_2200,N_2344);
nand U3615 (N_3615,N_2750,N_1894);
xnor U3616 (N_3616,N_2823,N_2738);
and U3617 (N_3617,N_2946,N_2301);
or U3618 (N_3618,N_2541,N_2638);
or U3619 (N_3619,N_2857,N_2795);
xor U3620 (N_3620,N_1921,N_2870);
nor U3621 (N_3621,N_2619,N_1788);
nor U3622 (N_3622,N_1799,N_2701);
xor U3623 (N_3623,N_1522,N_1749);
xnor U3624 (N_3624,N_2739,N_2829);
or U3625 (N_3625,N_2887,N_2625);
xor U3626 (N_3626,N_2223,N_2642);
nor U3627 (N_3627,N_2124,N_2404);
xnor U3628 (N_3628,N_2632,N_1653);
nor U3629 (N_3629,N_2804,N_1636);
and U3630 (N_3630,N_2552,N_2533);
and U3631 (N_3631,N_2176,N_2807);
nand U3632 (N_3632,N_1630,N_2074);
nor U3633 (N_3633,N_2143,N_2674);
and U3634 (N_3634,N_2706,N_2025);
or U3635 (N_3635,N_2070,N_2995);
nor U3636 (N_3636,N_2765,N_1993);
nor U3637 (N_3637,N_2770,N_2316);
and U3638 (N_3638,N_1824,N_2088);
nand U3639 (N_3639,N_1554,N_1963);
and U3640 (N_3640,N_2092,N_2718);
and U3641 (N_3641,N_1747,N_2277);
nor U3642 (N_3642,N_2792,N_2653);
nor U3643 (N_3643,N_2847,N_2127);
nand U3644 (N_3644,N_1772,N_1778);
and U3645 (N_3645,N_2633,N_1616);
nand U3646 (N_3646,N_1967,N_2949);
and U3647 (N_3647,N_2173,N_2611);
nand U3648 (N_3648,N_1821,N_2595);
nor U3649 (N_3649,N_1903,N_2357);
nor U3650 (N_3650,N_2842,N_2031);
nor U3651 (N_3651,N_2162,N_2166);
nand U3652 (N_3652,N_2982,N_2145);
nand U3653 (N_3653,N_2112,N_2839);
xnor U3654 (N_3654,N_2783,N_2869);
nand U3655 (N_3655,N_2154,N_2158);
nor U3656 (N_3656,N_2195,N_2460);
or U3657 (N_3657,N_2339,N_1606);
and U3658 (N_3658,N_2467,N_2630);
nor U3659 (N_3659,N_1669,N_2024);
or U3660 (N_3660,N_1775,N_2252);
xnor U3661 (N_3661,N_2111,N_2020);
nand U3662 (N_3662,N_1582,N_2749);
xor U3663 (N_3663,N_2398,N_2011);
xor U3664 (N_3664,N_2878,N_2698);
nor U3665 (N_3665,N_2321,N_2979);
and U3666 (N_3666,N_2437,N_1617);
nor U3667 (N_3667,N_2476,N_2043);
xor U3668 (N_3668,N_2153,N_2250);
or U3669 (N_3669,N_1859,N_1784);
or U3670 (N_3670,N_2319,N_2085);
xor U3671 (N_3671,N_1729,N_1510);
xor U3672 (N_3672,N_2963,N_2714);
xnor U3673 (N_3673,N_2372,N_2430);
nand U3674 (N_3674,N_2477,N_2505);
xnor U3675 (N_3675,N_2152,N_2182);
nand U3676 (N_3676,N_2447,N_2495);
or U3677 (N_3677,N_2131,N_1578);
xnor U3678 (N_3678,N_2912,N_1711);
or U3679 (N_3679,N_2214,N_2821);
xor U3680 (N_3680,N_2906,N_2513);
nor U3681 (N_3681,N_1938,N_2305);
nand U3682 (N_3682,N_1920,N_2257);
or U3683 (N_3683,N_1701,N_2753);
xor U3684 (N_3684,N_2051,N_1604);
and U3685 (N_3685,N_1628,N_2198);
xnor U3686 (N_3686,N_2566,N_1559);
and U3687 (N_3687,N_1989,N_1539);
nor U3688 (N_3688,N_1939,N_2685);
xor U3689 (N_3689,N_2411,N_2221);
nor U3690 (N_3690,N_2110,N_2942);
or U3691 (N_3691,N_1651,N_2636);
and U3692 (N_3692,N_2400,N_2272);
or U3693 (N_3693,N_1753,N_1812);
nor U3694 (N_3694,N_2836,N_2183);
xor U3695 (N_3695,N_1767,N_1566);
nand U3696 (N_3696,N_1942,N_2588);
and U3697 (N_3697,N_1816,N_2084);
nand U3698 (N_3698,N_1876,N_2977);
and U3699 (N_3699,N_2181,N_2893);
xor U3700 (N_3700,N_2230,N_2952);
xnor U3701 (N_3701,N_2038,N_2227);
and U3702 (N_3702,N_2347,N_2258);
and U3703 (N_3703,N_2248,N_2469);
and U3704 (N_3704,N_2609,N_1736);
or U3705 (N_3705,N_2289,N_2827);
nor U3706 (N_3706,N_2843,N_1956);
and U3707 (N_3707,N_1759,N_1657);
nor U3708 (N_3708,N_2978,N_1668);
xnor U3709 (N_3709,N_2966,N_2234);
nor U3710 (N_3710,N_2825,N_2100);
nand U3711 (N_3711,N_2983,N_2332);
and U3712 (N_3712,N_1916,N_1563);
nand U3713 (N_3713,N_2090,N_2904);
or U3714 (N_3714,N_1947,N_2389);
nor U3715 (N_3715,N_1953,N_2035);
xor U3716 (N_3716,N_2300,N_2553);
and U3717 (N_3717,N_2135,N_2058);
xnor U3718 (N_3718,N_1570,N_2849);
xor U3719 (N_3719,N_1771,N_1970);
nand U3720 (N_3720,N_2510,N_1849);
nor U3721 (N_3721,N_2498,N_1640);
xnor U3722 (N_3722,N_1673,N_1540);
and U3723 (N_3723,N_2067,N_1631);
xor U3724 (N_3724,N_1581,N_2647);
nor U3725 (N_3725,N_2748,N_1511);
xor U3726 (N_3726,N_1567,N_2844);
xor U3727 (N_3727,N_1843,N_1599);
xnor U3728 (N_3728,N_1835,N_2235);
and U3729 (N_3729,N_1537,N_1844);
and U3730 (N_3730,N_2122,N_1646);
nand U3731 (N_3731,N_2954,N_1837);
or U3732 (N_3732,N_1569,N_2856);
nor U3733 (N_3733,N_1721,N_1639);
nand U3734 (N_3734,N_1613,N_1800);
and U3735 (N_3735,N_2407,N_1737);
xor U3736 (N_3736,N_2962,N_2707);
or U3737 (N_3737,N_2228,N_2109);
xor U3738 (N_3738,N_2756,N_2524);
or U3739 (N_3739,N_2073,N_1516);
and U3740 (N_3740,N_2410,N_2367);
and U3741 (N_3741,N_2629,N_1777);
xnor U3742 (N_3742,N_1817,N_2314);
nand U3743 (N_3743,N_1555,N_1681);
and U3744 (N_3744,N_2586,N_1608);
xor U3745 (N_3745,N_2730,N_2290);
nor U3746 (N_3746,N_1645,N_2384);
nor U3747 (N_3747,N_2048,N_2568);
nand U3748 (N_3748,N_2457,N_1994);
or U3749 (N_3749,N_2972,N_1542);
xnor U3750 (N_3750,N_2146,N_1646);
nand U3751 (N_3751,N_2796,N_1870);
nor U3752 (N_3752,N_2788,N_2144);
and U3753 (N_3753,N_2936,N_2369);
or U3754 (N_3754,N_2749,N_2896);
and U3755 (N_3755,N_2718,N_1641);
nor U3756 (N_3756,N_2941,N_2001);
nand U3757 (N_3757,N_2568,N_2040);
nor U3758 (N_3758,N_2475,N_2097);
nor U3759 (N_3759,N_2092,N_1638);
and U3760 (N_3760,N_2123,N_2467);
xor U3761 (N_3761,N_2320,N_1820);
nor U3762 (N_3762,N_1687,N_1860);
and U3763 (N_3763,N_1828,N_1541);
nand U3764 (N_3764,N_1545,N_2883);
nor U3765 (N_3765,N_2847,N_2098);
nor U3766 (N_3766,N_2541,N_2138);
and U3767 (N_3767,N_2328,N_1793);
nand U3768 (N_3768,N_2118,N_2991);
and U3769 (N_3769,N_2410,N_2113);
nor U3770 (N_3770,N_2066,N_2163);
nand U3771 (N_3771,N_1928,N_2361);
xnor U3772 (N_3772,N_1971,N_2655);
nor U3773 (N_3773,N_2927,N_2124);
or U3774 (N_3774,N_1577,N_2195);
nor U3775 (N_3775,N_1669,N_2830);
xnor U3776 (N_3776,N_2212,N_2775);
xnor U3777 (N_3777,N_2950,N_2339);
nand U3778 (N_3778,N_1973,N_2748);
and U3779 (N_3779,N_2964,N_2470);
nor U3780 (N_3780,N_1577,N_1966);
nor U3781 (N_3781,N_2936,N_2857);
xor U3782 (N_3782,N_2836,N_2561);
and U3783 (N_3783,N_1649,N_1879);
or U3784 (N_3784,N_2695,N_1591);
nor U3785 (N_3785,N_2807,N_2644);
nor U3786 (N_3786,N_2781,N_1697);
xor U3787 (N_3787,N_2157,N_1807);
xnor U3788 (N_3788,N_2626,N_1712);
and U3789 (N_3789,N_1520,N_2353);
and U3790 (N_3790,N_1775,N_2124);
and U3791 (N_3791,N_2534,N_2706);
or U3792 (N_3792,N_2944,N_2531);
xor U3793 (N_3793,N_2524,N_1819);
nor U3794 (N_3794,N_2131,N_2643);
or U3795 (N_3795,N_2465,N_2893);
xor U3796 (N_3796,N_1960,N_2898);
nor U3797 (N_3797,N_2063,N_2565);
nand U3798 (N_3798,N_2622,N_2135);
and U3799 (N_3799,N_1786,N_2977);
or U3800 (N_3800,N_1641,N_1961);
and U3801 (N_3801,N_2897,N_2439);
or U3802 (N_3802,N_2675,N_2844);
or U3803 (N_3803,N_2686,N_2061);
xor U3804 (N_3804,N_1811,N_2197);
nor U3805 (N_3805,N_2779,N_2258);
nand U3806 (N_3806,N_2898,N_2658);
or U3807 (N_3807,N_2727,N_2690);
nand U3808 (N_3808,N_2178,N_2204);
nand U3809 (N_3809,N_2956,N_2242);
xnor U3810 (N_3810,N_2956,N_1523);
nor U3811 (N_3811,N_2938,N_2860);
and U3812 (N_3812,N_1859,N_2562);
or U3813 (N_3813,N_2856,N_2121);
nand U3814 (N_3814,N_2529,N_1901);
nor U3815 (N_3815,N_2060,N_2440);
and U3816 (N_3816,N_2268,N_2682);
xnor U3817 (N_3817,N_2997,N_1897);
nand U3818 (N_3818,N_1905,N_2786);
nor U3819 (N_3819,N_2794,N_2914);
nor U3820 (N_3820,N_1922,N_2444);
nand U3821 (N_3821,N_2931,N_2153);
nand U3822 (N_3822,N_2229,N_2922);
or U3823 (N_3823,N_2287,N_2898);
and U3824 (N_3824,N_2804,N_2260);
xor U3825 (N_3825,N_2717,N_2755);
nand U3826 (N_3826,N_2113,N_2547);
nand U3827 (N_3827,N_2793,N_1708);
xnor U3828 (N_3828,N_1668,N_2982);
xor U3829 (N_3829,N_2175,N_2351);
and U3830 (N_3830,N_2163,N_1933);
or U3831 (N_3831,N_2025,N_2456);
and U3832 (N_3832,N_2397,N_2737);
nor U3833 (N_3833,N_2551,N_2902);
xor U3834 (N_3834,N_1759,N_1768);
xor U3835 (N_3835,N_1726,N_2912);
nor U3836 (N_3836,N_2211,N_2358);
or U3837 (N_3837,N_1750,N_2879);
or U3838 (N_3838,N_1601,N_2695);
nor U3839 (N_3839,N_2117,N_2142);
xor U3840 (N_3840,N_2593,N_2298);
xnor U3841 (N_3841,N_2663,N_2302);
and U3842 (N_3842,N_2188,N_2766);
xnor U3843 (N_3843,N_2043,N_1515);
xor U3844 (N_3844,N_2542,N_2432);
xnor U3845 (N_3845,N_2161,N_2729);
xnor U3846 (N_3846,N_1573,N_1947);
and U3847 (N_3847,N_2311,N_1562);
xor U3848 (N_3848,N_2627,N_1859);
nor U3849 (N_3849,N_2694,N_1657);
and U3850 (N_3850,N_2699,N_1917);
and U3851 (N_3851,N_1557,N_1906);
and U3852 (N_3852,N_1853,N_2447);
or U3853 (N_3853,N_2801,N_2716);
or U3854 (N_3854,N_2515,N_2520);
and U3855 (N_3855,N_2214,N_1800);
and U3856 (N_3856,N_2563,N_1901);
xor U3857 (N_3857,N_2593,N_1814);
nor U3858 (N_3858,N_1851,N_1728);
nand U3859 (N_3859,N_2277,N_2960);
nand U3860 (N_3860,N_2207,N_1834);
and U3861 (N_3861,N_2084,N_2036);
or U3862 (N_3862,N_2849,N_1627);
or U3863 (N_3863,N_1961,N_2854);
nand U3864 (N_3864,N_2452,N_2272);
and U3865 (N_3865,N_2731,N_1847);
or U3866 (N_3866,N_2475,N_2497);
nand U3867 (N_3867,N_2874,N_2802);
nor U3868 (N_3868,N_1915,N_2411);
and U3869 (N_3869,N_1525,N_2725);
nor U3870 (N_3870,N_1636,N_1806);
and U3871 (N_3871,N_2905,N_1753);
nand U3872 (N_3872,N_2683,N_1569);
nor U3873 (N_3873,N_2367,N_2332);
or U3874 (N_3874,N_1765,N_2127);
and U3875 (N_3875,N_2307,N_1552);
xnor U3876 (N_3876,N_2917,N_2531);
and U3877 (N_3877,N_2480,N_1844);
xor U3878 (N_3878,N_1666,N_1557);
nor U3879 (N_3879,N_2871,N_2758);
nor U3880 (N_3880,N_2667,N_2119);
or U3881 (N_3881,N_1974,N_2730);
or U3882 (N_3882,N_2234,N_2616);
or U3883 (N_3883,N_2454,N_1963);
and U3884 (N_3884,N_2126,N_1672);
xor U3885 (N_3885,N_1782,N_2325);
and U3886 (N_3886,N_1926,N_1851);
nor U3887 (N_3887,N_2688,N_1642);
xor U3888 (N_3888,N_1898,N_2815);
nor U3889 (N_3889,N_1852,N_1757);
nand U3890 (N_3890,N_2930,N_2119);
or U3891 (N_3891,N_1973,N_2322);
xnor U3892 (N_3892,N_2343,N_2729);
or U3893 (N_3893,N_1943,N_2639);
nor U3894 (N_3894,N_2378,N_2214);
xnor U3895 (N_3895,N_1654,N_2552);
xor U3896 (N_3896,N_2601,N_2805);
or U3897 (N_3897,N_2041,N_1648);
or U3898 (N_3898,N_1876,N_2704);
xor U3899 (N_3899,N_2967,N_1959);
nand U3900 (N_3900,N_2463,N_1572);
nand U3901 (N_3901,N_2308,N_2541);
nand U3902 (N_3902,N_2678,N_2875);
or U3903 (N_3903,N_2000,N_2817);
or U3904 (N_3904,N_2685,N_2973);
or U3905 (N_3905,N_2795,N_2955);
and U3906 (N_3906,N_2140,N_1746);
nor U3907 (N_3907,N_2400,N_1848);
or U3908 (N_3908,N_2312,N_2576);
or U3909 (N_3909,N_1746,N_2735);
xor U3910 (N_3910,N_2340,N_2020);
and U3911 (N_3911,N_1853,N_1821);
nand U3912 (N_3912,N_2923,N_1529);
xor U3913 (N_3913,N_1801,N_1653);
and U3914 (N_3914,N_2104,N_2283);
or U3915 (N_3915,N_1890,N_2576);
or U3916 (N_3916,N_1762,N_1786);
xor U3917 (N_3917,N_2558,N_2576);
xor U3918 (N_3918,N_2178,N_1549);
xor U3919 (N_3919,N_2272,N_1578);
nor U3920 (N_3920,N_1994,N_2738);
nor U3921 (N_3921,N_2561,N_2083);
or U3922 (N_3922,N_2250,N_1507);
and U3923 (N_3923,N_2817,N_2833);
and U3924 (N_3924,N_2010,N_1999);
and U3925 (N_3925,N_2217,N_1717);
nor U3926 (N_3926,N_1564,N_2183);
xor U3927 (N_3927,N_2493,N_2332);
or U3928 (N_3928,N_2583,N_2054);
xor U3929 (N_3929,N_1752,N_2089);
and U3930 (N_3930,N_1542,N_2848);
nand U3931 (N_3931,N_2218,N_2628);
nor U3932 (N_3932,N_2349,N_1695);
and U3933 (N_3933,N_1506,N_2147);
nand U3934 (N_3934,N_2828,N_2655);
xnor U3935 (N_3935,N_1941,N_1682);
or U3936 (N_3936,N_2702,N_2552);
nand U3937 (N_3937,N_2465,N_2293);
nor U3938 (N_3938,N_2088,N_2915);
and U3939 (N_3939,N_2863,N_2656);
nor U3940 (N_3940,N_1993,N_2327);
or U3941 (N_3941,N_1872,N_2122);
and U3942 (N_3942,N_2127,N_2197);
nor U3943 (N_3943,N_2120,N_2220);
xor U3944 (N_3944,N_1814,N_2368);
xor U3945 (N_3945,N_2533,N_2625);
nor U3946 (N_3946,N_1766,N_1589);
and U3947 (N_3947,N_2270,N_2779);
nand U3948 (N_3948,N_1979,N_2766);
or U3949 (N_3949,N_1698,N_2163);
or U3950 (N_3950,N_2458,N_2770);
xor U3951 (N_3951,N_1873,N_1643);
or U3952 (N_3952,N_1571,N_2794);
nand U3953 (N_3953,N_2595,N_2429);
or U3954 (N_3954,N_1756,N_1933);
or U3955 (N_3955,N_2558,N_1686);
xnor U3956 (N_3956,N_1544,N_1623);
and U3957 (N_3957,N_2897,N_2903);
nor U3958 (N_3958,N_1531,N_2027);
nor U3959 (N_3959,N_1944,N_2343);
nor U3960 (N_3960,N_2023,N_2779);
xor U3961 (N_3961,N_2560,N_2465);
or U3962 (N_3962,N_2792,N_1839);
xnor U3963 (N_3963,N_2846,N_2847);
nand U3964 (N_3964,N_2010,N_2456);
xnor U3965 (N_3965,N_2603,N_2326);
and U3966 (N_3966,N_2745,N_2137);
nor U3967 (N_3967,N_2101,N_2127);
nand U3968 (N_3968,N_2688,N_2172);
xnor U3969 (N_3969,N_2753,N_2123);
nor U3970 (N_3970,N_2939,N_1547);
or U3971 (N_3971,N_2831,N_1912);
nor U3972 (N_3972,N_1975,N_2121);
nor U3973 (N_3973,N_1846,N_2395);
xor U3974 (N_3974,N_2887,N_2330);
xor U3975 (N_3975,N_2955,N_1757);
or U3976 (N_3976,N_1981,N_2100);
or U3977 (N_3977,N_2000,N_2329);
nor U3978 (N_3978,N_1650,N_1890);
or U3979 (N_3979,N_2493,N_2596);
or U3980 (N_3980,N_2230,N_2675);
and U3981 (N_3981,N_2276,N_2525);
nand U3982 (N_3982,N_1786,N_2943);
nand U3983 (N_3983,N_2480,N_2176);
nand U3984 (N_3984,N_1817,N_1876);
nor U3985 (N_3985,N_2498,N_2358);
and U3986 (N_3986,N_2025,N_2007);
xnor U3987 (N_3987,N_1928,N_2909);
xnor U3988 (N_3988,N_1678,N_1627);
xnor U3989 (N_3989,N_2606,N_2698);
nand U3990 (N_3990,N_2210,N_1629);
or U3991 (N_3991,N_1595,N_2548);
and U3992 (N_3992,N_2177,N_1862);
xor U3993 (N_3993,N_2399,N_1577);
and U3994 (N_3994,N_2370,N_1703);
or U3995 (N_3995,N_1872,N_2512);
nor U3996 (N_3996,N_1646,N_1798);
nand U3997 (N_3997,N_2876,N_2427);
xor U3998 (N_3998,N_1501,N_2984);
and U3999 (N_3999,N_2921,N_2843);
nand U4000 (N_4000,N_2237,N_2514);
and U4001 (N_4001,N_2309,N_2285);
xor U4002 (N_4002,N_1745,N_1917);
nor U4003 (N_4003,N_2813,N_2715);
or U4004 (N_4004,N_2237,N_2698);
and U4005 (N_4005,N_2714,N_2356);
nand U4006 (N_4006,N_1688,N_1720);
or U4007 (N_4007,N_1959,N_1612);
nand U4008 (N_4008,N_2760,N_2514);
nor U4009 (N_4009,N_1787,N_2735);
or U4010 (N_4010,N_2728,N_2131);
and U4011 (N_4011,N_1593,N_2269);
nand U4012 (N_4012,N_2501,N_2657);
nor U4013 (N_4013,N_1591,N_2126);
nor U4014 (N_4014,N_2665,N_2489);
nand U4015 (N_4015,N_2542,N_1546);
or U4016 (N_4016,N_1925,N_2570);
xor U4017 (N_4017,N_1612,N_2469);
or U4018 (N_4018,N_2047,N_1693);
nor U4019 (N_4019,N_1576,N_1721);
nand U4020 (N_4020,N_2687,N_2650);
nor U4021 (N_4021,N_2665,N_2031);
nor U4022 (N_4022,N_2463,N_1772);
and U4023 (N_4023,N_2103,N_1690);
or U4024 (N_4024,N_2299,N_2638);
or U4025 (N_4025,N_2451,N_1766);
xor U4026 (N_4026,N_2766,N_2380);
nor U4027 (N_4027,N_1685,N_2794);
and U4028 (N_4028,N_2387,N_1526);
nor U4029 (N_4029,N_1771,N_2792);
nand U4030 (N_4030,N_1990,N_2881);
and U4031 (N_4031,N_2366,N_2088);
or U4032 (N_4032,N_2630,N_2565);
or U4033 (N_4033,N_1502,N_1573);
nand U4034 (N_4034,N_1891,N_1783);
xor U4035 (N_4035,N_1972,N_2378);
xnor U4036 (N_4036,N_2048,N_2629);
xnor U4037 (N_4037,N_2951,N_2756);
nand U4038 (N_4038,N_1948,N_2122);
and U4039 (N_4039,N_2274,N_2170);
or U4040 (N_4040,N_2106,N_2113);
or U4041 (N_4041,N_2420,N_2556);
nand U4042 (N_4042,N_1973,N_2253);
or U4043 (N_4043,N_2533,N_2111);
nand U4044 (N_4044,N_1723,N_2174);
nor U4045 (N_4045,N_2944,N_1560);
and U4046 (N_4046,N_2556,N_2462);
or U4047 (N_4047,N_1636,N_2787);
nor U4048 (N_4048,N_1793,N_2908);
nor U4049 (N_4049,N_1644,N_1700);
nand U4050 (N_4050,N_2860,N_2541);
or U4051 (N_4051,N_1636,N_1581);
and U4052 (N_4052,N_1549,N_1683);
or U4053 (N_4053,N_2001,N_1750);
or U4054 (N_4054,N_1690,N_2094);
nand U4055 (N_4055,N_1542,N_1970);
xor U4056 (N_4056,N_1851,N_2667);
nand U4057 (N_4057,N_2402,N_1621);
and U4058 (N_4058,N_1638,N_2295);
and U4059 (N_4059,N_1514,N_2769);
xor U4060 (N_4060,N_1712,N_2826);
nand U4061 (N_4061,N_2614,N_2684);
or U4062 (N_4062,N_1855,N_2324);
xnor U4063 (N_4063,N_2898,N_2579);
nor U4064 (N_4064,N_1586,N_2251);
or U4065 (N_4065,N_2687,N_2601);
nor U4066 (N_4066,N_2487,N_2951);
nor U4067 (N_4067,N_2259,N_2407);
and U4068 (N_4068,N_2026,N_2048);
xor U4069 (N_4069,N_1598,N_2992);
nor U4070 (N_4070,N_2407,N_2524);
nand U4071 (N_4071,N_1988,N_2473);
nor U4072 (N_4072,N_2610,N_2066);
and U4073 (N_4073,N_2775,N_2671);
and U4074 (N_4074,N_1922,N_2551);
nand U4075 (N_4075,N_1866,N_2880);
xor U4076 (N_4076,N_2372,N_1923);
xor U4077 (N_4077,N_1620,N_2397);
nand U4078 (N_4078,N_2922,N_2576);
nor U4079 (N_4079,N_1831,N_1512);
and U4080 (N_4080,N_2998,N_2940);
nor U4081 (N_4081,N_1565,N_1855);
or U4082 (N_4082,N_2721,N_1745);
and U4083 (N_4083,N_1872,N_2572);
and U4084 (N_4084,N_1905,N_2135);
nand U4085 (N_4085,N_2259,N_2191);
or U4086 (N_4086,N_2918,N_1626);
or U4087 (N_4087,N_2153,N_2662);
xor U4088 (N_4088,N_2167,N_2507);
or U4089 (N_4089,N_2036,N_2045);
xor U4090 (N_4090,N_1505,N_1544);
or U4091 (N_4091,N_2456,N_2778);
xnor U4092 (N_4092,N_1591,N_2044);
or U4093 (N_4093,N_2584,N_1529);
or U4094 (N_4094,N_1510,N_2920);
and U4095 (N_4095,N_1936,N_2863);
xor U4096 (N_4096,N_1588,N_2044);
nor U4097 (N_4097,N_2625,N_2586);
nor U4098 (N_4098,N_2892,N_2731);
or U4099 (N_4099,N_2908,N_2072);
nor U4100 (N_4100,N_2596,N_2771);
nand U4101 (N_4101,N_2415,N_2435);
or U4102 (N_4102,N_1946,N_2262);
and U4103 (N_4103,N_2617,N_2390);
xor U4104 (N_4104,N_2812,N_2377);
nand U4105 (N_4105,N_2009,N_2449);
and U4106 (N_4106,N_2767,N_2645);
xor U4107 (N_4107,N_2308,N_1755);
nor U4108 (N_4108,N_2424,N_1989);
and U4109 (N_4109,N_2918,N_1903);
and U4110 (N_4110,N_1674,N_2039);
or U4111 (N_4111,N_2544,N_2998);
nand U4112 (N_4112,N_1831,N_2352);
and U4113 (N_4113,N_2816,N_2296);
nor U4114 (N_4114,N_2925,N_2597);
xnor U4115 (N_4115,N_2621,N_1947);
nand U4116 (N_4116,N_2663,N_1766);
or U4117 (N_4117,N_1560,N_1665);
xor U4118 (N_4118,N_2568,N_2070);
or U4119 (N_4119,N_2331,N_2793);
nand U4120 (N_4120,N_2475,N_2380);
nand U4121 (N_4121,N_2347,N_2408);
xnor U4122 (N_4122,N_1916,N_2047);
nor U4123 (N_4123,N_1990,N_2488);
and U4124 (N_4124,N_2180,N_1515);
or U4125 (N_4125,N_1924,N_1927);
nand U4126 (N_4126,N_1763,N_2616);
nor U4127 (N_4127,N_2348,N_2109);
nor U4128 (N_4128,N_2062,N_2298);
and U4129 (N_4129,N_2429,N_1547);
nor U4130 (N_4130,N_2227,N_2110);
xnor U4131 (N_4131,N_2103,N_2661);
nand U4132 (N_4132,N_2805,N_2878);
xor U4133 (N_4133,N_2931,N_1508);
and U4134 (N_4134,N_1689,N_2913);
and U4135 (N_4135,N_2248,N_2500);
and U4136 (N_4136,N_2093,N_2848);
and U4137 (N_4137,N_2879,N_2090);
nor U4138 (N_4138,N_1746,N_2297);
and U4139 (N_4139,N_2201,N_2687);
nor U4140 (N_4140,N_2750,N_2870);
nand U4141 (N_4141,N_2058,N_1610);
or U4142 (N_4142,N_2327,N_2847);
or U4143 (N_4143,N_2652,N_2854);
nand U4144 (N_4144,N_1824,N_2348);
xnor U4145 (N_4145,N_1914,N_2432);
and U4146 (N_4146,N_2231,N_1699);
and U4147 (N_4147,N_2071,N_1853);
or U4148 (N_4148,N_2778,N_2375);
nand U4149 (N_4149,N_1851,N_2337);
nand U4150 (N_4150,N_2653,N_2848);
xor U4151 (N_4151,N_1870,N_1545);
xor U4152 (N_4152,N_1773,N_2150);
or U4153 (N_4153,N_2467,N_2126);
nand U4154 (N_4154,N_2316,N_1836);
nor U4155 (N_4155,N_1939,N_2420);
xnor U4156 (N_4156,N_1618,N_2883);
and U4157 (N_4157,N_2516,N_1674);
xnor U4158 (N_4158,N_2679,N_2017);
or U4159 (N_4159,N_2894,N_2623);
nor U4160 (N_4160,N_1942,N_2421);
or U4161 (N_4161,N_2070,N_2796);
or U4162 (N_4162,N_2738,N_1568);
nand U4163 (N_4163,N_2437,N_1567);
nand U4164 (N_4164,N_2053,N_2139);
or U4165 (N_4165,N_2561,N_1691);
nor U4166 (N_4166,N_2823,N_2557);
nor U4167 (N_4167,N_2457,N_1714);
nand U4168 (N_4168,N_2218,N_2624);
xor U4169 (N_4169,N_2493,N_1525);
nand U4170 (N_4170,N_2646,N_1990);
and U4171 (N_4171,N_2671,N_2217);
nor U4172 (N_4172,N_2342,N_1831);
nor U4173 (N_4173,N_1526,N_2012);
or U4174 (N_4174,N_1653,N_2937);
nand U4175 (N_4175,N_2123,N_1527);
xor U4176 (N_4176,N_1557,N_2834);
nor U4177 (N_4177,N_2271,N_1739);
xnor U4178 (N_4178,N_2814,N_2964);
nand U4179 (N_4179,N_2692,N_2315);
xor U4180 (N_4180,N_1765,N_2080);
nand U4181 (N_4181,N_2617,N_1702);
xor U4182 (N_4182,N_2342,N_2617);
nand U4183 (N_4183,N_1690,N_2883);
xnor U4184 (N_4184,N_2401,N_2367);
nor U4185 (N_4185,N_2136,N_2938);
xor U4186 (N_4186,N_1842,N_2077);
and U4187 (N_4187,N_2837,N_1881);
nand U4188 (N_4188,N_2296,N_2592);
or U4189 (N_4189,N_2280,N_1578);
or U4190 (N_4190,N_1804,N_2164);
xnor U4191 (N_4191,N_1862,N_1661);
xor U4192 (N_4192,N_2950,N_2030);
xor U4193 (N_4193,N_2618,N_2849);
or U4194 (N_4194,N_1855,N_2597);
nand U4195 (N_4195,N_2755,N_2432);
nand U4196 (N_4196,N_2005,N_2196);
nand U4197 (N_4197,N_2447,N_2883);
xnor U4198 (N_4198,N_1771,N_2048);
xnor U4199 (N_4199,N_2915,N_2994);
or U4200 (N_4200,N_1750,N_2969);
xor U4201 (N_4201,N_1692,N_2855);
xor U4202 (N_4202,N_1647,N_1940);
or U4203 (N_4203,N_2011,N_2074);
nand U4204 (N_4204,N_1811,N_1942);
or U4205 (N_4205,N_2827,N_2589);
xnor U4206 (N_4206,N_2342,N_2221);
and U4207 (N_4207,N_1525,N_2249);
and U4208 (N_4208,N_1578,N_2968);
or U4209 (N_4209,N_2180,N_2106);
nor U4210 (N_4210,N_2854,N_2924);
or U4211 (N_4211,N_1696,N_2649);
xor U4212 (N_4212,N_1806,N_2971);
nand U4213 (N_4213,N_1520,N_1878);
or U4214 (N_4214,N_2546,N_2704);
nor U4215 (N_4215,N_2168,N_2524);
nor U4216 (N_4216,N_1622,N_1961);
xnor U4217 (N_4217,N_2972,N_1956);
or U4218 (N_4218,N_2406,N_2315);
nand U4219 (N_4219,N_1880,N_2064);
nand U4220 (N_4220,N_1701,N_1706);
nand U4221 (N_4221,N_2515,N_2196);
nor U4222 (N_4222,N_2285,N_2322);
xnor U4223 (N_4223,N_2897,N_2281);
or U4224 (N_4224,N_2965,N_2132);
xor U4225 (N_4225,N_1858,N_2597);
or U4226 (N_4226,N_2629,N_1522);
xnor U4227 (N_4227,N_2917,N_1550);
and U4228 (N_4228,N_1603,N_2845);
or U4229 (N_4229,N_2694,N_2584);
and U4230 (N_4230,N_2167,N_2809);
and U4231 (N_4231,N_2030,N_1617);
nand U4232 (N_4232,N_2812,N_2578);
and U4233 (N_4233,N_2200,N_2088);
nor U4234 (N_4234,N_1590,N_1733);
nand U4235 (N_4235,N_2514,N_1912);
nand U4236 (N_4236,N_2845,N_2800);
nand U4237 (N_4237,N_2080,N_2472);
or U4238 (N_4238,N_1876,N_2542);
nand U4239 (N_4239,N_2860,N_1810);
and U4240 (N_4240,N_2485,N_2853);
nand U4241 (N_4241,N_2642,N_2752);
and U4242 (N_4242,N_1941,N_2392);
nand U4243 (N_4243,N_1919,N_2378);
xnor U4244 (N_4244,N_2371,N_1576);
nor U4245 (N_4245,N_2318,N_2278);
and U4246 (N_4246,N_2885,N_2689);
nand U4247 (N_4247,N_2787,N_2916);
xor U4248 (N_4248,N_2205,N_2561);
or U4249 (N_4249,N_1753,N_1709);
nor U4250 (N_4250,N_2291,N_2072);
and U4251 (N_4251,N_2485,N_2818);
nor U4252 (N_4252,N_2802,N_2151);
nand U4253 (N_4253,N_2240,N_2906);
and U4254 (N_4254,N_2185,N_2440);
or U4255 (N_4255,N_2761,N_1511);
or U4256 (N_4256,N_2370,N_1820);
nand U4257 (N_4257,N_2842,N_2192);
and U4258 (N_4258,N_2112,N_2111);
xnor U4259 (N_4259,N_2794,N_2073);
and U4260 (N_4260,N_1989,N_2187);
xnor U4261 (N_4261,N_2914,N_2978);
and U4262 (N_4262,N_1982,N_1722);
or U4263 (N_4263,N_2221,N_2961);
and U4264 (N_4264,N_2239,N_2084);
or U4265 (N_4265,N_2597,N_2834);
or U4266 (N_4266,N_2360,N_2373);
or U4267 (N_4267,N_2816,N_2186);
nand U4268 (N_4268,N_1637,N_2480);
or U4269 (N_4269,N_2559,N_2476);
nand U4270 (N_4270,N_2395,N_1572);
nand U4271 (N_4271,N_2783,N_2432);
xor U4272 (N_4272,N_1641,N_2339);
nor U4273 (N_4273,N_1843,N_1940);
xor U4274 (N_4274,N_1889,N_1776);
and U4275 (N_4275,N_2106,N_2792);
nor U4276 (N_4276,N_1940,N_1752);
and U4277 (N_4277,N_1746,N_2370);
nand U4278 (N_4278,N_2131,N_1608);
and U4279 (N_4279,N_2497,N_2518);
or U4280 (N_4280,N_2321,N_1848);
nor U4281 (N_4281,N_1745,N_2848);
or U4282 (N_4282,N_2983,N_1621);
xnor U4283 (N_4283,N_2220,N_2147);
nand U4284 (N_4284,N_2451,N_1571);
or U4285 (N_4285,N_2511,N_1995);
nand U4286 (N_4286,N_1977,N_2535);
and U4287 (N_4287,N_2600,N_2082);
xor U4288 (N_4288,N_1944,N_2861);
xnor U4289 (N_4289,N_2078,N_2542);
xor U4290 (N_4290,N_1928,N_2816);
and U4291 (N_4291,N_2969,N_2169);
or U4292 (N_4292,N_2791,N_2809);
xor U4293 (N_4293,N_2771,N_1763);
nand U4294 (N_4294,N_2234,N_1782);
nand U4295 (N_4295,N_1811,N_2340);
nand U4296 (N_4296,N_2576,N_1918);
nor U4297 (N_4297,N_1909,N_2430);
nand U4298 (N_4298,N_2197,N_2807);
xor U4299 (N_4299,N_1746,N_1524);
nor U4300 (N_4300,N_2240,N_2420);
nand U4301 (N_4301,N_2812,N_2079);
nand U4302 (N_4302,N_1645,N_1750);
nand U4303 (N_4303,N_2088,N_2493);
nand U4304 (N_4304,N_2754,N_2958);
and U4305 (N_4305,N_2345,N_2356);
and U4306 (N_4306,N_2275,N_2476);
nor U4307 (N_4307,N_2884,N_2007);
or U4308 (N_4308,N_1810,N_1500);
nand U4309 (N_4309,N_1666,N_1711);
or U4310 (N_4310,N_1636,N_1900);
nor U4311 (N_4311,N_1518,N_2860);
and U4312 (N_4312,N_2068,N_2759);
xnor U4313 (N_4313,N_2291,N_1532);
and U4314 (N_4314,N_1601,N_2304);
nand U4315 (N_4315,N_2023,N_2743);
or U4316 (N_4316,N_2229,N_2122);
or U4317 (N_4317,N_1762,N_2526);
or U4318 (N_4318,N_2905,N_1938);
nand U4319 (N_4319,N_1615,N_2969);
and U4320 (N_4320,N_2442,N_1771);
xor U4321 (N_4321,N_2164,N_2454);
nor U4322 (N_4322,N_2358,N_1612);
nand U4323 (N_4323,N_2330,N_2169);
and U4324 (N_4324,N_2996,N_1853);
xnor U4325 (N_4325,N_1742,N_2224);
and U4326 (N_4326,N_2962,N_2277);
or U4327 (N_4327,N_1505,N_2705);
and U4328 (N_4328,N_1679,N_2653);
xnor U4329 (N_4329,N_2149,N_2464);
nor U4330 (N_4330,N_1802,N_1664);
and U4331 (N_4331,N_2479,N_1573);
or U4332 (N_4332,N_2303,N_2123);
xnor U4333 (N_4333,N_2236,N_2802);
and U4334 (N_4334,N_2607,N_2287);
xor U4335 (N_4335,N_1877,N_2022);
or U4336 (N_4336,N_1591,N_1509);
nand U4337 (N_4337,N_1990,N_2194);
and U4338 (N_4338,N_2343,N_2279);
nand U4339 (N_4339,N_2811,N_2985);
and U4340 (N_4340,N_1830,N_2502);
or U4341 (N_4341,N_2461,N_1755);
nand U4342 (N_4342,N_2541,N_1953);
and U4343 (N_4343,N_2720,N_2926);
xnor U4344 (N_4344,N_2773,N_2480);
nand U4345 (N_4345,N_2097,N_1703);
nand U4346 (N_4346,N_2645,N_2509);
and U4347 (N_4347,N_1816,N_2638);
and U4348 (N_4348,N_2080,N_2208);
and U4349 (N_4349,N_2806,N_2930);
and U4350 (N_4350,N_1586,N_2065);
nor U4351 (N_4351,N_2016,N_2362);
nand U4352 (N_4352,N_1555,N_2917);
nand U4353 (N_4353,N_2563,N_1858);
or U4354 (N_4354,N_2997,N_2861);
and U4355 (N_4355,N_2135,N_2571);
xor U4356 (N_4356,N_2616,N_2277);
or U4357 (N_4357,N_2848,N_2384);
xor U4358 (N_4358,N_2008,N_2916);
nand U4359 (N_4359,N_2829,N_1732);
or U4360 (N_4360,N_2398,N_2409);
and U4361 (N_4361,N_2885,N_2789);
nor U4362 (N_4362,N_1689,N_2324);
nand U4363 (N_4363,N_2502,N_2261);
xor U4364 (N_4364,N_1500,N_2596);
or U4365 (N_4365,N_2196,N_2338);
nor U4366 (N_4366,N_1877,N_1890);
and U4367 (N_4367,N_1989,N_2945);
or U4368 (N_4368,N_1700,N_2443);
or U4369 (N_4369,N_2954,N_2138);
nor U4370 (N_4370,N_1517,N_1972);
and U4371 (N_4371,N_1589,N_1559);
and U4372 (N_4372,N_2870,N_2286);
nand U4373 (N_4373,N_2903,N_2288);
nand U4374 (N_4374,N_2940,N_2108);
and U4375 (N_4375,N_1704,N_1964);
nor U4376 (N_4376,N_1830,N_2536);
xnor U4377 (N_4377,N_2467,N_2725);
nor U4378 (N_4378,N_2446,N_1936);
xnor U4379 (N_4379,N_2870,N_2669);
and U4380 (N_4380,N_2665,N_1602);
nand U4381 (N_4381,N_1787,N_2563);
nor U4382 (N_4382,N_2819,N_2931);
or U4383 (N_4383,N_1579,N_2178);
nand U4384 (N_4384,N_2930,N_1670);
nor U4385 (N_4385,N_2134,N_2756);
and U4386 (N_4386,N_2705,N_2944);
nand U4387 (N_4387,N_1543,N_2117);
xnor U4388 (N_4388,N_2504,N_2697);
xnor U4389 (N_4389,N_2679,N_2640);
nor U4390 (N_4390,N_1650,N_1683);
or U4391 (N_4391,N_2821,N_2001);
xor U4392 (N_4392,N_2489,N_2988);
and U4393 (N_4393,N_2535,N_2420);
xor U4394 (N_4394,N_2341,N_2804);
and U4395 (N_4395,N_1520,N_2239);
and U4396 (N_4396,N_2481,N_2292);
nor U4397 (N_4397,N_2110,N_2898);
or U4398 (N_4398,N_2690,N_1792);
nand U4399 (N_4399,N_1616,N_2854);
or U4400 (N_4400,N_2440,N_2147);
nor U4401 (N_4401,N_2577,N_2409);
and U4402 (N_4402,N_2049,N_2034);
nand U4403 (N_4403,N_2472,N_2487);
nor U4404 (N_4404,N_2444,N_1731);
xor U4405 (N_4405,N_2275,N_2650);
or U4406 (N_4406,N_2757,N_2870);
xor U4407 (N_4407,N_1739,N_2441);
nor U4408 (N_4408,N_1861,N_1501);
or U4409 (N_4409,N_2352,N_2127);
and U4410 (N_4410,N_2755,N_2157);
or U4411 (N_4411,N_2505,N_2235);
nand U4412 (N_4412,N_2563,N_1988);
xnor U4413 (N_4413,N_2310,N_2708);
and U4414 (N_4414,N_2272,N_1633);
xnor U4415 (N_4415,N_2254,N_2798);
and U4416 (N_4416,N_1805,N_1532);
nor U4417 (N_4417,N_2483,N_2861);
or U4418 (N_4418,N_2278,N_1534);
nand U4419 (N_4419,N_2456,N_2737);
xor U4420 (N_4420,N_1866,N_2294);
nor U4421 (N_4421,N_2495,N_1964);
nor U4422 (N_4422,N_2572,N_1662);
or U4423 (N_4423,N_2773,N_1543);
nor U4424 (N_4424,N_2271,N_2831);
or U4425 (N_4425,N_1980,N_2823);
or U4426 (N_4426,N_2449,N_2872);
nor U4427 (N_4427,N_1857,N_1689);
and U4428 (N_4428,N_1795,N_2551);
and U4429 (N_4429,N_1855,N_2231);
and U4430 (N_4430,N_2926,N_2532);
xnor U4431 (N_4431,N_2122,N_1925);
nand U4432 (N_4432,N_2000,N_1781);
or U4433 (N_4433,N_2099,N_1962);
nand U4434 (N_4434,N_2081,N_2510);
nor U4435 (N_4435,N_2588,N_1929);
nand U4436 (N_4436,N_1546,N_2206);
nor U4437 (N_4437,N_2148,N_2884);
or U4438 (N_4438,N_2913,N_2176);
nand U4439 (N_4439,N_2489,N_1929);
xor U4440 (N_4440,N_2867,N_1557);
or U4441 (N_4441,N_2862,N_2268);
xnor U4442 (N_4442,N_2583,N_1569);
nor U4443 (N_4443,N_2150,N_1935);
or U4444 (N_4444,N_1948,N_1572);
nand U4445 (N_4445,N_2276,N_2202);
xor U4446 (N_4446,N_1736,N_1754);
xor U4447 (N_4447,N_2398,N_2895);
or U4448 (N_4448,N_2037,N_1545);
and U4449 (N_4449,N_1532,N_1969);
and U4450 (N_4450,N_1697,N_1572);
and U4451 (N_4451,N_2304,N_1632);
nand U4452 (N_4452,N_1673,N_2397);
and U4453 (N_4453,N_2500,N_2902);
xor U4454 (N_4454,N_1559,N_2193);
nor U4455 (N_4455,N_1991,N_2112);
nor U4456 (N_4456,N_2400,N_1873);
or U4457 (N_4457,N_2293,N_1844);
xnor U4458 (N_4458,N_2025,N_2391);
nand U4459 (N_4459,N_2880,N_1677);
and U4460 (N_4460,N_1564,N_1879);
xor U4461 (N_4461,N_2604,N_2511);
xnor U4462 (N_4462,N_1519,N_1718);
xor U4463 (N_4463,N_2993,N_1647);
or U4464 (N_4464,N_2277,N_2409);
or U4465 (N_4465,N_1512,N_1832);
nor U4466 (N_4466,N_2316,N_1917);
nor U4467 (N_4467,N_2378,N_1838);
xnor U4468 (N_4468,N_1991,N_2411);
nand U4469 (N_4469,N_1545,N_2599);
xnor U4470 (N_4470,N_2731,N_1736);
nor U4471 (N_4471,N_1729,N_1611);
and U4472 (N_4472,N_1834,N_2097);
xnor U4473 (N_4473,N_2627,N_1655);
xnor U4474 (N_4474,N_2966,N_2004);
or U4475 (N_4475,N_2329,N_1536);
and U4476 (N_4476,N_1634,N_2276);
or U4477 (N_4477,N_2568,N_1960);
xnor U4478 (N_4478,N_1716,N_2612);
nor U4479 (N_4479,N_1800,N_1852);
nand U4480 (N_4480,N_1795,N_2068);
or U4481 (N_4481,N_1915,N_2458);
nor U4482 (N_4482,N_2367,N_2394);
nor U4483 (N_4483,N_2065,N_2867);
or U4484 (N_4484,N_1804,N_2351);
nor U4485 (N_4485,N_2229,N_2963);
nor U4486 (N_4486,N_2483,N_1708);
and U4487 (N_4487,N_2330,N_2703);
and U4488 (N_4488,N_2504,N_1748);
or U4489 (N_4489,N_2277,N_2235);
and U4490 (N_4490,N_2764,N_2459);
nand U4491 (N_4491,N_2578,N_2620);
nand U4492 (N_4492,N_1936,N_1934);
xnor U4493 (N_4493,N_1503,N_2324);
nor U4494 (N_4494,N_2576,N_1618);
nor U4495 (N_4495,N_2479,N_2758);
or U4496 (N_4496,N_1992,N_2968);
or U4497 (N_4497,N_1805,N_2347);
nand U4498 (N_4498,N_2497,N_2009);
or U4499 (N_4499,N_2363,N_2690);
xor U4500 (N_4500,N_3059,N_3646);
or U4501 (N_4501,N_3835,N_3204);
and U4502 (N_4502,N_4062,N_4267);
nor U4503 (N_4503,N_4346,N_4171);
nand U4504 (N_4504,N_4169,N_4233);
and U4505 (N_4505,N_3298,N_4475);
nor U4506 (N_4506,N_4286,N_4210);
nand U4507 (N_4507,N_3378,N_3147);
nor U4508 (N_4508,N_3719,N_4178);
xor U4509 (N_4509,N_3413,N_3087);
and U4510 (N_4510,N_4389,N_4331);
or U4511 (N_4511,N_4419,N_4111);
nand U4512 (N_4512,N_4247,N_4032);
nor U4513 (N_4513,N_4318,N_3911);
nor U4514 (N_4514,N_4234,N_3616);
xnor U4515 (N_4515,N_3258,N_4118);
nand U4516 (N_4516,N_4329,N_3385);
nor U4517 (N_4517,N_4063,N_3034);
and U4518 (N_4518,N_3778,N_3342);
nand U4519 (N_4519,N_4205,N_3815);
nand U4520 (N_4520,N_4020,N_4220);
xnor U4521 (N_4521,N_3964,N_3484);
nand U4522 (N_4522,N_4039,N_3775);
nor U4523 (N_4523,N_4384,N_3628);
nand U4524 (N_4524,N_3264,N_4117);
or U4525 (N_4525,N_3965,N_3121);
or U4526 (N_4526,N_3518,N_3916);
and U4527 (N_4527,N_3821,N_3467);
or U4528 (N_4528,N_4291,N_3115);
or U4529 (N_4529,N_3324,N_3767);
nor U4530 (N_4530,N_3496,N_4338);
or U4531 (N_4531,N_4200,N_3590);
and U4532 (N_4532,N_4036,N_3272);
nand U4533 (N_4533,N_3527,N_3520);
and U4534 (N_4534,N_3002,N_3776);
and U4535 (N_4535,N_3302,N_3828);
nand U4536 (N_4536,N_3555,N_3049);
xnor U4537 (N_4537,N_3470,N_3572);
or U4538 (N_4538,N_3387,N_3625);
nand U4539 (N_4539,N_4482,N_3933);
nor U4540 (N_4540,N_4236,N_3399);
nand U4541 (N_4541,N_4315,N_3037);
nor U4542 (N_4542,N_4383,N_3439);
and U4543 (N_4543,N_3537,N_4115);
xnor U4544 (N_4544,N_4425,N_3605);
nand U4545 (N_4545,N_3357,N_4268);
nand U4546 (N_4546,N_3603,N_3630);
nor U4547 (N_4547,N_3794,N_3089);
nand U4548 (N_4548,N_3065,N_4175);
nand U4549 (N_4549,N_3744,N_3491);
nand U4550 (N_4550,N_3701,N_3149);
and U4551 (N_4551,N_3931,N_4430);
xnor U4552 (N_4552,N_4015,N_3807);
xor U4553 (N_4553,N_3909,N_4370);
and U4554 (N_4554,N_3203,N_3486);
and U4555 (N_4555,N_4487,N_4124);
or U4556 (N_4556,N_3596,N_3266);
or U4557 (N_4557,N_3959,N_3655);
nand U4558 (N_4558,N_4305,N_4161);
or U4559 (N_4559,N_4104,N_3384);
nor U4560 (N_4560,N_3528,N_3732);
or U4561 (N_4561,N_3019,N_4049);
or U4562 (N_4562,N_4293,N_3440);
xor U4563 (N_4563,N_3245,N_3741);
nor U4564 (N_4564,N_3417,N_4427);
nand U4565 (N_4565,N_3010,N_4477);
xor U4566 (N_4566,N_3394,N_4071);
or U4567 (N_4567,N_3305,N_3313);
and U4568 (N_4568,N_4086,N_3334);
nor U4569 (N_4569,N_4326,N_3610);
nor U4570 (N_4570,N_4493,N_4371);
and U4571 (N_4571,N_3820,N_4146);
and U4572 (N_4572,N_3762,N_3722);
and U4573 (N_4573,N_4136,N_3580);
or U4574 (N_4574,N_4185,N_3934);
xnor U4575 (N_4575,N_4335,N_4177);
or U4576 (N_4576,N_4040,N_3338);
nand U4577 (N_4577,N_3045,N_3388);
or U4578 (N_4578,N_3228,N_3671);
xor U4579 (N_4579,N_4344,N_3866);
nor U4580 (N_4580,N_3371,N_4140);
xor U4581 (N_4581,N_3550,N_3173);
or U4582 (N_4582,N_3903,N_3875);
xnor U4583 (N_4583,N_4271,N_4207);
nand U4584 (N_4584,N_3494,N_3764);
or U4585 (N_4585,N_3252,N_3057);
and U4586 (N_4586,N_3006,N_3485);
or U4587 (N_4587,N_3030,N_3914);
and U4588 (N_4588,N_3627,N_3178);
and U4589 (N_4589,N_3641,N_3531);
or U4590 (N_4590,N_3919,N_3957);
and U4591 (N_4591,N_4466,N_3084);
xnor U4592 (N_4592,N_4021,N_3459);
and U4593 (N_4593,N_4273,N_4188);
xor U4594 (N_4594,N_3466,N_3331);
or U4595 (N_4595,N_3564,N_4376);
xor U4596 (N_4596,N_3237,N_3380);
nor U4597 (N_4597,N_4393,N_3111);
nand U4598 (N_4598,N_3644,N_4284);
and U4599 (N_4599,N_4102,N_3851);
and U4600 (N_4600,N_4132,N_3005);
xor U4601 (N_4601,N_3329,N_3020);
or U4602 (N_4602,N_3151,N_3437);
or U4603 (N_4603,N_3569,N_4302);
xor U4604 (N_4604,N_3672,N_3800);
nor U4605 (N_4605,N_3805,N_3694);
or U4606 (N_4606,N_3139,N_3219);
or U4607 (N_4607,N_4098,N_4467);
and U4608 (N_4608,N_3543,N_3103);
xnor U4609 (N_4609,N_4292,N_3392);
and U4610 (N_4610,N_3478,N_4099);
nand U4611 (N_4611,N_3925,N_3436);
nand U4612 (N_4612,N_4238,N_3735);
xor U4613 (N_4613,N_4130,N_3664);
nand U4614 (N_4614,N_3231,N_3877);
and U4615 (N_4615,N_4208,N_3487);
and U4616 (N_4616,N_4151,N_4013);
nand U4617 (N_4617,N_3122,N_3373);
or U4618 (N_4618,N_3765,N_3573);
nand U4619 (N_4619,N_3066,N_4119);
nand U4620 (N_4620,N_4141,N_3637);
xor U4621 (N_4621,N_3984,N_3678);
nand U4622 (N_4622,N_3215,N_3830);
nor U4623 (N_4623,N_4415,N_3771);
xor U4624 (N_4624,N_3202,N_3445);
and U4625 (N_4625,N_4374,N_3495);
or U4626 (N_4626,N_3987,N_4100);
and U4627 (N_4627,N_3442,N_3364);
nor U4628 (N_4628,N_3966,N_3177);
nor U4629 (N_4629,N_3856,N_3014);
or U4630 (N_4630,N_3663,N_3094);
and U4631 (N_4631,N_4321,N_4327);
and U4632 (N_4632,N_3554,N_4155);
nand U4633 (N_4633,N_4033,N_3549);
and U4634 (N_4634,N_3426,N_4193);
or U4635 (N_4635,N_3067,N_4088);
and U4636 (N_4636,N_4385,N_3904);
and U4637 (N_4637,N_3736,N_3761);
nor U4638 (N_4638,N_3235,N_3985);
and U4639 (N_4639,N_3261,N_3262);
and U4640 (N_4640,N_4229,N_3015);
or U4641 (N_4641,N_4281,N_3248);
nand U4642 (N_4642,N_4087,N_4241);
or U4643 (N_4643,N_4157,N_3451);
nor U4644 (N_4644,N_3568,N_3662);
nor U4645 (N_4645,N_4164,N_4445);
or U4646 (N_4646,N_3697,N_4495);
nor U4647 (N_4647,N_3131,N_3656);
nor U4648 (N_4648,N_3434,N_3839);
xor U4649 (N_4649,N_4413,N_3758);
nand U4650 (N_4650,N_3503,N_3499);
xor U4651 (N_4651,N_3941,N_3414);
or U4652 (N_4652,N_3947,N_3801);
xnor U4653 (N_4653,N_4257,N_3213);
or U4654 (N_4654,N_4070,N_3396);
nand U4655 (N_4655,N_3687,N_4462);
and U4656 (N_4656,N_3353,N_3469);
nor U4657 (N_4657,N_4242,N_3926);
nor U4658 (N_4658,N_4492,N_3560);
nor U4659 (N_4659,N_4019,N_3383);
nand U4660 (N_4660,N_4282,N_4198);
or U4661 (N_4661,N_3932,N_3593);
xor U4662 (N_4662,N_3545,N_3337);
xor U4663 (N_4663,N_3688,N_4323);
nor U4664 (N_4664,N_4187,N_3563);
and U4665 (N_4665,N_3330,N_4008);
xnor U4666 (N_4666,N_3120,N_3567);
nor U4667 (N_4667,N_4226,N_3128);
or U4668 (N_4668,N_3176,N_4011);
nor U4669 (N_4669,N_3074,N_3477);
and U4670 (N_4670,N_4190,N_3927);
and U4671 (N_4671,N_4397,N_3127);
nor U4672 (N_4672,N_4219,N_4322);
nor U4673 (N_4673,N_3431,N_3157);
and U4674 (N_4674,N_3083,N_3158);
or U4675 (N_4675,N_3649,N_3544);
or U4676 (N_4676,N_3058,N_3136);
xor U4677 (N_4677,N_3635,N_4172);
xor U4678 (N_4678,N_3940,N_3556);
and U4679 (N_4679,N_4356,N_3462);
nand U4680 (N_4680,N_3530,N_3297);
or U4681 (N_4681,N_3670,N_4084);
nor U4682 (N_4682,N_4095,N_3675);
or U4683 (N_4683,N_3340,N_3869);
or U4684 (N_4684,N_3042,N_4288);
nor U4685 (N_4685,N_3939,N_3133);
nor U4686 (N_4686,N_3779,N_3513);
nor U4687 (N_4687,N_3977,N_3367);
xor U4688 (N_4688,N_3587,N_4189);
and U4689 (N_4689,N_4368,N_3063);
and U4690 (N_4690,N_4054,N_3416);
nor U4691 (N_4691,N_3422,N_3016);
and U4692 (N_4692,N_3347,N_3910);
nor U4693 (N_4693,N_4264,N_3638);
nand U4694 (N_4694,N_4074,N_3608);
and U4695 (N_4695,N_3355,N_4114);
or U4696 (N_4696,N_3757,N_3197);
xor U4697 (N_4697,N_4160,N_3474);
nand U4698 (N_4698,N_3225,N_4352);
and U4699 (N_4699,N_3915,N_3583);
or U4700 (N_4700,N_3449,N_3277);
and U4701 (N_4701,N_4283,N_3892);
or U4702 (N_4702,N_4191,N_3328);
nand U4703 (N_4703,N_3960,N_3994);
xor U4704 (N_4704,N_4379,N_3379);
and U4705 (N_4705,N_3168,N_3322);
xor U4706 (N_4706,N_3706,N_4142);
and U4707 (N_4707,N_3148,N_4348);
or U4708 (N_4708,N_3541,N_3222);
and U4709 (N_4709,N_3551,N_4166);
nand U4710 (N_4710,N_4481,N_4307);
nand U4711 (N_4711,N_3818,N_4162);
and U4712 (N_4712,N_3288,N_4259);
xor U4713 (N_4713,N_3134,N_3260);
or U4714 (N_4714,N_4459,N_4055);
nand U4715 (N_4715,N_4051,N_3398);
nor U4716 (N_4716,N_3665,N_3185);
xor U4717 (N_4717,N_3812,N_3946);
and U4718 (N_4718,N_3035,N_4277);
or U4719 (N_4719,N_4382,N_3497);
nor U4720 (N_4720,N_4429,N_3810);
xor U4721 (N_4721,N_3412,N_4025);
nor U4722 (N_4722,N_4306,N_4056);
nand U4723 (N_4723,N_3244,N_4250);
nand U4724 (N_4724,N_3232,N_3923);
nor U4725 (N_4725,N_4176,N_4460);
xnor U4726 (N_4726,N_4399,N_3300);
and U4727 (N_4727,N_4245,N_4248);
nand U4728 (N_4728,N_3553,N_4464);
nand U4729 (N_4729,N_3924,N_3429);
or U4730 (N_4730,N_3072,N_3375);
and U4731 (N_4731,N_4333,N_4408);
xor U4732 (N_4732,N_3184,N_4002);
and U4733 (N_4733,N_3001,N_3256);
or U4734 (N_4734,N_3898,N_4167);
or U4735 (N_4735,N_3286,N_3634);
xor U4736 (N_4736,N_3377,N_3409);
and U4737 (N_4737,N_4499,N_3418);
and U4738 (N_4738,N_3629,N_4061);
nor U4739 (N_4739,N_3243,N_4005);
nor U4740 (N_4740,N_3315,N_3636);
nor U4741 (N_4741,N_3376,N_4228);
and U4742 (N_4742,N_3463,N_3310);
and U4743 (N_4743,N_4422,N_3425);
nand U4744 (N_4744,N_3335,N_3850);
or U4745 (N_4745,N_4179,N_3492);
nand U4746 (N_4746,N_3408,N_3404);
and U4747 (N_4747,N_3796,N_4443);
nand U4748 (N_4748,N_3673,N_3669);
nor U4749 (N_4749,N_3220,N_4361);
nand U4750 (N_4750,N_3088,N_3109);
nor U4751 (N_4751,N_4266,N_3196);
xor U4752 (N_4752,N_3716,N_3770);
and U4753 (N_4753,N_4375,N_3565);
or U4754 (N_4754,N_3129,N_4123);
nand U4755 (N_4755,N_3181,N_4249);
nor U4756 (N_4756,N_3751,N_4411);
xnor U4757 (N_4757,N_3318,N_3025);
xor U4758 (N_4758,N_3705,N_3652);
nor U4759 (N_4759,N_4280,N_3291);
nor U4760 (N_4760,N_3435,N_3532);
and U4761 (N_4761,N_3709,N_3427);
and U4762 (N_4762,N_4078,N_4022);
nand U4763 (N_4763,N_4092,N_3276);
xor U4764 (N_4764,N_4449,N_3843);
or U4765 (N_4765,N_3073,N_3577);
xnor U4766 (N_4766,N_3684,N_3117);
nand U4767 (N_4767,N_3996,N_4437);
nor U4768 (N_4768,N_4034,N_4143);
nor U4769 (N_4769,N_3842,N_3658);
xor U4770 (N_4770,N_3054,N_4096);
nor U4771 (N_4771,N_3853,N_3715);
nor U4772 (N_4772,N_3033,N_3165);
xor U4773 (N_4773,N_3112,N_4439);
xnor U4774 (N_4774,N_3356,N_3717);
or U4775 (N_4775,N_4479,N_4334);
xor U4776 (N_4776,N_4094,N_4258);
nor U4777 (N_4777,N_4209,N_3677);
nand U4778 (N_4778,N_4440,N_3113);
xor U4779 (N_4779,N_3078,N_3983);
or U4780 (N_4780,N_4369,N_4287);
and U4781 (N_4781,N_4030,N_3874);
and U4782 (N_4782,N_3246,N_3359);
and U4783 (N_4783,N_3743,N_3132);
and U4784 (N_4784,N_3858,N_3453);
or U4785 (N_4785,N_3692,N_3990);
and U4786 (N_4786,N_3540,N_3723);
and U4787 (N_4787,N_3118,N_4451);
and U4788 (N_4788,N_3742,N_4418);
or U4789 (N_4789,N_4478,N_3703);
and U4790 (N_4790,N_3847,N_3031);
or U4791 (N_4791,N_3609,N_3949);
and U4792 (N_4792,N_4065,N_3902);
nor U4793 (N_4793,N_4426,N_4497);
nand U4794 (N_4794,N_3307,N_3547);
nand U4795 (N_4795,N_3861,N_3979);
and U4796 (N_4796,N_3681,N_4239);
nand U4797 (N_4797,N_3040,N_3278);
xnor U4798 (N_4798,N_3819,N_3798);
nand U4799 (N_4799,N_3920,N_4489);
nor U4800 (N_4800,N_3490,N_3829);
nor U4801 (N_4801,N_3886,N_3548);
nor U4802 (N_4802,N_4058,N_3750);
nor U4803 (N_4803,N_3639,N_4077);
nand U4804 (N_4804,N_3039,N_3257);
and U4805 (N_4805,N_3802,N_3766);
xnor U4806 (N_4806,N_4355,N_3224);
and U4807 (N_4807,N_4007,N_4103);
nand U4808 (N_4808,N_3082,N_3186);
and U4809 (N_4809,N_3838,N_3622);
or U4810 (N_4810,N_3500,N_3623);
and U4811 (N_4811,N_3461,N_4309);
nand U4812 (N_4812,N_3529,N_3797);
or U4813 (N_4813,N_3188,N_3464);
xor U4814 (N_4814,N_3167,N_3574);
xor U4815 (N_4815,N_3183,N_3854);
and U4816 (N_4816,N_3009,N_3614);
and U4817 (N_4817,N_4133,N_4199);
nand U4818 (N_4818,N_4396,N_3400);
nor U4819 (N_4819,N_3973,N_3522);
or U4820 (N_4820,N_4028,N_4400);
or U4821 (N_4821,N_4488,N_3242);
nand U4822 (N_4822,N_3986,N_3410);
nor U4823 (N_4823,N_4137,N_3195);
and U4824 (N_4824,N_3907,N_3013);
nor U4825 (N_4825,N_3878,N_3607);
nor U4826 (N_4826,N_3651,N_3698);
xnor U4827 (N_4827,N_3411,N_3126);
or U4828 (N_4828,N_4223,N_3621);
or U4829 (N_4829,N_3021,N_4404);
and U4830 (N_4830,N_3963,N_4009);
nor U4831 (N_4831,N_4154,N_3980);
or U4832 (N_4832,N_3788,N_4476);
or U4833 (N_4833,N_4116,N_3227);
xnor U4834 (N_4834,N_3312,N_4206);
and U4835 (N_4835,N_4256,N_4064);
and U4836 (N_4836,N_3104,N_3138);
nor U4837 (N_4837,N_4079,N_3969);
nand U4838 (N_4838,N_4076,N_4173);
nor U4839 (N_4839,N_4147,N_3958);
or U4840 (N_4840,N_3626,N_3552);
or U4841 (N_4841,N_3840,N_3489);
and U4842 (N_4842,N_3504,N_4342);
and U4843 (N_4843,N_3535,N_3036);
nand U4844 (N_4844,N_4278,N_3793);
nand U4845 (N_4845,N_3795,N_4230);
and U4846 (N_4846,N_3817,N_3508);
nor U4847 (N_4847,N_3882,N_4217);
and U4848 (N_4848,N_4004,N_3598);
or U4849 (N_4849,N_3476,N_4276);
nand U4850 (N_4850,N_3447,N_3358);
nor U4851 (N_4851,N_3080,N_4109);
xor U4852 (N_4852,N_4072,N_4203);
nand U4853 (N_4853,N_3233,N_4201);
or U4854 (N_4854,N_3166,N_3424);
nor U4855 (N_4855,N_4269,N_4359);
xnor U4856 (N_4856,N_3632,N_3566);
or U4857 (N_4857,N_3201,N_4153);
xor U4858 (N_4858,N_4456,N_3950);
and U4859 (N_4859,N_4366,N_3473);
nor U4860 (N_4860,N_3061,N_4125);
xor U4861 (N_4861,N_3557,N_3514);
nand U4862 (N_4862,N_4463,N_3296);
nand U4863 (N_4863,N_3003,N_4377);
and U4864 (N_4864,N_3457,N_4149);
nand U4865 (N_4865,N_3441,N_4018);
xnor U4866 (N_4866,N_4044,N_3791);
and U4867 (N_4867,N_4452,N_3119);
nor U4868 (N_4868,N_4290,N_3667);
xnor U4869 (N_4869,N_3206,N_3200);
xnor U4870 (N_4870,N_4252,N_3747);
and U4871 (N_4871,N_4320,N_3279);
nor U4872 (N_4872,N_3975,N_3525);
nand U4873 (N_4873,N_3208,N_3323);
xnor U4874 (N_4874,N_4390,N_4192);
nand U4875 (N_4875,N_4120,N_3785);
or U4876 (N_4876,N_4165,N_4304);
nor U4877 (N_4877,N_3814,N_4373);
or U4878 (N_4878,N_3783,N_3690);
xnor U4879 (N_4879,N_4081,N_4336);
and U4880 (N_4880,N_3017,N_3695);
or U4881 (N_4881,N_3116,N_3606);
xor U4882 (N_4882,N_3961,N_4214);
and U4883 (N_4883,N_4386,N_3571);
or U4884 (N_4884,N_3602,N_4496);
nand U4885 (N_4885,N_4253,N_4353);
or U4886 (N_4886,N_3205,N_3935);
nor U4887 (N_4887,N_3595,N_3407);
and U4888 (N_4888,N_4038,N_4043);
nand U4889 (N_4889,N_3937,N_3406);
xnor U4890 (N_4890,N_3968,N_4244);
nor U4891 (N_4891,N_4423,N_3992);
nor U4892 (N_4892,N_4314,N_3686);
nor U4893 (N_4893,N_3523,N_3238);
or U4894 (N_4894,N_4484,N_4380);
or U4895 (N_4895,N_3189,N_3468);
xor U4896 (N_4896,N_3316,N_3953);
and U4897 (N_4897,N_4184,N_3803);
xor U4898 (N_4898,N_3710,N_3099);
and U4899 (N_4899,N_3075,N_4325);
nor U4900 (N_4900,N_4068,N_3852);
nor U4901 (N_4901,N_3945,N_3153);
xor U4902 (N_4902,N_3198,N_3069);
and U4903 (N_4903,N_4156,N_4026);
or U4904 (N_4904,N_3711,N_3619);
and U4905 (N_4905,N_3633,N_3420);
nand U4906 (N_4906,N_3226,N_3265);
nand U4907 (N_4907,N_4150,N_4468);
xor U4908 (N_4908,N_4204,N_4180);
xor U4909 (N_4909,N_3581,N_3648);
and U4910 (N_4910,N_3870,N_3836);
nor U4911 (N_4911,N_3970,N_3659);
xnor U4912 (N_4912,N_3682,N_3873);
nand U4913 (N_4913,N_3386,N_3570);
and U4914 (N_4914,N_4378,N_3860);
nand U4915 (N_4915,N_3831,N_4135);
or U4916 (N_4916,N_3773,N_4432);
xnor U4917 (N_4917,N_3993,N_3519);
or U4918 (N_4918,N_4388,N_3822);
or U4919 (N_4919,N_3085,N_3050);
nor U4920 (N_4920,N_3594,N_4101);
and U4921 (N_4921,N_3562,N_4406);
and U4922 (N_4922,N_4345,N_3026);
and U4923 (N_4923,N_3576,N_4360);
nor U4924 (N_4924,N_4045,N_3756);
or U4925 (N_4925,N_3921,N_3995);
nand U4926 (N_4926,N_3363,N_4202);
nor U4927 (N_4927,N_3209,N_4006);
nor U4928 (N_4928,N_3871,N_3433);
nand U4929 (N_4929,N_3772,N_3090);
nand U4930 (N_4930,N_4181,N_4299);
nand U4931 (N_4931,N_4225,N_3848);
or U4932 (N_4932,N_3319,N_3381);
nor U4933 (N_4933,N_4480,N_3150);
nor U4934 (N_4934,N_3967,N_3749);
or U4935 (N_4935,N_3917,N_3269);
nor U4936 (N_4936,N_4337,N_3267);
nor U4937 (N_4937,N_3739,N_4295);
nor U4938 (N_4938,N_3865,N_4213);
and U4939 (N_4939,N_4363,N_3056);
nor U4940 (N_4940,N_3509,N_3809);
xor U4941 (N_4941,N_4296,N_3730);
xnor U4942 (N_4942,N_3674,N_3273);
nand U4943 (N_4943,N_4474,N_3391);
and U4944 (N_4944,N_3448,N_3654);
nand U4945 (N_4945,N_3708,N_4401);
and U4946 (N_4946,N_3460,N_3929);
nor U4947 (N_4947,N_4075,N_3981);
and U4948 (N_4948,N_3345,N_3000);
xnor U4949 (N_4949,N_4362,N_4275);
and U4950 (N_4950,N_4319,N_3650);
nor U4951 (N_4951,N_4127,N_3559);
nand U4952 (N_4952,N_4428,N_3022);
or U4953 (N_4953,N_4231,N_3229);
nor U4954 (N_4954,N_3271,N_3214);
nand U4955 (N_4955,N_3901,N_3944);
xnor U4956 (N_4956,N_4126,N_3326);
and U4957 (N_4957,N_3867,N_4148);
or U4958 (N_4958,N_3458,N_3645);
and U4959 (N_4959,N_3734,N_3432);
nand U4960 (N_4960,N_3230,N_4170);
and U4961 (N_4961,N_3752,N_3978);
xor U4962 (N_4962,N_3806,N_3714);
nor U4963 (N_4963,N_3137,N_4131);
xnor U4964 (N_4964,N_4270,N_4310);
xnor U4965 (N_4965,N_3472,N_4372);
or U4966 (N_4966,N_4060,N_3982);
or U4967 (N_4967,N_4186,N_3270);
and U4968 (N_4968,N_3811,N_3780);
or U4969 (N_4969,N_3507,N_3471);
nor U4970 (N_4970,N_3689,N_4196);
nand U4971 (N_4971,N_3423,N_3787);
or U4972 (N_4972,N_3889,N_3790);
xnor U4973 (N_4973,N_4324,N_3539);
or U4974 (N_4974,N_3125,N_4243);
nor U4975 (N_4975,N_3038,N_4024);
or U4976 (N_4976,N_3287,N_3344);
or U4977 (N_4977,N_4235,N_4069);
nand U4978 (N_4978,N_3047,N_3382);
or U4979 (N_4979,N_3169,N_3857);
or U4980 (N_4980,N_3055,N_3465);
and U4981 (N_4981,N_3320,N_3446);
or U4982 (N_4982,N_3912,N_3832);
or U4983 (N_4983,N_3521,N_3533);
or U4984 (N_4984,N_3585,N_3044);
or U4985 (N_4985,N_3180,N_3163);
nor U4986 (N_4986,N_3360,N_4301);
xnor U4987 (N_4987,N_4224,N_3844);
and U4988 (N_4988,N_3100,N_3393);
nand U4989 (N_4989,N_3368,N_4272);
nor U4990 (N_4990,N_3737,N_3728);
nor U4991 (N_4991,N_3612,N_3259);
nor U4992 (N_4992,N_3365,N_4134);
or U4993 (N_4993,N_4097,N_4237);
and U4994 (N_4994,N_4289,N_4082);
xnor U4995 (N_4995,N_3043,N_4365);
or U4996 (N_4996,N_3156,N_3618);
nand U4997 (N_4997,N_3702,N_3754);
xnor U4998 (N_4998,N_3369,N_4311);
xor U4999 (N_4999,N_3299,N_3106);
or U5000 (N_5000,N_3881,N_3295);
nand U5001 (N_5001,N_3403,N_4398);
and U5002 (N_5002,N_3221,N_3501);
xnor U5003 (N_5003,N_4455,N_3223);
and U5004 (N_5004,N_3475,N_3366);
and U5005 (N_5005,N_3845,N_3098);
and U5006 (N_5006,N_4457,N_4139);
nor U5007 (N_5007,N_3479,N_4195);
and U5008 (N_5008,N_3211,N_3162);
xnor U5009 (N_5009,N_4351,N_3913);
or U5010 (N_5010,N_3604,N_4317);
or U5011 (N_5011,N_3588,N_3685);
nor U5012 (N_5012,N_4339,N_3012);
and U5013 (N_5013,N_4222,N_3624);
xor U5014 (N_5014,N_3951,N_4254);
xor U5015 (N_5015,N_3234,N_4387);
and U5016 (N_5016,N_3897,N_4073);
nor U5017 (N_5017,N_3430,N_4357);
nand U5018 (N_5018,N_3782,N_3774);
nand U5019 (N_5019,N_4122,N_3456);
nor U5020 (N_5020,N_3443,N_3175);
xnor U5021 (N_5021,N_4473,N_4444);
xor U5022 (N_5022,N_3046,N_3062);
nor U5023 (N_5023,N_3855,N_3647);
or U5024 (N_5024,N_3304,N_4297);
nand U5025 (N_5025,N_3023,N_4350);
and U5026 (N_5026,N_3834,N_3102);
or U5027 (N_5027,N_3586,N_3141);
xor U5028 (N_5028,N_3640,N_3438);
or U5029 (N_5029,N_4470,N_4498);
xor U5030 (N_5030,N_3859,N_3159);
xor U5031 (N_5031,N_3027,N_3962);
nand U5032 (N_5032,N_4128,N_3918);
xnor U5033 (N_5033,N_4194,N_3361);
nor U5034 (N_5034,N_3395,N_4298);
or U5035 (N_5035,N_3303,N_3160);
and U5036 (N_5036,N_3142,N_4262);
and U5037 (N_5037,N_3051,N_4471);
and U5038 (N_5038,N_3372,N_4340);
or U5039 (N_5039,N_3249,N_3683);
nand U5040 (N_5040,N_3239,N_3505);
nand U5041 (N_5041,N_4145,N_3254);
and U5042 (N_5042,N_4138,N_3879);
xor U5043 (N_5043,N_3140,N_3191);
xor U5044 (N_5044,N_4316,N_3086);
nand U5045 (N_5045,N_3972,N_3534);
and U5046 (N_5046,N_3899,N_4441);
xnor U5047 (N_5047,N_3611,N_3956);
nor U5048 (N_5048,N_3240,N_3110);
nand U5049 (N_5049,N_3064,N_3145);
nand U5050 (N_5050,N_4014,N_3247);
or U5051 (N_5051,N_4197,N_3081);
or U5052 (N_5052,N_4410,N_3642);
xnor U5053 (N_5053,N_3352,N_3155);
or U5054 (N_5054,N_4129,N_4240);
or U5055 (N_5055,N_3253,N_3024);
and U5056 (N_5056,N_4303,N_4436);
nor U5057 (N_5057,N_4080,N_3760);
or U5058 (N_5058,N_3060,N_3280);
xor U5059 (N_5059,N_3582,N_3895);
nand U5060 (N_5060,N_3428,N_4453);
nand U5061 (N_5061,N_3578,N_4108);
or U5062 (N_5062,N_3336,N_4448);
and U5063 (N_5063,N_3643,N_4431);
or U5064 (N_5064,N_3661,N_4472);
nand U5065 (N_5065,N_3693,N_3691);
xnor U5066 (N_5066,N_3070,N_3700);
or U5067 (N_5067,N_4091,N_3498);
or U5068 (N_5068,N_4212,N_3290);
or U5069 (N_5069,N_3011,N_3908);
or U5070 (N_5070,N_3263,N_4001);
nor U5071 (N_5071,N_3350,N_4434);
and U5072 (N_5072,N_4433,N_3346);
xnor U5073 (N_5073,N_3885,N_4261);
or U5074 (N_5074,N_3101,N_3952);
nand U5075 (N_5075,N_4405,N_3193);
nor U5076 (N_5076,N_3668,N_4093);
nor U5077 (N_5077,N_4152,N_3282);
or U5078 (N_5078,N_4435,N_3837);
nand U5079 (N_5079,N_4144,N_3849);
xnor U5080 (N_5080,N_4279,N_3421);
xnor U5081 (N_5081,N_3600,N_4041);
xnor U5082 (N_5082,N_3216,N_4424);
or U5083 (N_5083,N_4059,N_3726);
and U5084 (N_5084,N_3349,N_3405);
nand U5085 (N_5085,N_3283,N_3660);
and U5086 (N_5086,N_3890,N_3444);
and U5087 (N_5087,N_3746,N_3317);
nor U5088 (N_5088,N_4395,N_4227);
and U5089 (N_5089,N_3332,N_3942);
or U5090 (N_5090,N_3351,N_3930);
or U5091 (N_5091,N_4438,N_4182);
xor U5092 (N_5092,N_3592,N_3199);
xor U5093 (N_5093,N_4486,N_3989);
nor U5094 (N_5094,N_3900,N_4332);
and U5095 (N_5095,N_3763,N_3301);
xor U5096 (N_5096,N_3954,N_3928);
and U5097 (N_5097,N_3883,N_3721);
or U5098 (N_5098,N_3402,N_3096);
nor U5099 (N_5099,N_3091,N_3725);
and U5100 (N_5100,N_3187,N_3813);
xor U5101 (N_5101,N_3846,N_4048);
or U5102 (N_5102,N_4046,N_3327);
nor U5103 (N_5103,N_3863,N_3482);
and U5104 (N_5104,N_3631,N_3862);
xnor U5105 (N_5105,N_4367,N_3579);
or U5106 (N_5106,N_4042,N_3888);
nand U5107 (N_5107,N_3450,N_3241);
or U5108 (N_5108,N_4446,N_3348);
or U5109 (N_5109,N_3804,N_3207);
nand U5110 (N_5110,N_3362,N_3620);
xor U5111 (N_5111,N_3008,N_3179);
nand U5112 (N_5112,N_3955,N_3321);
xor U5113 (N_5113,N_4066,N_3792);
xnor U5114 (N_5114,N_4417,N_3905);
xor U5115 (N_5115,N_3731,N_4211);
nand U5116 (N_5116,N_4012,N_4251);
nand U5117 (N_5117,N_3745,N_3354);
or U5118 (N_5118,N_3251,N_3536);
xor U5119 (N_5119,N_4110,N_4000);
or U5120 (N_5120,N_4308,N_3894);
and U5121 (N_5121,N_4494,N_3048);
xor U5122 (N_5122,N_3130,N_3584);
nor U5123 (N_5123,N_3284,N_4246);
and U5124 (N_5124,N_4294,N_3052);
or U5125 (N_5125,N_3841,N_4232);
nor U5126 (N_5126,N_3512,N_3161);
or U5127 (N_5127,N_3210,N_3493);
nand U5128 (N_5128,N_3823,N_3816);
nor U5129 (N_5129,N_3943,N_4358);
xnor U5130 (N_5130,N_3615,N_3676);
or U5131 (N_5131,N_3341,N_4407);
nor U5132 (N_5132,N_3679,N_3007);
xor U5133 (N_5133,N_4416,N_3488);
nor U5134 (N_5134,N_3455,N_3991);
nor U5135 (N_5135,N_3154,N_3517);
or U5136 (N_5136,N_3028,N_3825);
xnor U5137 (N_5137,N_4085,N_3415);
xnor U5138 (N_5138,N_3135,N_3390);
xor U5139 (N_5139,N_3740,N_4031);
nand U5140 (N_5140,N_4260,N_4392);
and U5141 (N_5141,N_3748,N_4330);
xor U5142 (N_5142,N_4454,N_3755);
nor U5143 (N_5143,N_3389,N_3095);
nor U5144 (N_5144,N_3948,N_4053);
nor U5145 (N_5145,N_4215,N_4442);
and U5146 (N_5146,N_4490,N_4414);
nor U5147 (N_5147,N_3561,N_3309);
xnor U5148 (N_5148,N_4067,N_3143);
xor U5149 (N_5149,N_4016,N_4090);
nor U5150 (N_5150,N_4029,N_3076);
or U5151 (N_5151,N_3029,N_3032);
xor U5152 (N_5152,N_4491,N_4313);
and U5153 (N_5153,N_3510,N_3546);
nor U5154 (N_5154,N_4450,N_3506);
xnor U5155 (N_5155,N_3144,N_3194);
xor U5156 (N_5156,N_3053,N_3680);
or U5157 (N_5157,N_3077,N_3733);
and U5158 (N_5158,N_3936,N_3174);
or U5159 (N_5159,N_3452,N_3311);
xnor U5160 (N_5160,N_3777,N_3339);
xor U5161 (N_5161,N_3988,N_3666);
nand U5162 (N_5162,N_3868,N_3454);
xor U5163 (N_5163,N_4465,N_3827);
nand U5164 (N_5164,N_3597,N_3824);
nand U5165 (N_5165,N_3092,N_3876);
and U5166 (N_5166,N_3575,N_3768);
nand U5167 (N_5167,N_4341,N_4159);
or U5168 (N_5168,N_3884,N_3893);
nor U5169 (N_5169,N_3724,N_3502);
and U5170 (N_5170,N_3864,N_3524);
nand U5171 (N_5171,N_3784,N_4403);
or U5172 (N_5172,N_4274,N_3289);
nor U5173 (N_5173,N_3308,N_3123);
and U5174 (N_5174,N_4420,N_3097);
nand U5175 (N_5175,N_3325,N_4158);
and U5176 (N_5176,N_3617,N_3293);
and U5177 (N_5177,N_3192,N_4047);
nand U5178 (N_5178,N_3713,N_3653);
xnor U5179 (N_5179,N_4483,N_4107);
or U5180 (N_5180,N_3880,N_3004);
and U5181 (N_5181,N_3727,N_3707);
nand U5182 (N_5182,N_4381,N_3306);
xnor U5183 (N_5183,N_4255,N_3333);
xor U5184 (N_5184,N_4037,N_3896);
xor U5185 (N_5185,N_3190,N_3974);
nor U5186 (N_5186,N_3170,N_3511);
and U5187 (N_5187,N_4391,N_3294);
and U5188 (N_5188,N_3314,N_3704);
or U5189 (N_5189,N_3526,N_3292);
or U5190 (N_5190,N_4265,N_4050);
xor U5191 (N_5191,N_4023,N_4106);
nand U5192 (N_5192,N_4469,N_4035);
and U5193 (N_5193,N_3997,N_4121);
and U5194 (N_5194,N_4312,N_3938);
xnor U5195 (N_5195,N_4105,N_3599);
xor U5196 (N_5196,N_3872,N_3976);
nand U5197 (N_5197,N_4394,N_4113);
nor U5198 (N_5198,N_3281,N_3601);
and U5199 (N_5199,N_4216,N_3146);
nor U5200 (N_5200,N_4354,N_3999);
and U5201 (N_5201,N_3769,N_3906);
nand U5202 (N_5202,N_3613,N_3107);
nor U5203 (N_5203,N_3480,N_4089);
or U5204 (N_5204,N_3481,N_3789);
and U5205 (N_5205,N_3212,N_3738);
and U5206 (N_5206,N_3538,N_3236);
and U5207 (N_5207,N_3152,N_3079);
or U5208 (N_5208,N_4364,N_4421);
xnor U5209 (N_5209,N_4458,N_3171);
xnor U5210 (N_5210,N_4300,N_3164);
nand U5211 (N_5211,N_3274,N_3419);
nand U5212 (N_5212,N_3887,N_4447);
or U5213 (N_5213,N_3105,N_4349);
and U5214 (N_5214,N_3114,N_4027);
or U5215 (N_5215,N_4168,N_3397);
xor U5216 (N_5216,N_4402,N_3182);
xnor U5217 (N_5217,N_4409,N_3998);
xnor U5218 (N_5218,N_3071,N_4285);
or U5219 (N_5219,N_3591,N_4017);
xnor U5220 (N_5220,N_3018,N_4112);
or U5221 (N_5221,N_3068,N_3250);
and U5222 (N_5222,N_3833,N_4183);
or U5223 (N_5223,N_3799,N_3971);
or U5224 (N_5224,N_4218,N_4003);
xnor U5225 (N_5225,N_4052,N_3699);
xor U5226 (N_5226,N_3275,N_3589);
or U5227 (N_5227,N_3124,N_3922);
or U5228 (N_5228,N_4010,N_3720);
and U5229 (N_5229,N_3657,N_4174);
or U5230 (N_5230,N_3542,N_3753);
nor U5231 (N_5231,N_4343,N_3718);
xor U5232 (N_5232,N_3401,N_3729);
or U5233 (N_5233,N_3786,N_3108);
or U5234 (N_5234,N_3558,N_3041);
xor U5235 (N_5235,N_4221,N_3808);
or U5236 (N_5236,N_4347,N_3712);
and U5237 (N_5237,N_3093,N_3285);
nand U5238 (N_5238,N_3268,N_3370);
xnor U5239 (N_5239,N_3217,N_3759);
or U5240 (N_5240,N_4083,N_4328);
nor U5241 (N_5241,N_4412,N_4057);
nand U5242 (N_5242,N_3515,N_3516);
nand U5243 (N_5243,N_4461,N_3483);
nor U5244 (N_5244,N_4163,N_3696);
nand U5245 (N_5245,N_3891,N_3826);
nand U5246 (N_5246,N_4485,N_3343);
nand U5247 (N_5247,N_4263,N_3172);
or U5248 (N_5248,N_3255,N_3781);
xnor U5249 (N_5249,N_3374,N_3218);
nand U5250 (N_5250,N_3936,N_4409);
nor U5251 (N_5251,N_3902,N_3184);
nor U5252 (N_5252,N_3452,N_3964);
nor U5253 (N_5253,N_4019,N_3940);
or U5254 (N_5254,N_4354,N_3898);
nand U5255 (N_5255,N_4267,N_4431);
and U5256 (N_5256,N_3968,N_3632);
nor U5257 (N_5257,N_3538,N_4240);
nor U5258 (N_5258,N_4108,N_3801);
xnor U5259 (N_5259,N_3085,N_4032);
or U5260 (N_5260,N_3998,N_3837);
or U5261 (N_5261,N_3545,N_3665);
or U5262 (N_5262,N_4322,N_4080);
xnor U5263 (N_5263,N_3552,N_3085);
nor U5264 (N_5264,N_4462,N_3837);
and U5265 (N_5265,N_3247,N_3879);
nand U5266 (N_5266,N_3534,N_3516);
and U5267 (N_5267,N_4188,N_3704);
and U5268 (N_5268,N_3578,N_3515);
and U5269 (N_5269,N_4442,N_3912);
nor U5270 (N_5270,N_3089,N_4385);
nand U5271 (N_5271,N_3379,N_3999);
nor U5272 (N_5272,N_4414,N_3139);
and U5273 (N_5273,N_3349,N_4347);
nor U5274 (N_5274,N_3078,N_4032);
or U5275 (N_5275,N_3196,N_3163);
or U5276 (N_5276,N_3365,N_3502);
nor U5277 (N_5277,N_3434,N_3681);
and U5278 (N_5278,N_3488,N_3685);
or U5279 (N_5279,N_3731,N_3741);
nor U5280 (N_5280,N_3915,N_3385);
nor U5281 (N_5281,N_4246,N_4184);
or U5282 (N_5282,N_3320,N_4447);
or U5283 (N_5283,N_3171,N_4220);
nor U5284 (N_5284,N_4338,N_3254);
nand U5285 (N_5285,N_3785,N_4421);
and U5286 (N_5286,N_3297,N_3720);
nand U5287 (N_5287,N_3167,N_3046);
xnor U5288 (N_5288,N_4123,N_3124);
xor U5289 (N_5289,N_4018,N_3625);
and U5290 (N_5290,N_3649,N_4347);
and U5291 (N_5291,N_3896,N_3585);
and U5292 (N_5292,N_3398,N_4180);
and U5293 (N_5293,N_3862,N_3321);
or U5294 (N_5294,N_3108,N_3467);
nand U5295 (N_5295,N_3035,N_3977);
nor U5296 (N_5296,N_4235,N_4106);
xnor U5297 (N_5297,N_4101,N_3894);
xnor U5298 (N_5298,N_3413,N_4298);
or U5299 (N_5299,N_4276,N_3619);
or U5300 (N_5300,N_3594,N_4431);
nand U5301 (N_5301,N_3833,N_3942);
nor U5302 (N_5302,N_3397,N_3893);
nand U5303 (N_5303,N_3637,N_3421);
or U5304 (N_5304,N_4365,N_3387);
or U5305 (N_5305,N_3216,N_4147);
nor U5306 (N_5306,N_3290,N_3225);
and U5307 (N_5307,N_3798,N_3765);
or U5308 (N_5308,N_3183,N_3317);
nand U5309 (N_5309,N_3633,N_4066);
nand U5310 (N_5310,N_3893,N_3556);
and U5311 (N_5311,N_3726,N_3061);
nand U5312 (N_5312,N_3041,N_4378);
nand U5313 (N_5313,N_3201,N_4233);
or U5314 (N_5314,N_4238,N_4065);
nor U5315 (N_5315,N_3346,N_3311);
xnor U5316 (N_5316,N_3430,N_3418);
nand U5317 (N_5317,N_3428,N_3099);
nor U5318 (N_5318,N_3634,N_3937);
and U5319 (N_5319,N_4134,N_4056);
xor U5320 (N_5320,N_3974,N_3090);
nor U5321 (N_5321,N_3635,N_4295);
and U5322 (N_5322,N_4106,N_4307);
or U5323 (N_5323,N_4119,N_3419);
and U5324 (N_5324,N_3733,N_4088);
or U5325 (N_5325,N_3151,N_4083);
xnor U5326 (N_5326,N_3037,N_3721);
xnor U5327 (N_5327,N_3638,N_4267);
nor U5328 (N_5328,N_3134,N_3624);
nor U5329 (N_5329,N_3869,N_3233);
or U5330 (N_5330,N_3276,N_3480);
nand U5331 (N_5331,N_3152,N_3648);
or U5332 (N_5332,N_3629,N_4379);
xnor U5333 (N_5333,N_4103,N_3869);
nand U5334 (N_5334,N_4053,N_3989);
xnor U5335 (N_5335,N_3065,N_3703);
and U5336 (N_5336,N_3121,N_4292);
or U5337 (N_5337,N_3173,N_3053);
nand U5338 (N_5338,N_3429,N_3831);
xor U5339 (N_5339,N_3502,N_3842);
and U5340 (N_5340,N_3673,N_3836);
and U5341 (N_5341,N_4370,N_3713);
nor U5342 (N_5342,N_3492,N_4010);
nor U5343 (N_5343,N_3440,N_3811);
or U5344 (N_5344,N_3739,N_3207);
nand U5345 (N_5345,N_3322,N_3816);
nand U5346 (N_5346,N_3440,N_3599);
nand U5347 (N_5347,N_4233,N_3144);
nand U5348 (N_5348,N_3792,N_3759);
nand U5349 (N_5349,N_4429,N_3292);
or U5350 (N_5350,N_3162,N_3214);
nor U5351 (N_5351,N_3502,N_3659);
and U5352 (N_5352,N_4189,N_4374);
xor U5353 (N_5353,N_4105,N_3201);
nand U5354 (N_5354,N_3657,N_3159);
and U5355 (N_5355,N_3027,N_3834);
xor U5356 (N_5356,N_4340,N_3216);
or U5357 (N_5357,N_4423,N_3008);
and U5358 (N_5358,N_3745,N_4468);
nand U5359 (N_5359,N_4218,N_4354);
nand U5360 (N_5360,N_4001,N_4038);
and U5361 (N_5361,N_3391,N_4146);
or U5362 (N_5362,N_3511,N_3958);
nor U5363 (N_5363,N_3276,N_3394);
nor U5364 (N_5364,N_4291,N_4495);
xnor U5365 (N_5365,N_3308,N_4140);
and U5366 (N_5366,N_3522,N_4363);
xnor U5367 (N_5367,N_3043,N_3133);
xnor U5368 (N_5368,N_3341,N_3446);
xor U5369 (N_5369,N_3630,N_4323);
nand U5370 (N_5370,N_3152,N_3491);
nand U5371 (N_5371,N_3115,N_3431);
or U5372 (N_5372,N_3554,N_3337);
and U5373 (N_5373,N_3882,N_3838);
nor U5374 (N_5374,N_3367,N_4008);
or U5375 (N_5375,N_3008,N_4203);
xnor U5376 (N_5376,N_4394,N_3612);
nor U5377 (N_5377,N_3102,N_3111);
nor U5378 (N_5378,N_3268,N_3637);
and U5379 (N_5379,N_4022,N_3316);
or U5380 (N_5380,N_3917,N_3988);
nand U5381 (N_5381,N_3575,N_3548);
or U5382 (N_5382,N_4209,N_3331);
nand U5383 (N_5383,N_3691,N_3086);
nand U5384 (N_5384,N_3114,N_3055);
nand U5385 (N_5385,N_3091,N_4129);
nor U5386 (N_5386,N_4220,N_3180);
or U5387 (N_5387,N_3969,N_3931);
nand U5388 (N_5388,N_3497,N_3081);
and U5389 (N_5389,N_3196,N_3692);
xnor U5390 (N_5390,N_3690,N_3568);
or U5391 (N_5391,N_3266,N_3153);
or U5392 (N_5392,N_3486,N_3835);
nand U5393 (N_5393,N_3199,N_3663);
and U5394 (N_5394,N_3547,N_4090);
xnor U5395 (N_5395,N_3622,N_3823);
and U5396 (N_5396,N_3475,N_3026);
nand U5397 (N_5397,N_4484,N_3866);
and U5398 (N_5398,N_4093,N_3490);
nand U5399 (N_5399,N_3142,N_3438);
or U5400 (N_5400,N_4441,N_3977);
nand U5401 (N_5401,N_3863,N_3332);
and U5402 (N_5402,N_3599,N_4314);
nor U5403 (N_5403,N_3227,N_4357);
nand U5404 (N_5404,N_3980,N_4092);
and U5405 (N_5405,N_3241,N_3529);
and U5406 (N_5406,N_3669,N_3265);
xor U5407 (N_5407,N_3740,N_4158);
or U5408 (N_5408,N_3180,N_3124);
nand U5409 (N_5409,N_3260,N_3774);
xor U5410 (N_5410,N_4427,N_3839);
nand U5411 (N_5411,N_3476,N_3859);
nand U5412 (N_5412,N_3072,N_3565);
nor U5413 (N_5413,N_3473,N_3785);
nor U5414 (N_5414,N_4422,N_4363);
xor U5415 (N_5415,N_3590,N_3710);
xor U5416 (N_5416,N_4252,N_3284);
or U5417 (N_5417,N_4102,N_3147);
nor U5418 (N_5418,N_4005,N_4015);
nor U5419 (N_5419,N_3723,N_3611);
nor U5420 (N_5420,N_3577,N_4151);
or U5421 (N_5421,N_3822,N_3985);
xnor U5422 (N_5422,N_3433,N_3867);
xnor U5423 (N_5423,N_3643,N_3758);
nand U5424 (N_5424,N_3127,N_3578);
or U5425 (N_5425,N_3734,N_4007);
nand U5426 (N_5426,N_3543,N_3624);
or U5427 (N_5427,N_3035,N_3903);
and U5428 (N_5428,N_3536,N_4426);
xnor U5429 (N_5429,N_3181,N_4267);
nor U5430 (N_5430,N_3986,N_3279);
xor U5431 (N_5431,N_3754,N_3600);
or U5432 (N_5432,N_3712,N_4117);
and U5433 (N_5433,N_3584,N_4092);
nor U5434 (N_5434,N_4399,N_3586);
nor U5435 (N_5435,N_3742,N_3940);
and U5436 (N_5436,N_3623,N_3187);
or U5437 (N_5437,N_3839,N_3907);
nand U5438 (N_5438,N_3534,N_4478);
or U5439 (N_5439,N_3120,N_3149);
and U5440 (N_5440,N_3779,N_4389);
xnor U5441 (N_5441,N_3467,N_4172);
xor U5442 (N_5442,N_3113,N_3634);
xor U5443 (N_5443,N_4075,N_3764);
nand U5444 (N_5444,N_3692,N_4266);
xor U5445 (N_5445,N_3294,N_4427);
nor U5446 (N_5446,N_4451,N_3247);
nor U5447 (N_5447,N_4236,N_3400);
and U5448 (N_5448,N_3996,N_4226);
or U5449 (N_5449,N_3737,N_3536);
and U5450 (N_5450,N_3122,N_4326);
nand U5451 (N_5451,N_3581,N_3449);
nor U5452 (N_5452,N_3083,N_3190);
and U5453 (N_5453,N_3749,N_3897);
nor U5454 (N_5454,N_3224,N_3965);
nand U5455 (N_5455,N_4255,N_3181);
or U5456 (N_5456,N_3346,N_4299);
and U5457 (N_5457,N_3352,N_3471);
and U5458 (N_5458,N_4241,N_4061);
and U5459 (N_5459,N_4246,N_3447);
nor U5460 (N_5460,N_3093,N_4248);
and U5461 (N_5461,N_4036,N_4059);
nand U5462 (N_5462,N_3696,N_3561);
nand U5463 (N_5463,N_3734,N_3206);
or U5464 (N_5464,N_4234,N_3471);
and U5465 (N_5465,N_3063,N_4331);
nand U5466 (N_5466,N_4474,N_3577);
nor U5467 (N_5467,N_4164,N_4184);
nor U5468 (N_5468,N_3317,N_3574);
xor U5469 (N_5469,N_3571,N_3505);
and U5470 (N_5470,N_3599,N_3521);
or U5471 (N_5471,N_3074,N_3783);
or U5472 (N_5472,N_4265,N_4250);
or U5473 (N_5473,N_3995,N_3962);
and U5474 (N_5474,N_4495,N_3127);
or U5475 (N_5475,N_4449,N_3978);
nor U5476 (N_5476,N_3900,N_3343);
and U5477 (N_5477,N_4257,N_3104);
nor U5478 (N_5478,N_3025,N_3917);
nand U5479 (N_5479,N_4121,N_4222);
and U5480 (N_5480,N_3543,N_3374);
and U5481 (N_5481,N_3964,N_3702);
xor U5482 (N_5482,N_4008,N_3072);
nor U5483 (N_5483,N_4356,N_4446);
xor U5484 (N_5484,N_3050,N_4459);
xor U5485 (N_5485,N_4047,N_4213);
or U5486 (N_5486,N_3265,N_3036);
or U5487 (N_5487,N_4241,N_4178);
xnor U5488 (N_5488,N_3332,N_3182);
nor U5489 (N_5489,N_3625,N_4148);
xor U5490 (N_5490,N_3127,N_4183);
xor U5491 (N_5491,N_3365,N_3185);
nand U5492 (N_5492,N_3195,N_4001);
nand U5493 (N_5493,N_4171,N_3789);
nor U5494 (N_5494,N_3985,N_3366);
and U5495 (N_5495,N_3859,N_4037);
nor U5496 (N_5496,N_3613,N_3170);
xor U5497 (N_5497,N_3535,N_4099);
nor U5498 (N_5498,N_3750,N_3565);
nand U5499 (N_5499,N_3795,N_3502);
or U5500 (N_5500,N_3826,N_3661);
nor U5501 (N_5501,N_3167,N_3594);
xor U5502 (N_5502,N_4474,N_3769);
nor U5503 (N_5503,N_3564,N_3909);
nand U5504 (N_5504,N_3060,N_3189);
and U5505 (N_5505,N_3418,N_3382);
and U5506 (N_5506,N_3784,N_3041);
xor U5507 (N_5507,N_3388,N_3122);
nand U5508 (N_5508,N_3532,N_4081);
xor U5509 (N_5509,N_3493,N_3790);
or U5510 (N_5510,N_4017,N_3295);
and U5511 (N_5511,N_4394,N_3764);
xnor U5512 (N_5512,N_3148,N_4223);
nand U5513 (N_5513,N_3605,N_4193);
nor U5514 (N_5514,N_4269,N_3497);
xnor U5515 (N_5515,N_3870,N_3212);
xnor U5516 (N_5516,N_4125,N_3774);
nand U5517 (N_5517,N_4478,N_3345);
xor U5518 (N_5518,N_3736,N_4223);
xnor U5519 (N_5519,N_3937,N_3785);
and U5520 (N_5520,N_3821,N_3501);
and U5521 (N_5521,N_3299,N_3149);
and U5522 (N_5522,N_4167,N_3220);
xnor U5523 (N_5523,N_4315,N_4452);
xnor U5524 (N_5524,N_3039,N_3288);
nand U5525 (N_5525,N_4298,N_4216);
or U5526 (N_5526,N_3274,N_3300);
xnor U5527 (N_5527,N_3322,N_3998);
nand U5528 (N_5528,N_4098,N_3544);
xor U5529 (N_5529,N_4123,N_4191);
xor U5530 (N_5530,N_3055,N_3860);
or U5531 (N_5531,N_4115,N_3277);
or U5532 (N_5532,N_3874,N_4392);
xor U5533 (N_5533,N_4479,N_3572);
and U5534 (N_5534,N_3381,N_3814);
nand U5535 (N_5535,N_4010,N_3131);
and U5536 (N_5536,N_3412,N_3925);
nor U5537 (N_5537,N_4061,N_3036);
and U5538 (N_5538,N_3837,N_3092);
xnor U5539 (N_5539,N_3957,N_3103);
or U5540 (N_5540,N_3542,N_3935);
nor U5541 (N_5541,N_4129,N_3970);
xnor U5542 (N_5542,N_3960,N_3787);
or U5543 (N_5543,N_3028,N_3953);
nand U5544 (N_5544,N_4120,N_3950);
xor U5545 (N_5545,N_3052,N_3696);
or U5546 (N_5546,N_4413,N_3162);
and U5547 (N_5547,N_4434,N_3497);
and U5548 (N_5548,N_4385,N_4089);
nand U5549 (N_5549,N_3346,N_3970);
and U5550 (N_5550,N_3754,N_3418);
or U5551 (N_5551,N_4412,N_4354);
nor U5552 (N_5552,N_4172,N_3047);
nor U5553 (N_5553,N_4073,N_3667);
or U5554 (N_5554,N_3270,N_3864);
or U5555 (N_5555,N_3286,N_3192);
nor U5556 (N_5556,N_4071,N_3316);
xnor U5557 (N_5557,N_3151,N_4299);
or U5558 (N_5558,N_4012,N_3253);
nor U5559 (N_5559,N_3062,N_3380);
nor U5560 (N_5560,N_3084,N_4446);
nor U5561 (N_5561,N_4403,N_3673);
nor U5562 (N_5562,N_3817,N_3446);
and U5563 (N_5563,N_3916,N_3888);
nor U5564 (N_5564,N_3302,N_4397);
nand U5565 (N_5565,N_3261,N_4051);
nor U5566 (N_5566,N_3540,N_4246);
xnor U5567 (N_5567,N_3682,N_3673);
xor U5568 (N_5568,N_3623,N_3720);
or U5569 (N_5569,N_3070,N_3928);
nor U5570 (N_5570,N_3176,N_4235);
nor U5571 (N_5571,N_3665,N_3600);
xor U5572 (N_5572,N_3817,N_3411);
or U5573 (N_5573,N_3657,N_3276);
xnor U5574 (N_5574,N_4195,N_3191);
and U5575 (N_5575,N_3910,N_3469);
nand U5576 (N_5576,N_3043,N_4129);
nand U5577 (N_5577,N_4412,N_3167);
nor U5578 (N_5578,N_3206,N_3573);
nand U5579 (N_5579,N_3398,N_3561);
and U5580 (N_5580,N_3522,N_3927);
nand U5581 (N_5581,N_4029,N_3639);
nand U5582 (N_5582,N_3662,N_3234);
xor U5583 (N_5583,N_3316,N_4010);
or U5584 (N_5584,N_3011,N_3722);
and U5585 (N_5585,N_3090,N_4376);
or U5586 (N_5586,N_3511,N_3259);
nor U5587 (N_5587,N_3221,N_3197);
xor U5588 (N_5588,N_3567,N_4416);
nor U5589 (N_5589,N_4366,N_4079);
nor U5590 (N_5590,N_3437,N_3744);
nand U5591 (N_5591,N_3175,N_3345);
nand U5592 (N_5592,N_3405,N_3824);
or U5593 (N_5593,N_3254,N_3616);
nor U5594 (N_5594,N_3093,N_4355);
and U5595 (N_5595,N_3374,N_3076);
nor U5596 (N_5596,N_4094,N_4291);
nor U5597 (N_5597,N_3084,N_4390);
or U5598 (N_5598,N_3140,N_3980);
nor U5599 (N_5599,N_3868,N_4068);
xnor U5600 (N_5600,N_3632,N_4153);
or U5601 (N_5601,N_4443,N_3061);
nand U5602 (N_5602,N_4213,N_3451);
nand U5603 (N_5603,N_4195,N_3293);
and U5604 (N_5604,N_3350,N_3753);
nand U5605 (N_5605,N_4197,N_4188);
xnor U5606 (N_5606,N_3182,N_4207);
nor U5607 (N_5607,N_4241,N_4234);
or U5608 (N_5608,N_3988,N_3307);
xnor U5609 (N_5609,N_3971,N_4042);
and U5610 (N_5610,N_3179,N_3535);
or U5611 (N_5611,N_4111,N_4339);
nand U5612 (N_5612,N_4225,N_3438);
and U5613 (N_5613,N_4034,N_4001);
and U5614 (N_5614,N_3246,N_3545);
or U5615 (N_5615,N_4037,N_4382);
or U5616 (N_5616,N_4230,N_3188);
and U5617 (N_5617,N_3173,N_4202);
and U5618 (N_5618,N_3005,N_3741);
or U5619 (N_5619,N_3497,N_4043);
nand U5620 (N_5620,N_3944,N_4386);
xor U5621 (N_5621,N_4197,N_3982);
xnor U5622 (N_5622,N_3093,N_4104);
or U5623 (N_5623,N_4449,N_3378);
nand U5624 (N_5624,N_3398,N_3736);
nand U5625 (N_5625,N_4197,N_4450);
or U5626 (N_5626,N_4468,N_3502);
and U5627 (N_5627,N_4289,N_3983);
or U5628 (N_5628,N_3561,N_3444);
nand U5629 (N_5629,N_3417,N_3573);
nor U5630 (N_5630,N_3401,N_4289);
nor U5631 (N_5631,N_3979,N_3157);
and U5632 (N_5632,N_3107,N_3048);
nand U5633 (N_5633,N_3400,N_4032);
or U5634 (N_5634,N_3817,N_3445);
and U5635 (N_5635,N_4231,N_3071);
or U5636 (N_5636,N_3914,N_3729);
nor U5637 (N_5637,N_4314,N_4082);
xor U5638 (N_5638,N_3278,N_4464);
xnor U5639 (N_5639,N_4097,N_3115);
nor U5640 (N_5640,N_4444,N_4335);
xor U5641 (N_5641,N_4047,N_3426);
and U5642 (N_5642,N_3766,N_4079);
nor U5643 (N_5643,N_3184,N_4315);
nor U5644 (N_5644,N_4164,N_4317);
nor U5645 (N_5645,N_3731,N_4343);
and U5646 (N_5646,N_3800,N_3727);
xnor U5647 (N_5647,N_3197,N_3884);
or U5648 (N_5648,N_3806,N_3740);
nand U5649 (N_5649,N_3206,N_3744);
and U5650 (N_5650,N_3848,N_3956);
and U5651 (N_5651,N_3656,N_3468);
xor U5652 (N_5652,N_4333,N_4116);
and U5653 (N_5653,N_4385,N_3310);
xnor U5654 (N_5654,N_3792,N_3580);
and U5655 (N_5655,N_3770,N_4038);
xor U5656 (N_5656,N_3583,N_3251);
or U5657 (N_5657,N_4399,N_3963);
or U5658 (N_5658,N_3067,N_4097);
nor U5659 (N_5659,N_4466,N_4379);
and U5660 (N_5660,N_3237,N_4098);
nor U5661 (N_5661,N_3922,N_3446);
xor U5662 (N_5662,N_3639,N_3330);
or U5663 (N_5663,N_3052,N_3012);
nor U5664 (N_5664,N_3470,N_4261);
nand U5665 (N_5665,N_3735,N_3750);
nand U5666 (N_5666,N_3993,N_3419);
nor U5667 (N_5667,N_3518,N_3432);
nor U5668 (N_5668,N_3795,N_3126);
nor U5669 (N_5669,N_4280,N_3248);
nand U5670 (N_5670,N_3358,N_4121);
nor U5671 (N_5671,N_4368,N_4173);
and U5672 (N_5672,N_4180,N_3125);
xnor U5673 (N_5673,N_3866,N_3158);
xor U5674 (N_5674,N_3000,N_4031);
nand U5675 (N_5675,N_3555,N_4441);
or U5676 (N_5676,N_3510,N_4217);
nor U5677 (N_5677,N_3819,N_3257);
xnor U5678 (N_5678,N_4490,N_4454);
xor U5679 (N_5679,N_3867,N_4035);
xnor U5680 (N_5680,N_3405,N_3311);
and U5681 (N_5681,N_4105,N_3191);
nand U5682 (N_5682,N_4442,N_3974);
and U5683 (N_5683,N_3768,N_3917);
xnor U5684 (N_5684,N_3436,N_3861);
and U5685 (N_5685,N_3644,N_4285);
nand U5686 (N_5686,N_3302,N_4176);
and U5687 (N_5687,N_3605,N_4103);
xnor U5688 (N_5688,N_3757,N_3735);
nand U5689 (N_5689,N_3685,N_3781);
nor U5690 (N_5690,N_3164,N_3435);
xnor U5691 (N_5691,N_4293,N_3076);
and U5692 (N_5692,N_4249,N_3313);
or U5693 (N_5693,N_3440,N_3945);
nand U5694 (N_5694,N_3837,N_3186);
xnor U5695 (N_5695,N_3106,N_3752);
and U5696 (N_5696,N_3290,N_3965);
nand U5697 (N_5697,N_3307,N_4028);
nand U5698 (N_5698,N_3206,N_4159);
xnor U5699 (N_5699,N_3353,N_3672);
or U5700 (N_5700,N_3382,N_4475);
and U5701 (N_5701,N_3486,N_3601);
or U5702 (N_5702,N_4188,N_4267);
xnor U5703 (N_5703,N_3260,N_3462);
nor U5704 (N_5704,N_4040,N_3096);
xor U5705 (N_5705,N_4172,N_4399);
nand U5706 (N_5706,N_4453,N_3954);
and U5707 (N_5707,N_4101,N_4385);
or U5708 (N_5708,N_3547,N_3371);
nor U5709 (N_5709,N_4146,N_3989);
nand U5710 (N_5710,N_3038,N_4314);
or U5711 (N_5711,N_3481,N_3690);
and U5712 (N_5712,N_4089,N_4363);
nor U5713 (N_5713,N_4148,N_3327);
or U5714 (N_5714,N_3521,N_3054);
or U5715 (N_5715,N_3903,N_3793);
xnor U5716 (N_5716,N_3212,N_4243);
nor U5717 (N_5717,N_3216,N_4016);
and U5718 (N_5718,N_3517,N_3540);
nand U5719 (N_5719,N_3400,N_3790);
xnor U5720 (N_5720,N_3093,N_3458);
nor U5721 (N_5721,N_4284,N_4340);
or U5722 (N_5722,N_3323,N_3228);
xor U5723 (N_5723,N_3161,N_4368);
or U5724 (N_5724,N_3429,N_4240);
nand U5725 (N_5725,N_3575,N_3417);
nand U5726 (N_5726,N_3218,N_4237);
nor U5727 (N_5727,N_4476,N_3823);
nor U5728 (N_5728,N_4210,N_3417);
nand U5729 (N_5729,N_3659,N_3716);
or U5730 (N_5730,N_3399,N_3330);
or U5731 (N_5731,N_4288,N_4433);
nor U5732 (N_5732,N_3370,N_3651);
and U5733 (N_5733,N_3452,N_3739);
xor U5734 (N_5734,N_4084,N_4222);
nor U5735 (N_5735,N_4163,N_4400);
nor U5736 (N_5736,N_3632,N_3132);
or U5737 (N_5737,N_3824,N_3498);
or U5738 (N_5738,N_3741,N_3063);
or U5739 (N_5739,N_3629,N_3624);
or U5740 (N_5740,N_3227,N_3640);
or U5741 (N_5741,N_3824,N_3908);
nand U5742 (N_5742,N_4281,N_3829);
and U5743 (N_5743,N_3792,N_3431);
nand U5744 (N_5744,N_3060,N_3125);
or U5745 (N_5745,N_4088,N_3878);
and U5746 (N_5746,N_4083,N_4226);
and U5747 (N_5747,N_3962,N_3219);
or U5748 (N_5748,N_4065,N_3780);
nand U5749 (N_5749,N_3031,N_3005);
and U5750 (N_5750,N_3918,N_3247);
and U5751 (N_5751,N_3106,N_4152);
or U5752 (N_5752,N_4139,N_4455);
xnor U5753 (N_5753,N_4397,N_4319);
nand U5754 (N_5754,N_4354,N_4224);
nand U5755 (N_5755,N_3517,N_4401);
nand U5756 (N_5756,N_3713,N_3903);
nor U5757 (N_5757,N_4352,N_4357);
or U5758 (N_5758,N_3389,N_3519);
and U5759 (N_5759,N_3520,N_3086);
and U5760 (N_5760,N_3777,N_4480);
nor U5761 (N_5761,N_4131,N_4136);
xnor U5762 (N_5762,N_3602,N_3484);
nand U5763 (N_5763,N_3421,N_3564);
xnor U5764 (N_5764,N_4359,N_3842);
or U5765 (N_5765,N_4283,N_4133);
xor U5766 (N_5766,N_3874,N_3242);
xor U5767 (N_5767,N_4173,N_4391);
nand U5768 (N_5768,N_4349,N_3245);
nor U5769 (N_5769,N_3133,N_3993);
nor U5770 (N_5770,N_3295,N_3320);
or U5771 (N_5771,N_3311,N_3073);
xor U5772 (N_5772,N_4299,N_3311);
or U5773 (N_5773,N_4147,N_3228);
nand U5774 (N_5774,N_3951,N_3097);
xor U5775 (N_5775,N_3052,N_3583);
xnor U5776 (N_5776,N_3541,N_3773);
or U5777 (N_5777,N_3884,N_3828);
xor U5778 (N_5778,N_4308,N_3970);
nor U5779 (N_5779,N_3903,N_4145);
xor U5780 (N_5780,N_4363,N_4270);
or U5781 (N_5781,N_4449,N_4096);
or U5782 (N_5782,N_3270,N_3777);
nand U5783 (N_5783,N_3435,N_4387);
and U5784 (N_5784,N_3316,N_3237);
nor U5785 (N_5785,N_3447,N_4124);
and U5786 (N_5786,N_3469,N_3506);
nor U5787 (N_5787,N_4368,N_4074);
nand U5788 (N_5788,N_4452,N_3039);
nand U5789 (N_5789,N_3611,N_4282);
xor U5790 (N_5790,N_4476,N_4081);
or U5791 (N_5791,N_3322,N_3863);
and U5792 (N_5792,N_3696,N_4308);
or U5793 (N_5793,N_3292,N_3985);
nor U5794 (N_5794,N_3339,N_4175);
xnor U5795 (N_5795,N_4318,N_4388);
nand U5796 (N_5796,N_3691,N_3553);
nor U5797 (N_5797,N_3953,N_3158);
or U5798 (N_5798,N_4197,N_3425);
and U5799 (N_5799,N_3780,N_3764);
nand U5800 (N_5800,N_3920,N_3290);
nand U5801 (N_5801,N_4413,N_3602);
or U5802 (N_5802,N_4054,N_3920);
or U5803 (N_5803,N_4419,N_3650);
xnor U5804 (N_5804,N_3542,N_3087);
nand U5805 (N_5805,N_3715,N_4149);
xnor U5806 (N_5806,N_4262,N_3669);
and U5807 (N_5807,N_3308,N_4138);
or U5808 (N_5808,N_3948,N_3316);
or U5809 (N_5809,N_3541,N_3004);
nor U5810 (N_5810,N_4185,N_4195);
xor U5811 (N_5811,N_4242,N_3480);
nand U5812 (N_5812,N_3919,N_3366);
and U5813 (N_5813,N_3709,N_4169);
nor U5814 (N_5814,N_4171,N_4130);
and U5815 (N_5815,N_3822,N_3828);
xnor U5816 (N_5816,N_3724,N_3399);
or U5817 (N_5817,N_4175,N_3982);
or U5818 (N_5818,N_3498,N_4095);
and U5819 (N_5819,N_3573,N_3994);
nor U5820 (N_5820,N_3880,N_4373);
and U5821 (N_5821,N_3926,N_3951);
nand U5822 (N_5822,N_4327,N_4169);
or U5823 (N_5823,N_3714,N_4035);
nor U5824 (N_5824,N_3397,N_4296);
and U5825 (N_5825,N_4409,N_3980);
xnor U5826 (N_5826,N_4136,N_4031);
xor U5827 (N_5827,N_4016,N_3690);
xnor U5828 (N_5828,N_3853,N_3926);
and U5829 (N_5829,N_3845,N_3652);
nand U5830 (N_5830,N_3910,N_3283);
nor U5831 (N_5831,N_3099,N_3235);
and U5832 (N_5832,N_3348,N_4376);
nand U5833 (N_5833,N_4426,N_3514);
or U5834 (N_5834,N_3783,N_3765);
xor U5835 (N_5835,N_3536,N_3157);
and U5836 (N_5836,N_3130,N_4223);
or U5837 (N_5837,N_3262,N_3635);
and U5838 (N_5838,N_3090,N_4437);
nor U5839 (N_5839,N_4224,N_3383);
xnor U5840 (N_5840,N_3136,N_3534);
xor U5841 (N_5841,N_3775,N_4055);
and U5842 (N_5842,N_4454,N_4413);
and U5843 (N_5843,N_3329,N_4066);
nor U5844 (N_5844,N_3912,N_3775);
nand U5845 (N_5845,N_4196,N_3514);
xor U5846 (N_5846,N_3472,N_4119);
xnor U5847 (N_5847,N_4139,N_4134);
or U5848 (N_5848,N_4478,N_4210);
or U5849 (N_5849,N_4470,N_3952);
nand U5850 (N_5850,N_4371,N_4063);
nor U5851 (N_5851,N_3118,N_3558);
or U5852 (N_5852,N_3612,N_3744);
and U5853 (N_5853,N_3021,N_3402);
nand U5854 (N_5854,N_4207,N_3734);
and U5855 (N_5855,N_3042,N_3489);
xnor U5856 (N_5856,N_3420,N_3986);
xor U5857 (N_5857,N_3230,N_4416);
nor U5858 (N_5858,N_4054,N_4271);
or U5859 (N_5859,N_4370,N_3251);
xnor U5860 (N_5860,N_3673,N_3413);
nand U5861 (N_5861,N_3500,N_3301);
or U5862 (N_5862,N_3967,N_3275);
nor U5863 (N_5863,N_4005,N_3220);
nand U5864 (N_5864,N_4155,N_4438);
nand U5865 (N_5865,N_3515,N_4028);
nor U5866 (N_5866,N_4305,N_4478);
or U5867 (N_5867,N_4364,N_4228);
xor U5868 (N_5868,N_3052,N_4454);
xor U5869 (N_5869,N_4445,N_4117);
xor U5870 (N_5870,N_4163,N_4354);
xnor U5871 (N_5871,N_3996,N_3781);
nor U5872 (N_5872,N_4075,N_3946);
nand U5873 (N_5873,N_4451,N_3455);
and U5874 (N_5874,N_4425,N_4423);
xor U5875 (N_5875,N_4362,N_3804);
nor U5876 (N_5876,N_4185,N_3514);
and U5877 (N_5877,N_3798,N_4411);
nand U5878 (N_5878,N_4316,N_3477);
or U5879 (N_5879,N_3317,N_3200);
xnor U5880 (N_5880,N_4291,N_3220);
nor U5881 (N_5881,N_3838,N_3284);
nand U5882 (N_5882,N_4188,N_3139);
nor U5883 (N_5883,N_4368,N_4345);
nand U5884 (N_5884,N_4223,N_3589);
and U5885 (N_5885,N_3166,N_4301);
or U5886 (N_5886,N_3343,N_4271);
nor U5887 (N_5887,N_3843,N_4168);
and U5888 (N_5888,N_3557,N_4381);
nor U5889 (N_5889,N_4279,N_3637);
nor U5890 (N_5890,N_3147,N_3661);
or U5891 (N_5891,N_3778,N_3420);
nor U5892 (N_5892,N_3999,N_3814);
nor U5893 (N_5893,N_3735,N_4457);
and U5894 (N_5894,N_3613,N_3998);
xnor U5895 (N_5895,N_4468,N_3596);
and U5896 (N_5896,N_3489,N_3126);
nor U5897 (N_5897,N_3152,N_3260);
nor U5898 (N_5898,N_3457,N_4061);
xor U5899 (N_5899,N_3950,N_3796);
or U5900 (N_5900,N_3207,N_4055);
nand U5901 (N_5901,N_3068,N_4488);
nor U5902 (N_5902,N_3163,N_3798);
nor U5903 (N_5903,N_3522,N_3248);
nor U5904 (N_5904,N_3860,N_3453);
and U5905 (N_5905,N_3417,N_3477);
xor U5906 (N_5906,N_4049,N_4352);
nor U5907 (N_5907,N_3190,N_3960);
and U5908 (N_5908,N_4083,N_3213);
or U5909 (N_5909,N_3880,N_3164);
or U5910 (N_5910,N_3632,N_3465);
nand U5911 (N_5911,N_3205,N_3505);
and U5912 (N_5912,N_4182,N_3107);
nand U5913 (N_5913,N_3025,N_4319);
xnor U5914 (N_5914,N_4047,N_3302);
nor U5915 (N_5915,N_3336,N_3067);
xor U5916 (N_5916,N_3114,N_3097);
or U5917 (N_5917,N_4018,N_3733);
nor U5918 (N_5918,N_3894,N_3888);
xor U5919 (N_5919,N_3081,N_3411);
xor U5920 (N_5920,N_3861,N_3232);
and U5921 (N_5921,N_3197,N_4437);
nand U5922 (N_5922,N_3604,N_3531);
or U5923 (N_5923,N_3017,N_4281);
and U5924 (N_5924,N_3145,N_3458);
xnor U5925 (N_5925,N_3773,N_3300);
nor U5926 (N_5926,N_3152,N_3107);
nand U5927 (N_5927,N_3335,N_3778);
xnor U5928 (N_5928,N_4342,N_3033);
xnor U5929 (N_5929,N_4414,N_3526);
or U5930 (N_5930,N_3097,N_3504);
nand U5931 (N_5931,N_3656,N_3515);
nor U5932 (N_5932,N_4357,N_3151);
nand U5933 (N_5933,N_3821,N_3022);
nand U5934 (N_5934,N_4237,N_4400);
nand U5935 (N_5935,N_3476,N_3028);
and U5936 (N_5936,N_3803,N_3302);
or U5937 (N_5937,N_4206,N_3490);
and U5938 (N_5938,N_3889,N_3571);
or U5939 (N_5939,N_4188,N_3331);
xnor U5940 (N_5940,N_4452,N_3733);
nand U5941 (N_5941,N_4199,N_3575);
nor U5942 (N_5942,N_4179,N_4168);
or U5943 (N_5943,N_4367,N_4225);
nor U5944 (N_5944,N_3793,N_3114);
and U5945 (N_5945,N_4289,N_3975);
or U5946 (N_5946,N_4163,N_3631);
or U5947 (N_5947,N_3821,N_3635);
and U5948 (N_5948,N_4471,N_3211);
nand U5949 (N_5949,N_3704,N_3229);
or U5950 (N_5950,N_3954,N_3021);
xnor U5951 (N_5951,N_3306,N_4359);
nor U5952 (N_5952,N_3041,N_4157);
and U5953 (N_5953,N_3961,N_3657);
xor U5954 (N_5954,N_4401,N_3382);
nor U5955 (N_5955,N_3401,N_3271);
nand U5956 (N_5956,N_3189,N_4194);
xnor U5957 (N_5957,N_3505,N_3602);
nor U5958 (N_5958,N_4203,N_3739);
nor U5959 (N_5959,N_3829,N_3674);
and U5960 (N_5960,N_4193,N_3595);
xnor U5961 (N_5961,N_3047,N_3166);
or U5962 (N_5962,N_3127,N_3629);
nor U5963 (N_5963,N_3092,N_4481);
xor U5964 (N_5964,N_3294,N_3029);
xnor U5965 (N_5965,N_4300,N_3135);
and U5966 (N_5966,N_3352,N_4174);
nor U5967 (N_5967,N_3518,N_4022);
or U5968 (N_5968,N_3347,N_4245);
nor U5969 (N_5969,N_3125,N_3130);
nor U5970 (N_5970,N_4384,N_3073);
nor U5971 (N_5971,N_3935,N_3922);
xor U5972 (N_5972,N_3553,N_3100);
xnor U5973 (N_5973,N_4488,N_3925);
and U5974 (N_5974,N_3528,N_4216);
or U5975 (N_5975,N_4134,N_3096);
nand U5976 (N_5976,N_3134,N_4371);
or U5977 (N_5977,N_3959,N_3925);
nor U5978 (N_5978,N_3027,N_3680);
nor U5979 (N_5979,N_3755,N_3165);
nor U5980 (N_5980,N_4400,N_4289);
xnor U5981 (N_5981,N_3146,N_3890);
and U5982 (N_5982,N_3919,N_3336);
and U5983 (N_5983,N_4380,N_3270);
nand U5984 (N_5984,N_4083,N_3778);
nand U5985 (N_5985,N_3421,N_4455);
or U5986 (N_5986,N_3958,N_3310);
nand U5987 (N_5987,N_4438,N_3859);
or U5988 (N_5988,N_3943,N_3522);
nor U5989 (N_5989,N_3508,N_3309);
and U5990 (N_5990,N_4382,N_3996);
and U5991 (N_5991,N_3477,N_3128);
or U5992 (N_5992,N_3569,N_3120);
xnor U5993 (N_5993,N_3194,N_3666);
and U5994 (N_5994,N_3239,N_4324);
nor U5995 (N_5995,N_3643,N_3416);
nor U5996 (N_5996,N_4356,N_3648);
nand U5997 (N_5997,N_3024,N_3307);
xor U5998 (N_5998,N_3610,N_3428);
and U5999 (N_5999,N_3857,N_3437);
nand U6000 (N_6000,N_5251,N_5856);
nand U6001 (N_6001,N_5381,N_5294);
and U6002 (N_6002,N_5031,N_4585);
and U6003 (N_6003,N_5175,N_5731);
xnor U6004 (N_6004,N_5901,N_4850);
nand U6005 (N_6005,N_4939,N_5577);
or U6006 (N_6006,N_5763,N_4604);
or U6007 (N_6007,N_5448,N_5487);
nand U6008 (N_6008,N_4896,N_5304);
nor U6009 (N_6009,N_5380,N_5992);
xnor U6010 (N_6010,N_4520,N_5445);
xnor U6011 (N_6011,N_5660,N_4847);
and U6012 (N_6012,N_4812,N_4581);
nor U6013 (N_6013,N_5222,N_4566);
and U6014 (N_6014,N_4725,N_5208);
or U6015 (N_6015,N_5300,N_5833);
and U6016 (N_6016,N_5906,N_4663);
nand U6017 (N_6017,N_5132,N_5422);
and U6018 (N_6018,N_5002,N_5245);
nand U6019 (N_6019,N_4995,N_5799);
nor U6020 (N_6020,N_5198,N_4808);
or U6021 (N_6021,N_5551,N_4719);
nand U6022 (N_6022,N_5729,N_5685);
nand U6023 (N_6023,N_5370,N_5985);
nor U6024 (N_6024,N_5828,N_5835);
or U6025 (N_6025,N_5665,N_4662);
xnor U6026 (N_6026,N_5942,N_5193);
or U6027 (N_6027,N_5421,N_5553);
xor U6028 (N_6028,N_5213,N_5544);
or U6029 (N_6029,N_5368,N_5573);
xor U6030 (N_6030,N_5859,N_5273);
and U6031 (N_6031,N_5152,N_5975);
nor U6032 (N_6032,N_5072,N_4848);
xnor U6033 (N_6033,N_5201,N_4908);
nand U6034 (N_6034,N_5626,N_5686);
nor U6035 (N_6035,N_5321,N_5988);
and U6036 (N_6036,N_4723,N_4676);
nand U6037 (N_6037,N_5816,N_4509);
and U6038 (N_6038,N_5540,N_4521);
and U6039 (N_6039,N_4794,N_5563);
and U6040 (N_6040,N_5558,N_5583);
xnor U6041 (N_6041,N_5654,N_5397);
nand U6042 (N_6042,N_4568,N_5647);
and U6043 (N_6043,N_5025,N_4711);
xor U6044 (N_6044,N_5829,N_5052);
nor U6045 (N_6045,N_4539,N_5036);
xnor U6046 (N_6046,N_5454,N_5821);
xnor U6047 (N_6047,N_4636,N_4641);
nand U6048 (N_6048,N_4682,N_5373);
xor U6049 (N_6049,N_5332,N_4646);
nor U6050 (N_6050,N_4962,N_4635);
or U6051 (N_6051,N_5896,N_4872);
xor U6052 (N_6052,N_5032,N_4658);
and U6053 (N_6053,N_4652,N_4551);
nand U6054 (N_6054,N_4975,N_5240);
nand U6055 (N_6055,N_4846,N_4562);
nor U6056 (N_6056,N_4788,N_4906);
xor U6057 (N_6057,N_4919,N_5225);
and U6058 (N_6058,N_5409,N_5857);
nand U6059 (N_6059,N_5075,N_5008);
and U6060 (N_6060,N_5335,N_5897);
or U6061 (N_6061,N_5314,N_5532);
nor U6062 (N_6062,N_5705,N_5793);
nand U6063 (N_6063,N_5872,N_5131);
nand U6064 (N_6064,N_5268,N_4565);
and U6065 (N_6065,N_5775,N_5139);
nand U6066 (N_6066,N_5186,N_5880);
or U6067 (N_6067,N_4998,N_5642);
nand U6068 (N_6068,N_5952,N_5787);
nand U6069 (N_6069,N_5931,N_5400);
xor U6070 (N_6070,N_5961,N_5166);
nor U6071 (N_6071,N_5475,N_5702);
and U6072 (N_6072,N_5565,N_5112);
nor U6073 (N_6073,N_5029,N_4761);
or U6074 (N_6074,N_4835,N_5840);
nand U6075 (N_6075,N_4598,N_5003);
and U6076 (N_6076,N_5231,N_4976);
nand U6077 (N_6077,N_5493,N_4833);
and U6078 (N_6078,N_5651,N_4513);
nor U6079 (N_6079,N_5452,N_5444);
and U6080 (N_6080,N_4512,N_5734);
and U6081 (N_6081,N_5291,N_5242);
nor U6082 (N_6082,N_5441,N_5679);
and U6083 (N_6083,N_5286,N_4747);
and U6084 (N_6084,N_4997,N_4678);
or U6085 (N_6085,N_4697,N_5687);
xor U6086 (N_6086,N_5655,N_5778);
and U6087 (N_6087,N_5710,N_5056);
nor U6088 (N_6088,N_5983,N_4935);
or U6089 (N_6089,N_4904,N_5320);
nor U6090 (N_6090,N_4800,N_4642);
or U6091 (N_6091,N_5894,N_5841);
xor U6092 (N_6092,N_4510,N_5586);
and U6093 (N_6093,N_5416,N_5305);
and U6094 (N_6094,N_5481,N_5542);
nor U6095 (N_6095,N_4708,N_4967);
or U6096 (N_6096,N_5509,N_4882);
nor U6097 (N_6097,N_5955,N_5303);
nor U6098 (N_6098,N_5824,N_5570);
nand U6099 (N_6099,N_5216,N_5282);
nand U6100 (N_6100,N_4993,N_5261);
xnor U6101 (N_6101,N_4587,N_4557);
or U6102 (N_6102,N_5354,N_5330);
xor U6103 (N_6103,N_5333,N_4698);
or U6104 (N_6104,N_5228,N_4536);
and U6105 (N_6105,N_5666,N_5415);
and U6106 (N_6106,N_5044,N_5078);
nand U6107 (N_6107,N_5199,N_5383);
or U6108 (N_6108,N_5502,N_5735);
or U6109 (N_6109,N_5034,N_5226);
nor U6110 (N_6110,N_5065,N_4702);
or U6111 (N_6111,N_5969,N_4629);
nand U6112 (N_6112,N_5125,N_4790);
and U6113 (N_6113,N_5243,N_5535);
or U6114 (N_6114,N_4612,N_4755);
and U6115 (N_6115,N_5943,N_5604);
nand U6116 (N_6116,N_4673,N_5723);
or U6117 (N_6117,N_5158,N_5471);
xnor U6118 (N_6118,N_5108,N_5641);
and U6119 (N_6119,N_4506,N_5277);
and U6120 (N_6120,N_5879,N_4782);
or U6121 (N_6121,N_5499,N_5238);
and U6122 (N_6122,N_4945,N_5904);
nor U6123 (N_6123,N_4726,N_4897);
nand U6124 (N_6124,N_5007,N_5736);
xor U6125 (N_6125,N_4964,N_5803);
nand U6126 (N_6126,N_5770,N_4692);
and U6127 (N_6127,N_4783,N_5699);
or U6128 (N_6128,N_5755,N_5668);
or U6129 (N_6129,N_4579,N_4953);
or U6130 (N_6130,N_5730,N_5328);
nor U6131 (N_6131,N_5311,N_5965);
and U6132 (N_6132,N_4610,N_4648);
xnor U6133 (N_6133,N_5436,N_4672);
nor U6134 (N_6134,N_4900,N_4865);
nand U6135 (N_6135,N_4696,N_4826);
nor U6136 (N_6136,N_4877,N_4884);
and U6137 (N_6137,N_5628,N_5772);
nor U6138 (N_6138,N_5689,N_4963);
nand U6139 (N_6139,N_5086,N_4854);
nor U6140 (N_6140,N_4756,N_5254);
nand U6141 (N_6141,N_5620,N_5087);
nand U6142 (N_6142,N_5575,N_4784);
and U6143 (N_6143,N_4778,N_5554);
and U6144 (N_6144,N_5656,N_5667);
or U6145 (N_6145,N_5145,N_5653);
or U6146 (N_6146,N_5004,N_4855);
xnor U6147 (N_6147,N_4645,N_4816);
and U6148 (N_6148,N_5521,N_4737);
or U6149 (N_6149,N_5392,N_4627);
and U6150 (N_6150,N_4974,N_4739);
xor U6151 (N_6151,N_5283,N_5359);
and U6152 (N_6152,N_5148,N_5914);
xor U6153 (N_6153,N_5684,N_5116);
nor U6154 (N_6154,N_5083,N_4514);
and U6155 (N_6155,N_5114,N_5633);
nor U6156 (N_6156,N_4938,N_4991);
and U6157 (N_6157,N_5230,N_4720);
xnor U6158 (N_6158,N_5163,N_4954);
nand U6159 (N_6159,N_5886,N_4607);
nand U6160 (N_6160,N_4547,N_5141);
xor U6161 (N_6161,N_4825,N_5589);
xor U6162 (N_6162,N_4543,N_5253);
or U6163 (N_6163,N_4883,N_4528);
nor U6164 (N_6164,N_5149,N_5865);
xnor U6165 (N_6165,N_4928,N_5753);
xor U6166 (N_6166,N_4910,N_5657);
xor U6167 (N_6167,N_4631,N_4803);
nand U6168 (N_6168,N_4699,N_5534);
xor U6169 (N_6169,N_4859,N_5182);
and U6170 (N_6170,N_5260,N_5097);
and U6171 (N_6171,N_5105,N_5246);
xor U6172 (N_6172,N_4920,N_5062);
nor U6173 (N_6173,N_5150,N_4577);
and U6174 (N_6174,N_4622,N_5501);
nand U6175 (N_6175,N_5232,N_5109);
nor U6176 (N_6176,N_5255,N_4597);
or U6177 (N_6177,N_5754,N_4734);
and U6178 (N_6178,N_5122,N_5677);
nand U6179 (N_6179,N_5269,N_5119);
xnor U6180 (N_6180,N_5682,N_4594);
xnor U6181 (N_6181,N_4824,N_5142);
or U6182 (N_6182,N_4522,N_5627);
xnor U6183 (N_6183,N_4643,N_4606);
or U6184 (N_6184,N_5073,N_5808);
xnor U6185 (N_6185,N_5802,N_5401);
or U6186 (N_6186,N_5507,N_5398);
xor U6187 (N_6187,N_5010,N_5021);
xnor U6188 (N_6188,N_4628,N_5556);
xnor U6189 (N_6189,N_4950,N_5278);
nand U6190 (N_6190,N_5379,N_4608);
nand U6191 (N_6191,N_5130,N_5769);
and U6192 (N_6192,N_5997,N_5463);
xnor U6193 (N_6193,N_5630,N_5411);
nand U6194 (N_6194,N_4988,N_5746);
or U6195 (N_6195,N_4898,N_5531);
nor U6196 (N_6196,N_5176,N_4728);
xor U6197 (N_6197,N_4860,N_5767);
xnor U6198 (N_6198,N_5934,N_5618);
or U6199 (N_6199,N_5979,N_5805);
xor U6200 (N_6200,N_5870,N_5350);
or U6201 (N_6201,N_5779,N_5910);
nor U6202 (N_6202,N_5893,N_4637);
or U6203 (N_6203,N_5733,N_5066);
nor U6204 (N_6204,N_4574,N_5695);
or U6205 (N_6205,N_5171,N_5023);
and U6206 (N_6206,N_5966,N_4903);
xnor U6207 (N_6207,N_5822,N_5055);
nor U6208 (N_6208,N_5786,N_5764);
or U6209 (N_6209,N_5672,N_5727);
nor U6210 (N_6210,N_5536,N_4949);
xnor U6211 (N_6211,N_5784,N_4552);
and U6212 (N_6212,N_4902,N_5545);
or U6213 (N_6213,N_5909,N_5610);
xor U6214 (N_6214,N_5138,N_5587);
xnor U6215 (N_6215,N_5892,N_5584);
xor U6216 (N_6216,N_5898,N_5578);
and U6217 (N_6217,N_4504,N_5920);
xnor U6218 (N_6218,N_5325,N_5825);
nand U6219 (N_6219,N_5818,N_5203);
nand U6220 (N_6220,N_5938,N_5069);
nand U6221 (N_6221,N_4625,N_4852);
nor U6222 (N_6222,N_5718,N_4650);
nor U6223 (N_6223,N_5530,N_5771);
nor U6224 (N_6224,N_5991,N_4802);
nand U6225 (N_6225,N_5712,N_4655);
or U6226 (N_6226,N_4667,N_5624);
nor U6227 (N_6227,N_5696,N_5143);
and U6228 (N_6228,N_4817,N_5506);
xor U6229 (N_6229,N_4729,N_5479);
or U6230 (N_6230,N_4531,N_5751);
and U6231 (N_6231,N_5555,N_5981);
or U6232 (N_6232,N_5096,N_5498);
nor U6233 (N_6233,N_5067,N_5386);
or U6234 (N_6234,N_5206,N_5315);
or U6235 (N_6235,N_4986,N_5504);
nor U6236 (N_6236,N_4589,N_5413);
and U6237 (N_6237,N_5154,N_4789);
or U6238 (N_6238,N_5178,N_5744);
or U6239 (N_6239,N_4913,N_5982);
and U6240 (N_6240,N_5877,N_5738);
xor U6241 (N_6241,N_5172,N_4529);
nor U6242 (N_6242,N_5813,N_5862);
and U6243 (N_6243,N_4971,N_5399);
or U6244 (N_6244,N_4779,N_5622);
and U6245 (N_6245,N_5717,N_5423);
nand U6246 (N_6246,N_5839,N_5070);
nor U6247 (N_6247,N_5218,N_4685);
xnor U6248 (N_6248,N_5547,N_4660);
nand U6249 (N_6249,N_5963,N_5153);
xor U6250 (N_6250,N_5280,N_5976);
and U6251 (N_6251,N_5431,N_5136);
xnor U6252 (N_6252,N_4586,N_4942);
xor U6253 (N_6253,N_4982,N_5798);
xnor U6254 (N_6254,N_5357,N_5496);
xnor U6255 (N_6255,N_4588,N_5806);
nor U6256 (N_6256,N_5644,N_4544);
xor U6257 (N_6257,N_4752,N_5537);
nand U6258 (N_6258,N_5766,N_4841);
nand U6259 (N_6259,N_5941,N_5049);
and U6260 (N_6260,N_5579,N_5936);
and U6261 (N_6261,N_4787,N_4960);
or U6262 (N_6262,N_4909,N_5345);
nor U6263 (N_6263,N_5334,N_5944);
and U6264 (N_6264,N_4970,N_5815);
xor U6265 (N_6265,N_5722,N_4758);
nand U6266 (N_6266,N_5564,N_5640);
nand U6267 (N_6267,N_5758,N_5406);
nor U6268 (N_6268,N_5590,N_5180);
nor U6269 (N_6269,N_5292,N_5395);
xnor U6270 (N_6270,N_5249,N_5671);
nor U6271 (N_6271,N_5051,N_5876);
nand U6272 (N_6272,N_5608,N_4640);
and U6273 (N_6273,N_4844,N_5662);
nor U6274 (N_6274,N_4603,N_5494);
nor U6275 (N_6275,N_5410,N_4966);
or U6276 (N_6276,N_5500,N_4929);
xnor U6277 (N_6277,N_4893,N_4630);
and U6278 (N_6278,N_5472,N_5864);
nor U6279 (N_6279,N_5514,N_4717);
xor U6280 (N_6280,N_4500,N_5785);
and U6281 (N_6281,N_4767,N_4560);
and U6282 (N_6282,N_4714,N_5322);
and U6283 (N_6283,N_5019,N_4639);
xor U6284 (N_6284,N_4540,N_5510);
xnor U6285 (N_6285,N_4745,N_4766);
nand U6286 (N_6286,N_5937,N_5185);
xnor U6287 (N_6287,N_5792,N_5543);
nor U6288 (N_6288,N_4821,N_5670);
or U6289 (N_6289,N_5683,N_4669);
nor U6290 (N_6290,N_5404,N_5698);
or U6291 (N_6291,N_4918,N_4927);
and U6292 (N_6292,N_4831,N_5058);
xnor U6293 (N_6293,N_5375,N_5552);
nand U6294 (N_6294,N_5495,N_4980);
nor U6295 (N_6295,N_5313,N_5739);
nor U6296 (N_6296,N_5035,N_4861);
nor U6297 (N_6297,N_4815,N_4881);
xnor U6298 (N_6298,N_5337,N_4958);
or U6299 (N_6299,N_4677,N_4710);
xnor U6300 (N_6300,N_5252,N_5264);
xnor U6301 (N_6301,N_5884,N_5849);
xnor U6302 (N_6302,N_4600,N_4762);
nor U6303 (N_6303,N_5102,N_5486);
or U6304 (N_6304,N_4890,N_5371);
nand U6305 (N_6305,N_4839,N_5000);
nand U6306 (N_6306,N_5615,N_5440);
and U6307 (N_6307,N_4664,N_5492);
xor U6308 (N_6308,N_4917,N_5133);
xor U6309 (N_6309,N_5281,N_5110);
xnor U6310 (N_6310,N_5525,N_4749);
and U6311 (N_6311,N_5692,N_5024);
or U6312 (N_6312,N_5121,N_4754);
or U6313 (N_6313,N_5342,N_4932);
and U6314 (N_6314,N_5874,N_5939);
nand U6315 (N_6315,N_4675,N_5284);
nand U6316 (N_6316,N_4901,N_5188);
or U6317 (N_6317,N_5239,N_4743);
nand U6318 (N_6318,N_5810,N_5236);
nand U6319 (N_6319,N_4674,N_4773);
and U6320 (N_6320,N_5838,N_4501);
nand U6321 (N_6321,N_5706,N_4623);
or U6322 (N_6322,N_4799,N_5316);
or U6323 (N_6323,N_5990,N_5924);
nand U6324 (N_6324,N_4879,N_5609);
xor U6325 (N_6325,N_5998,N_5566);
xor U6326 (N_6326,N_4753,N_5956);
and U6327 (N_6327,N_5861,N_5889);
xnor U6328 (N_6328,N_5752,N_5945);
and U6329 (N_6329,N_5351,N_5974);
nand U6330 (N_6330,N_5204,N_5658);
nor U6331 (N_6331,N_5214,N_4617);
and U6332 (N_6332,N_5908,N_5290);
and U6333 (N_6333,N_5196,N_4615);
xor U6334 (N_6334,N_5928,N_5580);
nor U6335 (N_6335,N_4690,N_4680);
xor U6336 (N_6336,N_5104,N_5030);
nor U6337 (N_6337,N_5447,N_5327);
nor U6338 (N_6338,N_5437,N_4713);
xnor U6339 (N_6339,N_4687,N_5899);
nand U6340 (N_6340,N_5276,N_5643);
and U6341 (N_6341,N_5905,N_4820);
nor U6342 (N_6342,N_5635,N_4907);
nand U6343 (N_6343,N_5716,N_5549);
nor U6344 (N_6344,N_5266,N_5794);
xnor U6345 (N_6345,N_5299,N_4718);
xor U6346 (N_6346,N_4905,N_5688);
and U6347 (N_6347,N_4611,N_5593);
nand U6348 (N_6348,N_5996,N_5967);
and U6349 (N_6349,N_5572,N_5947);
or U6350 (N_6350,N_4797,N_4842);
xnor U6351 (N_6351,N_5092,N_4886);
nor U6352 (N_6352,N_4856,N_4810);
and U6353 (N_6353,N_5517,N_5680);
nand U6354 (N_6354,N_4780,N_4978);
nand U6355 (N_6355,N_5827,N_5174);
nor U6356 (N_6356,N_5124,N_4838);
nand U6357 (N_6357,N_4936,N_5013);
xnor U6358 (N_6358,N_5823,N_5037);
nand U6359 (N_6359,N_5361,N_4661);
nor U6360 (N_6360,N_4716,N_4804);
or U6361 (N_6361,N_4926,N_4837);
and U6362 (N_6362,N_5592,N_5724);
and U6363 (N_6363,N_4806,N_5179);
xor U6364 (N_6364,N_5458,N_4647);
nor U6365 (N_6365,N_4862,N_5617);
nor U6366 (N_6366,N_5557,N_5745);
xnor U6367 (N_6367,N_4946,N_5054);
nand U6368 (N_6368,N_4703,N_4613);
nor U6369 (N_6369,N_5011,N_5972);
nand U6370 (N_6370,N_5599,N_5546);
nand U6371 (N_6371,N_4840,N_5984);
and U6372 (N_6372,N_5467,N_5466);
xnor U6373 (N_6373,N_5989,N_4930);
and U6374 (N_6374,N_5167,N_5987);
and U6375 (N_6375,N_5272,N_5372);
nor U6376 (N_6376,N_5265,N_5215);
or U6377 (N_6377,N_5363,N_4965);
xor U6378 (N_6378,N_4638,N_5851);
nand U6379 (N_6379,N_5120,N_4880);
or U6380 (N_6380,N_5353,N_5523);
or U6381 (N_6381,N_4576,N_4757);
xor U6382 (N_6382,N_5860,N_5168);
and U6383 (N_6383,N_4569,N_4558);
and U6384 (N_6384,N_5650,N_5749);
xnor U6385 (N_6385,N_5484,N_5407);
nand U6386 (N_6386,N_4836,N_5776);
and U6387 (N_6387,N_4771,N_5659);
or U6388 (N_6388,N_4934,N_5100);
nand U6389 (N_6389,N_5594,N_5598);
or U6390 (N_6390,N_5297,N_5853);
nor U6391 (N_6391,N_5780,N_5039);
or U6392 (N_6392,N_5480,N_4770);
nand U6393 (N_6393,N_5878,N_5917);
xor U6394 (N_6394,N_5707,N_5888);
nor U6395 (N_6395,N_4873,N_4922);
and U6396 (N_6396,N_5747,N_4751);
xor U6397 (N_6397,N_4633,N_5224);
and U6398 (N_6398,N_4651,N_5637);
nor U6399 (N_6399,N_5804,N_5836);
xnor U6400 (N_6400,N_5863,N_5160);
or U6401 (N_6401,N_4869,N_4519);
or U6402 (N_6402,N_4538,N_5068);
nor U6403 (N_6403,N_5797,N_4781);
and U6404 (N_6404,N_4740,N_4634);
xnor U6405 (N_6405,N_4649,N_4549);
xnor U6406 (N_6406,N_5903,N_4666);
nor U6407 (N_6407,N_5693,N_5126);
xor U6408 (N_6408,N_5352,N_5567);
and U6409 (N_6409,N_5309,N_5288);
or U6410 (N_6410,N_4595,N_4537);
xor U6411 (N_6411,N_5519,N_5324);
and U6412 (N_6412,N_4503,N_5740);
and U6413 (N_6413,N_4834,N_5428);
and U6414 (N_6414,N_5895,N_5703);
xor U6415 (N_6415,N_4580,N_4525);
xor U6416 (N_6416,N_5429,N_5512);
nor U6417 (N_6417,N_4533,N_5192);
or U6418 (N_6418,N_4567,N_4596);
xor U6419 (N_6419,N_5935,N_4724);
and U6420 (N_6420,N_5631,N_5101);
or U6421 (N_6421,N_5602,N_5959);
or U6422 (N_6422,N_5923,N_5151);
xor U6423 (N_6423,N_5664,N_5845);
nand U6424 (N_6424,N_4731,N_4968);
or U6425 (N_6425,N_5814,N_5417);
xnor U6426 (N_6426,N_4868,N_5781);
nor U6427 (N_6427,N_4774,N_5875);
or U6428 (N_6428,N_4940,N_5508);
nand U6429 (N_6429,N_5562,N_5485);
and U6430 (N_6430,N_4727,N_5491);
nand U6431 (N_6431,N_4693,N_5473);
nor U6432 (N_6432,N_4684,N_4941);
nor U6433 (N_6433,N_5623,N_5801);
and U6434 (N_6434,N_5694,N_5164);
and U6435 (N_6435,N_5912,N_5950);
nand U6436 (N_6436,N_5219,N_4829);
and U6437 (N_6437,N_5047,N_4686);
nand U6438 (N_6438,N_5442,N_5930);
or U6439 (N_6439,N_5170,N_5128);
xor U6440 (N_6440,N_4760,N_5085);
nor U6441 (N_6441,N_4712,N_5184);
or U6442 (N_6442,N_5661,N_5451);
or U6443 (N_6443,N_5891,N_5190);
xor U6444 (N_6444,N_5871,N_4694);
nor U6445 (N_6445,N_4895,N_5307);
and U6446 (N_6446,N_4955,N_4990);
nand U6447 (N_6447,N_5369,N_5711);
and U6448 (N_6448,N_4924,N_5953);
or U6449 (N_6449,N_4811,N_5026);
or U6450 (N_6450,N_5980,N_5090);
and U6451 (N_6451,N_5223,N_4996);
and U6452 (N_6452,N_5425,N_5783);
nor U6453 (N_6453,N_5607,N_5256);
or U6454 (N_6454,N_5088,N_4818);
or U6455 (N_6455,N_4992,N_5343);
and U6456 (N_6456,N_5478,N_5949);
nand U6457 (N_6457,N_5629,N_5726);
xor U6458 (N_6458,N_5576,N_5446);
nand U6459 (N_6459,N_4987,N_4590);
or U6460 (N_6460,N_5326,N_5713);
and U6461 (N_6461,N_4591,N_5298);
or U6462 (N_6462,N_5355,N_4763);
nand U6463 (N_6463,N_5887,N_4527);
or U6464 (N_6464,N_4691,N_5384);
or U6465 (N_6465,N_5958,N_5443);
or U6466 (N_6466,N_4556,N_5459);
and U6467 (N_6467,N_5059,N_5162);
nand U6468 (N_6468,N_5367,N_4801);
or U6469 (N_6469,N_5962,N_5402);
nor U6470 (N_6470,N_5323,N_4542);
xor U6471 (N_6471,N_5331,N_5107);
nand U6472 (N_6472,N_4915,N_5414);
and U6473 (N_6473,N_4671,N_5227);
or U6474 (N_6474,N_4524,N_4973);
nor U6475 (N_6475,N_4916,N_5800);
and U6476 (N_6476,N_4866,N_5691);
xnor U6477 (N_6477,N_5135,N_4843);
and U6478 (N_6478,N_5079,N_4721);
nand U6479 (N_6479,N_4931,N_5559);
nor U6480 (N_6480,N_5202,N_5619);
or U6481 (N_6481,N_5348,N_5385);
nand U6482 (N_6482,N_5457,N_5312);
or U6483 (N_6483,N_5977,N_5922);
and U6484 (N_6484,N_5476,N_5205);
and U6485 (N_6485,N_4981,N_5807);
or U6486 (N_6486,N_5588,N_4746);
or U6487 (N_6487,N_5183,N_5714);
nand U6488 (N_6488,N_4937,N_5248);
nand U6489 (N_6489,N_5081,N_4807);
or U6490 (N_6490,N_5690,N_5568);
or U6491 (N_6491,N_5732,N_4626);
nor U6492 (N_6492,N_5830,N_5050);
and U6493 (N_6493,N_4668,N_5419);
or U6494 (N_6494,N_5819,N_5649);
nor U6495 (N_6495,N_5434,N_4592);
xnor U6496 (N_6496,N_5468,N_5165);
xor U6497 (N_6497,N_5111,N_4887);
or U6498 (N_6498,N_5533,N_4911);
and U6499 (N_6499,N_4601,N_5048);
and U6500 (N_6500,N_5634,N_5106);
nor U6501 (N_6501,N_5933,N_5041);
xor U6502 (N_6502,N_5720,N_5103);
nor U6503 (N_6503,N_4830,N_4785);
xor U6504 (N_6504,N_5709,N_5854);
and U6505 (N_6505,N_5389,N_5529);
nand U6506 (N_6506,N_5187,N_5489);
nor U6507 (N_6507,N_5140,N_5993);
nor U6508 (N_6508,N_5430,N_5970);
nor U6509 (N_6509,N_5289,N_5382);
nand U6510 (N_6510,N_4605,N_5663);
or U6511 (N_6511,N_4621,N_5306);
and U6512 (N_6512,N_5837,N_5700);
nand U6513 (N_6513,N_4517,N_4921);
nand U6514 (N_6514,N_5275,N_5220);
nand U6515 (N_6515,N_5009,N_4977);
xor U6516 (N_6516,N_5014,N_4944);
or U6517 (N_6517,N_5329,N_5270);
and U6518 (N_6518,N_5159,N_4742);
or U6519 (N_6519,N_5426,N_4867);
nor U6520 (N_6520,N_5200,N_4748);
and U6521 (N_6521,N_5789,N_5450);
and U6522 (N_6522,N_4914,N_5396);
nand U6523 (N_6523,N_4951,N_5708);
or U6524 (N_6524,N_4502,N_4515);
nor U6525 (N_6525,N_5018,N_4679);
xor U6526 (N_6526,N_5424,N_5221);
xor U6527 (N_6527,N_5907,N_5605);
xnor U6528 (N_6528,N_5317,N_5127);
or U6529 (N_6529,N_5082,N_5728);
or U6530 (N_6530,N_5274,N_5123);
nand U6531 (N_6531,N_4715,N_5788);
nand U6532 (N_6532,N_4750,N_4632);
nor U6533 (N_6533,N_4952,N_4947);
xor U6534 (N_6534,N_4857,N_5900);
nor U6535 (N_6535,N_5971,N_5229);
nand U6536 (N_6536,N_5882,N_4583);
and U6537 (N_6537,N_5469,N_5460);
nor U6538 (N_6538,N_5279,N_5646);
and U6539 (N_6539,N_5043,N_5453);
or U6540 (N_6540,N_5881,N_5173);
nand U6541 (N_6541,N_4796,N_4584);
and U6542 (N_6542,N_5020,N_4933);
nand U6543 (N_6543,N_5461,N_5574);
nor U6544 (N_6544,N_4688,N_5077);
xnor U6545 (N_6545,N_5267,N_4943);
and U6546 (N_6546,N_5391,N_4665);
and U6547 (N_6547,N_4984,N_5516);
nand U6548 (N_6548,N_5412,N_5497);
and U6549 (N_6549,N_4593,N_5462);
or U6550 (N_6550,N_5057,N_5625);
nor U6551 (N_6551,N_5217,N_5697);
nor U6552 (N_6552,N_5042,N_5347);
nand U6553 (N_6553,N_5606,N_5118);
and U6554 (N_6554,N_5520,N_5850);
nand U6555 (N_6555,N_5921,N_5597);
or U6556 (N_6556,N_4735,N_5774);
and U6557 (N_6557,N_4969,N_5181);
nand U6558 (N_6558,N_5341,N_5812);
nor U6559 (N_6559,N_5505,N_5873);
xnor U6560 (N_6560,N_5210,N_4814);
nor U6561 (N_6561,N_5017,N_4959);
and U6562 (N_6562,N_5465,N_5063);
nand U6563 (N_6563,N_4561,N_5913);
or U6564 (N_6564,N_4871,N_5117);
nand U6565 (N_6565,N_5986,N_5725);
nand U6566 (N_6566,N_5621,N_5015);
or U6567 (N_6567,N_5247,N_5259);
nor U6568 (N_6568,N_5524,N_4956);
or U6569 (N_6569,N_4523,N_5846);
and U6570 (N_6570,N_5515,N_4858);
nor U6571 (N_6571,N_5474,N_4983);
nand U6572 (N_6572,N_5890,N_5926);
xor U6573 (N_6573,N_4888,N_4985);
nand U6574 (N_6574,N_5743,N_5433);
xor U6575 (N_6575,N_4772,N_5005);
nor U6576 (N_6576,N_5080,N_5756);
nor U6577 (N_6577,N_5390,N_4849);
nand U6578 (N_6578,N_5374,N_5603);
nor U6579 (N_6579,N_5432,N_5585);
or U6580 (N_6580,N_4530,N_5675);
nor U6581 (N_6581,N_5701,N_5129);
or U6582 (N_6582,N_5339,N_4706);
xor U6583 (N_6583,N_5115,N_4738);
nor U6584 (N_6584,N_5995,N_5811);
and U6585 (N_6585,N_5681,N_5999);
nor U6586 (N_6586,N_5669,N_5777);
or U6587 (N_6587,N_5134,N_5338);
or U6588 (N_6588,N_4553,N_5296);
or U6589 (N_6589,N_5795,N_5061);
and U6590 (N_6590,N_5831,N_5356);
nand U6591 (N_6591,N_5582,N_5639);
or U6592 (N_6592,N_5157,N_5918);
and U6593 (N_6593,N_5099,N_4828);
xor U6594 (N_6594,N_5569,N_5522);
or U6595 (N_6595,N_5760,N_4823);
and U6596 (N_6596,N_5318,N_5832);
or U6597 (N_6597,N_5365,N_4578);
or U6598 (N_6598,N_5869,N_5155);
nand U6599 (N_6599,N_5089,N_5393);
or U6600 (N_6600,N_5834,N_4885);
and U6601 (N_6601,N_5156,N_5539);
nor U6602 (N_6602,N_4705,N_5209);
xnor U6603 (N_6603,N_4759,N_5006);
or U6604 (N_6604,N_5940,N_5211);
or U6605 (N_6605,N_5191,N_4573);
or U6606 (N_6606,N_4701,N_4793);
or U6607 (N_6607,N_5858,N_4805);
and U6608 (N_6608,N_5483,N_5957);
xor U6609 (N_6609,N_5001,N_5676);
nor U6610 (N_6610,N_5757,N_5782);
or U6611 (N_6611,N_5378,N_5076);
nand U6612 (N_6612,N_4526,N_5759);
nor U6613 (N_6613,N_5045,N_4508);
nor U6614 (N_6614,N_4853,N_4994);
nand U6615 (N_6615,N_4700,N_5405);
or U6616 (N_6616,N_5310,N_4653);
xnor U6617 (N_6617,N_5614,N_5340);
nand U6618 (N_6618,N_5868,N_4979);
or U6619 (N_6619,N_4507,N_4620);
xor U6620 (N_6620,N_5742,N_5377);
nor U6621 (N_6621,N_4809,N_4559);
xor U6622 (N_6622,N_5503,N_5852);
nand U6623 (N_6623,N_5349,N_5319);
and U6624 (N_6624,N_5302,N_4795);
nand U6625 (N_6625,N_5960,N_5449);
nand U6626 (N_6626,N_4736,N_5561);
nand U6627 (N_6627,N_5394,N_5600);
nor U6628 (N_6628,N_5638,N_5847);
or U6629 (N_6629,N_4709,N_5064);
or U6630 (N_6630,N_5144,N_4575);
xor U6631 (N_6631,N_4572,N_4957);
nand U6632 (N_6632,N_5817,N_5842);
xor U6633 (N_6633,N_5560,N_5147);
or U6634 (N_6634,N_4570,N_5826);
xor U6635 (N_6635,N_5946,N_4876);
nand U6636 (N_6636,N_5916,N_4863);
nor U6637 (N_6637,N_5978,N_4864);
nand U6638 (N_6638,N_4546,N_4776);
nand U6639 (N_6639,N_4791,N_4571);
xnor U6640 (N_6640,N_5262,N_5927);
or U6641 (N_6641,N_5177,N_5768);
and U6642 (N_6642,N_5376,N_5360);
or U6643 (N_6643,N_4827,N_5809);
or U6644 (N_6644,N_5094,N_4564);
xnor U6645 (N_6645,N_4870,N_5233);
xnor U6646 (N_6646,N_5362,N_5113);
xnor U6647 (N_6647,N_5591,N_4744);
nand U6648 (N_6648,N_5053,N_4961);
nor U6649 (N_6649,N_5212,N_5883);
xor U6650 (N_6650,N_5773,N_5948);
or U6651 (N_6651,N_4813,N_5636);
or U6652 (N_6652,N_4670,N_5673);
nor U6653 (N_6653,N_5388,N_5737);
xor U6654 (N_6654,N_4541,N_5093);
nand U6655 (N_6655,N_5146,N_4614);
and U6656 (N_6656,N_5538,N_5721);
xor U6657 (N_6657,N_4733,N_4554);
or U6658 (N_6658,N_5366,N_5902);
nand U6659 (N_6659,N_5550,N_5790);
nand U6660 (N_6660,N_5613,N_5527);
xnor U6661 (N_6661,N_5678,N_5263);
or U6662 (N_6662,N_5456,N_5541);
xor U6663 (N_6663,N_4624,N_5420);
nor U6664 (N_6664,N_5091,N_5765);
or U6665 (N_6665,N_5762,N_5244);
and U6666 (N_6666,N_5040,N_5295);
and U6667 (N_6667,N_5866,N_5951);
xor U6668 (N_6668,N_4912,N_4899);
xor U6669 (N_6669,N_5346,N_4775);
nand U6670 (N_6670,N_4822,N_4656);
nor U6671 (N_6671,N_5301,N_5344);
nand U6672 (N_6672,N_5919,N_5968);
or U6673 (N_6673,N_5074,N_5195);
and U6674 (N_6674,N_5022,N_5581);
or U6675 (N_6675,N_5207,N_5964);
nor U6676 (N_6676,N_5848,N_4707);
and U6677 (N_6677,N_5954,N_5038);
nor U6678 (N_6678,N_4769,N_4819);
or U6679 (N_6679,N_4654,N_4999);
or U6680 (N_6680,N_5715,N_4582);
and U6681 (N_6681,N_4765,N_5308);
nand U6682 (N_6682,N_5994,N_5137);
nand U6683 (N_6683,N_5932,N_5287);
or U6684 (N_6684,N_5488,N_5033);
and U6685 (N_6685,N_4511,N_5364);
nand U6686 (N_6686,N_5704,N_5387);
xor U6687 (N_6687,N_5234,N_4550);
or U6688 (N_6688,N_5674,N_5235);
or U6689 (N_6689,N_5595,N_4878);
nand U6690 (N_6690,N_4619,N_5748);
nor U6691 (N_6691,N_4704,N_5189);
or U6692 (N_6692,N_5645,N_5250);
or U6693 (N_6693,N_5439,N_4681);
nor U6694 (N_6694,N_5241,N_4875);
or U6695 (N_6695,N_5548,N_4609);
and U6696 (N_6696,N_5455,N_5611);
nor U6697 (N_6697,N_5490,N_4874);
or U6698 (N_6698,N_4657,N_5843);
nand U6699 (N_6699,N_4695,N_4545);
nor U6700 (N_6700,N_4948,N_5632);
or U6701 (N_6701,N_5616,N_5612);
or U6702 (N_6702,N_4777,N_5796);
xnor U6703 (N_6703,N_5271,N_5012);
and U6704 (N_6704,N_5648,N_5027);
or U6705 (N_6705,N_5511,N_5526);
nor U6706 (N_6706,N_4792,N_4518);
xor U6707 (N_6707,N_5929,N_5358);
and U6708 (N_6708,N_5071,N_4832);
nand U6709 (N_6709,N_4786,N_5477);
nor U6710 (N_6710,N_4516,N_5652);
or U6711 (N_6711,N_4989,N_5482);
and U6712 (N_6712,N_4535,N_4972);
nand U6713 (N_6713,N_4548,N_5855);
and U6714 (N_6714,N_4722,N_4532);
and U6715 (N_6715,N_4891,N_5761);
nor U6716 (N_6716,N_4730,N_5237);
nand U6717 (N_6717,N_4845,N_4851);
and U6718 (N_6718,N_5408,N_5095);
nand U6719 (N_6719,N_5750,N_4534);
or U6720 (N_6720,N_4925,N_5470);
xnor U6721 (N_6721,N_5098,N_4732);
nor U6722 (N_6722,N_5571,N_5464);
or U6723 (N_6723,N_5194,N_5169);
nor U6724 (N_6724,N_5719,N_4659);
or U6725 (N_6725,N_4683,N_4602);
nor U6726 (N_6726,N_5016,N_4689);
and U6727 (N_6727,N_5161,N_4741);
or U6728 (N_6728,N_5293,N_4505);
nor U6729 (N_6729,N_5257,N_5528);
nor U6730 (N_6730,N_5438,N_5427);
and U6731 (N_6731,N_5084,N_5791);
or U6732 (N_6732,N_5513,N_5028);
and U6733 (N_6733,N_5418,N_5197);
and U6734 (N_6734,N_5885,N_5285);
xnor U6735 (N_6735,N_5867,N_5911);
nand U6736 (N_6736,N_5844,N_4889);
nor U6737 (N_6737,N_5820,N_4768);
nor U6738 (N_6738,N_5435,N_5336);
nor U6739 (N_6739,N_4644,N_4764);
nand U6740 (N_6740,N_5403,N_4599);
xor U6741 (N_6741,N_5741,N_4618);
nand U6742 (N_6742,N_5518,N_4555);
nor U6743 (N_6743,N_5925,N_4892);
and U6744 (N_6744,N_5973,N_4616);
nand U6745 (N_6745,N_5046,N_4798);
nor U6746 (N_6746,N_4894,N_5915);
and U6747 (N_6747,N_5601,N_5060);
or U6748 (N_6748,N_4923,N_4563);
xnor U6749 (N_6749,N_5596,N_5258);
xor U6750 (N_6750,N_4523,N_5265);
nor U6751 (N_6751,N_4816,N_5628);
or U6752 (N_6752,N_5272,N_5158);
or U6753 (N_6753,N_5867,N_5055);
and U6754 (N_6754,N_4644,N_5521);
and U6755 (N_6755,N_5465,N_5516);
or U6756 (N_6756,N_5567,N_5175);
and U6757 (N_6757,N_5057,N_5638);
nand U6758 (N_6758,N_4753,N_4721);
nor U6759 (N_6759,N_4539,N_5074);
or U6760 (N_6760,N_4577,N_5770);
and U6761 (N_6761,N_5705,N_5606);
xor U6762 (N_6762,N_4752,N_5197);
xor U6763 (N_6763,N_5738,N_4559);
and U6764 (N_6764,N_4939,N_4909);
nand U6765 (N_6765,N_5047,N_4708);
and U6766 (N_6766,N_4507,N_4983);
and U6767 (N_6767,N_4568,N_5249);
nand U6768 (N_6768,N_4504,N_5214);
or U6769 (N_6769,N_4694,N_5655);
nand U6770 (N_6770,N_4639,N_4648);
xnor U6771 (N_6771,N_4697,N_5077);
or U6772 (N_6772,N_5597,N_4505);
nand U6773 (N_6773,N_4833,N_5719);
and U6774 (N_6774,N_5949,N_5247);
xor U6775 (N_6775,N_5928,N_5938);
nand U6776 (N_6776,N_5905,N_5893);
and U6777 (N_6777,N_4607,N_5359);
nor U6778 (N_6778,N_5546,N_5071);
or U6779 (N_6779,N_5462,N_5381);
nand U6780 (N_6780,N_5787,N_5595);
and U6781 (N_6781,N_4581,N_4504);
nor U6782 (N_6782,N_5896,N_5364);
nand U6783 (N_6783,N_4945,N_4620);
xor U6784 (N_6784,N_5104,N_5576);
xor U6785 (N_6785,N_5081,N_4591);
xor U6786 (N_6786,N_5108,N_5357);
nor U6787 (N_6787,N_5710,N_5385);
nor U6788 (N_6788,N_5219,N_4822);
nand U6789 (N_6789,N_4531,N_5569);
and U6790 (N_6790,N_5133,N_4602);
nor U6791 (N_6791,N_4706,N_5613);
and U6792 (N_6792,N_5929,N_4618);
xor U6793 (N_6793,N_5538,N_4605);
and U6794 (N_6794,N_5685,N_5888);
xor U6795 (N_6795,N_5350,N_4615);
xnor U6796 (N_6796,N_5732,N_5059);
and U6797 (N_6797,N_4993,N_5899);
and U6798 (N_6798,N_5440,N_4913);
nor U6799 (N_6799,N_5556,N_4918);
nor U6800 (N_6800,N_5032,N_5489);
and U6801 (N_6801,N_5749,N_4849);
or U6802 (N_6802,N_5383,N_4957);
or U6803 (N_6803,N_5030,N_5777);
nor U6804 (N_6804,N_4987,N_5626);
nand U6805 (N_6805,N_4923,N_4962);
xnor U6806 (N_6806,N_5742,N_4843);
xnor U6807 (N_6807,N_5602,N_4790);
and U6808 (N_6808,N_5925,N_4558);
xor U6809 (N_6809,N_4898,N_5897);
nor U6810 (N_6810,N_4846,N_5885);
nor U6811 (N_6811,N_5837,N_5010);
nand U6812 (N_6812,N_5236,N_4590);
nand U6813 (N_6813,N_5223,N_5839);
nor U6814 (N_6814,N_5811,N_5132);
or U6815 (N_6815,N_4942,N_5398);
and U6816 (N_6816,N_5007,N_4541);
nor U6817 (N_6817,N_5289,N_5350);
nor U6818 (N_6818,N_5437,N_5592);
nand U6819 (N_6819,N_5236,N_4695);
nand U6820 (N_6820,N_5674,N_4915);
and U6821 (N_6821,N_5912,N_5749);
nand U6822 (N_6822,N_5946,N_5904);
or U6823 (N_6823,N_4711,N_4677);
and U6824 (N_6824,N_4761,N_5134);
and U6825 (N_6825,N_5349,N_5290);
and U6826 (N_6826,N_4518,N_4967);
and U6827 (N_6827,N_5936,N_5495);
and U6828 (N_6828,N_5126,N_4644);
or U6829 (N_6829,N_5895,N_4572);
and U6830 (N_6830,N_5595,N_5364);
xnor U6831 (N_6831,N_5514,N_4881);
xnor U6832 (N_6832,N_5342,N_4959);
or U6833 (N_6833,N_5556,N_5037);
xor U6834 (N_6834,N_5889,N_4811);
and U6835 (N_6835,N_4582,N_5849);
and U6836 (N_6836,N_5277,N_4688);
and U6837 (N_6837,N_5994,N_5702);
and U6838 (N_6838,N_5915,N_4611);
or U6839 (N_6839,N_5497,N_5052);
xor U6840 (N_6840,N_4919,N_4719);
nor U6841 (N_6841,N_5175,N_4864);
or U6842 (N_6842,N_4582,N_4998);
xnor U6843 (N_6843,N_5364,N_5008);
nor U6844 (N_6844,N_5938,N_4927);
xor U6845 (N_6845,N_4546,N_5515);
nand U6846 (N_6846,N_4893,N_5847);
nor U6847 (N_6847,N_4779,N_5862);
nor U6848 (N_6848,N_5845,N_5942);
or U6849 (N_6849,N_4960,N_5002);
nor U6850 (N_6850,N_5339,N_5072);
and U6851 (N_6851,N_4782,N_5754);
xnor U6852 (N_6852,N_5224,N_5298);
nand U6853 (N_6853,N_5733,N_5876);
or U6854 (N_6854,N_5372,N_5059);
xor U6855 (N_6855,N_5493,N_4630);
nand U6856 (N_6856,N_5793,N_4982);
xor U6857 (N_6857,N_4956,N_5720);
nand U6858 (N_6858,N_4671,N_4589);
or U6859 (N_6859,N_5548,N_5029);
xor U6860 (N_6860,N_4797,N_4834);
nand U6861 (N_6861,N_5673,N_4788);
xnor U6862 (N_6862,N_5639,N_5913);
nand U6863 (N_6863,N_5645,N_5839);
or U6864 (N_6864,N_5342,N_5046);
nand U6865 (N_6865,N_5350,N_4863);
nand U6866 (N_6866,N_5400,N_5589);
or U6867 (N_6867,N_5504,N_5451);
nand U6868 (N_6868,N_5536,N_5970);
and U6869 (N_6869,N_5933,N_5287);
or U6870 (N_6870,N_5967,N_5780);
nand U6871 (N_6871,N_5038,N_5170);
or U6872 (N_6872,N_5602,N_4665);
nand U6873 (N_6873,N_5093,N_5107);
xor U6874 (N_6874,N_4513,N_4952);
nand U6875 (N_6875,N_5690,N_5749);
or U6876 (N_6876,N_4898,N_5875);
and U6877 (N_6877,N_4630,N_5858);
or U6878 (N_6878,N_4790,N_4936);
and U6879 (N_6879,N_5209,N_4625);
xor U6880 (N_6880,N_4870,N_5155);
nor U6881 (N_6881,N_4973,N_4775);
xor U6882 (N_6882,N_5614,N_5966);
or U6883 (N_6883,N_5010,N_4959);
and U6884 (N_6884,N_4704,N_5369);
or U6885 (N_6885,N_4986,N_4595);
nand U6886 (N_6886,N_5562,N_5759);
nand U6887 (N_6887,N_5967,N_5011);
and U6888 (N_6888,N_5606,N_4790);
nor U6889 (N_6889,N_4538,N_4784);
nor U6890 (N_6890,N_5048,N_5619);
xor U6891 (N_6891,N_5016,N_5810);
xor U6892 (N_6892,N_5790,N_5431);
and U6893 (N_6893,N_5023,N_4962);
or U6894 (N_6894,N_5074,N_4771);
nand U6895 (N_6895,N_5425,N_5179);
nand U6896 (N_6896,N_4603,N_4553);
and U6897 (N_6897,N_5574,N_5288);
xor U6898 (N_6898,N_5098,N_5179);
nor U6899 (N_6899,N_4811,N_5327);
or U6900 (N_6900,N_5515,N_5555);
nand U6901 (N_6901,N_5713,N_5318);
and U6902 (N_6902,N_4798,N_5136);
or U6903 (N_6903,N_4855,N_4576);
nor U6904 (N_6904,N_5375,N_5512);
and U6905 (N_6905,N_4998,N_5162);
or U6906 (N_6906,N_5579,N_5961);
or U6907 (N_6907,N_5021,N_4748);
and U6908 (N_6908,N_5821,N_5827);
and U6909 (N_6909,N_5524,N_5649);
and U6910 (N_6910,N_5729,N_5612);
nor U6911 (N_6911,N_4599,N_5867);
and U6912 (N_6912,N_5629,N_4640);
nand U6913 (N_6913,N_5790,N_5347);
xnor U6914 (N_6914,N_5215,N_5734);
nand U6915 (N_6915,N_4827,N_5252);
or U6916 (N_6916,N_5442,N_5731);
or U6917 (N_6917,N_5752,N_5541);
xor U6918 (N_6918,N_4614,N_5391);
nand U6919 (N_6919,N_5215,N_5806);
nand U6920 (N_6920,N_5210,N_4555);
nor U6921 (N_6921,N_5189,N_4924);
nor U6922 (N_6922,N_5267,N_5758);
nand U6923 (N_6923,N_5287,N_5264);
xnor U6924 (N_6924,N_4756,N_4853);
nor U6925 (N_6925,N_5526,N_5557);
or U6926 (N_6926,N_5471,N_5005);
or U6927 (N_6927,N_4660,N_4934);
xnor U6928 (N_6928,N_5398,N_5780);
nor U6929 (N_6929,N_5137,N_5579);
nand U6930 (N_6930,N_5383,N_4815);
and U6931 (N_6931,N_5242,N_5470);
and U6932 (N_6932,N_4841,N_4877);
nand U6933 (N_6933,N_4717,N_5008);
or U6934 (N_6934,N_5329,N_5301);
nor U6935 (N_6935,N_5348,N_5554);
and U6936 (N_6936,N_5246,N_4977);
nand U6937 (N_6937,N_5048,N_5773);
xnor U6938 (N_6938,N_5486,N_5481);
and U6939 (N_6939,N_5843,N_5735);
nor U6940 (N_6940,N_5109,N_5399);
or U6941 (N_6941,N_5197,N_5395);
nand U6942 (N_6942,N_5730,N_5593);
nor U6943 (N_6943,N_5363,N_4782);
nor U6944 (N_6944,N_5984,N_5509);
nand U6945 (N_6945,N_5209,N_5002);
nor U6946 (N_6946,N_5834,N_4746);
nor U6947 (N_6947,N_5651,N_5581);
or U6948 (N_6948,N_5018,N_4782);
nand U6949 (N_6949,N_4641,N_5726);
nor U6950 (N_6950,N_5117,N_4530);
nor U6951 (N_6951,N_5090,N_5481);
xnor U6952 (N_6952,N_5590,N_5730);
nand U6953 (N_6953,N_5890,N_5817);
nand U6954 (N_6954,N_5571,N_5311);
xor U6955 (N_6955,N_4947,N_4526);
nor U6956 (N_6956,N_5999,N_5115);
or U6957 (N_6957,N_5679,N_5234);
nand U6958 (N_6958,N_5916,N_5594);
nor U6959 (N_6959,N_4711,N_4810);
or U6960 (N_6960,N_4645,N_5480);
and U6961 (N_6961,N_5897,N_5882);
nor U6962 (N_6962,N_4628,N_4990);
xor U6963 (N_6963,N_5605,N_5880);
nor U6964 (N_6964,N_5517,N_5030);
nor U6965 (N_6965,N_5962,N_5089);
and U6966 (N_6966,N_5075,N_4683);
or U6967 (N_6967,N_4598,N_5896);
and U6968 (N_6968,N_5577,N_5924);
xor U6969 (N_6969,N_5024,N_4633);
nor U6970 (N_6970,N_5939,N_5652);
nand U6971 (N_6971,N_4566,N_5165);
or U6972 (N_6972,N_4832,N_5093);
or U6973 (N_6973,N_5750,N_5640);
or U6974 (N_6974,N_5574,N_4927);
nand U6975 (N_6975,N_5003,N_4705);
or U6976 (N_6976,N_4781,N_5396);
nor U6977 (N_6977,N_4742,N_5226);
xor U6978 (N_6978,N_5097,N_5424);
and U6979 (N_6979,N_5575,N_5365);
or U6980 (N_6980,N_4590,N_4985);
nand U6981 (N_6981,N_4732,N_5989);
nor U6982 (N_6982,N_5434,N_4964);
nor U6983 (N_6983,N_4613,N_5461);
nand U6984 (N_6984,N_5011,N_5785);
and U6985 (N_6985,N_4833,N_4904);
xor U6986 (N_6986,N_5159,N_4978);
nand U6987 (N_6987,N_5305,N_4663);
xor U6988 (N_6988,N_4640,N_5369);
and U6989 (N_6989,N_4945,N_5456);
nand U6990 (N_6990,N_5186,N_5727);
nand U6991 (N_6991,N_5049,N_5834);
xnor U6992 (N_6992,N_4659,N_5877);
and U6993 (N_6993,N_5454,N_5496);
or U6994 (N_6994,N_5588,N_4889);
or U6995 (N_6995,N_5406,N_5038);
or U6996 (N_6996,N_4824,N_5090);
xor U6997 (N_6997,N_5104,N_5388);
and U6998 (N_6998,N_4934,N_5584);
xor U6999 (N_6999,N_5666,N_5568);
and U7000 (N_7000,N_5596,N_5150);
and U7001 (N_7001,N_4683,N_4897);
xor U7002 (N_7002,N_5721,N_5329);
nor U7003 (N_7003,N_4848,N_4802);
nor U7004 (N_7004,N_5126,N_5534);
or U7005 (N_7005,N_4997,N_5727);
and U7006 (N_7006,N_4688,N_5359);
nor U7007 (N_7007,N_4988,N_5477);
xor U7008 (N_7008,N_5187,N_4600);
xnor U7009 (N_7009,N_4943,N_4516);
and U7010 (N_7010,N_5872,N_5683);
xor U7011 (N_7011,N_5134,N_4671);
xor U7012 (N_7012,N_4876,N_5959);
xor U7013 (N_7013,N_5546,N_5240);
nor U7014 (N_7014,N_5451,N_4805);
or U7015 (N_7015,N_5531,N_5071);
nor U7016 (N_7016,N_5713,N_5608);
xor U7017 (N_7017,N_5946,N_5842);
nor U7018 (N_7018,N_4575,N_5795);
nand U7019 (N_7019,N_5217,N_5161);
or U7020 (N_7020,N_5297,N_5349);
nand U7021 (N_7021,N_5813,N_5804);
and U7022 (N_7022,N_5977,N_4832);
or U7023 (N_7023,N_5190,N_5946);
or U7024 (N_7024,N_5629,N_5711);
nor U7025 (N_7025,N_5983,N_4823);
nand U7026 (N_7026,N_5854,N_4787);
or U7027 (N_7027,N_5550,N_4616);
nor U7028 (N_7028,N_5762,N_5643);
nor U7029 (N_7029,N_5402,N_5027);
or U7030 (N_7030,N_5156,N_5586);
xor U7031 (N_7031,N_5617,N_4653);
nor U7032 (N_7032,N_5173,N_4804);
and U7033 (N_7033,N_5214,N_4681);
or U7034 (N_7034,N_5843,N_4804);
and U7035 (N_7035,N_5781,N_5527);
nand U7036 (N_7036,N_4685,N_4562);
nand U7037 (N_7037,N_5670,N_4690);
nand U7038 (N_7038,N_5589,N_5984);
nand U7039 (N_7039,N_5104,N_5877);
xor U7040 (N_7040,N_5972,N_5410);
xnor U7041 (N_7041,N_5357,N_5169);
nor U7042 (N_7042,N_5816,N_4548);
and U7043 (N_7043,N_5365,N_5584);
or U7044 (N_7044,N_4554,N_5907);
and U7045 (N_7045,N_5670,N_5674);
xnor U7046 (N_7046,N_5280,N_5049);
nand U7047 (N_7047,N_4642,N_5247);
or U7048 (N_7048,N_4834,N_5427);
and U7049 (N_7049,N_5127,N_5998);
nor U7050 (N_7050,N_5195,N_5612);
and U7051 (N_7051,N_5748,N_5062);
xor U7052 (N_7052,N_4886,N_5411);
xor U7053 (N_7053,N_4628,N_4541);
and U7054 (N_7054,N_4861,N_5406);
or U7055 (N_7055,N_4616,N_5826);
xnor U7056 (N_7056,N_5736,N_5542);
and U7057 (N_7057,N_4668,N_4792);
xnor U7058 (N_7058,N_5966,N_5244);
or U7059 (N_7059,N_5615,N_5296);
xor U7060 (N_7060,N_4579,N_4968);
nand U7061 (N_7061,N_4681,N_5820);
nor U7062 (N_7062,N_5502,N_4512);
nand U7063 (N_7063,N_4569,N_4568);
nor U7064 (N_7064,N_4733,N_5138);
and U7065 (N_7065,N_5584,N_5066);
and U7066 (N_7066,N_5987,N_5811);
or U7067 (N_7067,N_5809,N_4857);
and U7068 (N_7068,N_5490,N_5265);
xor U7069 (N_7069,N_5065,N_4560);
and U7070 (N_7070,N_4529,N_5078);
xor U7071 (N_7071,N_4623,N_4882);
xor U7072 (N_7072,N_5996,N_5549);
xnor U7073 (N_7073,N_5603,N_5870);
or U7074 (N_7074,N_4632,N_4740);
and U7075 (N_7075,N_5669,N_4614);
nor U7076 (N_7076,N_4758,N_5569);
nor U7077 (N_7077,N_4684,N_5800);
nor U7078 (N_7078,N_5574,N_4797);
nand U7079 (N_7079,N_4508,N_5308);
nand U7080 (N_7080,N_5217,N_4705);
xnor U7081 (N_7081,N_5391,N_5285);
nor U7082 (N_7082,N_5548,N_5733);
nor U7083 (N_7083,N_5550,N_5350);
nand U7084 (N_7084,N_4580,N_5742);
xnor U7085 (N_7085,N_4666,N_5475);
or U7086 (N_7086,N_4962,N_5140);
nor U7087 (N_7087,N_5511,N_4511);
nor U7088 (N_7088,N_5697,N_5205);
nand U7089 (N_7089,N_5835,N_5472);
nand U7090 (N_7090,N_4726,N_5288);
nor U7091 (N_7091,N_5553,N_5704);
nand U7092 (N_7092,N_4694,N_5747);
nor U7093 (N_7093,N_5883,N_5452);
xnor U7094 (N_7094,N_5486,N_5621);
or U7095 (N_7095,N_4653,N_5739);
and U7096 (N_7096,N_5365,N_5384);
and U7097 (N_7097,N_4680,N_5437);
nand U7098 (N_7098,N_4949,N_5557);
nand U7099 (N_7099,N_4635,N_4908);
xnor U7100 (N_7100,N_5793,N_4780);
and U7101 (N_7101,N_5475,N_5135);
nor U7102 (N_7102,N_5452,N_5865);
or U7103 (N_7103,N_5167,N_5212);
and U7104 (N_7104,N_5368,N_4613);
xor U7105 (N_7105,N_4799,N_4687);
nand U7106 (N_7106,N_4757,N_5190);
nand U7107 (N_7107,N_5997,N_5836);
nor U7108 (N_7108,N_5729,N_5466);
nand U7109 (N_7109,N_4532,N_5883);
nor U7110 (N_7110,N_5902,N_4632);
and U7111 (N_7111,N_4637,N_5333);
nand U7112 (N_7112,N_5914,N_4939);
and U7113 (N_7113,N_5447,N_5809);
nand U7114 (N_7114,N_5588,N_4885);
nand U7115 (N_7115,N_5830,N_4922);
and U7116 (N_7116,N_4703,N_5188);
and U7117 (N_7117,N_5997,N_5056);
nor U7118 (N_7118,N_5260,N_5820);
and U7119 (N_7119,N_4572,N_5024);
nand U7120 (N_7120,N_5536,N_5394);
nor U7121 (N_7121,N_5914,N_4650);
nor U7122 (N_7122,N_5542,N_5056);
and U7123 (N_7123,N_4828,N_5169);
or U7124 (N_7124,N_5350,N_5285);
or U7125 (N_7125,N_4819,N_5421);
nand U7126 (N_7126,N_5472,N_4592);
nor U7127 (N_7127,N_5509,N_4874);
or U7128 (N_7128,N_5532,N_5015);
nand U7129 (N_7129,N_5168,N_5478);
and U7130 (N_7130,N_5229,N_5549);
xnor U7131 (N_7131,N_4773,N_4995);
xnor U7132 (N_7132,N_5011,N_5451);
nor U7133 (N_7133,N_4926,N_5545);
or U7134 (N_7134,N_5981,N_5824);
or U7135 (N_7135,N_5219,N_5586);
nand U7136 (N_7136,N_5398,N_5142);
nand U7137 (N_7137,N_4685,N_4789);
xnor U7138 (N_7138,N_5595,N_5998);
and U7139 (N_7139,N_5466,N_4639);
xor U7140 (N_7140,N_5192,N_5896);
nand U7141 (N_7141,N_4725,N_4747);
or U7142 (N_7142,N_4800,N_4968);
or U7143 (N_7143,N_5559,N_5976);
or U7144 (N_7144,N_5560,N_5182);
nor U7145 (N_7145,N_5496,N_5148);
and U7146 (N_7146,N_4992,N_4646);
nand U7147 (N_7147,N_4597,N_5650);
nor U7148 (N_7148,N_5219,N_4848);
nor U7149 (N_7149,N_5644,N_4801);
or U7150 (N_7150,N_4740,N_4715);
nor U7151 (N_7151,N_4828,N_5088);
or U7152 (N_7152,N_5280,N_4604);
or U7153 (N_7153,N_4843,N_4681);
nand U7154 (N_7154,N_5702,N_4794);
and U7155 (N_7155,N_4559,N_5796);
xor U7156 (N_7156,N_4939,N_5800);
and U7157 (N_7157,N_5513,N_4901);
and U7158 (N_7158,N_5609,N_5805);
and U7159 (N_7159,N_5093,N_5372);
nor U7160 (N_7160,N_5459,N_5764);
and U7161 (N_7161,N_4596,N_5165);
nand U7162 (N_7162,N_4707,N_5068);
or U7163 (N_7163,N_5750,N_5838);
nand U7164 (N_7164,N_5572,N_4728);
and U7165 (N_7165,N_5578,N_5756);
or U7166 (N_7166,N_5370,N_5202);
xor U7167 (N_7167,N_4870,N_5377);
nand U7168 (N_7168,N_5129,N_5838);
and U7169 (N_7169,N_5498,N_4804);
nand U7170 (N_7170,N_5780,N_4758);
or U7171 (N_7171,N_4980,N_5076);
nor U7172 (N_7172,N_4901,N_5716);
and U7173 (N_7173,N_5919,N_5900);
and U7174 (N_7174,N_4624,N_5503);
or U7175 (N_7175,N_5586,N_4994);
or U7176 (N_7176,N_4925,N_5380);
xor U7177 (N_7177,N_5046,N_4963);
nand U7178 (N_7178,N_5611,N_4711);
nor U7179 (N_7179,N_4697,N_5940);
nor U7180 (N_7180,N_5974,N_5013);
nand U7181 (N_7181,N_5505,N_5172);
or U7182 (N_7182,N_5877,N_4621);
and U7183 (N_7183,N_5884,N_5118);
xnor U7184 (N_7184,N_5550,N_5767);
nand U7185 (N_7185,N_5375,N_4875);
or U7186 (N_7186,N_4632,N_5027);
nand U7187 (N_7187,N_5493,N_5161);
nand U7188 (N_7188,N_5382,N_5902);
and U7189 (N_7189,N_5246,N_5313);
xor U7190 (N_7190,N_5808,N_5008);
or U7191 (N_7191,N_5471,N_5059);
nand U7192 (N_7192,N_4579,N_5376);
or U7193 (N_7193,N_5029,N_5203);
or U7194 (N_7194,N_5325,N_5398);
xor U7195 (N_7195,N_4654,N_5024);
and U7196 (N_7196,N_5600,N_5902);
and U7197 (N_7197,N_5011,N_5505);
nor U7198 (N_7198,N_4932,N_5678);
nand U7199 (N_7199,N_5080,N_4986);
nor U7200 (N_7200,N_5046,N_5843);
nor U7201 (N_7201,N_4504,N_4520);
or U7202 (N_7202,N_4643,N_5779);
or U7203 (N_7203,N_5105,N_5243);
xnor U7204 (N_7204,N_5731,N_4725);
and U7205 (N_7205,N_5576,N_5997);
nand U7206 (N_7206,N_5596,N_4692);
nor U7207 (N_7207,N_5434,N_5460);
or U7208 (N_7208,N_5379,N_4721);
nor U7209 (N_7209,N_5836,N_5343);
nor U7210 (N_7210,N_4554,N_4851);
nand U7211 (N_7211,N_4747,N_5342);
xor U7212 (N_7212,N_4780,N_4831);
xnor U7213 (N_7213,N_5871,N_5098);
or U7214 (N_7214,N_4996,N_4575);
nor U7215 (N_7215,N_5535,N_5791);
nor U7216 (N_7216,N_4531,N_4771);
xnor U7217 (N_7217,N_5512,N_4704);
xor U7218 (N_7218,N_4891,N_4949);
and U7219 (N_7219,N_5409,N_5362);
nor U7220 (N_7220,N_5924,N_5419);
and U7221 (N_7221,N_5628,N_5991);
and U7222 (N_7222,N_4905,N_5275);
and U7223 (N_7223,N_5186,N_5005);
nand U7224 (N_7224,N_4536,N_4550);
and U7225 (N_7225,N_4900,N_4716);
or U7226 (N_7226,N_5468,N_5959);
or U7227 (N_7227,N_5712,N_5054);
nor U7228 (N_7228,N_4950,N_5490);
xor U7229 (N_7229,N_5870,N_4598);
and U7230 (N_7230,N_4528,N_4645);
nand U7231 (N_7231,N_5547,N_5914);
nand U7232 (N_7232,N_5413,N_5083);
xnor U7233 (N_7233,N_5078,N_5907);
or U7234 (N_7234,N_4619,N_5032);
and U7235 (N_7235,N_4964,N_5922);
nand U7236 (N_7236,N_5449,N_5465);
xor U7237 (N_7237,N_4662,N_4518);
and U7238 (N_7238,N_5526,N_5643);
or U7239 (N_7239,N_5303,N_4627);
or U7240 (N_7240,N_4655,N_4925);
nand U7241 (N_7241,N_5118,N_4712);
or U7242 (N_7242,N_5411,N_4574);
nor U7243 (N_7243,N_5619,N_5072);
or U7244 (N_7244,N_5890,N_5871);
nand U7245 (N_7245,N_5039,N_5787);
or U7246 (N_7246,N_5324,N_5600);
xnor U7247 (N_7247,N_5382,N_4742);
nor U7248 (N_7248,N_5526,N_5161);
nor U7249 (N_7249,N_4993,N_4956);
nand U7250 (N_7250,N_5233,N_4598);
nand U7251 (N_7251,N_5813,N_5845);
nand U7252 (N_7252,N_5018,N_5451);
or U7253 (N_7253,N_5398,N_5024);
and U7254 (N_7254,N_5107,N_5414);
nor U7255 (N_7255,N_4928,N_5943);
xnor U7256 (N_7256,N_4677,N_4514);
and U7257 (N_7257,N_4586,N_5573);
nand U7258 (N_7258,N_4649,N_5301);
and U7259 (N_7259,N_4618,N_4859);
xor U7260 (N_7260,N_5991,N_4681);
and U7261 (N_7261,N_5421,N_5033);
or U7262 (N_7262,N_4639,N_5710);
xor U7263 (N_7263,N_5030,N_4982);
xor U7264 (N_7264,N_5116,N_4778);
xor U7265 (N_7265,N_5871,N_5948);
or U7266 (N_7266,N_5076,N_5910);
and U7267 (N_7267,N_5373,N_4642);
nand U7268 (N_7268,N_5641,N_4645);
and U7269 (N_7269,N_4506,N_4681);
or U7270 (N_7270,N_5546,N_5289);
nand U7271 (N_7271,N_4967,N_5900);
nor U7272 (N_7272,N_5737,N_5069);
xor U7273 (N_7273,N_5972,N_5117);
nor U7274 (N_7274,N_5427,N_5071);
xnor U7275 (N_7275,N_5824,N_4851);
or U7276 (N_7276,N_5443,N_4920);
or U7277 (N_7277,N_5054,N_5686);
or U7278 (N_7278,N_4518,N_5040);
nor U7279 (N_7279,N_5423,N_4821);
and U7280 (N_7280,N_4932,N_5256);
nand U7281 (N_7281,N_4647,N_5013);
and U7282 (N_7282,N_4551,N_5830);
or U7283 (N_7283,N_5447,N_5358);
or U7284 (N_7284,N_5602,N_4773);
or U7285 (N_7285,N_5304,N_5462);
and U7286 (N_7286,N_5272,N_5346);
or U7287 (N_7287,N_5233,N_4854);
or U7288 (N_7288,N_5341,N_5378);
nor U7289 (N_7289,N_5843,N_4747);
xnor U7290 (N_7290,N_5162,N_5629);
and U7291 (N_7291,N_5817,N_5982);
and U7292 (N_7292,N_5499,N_5674);
nand U7293 (N_7293,N_5632,N_5338);
nor U7294 (N_7294,N_5835,N_5050);
xnor U7295 (N_7295,N_4598,N_5011);
nor U7296 (N_7296,N_5094,N_5332);
xnor U7297 (N_7297,N_5204,N_5350);
nand U7298 (N_7298,N_4758,N_5388);
xnor U7299 (N_7299,N_5643,N_5833);
and U7300 (N_7300,N_4976,N_5853);
and U7301 (N_7301,N_4645,N_5563);
and U7302 (N_7302,N_5534,N_5752);
and U7303 (N_7303,N_4700,N_5230);
and U7304 (N_7304,N_5337,N_4817);
and U7305 (N_7305,N_4960,N_4669);
nor U7306 (N_7306,N_4626,N_4672);
or U7307 (N_7307,N_4507,N_5028);
nor U7308 (N_7308,N_5442,N_5408);
xnor U7309 (N_7309,N_5036,N_5792);
xor U7310 (N_7310,N_5580,N_5213);
nor U7311 (N_7311,N_5006,N_5747);
and U7312 (N_7312,N_4670,N_5314);
and U7313 (N_7313,N_5162,N_4656);
and U7314 (N_7314,N_5532,N_4508);
and U7315 (N_7315,N_5223,N_5506);
or U7316 (N_7316,N_4638,N_5012);
or U7317 (N_7317,N_5354,N_4614);
nand U7318 (N_7318,N_4817,N_4522);
nand U7319 (N_7319,N_4889,N_4746);
xnor U7320 (N_7320,N_4702,N_5288);
nand U7321 (N_7321,N_5715,N_5064);
or U7322 (N_7322,N_5930,N_4819);
nor U7323 (N_7323,N_5804,N_5817);
nor U7324 (N_7324,N_5519,N_4966);
nand U7325 (N_7325,N_5990,N_4543);
nand U7326 (N_7326,N_4919,N_5713);
nor U7327 (N_7327,N_4998,N_5294);
nand U7328 (N_7328,N_5616,N_5283);
xor U7329 (N_7329,N_5592,N_5359);
or U7330 (N_7330,N_4858,N_5490);
nand U7331 (N_7331,N_4508,N_5978);
xnor U7332 (N_7332,N_5167,N_5257);
xnor U7333 (N_7333,N_5720,N_4568);
and U7334 (N_7334,N_5223,N_5617);
and U7335 (N_7335,N_5467,N_5296);
nor U7336 (N_7336,N_4984,N_5743);
or U7337 (N_7337,N_5041,N_5872);
and U7338 (N_7338,N_5400,N_5787);
xor U7339 (N_7339,N_5849,N_5148);
nor U7340 (N_7340,N_4532,N_4696);
nor U7341 (N_7341,N_5408,N_5356);
and U7342 (N_7342,N_4607,N_5075);
nand U7343 (N_7343,N_5813,N_5494);
xnor U7344 (N_7344,N_5945,N_4919);
nand U7345 (N_7345,N_5004,N_5600);
or U7346 (N_7346,N_4945,N_5461);
xnor U7347 (N_7347,N_4606,N_5273);
nand U7348 (N_7348,N_4940,N_5647);
and U7349 (N_7349,N_5482,N_4531);
nand U7350 (N_7350,N_5259,N_4508);
and U7351 (N_7351,N_5734,N_4803);
nor U7352 (N_7352,N_5703,N_4975);
and U7353 (N_7353,N_5962,N_5038);
nand U7354 (N_7354,N_5767,N_4798);
nand U7355 (N_7355,N_5625,N_5750);
nor U7356 (N_7356,N_5587,N_5459);
and U7357 (N_7357,N_5177,N_4680);
xnor U7358 (N_7358,N_5540,N_5175);
nand U7359 (N_7359,N_5618,N_5406);
and U7360 (N_7360,N_5892,N_5586);
nor U7361 (N_7361,N_4742,N_5077);
and U7362 (N_7362,N_5213,N_4548);
and U7363 (N_7363,N_5271,N_4959);
or U7364 (N_7364,N_5739,N_5005);
and U7365 (N_7365,N_4583,N_5766);
nor U7366 (N_7366,N_5910,N_5185);
or U7367 (N_7367,N_5702,N_4743);
and U7368 (N_7368,N_5543,N_4689);
nand U7369 (N_7369,N_5888,N_5453);
xnor U7370 (N_7370,N_5341,N_4764);
nand U7371 (N_7371,N_4522,N_4699);
nor U7372 (N_7372,N_5430,N_5571);
and U7373 (N_7373,N_5828,N_5626);
and U7374 (N_7374,N_4862,N_4874);
and U7375 (N_7375,N_4593,N_5316);
and U7376 (N_7376,N_5949,N_5784);
nor U7377 (N_7377,N_5256,N_5465);
nand U7378 (N_7378,N_4921,N_5294);
nand U7379 (N_7379,N_5988,N_4598);
and U7380 (N_7380,N_4652,N_5299);
and U7381 (N_7381,N_4566,N_5043);
and U7382 (N_7382,N_5889,N_4912);
or U7383 (N_7383,N_4782,N_5815);
nand U7384 (N_7384,N_4950,N_4764);
and U7385 (N_7385,N_5841,N_5605);
and U7386 (N_7386,N_5707,N_4864);
or U7387 (N_7387,N_5164,N_4960);
xor U7388 (N_7388,N_5697,N_5970);
nand U7389 (N_7389,N_5878,N_5430);
xor U7390 (N_7390,N_4974,N_5377);
and U7391 (N_7391,N_5958,N_4539);
or U7392 (N_7392,N_4806,N_5574);
xnor U7393 (N_7393,N_5215,N_4866);
nand U7394 (N_7394,N_4768,N_5179);
or U7395 (N_7395,N_5570,N_4697);
xor U7396 (N_7396,N_5750,N_5965);
and U7397 (N_7397,N_5104,N_4868);
nand U7398 (N_7398,N_5446,N_5298);
or U7399 (N_7399,N_5455,N_5438);
nor U7400 (N_7400,N_4845,N_5426);
and U7401 (N_7401,N_5324,N_5177);
and U7402 (N_7402,N_4532,N_4931);
nor U7403 (N_7403,N_5383,N_5900);
xor U7404 (N_7404,N_5452,N_5926);
and U7405 (N_7405,N_5351,N_4506);
or U7406 (N_7406,N_5383,N_5430);
nand U7407 (N_7407,N_5777,N_5918);
and U7408 (N_7408,N_4675,N_5766);
nand U7409 (N_7409,N_4904,N_5071);
and U7410 (N_7410,N_4595,N_5437);
and U7411 (N_7411,N_5902,N_4602);
and U7412 (N_7412,N_4959,N_4649);
xor U7413 (N_7413,N_4500,N_4917);
or U7414 (N_7414,N_4791,N_5553);
or U7415 (N_7415,N_5250,N_4920);
nor U7416 (N_7416,N_4894,N_5667);
nor U7417 (N_7417,N_5252,N_5192);
nor U7418 (N_7418,N_5978,N_5634);
xnor U7419 (N_7419,N_5523,N_5744);
nor U7420 (N_7420,N_5302,N_5803);
nand U7421 (N_7421,N_5817,N_5427);
and U7422 (N_7422,N_5139,N_4567);
xor U7423 (N_7423,N_5073,N_5024);
or U7424 (N_7424,N_5537,N_5869);
and U7425 (N_7425,N_5688,N_5318);
and U7426 (N_7426,N_4753,N_5211);
nand U7427 (N_7427,N_4521,N_4669);
or U7428 (N_7428,N_4554,N_4813);
nand U7429 (N_7429,N_5273,N_5942);
and U7430 (N_7430,N_4923,N_4579);
nand U7431 (N_7431,N_4715,N_5957);
nor U7432 (N_7432,N_5509,N_4741);
nor U7433 (N_7433,N_5198,N_4728);
or U7434 (N_7434,N_4549,N_5223);
or U7435 (N_7435,N_4572,N_5364);
and U7436 (N_7436,N_5696,N_4971);
xnor U7437 (N_7437,N_5384,N_5694);
nand U7438 (N_7438,N_5573,N_4710);
xnor U7439 (N_7439,N_4873,N_5243);
and U7440 (N_7440,N_5582,N_5579);
nand U7441 (N_7441,N_5626,N_4781);
nor U7442 (N_7442,N_5785,N_5846);
or U7443 (N_7443,N_4963,N_4676);
or U7444 (N_7444,N_5760,N_5939);
nor U7445 (N_7445,N_4694,N_4801);
nand U7446 (N_7446,N_5692,N_5491);
nand U7447 (N_7447,N_4947,N_5728);
nor U7448 (N_7448,N_5955,N_5508);
nand U7449 (N_7449,N_4930,N_4564);
nor U7450 (N_7450,N_5230,N_4751);
xor U7451 (N_7451,N_5744,N_4996);
or U7452 (N_7452,N_5935,N_5619);
nand U7453 (N_7453,N_5658,N_5547);
xor U7454 (N_7454,N_5867,N_4550);
nand U7455 (N_7455,N_4605,N_4987);
xnor U7456 (N_7456,N_5411,N_5068);
nand U7457 (N_7457,N_4719,N_4548);
and U7458 (N_7458,N_5469,N_5429);
or U7459 (N_7459,N_4880,N_5201);
or U7460 (N_7460,N_5291,N_4835);
nand U7461 (N_7461,N_5194,N_5739);
nand U7462 (N_7462,N_5233,N_5369);
nor U7463 (N_7463,N_5821,N_4934);
nand U7464 (N_7464,N_4761,N_5699);
xor U7465 (N_7465,N_4685,N_5305);
nand U7466 (N_7466,N_5138,N_5819);
and U7467 (N_7467,N_5683,N_4650);
and U7468 (N_7468,N_5715,N_5719);
nor U7469 (N_7469,N_4909,N_4507);
nor U7470 (N_7470,N_4559,N_5706);
xor U7471 (N_7471,N_5641,N_5191);
and U7472 (N_7472,N_4691,N_5009);
nand U7473 (N_7473,N_4788,N_5757);
or U7474 (N_7474,N_5936,N_4935);
or U7475 (N_7475,N_4607,N_5828);
nand U7476 (N_7476,N_4595,N_5278);
and U7477 (N_7477,N_4667,N_4975);
xor U7478 (N_7478,N_5029,N_4585);
or U7479 (N_7479,N_4751,N_5062);
nand U7480 (N_7480,N_5269,N_5550);
and U7481 (N_7481,N_5380,N_4702);
xnor U7482 (N_7482,N_5615,N_5094);
xnor U7483 (N_7483,N_4869,N_5518);
nor U7484 (N_7484,N_5487,N_4898);
xnor U7485 (N_7485,N_5403,N_5201);
xnor U7486 (N_7486,N_5779,N_5224);
nor U7487 (N_7487,N_5096,N_5525);
or U7488 (N_7488,N_4770,N_5970);
nand U7489 (N_7489,N_4517,N_4969);
or U7490 (N_7490,N_4970,N_4646);
nor U7491 (N_7491,N_4626,N_5924);
xnor U7492 (N_7492,N_4939,N_5480);
nand U7493 (N_7493,N_4672,N_5842);
or U7494 (N_7494,N_5247,N_5147);
nand U7495 (N_7495,N_5749,N_4736);
or U7496 (N_7496,N_5621,N_5126);
nand U7497 (N_7497,N_5333,N_5928);
nand U7498 (N_7498,N_5740,N_5447);
or U7499 (N_7499,N_5736,N_5764);
or U7500 (N_7500,N_6927,N_6415);
nor U7501 (N_7501,N_7138,N_7122);
or U7502 (N_7502,N_7297,N_6599);
nor U7503 (N_7503,N_6030,N_6162);
nor U7504 (N_7504,N_7086,N_7144);
or U7505 (N_7505,N_6330,N_6409);
and U7506 (N_7506,N_6410,N_6047);
or U7507 (N_7507,N_7043,N_6395);
and U7508 (N_7508,N_6314,N_7464);
nand U7509 (N_7509,N_6480,N_7084);
nor U7510 (N_7510,N_7188,N_6851);
nand U7511 (N_7511,N_6186,N_6348);
and U7512 (N_7512,N_6816,N_6973);
or U7513 (N_7513,N_6828,N_7382);
nor U7514 (N_7514,N_7284,N_6227);
or U7515 (N_7515,N_7456,N_7078);
nand U7516 (N_7516,N_6610,N_7291);
xnor U7517 (N_7517,N_6834,N_7332);
xor U7518 (N_7518,N_6905,N_6475);
nand U7519 (N_7519,N_7412,N_6858);
or U7520 (N_7520,N_6190,N_6678);
or U7521 (N_7521,N_6433,N_6767);
nor U7522 (N_7522,N_6950,N_6308);
and U7523 (N_7523,N_6142,N_6929);
xor U7524 (N_7524,N_6467,N_7421);
xnor U7525 (N_7525,N_7450,N_6645);
and U7526 (N_7526,N_6488,N_6800);
nand U7527 (N_7527,N_6920,N_6882);
or U7528 (N_7528,N_7157,N_6965);
nand U7529 (N_7529,N_6481,N_6210);
xnor U7530 (N_7530,N_6299,N_6473);
nand U7531 (N_7531,N_6984,N_6734);
nor U7532 (N_7532,N_6563,N_6655);
or U7533 (N_7533,N_6668,N_6328);
nor U7534 (N_7534,N_6810,N_7329);
xor U7535 (N_7535,N_6518,N_7311);
xnor U7536 (N_7536,N_6757,N_7184);
and U7537 (N_7537,N_6266,N_6750);
xnor U7538 (N_7538,N_6438,N_7040);
xor U7539 (N_7539,N_6795,N_6262);
xnor U7540 (N_7540,N_7098,N_6818);
nor U7541 (N_7541,N_6674,N_7136);
xnor U7542 (N_7542,N_7003,N_6303);
nand U7543 (N_7543,N_6201,N_6390);
xor U7544 (N_7544,N_6630,N_7493);
xor U7545 (N_7545,N_6222,N_6325);
nand U7546 (N_7546,N_6611,N_7015);
nor U7547 (N_7547,N_6393,N_7177);
xnor U7548 (N_7548,N_7099,N_7226);
xnor U7549 (N_7549,N_6284,N_7167);
and U7550 (N_7550,N_7025,N_6682);
or U7551 (N_7551,N_7163,N_7404);
xnor U7552 (N_7552,N_6392,N_7400);
nor U7553 (N_7553,N_6355,N_7439);
or U7554 (N_7554,N_6283,N_6461);
xnor U7555 (N_7555,N_6051,N_7055);
nand U7556 (N_7556,N_6896,N_6510);
or U7557 (N_7557,N_7491,N_6492);
xor U7558 (N_7558,N_6228,N_6379);
or U7559 (N_7559,N_6163,N_6145);
nor U7560 (N_7560,N_6629,N_7183);
xor U7561 (N_7561,N_6369,N_6136);
xnor U7562 (N_7562,N_6822,N_7394);
and U7563 (N_7563,N_6447,N_7125);
nand U7564 (N_7564,N_6759,N_6726);
or U7565 (N_7565,N_7186,N_7061);
and U7566 (N_7566,N_6383,N_6647);
and U7567 (N_7567,N_7073,N_6548);
nor U7568 (N_7568,N_6043,N_7492);
nor U7569 (N_7569,N_6496,N_6126);
nand U7570 (N_7570,N_6000,N_6663);
nor U7571 (N_7571,N_7093,N_7090);
xnor U7572 (N_7572,N_6368,N_6890);
xnor U7573 (N_7573,N_6309,N_6343);
or U7574 (N_7574,N_7216,N_6997);
and U7575 (N_7575,N_6034,N_6517);
or U7576 (N_7576,N_7010,N_7000);
and U7577 (N_7577,N_7262,N_7320);
nor U7578 (N_7578,N_6493,N_6741);
or U7579 (N_7579,N_7447,N_6195);
or U7580 (N_7580,N_7178,N_6707);
or U7581 (N_7581,N_6524,N_7198);
xnor U7582 (N_7582,N_6371,N_7156);
nor U7583 (N_7583,N_6298,N_6806);
xnor U7584 (N_7584,N_6280,N_7384);
xor U7585 (N_7585,N_7244,N_6605);
nor U7586 (N_7586,N_7154,N_6826);
nand U7587 (N_7587,N_6456,N_7294);
or U7588 (N_7588,N_7009,N_6646);
nand U7589 (N_7589,N_6585,N_6787);
or U7590 (N_7590,N_7429,N_7030);
and U7591 (N_7591,N_7190,N_6442);
nand U7592 (N_7592,N_6264,N_6792);
or U7593 (N_7593,N_7380,N_6286);
or U7594 (N_7594,N_7327,N_7295);
xor U7595 (N_7595,N_7426,N_6650);
and U7596 (N_7596,N_7259,N_7410);
xor U7597 (N_7597,N_6840,N_6260);
xnor U7598 (N_7598,N_6762,N_6515);
or U7599 (N_7599,N_6705,N_7109);
or U7600 (N_7600,N_6188,N_6231);
nand U7601 (N_7601,N_7155,N_6472);
or U7602 (N_7602,N_6704,N_6131);
and U7603 (N_7603,N_7418,N_6935);
or U7604 (N_7604,N_7103,N_6437);
nor U7605 (N_7605,N_6115,N_6909);
or U7606 (N_7606,N_6076,N_6633);
nand U7607 (N_7607,N_6577,N_6334);
nor U7608 (N_7608,N_6556,N_6153);
and U7609 (N_7609,N_7142,N_6995);
nor U7610 (N_7610,N_6638,N_7462);
and U7611 (N_7611,N_6578,N_7308);
nand U7612 (N_7612,N_6217,N_7046);
nor U7613 (N_7613,N_7200,N_7014);
nand U7614 (N_7614,N_6765,N_6823);
and U7615 (N_7615,N_6321,N_6275);
nand U7616 (N_7616,N_6972,N_7048);
and U7617 (N_7617,N_7466,N_7470);
nor U7618 (N_7618,N_6109,N_6513);
and U7619 (N_7619,N_6057,N_7346);
and U7620 (N_7620,N_6535,N_6135);
or U7621 (N_7621,N_7298,N_7207);
nor U7622 (N_7622,N_7067,N_7191);
nand U7623 (N_7623,N_6281,N_6593);
nor U7624 (N_7624,N_7088,N_6484);
or U7625 (N_7625,N_6466,N_6237);
xor U7626 (N_7626,N_7052,N_6620);
xnor U7627 (N_7627,N_7266,N_6970);
nor U7628 (N_7628,N_6170,N_7425);
nand U7629 (N_7629,N_6134,N_6656);
or U7630 (N_7630,N_6374,N_6534);
nand U7631 (N_7631,N_6315,N_7481);
nand U7632 (N_7632,N_6684,N_6127);
nand U7633 (N_7633,N_7045,N_7221);
and U7634 (N_7634,N_7085,N_6440);
and U7635 (N_7635,N_6837,N_7037);
nor U7636 (N_7636,N_7387,N_6066);
or U7637 (N_7637,N_6282,N_6717);
nand U7638 (N_7638,N_6602,N_7006);
nor U7639 (N_7639,N_7172,N_6336);
or U7640 (N_7640,N_6895,N_7457);
or U7641 (N_7641,N_6416,N_6868);
xor U7642 (N_7642,N_7119,N_6418);
xnor U7643 (N_7643,N_7406,N_6312);
xnor U7644 (N_7644,N_6317,N_6304);
or U7645 (N_7645,N_7047,N_7137);
nor U7646 (N_7646,N_6294,N_6412);
nor U7647 (N_7647,N_7145,N_6293);
or U7648 (N_7648,N_6016,N_6539);
nand U7649 (N_7649,N_6587,N_6154);
and U7650 (N_7650,N_7407,N_7101);
nand U7651 (N_7651,N_6872,N_7240);
and U7652 (N_7652,N_6009,N_6408);
xnor U7653 (N_7653,N_6221,N_6146);
and U7654 (N_7654,N_6226,N_6081);
or U7655 (N_7655,N_7293,N_7095);
and U7656 (N_7656,N_6071,N_7082);
nor U7657 (N_7657,N_6313,N_7299);
nor U7658 (N_7658,N_6983,N_7041);
nand U7659 (N_7659,N_7247,N_7401);
xnor U7660 (N_7660,N_6223,N_6160);
nor U7661 (N_7661,N_6627,N_6857);
nor U7662 (N_7662,N_6966,N_6653);
nand U7663 (N_7663,N_7202,N_6428);
and U7664 (N_7664,N_6786,N_6566);
xnor U7665 (N_7665,N_7397,N_7150);
nor U7666 (N_7666,N_6747,N_6485);
xnor U7667 (N_7667,N_7289,N_6665);
nor U7668 (N_7668,N_6628,N_6601);
and U7669 (N_7669,N_6659,N_6527);
or U7670 (N_7670,N_6967,N_6907);
nand U7671 (N_7671,N_7455,N_6797);
or U7672 (N_7672,N_6469,N_6088);
xor U7673 (N_7673,N_6660,N_6964);
and U7674 (N_7674,N_7353,N_6185);
or U7675 (N_7675,N_6434,N_6179);
nor U7676 (N_7676,N_6441,N_6006);
nand U7677 (N_7677,N_6214,N_6119);
nor U7678 (N_7678,N_6417,N_6435);
and U7679 (N_7679,N_6340,N_6094);
nand U7680 (N_7680,N_6411,N_6327);
xor U7681 (N_7681,N_6827,N_6498);
nor U7682 (N_7682,N_6565,N_7131);
nand U7683 (N_7683,N_6956,N_6528);
or U7684 (N_7684,N_6575,N_6087);
nor U7685 (N_7685,N_6132,N_7168);
xnor U7686 (N_7686,N_6452,N_7497);
xor U7687 (N_7687,N_6031,N_6853);
nor U7688 (N_7688,N_6039,N_7452);
xnor U7689 (N_7689,N_7104,N_7126);
xnor U7690 (N_7690,N_6265,N_7120);
xnor U7691 (N_7691,N_6380,N_6596);
nand U7692 (N_7692,N_6648,N_6960);
and U7693 (N_7693,N_6772,N_6864);
or U7694 (N_7694,N_6600,N_7166);
nand U7695 (N_7695,N_6919,N_6150);
nor U7696 (N_7696,N_6932,N_6497);
and U7697 (N_7697,N_7393,N_6893);
or U7698 (N_7698,N_6114,N_6061);
and U7699 (N_7699,N_7158,N_7370);
nor U7700 (N_7700,N_6885,N_6037);
nor U7701 (N_7701,N_6229,N_7049);
or U7702 (N_7702,N_7362,N_7013);
and U7703 (N_7703,N_6375,N_6451);
nand U7704 (N_7704,N_7286,N_6632);
and U7705 (N_7705,N_6789,N_6623);
and U7706 (N_7706,N_7449,N_6397);
xnor U7707 (N_7707,N_7129,N_6479);
or U7708 (N_7708,N_6486,N_7081);
nand U7709 (N_7709,N_6553,N_6886);
nand U7710 (N_7710,N_6879,N_6183);
and U7711 (N_7711,N_6576,N_6733);
or U7712 (N_7712,N_6306,N_6948);
or U7713 (N_7713,N_7375,N_6860);
nand U7714 (N_7714,N_6613,N_6062);
or U7715 (N_7715,N_6407,N_6875);
xor U7716 (N_7716,N_6233,N_6019);
xor U7717 (N_7717,N_7070,N_6844);
and U7718 (N_7718,N_6999,N_7110);
and U7719 (N_7719,N_6029,N_6590);
and U7720 (N_7720,N_6666,N_6508);
xor U7721 (N_7721,N_6918,N_7372);
nand U7722 (N_7722,N_6300,N_7253);
and U7723 (N_7723,N_7337,N_7420);
or U7724 (N_7724,N_6028,N_6873);
xor U7725 (N_7725,N_7258,N_6147);
nor U7726 (N_7726,N_6691,N_6606);
nor U7727 (N_7727,N_6715,N_6702);
xor U7728 (N_7728,N_6139,N_7066);
nand U7729 (N_7729,N_7152,N_6752);
nor U7730 (N_7730,N_7442,N_6544);
nand U7731 (N_7731,N_6156,N_6248);
nor U7732 (N_7732,N_6945,N_6838);
nand U7733 (N_7733,N_6813,N_6677);
and U7734 (N_7734,N_6570,N_6764);
and U7735 (N_7735,N_6808,N_6760);
nor U7736 (N_7736,N_7097,N_7318);
nor U7737 (N_7737,N_6211,N_6794);
nor U7738 (N_7738,N_6658,N_6982);
nor U7739 (N_7739,N_6523,N_6063);
and U7740 (N_7740,N_6198,N_6531);
xor U7741 (N_7741,N_6985,N_6084);
or U7742 (N_7742,N_7272,N_6654);
nor U7743 (N_7743,N_7121,N_7012);
nor U7744 (N_7744,N_6250,N_6520);
or U7745 (N_7745,N_6376,N_6345);
xor U7746 (N_7746,N_7193,N_6219);
nand U7747 (N_7747,N_6419,N_7091);
or U7748 (N_7748,N_7044,N_7023);
and U7749 (N_7749,N_6562,N_6096);
nor U7750 (N_7750,N_6100,N_6207);
nor U7751 (N_7751,N_6941,N_6450);
or U7752 (N_7752,N_7056,N_7367);
nand U7753 (N_7753,N_6561,N_6942);
nor U7754 (N_7754,N_7288,N_6507);
nand U7755 (N_7755,N_6884,N_6120);
nor U7756 (N_7756,N_7199,N_7227);
or U7757 (N_7757,N_7445,N_6268);
or U7758 (N_7758,N_7479,N_6270);
and U7759 (N_7759,N_6790,N_6050);
or U7760 (N_7760,N_6846,N_6400);
nor U7761 (N_7761,N_6737,N_6778);
and U7762 (N_7762,N_7241,N_6607);
and U7763 (N_7763,N_6706,N_6987);
and U7764 (N_7764,N_6898,N_7132);
nor U7765 (N_7765,N_6644,N_7399);
nand U7766 (N_7766,N_7151,N_6391);
nor U7767 (N_7767,N_7135,N_6549);
xnor U7768 (N_7768,N_6912,N_6316);
xnor U7769 (N_7769,N_6436,N_6954);
or U7770 (N_7770,N_6098,N_6996);
nand U7771 (N_7771,N_7143,N_7275);
xor U7772 (N_7772,N_6238,N_6962);
xor U7773 (N_7773,N_6651,N_7064);
nor U7774 (N_7774,N_7279,N_6239);
and U7775 (N_7775,N_7035,N_7225);
nand U7776 (N_7776,N_6568,N_7027);
or U7777 (N_7777,N_6708,N_6140);
and U7778 (N_7778,N_6110,N_6724);
or U7779 (N_7779,N_6526,N_6722);
and U7780 (N_7780,N_7222,N_6187);
xnor U7781 (N_7781,N_6637,N_7063);
nand U7782 (N_7782,N_6107,N_7071);
xnor U7783 (N_7783,N_6197,N_6487);
nand U7784 (N_7784,N_7274,N_6193);
nand U7785 (N_7785,N_6149,N_6641);
nor U7786 (N_7786,N_7499,N_7260);
nor U7787 (N_7787,N_6326,N_6113);
nor U7788 (N_7788,N_7252,N_6713);
or U7789 (N_7789,N_7153,N_6387);
nor U7790 (N_7790,N_7039,N_6324);
nand U7791 (N_7791,N_7366,N_6020);
nor U7792 (N_7792,N_6425,N_6928);
and U7793 (N_7793,N_7194,N_6514);
nand U7794 (N_7794,N_6274,N_6449);
xnor U7795 (N_7795,N_6843,N_6247);
nand U7796 (N_7796,N_6199,N_6471);
or U7797 (N_7797,N_6791,N_6554);
nor U7798 (N_7798,N_6196,N_6070);
and U7799 (N_7799,N_6095,N_6992);
nand U7800 (N_7800,N_6617,N_7278);
nor U7801 (N_7801,N_6824,N_6732);
nor U7802 (N_7802,N_6249,N_6571);
xnor U7803 (N_7803,N_6855,N_6714);
nor U7804 (N_7804,N_6405,N_6835);
and U7805 (N_7805,N_6728,N_6253);
nand U7806 (N_7806,N_6924,N_7360);
or U7807 (N_7807,N_6008,N_7422);
nor U7808 (N_7808,N_6333,N_7133);
nor U7809 (N_7809,N_7377,N_6118);
nand U7810 (N_7810,N_7127,N_7001);
or U7811 (N_7811,N_6742,N_6738);
nand U7812 (N_7812,N_6761,N_7267);
or U7813 (N_7813,N_6968,N_6547);
or U7814 (N_7814,N_6463,N_7160);
xor U7815 (N_7815,N_7218,N_6673);
or U7816 (N_7816,N_7114,N_7363);
or U7817 (N_7817,N_7165,N_6955);
nor U7818 (N_7818,N_7182,N_6168);
nor U7819 (N_7819,N_6703,N_6460);
and U7820 (N_7820,N_7077,N_6529);
xnor U7821 (N_7821,N_6388,N_6502);
or U7822 (N_7822,N_7074,N_6216);
nor U7823 (N_7823,N_7437,N_7477);
xor U7824 (N_7824,N_6494,N_6205);
xor U7825 (N_7825,N_6427,N_6358);
nand U7826 (N_7826,N_6719,N_6279);
nand U7827 (N_7827,N_7196,N_6811);
nor U7828 (N_7828,N_6181,N_6122);
or U7829 (N_7829,N_6065,N_6963);
and U7830 (N_7830,N_6692,N_7148);
or U7831 (N_7831,N_6432,N_7321);
nand U7832 (N_7832,N_7220,N_7029);
and U7833 (N_7833,N_7238,N_6086);
nor U7834 (N_7834,N_7460,N_6642);
xnor U7835 (N_7835,N_6116,N_6335);
nand U7836 (N_7836,N_6230,N_6667);
nand U7837 (N_7837,N_6064,N_7303);
and U7838 (N_7838,N_7036,N_6586);
or U7839 (N_7839,N_7304,N_7263);
or U7840 (N_7840,N_7391,N_7228);
and U7841 (N_7841,N_6777,N_6033);
or U7842 (N_7842,N_6338,N_6915);
nand U7843 (N_7843,N_6783,N_6579);
and U7844 (N_7844,N_6241,N_6874);
or U7845 (N_7845,N_6906,N_6232);
or U7846 (N_7846,N_6871,N_6079);
nor U7847 (N_7847,N_7356,N_6117);
xor U7848 (N_7848,N_6297,N_6091);
nor U7849 (N_7849,N_6640,N_6774);
and U7850 (N_7850,N_6903,N_6049);
nor U7851 (N_7851,N_6194,N_6024);
and U7852 (N_7852,N_6491,N_6277);
nand U7853 (N_7853,N_6842,N_7096);
xnor U7854 (N_7854,N_7433,N_7038);
and U7855 (N_7855,N_7487,N_7239);
and U7856 (N_7856,N_6060,N_6075);
and U7857 (N_7857,N_7306,N_6621);
nor U7858 (N_7858,N_6121,N_6725);
and U7859 (N_7859,N_6421,N_6781);
nand U7860 (N_7860,N_6396,N_7444);
nor U7861 (N_7861,N_6989,N_7243);
or U7862 (N_7862,N_7374,N_6836);
nand U7863 (N_7863,N_7232,N_6311);
or U7864 (N_7864,N_6423,N_7484);
nand U7865 (N_7865,N_6189,N_6657);
and U7866 (N_7866,N_7409,N_6543);
and U7867 (N_7867,N_7416,N_6093);
or U7868 (N_7868,N_7250,N_6910);
nand U7869 (N_7869,N_6490,N_6360);
xnor U7870 (N_7870,N_7358,N_6603);
nand U7871 (N_7871,N_7364,N_6739);
xnor U7872 (N_7872,N_6511,N_7195);
or U7873 (N_7873,N_6242,N_7371);
nor U7874 (N_7874,N_7476,N_6749);
and U7875 (N_7875,N_6468,N_6779);
nand U7876 (N_7876,N_6943,N_7341);
and U7877 (N_7877,N_7310,N_7435);
nor U7878 (N_7878,N_7231,N_6384);
or U7879 (N_7879,N_7234,N_6537);
or U7880 (N_7880,N_7201,N_7495);
and U7881 (N_7881,N_7105,N_7330);
xnor U7882 (N_7882,N_6448,N_7065);
xnor U7883 (N_7883,N_6977,N_6404);
nand U7884 (N_7884,N_6372,N_6164);
or U7885 (N_7885,N_7348,N_6574);
or U7886 (N_7886,N_6103,N_7254);
and U7887 (N_7887,N_6830,N_7256);
and U7888 (N_7888,N_6730,N_7233);
and U7889 (N_7889,N_6723,N_6720);
nand U7890 (N_7890,N_7345,N_6295);
or U7891 (N_7891,N_6124,N_7463);
nand U7892 (N_7892,N_6445,N_7032);
nand U7893 (N_7893,N_7331,N_7474);
nor U7894 (N_7894,N_6097,N_7428);
nand U7895 (N_7895,N_7203,N_6540);
nor U7896 (N_7896,N_6257,N_7205);
or U7897 (N_7897,N_6917,N_6986);
and U7898 (N_7898,N_7402,N_6624);
nand U7899 (N_7899,N_7079,N_6814);
nor U7900 (N_7900,N_7209,N_6625);
xnor U7901 (N_7901,N_6478,N_6676);
xor U7902 (N_7902,N_6220,N_6329);
or U7903 (N_7903,N_7057,N_7296);
and U7904 (N_7904,N_6133,N_6042);
nand U7905 (N_7905,N_6353,N_6015);
and U7906 (N_7906,N_6026,N_6569);
and U7907 (N_7907,N_7271,N_6359);
xor U7908 (N_7908,N_7042,N_7002);
and U7909 (N_7909,N_6729,N_6595);
and U7910 (N_7910,N_7219,N_7316);
and U7911 (N_7911,N_7257,N_6696);
nor U7912 (N_7912,N_6208,N_6204);
or U7913 (N_7913,N_6564,N_6690);
xor U7914 (N_7914,N_6542,N_6011);
nor U7915 (N_7915,N_6850,N_6519);
and U7916 (N_7916,N_6994,N_7312);
xnor U7917 (N_7917,N_6947,N_6092);
xnor U7918 (N_7918,N_6591,N_7223);
nor U7919 (N_7919,N_6272,N_6038);
nand U7920 (N_7920,N_7072,N_6344);
or U7921 (N_7921,N_7381,N_6495);
nand U7922 (N_7922,N_7368,N_6670);
nor U7923 (N_7923,N_7060,N_6784);
nand U7924 (N_7924,N_7488,N_6716);
nand U7925 (N_7925,N_7255,N_6863);
nand U7926 (N_7926,N_6809,N_6269);
and U7927 (N_7927,N_6971,N_6618);
and U7928 (N_7928,N_6206,N_6793);
or U7929 (N_7929,N_7408,N_6341);
xor U7930 (N_7930,N_7212,N_6856);
nor U7931 (N_7931,N_7436,N_7379);
nand U7932 (N_7932,N_7192,N_7403);
or U7933 (N_7933,N_6399,N_6414);
and U7934 (N_7934,N_6815,N_7319);
and U7935 (N_7935,N_6652,N_6111);
and U7936 (N_7936,N_7351,N_7111);
nand U7937 (N_7937,N_6273,N_7117);
nor U7938 (N_7938,N_6981,N_6536);
xnor U7939 (N_7939,N_6776,N_7051);
and U7940 (N_7940,N_7485,N_6161);
xor U7941 (N_7941,N_7369,N_6572);
nand U7942 (N_7942,N_6054,N_6259);
and U7943 (N_7943,N_6718,N_7069);
and U7944 (N_7944,N_6177,N_6010);
nor U7945 (N_7945,N_7432,N_7058);
nor U7946 (N_7946,N_6735,N_6916);
and U7947 (N_7947,N_6243,N_6128);
nor U7948 (N_7948,N_7235,N_7140);
nor U7949 (N_7949,N_7115,N_7080);
and U7950 (N_7950,N_6788,N_7336);
or U7951 (N_7951,N_6209,N_6056);
xnor U7952 (N_7952,N_7438,N_7313);
nor U7953 (N_7953,N_7325,N_6158);
and U7954 (N_7954,N_6366,N_6686);
nand U7955 (N_7955,N_7324,N_7333);
nand U7956 (N_7956,N_6278,N_6256);
nand U7957 (N_7957,N_6608,N_7472);
or U7958 (N_7958,N_6155,N_7017);
xnor U7959 (N_7959,N_6083,N_7283);
and U7960 (N_7960,N_6455,N_7378);
or U7961 (N_7961,N_6255,N_6758);
or U7962 (N_7962,N_6959,N_7011);
nor U7963 (N_7963,N_6426,N_6018);
nand U7964 (N_7964,N_6148,N_6365);
nor U7965 (N_7965,N_6501,N_6271);
xnor U7966 (N_7966,N_6891,N_7076);
and U7967 (N_7967,N_7280,N_6699);
xor U7968 (N_7968,N_7197,N_6377);
or U7969 (N_7969,N_6499,N_6894);
nor U7970 (N_7970,N_7008,N_7176);
and U7971 (N_7971,N_7031,N_7467);
nand U7972 (N_7972,N_7419,N_6869);
nand U7973 (N_7973,N_6887,N_6058);
or U7974 (N_7974,N_6934,N_7465);
xnor U7975 (N_7975,N_7392,N_7185);
nand U7976 (N_7976,N_7159,N_6429);
and U7977 (N_7977,N_6143,N_7423);
xor U7978 (N_7978,N_6001,N_7498);
nand U7979 (N_7979,N_6635,N_7034);
and U7980 (N_7980,N_6512,N_7092);
and U7981 (N_7981,N_6939,N_7141);
nor U7982 (N_7982,N_6339,N_7482);
xnor U7983 (N_7983,N_6978,N_6751);
or U7984 (N_7984,N_6180,N_6626);
or U7985 (N_7985,N_7305,N_7128);
xor U7986 (N_7986,N_6483,N_6953);
and U7987 (N_7987,N_7075,N_6482);
xnor U7988 (N_7988,N_7446,N_6930);
nor U7989 (N_7989,N_6212,N_7026);
or U7990 (N_7990,N_6675,N_7230);
and U7991 (N_7991,N_7451,N_6922);
nor U7992 (N_7992,N_7453,N_6218);
nand U7993 (N_7993,N_7471,N_6251);
and U7994 (N_7994,N_7405,N_6541);
or U7995 (N_7995,N_7123,N_6235);
or U7996 (N_7996,N_6246,N_6521);
xor U7997 (N_7997,N_7189,N_6866);
or U7998 (N_7998,N_7338,N_7350);
xnor U7999 (N_7999,N_6245,N_6546);
nor U8000 (N_8000,N_7208,N_6763);
nand U8001 (N_8001,N_7007,N_6036);
or U8002 (N_8002,N_6477,N_7248);
nor U8003 (N_8003,N_6768,N_6055);
nor U8004 (N_8004,N_6166,N_6394);
xor U8005 (N_8005,N_7113,N_6865);
nand U8006 (N_8006,N_6545,N_7089);
and U8007 (N_8007,N_6267,N_6263);
nand U8008 (N_8008,N_6649,N_7292);
and U8009 (N_8009,N_7287,N_7175);
xor U8010 (N_8010,N_6588,N_7424);
nand U8011 (N_8011,N_6004,N_7483);
nor U8012 (N_8012,N_7411,N_6288);
xnor U8013 (N_8013,N_6883,N_6080);
xnor U8014 (N_8014,N_6402,N_6662);
or U8015 (N_8015,N_6619,N_6700);
or U8016 (N_8016,N_6302,N_6462);
nor U8017 (N_8017,N_6305,N_7314);
and U8018 (N_8018,N_7343,N_6701);
or U8019 (N_8019,N_7359,N_6581);
and U8020 (N_8020,N_6059,N_6240);
nor U8021 (N_8021,N_6852,N_6573);
xor U8022 (N_8022,N_7134,N_6748);
xor U8023 (N_8023,N_7213,N_6862);
nand U8024 (N_8024,N_7116,N_6839);
nor U8025 (N_8025,N_6592,N_6077);
nor U8026 (N_8026,N_6378,N_6078);
xor U8027 (N_8027,N_6500,N_6443);
or U8028 (N_8028,N_6192,N_7217);
nand U8029 (N_8029,N_7398,N_6474);
nor U8030 (N_8030,N_6354,N_6252);
or U8031 (N_8031,N_6693,N_7326);
and U8032 (N_8032,N_6307,N_6988);
nor U8033 (N_8033,N_6867,N_6812);
xnor U8034 (N_8034,N_6291,N_6357);
nand U8035 (N_8035,N_6046,N_7430);
and U8036 (N_8036,N_6234,N_7229);
xor U8037 (N_8037,N_7443,N_7242);
and U8038 (N_8038,N_6385,N_6332);
xnor U8039 (N_8039,N_6616,N_6754);
nand U8040 (N_8040,N_6925,N_6301);
or U8041 (N_8041,N_7340,N_6173);
xnor U8042 (N_8042,N_6597,N_6072);
nor U8043 (N_8043,N_7161,N_6957);
nor U8044 (N_8044,N_6848,N_6151);
xnor U8045 (N_8045,N_6053,N_6174);
xor U8046 (N_8046,N_6598,N_7022);
and U8047 (N_8047,N_6191,N_6007);
nor U8048 (N_8048,N_6615,N_7162);
or U8049 (N_8049,N_6224,N_6913);
nand U8050 (N_8050,N_6990,N_6171);
xor U8051 (N_8051,N_6847,N_7224);
and U8052 (N_8052,N_6525,N_7458);
or U8053 (N_8053,N_6825,N_6203);
nand U8054 (N_8054,N_6952,N_6176);
nand U8055 (N_8055,N_6877,N_6458);
xnor U8056 (N_8056,N_6604,N_6337);
nor U8057 (N_8057,N_7335,N_6744);
or U8058 (N_8058,N_6631,N_6319);
nand U8059 (N_8059,N_6108,N_7431);
xnor U8060 (N_8060,N_6144,N_6555);
nor U8061 (N_8061,N_6090,N_7277);
and U8062 (N_8062,N_6773,N_6424);
and U8063 (N_8063,N_7469,N_7094);
xnor U8064 (N_8064,N_6841,N_7174);
nor U8065 (N_8065,N_6202,N_6200);
nand U8066 (N_8066,N_6664,N_7468);
xnor U8067 (N_8067,N_6861,N_7434);
nor U8068 (N_8068,N_7454,N_6557);
or U8069 (N_8069,N_6589,N_6516);
or U8070 (N_8070,N_6711,N_6362);
or U8071 (N_8071,N_7461,N_6041);
and U8072 (N_8072,N_6756,N_6636);
and U8073 (N_8073,N_7342,N_6323);
xor U8074 (N_8074,N_6859,N_7373);
nand U8075 (N_8075,N_7300,N_7206);
or U8076 (N_8076,N_6048,N_6745);
or U8077 (N_8077,N_6005,N_6082);
xor U8078 (N_8078,N_6331,N_6112);
nand U8079 (N_8079,N_6476,N_7269);
xnor U8080 (N_8080,N_6612,N_6138);
nand U8081 (N_8081,N_6782,N_7285);
nand U8082 (N_8082,N_6911,N_6254);
nand U8083 (N_8083,N_7204,N_7211);
nor U8084 (N_8084,N_7315,N_7496);
nor U8085 (N_8085,N_7268,N_6032);
nor U8086 (N_8086,N_7261,N_6899);
nor U8087 (N_8087,N_6904,N_7339);
xnor U8088 (N_8088,N_6413,N_6261);
or U8089 (N_8089,N_7489,N_6382);
nand U8090 (N_8090,N_6805,N_6225);
nor U8091 (N_8091,N_6430,N_6398);
xor U8092 (N_8092,N_7146,N_7413);
nand U8093 (N_8093,N_6689,N_6125);
nand U8094 (N_8094,N_6923,N_6558);
nor U8095 (N_8095,N_6634,N_6946);
and U8096 (N_8096,N_7028,N_6672);
xnor U8097 (N_8097,N_6023,N_7016);
xnor U8098 (N_8098,N_6914,N_6067);
xor U8099 (N_8099,N_7389,N_6594);
or U8100 (N_8100,N_7365,N_6178);
and U8101 (N_8101,N_7301,N_6351);
nor U8102 (N_8102,N_7118,N_6580);
nand U8103 (N_8103,N_6785,N_6137);
xor U8104 (N_8104,N_7290,N_7130);
nor U8105 (N_8105,N_6439,N_6969);
or U8106 (N_8106,N_6373,N_7440);
nand U8107 (N_8107,N_6694,N_6958);
and U8108 (N_8108,N_6364,N_6532);
nor U8109 (N_8109,N_6892,N_6802);
xor U8110 (N_8110,N_6453,N_6215);
nor U8111 (N_8111,N_7273,N_6993);
nand U8112 (N_8112,N_7270,N_6184);
and U8113 (N_8113,N_6731,N_6736);
and U8114 (N_8114,N_7087,N_6165);
or U8115 (N_8115,N_6287,N_7282);
and U8116 (N_8116,N_7024,N_6003);
and U8117 (N_8117,N_7494,N_6454);
and U8118 (N_8118,N_6289,N_6849);
nor U8119 (N_8119,N_6504,N_7033);
nand U8120 (N_8120,N_6991,N_6014);
nor U8121 (N_8121,N_6401,N_6175);
xnor U8122 (N_8122,N_6926,N_6721);
or U8123 (N_8123,N_6213,N_6901);
nand U8124 (N_8124,N_6807,N_6817);
and U8125 (N_8125,N_6102,N_7344);
nor U8126 (N_8126,N_7139,N_6908);
nand U8127 (N_8127,N_7354,N_6074);
xnor U8128 (N_8128,N_6017,N_6780);
or U8129 (N_8129,N_7386,N_7361);
xor U8130 (N_8130,N_6182,N_7018);
and U8131 (N_8131,N_6888,N_6167);
nor U8132 (N_8132,N_7417,N_7427);
and U8133 (N_8133,N_6582,N_7265);
xnor U8134 (N_8134,N_7237,N_6880);
or U8135 (N_8135,N_7328,N_7053);
xnor U8136 (N_8136,N_6157,N_7414);
or U8137 (N_8137,N_7050,N_6900);
and U8138 (N_8138,N_6104,N_7054);
or U8139 (N_8139,N_7281,N_6609);
xnor U8140 (N_8140,N_6044,N_6974);
xnor U8141 (N_8141,N_6290,N_6129);
or U8142 (N_8142,N_6870,N_6370);
nor U8143 (N_8143,N_6979,N_7251);
nor U8144 (N_8144,N_6099,N_6422);
or U8145 (N_8145,N_6236,N_7180);
xnor U8146 (N_8146,N_6975,N_7147);
nor U8147 (N_8147,N_7215,N_7083);
nand U8148 (N_8148,N_6322,N_6889);
and U8149 (N_8149,N_6296,N_6669);
and U8150 (N_8150,N_6320,N_6420);
nor U8151 (N_8151,N_7309,N_6951);
and U8152 (N_8152,N_7210,N_7021);
nor U8153 (N_8153,N_6258,N_6639);
xnor U8154 (N_8154,N_6444,N_6998);
xnor U8155 (N_8155,N_7169,N_6680);
xnor U8156 (N_8156,N_6069,N_7390);
xnor U8157 (N_8157,N_6350,N_6538);
nand U8158 (N_8158,N_6819,N_6881);
nand U8159 (N_8159,N_6552,N_7068);
nor U8160 (N_8160,N_6933,N_6876);
nor U8161 (N_8161,N_6470,N_6035);
nand U8162 (N_8162,N_6386,N_6746);
nand U8163 (N_8163,N_7173,N_7106);
nor U8164 (N_8164,N_7181,N_6940);
or U8165 (N_8165,N_7334,N_7490);
nand U8166 (N_8166,N_6803,N_6446);
xnor U8167 (N_8167,N_6550,N_6431);
and U8168 (N_8168,N_6346,N_6832);
and U8169 (N_8169,N_6796,N_7100);
nor U8170 (N_8170,N_6347,N_6687);
nor U8171 (N_8171,N_6698,N_6829);
nor U8172 (N_8172,N_6938,N_6085);
and U8173 (N_8173,N_7395,N_6766);
xor U8174 (N_8174,N_7187,N_7478);
xnor U8175 (N_8175,N_6695,N_6551);
or U8176 (N_8176,N_7062,N_6949);
xnor U8177 (N_8177,N_6021,N_7322);
nand U8178 (N_8178,N_7164,N_6614);
nor U8179 (N_8179,N_6002,N_7102);
xnor U8180 (N_8180,N_7352,N_7124);
nand U8181 (N_8181,N_7149,N_6921);
nand U8182 (N_8182,N_6740,N_7317);
nor U8183 (N_8183,N_6318,N_6878);
or U8184 (N_8184,N_6743,N_6013);
nand U8185 (N_8185,N_6244,N_6172);
nand U8186 (N_8186,N_6152,N_6770);
xor U8187 (N_8187,N_6105,N_7179);
or U8188 (N_8188,N_6902,N_6381);
xor U8189 (N_8189,N_6403,N_7347);
xor U8190 (N_8190,N_6276,N_6688);
xor U8191 (N_8191,N_7307,N_6169);
xor U8192 (N_8192,N_6685,N_6798);
xor U8193 (N_8193,N_7480,N_6406);
or U8194 (N_8194,N_6073,N_6101);
or U8195 (N_8195,N_6804,N_6709);
nand U8196 (N_8196,N_6068,N_6799);
and U8197 (N_8197,N_6697,N_6489);
xnor U8198 (N_8198,N_6671,N_6292);
and U8199 (N_8199,N_7107,N_6976);
xor U8200 (N_8200,N_6683,N_6755);
or U8201 (N_8201,N_7004,N_6045);
nand U8202 (N_8202,N_6775,N_6089);
or U8203 (N_8203,N_7388,N_7245);
nand U8204 (N_8204,N_6821,N_6560);
and U8205 (N_8205,N_6712,N_6285);
nand U8206 (N_8206,N_6342,N_6464);
or U8207 (N_8207,N_6931,N_6025);
nand U8208 (N_8208,N_6936,N_6854);
or U8209 (N_8209,N_6141,N_6052);
xor U8210 (N_8210,N_6961,N_6389);
and U8211 (N_8211,N_7349,N_7376);
and U8212 (N_8212,N_6980,N_6681);
and U8213 (N_8213,N_6457,N_6361);
nand U8214 (N_8214,N_6130,N_7448);
nor U8215 (N_8215,N_7473,N_7005);
nand U8216 (N_8216,N_6506,N_7415);
or U8217 (N_8217,N_7459,N_6833);
or U8218 (N_8218,N_6459,N_7112);
nand U8219 (N_8219,N_6567,N_7396);
nor U8220 (N_8220,N_6159,N_6465);
and U8221 (N_8221,N_6022,N_6522);
or U8222 (N_8222,N_6897,N_6727);
or U8223 (N_8223,N_7276,N_7019);
or U8224 (N_8224,N_7355,N_6363);
and U8225 (N_8225,N_7170,N_7059);
nand U8226 (N_8226,N_6027,N_6349);
or U8227 (N_8227,N_6559,N_6820);
and U8228 (N_8228,N_6352,N_7246);
and U8229 (N_8229,N_6310,N_6012);
or U8230 (N_8230,N_7441,N_6509);
xor U8231 (N_8231,N_6944,N_6584);
and U8232 (N_8232,N_7249,N_7385);
nand U8233 (N_8233,N_7171,N_7020);
and U8234 (N_8234,N_6845,N_6123);
and U8235 (N_8235,N_7323,N_6533);
nand U8236 (N_8236,N_7236,N_6583);
and U8237 (N_8237,N_6622,N_6937);
nor U8238 (N_8238,N_7302,N_6356);
nor U8239 (N_8239,N_7264,N_7357);
nor U8240 (N_8240,N_7486,N_6367);
xor U8241 (N_8241,N_7475,N_6643);
nor U8242 (N_8242,N_6753,N_6106);
and U8243 (N_8243,N_6661,N_6710);
nand U8244 (N_8244,N_6040,N_6769);
or U8245 (N_8245,N_6530,N_7108);
nor U8246 (N_8246,N_7383,N_6831);
or U8247 (N_8247,N_6505,N_7214);
nor U8248 (N_8248,N_6771,N_6801);
or U8249 (N_8249,N_6679,N_6503);
nor U8250 (N_8250,N_7368,N_7161);
xnor U8251 (N_8251,N_6123,N_7087);
xnor U8252 (N_8252,N_7107,N_6679);
xor U8253 (N_8253,N_7456,N_6622);
nor U8254 (N_8254,N_6176,N_7042);
xnor U8255 (N_8255,N_6216,N_6640);
nor U8256 (N_8256,N_6597,N_6378);
nand U8257 (N_8257,N_6590,N_7287);
or U8258 (N_8258,N_7481,N_7054);
xor U8259 (N_8259,N_6798,N_7108);
nand U8260 (N_8260,N_6964,N_6231);
nand U8261 (N_8261,N_6394,N_7448);
and U8262 (N_8262,N_6585,N_6373);
nand U8263 (N_8263,N_6189,N_6832);
nand U8264 (N_8264,N_7494,N_6080);
nor U8265 (N_8265,N_6733,N_6404);
nor U8266 (N_8266,N_6408,N_6728);
and U8267 (N_8267,N_6836,N_6502);
and U8268 (N_8268,N_6052,N_6404);
or U8269 (N_8269,N_7347,N_6369);
and U8270 (N_8270,N_7072,N_6656);
nand U8271 (N_8271,N_6820,N_7122);
nor U8272 (N_8272,N_6978,N_6320);
and U8273 (N_8273,N_7243,N_7430);
or U8274 (N_8274,N_7261,N_6677);
or U8275 (N_8275,N_7240,N_6328);
xor U8276 (N_8276,N_7318,N_6112);
nor U8277 (N_8277,N_6393,N_7392);
or U8278 (N_8278,N_6941,N_7098);
or U8279 (N_8279,N_7335,N_7030);
xnor U8280 (N_8280,N_6740,N_6951);
or U8281 (N_8281,N_7385,N_7466);
and U8282 (N_8282,N_6916,N_6661);
and U8283 (N_8283,N_6864,N_7138);
or U8284 (N_8284,N_6069,N_7405);
and U8285 (N_8285,N_6355,N_6466);
xnor U8286 (N_8286,N_6003,N_6913);
and U8287 (N_8287,N_6672,N_7152);
nand U8288 (N_8288,N_7377,N_7410);
and U8289 (N_8289,N_6451,N_6753);
nand U8290 (N_8290,N_6089,N_7257);
nor U8291 (N_8291,N_6696,N_6531);
or U8292 (N_8292,N_6516,N_6156);
xor U8293 (N_8293,N_7142,N_6922);
nand U8294 (N_8294,N_6440,N_7027);
or U8295 (N_8295,N_6516,N_7491);
nand U8296 (N_8296,N_7212,N_6638);
nor U8297 (N_8297,N_6139,N_6654);
and U8298 (N_8298,N_6303,N_6332);
xor U8299 (N_8299,N_7393,N_6270);
nand U8300 (N_8300,N_6821,N_6399);
nor U8301 (N_8301,N_6523,N_6234);
xor U8302 (N_8302,N_6836,N_6819);
or U8303 (N_8303,N_6427,N_6095);
xor U8304 (N_8304,N_7152,N_7153);
nand U8305 (N_8305,N_6252,N_7489);
nand U8306 (N_8306,N_6147,N_7067);
nor U8307 (N_8307,N_7024,N_6713);
xnor U8308 (N_8308,N_6349,N_7444);
xor U8309 (N_8309,N_6329,N_6258);
and U8310 (N_8310,N_6930,N_7032);
or U8311 (N_8311,N_6368,N_6899);
and U8312 (N_8312,N_6577,N_7456);
or U8313 (N_8313,N_6144,N_6285);
and U8314 (N_8314,N_6924,N_6096);
xor U8315 (N_8315,N_6226,N_7071);
or U8316 (N_8316,N_6970,N_7462);
and U8317 (N_8317,N_6557,N_7347);
nand U8318 (N_8318,N_6197,N_6312);
and U8319 (N_8319,N_6824,N_6837);
and U8320 (N_8320,N_6090,N_6979);
nor U8321 (N_8321,N_6549,N_6966);
xnor U8322 (N_8322,N_6671,N_6409);
xor U8323 (N_8323,N_6254,N_7364);
nor U8324 (N_8324,N_6287,N_6032);
or U8325 (N_8325,N_6279,N_7307);
nand U8326 (N_8326,N_7214,N_6311);
nand U8327 (N_8327,N_6937,N_6540);
xor U8328 (N_8328,N_6601,N_6886);
nor U8329 (N_8329,N_6064,N_6703);
nand U8330 (N_8330,N_7243,N_7197);
nand U8331 (N_8331,N_6294,N_6077);
nand U8332 (N_8332,N_6511,N_6468);
or U8333 (N_8333,N_7177,N_6905);
xor U8334 (N_8334,N_6486,N_6810);
nand U8335 (N_8335,N_7359,N_6184);
and U8336 (N_8336,N_6672,N_6791);
nand U8337 (N_8337,N_7436,N_6123);
or U8338 (N_8338,N_6602,N_6839);
or U8339 (N_8339,N_7434,N_7156);
xnor U8340 (N_8340,N_6139,N_6023);
and U8341 (N_8341,N_6891,N_6573);
nand U8342 (N_8342,N_7212,N_6286);
and U8343 (N_8343,N_7001,N_6846);
xor U8344 (N_8344,N_6927,N_7431);
and U8345 (N_8345,N_6348,N_6477);
and U8346 (N_8346,N_7026,N_6986);
xor U8347 (N_8347,N_6128,N_7102);
or U8348 (N_8348,N_7497,N_7166);
nand U8349 (N_8349,N_6988,N_7440);
xor U8350 (N_8350,N_6097,N_7022);
nand U8351 (N_8351,N_7006,N_6596);
xor U8352 (N_8352,N_6960,N_6847);
nor U8353 (N_8353,N_6418,N_6250);
nand U8354 (N_8354,N_6389,N_7470);
nor U8355 (N_8355,N_6472,N_6204);
nand U8356 (N_8356,N_6275,N_7407);
xor U8357 (N_8357,N_6814,N_7423);
nand U8358 (N_8358,N_7334,N_7256);
xnor U8359 (N_8359,N_7160,N_6653);
and U8360 (N_8360,N_6752,N_6086);
or U8361 (N_8361,N_6450,N_6877);
and U8362 (N_8362,N_6514,N_7493);
nand U8363 (N_8363,N_6247,N_6754);
xor U8364 (N_8364,N_6742,N_6343);
and U8365 (N_8365,N_6895,N_7070);
or U8366 (N_8366,N_6005,N_6206);
xnor U8367 (N_8367,N_6603,N_6498);
nor U8368 (N_8368,N_6424,N_6168);
xor U8369 (N_8369,N_7068,N_6971);
or U8370 (N_8370,N_6848,N_6182);
and U8371 (N_8371,N_7056,N_6998);
nor U8372 (N_8372,N_6876,N_6986);
xnor U8373 (N_8373,N_6370,N_6626);
nand U8374 (N_8374,N_6481,N_7265);
nand U8375 (N_8375,N_6584,N_7419);
xnor U8376 (N_8376,N_6807,N_6756);
and U8377 (N_8377,N_7239,N_6583);
or U8378 (N_8378,N_6892,N_7465);
and U8379 (N_8379,N_7293,N_6372);
or U8380 (N_8380,N_6450,N_6891);
and U8381 (N_8381,N_6489,N_7277);
xor U8382 (N_8382,N_6994,N_6866);
or U8383 (N_8383,N_6119,N_6720);
nor U8384 (N_8384,N_6597,N_7315);
or U8385 (N_8385,N_7323,N_6949);
or U8386 (N_8386,N_6954,N_6968);
xor U8387 (N_8387,N_6651,N_6399);
xnor U8388 (N_8388,N_6013,N_6090);
xnor U8389 (N_8389,N_7173,N_6706);
nand U8390 (N_8390,N_7347,N_6116);
or U8391 (N_8391,N_6739,N_6173);
or U8392 (N_8392,N_7266,N_7461);
nor U8393 (N_8393,N_6865,N_6015);
or U8394 (N_8394,N_6921,N_7276);
or U8395 (N_8395,N_6294,N_7319);
or U8396 (N_8396,N_6320,N_6143);
and U8397 (N_8397,N_7126,N_6080);
xnor U8398 (N_8398,N_6244,N_6557);
or U8399 (N_8399,N_6371,N_7348);
nor U8400 (N_8400,N_6367,N_6697);
xor U8401 (N_8401,N_7403,N_7185);
or U8402 (N_8402,N_7116,N_7067);
xnor U8403 (N_8403,N_6979,N_6458);
xnor U8404 (N_8404,N_7213,N_6110);
xor U8405 (N_8405,N_6045,N_6131);
xnor U8406 (N_8406,N_6310,N_6451);
nand U8407 (N_8407,N_6412,N_6127);
or U8408 (N_8408,N_7327,N_6850);
and U8409 (N_8409,N_6314,N_6068);
or U8410 (N_8410,N_7265,N_6009);
nand U8411 (N_8411,N_6275,N_6672);
or U8412 (N_8412,N_6543,N_7238);
and U8413 (N_8413,N_7259,N_7124);
nand U8414 (N_8414,N_6646,N_6545);
nor U8415 (N_8415,N_6390,N_7326);
xnor U8416 (N_8416,N_6035,N_6791);
and U8417 (N_8417,N_7077,N_6459);
and U8418 (N_8418,N_6914,N_6320);
nor U8419 (N_8419,N_6859,N_6359);
nand U8420 (N_8420,N_6269,N_6826);
or U8421 (N_8421,N_7485,N_7476);
and U8422 (N_8422,N_7146,N_6628);
nor U8423 (N_8423,N_6156,N_6578);
and U8424 (N_8424,N_6028,N_6286);
xnor U8425 (N_8425,N_6083,N_7022);
xnor U8426 (N_8426,N_7177,N_6991);
nand U8427 (N_8427,N_6391,N_7160);
or U8428 (N_8428,N_6780,N_7226);
and U8429 (N_8429,N_6802,N_6169);
nor U8430 (N_8430,N_6723,N_6968);
nor U8431 (N_8431,N_6355,N_6527);
nor U8432 (N_8432,N_6760,N_7364);
nor U8433 (N_8433,N_6860,N_7484);
or U8434 (N_8434,N_7114,N_6951);
and U8435 (N_8435,N_7473,N_6246);
nor U8436 (N_8436,N_6525,N_6499);
and U8437 (N_8437,N_6991,N_7203);
nor U8438 (N_8438,N_6844,N_7097);
and U8439 (N_8439,N_6754,N_7452);
and U8440 (N_8440,N_6510,N_6354);
nand U8441 (N_8441,N_7169,N_6980);
or U8442 (N_8442,N_7003,N_7301);
nand U8443 (N_8443,N_6192,N_6826);
nand U8444 (N_8444,N_6212,N_6933);
and U8445 (N_8445,N_7256,N_7337);
xnor U8446 (N_8446,N_6067,N_7379);
nor U8447 (N_8447,N_6719,N_7183);
or U8448 (N_8448,N_6676,N_6211);
and U8449 (N_8449,N_6858,N_7066);
nor U8450 (N_8450,N_6706,N_6687);
and U8451 (N_8451,N_7246,N_7362);
and U8452 (N_8452,N_7399,N_6878);
xor U8453 (N_8453,N_7095,N_6141);
xor U8454 (N_8454,N_6837,N_6334);
and U8455 (N_8455,N_7083,N_6791);
nor U8456 (N_8456,N_6465,N_6886);
nand U8457 (N_8457,N_6703,N_7328);
or U8458 (N_8458,N_6920,N_6528);
and U8459 (N_8459,N_6926,N_6956);
or U8460 (N_8460,N_6196,N_6222);
nor U8461 (N_8461,N_6017,N_6556);
nor U8462 (N_8462,N_7430,N_6084);
or U8463 (N_8463,N_7475,N_6956);
nand U8464 (N_8464,N_6652,N_7074);
nand U8465 (N_8465,N_6966,N_7041);
and U8466 (N_8466,N_7442,N_7413);
nand U8467 (N_8467,N_6313,N_6805);
or U8468 (N_8468,N_6127,N_7313);
xor U8469 (N_8469,N_6766,N_6107);
or U8470 (N_8470,N_6762,N_6587);
and U8471 (N_8471,N_6996,N_6573);
or U8472 (N_8472,N_6582,N_6744);
nor U8473 (N_8473,N_7212,N_6329);
and U8474 (N_8474,N_6621,N_7067);
xnor U8475 (N_8475,N_6687,N_6437);
nand U8476 (N_8476,N_6761,N_6413);
and U8477 (N_8477,N_6637,N_6558);
and U8478 (N_8478,N_6283,N_6562);
xnor U8479 (N_8479,N_7174,N_7380);
and U8480 (N_8480,N_6987,N_7076);
nor U8481 (N_8481,N_6939,N_7435);
or U8482 (N_8482,N_6809,N_6659);
or U8483 (N_8483,N_6026,N_6435);
or U8484 (N_8484,N_6119,N_7141);
and U8485 (N_8485,N_6210,N_6726);
nand U8486 (N_8486,N_6795,N_7332);
or U8487 (N_8487,N_7387,N_7294);
xnor U8488 (N_8488,N_7468,N_6727);
xor U8489 (N_8489,N_6211,N_6092);
and U8490 (N_8490,N_7021,N_6502);
or U8491 (N_8491,N_6289,N_6864);
and U8492 (N_8492,N_7204,N_6468);
nor U8493 (N_8493,N_6135,N_6317);
or U8494 (N_8494,N_6181,N_6705);
and U8495 (N_8495,N_7224,N_6628);
and U8496 (N_8496,N_7074,N_6584);
nor U8497 (N_8497,N_6813,N_7071);
xor U8498 (N_8498,N_6770,N_6796);
or U8499 (N_8499,N_6184,N_7376);
nand U8500 (N_8500,N_6656,N_6731);
nor U8501 (N_8501,N_6409,N_6307);
or U8502 (N_8502,N_6351,N_6282);
xor U8503 (N_8503,N_7329,N_7430);
and U8504 (N_8504,N_7086,N_7251);
nor U8505 (N_8505,N_7004,N_6925);
xnor U8506 (N_8506,N_7185,N_6638);
nor U8507 (N_8507,N_6741,N_7241);
or U8508 (N_8508,N_7022,N_6539);
nand U8509 (N_8509,N_6920,N_6618);
or U8510 (N_8510,N_6016,N_6063);
xnor U8511 (N_8511,N_6535,N_6056);
and U8512 (N_8512,N_6853,N_7313);
xnor U8513 (N_8513,N_6475,N_7380);
and U8514 (N_8514,N_6775,N_7412);
xor U8515 (N_8515,N_7474,N_6546);
and U8516 (N_8516,N_7270,N_7100);
nand U8517 (N_8517,N_6573,N_6747);
and U8518 (N_8518,N_7107,N_6776);
or U8519 (N_8519,N_6378,N_6091);
or U8520 (N_8520,N_6142,N_7102);
xnor U8521 (N_8521,N_7195,N_6842);
and U8522 (N_8522,N_6436,N_6006);
and U8523 (N_8523,N_7066,N_6381);
nand U8524 (N_8524,N_6560,N_6926);
and U8525 (N_8525,N_6444,N_7344);
nand U8526 (N_8526,N_6652,N_7027);
xnor U8527 (N_8527,N_6289,N_6228);
xor U8528 (N_8528,N_6938,N_6326);
nand U8529 (N_8529,N_7286,N_7351);
nand U8530 (N_8530,N_6576,N_6802);
or U8531 (N_8531,N_6829,N_7292);
xnor U8532 (N_8532,N_6976,N_6276);
nand U8533 (N_8533,N_6955,N_6787);
or U8534 (N_8534,N_6154,N_7358);
or U8535 (N_8535,N_6355,N_6554);
or U8536 (N_8536,N_7368,N_6803);
or U8537 (N_8537,N_6073,N_7340);
xor U8538 (N_8538,N_6781,N_6736);
nand U8539 (N_8539,N_7490,N_7021);
and U8540 (N_8540,N_6160,N_6520);
and U8541 (N_8541,N_6109,N_7008);
and U8542 (N_8542,N_6987,N_6460);
and U8543 (N_8543,N_6760,N_6637);
nand U8544 (N_8544,N_7011,N_7141);
nand U8545 (N_8545,N_6538,N_7459);
and U8546 (N_8546,N_7076,N_7167);
or U8547 (N_8547,N_6384,N_6978);
nand U8548 (N_8548,N_7234,N_6774);
xnor U8549 (N_8549,N_6677,N_6094);
or U8550 (N_8550,N_7385,N_6248);
nor U8551 (N_8551,N_6550,N_6808);
nand U8552 (N_8552,N_7264,N_7303);
nor U8553 (N_8553,N_7412,N_6268);
nor U8554 (N_8554,N_6998,N_6580);
nor U8555 (N_8555,N_6065,N_6077);
nor U8556 (N_8556,N_6627,N_6639);
or U8557 (N_8557,N_6227,N_6584);
nor U8558 (N_8558,N_6516,N_6102);
nor U8559 (N_8559,N_6179,N_7187);
nand U8560 (N_8560,N_6688,N_6800);
or U8561 (N_8561,N_7441,N_6611);
nand U8562 (N_8562,N_7383,N_6845);
nand U8563 (N_8563,N_6822,N_6295);
xnor U8564 (N_8564,N_6256,N_7023);
nor U8565 (N_8565,N_6477,N_6511);
nor U8566 (N_8566,N_7146,N_6765);
xnor U8567 (N_8567,N_7382,N_6260);
nand U8568 (N_8568,N_7451,N_6938);
or U8569 (N_8569,N_6968,N_6882);
xnor U8570 (N_8570,N_6692,N_6119);
or U8571 (N_8571,N_6937,N_6608);
and U8572 (N_8572,N_6006,N_6586);
and U8573 (N_8573,N_7287,N_6796);
and U8574 (N_8574,N_6163,N_7039);
or U8575 (N_8575,N_6675,N_6224);
xnor U8576 (N_8576,N_6389,N_6844);
or U8577 (N_8577,N_6293,N_6973);
nor U8578 (N_8578,N_7018,N_6817);
nand U8579 (N_8579,N_7164,N_6611);
or U8580 (N_8580,N_6003,N_6926);
nand U8581 (N_8581,N_6256,N_6140);
or U8582 (N_8582,N_6280,N_6301);
xor U8583 (N_8583,N_6055,N_6480);
nand U8584 (N_8584,N_6058,N_6997);
nor U8585 (N_8585,N_6560,N_7026);
and U8586 (N_8586,N_7295,N_7345);
nor U8587 (N_8587,N_6510,N_7350);
nor U8588 (N_8588,N_6653,N_6204);
and U8589 (N_8589,N_6531,N_7234);
nor U8590 (N_8590,N_6860,N_6988);
xnor U8591 (N_8591,N_6278,N_7162);
xor U8592 (N_8592,N_6540,N_6273);
and U8593 (N_8593,N_6456,N_7184);
or U8594 (N_8594,N_6500,N_6441);
xnor U8595 (N_8595,N_6544,N_6248);
and U8596 (N_8596,N_7090,N_7200);
nor U8597 (N_8597,N_6486,N_7023);
xor U8598 (N_8598,N_7117,N_6523);
or U8599 (N_8599,N_7389,N_7137);
xor U8600 (N_8600,N_6341,N_7145);
nand U8601 (N_8601,N_6322,N_6430);
xnor U8602 (N_8602,N_7393,N_6456);
nor U8603 (N_8603,N_6556,N_7438);
nor U8604 (N_8604,N_7225,N_6293);
nor U8605 (N_8605,N_6514,N_6402);
xor U8606 (N_8606,N_6157,N_6941);
and U8607 (N_8607,N_7213,N_6335);
and U8608 (N_8608,N_6359,N_6232);
nand U8609 (N_8609,N_7157,N_6061);
or U8610 (N_8610,N_7089,N_7239);
xor U8611 (N_8611,N_7372,N_6742);
nand U8612 (N_8612,N_6737,N_6118);
xnor U8613 (N_8613,N_6107,N_6922);
nor U8614 (N_8614,N_6283,N_7339);
or U8615 (N_8615,N_7360,N_6239);
xor U8616 (N_8616,N_7085,N_7064);
nor U8617 (N_8617,N_7089,N_7173);
nand U8618 (N_8618,N_6455,N_7355);
nor U8619 (N_8619,N_6502,N_7478);
xor U8620 (N_8620,N_7276,N_6239);
xor U8621 (N_8621,N_6933,N_7137);
nor U8622 (N_8622,N_6275,N_7421);
nor U8623 (N_8623,N_6936,N_6480);
nand U8624 (N_8624,N_6078,N_6616);
or U8625 (N_8625,N_7083,N_6510);
nor U8626 (N_8626,N_7189,N_6497);
nor U8627 (N_8627,N_6698,N_6528);
or U8628 (N_8628,N_6989,N_6467);
nor U8629 (N_8629,N_6636,N_6986);
nor U8630 (N_8630,N_6677,N_6336);
and U8631 (N_8631,N_7020,N_6949);
xor U8632 (N_8632,N_7466,N_6117);
or U8633 (N_8633,N_7253,N_7151);
nand U8634 (N_8634,N_7276,N_6188);
nand U8635 (N_8635,N_6341,N_6688);
or U8636 (N_8636,N_6011,N_7130);
xor U8637 (N_8637,N_6171,N_6203);
or U8638 (N_8638,N_7169,N_7078);
and U8639 (N_8639,N_6648,N_6335);
xor U8640 (N_8640,N_6093,N_6328);
or U8641 (N_8641,N_6889,N_6296);
xor U8642 (N_8642,N_6252,N_6085);
or U8643 (N_8643,N_7377,N_7165);
or U8644 (N_8644,N_7332,N_6877);
or U8645 (N_8645,N_6966,N_6630);
xor U8646 (N_8646,N_6843,N_6635);
and U8647 (N_8647,N_6978,N_6589);
nor U8648 (N_8648,N_7355,N_6592);
nand U8649 (N_8649,N_6310,N_6919);
and U8650 (N_8650,N_6574,N_6486);
and U8651 (N_8651,N_6053,N_7117);
or U8652 (N_8652,N_7187,N_6424);
or U8653 (N_8653,N_7262,N_6888);
and U8654 (N_8654,N_6052,N_7311);
xor U8655 (N_8655,N_7350,N_6575);
or U8656 (N_8656,N_7046,N_7116);
or U8657 (N_8657,N_6548,N_6210);
xor U8658 (N_8658,N_7447,N_6679);
and U8659 (N_8659,N_7145,N_7030);
and U8660 (N_8660,N_6494,N_7041);
xor U8661 (N_8661,N_6613,N_6148);
or U8662 (N_8662,N_7174,N_6755);
nor U8663 (N_8663,N_6394,N_6677);
xor U8664 (N_8664,N_6010,N_7139);
xor U8665 (N_8665,N_6468,N_7020);
nor U8666 (N_8666,N_6209,N_6093);
xnor U8667 (N_8667,N_7085,N_6928);
nor U8668 (N_8668,N_6854,N_6780);
nor U8669 (N_8669,N_6339,N_7351);
xnor U8670 (N_8670,N_6415,N_7018);
or U8671 (N_8671,N_7456,N_6857);
nor U8672 (N_8672,N_6733,N_6570);
xor U8673 (N_8673,N_6064,N_6469);
xor U8674 (N_8674,N_6804,N_7277);
and U8675 (N_8675,N_6107,N_6969);
and U8676 (N_8676,N_6698,N_6986);
or U8677 (N_8677,N_6551,N_6624);
nand U8678 (N_8678,N_6739,N_7104);
nor U8679 (N_8679,N_7332,N_6924);
nand U8680 (N_8680,N_6418,N_6210);
and U8681 (N_8681,N_6508,N_6310);
or U8682 (N_8682,N_6270,N_7241);
or U8683 (N_8683,N_6464,N_6179);
nor U8684 (N_8684,N_7380,N_7162);
or U8685 (N_8685,N_7043,N_6231);
xor U8686 (N_8686,N_6364,N_6984);
or U8687 (N_8687,N_7456,N_6240);
or U8688 (N_8688,N_6038,N_6181);
xor U8689 (N_8689,N_6629,N_6090);
or U8690 (N_8690,N_7024,N_6324);
nor U8691 (N_8691,N_6048,N_6616);
nor U8692 (N_8692,N_7491,N_6369);
or U8693 (N_8693,N_6622,N_6242);
nor U8694 (N_8694,N_6079,N_7468);
nand U8695 (N_8695,N_7351,N_6271);
and U8696 (N_8696,N_6061,N_7015);
and U8697 (N_8697,N_7336,N_6814);
nand U8698 (N_8698,N_7219,N_6153);
xnor U8699 (N_8699,N_6890,N_6279);
and U8700 (N_8700,N_6692,N_6971);
nor U8701 (N_8701,N_6597,N_6422);
xor U8702 (N_8702,N_6380,N_6385);
xnor U8703 (N_8703,N_7359,N_6145);
xor U8704 (N_8704,N_6331,N_7446);
and U8705 (N_8705,N_6670,N_6008);
and U8706 (N_8706,N_6521,N_7137);
nor U8707 (N_8707,N_7244,N_7485);
and U8708 (N_8708,N_6046,N_6370);
nor U8709 (N_8709,N_6959,N_6565);
xnor U8710 (N_8710,N_7478,N_6901);
xnor U8711 (N_8711,N_7104,N_6789);
xnor U8712 (N_8712,N_7280,N_6043);
nor U8713 (N_8713,N_7422,N_6900);
nor U8714 (N_8714,N_6937,N_7071);
or U8715 (N_8715,N_6095,N_6039);
nand U8716 (N_8716,N_6866,N_7259);
and U8717 (N_8717,N_6649,N_7051);
nor U8718 (N_8718,N_6683,N_6081);
nand U8719 (N_8719,N_7401,N_7246);
and U8720 (N_8720,N_6603,N_7473);
nand U8721 (N_8721,N_6563,N_6951);
xnor U8722 (N_8722,N_6272,N_6723);
or U8723 (N_8723,N_6029,N_6540);
or U8724 (N_8724,N_7061,N_6981);
xnor U8725 (N_8725,N_6392,N_7388);
nor U8726 (N_8726,N_7431,N_6969);
or U8727 (N_8727,N_6327,N_7052);
nand U8728 (N_8728,N_6059,N_6161);
nor U8729 (N_8729,N_7238,N_6534);
or U8730 (N_8730,N_6346,N_6469);
and U8731 (N_8731,N_7456,N_7459);
nand U8732 (N_8732,N_7086,N_6768);
nand U8733 (N_8733,N_6499,N_7296);
and U8734 (N_8734,N_6525,N_6102);
nand U8735 (N_8735,N_7341,N_6496);
or U8736 (N_8736,N_6372,N_6683);
nor U8737 (N_8737,N_7212,N_7310);
and U8738 (N_8738,N_7411,N_6194);
xnor U8739 (N_8739,N_6515,N_7479);
nor U8740 (N_8740,N_6874,N_7304);
xnor U8741 (N_8741,N_7114,N_6580);
and U8742 (N_8742,N_6543,N_7279);
or U8743 (N_8743,N_7259,N_6301);
and U8744 (N_8744,N_6618,N_7004);
xnor U8745 (N_8745,N_7394,N_7451);
and U8746 (N_8746,N_6751,N_6533);
nand U8747 (N_8747,N_6135,N_6310);
xor U8748 (N_8748,N_7317,N_6566);
xor U8749 (N_8749,N_6234,N_6547);
nand U8750 (N_8750,N_6713,N_6757);
or U8751 (N_8751,N_7006,N_6769);
nand U8752 (N_8752,N_6600,N_7060);
nor U8753 (N_8753,N_6342,N_6382);
nor U8754 (N_8754,N_6583,N_6261);
nand U8755 (N_8755,N_6720,N_7358);
or U8756 (N_8756,N_6571,N_6320);
nor U8757 (N_8757,N_6354,N_7484);
or U8758 (N_8758,N_7126,N_6609);
nor U8759 (N_8759,N_6230,N_6914);
nor U8760 (N_8760,N_7424,N_7412);
nor U8761 (N_8761,N_7016,N_6603);
nand U8762 (N_8762,N_6065,N_6351);
nor U8763 (N_8763,N_6846,N_7037);
nand U8764 (N_8764,N_7335,N_6027);
nor U8765 (N_8765,N_7296,N_6991);
xnor U8766 (N_8766,N_7039,N_6474);
and U8767 (N_8767,N_6609,N_7480);
and U8768 (N_8768,N_7316,N_7260);
xor U8769 (N_8769,N_7026,N_6532);
nor U8770 (N_8770,N_6265,N_6477);
or U8771 (N_8771,N_6412,N_7433);
nor U8772 (N_8772,N_6466,N_6879);
nand U8773 (N_8773,N_6590,N_6777);
nand U8774 (N_8774,N_7189,N_6370);
nand U8775 (N_8775,N_6162,N_6103);
nor U8776 (N_8776,N_7407,N_7392);
or U8777 (N_8777,N_6968,N_7310);
nand U8778 (N_8778,N_7233,N_6137);
nor U8779 (N_8779,N_6753,N_6493);
or U8780 (N_8780,N_6198,N_6544);
xnor U8781 (N_8781,N_6398,N_7049);
nand U8782 (N_8782,N_7173,N_7102);
and U8783 (N_8783,N_6774,N_6217);
nand U8784 (N_8784,N_6345,N_6605);
xnor U8785 (N_8785,N_6970,N_6554);
xnor U8786 (N_8786,N_7297,N_6918);
and U8787 (N_8787,N_6394,N_7444);
nand U8788 (N_8788,N_6302,N_7265);
or U8789 (N_8789,N_6920,N_7186);
nand U8790 (N_8790,N_6150,N_7415);
xnor U8791 (N_8791,N_7206,N_6060);
xor U8792 (N_8792,N_6796,N_7052);
nand U8793 (N_8793,N_6148,N_6466);
or U8794 (N_8794,N_7370,N_7433);
xnor U8795 (N_8795,N_7296,N_6391);
nand U8796 (N_8796,N_7370,N_6517);
nor U8797 (N_8797,N_6959,N_6858);
xnor U8798 (N_8798,N_6669,N_6586);
nor U8799 (N_8799,N_6787,N_6342);
and U8800 (N_8800,N_6636,N_7412);
xor U8801 (N_8801,N_7476,N_6498);
nand U8802 (N_8802,N_6047,N_6418);
and U8803 (N_8803,N_6388,N_7182);
nand U8804 (N_8804,N_7237,N_6910);
or U8805 (N_8805,N_6534,N_6723);
nor U8806 (N_8806,N_6714,N_7286);
xnor U8807 (N_8807,N_7497,N_7146);
and U8808 (N_8808,N_6222,N_6693);
xnor U8809 (N_8809,N_6471,N_7120);
nor U8810 (N_8810,N_6840,N_6456);
or U8811 (N_8811,N_7233,N_6302);
xnor U8812 (N_8812,N_7037,N_7059);
or U8813 (N_8813,N_7176,N_7250);
or U8814 (N_8814,N_7458,N_6147);
or U8815 (N_8815,N_6197,N_6779);
xor U8816 (N_8816,N_6973,N_7017);
nor U8817 (N_8817,N_6910,N_7085);
nor U8818 (N_8818,N_7084,N_6893);
nand U8819 (N_8819,N_6348,N_6746);
and U8820 (N_8820,N_7061,N_6177);
and U8821 (N_8821,N_6190,N_7271);
nand U8822 (N_8822,N_7335,N_6900);
xnor U8823 (N_8823,N_6390,N_7466);
nand U8824 (N_8824,N_6796,N_7479);
xnor U8825 (N_8825,N_6159,N_7395);
xnor U8826 (N_8826,N_7493,N_7283);
or U8827 (N_8827,N_6321,N_6349);
nor U8828 (N_8828,N_6421,N_6263);
and U8829 (N_8829,N_6772,N_7234);
or U8830 (N_8830,N_7135,N_6512);
or U8831 (N_8831,N_6876,N_6961);
xor U8832 (N_8832,N_6057,N_7284);
nor U8833 (N_8833,N_7227,N_6828);
nor U8834 (N_8834,N_7372,N_6320);
nor U8835 (N_8835,N_6915,N_6379);
or U8836 (N_8836,N_7123,N_7054);
and U8837 (N_8837,N_6000,N_6882);
or U8838 (N_8838,N_6827,N_6800);
or U8839 (N_8839,N_7106,N_7414);
nor U8840 (N_8840,N_7115,N_7485);
or U8841 (N_8841,N_7413,N_6641);
xor U8842 (N_8842,N_6414,N_6867);
nor U8843 (N_8843,N_6781,N_7249);
nor U8844 (N_8844,N_6532,N_6963);
or U8845 (N_8845,N_6530,N_6684);
xnor U8846 (N_8846,N_6549,N_6148);
xor U8847 (N_8847,N_7102,N_7026);
nand U8848 (N_8848,N_6949,N_6217);
or U8849 (N_8849,N_7009,N_6422);
and U8850 (N_8850,N_7203,N_7058);
and U8851 (N_8851,N_7069,N_7236);
or U8852 (N_8852,N_6228,N_6243);
nor U8853 (N_8853,N_6978,N_7469);
and U8854 (N_8854,N_6483,N_6343);
nor U8855 (N_8855,N_6836,N_6051);
or U8856 (N_8856,N_7311,N_6294);
and U8857 (N_8857,N_6865,N_6261);
or U8858 (N_8858,N_6623,N_7061);
or U8859 (N_8859,N_7476,N_6955);
or U8860 (N_8860,N_7494,N_6094);
xnor U8861 (N_8861,N_6866,N_6396);
and U8862 (N_8862,N_6492,N_6669);
and U8863 (N_8863,N_7473,N_7165);
nand U8864 (N_8864,N_6822,N_6556);
nand U8865 (N_8865,N_6800,N_6907);
or U8866 (N_8866,N_7200,N_6405);
nand U8867 (N_8867,N_6544,N_7385);
or U8868 (N_8868,N_7163,N_6346);
nor U8869 (N_8869,N_7162,N_6746);
xnor U8870 (N_8870,N_6111,N_7287);
and U8871 (N_8871,N_7412,N_7388);
xor U8872 (N_8872,N_6662,N_6460);
or U8873 (N_8873,N_6047,N_7076);
nor U8874 (N_8874,N_6817,N_6156);
nor U8875 (N_8875,N_6182,N_6485);
and U8876 (N_8876,N_6317,N_6851);
nor U8877 (N_8877,N_6199,N_7311);
xor U8878 (N_8878,N_7086,N_6875);
or U8879 (N_8879,N_6753,N_6601);
nand U8880 (N_8880,N_6532,N_7379);
or U8881 (N_8881,N_7371,N_6723);
and U8882 (N_8882,N_7285,N_6899);
nor U8883 (N_8883,N_7190,N_7315);
or U8884 (N_8884,N_7388,N_6867);
xnor U8885 (N_8885,N_6373,N_6983);
xor U8886 (N_8886,N_7206,N_7024);
or U8887 (N_8887,N_7415,N_6515);
and U8888 (N_8888,N_7329,N_6019);
and U8889 (N_8889,N_6481,N_7256);
nand U8890 (N_8890,N_7443,N_6970);
nor U8891 (N_8891,N_7200,N_6306);
nor U8892 (N_8892,N_6343,N_6708);
nand U8893 (N_8893,N_7027,N_6619);
xnor U8894 (N_8894,N_6750,N_6111);
nand U8895 (N_8895,N_7046,N_6613);
and U8896 (N_8896,N_6451,N_7062);
nand U8897 (N_8897,N_7209,N_6463);
nand U8898 (N_8898,N_6103,N_6606);
and U8899 (N_8899,N_6464,N_6973);
nand U8900 (N_8900,N_6990,N_6485);
and U8901 (N_8901,N_6462,N_7142);
nor U8902 (N_8902,N_6914,N_7474);
or U8903 (N_8903,N_6038,N_7315);
nor U8904 (N_8904,N_6864,N_6514);
nand U8905 (N_8905,N_7426,N_6251);
xor U8906 (N_8906,N_7097,N_6205);
nand U8907 (N_8907,N_6703,N_6955);
and U8908 (N_8908,N_7393,N_6443);
or U8909 (N_8909,N_7217,N_6803);
nand U8910 (N_8910,N_6469,N_6850);
and U8911 (N_8911,N_6076,N_7286);
nor U8912 (N_8912,N_6643,N_6411);
nand U8913 (N_8913,N_7491,N_6342);
xor U8914 (N_8914,N_7132,N_7440);
and U8915 (N_8915,N_7052,N_6495);
and U8916 (N_8916,N_6464,N_6498);
xor U8917 (N_8917,N_7238,N_6403);
xor U8918 (N_8918,N_6604,N_7137);
or U8919 (N_8919,N_6800,N_6307);
nor U8920 (N_8920,N_6641,N_6955);
and U8921 (N_8921,N_7080,N_6486);
or U8922 (N_8922,N_6233,N_6207);
or U8923 (N_8923,N_6190,N_7468);
or U8924 (N_8924,N_6165,N_7106);
or U8925 (N_8925,N_6563,N_6228);
and U8926 (N_8926,N_6464,N_6985);
and U8927 (N_8927,N_6497,N_6897);
xor U8928 (N_8928,N_6431,N_7220);
xor U8929 (N_8929,N_6527,N_6182);
and U8930 (N_8930,N_6047,N_6513);
nor U8931 (N_8931,N_7006,N_6459);
or U8932 (N_8932,N_6100,N_6369);
and U8933 (N_8933,N_6293,N_6688);
nor U8934 (N_8934,N_6049,N_6460);
and U8935 (N_8935,N_7289,N_6450);
and U8936 (N_8936,N_6101,N_6694);
nand U8937 (N_8937,N_7048,N_6826);
nor U8938 (N_8938,N_7050,N_7179);
nand U8939 (N_8939,N_6742,N_7200);
and U8940 (N_8940,N_6197,N_6904);
nor U8941 (N_8941,N_6422,N_7497);
nor U8942 (N_8942,N_6954,N_6812);
xnor U8943 (N_8943,N_6295,N_6071);
xor U8944 (N_8944,N_7223,N_6222);
nand U8945 (N_8945,N_7201,N_6241);
and U8946 (N_8946,N_6488,N_6028);
or U8947 (N_8947,N_7228,N_6873);
nand U8948 (N_8948,N_6748,N_6478);
xnor U8949 (N_8949,N_7361,N_6751);
nand U8950 (N_8950,N_6023,N_7141);
and U8951 (N_8951,N_7294,N_6371);
and U8952 (N_8952,N_6464,N_6538);
xor U8953 (N_8953,N_7069,N_6157);
or U8954 (N_8954,N_6647,N_7189);
and U8955 (N_8955,N_6979,N_7471);
nor U8956 (N_8956,N_6588,N_6512);
or U8957 (N_8957,N_6079,N_6052);
xor U8958 (N_8958,N_6489,N_7362);
and U8959 (N_8959,N_6229,N_6007);
xor U8960 (N_8960,N_6124,N_6095);
or U8961 (N_8961,N_6744,N_6999);
and U8962 (N_8962,N_6473,N_6953);
or U8963 (N_8963,N_6094,N_6396);
or U8964 (N_8964,N_6081,N_6162);
and U8965 (N_8965,N_6787,N_7327);
and U8966 (N_8966,N_6538,N_7488);
xor U8967 (N_8967,N_7288,N_7375);
and U8968 (N_8968,N_7397,N_6305);
nand U8969 (N_8969,N_6363,N_6622);
nand U8970 (N_8970,N_6417,N_6968);
xnor U8971 (N_8971,N_6397,N_6616);
nand U8972 (N_8972,N_7437,N_7495);
or U8973 (N_8973,N_7188,N_6317);
nand U8974 (N_8974,N_6162,N_6792);
and U8975 (N_8975,N_6082,N_7235);
or U8976 (N_8976,N_7119,N_7238);
nor U8977 (N_8977,N_7059,N_7277);
nor U8978 (N_8978,N_6645,N_7492);
xnor U8979 (N_8979,N_7340,N_6194);
xor U8980 (N_8980,N_6072,N_6496);
or U8981 (N_8981,N_7296,N_7288);
nand U8982 (N_8982,N_7205,N_7410);
nor U8983 (N_8983,N_7393,N_6021);
nand U8984 (N_8984,N_6426,N_7200);
nor U8985 (N_8985,N_7328,N_6257);
xnor U8986 (N_8986,N_6732,N_6149);
nand U8987 (N_8987,N_6575,N_6459);
nor U8988 (N_8988,N_6340,N_6317);
or U8989 (N_8989,N_6403,N_6686);
or U8990 (N_8990,N_6224,N_7346);
xnor U8991 (N_8991,N_7022,N_7399);
nand U8992 (N_8992,N_6252,N_7333);
xnor U8993 (N_8993,N_7388,N_7480);
nor U8994 (N_8994,N_6816,N_6513);
and U8995 (N_8995,N_7398,N_6793);
or U8996 (N_8996,N_6926,N_6211);
nand U8997 (N_8997,N_6666,N_7258);
nand U8998 (N_8998,N_7239,N_6124);
and U8999 (N_8999,N_6141,N_7464);
xor U9000 (N_9000,N_8206,N_7761);
nor U9001 (N_9001,N_8768,N_8657);
or U9002 (N_9002,N_8782,N_8746);
and U9003 (N_9003,N_8940,N_8813);
or U9004 (N_9004,N_8776,N_7810);
nand U9005 (N_9005,N_8750,N_8620);
nand U9006 (N_9006,N_7532,N_8505);
or U9007 (N_9007,N_8141,N_8994);
nor U9008 (N_9008,N_8823,N_8723);
nor U9009 (N_9009,N_8937,N_8644);
and U9010 (N_9010,N_8203,N_8373);
nand U9011 (N_9011,N_7704,N_8951);
or U9012 (N_9012,N_8862,N_7571);
or U9013 (N_9013,N_8988,N_8891);
nand U9014 (N_9014,N_8794,N_8114);
or U9015 (N_9015,N_8336,N_8310);
and U9016 (N_9016,N_8643,N_7832);
nor U9017 (N_9017,N_8322,N_8893);
nand U9018 (N_9018,N_8273,N_8137);
and U9019 (N_9019,N_7986,N_8866);
and U9020 (N_9020,N_8457,N_8412);
nor U9021 (N_9021,N_8555,N_7894);
nor U9022 (N_9022,N_8180,N_7950);
or U9023 (N_9023,N_7839,N_8035);
xor U9024 (N_9024,N_8223,N_8297);
or U9025 (N_9025,N_7682,N_8616);
nand U9026 (N_9026,N_7599,N_8199);
or U9027 (N_9027,N_8672,N_7664);
nor U9028 (N_9028,N_8158,N_7988);
or U9029 (N_9029,N_7779,N_7711);
nand U9030 (N_9030,N_8943,N_7521);
xnor U9031 (N_9031,N_7617,N_8701);
nand U9032 (N_9032,N_8634,N_7840);
or U9033 (N_9033,N_8175,N_8173);
xor U9034 (N_9034,N_8346,N_7981);
xor U9035 (N_9035,N_8513,N_8838);
nor U9036 (N_9036,N_7960,N_7838);
or U9037 (N_9037,N_8999,N_8392);
nor U9038 (N_9038,N_8081,N_7557);
xor U9039 (N_9039,N_8380,N_8969);
and U9040 (N_9040,N_8185,N_8564);
nor U9041 (N_9041,N_7511,N_7502);
and U9042 (N_9042,N_8984,N_7646);
xnor U9043 (N_9043,N_8692,N_7588);
or U9044 (N_9044,N_8883,N_7519);
or U9045 (N_9045,N_7522,N_8834);
and U9046 (N_9046,N_8339,N_8626);
or U9047 (N_9047,N_8451,N_8635);
nor U9048 (N_9048,N_8302,N_8758);
or U9049 (N_9049,N_7825,N_8464);
xor U9050 (N_9050,N_8831,N_8183);
or U9051 (N_9051,N_8415,N_8358);
nor U9052 (N_9052,N_8975,N_8507);
xnor U9053 (N_9053,N_8209,N_7737);
and U9054 (N_9054,N_7805,N_8836);
xor U9055 (N_9055,N_8193,N_8021);
nand U9056 (N_9056,N_8724,N_8720);
and U9057 (N_9057,N_7724,N_8145);
xnor U9058 (N_9058,N_7830,N_7590);
and U9059 (N_9059,N_8688,N_8664);
nand U9060 (N_9060,N_7964,N_8265);
nor U9061 (N_9061,N_8808,N_8015);
or U9062 (N_9062,N_8916,N_7924);
and U9063 (N_9063,N_8337,N_7996);
and U9064 (N_9064,N_8810,N_8868);
and U9065 (N_9065,N_8234,N_7655);
or U9066 (N_9066,N_7931,N_8286);
xor U9067 (N_9067,N_8689,N_7645);
or U9068 (N_9068,N_7944,N_8170);
nand U9069 (N_9069,N_8045,N_7970);
nand U9070 (N_9070,N_8540,N_8806);
or U9071 (N_9071,N_7824,N_7992);
or U9072 (N_9072,N_8097,N_8636);
xnor U9073 (N_9073,N_8867,N_8556);
nand U9074 (N_9074,N_7712,N_8453);
nor U9075 (N_9075,N_8211,N_7940);
or U9076 (N_9076,N_8587,N_8928);
nand U9077 (N_9077,N_8744,N_7624);
or U9078 (N_9078,N_7629,N_7754);
nand U9079 (N_9079,N_7886,N_8563);
nand U9080 (N_9080,N_7878,N_7551);
nand U9081 (N_9081,N_8870,N_7989);
xor U9082 (N_9082,N_8638,N_8532);
xnor U9083 (N_9083,N_7622,N_8172);
nor U9084 (N_9084,N_7549,N_8174);
xnor U9085 (N_9085,N_7735,N_8477);
xor U9086 (N_9086,N_8125,N_8245);
nor U9087 (N_9087,N_7969,N_7937);
and U9088 (N_9088,N_8352,N_8233);
xnor U9089 (N_9089,N_7841,N_8295);
and U9090 (N_9090,N_8013,N_7790);
nand U9091 (N_9091,N_8882,N_8987);
xnor U9092 (N_9092,N_8703,N_7560);
and U9093 (N_9093,N_8872,N_7956);
or U9094 (N_9094,N_8331,N_8287);
and U9095 (N_9095,N_7670,N_8506);
nor U9096 (N_9096,N_7884,N_8896);
nand U9097 (N_9097,N_8488,N_7581);
xor U9098 (N_9098,N_8349,N_8714);
or U9099 (N_9099,N_8379,N_7531);
nor U9100 (N_9100,N_7872,N_8027);
nand U9101 (N_9101,N_7852,N_8765);
nor U9102 (N_9102,N_8921,N_8117);
xnor U9103 (N_9103,N_7800,N_7829);
or U9104 (N_9104,N_8468,N_8847);
nand U9105 (N_9105,N_8875,N_7558);
or U9106 (N_9106,N_8908,N_8989);
or U9107 (N_9107,N_8001,N_8553);
nor U9108 (N_9108,N_7579,N_8702);
nor U9109 (N_9109,N_8600,N_8279);
xor U9110 (N_9110,N_7882,N_8930);
and U9111 (N_9111,N_8962,N_8923);
nand U9112 (N_9112,N_7782,N_8361);
nand U9113 (N_9113,N_7803,N_8374);
nor U9114 (N_9114,N_8881,N_7763);
and U9115 (N_9115,N_8727,N_7845);
and U9116 (N_9116,N_7576,N_8321);
and U9117 (N_9117,N_8046,N_7788);
and U9118 (N_9118,N_8026,N_8411);
or U9119 (N_9119,N_8278,N_8157);
or U9120 (N_9120,N_7921,N_7898);
xor U9121 (N_9121,N_7503,N_8742);
xor U9122 (N_9122,N_7536,N_8101);
nand U9123 (N_9123,N_8343,N_7636);
or U9124 (N_9124,N_8621,N_8116);
xnor U9125 (N_9125,N_8582,N_8828);
nor U9126 (N_9126,N_8285,N_8499);
xnor U9127 (N_9127,N_7934,N_7775);
and U9128 (N_9128,N_8455,N_8096);
and U9129 (N_9129,N_7923,N_7809);
and U9130 (N_9130,N_7768,N_8127);
xnor U9131 (N_9131,N_8409,N_7745);
and U9132 (N_9132,N_8382,N_7637);
nor U9133 (N_9133,N_8433,N_8238);
nand U9134 (N_9134,N_8603,N_8167);
xor U9135 (N_9135,N_8252,N_8601);
nor U9136 (N_9136,N_7807,N_7619);
and U9137 (N_9137,N_8003,N_8741);
nor U9138 (N_9138,N_8069,N_7595);
and U9139 (N_9139,N_7731,N_8375);
nand U9140 (N_9140,N_8461,N_7568);
nor U9141 (N_9141,N_8441,N_7669);
nand U9142 (N_9142,N_8973,N_8501);
nand U9143 (N_9143,N_7978,N_8598);
and U9144 (N_9144,N_7675,N_7747);
nor U9145 (N_9145,N_7570,N_7842);
nand U9146 (N_9146,N_8927,N_7866);
nand U9147 (N_9147,N_7974,N_8807);
or U9148 (N_9148,N_8777,N_8687);
nor U9149 (N_9149,N_7834,N_8931);
and U9150 (N_9150,N_8450,N_7612);
or U9151 (N_9151,N_8795,N_7527);
or U9152 (N_9152,N_8316,N_8067);
nand U9153 (N_9153,N_7723,N_7831);
xnor U9154 (N_9154,N_8200,N_8821);
nand U9155 (N_9155,N_8306,N_8985);
nand U9156 (N_9156,N_7792,N_8251);
and U9157 (N_9157,N_8159,N_8259);
or U9158 (N_9158,N_8722,N_8752);
nand U9159 (N_9159,N_8559,N_8960);
or U9160 (N_9160,N_8949,N_8475);
nor U9161 (N_9161,N_8978,N_8078);
xnor U9162 (N_9162,N_7601,N_8619);
xnor U9163 (N_9163,N_8088,N_8016);
and U9164 (N_9164,N_7739,N_8536);
xor U9165 (N_9165,N_7501,N_8524);
or U9166 (N_9166,N_7685,N_8425);
nor U9167 (N_9167,N_8263,N_8284);
or U9168 (N_9168,N_8844,N_7925);
nand U9169 (N_9169,N_8084,N_8493);
xnor U9170 (N_9170,N_8036,N_8121);
nor U9171 (N_9171,N_8188,N_8066);
nor U9172 (N_9172,N_8945,N_7856);
and U9173 (N_9173,N_8684,N_7574);
nor U9174 (N_9174,N_8229,N_8272);
and U9175 (N_9175,N_7600,N_8696);
nor U9176 (N_9176,N_8226,N_8602);
nand U9177 (N_9177,N_8571,N_8826);
nor U9178 (N_9178,N_8083,N_7941);
nor U9179 (N_9179,N_7722,N_8897);
or U9180 (N_9180,N_8000,N_7887);
or U9181 (N_9181,N_8064,N_7690);
nand U9182 (N_9182,N_8691,N_8557);
nand U9183 (N_9183,N_8712,N_7835);
nand U9184 (N_9184,N_8535,N_8715);
or U9185 (N_9185,N_7733,N_8543);
and U9186 (N_9186,N_8261,N_8394);
and U9187 (N_9187,N_7772,N_8965);
xor U9188 (N_9188,N_7597,N_7848);
or U9189 (N_9189,N_8890,N_7984);
or U9190 (N_9190,N_7708,N_8799);
and U9191 (N_9191,N_8319,N_8658);
and U9192 (N_9192,N_8198,N_7961);
xnor U9193 (N_9193,N_8822,N_8056);
nand U9194 (N_9194,N_8366,N_8055);
xor U9195 (N_9195,N_8248,N_8150);
or U9196 (N_9196,N_8661,N_8630);
xor U9197 (N_9197,N_8182,N_8397);
xnor U9198 (N_9198,N_8197,N_8177);
and U9199 (N_9199,N_8859,N_8797);
nor U9200 (N_9200,N_8617,N_8698);
or U9201 (N_9201,N_7959,N_7979);
xnor U9202 (N_9202,N_8075,N_8993);
nand U9203 (N_9203,N_8342,N_8113);
or U9204 (N_9204,N_8122,N_8291);
xnor U9205 (N_9205,N_8805,N_7710);
or U9206 (N_9206,N_8809,N_8649);
xnor U9207 (N_9207,N_8335,N_8710);
xnor U9208 (N_9208,N_8856,N_8749);
nor U9209 (N_9209,N_7677,N_7762);
or U9210 (N_9210,N_8640,N_8456);
nor U9211 (N_9211,N_8574,N_8376);
and U9212 (N_9212,N_8675,N_7982);
nand U9213 (N_9213,N_7876,N_7630);
xor U9214 (N_9214,N_8094,N_8262);
or U9215 (N_9215,N_8398,N_8944);
nand U9216 (N_9216,N_8019,N_8190);
and U9217 (N_9217,N_8326,N_7505);
nor U9218 (N_9218,N_8093,N_8857);
nand U9219 (N_9219,N_8186,N_8155);
xnor U9220 (N_9220,N_8663,N_8618);
xor U9221 (N_9221,N_8439,N_8538);
and U9222 (N_9222,N_8011,N_7973);
nand U9223 (N_9223,N_8947,N_8775);
nor U9224 (N_9224,N_7653,N_8932);
nor U9225 (N_9225,N_7820,N_8963);
nand U9226 (N_9226,N_7865,N_8469);
nand U9227 (N_9227,N_8476,N_7935);
or U9228 (N_9228,N_8133,N_8982);
nor U9229 (N_9229,N_7555,N_8588);
and U9230 (N_9230,N_8474,N_8929);
xor U9231 (N_9231,N_7948,N_8979);
nand U9232 (N_9232,N_8637,N_7525);
and U9233 (N_9233,N_8440,N_8381);
nor U9234 (N_9234,N_8490,N_8552);
nor U9235 (N_9235,N_8227,N_7823);
and U9236 (N_9236,N_8938,N_8508);
and U9237 (N_9237,N_8156,N_7847);
nand U9238 (N_9238,N_8424,N_8678);
and U9239 (N_9239,N_7691,N_7638);
or U9240 (N_9240,N_8918,N_7618);
nor U9241 (N_9241,N_8268,N_8589);
and U9242 (N_9242,N_7596,N_8176);
nor U9243 (N_9243,N_8841,N_8860);
nand U9244 (N_9244,N_7680,N_8232);
nor U9245 (N_9245,N_8357,N_8920);
and U9246 (N_9246,N_8560,N_7626);
xnor U9247 (N_9247,N_8915,N_7631);
xor U9248 (N_9248,N_7889,N_8120);
nor U9249 (N_9249,N_7849,N_8955);
and U9250 (N_9250,N_7694,N_8079);
nand U9251 (N_9251,N_7783,N_8010);
nand U9252 (N_9252,N_8403,N_8107);
xnor U9253 (N_9253,N_8344,N_7874);
and U9254 (N_9254,N_7954,N_7938);
and U9255 (N_9255,N_7652,N_8610);
nand U9256 (N_9256,N_8431,N_8144);
nor U9257 (N_9257,N_8416,N_8400);
and U9258 (N_9258,N_8801,N_8271);
nor U9259 (N_9259,N_8814,N_8816);
and U9260 (N_9260,N_7512,N_8449);
nand U9261 (N_9261,N_7905,N_8849);
or U9262 (N_9262,N_7804,N_7688);
or U9263 (N_9263,N_8966,N_7813);
or U9264 (N_9264,N_7707,N_8423);
xnor U9265 (N_9265,N_8737,N_8407);
and U9266 (N_9266,N_8130,N_8537);
nand U9267 (N_9267,N_7529,N_7523);
nor U9268 (N_9268,N_7985,N_7806);
nor U9269 (N_9269,N_8235,N_7795);
nand U9270 (N_9270,N_8851,N_8562);
or U9271 (N_9271,N_8654,N_8941);
xnor U9272 (N_9272,N_7860,N_8767);
or U9273 (N_9273,N_8260,N_8024);
nor U9274 (N_9274,N_8991,N_8502);
nor U9275 (N_9275,N_7915,N_8334);
and U9276 (N_9276,N_8074,N_8061);
nor U9277 (N_9277,N_8042,N_8443);
nand U9278 (N_9278,N_8249,N_8485);
nand U9279 (N_9279,N_7955,N_8787);
xor U9280 (N_9280,N_7586,N_8578);
nor U9281 (N_9281,N_8406,N_8512);
or U9282 (N_9282,N_8731,N_7506);
nor U9283 (N_9283,N_8914,N_8364);
nor U9284 (N_9284,N_8189,N_7963);
nand U9285 (N_9285,N_7720,N_8494);
and U9286 (N_9286,N_8585,N_8668);
xnor U9287 (N_9287,N_7896,N_8781);
and U9288 (N_9288,N_7651,N_8550);
xnor U9289 (N_9289,N_8832,N_8037);
xor U9290 (N_9290,N_8244,N_8030);
xnor U9291 (N_9291,N_8926,N_8526);
and U9292 (N_9292,N_7728,N_8653);
and U9293 (N_9293,N_8025,N_8481);
nor U9294 (N_9294,N_8429,N_8242);
nor U9295 (N_9295,N_8818,N_8002);
or U9296 (N_9296,N_7572,N_8467);
or U9297 (N_9297,N_7573,N_7995);
and U9298 (N_9298,N_7787,N_8936);
and U9299 (N_9299,N_8372,N_8216);
and U9300 (N_9300,N_8509,N_8325);
nor U9301 (N_9301,N_8996,N_8704);
and U9302 (N_9302,N_7513,N_8707);
and U9303 (N_9303,N_8759,N_7643);
and U9304 (N_9304,N_8539,N_7911);
xnor U9305 (N_9305,N_8837,N_8530);
nand U9306 (N_9306,N_8395,N_7952);
xor U9307 (N_9307,N_7533,N_8280);
nand U9308 (N_9308,N_7867,N_7880);
nand U9309 (N_9309,N_7908,N_8089);
xor U9310 (N_9310,N_7858,N_7583);
and U9311 (N_9311,N_8910,N_7546);
xor U9312 (N_9312,N_7801,N_7966);
nor U9313 (N_9313,N_7530,N_8545);
or U9314 (N_9314,N_7584,N_8317);
or U9315 (N_9315,N_8052,N_8566);
and U9316 (N_9316,N_7564,N_8895);
xor U9317 (N_9317,N_8480,N_8236);
or U9318 (N_9318,N_8038,N_8575);
nand U9319 (N_9319,N_8264,N_8134);
nand U9320 (N_9320,N_8212,N_8419);
nor U9321 (N_9321,N_8596,N_8631);
or U9322 (N_9322,N_7817,N_8080);
nor U9323 (N_9323,N_8031,N_8817);
xor U9324 (N_9324,N_8105,N_7854);
xor U9325 (N_9325,N_8700,N_8925);
nand U9326 (N_9326,N_7671,N_7883);
or U9327 (N_9327,N_8980,N_8783);
nand U9328 (N_9328,N_7500,N_7547);
or U9329 (N_9329,N_8528,N_8580);
nand U9330 (N_9330,N_8140,N_8472);
or U9331 (N_9331,N_8544,N_8732);
or U9332 (N_9332,N_8139,N_8320);
or U9333 (N_9333,N_8018,N_8681);
nor U9334 (N_9334,N_8676,N_7930);
nor U9335 (N_9335,N_8300,N_8593);
or U9336 (N_9336,N_7641,N_7649);
and U9337 (N_9337,N_7709,N_8099);
nor U9338 (N_9338,N_8459,N_8142);
and U9339 (N_9339,N_7700,N_8465);
nor U9340 (N_9340,N_7687,N_7696);
xor U9341 (N_9341,N_8231,N_8225);
nand U9342 (N_9342,N_8281,N_7580);
or U9343 (N_9343,N_8179,N_8674);
nand U9344 (N_9344,N_8774,N_8169);
nand U9345 (N_9345,N_8006,N_8109);
nor U9346 (N_9346,N_7912,N_8864);
nor U9347 (N_9347,N_7871,N_8132);
nand U9348 (N_9348,N_8491,N_8716);
or U9349 (N_9349,N_8110,N_8303);
or U9350 (N_9350,N_8377,N_7589);
nand U9351 (N_9351,N_7833,N_7881);
nor U9352 (N_9352,N_7818,N_8308);
and U9353 (N_9353,N_8420,N_7776);
and U9354 (N_9354,N_7877,N_7697);
xor U9355 (N_9355,N_7802,N_8143);
xor U9356 (N_9356,N_8386,N_8623);
nand U9357 (N_9357,N_8869,N_8168);
nand U9358 (N_9358,N_8187,N_7774);
xnor U9359 (N_9359,N_8679,N_8126);
nand U9360 (N_9360,N_7910,N_7765);
nand U9361 (N_9361,N_8964,N_8487);
or U9362 (N_9362,N_8426,N_8913);
or U9363 (N_9363,N_8523,N_8181);
or U9364 (N_9364,N_8733,N_8785);
nand U9365 (N_9365,N_8656,N_7543);
xor U9366 (N_9366,N_7900,N_7695);
or U9367 (N_9367,N_7642,N_8855);
and U9368 (N_9368,N_8390,N_8028);
and U9369 (N_9369,N_8436,N_8497);
and U9370 (N_9370,N_7702,N_8815);
xor U9371 (N_9371,N_8250,N_8332);
nor U9372 (N_9372,N_8854,N_7859);
nand U9373 (N_9373,N_7918,N_7821);
nor U9374 (N_9374,N_8218,N_8062);
and U9375 (N_9375,N_8473,N_8546);
and U9376 (N_9376,N_8511,N_7508);
xor U9377 (N_9377,N_8569,N_7784);
nor U9378 (N_9378,N_7851,N_7509);
or U9379 (N_9379,N_8370,N_8811);
xor U9380 (N_9380,N_8004,N_8292);
nand U9381 (N_9381,N_7693,N_8651);
or U9382 (N_9382,N_7759,N_8484);
and U9383 (N_9383,N_8830,N_8986);
nor U9384 (N_9384,N_8410,N_8492);
xor U9385 (N_9385,N_8106,N_7991);
xor U9386 (N_9386,N_8442,N_7604);
nor U9387 (N_9387,N_7556,N_7791);
or U9388 (N_9388,N_8953,N_7658);
xnor U9389 (N_9389,N_8434,N_7625);
nand U9390 (N_9390,N_8887,N_7518);
and U9391 (N_9391,N_8324,N_7798);
nor U9392 (N_9392,N_8213,N_8894);
nand U9393 (N_9393,N_8389,N_8751);
and U9394 (N_9394,N_8454,N_7901);
and U9395 (N_9395,N_8622,N_8470);
and U9396 (N_9396,N_8153,N_8665);
nor U9397 (N_9397,N_7785,N_8873);
nand U9398 (N_9398,N_8874,N_8763);
nand U9399 (N_9399,N_8572,N_8147);
xor U9400 (N_9400,N_7786,N_8118);
nand U9401 (N_9401,N_7706,N_8276);
nand U9402 (N_9402,N_8911,N_8008);
or U9403 (N_9403,N_8972,N_8648);
nand U9404 (N_9404,N_8353,N_8871);
and U9405 (N_9405,N_8422,N_7717);
or U9406 (N_9406,N_8779,N_8333);
or U9407 (N_9407,N_8705,N_8633);
nor U9408 (N_9408,N_8581,N_8592);
nor U9409 (N_9409,N_8729,N_8086);
nor U9410 (N_9410,N_8686,N_8812);
or U9411 (N_9411,N_8269,N_8309);
or U9412 (N_9412,N_7951,N_7705);
nand U9413 (N_9413,N_7741,N_7958);
xor U9414 (N_9414,N_8906,N_8059);
or U9415 (N_9415,N_8102,N_8076);
nor U9416 (N_9416,N_8047,N_7819);
and U9417 (N_9417,N_8071,N_7567);
and U9418 (N_9418,N_8256,N_7744);
and U9419 (N_9419,N_8104,N_7541);
or U9420 (N_9420,N_8728,N_8625);
or U9421 (N_9421,N_7827,N_8313);
nand U9422 (N_9422,N_7507,N_7668);
or U9423 (N_9423,N_7967,N_7539);
xnor U9424 (N_9424,N_8525,N_7528);
and U9425 (N_9425,N_7767,N_8583);
and U9426 (N_9426,N_7766,N_8356);
xnor U9427 (N_9427,N_8825,N_8095);
or U9428 (N_9428,N_8802,N_7701);
nor U9429 (N_9429,N_7561,N_8878);
and U9430 (N_9430,N_7692,N_8627);
nor U9431 (N_9431,N_7594,N_8057);
nand U9432 (N_9432,N_8541,N_8995);
xnor U9433 (N_9433,N_8877,N_8736);
nor U9434 (N_9434,N_7965,N_7535);
or U9435 (N_9435,N_7993,N_8243);
and U9436 (N_9436,N_7566,N_8747);
or U9437 (N_9437,N_8032,N_8208);
and U9438 (N_9438,N_8378,N_8152);
and U9439 (N_9439,N_8632,N_7603);
nor U9440 (N_9440,N_7748,N_8609);
xnor U9441 (N_9441,N_7730,N_7605);
nand U9442 (N_9442,N_8444,N_8458);
or U9443 (N_9443,N_7678,N_7907);
nand U9444 (N_9444,N_7927,N_8753);
and U9445 (N_9445,N_8605,N_8554);
nor U9446 (N_9446,N_8848,N_8967);
and U9447 (N_9447,N_8933,N_7746);
nor U9448 (N_9448,N_7773,N_8974);
nand U9449 (N_9449,N_7976,N_8519);
and U9450 (N_9450,N_7913,N_8773);
xnor U9451 (N_9451,N_8496,N_7822);
xor U9452 (N_9452,N_8624,N_8903);
nand U9453 (N_9453,N_8217,N_8757);
xnor U9454 (N_9454,N_8085,N_8956);
or U9455 (N_9455,N_8463,N_8642);
and U9456 (N_9456,N_8100,N_8072);
nand U9457 (N_9457,N_7752,N_8981);
and U9458 (N_9458,N_8160,N_8148);
or U9459 (N_9459,N_7777,N_8901);
nand U9460 (N_9460,N_8889,N_7957);
xor U9461 (N_9461,N_8149,N_8437);
xor U9462 (N_9462,N_7794,N_7756);
xnor U9463 (N_9463,N_8258,N_8820);
nor U9464 (N_9464,N_8123,N_8452);
or U9465 (N_9465,N_8693,N_8124);
nand U9466 (N_9466,N_7554,N_8629);
nor U9467 (N_9467,N_8840,N_7633);
nor U9468 (N_9468,N_8842,N_8796);
or U9469 (N_9469,N_8892,N_7844);
xnor U9470 (N_9470,N_7760,N_7514);
or U9471 (N_9471,N_8222,N_7749);
or U9472 (N_9472,N_8219,N_7758);
and U9473 (N_9473,N_8023,N_7743);
nand U9474 (N_9474,N_8853,N_7909);
or U9475 (N_9475,N_7879,N_8880);
or U9476 (N_9476,N_8171,N_8007);
and U9477 (N_9477,N_8743,N_8129);
or U9478 (N_9478,N_7623,N_8958);
xnor U9479 (N_9479,N_8510,N_8043);
or U9480 (N_9480,N_8561,N_7975);
nand U9481 (N_9481,N_7899,N_8946);
nor U9482 (N_9482,N_7738,N_8330);
or U9483 (N_9483,N_7537,N_8367);
nor U9484 (N_9484,N_7983,N_7681);
xnor U9485 (N_9485,N_8597,N_8611);
and U9486 (N_9486,N_7721,N_8748);
nand U9487 (N_9487,N_7644,N_8103);
and U9488 (N_9488,N_8858,N_8471);
nand U9489 (N_9489,N_8639,N_7917);
xor U9490 (N_9490,N_8246,N_8329);
and U9491 (N_9491,N_8876,N_8387);
nand U9492 (N_9492,N_8201,N_7666);
nor U9493 (N_9493,N_7593,N_7620);
nand U9494 (N_9494,N_8014,N_8971);
and U9495 (N_9495,N_8119,N_8338);
or U9496 (N_9496,N_7640,N_8961);
or U9497 (N_9497,N_8548,N_8270);
xnor U9498 (N_9498,N_7591,N_8899);
and U9499 (N_9499,N_8551,N_8290);
nor U9500 (N_9500,N_8756,N_8682);
nand U9501 (N_9501,N_8983,N_7812);
or U9502 (N_9502,N_7582,N_7769);
nand U9503 (N_9503,N_8486,N_7771);
nor U9504 (N_9504,N_8520,N_7936);
nand U9505 (N_9505,N_8586,N_8531);
nand U9506 (N_9506,N_7815,N_8900);
nor U9507 (N_9507,N_7949,N_8888);
nand U9508 (N_9508,N_8504,N_8073);
nand U9509 (N_9509,N_8401,N_7888);
nor U9510 (N_9510,N_7716,N_8518);
xnor U9511 (N_9511,N_8228,N_8054);
and U9512 (N_9512,N_7713,N_7578);
or U9513 (N_9513,N_7524,N_7628);
and U9514 (N_9514,N_7602,N_8296);
or U9515 (N_9515,N_8614,N_7718);
nand U9516 (N_9516,N_8068,N_7719);
or U9517 (N_9517,N_8063,N_7793);
nand U9518 (N_9518,N_8495,N_8591);
xor U9519 (N_9519,N_8954,N_7897);
nand U9520 (N_9520,N_8770,N_7727);
and U9521 (N_9521,N_7861,N_7587);
and U9522 (N_9522,N_7656,N_8907);
xor U9523 (N_9523,N_8202,N_8740);
and U9524 (N_9524,N_8070,N_8294);
nand U9525 (N_9525,N_7892,N_8791);
xor U9526 (N_9526,N_8761,N_8824);
nor U9527 (N_9527,N_8514,N_8041);
or U9528 (N_9528,N_8584,N_8350);
xor U9529 (N_9529,N_8789,N_8288);
and U9530 (N_9530,N_8413,N_8482);
nand U9531 (N_9531,N_7780,N_8922);
nand U9532 (N_9532,N_8863,N_8348);
xnor U9533 (N_9533,N_8612,N_7699);
nor U9534 (N_9534,N_7904,N_8718);
nor U9535 (N_9535,N_7621,N_8769);
nand U9536 (N_9536,N_8060,N_8959);
nor U9537 (N_9537,N_8039,N_8690);
nor U9538 (N_9538,N_8369,N_8466);
xnor U9539 (N_9539,N_8220,N_8709);
or U9540 (N_9540,N_8950,N_8050);
xnor U9541 (N_9541,N_8368,N_7608);
nor U9542 (N_9542,N_8590,N_7863);
and U9543 (N_9543,N_8579,N_8230);
xnor U9544 (N_9544,N_8576,N_7864);
or U9545 (N_9545,N_7665,N_7614);
nor U9546 (N_9546,N_8438,N_7676);
or U9547 (N_9547,N_8565,N_7736);
and U9548 (N_9548,N_8607,N_8968);
and U9549 (N_9549,N_7715,N_8305);
or U9550 (N_9550,N_8852,N_7526);
nor U9551 (N_9551,N_8210,N_8721);
nand U9552 (N_9552,N_7650,N_8719);
or U9553 (N_9553,N_7799,N_8051);
nand U9554 (N_9554,N_8257,N_8745);
and U9555 (N_9555,N_8293,N_8393);
or U9556 (N_9556,N_8628,N_7661);
nor U9557 (N_9557,N_8846,N_7939);
or U9558 (N_9558,N_8146,N_8058);
and U9559 (N_9559,N_8462,N_8670);
nor U9560 (N_9560,N_8594,N_8087);
and U9561 (N_9561,N_8646,N_8098);
and U9562 (N_9562,N_8939,N_8363);
nand U9563 (N_9563,N_7504,N_8677);
or U9564 (N_9564,N_8766,N_8726);
or U9565 (N_9565,N_7943,N_7932);
and U9566 (N_9566,N_7598,N_8267);
or U9567 (N_9567,N_8253,N_8012);
and U9568 (N_9568,N_7544,N_8447);
xor U9569 (N_9569,N_8274,N_8077);
xor U9570 (N_9570,N_8044,N_7928);
or U9571 (N_9571,N_8717,N_7903);
nand U9572 (N_9572,N_8207,N_8166);
and U9573 (N_9573,N_8659,N_8347);
or U9574 (N_9574,N_7945,N_8780);
nor U9575 (N_9575,N_7808,N_7635);
nor U9576 (N_9576,N_8240,N_7703);
nand U9577 (N_9577,N_8115,N_8827);
nand U9578 (N_9578,N_8029,N_8040);
and U9579 (N_9579,N_8912,N_7919);
and U9580 (N_9580,N_8697,N_8568);
or U9581 (N_9581,N_8604,N_8221);
nand U9582 (N_9582,N_7616,N_7994);
and U9583 (N_9583,N_8017,N_8384);
or U9584 (N_9584,N_7550,N_8355);
nor U9585 (N_9585,N_8215,N_8204);
or U9586 (N_9586,N_8399,N_8247);
or U9587 (N_9587,N_7757,N_8608);
or U9588 (N_9588,N_8503,N_7673);
or U9589 (N_9589,N_8112,N_7698);
nand U9590 (N_9590,N_8053,N_8652);
nand U9591 (N_9591,N_8529,N_8613);
and U9592 (N_9592,N_8266,N_7607);
xor U9593 (N_9593,N_7534,N_8885);
nand U9594 (N_9594,N_7683,N_8713);
nor U9595 (N_9595,N_7953,N_8318);
and U9596 (N_9596,N_7545,N_8755);
nor U9597 (N_9597,N_7853,N_8904);
nor U9598 (N_9598,N_8843,N_8314);
xnor U9599 (N_9599,N_7609,N_7634);
or U9600 (N_9600,N_8323,N_8304);
or U9601 (N_9601,N_8090,N_8391);
xnor U9602 (N_9602,N_8020,N_8500);
or U9603 (N_9603,N_8845,N_8163);
and U9604 (N_9604,N_8754,N_8517);
or U9605 (N_9605,N_8091,N_7855);
nor U9606 (N_9606,N_8427,N_8778);
nand U9607 (N_9607,N_8673,N_8136);
and U9608 (N_9608,N_7686,N_7968);
xnor U9609 (N_9609,N_8282,N_7732);
or U9610 (N_9610,N_8666,N_7778);
nand U9611 (N_9611,N_8298,N_8404);
nand U9612 (N_9612,N_8283,N_8408);
xor U9613 (N_9613,N_7540,N_7559);
or U9614 (N_9614,N_8178,N_8345);
or U9615 (N_9615,N_8680,N_7662);
or U9616 (N_9616,N_7647,N_7962);
nor U9617 (N_9617,N_8428,N_7972);
and U9618 (N_9618,N_8730,N_7592);
nor U9619 (N_9619,N_7843,N_7714);
or U9620 (N_9620,N_8886,N_8446);
nor U9621 (N_9621,N_7672,N_7734);
or U9622 (N_9622,N_7684,N_7742);
xor U9623 (N_9623,N_7797,N_8647);
or U9624 (N_9624,N_7875,N_7781);
xor U9625 (N_9625,N_7873,N_8935);
nand U9626 (N_9626,N_7796,N_8917);
nor U9627 (N_9627,N_8092,N_8685);
nor U9628 (N_9628,N_8521,N_8022);
nor U9629 (N_9629,N_8421,N_8924);
and U9630 (N_9630,N_8196,N_7565);
xnor U9631 (N_9631,N_7552,N_7575);
xnor U9632 (N_9632,N_7947,N_7577);
xor U9633 (N_9633,N_8255,N_7828);
xnor U9634 (N_9634,N_8432,N_8341);
and U9635 (N_9635,N_7902,N_8224);
nor U9636 (N_9636,N_8711,N_8599);
and U9637 (N_9637,N_8738,N_8489);
or U9638 (N_9638,N_7674,N_7895);
or U9639 (N_9639,N_7726,N_8819);
or U9640 (N_9640,N_8549,N_8301);
xor U9641 (N_9641,N_8977,N_7515);
and U9642 (N_9642,N_8577,N_8483);
nand U9643 (N_9643,N_8195,N_8662);
xnor U9644 (N_9644,N_7542,N_8135);
xor U9645 (N_9645,N_7517,N_8184);
and U9646 (N_9646,N_8957,N_8448);
nand U9647 (N_9647,N_8194,N_8645);
nor U9648 (N_9648,N_8522,N_7657);
or U9649 (N_9649,N_7627,N_7998);
nand U9650 (N_9650,N_7837,N_8793);
xor U9651 (N_9651,N_7548,N_7836);
xnor U9652 (N_9652,N_7516,N_8034);
and U9653 (N_9653,N_8762,N_8942);
xnor U9654 (N_9654,N_7679,N_8418);
or U9655 (N_9655,N_7891,N_8214);
or U9656 (N_9656,N_8049,N_7615);
nor U9657 (N_9657,N_7725,N_8371);
nor U9658 (N_9658,N_8997,N_8328);
or U9659 (N_9659,N_8311,N_7606);
xor U9660 (N_9660,N_8570,N_7826);
nor U9661 (N_9661,N_7569,N_7654);
nor U9662 (N_9662,N_7632,N_7751);
or U9663 (N_9663,N_8516,N_8547);
or U9664 (N_9664,N_8660,N_8340);
xnor U9665 (N_9665,N_8695,N_8992);
nand U9666 (N_9666,N_7689,N_8641);
nor U9667 (N_9667,N_8735,N_8478);
xor U9668 (N_9668,N_8567,N_7922);
or U9669 (N_9669,N_8205,N_8706);
nor U9670 (N_9670,N_7929,N_7869);
and U9671 (N_9671,N_8976,N_7862);
or U9672 (N_9672,N_8671,N_8998);
or U9673 (N_9673,N_8239,N_7868);
or U9674 (N_9674,N_8033,N_7764);
nor U9675 (N_9675,N_8734,N_8764);
or U9676 (N_9676,N_8615,N_8165);
or U9677 (N_9677,N_8162,N_8275);
and U9678 (N_9678,N_8879,N_8669);
nand U9679 (N_9679,N_8312,N_8254);
and U9680 (N_9680,N_8479,N_8414);
xnor U9681 (N_9681,N_8108,N_8667);
nand U9682 (N_9682,N_8138,N_8784);
xnor U9683 (N_9683,N_8786,N_7906);
nor U9684 (N_9684,N_8788,N_7990);
and U9685 (N_9685,N_8362,N_8558);
nand U9686 (N_9686,N_8315,N_8241);
xor U9687 (N_9687,N_8909,N_7971);
xnor U9688 (N_9688,N_8277,N_7667);
and U9689 (N_9689,N_8402,N_8515);
nor U9690 (N_9690,N_7942,N_8835);
nand U9691 (N_9691,N_7885,N_8359);
nand U9692 (N_9692,N_8498,N_7648);
nand U9693 (N_9693,N_7610,N_8354);
xnor U9694 (N_9694,N_7980,N_8804);
xor U9695 (N_9695,N_7893,N_8161);
nor U9696 (N_9696,N_8534,N_7770);
xnor U9697 (N_9697,N_8430,N_8445);
nand U9698 (N_9698,N_8884,N_8383);
and U9699 (N_9699,N_7729,N_8405);
and U9700 (N_9700,N_8385,N_8460);
nand U9701 (N_9701,N_7933,N_8798);
nand U9702 (N_9702,N_8351,N_8009);
xor U9703 (N_9703,N_8327,N_7914);
nor U9704 (N_9704,N_8850,N_8952);
xnor U9705 (N_9705,N_8699,N_8934);
xnor U9706 (N_9706,N_8595,N_8237);
or U9707 (N_9707,N_8289,N_8606);
xor U9708 (N_9708,N_8829,N_8990);
nor U9709 (N_9709,N_7740,N_7816);
nand U9710 (N_9710,N_7987,N_8154);
and U9711 (N_9711,N_8694,N_7553);
and U9712 (N_9712,N_7997,N_8082);
or U9713 (N_9713,N_8048,N_8111);
and U9714 (N_9714,N_7563,N_8191);
or U9715 (N_9715,N_7611,N_8573);
or U9716 (N_9716,N_8800,N_7753);
nand U9717 (N_9717,N_7663,N_8861);
and U9718 (N_9718,N_7520,N_8650);
or U9719 (N_9719,N_8865,N_8360);
xor U9720 (N_9720,N_8131,N_8533);
xnor U9721 (N_9721,N_8396,N_7999);
or U9722 (N_9722,N_7811,N_7538);
or U9723 (N_9723,N_8164,N_7585);
nor U9724 (N_9724,N_7926,N_7755);
and U9725 (N_9725,N_7659,N_8772);
nor U9726 (N_9726,N_8898,N_8435);
xnor U9727 (N_9727,N_8919,N_7789);
nor U9728 (N_9728,N_7850,N_8655);
nand U9729 (N_9729,N_7870,N_8527);
nor U9730 (N_9730,N_8683,N_8905);
nor U9731 (N_9731,N_7660,N_7562);
nand U9732 (N_9732,N_8388,N_7846);
and U9733 (N_9733,N_8790,N_8948);
and U9734 (N_9734,N_8970,N_8005);
xor U9735 (N_9735,N_7613,N_8739);
or U9736 (N_9736,N_7750,N_7977);
xor U9737 (N_9737,N_8771,N_8803);
nor U9738 (N_9738,N_8833,N_8417);
xor U9739 (N_9739,N_8365,N_8708);
nor U9740 (N_9740,N_8542,N_8192);
or U9741 (N_9741,N_8065,N_7916);
nand U9742 (N_9742,N_7920,N_8307);
or U9743 (N_9743,N_7857,N_8151);
or U9744 (N_9744,N_8839,N_8902);
or U9745 (N_9745,N_7510,N_8725);
nand U9746 (N_9746,N_8299,N_8760);
xnor U9747 (N_9747,N_7946,N_7814);
and U9748 (N_9748,N_7639,N_7890);
or U9749 (N_9749,N_8128,N_8792);
nor U9750 (N_9750,N_8824,N_8594);
and U9751 (N_9751,N_8806,N_8001);
nor U9752 (N_9752,N_8925,N_8285);
xor U9753 (N_9753,N_7554,N_8111);
or U9754 (N_9754,N_8485,N_8912);
nor U9755 (N_9755,N_7749,N_8216);
and U9756 (N_9756,N_7630,N_7862);
or U9757 (N_9757,N_7873,N_8012);
nand U9758 (N_9758,N_7680,N_8031);
nand U9759 (N_9759,N_8107,N_8888);
or U9760 (N_9760,N_8477,N_8175);
or U9761 (N_9761,N_8672,N_8574);
and U9762 (N_9762,N_8368,N_7522);
nor U9763 (N_9763,N_7983,N_7608);
xnor U9764 (N_9764,N_7873,N_7778);
and U9765 (N_9765,N_8554,N_8713);
nand U9766 (N_9766,N_8986,N_8487);
or U9767 (N_9767,N_8094,N_7904);
or U9768 (N_9768,N_8905,N_7977);
xor U9769 (N_9769,N_7938,N_7509);
nor U9770 (N_9770,N_8467,N_7975);
nand U9771 (N_9771,N_8302,N_8745);
or U9772 (N_9772,N_7528,N_8100);
nand U9773 (N_9773,N_8517,N_8360);
nand U9774 (N_9774,N_8711,N_8966);
nand U9775 (N_9775,N_7548,N_8000);
xor U9776 (N_9776,N_8704,N_8764);
and U9777 (N_9777,N_8124,N_7549);
and U9778 (N_9778,N_8439,N_7700);
and U9779 (N_9779,N_8798,N_7744);
and U9780 (N_9780,N_7994,N_7535);
xnor U9781 (N_9781,N_8806,N_8285);
or U9782 (N_9782,N_8786,N_7703);
or U9783 (N_9783,N_8118,N_7788);
and U9784 (N_9784,N_7728,N_8036);
xnor U9785 (N_9785,N_8970,N_8667);
nand U9786 (N_9786,N_8928,N_8615);
xnor U9787 (N_9787,N_8892,N_7851);
and U9788 (N_9788,N_8601,N_8063);
or U9789 (N_9789,N_7708,N_7771);
or U9790 (N_9790,N_8614,N_8625);
nor U9791 (N_9791,N_8636,N_8724);
nand U9792 (N_9792,N_7894,N_8427);
nand U9793 (N_9793,N_7649,N_7584);
or U9794 (N_9794,N_8549,N_7669);
xor U9795 (N_9795,N_8444,N_8024);
nor U9796 (N_9796,N_8382,N_8417);
xor U9797 (N_9797,N_8627,N_8485);
nor U9798 (N_9798,N_8004,N_7593);
xor U9799 (N_9799,N_8979,N_8144);
or U9800 (N_9800,N_7872,N_7899);
or U9801 (N_9801,N_7709,N_7886);
nor U9802 (N_9802,N_8067,N_8481);
nand U9803 (N_9803,N_7573,N_8591);
nor U9804 (N_9804,N_7618,N_7632);
nand U9805 (N_9805,N_7861,N_8250);
and U9806 (N_9806,N_8054,N_8598);
and U9807 (N_9807,N_7802,N_8818);
and U9808 (N_9808,N_8899,N_7667);
nor U9809 (N_9809,N_8139,N_7680);
nand U9810 (N_9810,N_8814,N_8178);
or U9811 (N_9811,N_8387,N_7612);
nor U9812 (N_9812,N_7667,N_7694);
nor U9813 (N_9813,N_7541,N_8332);
or U9814 (N_9814,N_7755,N_7973);
or U9815 (N_9815,N_8889,N_8393);
and U9816 (N_9816,N_8483,N_7766);
nor U9817 (N_9817,N_8736,N_7583);
nor U9818 (N_9818,N_8986,N_7768);
nor U9819 (N_9819,N_8155,N_8513);
xor U9820 (N_9820,N_8328,N_7593);
nor U9821 (N_9821,N_8999,N_7542);
and U9822 (N_9822,N_8982,N_8693);
and U9823 (N_9823,N_7878,N_8115);
or U9824 (N_9824,N_8389,N_8683);
xnor U9825 (N_9825,N_7572,N_7833);
xnor U9826 (N_9826,N_7504,N_7608);
and U9827 (N_9827,N_7508,N_7786);
nand U9828 (N_9828,N_7874,N_8063);
or U9829 (N_9829,N_8488,N_8400);
nand U9830 (N_9830,N_8007,N_8524);
nand U9831 (N_9831,N_8172,N_8969);
xor U9832 (N_9832,N_8784,N_8585);
xor U9833 (N_9833,N_8930,N_7563);
and U9834 (N_9834,N_7894,N_8627);
nand U9835 (N_9835,N_7649,N_7518);
and U9836 (N_9836,N_8704,N_7743);
nand U9837 (N_9837,N_8208,N_8054);
nand U9838 (N_9838,N_8437,N_8851);
or U9839 (N_9839,N_8593,N_7880);
xnor U9840 (N_9840,N_8188,N_8189);
xnor U9841 (N_9841,N_8508,N_7520);
xor U9842 (N_9842,N_8119,N_8751);
or U9843 (N_9843,N_8246,N_8853);
nand U9844 (N_9844,N_7676,N_8297);
and U9845 (N_9845,N_8504,N_7931);
or U9846 (N_9846,N_8843,N_8881);
and U9847 (N_9847,N_8110,N_8502);
xor U9848 (N_9848,N_7805,N_8150);
or U9849 (N_9849,N_7866,N_8396);
or U9850 (N_9850,N_8917,N_7749);
or U9851 (N_9851,N_8561,N_7956);
xnor U9852 (N_9852,N_8601,N_8104);
nand U9853 (N_9853,N_8057,N_7592);
nor U9854 (N_9854,N_8068,N_8511);
and U9855 (N_9855,N_8375,N_7938);
xnor U9856 (N_9856,N_8455,N_7577);
and U9857 (N_9857,N_7528,N_8863);
nor U9858 (N_9858,N_8402,N_8830);
nand U9859 (N_9859,N_8188,N_8395);
and U9860 (N_9860,N_7673,N_7602);
nand U9861 (N_9861,N_8327,N_7877);
or U9862 (N_9862,N_7509,N_8370);
xnor U9863 (N_9863,N_8798,N_7785);
nor U9864 (N_9864,N_7904,N_8449);
nor U9865 (N_9865,N_7765,N_8524);
nor U9866 (N_9866,N_7579,N_8707);
nand U9867 (N_9867,N_8030,N_8510);
nand U9868 (N_9868,N_8347,N_8066);
nand U9869 (N_9869,N_8937,N_8617);
nand U9870 (N_9870,N_8468,N_8861);
nor U9871 (N_9871,N_8999,N_8813);
xnor U9872 (N_9872,N_8961,N_8830);
xnor U9873 (N_9873,N_7515,N_7887);
nor U9874 (N_9874,N_7806,N_7547);
nor U9875 (N_9875,N_7814,N_8605);
and U9876 (N_9876,N_8214,N_8567);
and U9877 (N_9877,N_8008,N_8293);
xor U9878 (N_9878,N_7821,N_8952);
xnor U9879 (N_9879,N_7604,N_8712);
or U9880 (N_9880,N_7764,N_8579);
nand U9881 (N_9881,N_8927,N_8214);
or U9882 (N_9882,N_8444,N_7611);
nand U9883 (N_9883,N_7669,N_8326);
nand U9884 (N_9884,N_8007,N_8670);
and U9885 (N_9885,N_8082,N_8501);
nor U9886 (N_9886,N_8185,N_7556);
and U9887 (N_9887,N_7682,N_8743);
or U9888 (N_9888,N_8014,N_8769);
xor U9889 (N_9889,N_8860,N_8944);
nand U9890 (N_9890,N_8536,N_8495);
or U9891 (N_9891,N_8152,N_7793);
nor U9892 (N_9892,N_7670,N_8835);
xor U9893 (N_9893,N_8545,N_7977);
nor U9894 (N_9894,N_8185,N_8369);
and U9895 (N_9895,N_7774,N_8801);
or U9896 (N_9896,N_8920,N_8696);
xnor U9897 (N_9897,N_8684,N_7501);
and U9898 (N_9898,N_8523,N_8600);
xnor U9899 (N_9899,N_7850,N_8200);
and U9900 (N_9900,N_8491,N_7919);
and U9901 (N_9901,N_7702,N_7976);
nor U9902 (N_9902,N_8331,N_7641);
or U9903 (N_9903,N_8139,N_8959);
nor U9904 (N_9904,N_7675,N_8714);
and U9905 (N_9905,N_8474,N_8006);
xnor U9906 (N_9906,N_8404,N_8008);
xor U9907 (N_9907,N_7512,N_8259);
nand U9908 (N_9908,N_8814,N_8370);
and U9909 (N_9909,N_7846,N_7500);
or U9910 (N_9910,N_8838,N_8921);
or U9911 (N_9911,N_8106,N_8000);
or U9912 (N_9912,N_7536,N_8171);
nor U9913 (N_9913,N_8204,N_7599);
or U9914 (N_9914,N_8736,N_7822);
nand U9915 (N_9915,N_7586,N_8396);
and U9916 (N_9916,N_8903,N_8206);
nand U9917 (N_9917,N_7588,N_7818);
nor U9918 (N_9918,N_8987,N_7829);
xnor U9919 (N_9919,N_8429,N_7944);
nand U9920 (N_9920,N_7924,N_8821);
and U9921 (N_9921,N_7767,N_8480);
xnor U9922 (N_9922,N_8897,N_8933);
nor U9923 (N_9923,N_8992,N_8198);
and U9924 (N_9924,N_7744,N_8115);
nor U9925 (N_9925,N_8237,N_8594);
or U9926 (N_9926,N_8421,N_7644);
xnor U9927 (N_9927,N_8702,N_8704);
or U9928 (N_9928,N_8247,N_8718);
xor U9929 (N_9929,N_7700,N_8143);
and U9930 (N_9930,N_8344,N_8789);
or U9931 (N_9931,N_8504,N_8305);
xor U9932 (N_9932,N_8614,N_8455);
and U9933 (N_9933,N_8703,N_8543);
and U9934 (N_9934,N_8318,N_8795);
xor U9935 (N_9935,N_8858,N_8097);
nor U9936 (N_9936,N_8074,N_8444);
nor U9937 (N_9937,N_8677,N_8616);
xor U9938 (N_9938,N_7650,N_8983);
or U9939 (N_9939,N_7505,N_8769);
or U9940 (N_9940,N_8451,N_8230);
nand U9941 (N_9941,N_8364,N_7584);
and U9942 (N_9942,N_8241,N_8565);
nor U9943 (N_9943,N_7845,N_8853);
or U9944 (N_9944,N_7846,N_8644);
nor U9945 (N_9945,N_8348,N_8360);
xor U9946 (N_9946,N_8363,N_8124);
xor U9947 (N_9947,N_8719,N_8756);
and U9948 (N_9948,N_8541,N_8751);
nand U9949 (N_9949,N_8308,N_8675);
and U9950 (N_9950,N_7500,N_7570);
nor U9951 (N_9951,N_8339,N_7925);
nor U9952 (N_9952,N_8582,N_8111);
nor U9953 (N_9953,N_7806,N_7559);
or U9954 (N_9954,N_7504,N_8991);
nand U9955 (N_9955,N_8520,N_8977);
nor U9956 (N_9956,N_8681,N_8452);
xnor U9957 (N_9957,N_8225,N_8174);
and U9958 (N_9958,N_8802,N_8567);
xor U9959 (N_9959,N_8432,N_7646);
nor U9960 (N_9960,N_8248,N_7576);
xor U9961 (N_9961,N_8506,N_8020);
xor U9962 (N_9962,N_8233,N_8804);
or U9963 (N_9963,N_8049,N_8067);
and U9964 (N_9964,N_8731,N_8646);
nand U9965 (N_9965,N_7726,N_7879);
nand U9966 (N_9966,N_7568,N_8559);
and U9967 (N_9967,N_8979,N_7742);
or U9968 (N_9968,N_7772,N_8953);
xor U9969 (N_9969,N_7534,N_7643);
or U9970 (N_9970,N_8853,N_8889);
or U9971 (N_9971,N_7828,N_8748);
or U9972 (N_9972,N_8136,N_8430);
xnor U9973 (N_9973,N_8148,N_8143);
nand U9974 (N_9974,N_7902,N_8261);
or U9975 (N_9975,N_7577,N_7641);
nor U9976 (N_9976,N_7657,N_8558);
and U9977 (N_9977,N_8787,N_8921);
and U9978 (N_9978,N_8626,N_8703);
xor U9979 (N_9979,N_7848,N_8056);
and U9980 (N_9980,N_8028,N_8255);
nor U9981 (N_9981,N_8991,N_8041);
nor U9982 (N_9982,N_8195,N_7523);
or U9983 (N_9983,N_8592,N_8140);
xor U9984 (N_9984,N_8625,N_8955);
and U9985 (N_9985,N_8283,N_8371);
and U9986 (N_9986,N_8528,N_7686);
or U9987 (N_9987,N_7727,N_7620);
xnor U9988 (N_9988,N_8522,N_8878);
and U9989 (N_9989,N_7688,N_8921);
xnor U9990 (N_9990,N_8139,N_8332);
nor U9991 (N_9991,N_8046,N_7886);
nor U9992 (N_9992,N_8157,N_8203);
and U9993 (N_9993,N_7570,N_8375);
xor U9994 (N_9994,N_7597,N_8856);
nor U9995 (N_9995,N_7727,N_8407);
and U9996 (N_9996,N_8552,N_7914);
or U9997 (N_9997,N_8745,N_7962);
or U9998 (N_9998,N_7863,N_8783);
nor U9999 (N_9999,N_8365,N_8149);
nand U10000 (N_10000,N_8944,N_7502);
xnor U10001 (N_10001,N_8030,N_7974);
xnor U10002 (N_10002,N_8979,N_8978);
and U10003 (N_10003,N_8864,N_8551);
or U10004 (N_10004,N_8335,N_7778);
nor U10005 (N_10005,N_7534,N_7758);
and U10006 (N_10006,N_7530,N_8980);
or U10007 (N_10007,N_8169,N_8948);
and U10008 (N_10008,N_7977,N_8254);
and U10009 (N_10009,N_7571,N_8513);
and U10010 (N_10010,N_8685,N_8293);
nor U10011 (N_10011,N_7639,N_8879);
nand U10012 (N_10012,N_8922,N_8721);
and U10013 (N_10013,N_8358,N_8246);
nand U10014 (N_10014,N_8276,N_8360);
xor U10015 (N_10015,N_8720,N_8604);
and U10016 (N_10016,N_8959,N_7506);
nor U10017 (N_10017,N_7859,N_7887);
and U10018 (N_10018,N_7623,N_7726);
or U10019 (N_10019,N_8493,N_8269);
nand U10020 (N_10020,N_7522,N_8754);
or U10021 (N_10021,N_8131,N_7669);
xnor U10022 (N_10022,N_7825,N_8727);
or U10023 (N_10023,N_8277,N_7677);
or U10024 (N_10024,N_8754,N_8021);
and U10025 (N_10025,N_8776,N_8956);
xnor U10026 (N_10026,N_8619,N_7597);
nand U10027 (N_10027,N_8974,N_7588);
xnor U10028 (N_10028,N_8491,N_7944);
nor U10029 (N_10029,N_7912,N_8313);
and U10030 (N_10030,N_7571,N_7946);
xnor U10031 (N_10031,N_8600,N_8596);
and U10032 (N_10032,N_8114,N_7650);
and U10033 (N_10033,N_8729,N_8245);
nor U10034 (N_10034,N_8506,N_8012);
nor U10035 (N_10035,N_7773,N_8645);
and U10036 (N_10036,N_8322,N_7763);
and U10037 (N_10037,N_8420,N_7543);
nand U10038 (N_10038,N_8877,N_7692);
and U10039 (N_10039,N_8887,N_7672);
xnor U10040 (N_10040,N_8006,N_8042);
nor U10041 (N_10041,N_8863,N_8428);
nand U10042 (N_10042,N_7740,N_8855);
nand U10043 (N_10043,N_8232,N_8116);
xnor U10044 (N_10044,N_8789,N_8384);
xor U10045 (N_10045,N_7623,N_7860);
or U10046 (N_10046,N_8775,N_7681);
and U10047 (N_10047,N_7880,N_7956);
nor U10048 (N_10048,N_8348,N_7703);
nor U10049 (N_10049,N_8082,N_8188);
or U10050 (N_10050,N_7796,N_8852);
nor U10051 (N_10051,N_8740,N_8661);
nand U10052 (N_10052,N_8629,N_8751);
or U10053 (N_10053,N_8184,N_7671);
nand U10054 (N_10054,N_8686,N_8075);
or U10055 (N_10055,N_8953,N_7882);
and U10056 (N_10056,N_7944,N_8127);
or U10057 (N_10057,N_7992,N_7615);
xor U10058 (N_10058,N_8589,N_8272);
and U10059 (N_10059,N_7557,N_7524);
and U10060 (N_10060,N_7734,N_7504);
nand U10061 (N_10061,N_8646,N_8537);
and U10062 (N_10062,N_7755,N_7786);
nand U10063 (N_10063,N_7602,N_8906);
nor U10064 (N_10064,N_8177,N_7526);
and U10065 (N_10065,N_7715,N_8523);
nand U10066 (N_10066,N_8109,N_8042);
nor U10067 (N_10067,N_8665,N_8609);
or U10068 (N_10068,N_8184,N_8122);
or U10069 (N_10069,N_7833,N_8236);
xor U10070 (N_10070,N_8695,N_8180);
xor U10071 (N_10071,N_8437,N_7764);
and U10072 (N_10072,N_8164,N_8622);
nand U10073 (N_10073,N_8887,N_8102);
xor U10074 (N_10074,N_8623,N_8566);
xor U10075 (N_10075,N_8191,N_7577);
xor U10076 (N_10076,N_8976,N_7834);
nand U10077 (N_10077,N_7862,N_7639);
or U10078 (N_10078,N_8396,N_8734);
xor U10079 (N_10079,N_7828,N_8471);
nand U10080 (N_10080,N_8372,N_8743);
nor U10081 (N_10081,N_8575,N_8028);
and U10082 (N_10082,N_8850,N_7626);
nand U10083 (N_10083,N_8188,N_8884);
or U10084 (N_10084,N_8753,N_7730);
or U10085 (N_10085,N_8810,N_8255);
and U10086 (N_10086,N_8939,N_7843);
or U10087 (N_10087,N_8215,N_7882);
and U10088 (N_10088,N_8694,N_7504);
nor U10089 (N_10089,N_7562,N_7841);
and U10090 (N_10090,N_8434,N_8568);
or U10091 (N_10091,N_8621,N_7991);
nand U10092 (N_10092,N_8076,N_8395);
nand U10093 (N_10093,N_8301,N_8290);
and U10094 (N_10094,N_8586,N_7864);
nand U10095 (N_10095,N_8776,N_7772);
nor U10096 (N_10096,N_7661,N_7691);
or U10097 (N_10097,N_8236,N_8462);
xnor U10098 (N_10098,N_8209,N_8598);
nor U10099 (N_10099,N_7662,N_7939);
nand U10100 (N_10100,N_7982,N_8011);
xor U10101 (N_10101,N_7750,N_8647);
and U10102 (N_10102,N_7889,N_8516);
xnor U10103 (N_10103,N_7719,N_7909);
and U10104 (N_10104,N_7765,N_8436);
or U10105 (N_10105,N_7994,N_8702);
or U10106 (N_10106,N_8887,N_7510);
xnor U10107 (N_10107,N_7554,N_8624);
nand U10108 (N_10108,N_7992,N_8919);
xnor U10109 (N_10109,N_8229,N_8120);
and U10110 (N_10110,N_8827,N_8934);
and U10111 (N_10111,N_8122,N_8311);
nor U10112 (N_10112,N_8746,N_8849);
or U10113 (N_10113,N_7754,N_8214);
nand U10114 (N_10114,N_7821,N_8372);
nor U10115 (N_10115,N_8939,N_7689);
and U10116 (N_10116,N_7671,N_8776);
and U10117 (N_10117,N_8724,N_8046);
and U10118 (N_10118,N_8465,N_8976);
xor U10119 (N_10119,N_7895,N_8507);
or U10120 (N_10120,N_8063,N_8772);
nand U10121 (N_10121,N_8649,N_8991);
xnor U10122 (N_10122,N_7576,N_7777);
nand U10123 (N_10123,N_8533,N_8331);
xnor U10124 (N_10124,N_8823,N_7847);
and U10125 (N_10125,N_8770,N_7823);
and U10126 (N_10126,N_7870,N_8752);
and U10127 (N_10127,N_8329,N_8706);
nand U10128 (N_10128,N_8627,N_7640);
nor U10129 (N_10129,N_8976,N_7641);
nor U10130 (N_10130,N_8528,N_7898);
nand U10131 (N_10131,N_8012,N_7560);
and U10132 (N_10132,N_8134,N_7743);
xor U10133 (N_10133,N_7889,N_7902);
or U10134 (N_10134,N_8332,N_8541);
or U10135 (N_10135,N_8031,N_7687);
and U10136 (N_10136,N_8469,N_8723);
nand U10137 (N_10137,N_8531,N_8259);
nand U10138 (N_10138,N_8823,N_8925);
and U10139 (N_10139,N_7882,N_8231);
nor U10140 (N_10140,N_7991,N_8636);
nand U10141 (N_10141,N_7639,N_8662);
xnor U10142 (N_10142,N_8799,N_8230);
and U10143 (N_10143,N_8577,N_8922);
nor U10144 (N_10144,N_8542,N_8880);
xnor U10145 (N_10145,N_8996,N_8213);
nor U10146 (N_10146,N_7673,N_7999);
and U10147 (N_10147,N_7846,N_7575);
and U10148 (N_10148,N_8790,N_7929);
and U10149 (N_10149,N_7970,N_8302);
and U10150 (N_10150,N_8698,N_7776);
xnor U10151 (N_10151,N_8355,N_8784);
nor U10152 (N_10152,N_8386,N_8489);
and U10153 (N_10153,N_7732,N_8781);
nand U10154 (N_10154,N_7613,N_8701);
or U10155 (N_10155,N_8312,N_8049);
nor U10156 (N_10156,N_8854,N_8568);
nand U10157 (N_10157,N_8639,N_8088);
xor U10158 (N_10158,N_8285,N_8431);
or U10159 (N_10159,N_7864,N_7592);
xnor U10160 (N_10160,N_8438,N_7811);
or U10161 (N_10161,N_7795,N_8849);
and U10162 (N_10162,N_7510,N_7909);
nor U10163 (N_10163,N_8335,N_8870);
xor U10164 (N_10164,N_7908,N_8986);
or U10165 (N_10165,N_7507,N_8054);
xor U10166 (N_10166,N_8403,N_8513);
and U10167 (N_10167,N_8050,N_8900);
nor U10168 (N_10168,N_8973,N_8913);
nor U10169 (N_10169,N_7699,N_8762);
nor U10170 (N_10170,N_8846,N_7608);
xnor U10171 (N_10171,N_8568,N_7940);
xnor U10172 (N_10172,N_8157,N_8844);
nor U10173 (N_10173,N_8886,N_8490);
nor U10174 (N_10174,N_7545,N_8605);
or U10175 (N_10175,N_8243,N_8740);
xor U10176 (N_10176,N_7715,N_8013);
nor U10177 (N_10177,N_7841,N_8231);
or U10178 (N_10178,N_8379,N_7950);
or U10179 (N_10179,N_8120,N_8007);
nand U10180 (N_10180,N_8044,N_8714);
nand U10181 (N_10181,N_8881,N_8324);
nand U10182 (N_10182,N_8158,N_8161);
nand U10183 (N_10183,N_7751,N_8891);
nand U10184 (N_10184,N_8840,N_8253);
nand U10185 (N_10185,N_8391,N_8624);
nand U10186 (N_10186,N_8457,N_7944);
or U10187 (N_10187,N_8490,N_7540);
xnor U10188 (N_10188,N_8853,N_8812);
or U10189 (N_10189,N_7810,N_8213);
nor U10190 (N_10190,N_7975,N_7758);
nor U10191 (N_10191,N_7859,N_8538);
or U10192 (N_10192,N_8372,N_8339);
xnor U10193 (N_10193,N_8747,N_8733);
and U10194 (N_10194,N_8254,N_7783);
or U10195 (N_10195,N_8796,N_7975);
or U10196 (N_10196,N_8958,N_8348);
and U10197 (N_10197,N_8481,N_7747);
nor U10198 (N_10198,N_8639,N_8849);
xor U10199 (N_10199,N_8539,N_8822);
nand U10200 (N_10200,N_8259,N_8641);
nor U10201 (N_10201,N_7965,N_8170);
xnor U10202 (N_10202,N_7913,N_7871);
nand U10203 (N_10203,N_8177,N_8267);
nand U10204 (N_10204,N_7852,N_8361);
and U10205 (N_10205,N_7559,N_7720);
and U10206 (N_10206,N_8513,N_8083);
xor U10207 (N_10207,N_8852,N_8033);
nand U10208 (N_10208,N_7825,N_8580);
or U10209 (N_10209,N_8105,N_8903);
nor U10210 (N_10210,N_8658,N_8871);
nand U10211 (N_10211,N_8247,N_7569);
or U10212 (N_10212,N_7966,N_8958);
or U10213 (N_10213,N_7886,N_8567);
or U10214 (N_10214,N_7854,N_8397);
or U10215 (N_10215,N_8948,N_8040);
xnor U10216 (N_10216,N_7851,N_8959);
xnor U10217 (N_10217,N_8812,N_7719);
or U10218 (N_10218,N_8193,N_8384);
or U10219 (N_10219,N_7567,N_7644);
nand U10220 (N_10220,N_7737,N_7626);
xor U10221 (N_10221,N_7855,N_8578);
and U10222 (N_10222,N_8442,N_8719);
nor U10223 (N_10223,N_8169,N_8411);
nor U10224 (N_10224,N_8369,N_8843);
nand U10225 (N_10225,N_8224,N_8728);
or U10226 (N_10226,N_8110,N_8949);
nand U10227 (N_10227,N_8752,N_8195);
and U10228 (N_10228,N_7833,N_7607);
xnor U10229 (N_10229,N_7559,N_8234);
nand U10230 (N_10230,N_7551,N_8754);
or U10231 (N_10231,N_7670,N_8500);
xnor U10232 (N_10232,N_8111,N_8590);
and U10233 (N_10233,N_8015,N_7532);
nor U10234 (N_10234,N_8536,N_8908);
or U10235 (N_10235,N_7731,N_8237);
nand U10236 (N_10236,N_8144,N_7815);
nand U10237 (N_10237,N_7580,N_8810);
and U10238 (N_10238,N_7510,N_7783);
nand U10239 (N_10239,N_8305,N_8932);
xor U10240 (N_10240,N_8583,N_7585);
nand U10241 (N_10241,N_8701,N_7937);
nor U10242 (N_10242,N_8136,N_8239);
and U10243 (N_10243,N_7589,N_8564);
xor U10244 (N_10244,N_7552,N_8152);
nor U10245 (N_10245,N_8951,N_8870);
and U10246 (N_10246,N_7879,N_7605);
or U10247 (N_10247,N_7536,N_8435);
and U10248 (N_10248,N_7882,N_8504);
or U10249 (N_10249,N_7571,N_7668);
or U10250 (N_10250,N_8280,N_8614);
or U10251 (N_10251,N_8627,N_8491);
or U10252 (N_10252,N_8878,N_8834);
or U10253 (N_10253,N_7507,N_8857);
xor U10254 (N_10254,N_8413,N_7918);
or U10255 (N_10255,N_8082,N_8298);
nor U10256 (N_10256,N_8767,N_8033);
nand U10257 (N_10257,N_7582,N_8513);
xnor U10258 (N_10258,N_8829,N_7897);
nor U10259 (N_10259,N_8346,N_8381);
xor U10260 (N_10260,N_7991,N_8003);
or U10261 (N_10261,N_7837,N_8039);
nor U10262 (N_10262,N_8515,N_8811);
or U10263 (N_10263,N_7846,N_8442);
nor U10264 (N_10264,N_8964,N_7528);
nand U10265 (N_10265,N_7515,N_8528);
nor U10266 (N_10266,N_8996,N_8222);
nand U10267 (N_10267,N_7636,N_7907);
or U10268 (N_10268,N_8112,N_8885);
or U10269 (N_10269,N_8416,N_7986);
and U10270 (N_10270,N_8153,N_7682);
nand U10271 (N_10271,N_8633,N_7883);
xor U10272 (N_10272,N_7787,N_7828);
or U10273 (N_10273,N_8247,N_8212);
nor U10274 (N_10274,N_8389,N_8947);
and U10275 (N_10275,N_8756,N_8277);
nand U10276 (N_10276,N_8346,N_8843);
nand U10277 (N_10277,N_7919,N_8726);
and U10278 (N_10278,N_8741,N_8951);
xor U10279 (N_10279,N_8326,N_8477);
nand U10280 (N_10280,N_8808,N_8041);
nor U10281 (N_10281,N_8578,N_7799);
and U10282 (N_10282,N_8310,N_8248);
and U10283 (N_10283,N_7703,N_8150);
nand U10284 (N_10284,N_7688,N_8202);
xor U10285 (N_10285,N_8078,N_8585);
nor U10286 (N_10286,N_7652,N_8688);
or U10287 (N_10287,N_8047,N_8641);
nand U10288 (N_10288,N_8792,N_8920);
or U10289 (N_10289,N_8282,N_7672);
xnor U10290 (N_10290,N_8267,N_7652);
and U10291 (N_10291,N_7538,N_8362);
or U10292 (N_10292,N_7896,N_8750);
nor U10293 (N_10293,N_8869,N_8612);
xnor U10294 (N_10294,N_7897,N_8992);
and U10295 (N_10295,N_7699,N_8645);
and U10296 (N_10296,N_7809,N_7552);
xnor U10297 (N_10297,N_8675,N_8142);
nand U10298 (N_10298,N_8155,N_7626);
nor U10299 (N_10299,N_8895,N_8890);
xnor U10300 (N_10300,N_7993,N_7922);
nor U10301 (N_10301,N_7740,N_7802);
or U10302 (N_10302,N_7616,N_8827);
and U10303 (N_10303,N_8965,N_8125);
and U10304 (N_10304,N_8349,N_8436);
nor U10305 (N_10305,N_8467,N_8686);
and U10306 (N_10306,N_8942,N_7608);
xor U10307 (N_10307,N_7732,N_7877);
nor U10308 (N_10308,N_8027,N_7855);
nand U10309 (N_10309,N_8899,N_8023);
or U10310 (N_10310,N_7992,N_8709);
and U10311 (N_10311,N_8273,N_8575);
or U10312 (N_10312,N_7551,N_8756);
or U10313 (N_10313,N_7750,N_8737);
or U10314 (N_10314,N_7664,N_7592);
and U10315 (N_10315,N_8451,N_7768);
and U10316 (N_10316,N_8892,N_8253);
nor U10317 (N_10317,N_8068,N_8142);
and U10318 (N_10318,N_8752,N_8029);
and U10319 (N_10319,N_7633,N_7501);
or U10320 (N_10320,N_8172,N_8530);
nor U10321 (N_10321,N_8073,N_8663);
nor U10322 (N_10322,N_8422,N_8008);
nor U10323 (N_10323,N_8154,N_7776);
and U10324 (N_10324,N_7980,N_7918);
and U10325 (N_10325,N_8912,N_7623);
nor U10326 (N_10326,N_8113,N_8941);
and U10327 (N_10327,N_8930,N_8411);
xnor U10328 (N_10328,N_7815,N_8512);
or U10329 (N_10329,N_8996,N_7749);
nand U10330 (N_10330,N_8567,N_8038);
and U10331 (N_10331,N_8347,N_8085);
xnor U10332 (N_10332,N_8494,N_8181);
or U10333 (N_10333,N_7689,N_8191);
nand U10334 (N_10334,N_8389,N_8141);
nand U10335 (N_10335,N_7960,N_8586);
or U10336 (N_10336,N_8577,N_8802);
and U10337 (N_10337,N_7759,N_8797);
nor U10338 (N_10338,N_8960,N_8605);
or U10339 (N_10339,N_7906,N_8947);
or U10340 (N_10340,N_8515,N_7525);
and U10341 (N_10341,N_7769,N_8322);
nand U10342 (N_10342,N_8121,N_8506);
nor U10343 (N_10343,N_8021,N_8462);
xor U10344 (N_10344,N_8229,N_8296);
nor U10345 (N_10345,N_8500,N_7726);
or U10346 (N_10346,N_8105,N_8006);
nand U10347 (N_10347,N_8095,N_7638);
nand U10348 (N_10348,N_8691,N_8898);
nand U10349 (N_10349,N_8510,N_7874);
xnor U10350 (N_10350,N_8324,N_8928);
and U10351 (N_10351,N_8224,N_8380);
nand U10352 (N_10352,N_8679,N_7521);
nand U10353 (N_10353,N_7683,N_8740);
and U10354 (N_10354,N_8192,N_7726);
nand U10355 (N_10355,N_7950,N_8245);
and U10356 (N_10356,N_7555,N_8140);
nand U10357 (N_10357,N_8697,N_7502);
xor U10358 (N_10358,N_8092,N_8664);
nor U10359 (N_10359,N_8181,N_7577);
xor U10360 (N_10360,N_8308,N_8986);
xnor U10361 (N_10361,N_8198,N_8160);
or U10362 (N_10362,N_7626,N_7850);
and U10363 (N_10363,N_8201,N_7557);
nand U10364 (N_10364,N_8048,N_8717);
nand U10365 (N_10365,N_7507,N_7757);
nor U10366 (N_10366,N_7660,N_8746);
nor U10367 (N_10367,N_7558,N_7764);
nand U10368 (N_10368,N_8487,N_8205);
or U10369 (N_10369,N_8040,N_8938);
or U10370 (N_10370,N_8207,N_8575);
and U10371 (N_10371,N_8259,N_7974);
or U10372 (N_10372,N_8377,N_7997);
xnor U10373 (N_10373,N_8392,N_8884);
xor U10374 (N_10374,N_8266,N_7502);
xnor U10375 (N_10375,N_8517,N_7526);
or U10376 (N_10376,N_8867,N_8839);
xnor U10377 (N_10377,N_8659,N_7772);
or U10378 (N_10378,N_7569,N_7844);
nor U10379 (N_10379,N_8585,N_8849);
or U10380 (N_10380,N_8407,N_8710);
and U10381 (N_10381,N_8817,N_8546);
xnor U10382 (N_10382,N_7949,N_8441);
xor U10383 (N_10383,N_8556,N_8346);
nand U10384 (N_10384,N_7880,N_7707);
and U10385 (N_10385,N_7577,N_7874);
nor U10386 (N_10386,N_8652,N_7845);
nor U10387 (N_10387,N_7921,N_8870);
xnor U10388 (N_10388,N_8393,N_8021);
nand U10389 (N_10389,N_8946,N_8227);
xnor U10390 (N_10390,N_7548,N_8257);
nand U10391 (N_10391,N_8083,N_8830);
nor U10392 (N_10392,N_8954,N_8766);
xor U10393 (N_10393,N_8673,N_8131);
nand U10394 (N_10394,N_8914,N_8936);
or U10395 (N_10395,N_8830,N_8230);
xnor U10396 (N_10396,N_7946,N_8240);
nor U10397 (N_10397,N_8487,N_8530);
xor U10398 (N_10398,N_8692,N_8025);
nand U10399 (N_10399,N_8972,N_8430);
xnor U10400 (N_10400,N_8507,N_8429);
xor U10401 (N_10401,N_8769,N_8266);
nand U10402 (N_10402,N_8877,N_8579);
nor U10403 (N_10403,N_7582,N_7834);
nor U10404 (N_10404,N_8012,N_7809);
and U10405 (N_10405,N_7914,N_7534);
and U10406 (N_10406,N_7890,N_7657);
nor U10407 (N_10407,N_8707,N_8508);
or U10408 (N_10408,N_7709,N_8030);
xor U10409 (N_10409,N_8675,N_8328);
nor U10410 (N_10410,N_8394,N_8869);
and U10411 (N_10411,N_7914,N_8402);
nor U10412 (N_10412,N_8662,N_8132);
or U10413 (N_10413,N_7991,N_8944);
and U10414 (N_10414,N_8969,N_8873);
xnor U10415 (N_10415,N_8199,N_8808);
nor U10416 (N_10416,N_7665,N_8830);
nor U10417 (N_10417,N_8507,N_8649);
xor U10418 (N_10418,N_8732,N_8241);
xnor U10419 (N_10419,N_8828,N_8348);
or U10420 (N_10420,N_8728,N_8718);
xor U10421 (N_10421,N_8149,N_8181);
nor U10422 (N_10422,N_8144,N_8091);
nor U10423 (N_10423,N_8930,N_8943);
nand U10424 (N_10424,N_7780,N_7965);
nor U10425 (N_10425,N_8103,N_8385);
and U10426 (N_10426,N_8669,N_7782);
and U10427 (N_10427,N_8557,N_8192);
and U10428 (N_10428,N_8023,N_8169);
or U10429 (N_10429,N_7630,N_8063);
and U10430 (N_10430,N_7773,N_8893);
and U10431 (N_10431,N_7703,N_8993);
and U10432 (N_10432,N_8622,N_7757);
nor U10433 (N_10433,N_8354,N_8686);
xor U10434 (N_10434,N_8204,N_8113);
or U10435 (N_10435,N_7986,N_7571);
nand U10436 (N_10436,N_8288,N_7671);
nor U10437 (N_10437,N_8683,N_8114);
nand U10438 (N_10438,N_8383,N_8945);
xnor U10439 (N_10439,N_8601,N_7559);
or U10440 (N_10440,N_7732,N_7710);
xor U10441 (N_10441,N_7693,N_7648);
nor U10442 (N_10442,N_8649,N_7632);
xnor U10443 (N_10443,N_8691,N_8538);
or U10444 (N_10444,N_8942,N_7954);
nor U10445 (N_10445,N_7972,N_7851);
xnor U10446 (N_10446,N_8610,N_8686);
nor U10447 (N_10447,N_8350,N_8790);
nand U10448 (N_10448,N_7613,N_8886);
nor U10449 (N_10449,N_8932,N_8351);
nor U10450 (N_10450,N_8393,N_8717);
and U10451 (N_10451,N_8430,N_7636);
nor U10452 (N_10452,N_7517,N_8802);
and U10453 (N_10453,N_7776,N_7595);
or U10454 (N_10454,N_8495,N_8519);
nand U10455 (N_10455,N_7714,N_7702);
nor U10456 (N_10456,N_8652,N_7584);
nand U10457 (N_10457,N_8295,N_8114);
or U10458 (N_10458,N_8428,N_8217);
nor U10459 (N_10459,N_8222,N_7717);
or U10460 (N_10460,N_8271,N_8305);
nor U10461 (N_10461,N_8636,N_7847);
or U10462 (N_10462,N_7742,N_7909);
nand U10463 (N_10463,N_8041,N_7853);
nand U10464 (N_10464,N_8144,N_8556);
and U10465 (N_10465,N_8743,N_8276);
nand U10466 (N_10466,N_7944,N_7994);
nor U10467 (N_10467,N_8316,N_8560);
and U10468 (N_10468,N_7773,N_8532);
nor U10469 (N_10469,N_8055,N_8016);
xnor U10470 (N_10470,N_8471,N_8928);
nor U10471 (N_10471,N_7628,N_7920);
and U10472 (N_10472,N_8544,N_8089);
or U10473 (N_10473,N_8793,N_7809);
nand U10474 (N_10474,N_8605,N_7966);
nand U10475 (N_10475,N_7702,N_7701);
and U10476 (N_10476,N_8190,N_8914);
nor U10477 (N_10477,N_7522,N_8512);
or U10478 (N_10478,N_8753,N_8736);
or U10479 (N_10479,N_8112,N_8880);
nand U10480 (N_10480,N_7613,N_8756);
xnor U10481 (N_10481,N_8372,N_8340);
or U10482 (N_10482,N_8706,N_8292);
nor U10483 (N_10483,N_7547,N_8952);
and U10484 (N_10484,N_8653,N_8013);
and U10485 (N_10485,N_8616,N_8132);
or U10486 (N_10486,N_7551,N_8562);
xnor U10487 (N_10487,N_7612,N_8243);
nor U10488 (N_10488,N_8594,N_8438);
or U10489 (N_10489,N_8939,N_8096);
nand U10490 (N_10490,N_8538,N_7648);
nor U10491 (N_10491,N_7806,N_7637);
and U10492 (N_10492,N_7747,N_7786);
and U10493 (N_10493,N_7595,N_7675);
and U10494 (N_10494,N_7965,N_7503);
xnor U10495 (N_10495,N_7724,N_8031);
or U10496 (N_10496,N_8952,N_7894);
or U10497 (N_10497,N_8841,N_7800);
nand U10498 (N_10498,N_7829,N_8652);
and U10499 (N_10499,N_8116,N_8752);
or U10500 (N_10500,N_9875,N_9641);
or U10501 (N_10501,N_9706,N_10355);
and U10502 (N_10502,N_9014,N_9694);
nor U10503 (N_10503,N_9374,N_10027);
and U10504 (N_10504,N_10286,N_10256);
xnor U10505 (N_10505,N_9792,N_9921);
nor U10506 (N_10506,N_9034,N_9254);
or U10507 (N_10507,N_9478,N_10270);
xor U10508 (N_10508,N_10324,N_10337);
nand U10509 (N_10509,N_10320,N_10438);
or U10510 (N_10510,N_9639,N_10087);
nand U10511 (N_10511,N_9215,N_9811);
nor U10512 (N_10512,N_9889,N_10301);
and U10513 (N_10513,N_9128,N_9633);
nor U10514 (N_10514,N_10460,N_10002);
nor U10515 (N_10515,N_9810,N_9760);
xor U10516 (N_10516,N_10451,N_9319);
xor U10517 (N_10517,N_9955,N_9020);
nor U10518 (N_10518,N_9076,N_10360);
and U10519 (N_10519,N_9525,N_9184);
or U10520 (N_10520,N_9189,N_10445);
or U10521 (N_10521,N_10261,N_9912);
and U10522 (N_10522,N_10212,N_9164);
or U10523 (N_10523,N_9488,N_9375);
xnor U10524 (N_10524,N_10044,N_9703);
and U10525 (N_10525,N_9585,N_9961);
or U10526 (N_10526,N_9172,N_10478);
nand U10527 (N_10527,N_10412,N_10466);
nand U10528 (N_10528,N_9753,N_9312);
nand U10529 (N_10529,N_9834,N_9166);
nand U10530 (N_10530,N_9995,N_9013);
nor U10531 (N_10531,N_10119,N_9502);
or U10532 (N_10532,N_10312,N_10202);
nand U10533 (N_10533,N_9770,N_9876);
nand U10534 (N_10534,N_9016,N_9945);
and U10535 (N_10535,N_10384,N_9039);
xnor U10536 (N_10536,N_10158,N_10439);
or U10537 (N_10537,N_9964,N_9606);
and U10538 (N_10538,N_10229,N_9984);
nor U10539 (N_10539,N_9649,N_9009);
nand U10540 (N_10540,N_9863,N_10054);
and U10541 (N_10541,N_10469,N_10463);
nand U10542 (N_10542,N_9381,N_10447);
or U10543 (N_10543,N_9569,N_10170);
nor U10544 (N_10544,N_9089,N_9594);
and U10545 (N_10545,N_10051,N_10189);
or U10546 (N_10546,N_9030,N_9890);
nor U10547 (N_10547,N_9678,N_9506);
nand U10548 (N_10548,N_9924,N_9808);
and U10549 (N_10549,N_10375,N_10306);
nor U10550 (N_10550,N_9860,N_9887);
xor U10551 (N_10551,N_9690,N_9870);
and U10552 (N_10552,N_9718,N_9747);
and U10553 (N_10553,N_9994,N_9864);
nand U10554 (N_10554,N_10258,N_9960);
xnor U10555 (N_10555,N_9515,N_9754);
xnor U10556 (N_10556,N_9247,N_9777);
nor U10557 (N_10557,N_9390,N_9714);
or U10558 (N_10558,N_9930,N_9445);
and U10559 (N_10559,N_9812,N_9993);
nor U10560 (N_10560,N_9534,N_9681);
xor U10561 (N_10561,N_9807,N_9441);
nand U10562 (N_10562,N_9361,N_9093);
and U10563 (N_10563,N_9310,N_9943);
xor U10564 (N_10564,N_9198,N_10461);
or U10565 (N_10565,N_9308,N_9344);
nor U10566 (N_10566,N_10369,N_9692);
nor U10567 (N_10567,N_10347,N_10486);
and U10568 (N_10568,N_9821,N_9384);
and U10569 (N_10569,N_9495,N_9952);
nand U10570 (N_10570,N_9556,N_9303);
xnor U10571 (N_10571,N_10275,N_9951);
or U10572 (N_10572,N_10175,N_10210);
and U10573 (N_10573,N_10146,N_10323);
and U10574 (N_10574,N_9925,N_9904);
xor U10575 (N_10575,N_9135,N_9200);
and U10576 (N_10576,N_9221,N_10017);
and U10577 (N_10577,N_9096,N_9829);
nor U10578 (N_10578,N_9919,N_10191);
nor U10579 (N_10579,N_9377,N_9241);
nor U10580 (N_10580,N_9800,N_9064);
and U10581 (N_10581,N_9433,N_9684);
xor U10582 (N_10582,N_10333,N_10030);
nand U10583 (N_10583,N_10271,N_9315);
nor U10584 (N_10584,N_9090,N_9607);
nand U10585 (N_10585,N_9263,N_9899);
or U10586 (N_10586,N_9918,N_9902);
and U10587 (N_10587,N_9956,N_9366);
and U10588 (N_10588,N_10183,N_9066);
and U10589 (N_10589,N_9163,N_10186);
and U10590 (N_10590,N_10105,N_9970);
and U10591 (N_10591,N_9405,N_10096);
nor U10592 (N_10592,N_9783,N_10366);
xnor U10593 (N_10593,N_9977,N_9492);
and U10594 (N_10594,N_9068,N_10276);
and U10595 (N_10595,N_9053,N_9493);
and U10596 (N_10596,N_10063,N_9469);
nor U10597 (N_10597,N_9350,N_10015);
or U10598 (N_10598,N_10321,N_9392);
and U10599 (N_10599,N_10381,N_9538);
and U10600 (N_10600,N_9679,N_9387);
or U10601 (N_10601,N_10200,N_10325);
nor U10602 (N_10602,N_9178,N_9192);
xnor U10603 (N_10603,N_9149,N_9815);
and U10604 (N_10604,N_9072,N_9612);
nor U10605 (N_10605,N_10101,N_10454);
or U10606 (N_10606,N_9082,N_9285);
nor U10607 (N_10607,N_10084,N_10185);
or U10608 (N_10608,N_9572,N_9954);
nor U10609 (N_10609,N_9471,N_9797);
nor U10610 (N_10610,N_10477,N_9443);
or U10611 (N_10611,N_9512,N_10058);
or U10612 (N_10612,N_9736,N_9647);
and U10613 (N_10613,N_9845,N_9982);
nor U10614 (N_10614,N_9081,N_10045);
nand U10615 (N_10615,N_9154,N_9903);
nand U10616 (N_10616,N_9909,N_9841);
nor U10617 (N_10617,N_9793,N_9541);
or U10618 (N_10618,N_10040,N_9202);
nand U10619 (N_10619,N_10340,N_9322);
nor U10620 (N_10620,N_9717,N_9171);
xor U10621 (N_10621,N_9865,N_9219);
nor U10622 (N_10622,N_9661,N_10223);
nand U10623 (N_10623,N_9599,N_9965);
xor U10624 (N_10624,N_10269,N_10348);
nand U10625 (N_10625,N_9332,N_9849);
or U10626 (N_10626,N_10442,N_9508);
or U10627 (N_10627,N_9179,N_10374);
and U10628 (N_10628,N_9734,N_10459);
and U10629 (N_10629,N_9153,N_9240);
xor U10630 (N_10630,N_9075,N_9762);
and U10631 (N_10631,N_9077,N_10211);
xnor U10632 (N_10632,N_9728,N_9839);
xor U10633 (N_10633,N_10273,N_9278);
xnor U10634 (N_10634,N_10310,N_9624);
nand U10635 (N_10635,N_10283,N_9386);
nor U10636 (N_10636,N_9522,N_9788);
nor U10637 (N_10637,N_9942,N_10471);
xor U10638 (N_10638,N_9722,N_9781);
and U10639 (N_10639,N_9050,N_10187);
and U10640 (N_10640,N_10007,N_10006);
xor U10641 (N_10641,N_9558,N_9414);
nand U10642 (N_10642,N_10025,N_10339);
nor U10643 (N_10643,N_9476,N_9527);
nor U10644 (N_10644,N_9677,N_9329);
xnor U10645 (N_10645,N_9004,N_10201);
nor U10646 (N_10646,N_10026,N_9091);
nor U10647 (N_10647,N_9699,N_9608);
xnor U10648 (N_10648,N_10431,N_9475);
and U10649 (N_10649,N_9877,N_9609);
xor U10650 (N_10650,N_10316,N_9098);
or U10651 (N_10651,N_10184,N_9395);
nor U10652 (N_10652,N_10385,N_9411);
nand U10653 (N_10653,N_9357,N_10497);
or U10654 (N_10654,N_9462,N_9022);
and U10655 (N_10655,N_9434,N_10233);
nor U10656 (N_10656,N_9500,N_10473);
xor U10657 (N_10657,N_9047,N_9752);
xnor U10658 (N_10658,N_10443,N_9638);
nand U10659 (N_10659,N_10068,N_9108);
or U10660 (N_10660,N_9321,N_10124);
nand U10661 (N_10661,N_9467,N_9258);
or U10662 (N_10662,N_10219,N_9518);
nand U10663 (N_10663,N_9397,N_9740);
nor U10664 (N_10664,N_9353,N_10050);
nor U10665 (N_10665,N_10126,N_9186);
or U10666 (N_10666,N_9057,N_9604);
xor U10667 (N_10667,N_10110,N_9819);
nand U10668 (N_10668,N_9209,N_10097);
xor U10669 (N_10669,N_10290,N_9528);
xnor U10670 (N_10670,N_9205,N_10246);
xor U10671 (N_10671,N_9517,N_10239);
and U10672 (N_10672,N_10247,N_9835);
nand U10673 (N_10673,N_9698,N_9972);
or U10674 (N_10674,N_9729,N_10484);
and U10675 (N_10675,N_9922,N_9360);
or U10676 (N_10676,N_10071,N_10254);
nor U10677 (N_10677,N_10047,N_9157);
and U10678 (N_10678,N_10335,N_10330);
and U10679 (N_10679,N_10091,N_10417);
or U10680 (N_10680,N_9891,N_9425);
nor U10681 (N_10681,N_9822,N_10259);
nor U10682 (N_10682,N_9803,N_10480);
xor U10683 (N_10683,N_9051,N_10425);
and U10684 (N_10684,N_10309,N_9006);
xnor U10685 (N_10685,N_9437,N_10117);
nor U10686 (N_10686,N_9228,N_10498);
nor U10687 (N_10687,N_10268,N_9653);
and U10688 (N_10688,N_9695,N_10193);
xor U10689 (N_10689,N_9813,N_9300);
or U10690 (N_10690,N_9622,N_10305);
and U10691 (N_10691,N_10428,N_9073);
or U10692 (N_10692,N_9011,N_9503);
nand U10693 (N_10693,N_9957,N_10038);
or U10694 (N_10694,N_9243,N_9393);
and U10695 (N_10695,N_9447,N_10372);
and U10696 (N_10696,N_10150,N_9814);
or U10697 (N_10697,N_9261,N_9646);
nand U10698 (N_10698,N_9148,N_9652);
xor U10699 (N_10699,N_10159,N_9620);
nor U10700 (N_10700,N_10132,N_10345);
or U10701 (N_10701,N_9268,N_10289);
nor U10702 (N_10702,N_9272,N_9771);
or U10703 (N_10703,N_9539,N_9174);
or U10704 (N_10704,N_9298,N_10382);
and U10705 (N_10705,N_9979,N_9496);
and U10706 (N_10706,N_9524,N_9432);
xnor U10707 (N_10707,N_9364,N_9936);
and U10708 (N_10708,N_9767,N_9037);
nor U10709 (N_10709,N_10231,N_10089);
xor U10710 (N_10710,N_10456,N_10476);
nand U10711 (N_10711,N_9005,N_9831);
and U10712 (N_10712,N_9547,N_9160);
xor U10713 (N_10713,N_9636,N_9761);
nand U10714 (N_10714,N_10238,N_9802);
nor U10715 (N_10715,N_9832,N_9230);
nand U10716 (N_10716,N_10147,N_9341);
nor U10717 (N_10717,N_9290,N_9061);
nor U10718 (N_10718,N_10332,N_9763);
nand U10719 (N_10719,N_9583,N_10216);
and U10720 (N_10720,N_10267,N_10465);
or U10721 (N_10721,N_9537,N_10042);
xor U10722 (N_10722,N_9029,N_9297);
nand U10723 (N_10723,N_9409,N_9289);
nor U10724 (N_10724,N_10169,N_9271);
nand U10725 (N_10725,N_9573,N_9378);
and U10726 (N_10726,N_9264,N_9826);
xor U10727 (N_10727,N_9025,N_10297);
nand U10728 (N_10728,N_9339,N_9670);
or U10729 (N_10729,N_9920,N_10397);
and U10730 (N_10730,N_10279,N_9246);
xnor U10731 (N_10731,N_9110,N_10336);
xor U10732 (N_10732,N_9233,N_9857);
nand U10733 (N_10733,N_9631,N_10052);
xnor U10734 (N_10734,N_9696,N_10444);
and U10735 (N_10735,N_9299,N_9749);
or U10736 (N_10736,N_9712,N_10421);
and U10737 (N_10737,N_9660,N_9349);
and U10738 (N_10738,N_10370,N_9355);
and U10739 (N_10739,N_9520,N_9719);
xor U10740 (N_10740,N_9133,N_9359);
nor U10741 (N_10741,N_9746,N_9852);
or U10742 (N_10742,N_9439,N_9844);
xor U10743 (N_10743,N_9766,N_9101);
and U10744 (N_10744,N_9223,N_9062);
and U10745 (N_10745,N_9112,N_10069);
xor U10746 (N_10746,N_9118,N_9182);
and U10747 (N_10747,N_9197,N_9893);
nor U10748 (N_10748,N_9309,N_9262);
xor U10749 (N_10749,N_10318,N_10149);
nor U10750 (N_10750,N_9369,N_9531);
and U10751 (N_10751,N_9060,N_10176);
or U10752 (N_10752,N_10075,N_9643);
or U10753 (N_10753,N_9741,N_9199);
xnor U10754 (N_10754,N_9545,N_10155);
nor U10755 (N_10755,N_9406,N_9083);
nand U10756 (N_10756,N_10224,N_9400);
and U10757 (N_10757,N_9046,N_9280);
xor U10758 (N_10758,N_9532,N_10489);
nand U10759 (N_10759,N_9867,N_9941);
xor U10760 (N_10760,N_9466,N_9778);
and U10761 (N_10761,N_9963,N_9743);
nand U10762 (N_10762,N_9824,N_9707);
nand U10763 (N_10763,N_9644,N_9235);
nand U10764 (N_10764,N_9126,N_9911);
xor U10765 (N_10765,N_9521,N_10319);
nand U10766 (N_10766,N_9551,N_10048);
or U10767 (N_10767,N_9983,N_10434);
nor U10768 (N_10768,N_9586,N_10103);
and U10769 (N_10769,N_9194,N_9627);
nor U10770 (N_10770,N_9772,N_9419);
nor U10771 (N_10771,N_9155,N_9931);
and U10772 (N_10772,N_9131,N_9894);
and U10773 (N_10773,N_9279,N_9104);
nor U10774 (N_10774,N_9914,N_9480);
and U10775 (N_10775,N_9146,N_10393);
nor U10776 (N_10776,N_9000,N_9313);
nand U10777 (N_10777,N_10144,N_10253);
and U10778 (N_10778,N_10196,N_9579);
nor U10779 (N_10779,N_9173,N_9474);
and U10780 (N_10780,N_9327,N_9837);
xnor U10781 (N_10781,N_10353,N_9785);
or U10782 (N_10782,N_9170,N_9769);
nor U10783 (N_10783,N_9431,N_9465);
or U10784 (N_10784,N_9328,N_9751);
or U10785 (N_10785,N_9630,N_10034);
nor U10786 (N_10786,N_10338,N_10359);
or U10787 (N_10787,N_9568,N_9702);
xor U10788 (N_10788,N_9600,N_9564);
and U10789 (N_10789,N_9727,N_10475);
and U10790 (N_10790,N_9152,N_9513);
or U10791 (N_10791,N_9723,N_9549);
or U10792 (N_10792,N_9017,N_10401);
xor U10793 (N_10793,N_9966,N_9129);
and U10794 (N_10794,N_9275,N_9122);
nor U10795 (N_10795,N_9428,N_10467);
and U10796 (N_10796,N_10221,N_9078);
and U10797 (N_10797,N_9204,N_10130);
and U10798 (N_10798,N_9358,N_9113);
and U10799 (N_10799,N_10298,N_10230);
and U10800 (N_10800,N_10127,N_10357);
nor U10801 (N_10801,N_10274,N_9097);
and U10802 (N_10802,N_9343,N_9399);
nor U10803 (N_10803,N_9255,N_9602);
xnor U10804 (N_10804,N_9658,N_9094);
or U10805 (N_10805,N_10423,N_9284);
nor U10806 (N_10806,N_9207,N_9331);
nor U10807 (N_10807,N_9473,N_10215);
or U10808 (N_10808,N_10013,N_9523);
or U10809 (N_10809,N_10361,N_10039);
and U10810 (N_10810,N_9711,N_9305);
xnor U10811 (N_10811,N_9337,N_10053);
nor U10812 (N_10812,N_10213,N_9950);
and U10813 (N_10813,N_9069,N_10161);
and U10814 (N_10814,N_9773,N_9861);
xnor U10815 (N_10815,N_9468,N_9107);
nor U10816 (N_10816,N_9806,N_9479);
and U10817 (N_10817,N_9725,N_10195);
xor U10818 (N_10818,N_9992,N_9898);
xor U10819 (N_10819,N_9838,N_10386);
nand U10820 (N_10820,N_10373,N_9637);
and U10821 (N_10821,N_10457,N_9906);
xnor U10822 (N_10822,N_10148,N_9888);
nand U10823 (N_10823,N_10118,N_9933);
xor U10824 (N_10824,N_10172,N_9124);
or U10825 (N_10825,N_10344,N_10018);
nor U10826 (N_10826,N_9043,N_9978);
or U10827 (N_10827,N_9997,N_9775);
nor U10828 (N_10828,N_9611,N_9333);
nor U10829 (N_10829,N_10019,N_9833);
and U10830 (N_10830,N_9851,N_9033);
and U10831 (N_10831,N_10171,N_10280);
xnor U10832 (N_10832,N_9916,N_9302);
nor U10833 (N_10833,N_9394,N_10303);
xor U10834 (N_10834,N_9932,N_10395);
nand U10835 (N_10835,N_10479,N_9042);
xor U10836 (N_10836,N_9231,N_9555);
nand U10837 (N_10837,N_9292,N_9372);
or U10838 (N_10838,N_10060,N_10099);
nand U10839 (N_10839,N_9985,N_10113);
xor U10840 (N_10840,N_10079,N_9563);
xnor U10841 (N_10841,N_10308,N_9910);
or U10842 (N_10842,N_9482,N_9974);
nand U10843 (N_10843,N_9580,N_9576);
and U10844 (N_10844,N_9915,N_9396);
nor U10845 (N_10845,N_9454,N_9415);
nand U10846 (N_10846,N_9288,N_9161);
and U10847 (N_10847,N_10046,N_10365);
nor U10848 (N_10848,N_9283,N_9382);
nor U10849 (N_10849,N_10227,N_9732);
nand U10850 (N_10850,N_9998,N_9413);
and U10851 (N_10851,N_9048,N_9176);
nand U10852 (N_10852,N_10173,N_10011);
and U10853 (N_10853,N_10236,N_9481);
nand U10854 (N_10854,N_10031,N_9085);
nand U10855 (N_10855,N_9621,N_9591);
nand U10856 (N_10856,N_9615,N_10432);
and U10857 (N_10857,N_9790,N_9351);
nand U10858 (N_10858,N_10426,N_10402);
nor U10859 (N_10859,N_9610,N_9947);
and U10860 (N_10860,N_9301,N_9429);
xor U10861 (N_10861,N_10093,N_10152);
or U10862 (N_10862,N_10495,N_9858);
or U10863 (N_10863,N_9407,N_9354);
or U10864 (N_10864,N_10488,N_9756);
or U10865 (N_10865,N_10419,N_10151);
or U10866 (N_10866,N_9566,N_10483);
and U10867 (N_10867,N_9656,N_9330);
xnor U10868 (N_10868,N_9973,N_9968);
and U10869 (N_10869,N_9487,N_9134);
or U10870 (N_10870,N_9498,N_9367);
xnor U10871 (N_10871,N_10367,N_9404);
xnor U10872 (N_10872,N_9457,N_10218);
or U10873 (N_10873,N_9137,N_10368);
nor U10874 (N_10874,N_10157,N_10041);
xnor U10875 (N_10875,N_10326,N_10288);
and U10876 (N_10876,N_10192,N_9926);
or U10877 (N_10877,N_9464,N_9071);
and U10878 (N_10878,N_9632,N_10278);
and U10879 (N_10879,N_9106,N_10154);
and U10880 (N_10880,N_9370,N_9165);
xor U10881 (N_10881,N_9680,N_9483);
nor U10882 (N_10882,N_9505,N_9765);
xnor U10883 (N_10883,N_9111,N_9217);
nand U10884 (N_10884,N_9939,N_9102);
and U10885 (N_10885,N_10204,N_9895);
and U10886 (N_10886,N_10086,N_9958);
or U10887 (N_10887,N_10115,N_9676);
xor U10888 (N_10888,N_9817,N_9206);
nand U10889 (N_10889,N_9195,N_9138);
or U10890 (N_10890,N_9969,N_10009);
or U10891 (N_10891,N_9590,N_9776);
and U10892 (N_10892,N_9981,N_10464);
or U10893 (N_10893,N_9614,N_9686);
nor U10894 (N_10894,N_9989,N_9444);
and U10895 (N_10895,N_9260,N_10028);
xnor U10896 (N_10896,N_9587,N_9224);
xor U10897 (N_10897,N_9873,N_9203);
xnor U10898 (N_10898,N_10265,N_10100);
nand U10899 (N_10899,N_9559,N_9052);
and U10900 (N_10900,N_9976,N_9099);
nor U10901 (N_10901,N_10036,N_9024);
nor U10902 (N_10902,N_10016,N_9946);
and U10903 (N_10903,N_10207,N_10410);
nand U10904 (N_10904,N_9724,N_10095);
or U10905 (N_10905,N_9323,N_9582);
and U10906 (N_10906,N_10424,N_9704);
nor U10907 (N_10907,N_9248,N_9459);
or U10908 (N_10908,N_9613,N_9581);
or U10909 (N_10909,N_9320,N_9818);
or U10910 (N_10910,N_10220,N_10356);
or U10911 (N_10911,N_10153,N_10134);
or U10912 (N_10912,N_9856,N_9509);
xor U10913 (N_10913,N_9150,N_9588);
or U10914 (N_10914,N_9533,N_9672);
nor U10915 (N_10915,N_9616,N_9340);
nor U10916 (N_10916,N_10263,N_9245);
nor U10917 (N_10917,N_10494,N_9356);
xor U10918 (N_10918,N_9380,N_9971);
or U10919 (N_10919,N_9028,N_9035);
xnor U10920 (N_10920,N_9901,N_10418);
nand U10921 (N_10921,N_9088,N_10329);
or U10922 (N_10922,N_9510,N_9570);
and U10923 (N_10923,N_9267,N_9561);
or U10924 (N_10924,N_9900,N_9731);
nand U10925 (N_10925,N_10379,N_9715);
nand U10926 (N_10926,N_10055,N_9748);
nand U10927 (N_10927,N_9416,N_9440);
or U10928 (N_10928,N_9368,N_10142);
or U10929 (N_10929,N_9940,N_9923);
xnor U10930 (N_10930,N_9234,N_10065);
xnor U10931 (N_10931,N_9764,N_10021);
and U10932 (N_10932,N_9125,N_9687);
nand U10933 (N_10933,N_9226,N_10123);
nor U10934 (N_10934,N_10299,N_9239);
nand U10935 (N_10935,N_10203,N_10088);
xnor U10936 (N_10936,N_10449,N_10394);
xor U10937 (N_10937,N_10435,N_10346);
and U10938 (N_10938,N_9352,N_9501);
or U10939 (N_10939,N_10217,N_9675);
and U10940 (N_10940,N_10328,N_9683);
or U10941 (N_10941,N_9140,N_9705);
or U10942 (N_10942,N_9874,N_10197);
xnor U10943 (N_10943,N_9143,N_10433);
nand U10944 (N_10944,N_9449,N_9557);
and U10945 (N_10945,N_9023,N_9169);
and U10946 (N_10946,N_9012,N_9634);
and U10947 (N_10947,N_10413,N_9371);
xor U10948 (N_10948,N_9281,N_9823);
nor U10949 (N_10949,N_9674,N_9688);
and U10950 (N_10950,N_9529,N_10237);
or U10951 (N_10951,N_10085,N_10057);
and U10952 (N_10952,N_10104,N_10090);
xor U10953 (N_10953,N_9002,N_9345);
or U10954 (N_10954,N_9026,N_9571);
nor U10955 (N_10955,N_9780,N_9121);
nand U10956 (N_10956,N_10094,N_10188);
nand U10957 (N_10957,N_10262,N_9036);
nand U10958 (N_10958,N_9848,N_9187);
and U10959 (N_10959,N_10129,N_9786);
or U10960 (N_10960,N_10436,N_9908);
xnor U10961 (N_10961,N_9058,N_9391);
or U10962 (N_10962,N_9490,N_9259);
and U10963 (N_10963,N_9768,N_9991);
nor U10964 (N_10964,N_10241,N_9750);
nand U10965 (N_10965,N_9123,N_10168);
xnor U10966 (N_10966,N_9436,N_9809);
and U10967 (N_10967,N_10005,N_9342);
nor U10968 (N_10968,N_10307,N_9842);
nand U10969 (N_10969,N_10448,N_9779);
xor U10970 (N_10970,N_9516,N_9801);
xnor U10971 (N_10971,N_9491,N_10264);
nand U10972 (N_10972,N_9190,N_9304);
or U10973 (N_10973,N_9990,N_9866);
nor U10974 (N_10974,N_9376,N_10351);
nand U10975 (N_10975,N_10214,N_10266);
nand U10976 (N_10976,N_9544,N_10177);
xor U10977 (N_10977,N_9162,N_10180);
or U10978 (N_10978,N_10243,N_9645);
nand U10979 (N_10979,N_9147,N_9663);
nor U10980 (N_10980,N_9257,N_10371);
or U10981 (N_10981,N_9054,N_10121);
xnor U10982 (N_10982,N_9074,N_9132);
xnor U10983 (N_10983,N_10491,N_9212);
and U10984 (N_10984,N_9237,N_9536);
and U10985 (N_10985,N_9913,N_10092);
xor U10986 (N_10986,N_9010,N_10114);
or U10987 (N_10987,N_9167,N_9063);
nor U10988 (N_10988,N_9252,N_9242);
xor U10989 (N_10989,N_9774,N_10206);
and U10990 (N_10990,N_9499,N_9458);
xor U10991 (N_10991,N_9019,N_10455);
nor U10992 (N_10992,N_9548,N_9603);
xor U10993 (N_10993,N_9791,N_9697);
nand U10994 (N_10994,N_9408,N_9338);
nor U10995 (N_10995,N_9735,N_9648);
xnor U10996 (N_10996,N_10076,N_9363);
nand U10997 (N_10997,N_10074,N_9759);
nor U10998 (N_10998,N_9862,N_9015);
xnor U10999 (N_10999,N_9032,N_9999);
and U11000 (N_11000,N_10285,N_9287);
nor U11001 (N_11001,N_10391,N_9794);
nand U11002 (N_11002,N_9145,N_9045);
nand U11003 (N_11003,N_9084,N_9623);
nand U11004 (N_11004,N_10139,N_9196);
and U11005 (N_11005,N_10077,N_9070);
nor U11006 (N_11006,N_10392,N_9949);
nor U11007 (N_11007,N_9494,N_9018);
or U11008 (N_11008,N_9412,N_9087);
or U11009 (N_11009,N_9141,N_9871);
nand U11010 (N_11010,N_9185,N_9882);
nand U11011 (N_11011,N_9424,N_9701);
xor U11012 (N_11012,N_9673,N_9847);
nor U11013 (N_11013,N_10378,N_9250);
nand U11014 (N_11014,N_10472,N_9136);
nand U11015 (N_11015,N_10295,N_10403);
or U11016 (N_11016,N_10458,N_9008);
and U11017 (N_11017,N_9535,N_9626);
nand U11018 (N_11018,N_10341,N_9448);
and U11019 (N_11019,N_9193,N_9804);
and U11020 (N_11020,N_9745,N_9593);
or U11021 (N_11021,N_9177,N_9709);
xor U11022 (N_11022,N_9755,N_9489);
or U11023 (N_11023,N_9619,N_9886);
or U11024 (N_11024,N_9067,N_9757);
nand U11025 (N_11025,N_9092,N_10416);
nand U11026 (N_11026,N_9325,N_10492);
nand U11027 (N_11027,N_10125,N_9244);
and U11028 (N_11028,N_10493,N_9552);
xor U11029 (N_11029,N_9827,N_9530);
xnor U11030 (N_11030,N_9859,N_9805);
xor U11031 (N_11031,N_9151,N_10317);
nor U11032 (N_11032,N_10427,N_9317);
xor U11033 (N_11033,N_10001,N_10066);
nor U11034 (N_11034,N_9100,N_10122);
or U11035 (N_11035,N_9843,N_10205);
and U11036 (N_11036,N_9335,N_9987);
or U11037 (N_11037,N_9980,N_9456);
and U11038 (N_11038,N_9739,N_9389);
or U11039 (N_11039,N_10240,N_9651);
and U11040 (N_11040,N_9055,N_10165);
xor U11041 (N_11041,N_9159,N_9846);
or U11042 (N_11042,N_9575,N_9379);
and U11043 (N_11043,N_9210,N_10225);
or U11044 (N_11044,N_9038,N_9383);
nand U11045 (N_11045,N_9975,N_10334);
xnor U11046 (N_11046,N_9659,N_10198);
nor U11047 (N_11047,N_9540,N_10049);
nand U11048 (N_11048,N_10004,N_9472);
xor U11049 (N_11049,N_10342,N_10377);
and U11050 (N_11050,N_9546,N_9056);
xnor U11051 (N_11051,N_10160,N_9708);
or U11052 (N_11052,N_10422,N_10112);
or U11053 (N_11053,N_9795,N_10429);
nand U11054 (N_11054,N_9507,N_10081);
nor U11055 (N_11055,N_10404,N_10181);
and U11056 (N_11056,N_10242,N_9435);
xor U11057 (N_11057,N_10248,N_9021);
and U11058 (N_11058,N_10228,N_9286);
or U11059 (N_11059,N_10327,N_9721);
and U11060 (N_11060,N_10078,N_10499);
or U11061 (N_11061,N_9276,N_9742);
or U11062 (N_11062,N_9666,N_9825);
xor U11063 (N_11063,N_9334,N_9744);
or U11064 (N_11064,N_9884,N_10226);
nor U11065 (N_11065,N_9324,N_9988);
or U11066 (N_11066,N_10272,N_10490);
xor U11067 (N_11067,N_9589,N_9403);
or U11068 (N_11068,N_9117,N_10029);
and U11069 (N_11069,N_10362,N_9455);
or U11070 (N_11070,N_10293,N_9617);
or U11071 (N_11071,N_10302,N_9927);
or U11072 (N_11072,N_9928,N_10108);
nand U11073 (N_11073,N_10363,N_9907);
and U11074 (N_11074,N_9139,N_9421);
nor U11075 (N_11075,N_9080,N_10143);
and U11076 (N_11076,N_9295,N_9574);
or U11077 (N_11077,N_10440,N_10389);
nor U11078 (N_11078,N_10138,N_9664);
xnor U11079 (N_11079,N_10311,N_9840);
nor U11080 (N_11080,N_10080,N_9935);
or U11081 (N_11081,N_9450,N_9385);
xor U11082 (N_11082,N_10485,N_10407);
nor U11083 (N_11083,N_9642,N_9282);
and U11084 (N_11084,N_9417,N_10234);
nor U11085 (N_11085,N_9142,N_9402);
and U11086 (N_11086,N_10481,N_9578);
nor U11087 (N_11087,N_10315,N_9365);
nand U11088 (N_11088,N_9269,N_9655);
nand U11089 (N_11089,N_10010,N_9040);
or U11090 (N_11090,N_9650,N_9461);
xnor U11091 (N_11091,N_9597,N_10178);
or U11092 (N_11092,N_9996,N_9986);
nor U11093 (N_11093,N_10167,N_9225);
xor U11094 (N_11094,N_10387,N_9562);
nand U11095 (N_11095,N_9962,N_9306);
nor U11096 (N_11096,N_10163,N_10136);
xor U11097 (N_11097,N_9291,N_10462);
nand U11098 (N_11098,N_9191,N_9789);
or U11099 (N_11099,N_9730,N_10061);
xnor U11100 (N_11100,N_9253,N_9486);
or U11101 (N_11101,N_9892,N_9662);
or U11102 (N_11102,N_9446,N_10352);
nor U11103 (N_11103,N_10414,N_9116);
and U11104 (N_11104,N_9896,N_10450);
xnor U11105 (N_11105,N_9318,N_9592);
nor U11106 (N_11106,N_10287,N_9959);
and U11107 (N_11107,N_9307,N_9553);
nand U11108 (N_11108,N_10383,N_9868);
nor U11109 (N_11109,N_9629,N_10400);
or U11110 (N_11110,N_10420,N_10037);
xnor U11111 (N_11111,N_9693,N_9504);
nand U11112 (N_11112,N_9216,N_10260);
or U11113 (N_11113,N_9640,N_9869);
nand U11114 (N_11114,N_10453,N_9422);
or U11115 (N_11115,N_9336,N_9249);
and U11116 (N_11116,N_9878,N_9273);
xnor U11117 (N_11117,N_10070,N_9758);
nor U11118 (N_11118,N_10067,N_9463);
and U11119 (N_11119,N_10406,N_10174);
nand U11120 (N_11120,N_10032,N_9682);
xor U11121 (N_11121,N_9885,N_10282);
nor U11122 (N_11122,N_9526,N_10331);
or U11123 (N_11123,N_9452,N_9836);
nor U11124 (N_11124,N_10194,N_10082);
xor U11125 (N_11125,N_9671,N_10249);
xor U11126 (N_11126,N_10141,N_9850);
xor U11127 (N_11127,N_10250,N_9897);
xor U11128 (N_11128,N_10468,N_10222);
or U11129 (N_11129,N_10380,N_9872);
and U11130 (N_11130,N_10043,N_9917);
or U11131 (N_11131,N_9944,N_9181);
nor U11132 (N_11132,N_9460,N_10140);
nand U11133 (N_11133,N_9420,N_10452);
or U11134 (N_11134,N_9348,N_9514);
xor U11135 (N_11135,N_9737,N_10376);
or U11136 (N_11136,N_9543,N_10496);
nand U11137 (N_11137,N_9266,N_10209);
or U11138 (N_11138,N_9109,N_9937);
and U11139 (N_11139,N_9733,N_9044);
nand U11140 (N_11140,N_9086,N_9625);
and U11141 (N_11141,N_10350,N_10343);
nand U11142 (N_11142,N_10245,N_9426);
nand U11143 (N_11143,N_10145,N_9628);
or U11144 (N_11144,N_10251,N_10291);
or U11145 (N_11145,N_9059,N_9183);
or U11146 (N_11146,N_10137,N_9427);
or U11147 (N_11147,N_9373,N_10014);
and U11148 (N_11148,N_9784,N_9880);
xnor U11149 (N_11149,N_9031,N_9550);
xor U11150 (N_11150,N_9713,N_10128);
and U11151 (N_11151,N_10304,N_9601);
xnor U11152 (N_11152,N_10277,N_9554);
or U11153 (N_11153,N_9314,N_9477);
or U11154 (N_11154,N_10441,N_9595);
xnor U11155 (N_11155,N_10257,N_10179);
nor U11156 (N_11156,N_9883,N_10244);
and U11157 (N_11157,N_10072,N_9401);
nand U11158 (N_11158,N_10358,N_10411);
nand U11159 (N_11159,N_9929,N_10232);
xor U11160 (N_11160,N_9236,N_9855);
xnor U11161 (N_11161,N_10296,N_9738);
nor U11162 (N_11162,N_9214,N_10349);
or U11163 (N_11163,N_10156,N_10023);
nand U11164 (N_11164,N_9201,N_10199);
nand U11165 (N_11165,N_9953,N_9103);
nor U11166 (N_11166,N_10064,N_10252);
or U11167 (N_11167,N_10281,N_9618);
xor U11168 (N_11168,N_9438,N_9423);
nor U11169 (N_11169,N_9685,N_9665);
xnor U11170 (N_11170,N_10408,N_9222);
or U11171 (N_11171,N_10059,N_10003);
nor U11172 (N_11172,N_9451,N_9229);
and U11173 (N_11173,N_10398,N_9798);
xor U11174 (N_11174,N_10182,N_9347);
xnor U11175 (N_11175,N_9605,N_9114);
or U11176 (N_11176,N_9854,N_9079);
nor U11177 (N_11177,N_9565,N_9277);
xor U11178 (N_11178,N_9001,N_10482);
and U11179 (N_11179,N_9716,N_9519);
xor U11180 (N_11180,N_9938,N_9232);
or U11181 (N_11181,N_10020,N_9208);
or U11182 (N_11182,N_9567,N_9720);
nand U11183 (N_11183,N_9796,N_10396);
and U11184 (N_11184,N_9657,N_9596);
or U11185 (N_11185,N_9294,N_10409);
and U11186 (N_11186,N_9027,N_10111);
xor U11187 (N_11187,N_9710,N_10035);
or U11188 (N_11188,N_9853,N_9828);
nand U11189 (N_11189,N_9691,N_10284);
or U11190 (N_11190,N_9388,N_10133);
or U11191 (N_11191,N_9003,N_10000);
or U11192 (N_11192,N_10388,N_9346);
or U11193 (N_11193,N_10313,N_9293);
nor U11194 (N_11194,N_10116,N_9584);
nor U11195 (N_11195,N_10109,N_9256);
and U11196 (N_11196,N_10437,N_9296);
nor U11197 (N_11197,N_9485,N_10107);
nand U11198 (N_11198,N_9180,N_9635);
nor U11199 (N_11199,N_10430,N_10131);
and U11200 (N_11200,N_10073,N_10390);
nand U11201 (N_11201,N_9654,N_9948);
nand U11202 (N_11202,N_9442,N_9453);
or U11203 (N_11203,N_9158,N_9667);
nand U11204 (N_11204,N_10314,N_9238);
or U11205 (N_11205,N_9119,N_10405);
xor U11206 (N_11206,N_9065,N_9816);
or U11207 (N_11207,N_10208,N_9049);
and U11208 (N_11208,N_10294,N_10012);
xor U11209 (N_11209,N_10102,N_9095);
nand U11210 (N_11210,N_9175,N_9218);
nand U11211 (N_11211,N_9041,N_9311);
nor U11212 (N_11212,N_10292,N_9115);
and U11213 (N_11213,N_9007,N_10033);
xor U11214 (N_11214,N_9220,N_10487);
xnor U11215 (N_11215,N_9362,N_10166);
xor U11216 (N_11216,N_10354,N_9787);
and U11217 (N_11217,N_10008,N_9251);
xnor U11218 (N_11218,N_9211,N_9398);
nand U11219 (N_11219,N_9484,N_9726);
xor U11220 (N_11220,N_9120,N_9410);
nand U11221 (N_11221,N_9270,N_10056);
nand U11222 (N_11222,N_9188,N_9577);
xnor U11223 (N_11223,N_9669,N_10446);
nand U11224 (N_11224,N_9967,N_9497);
nand U11225 (N_11225,N_9156,N_10190);
nand U11226 (N_11226,N_10024,N_10098);
xor U11227 (N_11227,N_9144,N_9881);
nand U11228 (N_11228,N_10364,N_9274);
xor U11229 (N_11229,N_9905,N_9168);
nand U11230 (N_11230,N_9418,N_9830);
nor U11231 (N_11231,N_9227,N_9130);
or U11232 (N_11232,N_9668,N_9470);
xnor U11233 (N_11233,N_9879,N_10022);
nand U11234 (N_11234,N_10120,N_10415);
and U11235 (N_11235,N_10083,N_9265);
nor U11236 (N_11236,N_9560,N_9213);
nand U11237 (N_11237,N_10162,N_10300);
or U11238 (N_11238,N_9598,N_9127);
nor U11239 (N_11239,N_10470,N_9782);
and U11240 (N_11240,N_10062,N_10322);
or U11241 (N_11241,N_9316,N_9326);
xnor U11242 (N_11242,N_10135,N_9542);
xor U11243 (N_11243,N_9700,N_10106);
xnor U11244 (N_11244,N_10235,N_9511);
nor U11245 (N_11245,N_10474,N_9430);
nor U11246 (N_11246,N_9799,N_9934);
xor U11247 (N_11247,N_10164,N_9820);
xnor U11248 (N_11248,N_9689,N_10255);
nor U11249 (N_11249,N_9105,N_10399);
and U11250 (N_11250,N_9125,N_10307);
nand U11251 (N_11251,N_10468,N_9195);
nor U11252 (N_11252,N_9564,N_9782);
and U11253 (N_11253,N_10199,N_9675);
or U11254 (N_11254,N_10395,N_9473);
and U11255 (N_11255,N_9666,N_9145);
or U11256 (N_11256,N_9768,N_10393);
nand U11257 (N_11257,N_9147,N_9595);
xnor U11258 (N_11258,N_9298,N_10153);
xnor U11259 (N_11259,N_9610,N_10217);
xor U11260 (N_11260,N_9485,N_9284);
nor U11261 (N_11261,N_9967,N_9407);
nand U11262 (N_11262,N_9106,N_9000);
or U11263 (N_11263,N_9567,N_10305);
nor U11264 (N_11264,N_10002,N_9320);
and U11265 (N_11265,N_10240,N_9365);
nor U11266 (N_11266,N_10108,N_9263);
nor U11267 (N_11267,N_9031,N_9036);
nand U11268 (N_11268,N_10470,N_10012);
nor U11269 (N_11269,N_9859,N_10419);
xor U11270 (N_11270,N_9703,N_9739);
nand U11271 (N_11271,N_9419,N_9520);
or U11272 (N_11272,N_9470,N_9619);
xor U11273 (N_11273,N_10391,N_9945);
xnor U11274 (N_11274,N_9536,N_9439);
nor U11275 (N_11275,N_10050,N_10464);
or U11276 (N_11276,N_9899,N_10353);
nor U11277 (N_11277,N_10244,N_10229);
nand U11278 (N_11278,N_9898,N_10205);
nor U11279 (N_11279,N_10436,N_9679);
nand U11280 (N_11280,N_9264,N_9102);
nor U11281 (N_11281,N_10282,N_10443);
nand U11282 (N_11282,N_9999,N_10392);
nand U11283 (N_11283,N_9799,N_10442);
and U11284 (N_11284,N_10487,N_10330);
nand U11285 (N_11285,N_10318,N_9882);
and U11286 (N_11286,N_9027,N_10041);
nand U11287 (N_11287,N_9655,N_9517);
and U11288 (N_11288,N_9302,N_10452);
and U11289 (N_11289,N_10317,N_9720);
or U11290 (N_11290,N_9031,N_9859);
or U11291 (N_11291,N_9260,N_9131);
nand U11292 (N_11292,N_9627,N_9150);
nand U11293 (N_11293,N_10464,N_10467);
xor U11294 (N_11294,N_10496,N_10163);
xor U11295 (N_11295,N_9577,N_10404);
nor U11296 (N_11296,N_9948,N_10274);
nand U11297 (N_11297,N_9460,N_9534);
or U11298 (N_11298,N_9568,N_9312);
nand U11299 (N_11299,N_9794,N_9155);
or U11300 (N_11300,N_10208,N_9408);
nand U11301 (N_11301,N_10188,N_9752);
or U11302 (N_11302,N_9049,N_9937);
or U11303 (N_11303,N_10316,N_9775);
or U11304 (N_11304,N_10057,N_9845);
nor U11305 (N_11305,N_9899,N_10180);
xor U11306 (N_11306,N_10078,N_10406);
xnor U11307 (N_11307,N_9209,N_9656);
nor U11308 (N_11308,N_9392,N_10446);
nand U11309 (N_11309,N_9251,N_10346);
nand U11310 (N_11310,N_9420,N_10276);
or U11311 (N_11311,N_9965,N_10212);
nand U11312 (N_11312,N_10472,N_10157);
and U11313 (N_11313,N_9864,N_9858);
and U11314 (N_11314,N_9624,N_9670);
and U11315 (N_11315,N_10328,N_9648);
nor U11316 (N_11316,N_9541,N_9154);
and U11317 (N_11317,N_10294,N_10309);
nand U11318 (N_11318,N_9782,N_9755);
nor U11319 (N_11319,N_9861,N_9016);
and U11320 (N_11320,N_10059,N_9928);
nand U11321 (N_11321,N_9204,N_10068);
xor U11322 (N_11322,N_9637,N_9631);
nor U11323 (N_11323,N_9344,N_10168);
xnor U11324 (N_11324,N_9261,N_9766);
and U11325 (N_11325,N_9280,N_9571);
nor U11326 (N_11326,N_9386,N_9288);
nor U11327 (N_11327,N_9869,N_9475);
nor U11328 (N_11328,N_10157,N_10119);
and U11329 (N_11329,N_9457,N_9894);
nor U11330 (N_11330,N_9960,N_10043);
and U11331 (N_11331,N_9052,N_9084);
and U11332 (N_11332,N_10124,N_10232);
nor U11333 (N_11333,N_9045,N_10236);
nand U11334 (N_11334,N_9144,N_9773);
nor U11335 (N_11335,N_9670,N_9146);
xor U11336 (N_11336,N_9632,N_9124);
or U11337 (N_11337,N_9168,N_10486);
xnor U11338 (N_11338,N_9486,N_10147);
or U11339 (N_11339,N_10251,N_9566);
nand U11340 (N_11340,N_9013,N_9466);
and U11341 (N_11341,N_9143,N_9509);
and U11342 (N_11342,N_10287,N_9804);
nand U11343 (N_11343,N_10227,N_9375);
nor U11344 (N_11344,N_9217,N_9175);
nor U11345 (N_11345,N_9675,N_9523);
nor U11346 (N_11346,N_9985,N_10218);
and U11347 (N_11347,N_9108,N_9780);
xnor U11348 (N_11348,N_9210,N_9791);
nand U11349 (N_11349,N_9381,N_9177);
or U11350 (N_11350,N_9326,N_9451);
xor U11351 (N_11351,N_9785,N_10481);
xor U11352 (N_11352,N_9586,N_9140);
or U11353 (N_11353,N_10272,N_9289);
xnor U11354 (N_11354,N_9806,N_9800);
nor U11355 (N_11355,N_9148,N_10091);
and U11356 (N_11356,N_10348,N_9578);
xnor U11357 (N_11357,N_9181,N_9652);
xor U11358 (N_11358,N_9089,N_9442);
nand U11359 (N_11359,N_10141,N_9392);
xnor U11360 (N_11360,N_9566,N_9184);
nor U11361 (N_11361,N_9131,N_10061);
or U11362 (N_11362,N_9838,N_9757);
and U11363 (N_11363,N_9039,N_9964);
or U11364 (N_11364,N_9154,N_10069);
nor U11365 (N_11365,N_10299,N_9001);
and U11366 (N_11366,N_10062,N_9031);
and U11367 (N_11367,N_9782,N_9327);
nor U11368 (N_11368,N_10243,N_9948);
or U11369 (N_11369,N_9807,N_9561);
or U11370 (N_11370,N_9898,N_9924);
xor U11371 (N_11371,N_9312,N_10422);
or U11372 (N_11372,N_9910,N_9783);
nand U11373 (N_11373,N_9622,N_10243);
xnor U11374 (N_11374,N_10087,N_9423);
xnor U11375 (N_11375,N_9223,N_9274);
nand U11376 (N_11376,N_9095,N_9987);
xor U11377 (N_11377,N_9567,N_9328);
and U11378 (N_11378,N_10231,N_9012);
nand U11379 (N_11379,N_9526,N_10056);
and U11380 (N_11380,N_9651,N_10017);
or U11381 (N_11381,N_9173,N_10194);
nor U11382 (N_11382,N_9104,N_10297);
nand U11383 (N_11383,N_9722,N_10078);
nor U11384 (N_11384,N_9390,N_9305);
and U11385 (N_11385,N_10226,N_9381);
nor U11386 (N_11386,N_10015,N_9314);
nand U11387 (N_11387,N_9310,N_9256);
nor U11388 (N_11388,N_9142,N_9810);
nor U11389 (N_11389,N_10168,N_9134);
xnor U11390 (N_11390,N_9313,N_10159);
or U11391 (N_11391,N_9731,N_9089);
nor U11392 (N_11392,N_10456,N_9958);
and U11393 (N_11393,N_9232,N_9337);
nor U11394 (N_11394,N_10287,N_10251);
xor U11395 (N_11395,N_9090,N_10403);
xnor U11396 (N_11396,N_9569,N_9407);
nor U11397 (N_11397,N_10403,N_10046);
or U11398 (N_11398,N_9033,N_10413);
xnor U11399 (N_11399,N_9559,N_9530);
xor U11400 (N_11400,N_9254,N_9136);
nor U11401 (N_11401,N_9796,N_9686);
nor U11402 (N_11402,N_10275,N_10186);
nand U11403 (N_11403,N_10192,N_10168);
nor U11404 (N_11404,N_9881,N_9406);
xnor U11405 (N_11405,N_9421,N_10491);
xor U11406 (N_11406,N_10151,N_9152);
xor U11407 (N_11407,N_9957,N_9624);
and U11408 (N_11408,N_9920,N_9124);
nand U11409 (N_11409,N_10473,N_9085);
or U11410 (N_11410,N_9177,N_9388);
xnor U11411 (N_11411,N_9325,N_10463);
nand U11412 (N_11412,N_9081,N_9556);
and U11413 (N_11413,N_9613,N_9491);
nor U11414 (N_11414,N_10219,N_10445);
nand U11415 (N_11415,N_9649,N_9761);
nand U11416 (N_11416,N_9103,N_9964);
or U11417 (N_11417,N_10359,N_9787);
and U11418 (N_11418,N_10216,N_10359);
xor U11419 (N_11419,N_9984,N_9739);
nor U11420 (N_11420,N_9892,N_9792);
nor U11421 (N_11421,N_10261,N_9186);
nand U11422 (N_11422,N_9879,N_10485);
or U11423 (N_11423,N_9704,N_10375);
nand U11424 (N_11424,N_9532,N_10140);
nor U11425 (N_11425,N_9635,N_9684);
nor U11426 (N_11426,N_9020,N_9162);
or U11427 (N_11427,N_9373,N_9441);
xor U11428 (N_11428,N_10415,N_9799);
and U11429 (N_11429,N_10378,N_10192);
and U11430 (N_11430,N_9306,N_10261);
and U11431 (N_11431,N_9421,N_9852);
or U11432 (N_11432,N_9934,N_9105);
or U11433 (N_11433,N_9822,N_10394);
or U11434 (N_11434,N_9362,N_9676);
and U11435 (N_11435,N_9335,N_10470);
nand U11436 (N_11436,N_10219,N_9496);
xor U11437 (N_11437,N_10123,N_9623);
and U11438 (N_11438,N_9426,N_10322);
xor U11439 (N_11439,N_9234,N_10486);
or U11440 (N_11440,N_9897,N_9733);
or U11441 (N_11441,N_10312,N_9980);
nand U11442 (N_11442,N_10175,N_9415);
or U11443 (N_11443,N_10274,N_10126);
nand U11444 (N_11444,N_9278,N_10303);
xnor U11445 (N_11445,N_10446,N_10493);
and U11446 (N_11446,N_9277,N_10472);
or U11447 (N_11447,N_9174,N_9762);
and U11448 (N_11448,N_10418,N_10140);
xnor U11449 (N_11449,N_9334,N_9093);
and U11450 (N_11450,N_9117,N_9014);
or U11451 (N_11451,N_9933,N_9178);
nand U11452 (N_11452,N_9202,N_9383);
and U11453 (N_11453,N_9830,N_10465);
nand U11454 (N_11454,N_9981,N_10371);
nand U11455 (N_11455,N_10213,N_9674);
nand U11456 (N_11456,N_9040,N_9202);
nor U11457 (N_11457,N_9117,N_10108);
and U11458 (N_11458,N_9363,N_9634);
nor U11459 (N_11459,N_9470,N_10155);
or U11460 (N_11460,N_10161,N_9712);
and U11461 (N_11461,N_10256,N_9513);
nor U11462 (N_11462,N_9151,N_9318);
xnor U11463 (N_11463,N_9350,N_10300);
nand U11464 (N_11464,N_10158,N_9533);
nor U11465 (N_11465,N_10273,N_9912);
and U11466 (N_11466,N_10274,N_9048);
xor U11467 (N_11467,N_9653,N_9135);
and U11468 (N_11468,N_9746,N_9323);
and U11469 (N_11469,N_9310,N_10050);
and U11470 (N_11470,N_9074,N_9264);
xor U11471 (N_11471,N_9786,N_9924);
xor U11472 (N_11472,N_10216,N_9911);
or U11473 (N_11473,N_9802,N_9979);
or U11474 (N_11474,N_9087,N_9409);
xnor U11475 (N_11475,N_9132,N_9337);
nor U11476 (N_11476,N_9600,N_9966);
nor U11477 (N_11477,N_9168,N_10098);
nand U11478 (N_11478,N_9562,N_9045);
nor U11479 (N_11479,N_10048,N_10262);
nand U11480 (N_11480,N_10008,N_9681);
xnor U11481 (N_11481,N_9019,N_9795);
or U11482 (N_11482,N_9878,N_10006);
nand U11483 (N_11483,N_10291,N_9840);
xnor U11484 (N_11484,N_10271,N_9735);
or U11485 (N_11485,N_9319,N_9160);
or U11486 (N_11486,N_10205,N_9974);
and U11487 (N_11487,N_9732,N_10020);
nor U11488 (N_11488,N_10379,N_10326);
nand U11489 (N_11489,N_9015,N_9505);
nand U11490 (N_11490,N_10221,N_9669);
nand U11491 (N_11491,N_10028,N_10061);
xnor U11492 (N_11492,N_9901,N_9845);
and U11493 (N_11493,N_9602,N_9935);
nand U11494 (N_11494,N_10145,N_10140);
or U11495 (N_11495,N_9333,N_10121);
xor U11496 (N_11496,N_10199,N_9396);
or U11497 (N_11497,N_9269,N_9457);
nand U11498 (N_11498,N_9510,N_9110);
xnor U11499 (N_11499,N_9357,N_9562);
xnor U11500 (N_11500,N_9418,N_9643);
or U11501 (N_11501,N_10243,N_10060);
and U11502 (N_11502,N_10171,N_10083);
xnor U11503 (N_11503,N_10252,N_9008);
or U11504 (N_11504,N_10062,N_10323);
and U11505 (N_11505,N_10037,N_9965);
nand U11506 (N_11506,N_10354,N_9244);
and U11507 (N_11507,N_9402,N_9981);
xor U11508 (N_11508,N_9638,N_9195);
or U11509 (N_11509,N_10284,N_9966);
and U11510 (N_11510,N_9535,N_10218);
nand U11511 (N_11511,N_9496,N_10245);
and U11512 (N_11512,N_10349,N_10075);
nand U11513 (N_11513,N_9677,N_9373);
or U11514 (N_11514,N_9784,N_9401);
or U11515 (N_11515,N_10146,N_9855);
nand U11516 (N_11516,N_9295,N_9668);
or U11517 (N_11517,N_10350,N_9435);
or U11518 (N_11518,N_9571,N_9650);
and U11519 (N_11519,N_9697,N_10381);
nand U11520 (N_11520,N_9466,N_10166);
and U11521 (N_11521,N_10476,N_10109);
nand U11522 (N_11522,N_10089,N_9131);
xor U11523 (N_11523,N_9736,N_9799);
and U11524 (N_11524,N_10092,N_9127);
and U11525 (N_11525,N_9584,N_10320);
or U11526 (N_11526,N_9645,N_10372);
nand U11527 (N_11527,N_9646,N_9803);
xor U11528 (N_11528,N_9151,N_10298);
xnor U11529 (N_11529,N_9839,N_9732);
nand U11530 (N_11530,N_9044,N_9900);
nand U11531 (N_11531,N_9298,N_10085);
nand U11532 (N_11532,N_9834,N_9892);
and U11533 (N_11533,N_9672,N_9519);
and U11534 (N_11534,N_9678,N_10274);
nand U11535 (N_11535,N_9721,N_9860);
xor U11536 (N_11536,N_9471,N_9380);
nor U11537 (N_11537,N_9280,N_9750);
nor U11538 (N_11538,N_9645,N_10384);
or U11539 (N_11539,N_9294,N_10011);
nor U11540 (N_11540,N_9708,N_9175);
or U11541 (N_11541,N_9215,N_10397);
or U11542 (N_11542,N_9158,N_9278);
xnor U11543 (N_11543,N_10299,N_9834);
nand U11544 (N_11544,N_9358,N_9521);
nand U11545 (N_11545,N_10431,N_9880);
nor U11546 (N_11546,N_9651,N_9148);
and U11547 (N_11547,N_9373,N_9619);
xnor U11548 (N_11548,N_9434,N_9325);
xor U11549 (N_11549,N_9010,N_9572);
xor U11550 (N_11550,N_9829,N_10240);
xnor U11551 (N_11551,N_9323,N_9125);
nor U11552 (N_11552,N_10146,N_9211);
nand U11553 (N_11553,N_10247,N_10477);
and U11554 (N_11554,N_10411,N_9197);
or U11555 (N_11555,N_10264,N_9275);
or U11556 (N_11556,N_9412,N_9295);
nand U11557 (N_11557,N_9168,N_10456);
nand U11558 (N_11558,N_9602,N_9632);
nor U11559 (N_11559,N_10264,N_9895);
and U11560 (N_11560,N_9243,N_9569);
and U11561 (N_11561,N_10330,N_9478);
nand U11562 (N_11562,N_10081,N_9131);
or U11563 (N_11563,N_9047,N_9529);
and U11564 (N_11564,N_9255,N_10373);
and U11565 (N_11565,N_9996,N_9615);
nor U11566 (N_11566,N_9017,N_10202);
nand U11567 (N_11567,N_9248,N_10230);
xor U11568 (N_11568,N_9134,N_10440);
or U11569 (N_11569,N_9771,N_10384);
nand U11570 (N_11570,N_9813,N_10158);
nand U11571 (N_11571,N_10275,N_10138);
and U11572 (N_11572,N_10477,N_9732);
and U11573 (N_11573,N_9477,N_10319);
nor U11574 (N_11574,N_9414,N_9224);
nand U11575 (N_11575,N_10141,N_9913);
or U11576 (N_11576,N_9092,N_9401);
or U11577 (N_11577,N_9550,N_10073);
nand U11578 (N_11578,N_10360,N_10033);
nand U11579 (N_11579,N_10400,N_9913);
nand U11580 (N_11580,N_9884,N_9719);
xnor U11581 (N_11581,N_9751,N_9533);
and U11582 (N_11582,N_10216,N_9393);
xnor U11583 (N_11583,N_9744,N_9080);
xor U11584 (N_11584,N_10304,N_9525);
nand U11585 (N_11585,N_9588,N_9130);
nand U11586 (N_11586,N_9574,N_9379);
and U11587 (N_11587,N_10068,N_9139);
nand U11588 (N_11588,N_9028,N_9555);
nand U11589 (N_11589,N_9408,N_9772);
nand U11590 (N_11590,N_10016,N_10189);
or U11591 (N_11591,N_9533,N_10115);
nand U11592 (N_11592,N_9128,N_9150);
xnor U11593 (N_11593,N_9109,N_9060);
or U11594 (N_11594,N_10169,N_9134);
and U11595 (N_11595,N_10441,N_9584);
xor U11596 (N_11596,N_9204,N_9061);
and U11597 (N_11597,N_10313,N_9438);
or U11598 (N_11598,N_9750,N_10270);
nor U11599 (N_11599,N_9370,N_9970);
xor U11600 (N_11600,N_9048,N_9018);
xor U11601 (N_11601,N_10025,N_9262);
xnor U11602 (N_11602,N_9426,N_10180);
and U11603 (N_11603,N_9001,N_10214);
or U11604 (N_11604,N_10331,N_9652);
and U11605 (N_11605,N_10433,N_9860);
nor U11606 (N_11606,N_10226,N_9301);
xor U11607 (N_11607,N_9121,N_10148);
xnor U11608 (N_11608,N_10066,N_9541);
xor U11609 (N_11609,N_9294,N_9466);
and U11610 (N_11610,N_10490,N_10211);
nor U11611 (N_11611,N_10191,N_9987);
or U11612 (N_11612,N_9755,N_9875);
nor U11613 (N_11613,N_10128,N_9563);
xnor U11614 (N_11614,N_10095,N_10131);
or U11615 (N_11615,N_9821,N_10433);
nor U11616 (N_11616,N_9453,N_9993);
nor U11617 (N_11617,N_9546,N_9016);
and U11618 (N_11618,N_9497,N_10116);
nor U11619 (N_11619,N_9556,N_9449);
nor U11620 (N_11620,N_9264,N_10143);
nand U11621 (N_11621,N_10044,N_9891);
xor U11622 (N_11622,N_10326,N_10200);
nor U11623 (N_11623,N_10452,N_10095);
nand U11624 (N_11624,N_10164,N_9080);
and U11625 (N_11625,N_9315,N_9753);
and U11626 (N_11626,N_10148,N_9574);
or U11627 (N_11627,N_10495,N_10000);
xnor U11628 (N_11628,N_10412,N_9992);
and U11629 (N_11629,N_9063,N_9238);
or U11630 (N_11630,N_9037,N_9931);
nand U11631 (N_11631,N_9714,N_9729);
nor U11632 (N_11632,N_9067,N_9360);
xnor U11633 (N_11633,N_9169,N_9809);
nor U11634 (N_11634,N_10434,N_9200);
xnor U11635 (N_11635,N_9758,N_9720);
nor U11636 (N_11636,N_9585,N_10140);
or U11637 (N_11637,N_10114,N_10014);
or U11638 (N_11638,N_10264,N_10184);
or U11639 (N_11639,N_9755,N_9473);
xor U11640 (N_11640,N_9211,N_9544);
or U11641 (N_11641,N_9400,N_9869);
nand U11642 (N_11642,N_9959,N_10049);
nor U11643 (N_11643,N_9915,N_9594);
xor U11644 (N_11644,N_9565,N_9322);
and U11645 (N_11645,N_10481,N_9272);
nor U11646 (N_11646,N_9929,N_9062);
nor U11647 (N_11647,N_9085,N_9396);
and U11648 (N_11648,N_9976,N_9384);
or U11649 (N_11649,N_9164,N_10130);
nor U11650 (N_11650,N_10360,N_9577);
nor U11651 (N_11651,N_9539,N_9477);
xnor U11652 (N_11652,N_10473,N_10101);
nand U11653 (N_11653,N_10237,N_9991);
xnor U11654 (N_11654,N_9320,N_9906);
nand U11655 (N_11655,N_10378,N_9918);
xnor U11656 (N_11656,N_9706,N_10211);
nor U11657 (N_11657,N_9816,N_10474);
xnor U11658 (N_11658,N_9341,N_10335);
nor U11659 (N_11659,N_9250,N_10138);
nor U11660 (N_11660,N_10287,N_9169);
and U11661 (N_11661,N_9376,N_9853);
nand U11662 (N_11662,N_9609,N_10468);
and U11663 (N_11663,N_10198,N_9684);
or U11664 (N_11664,N_9922,N_9093);
and U11665 (N_11665,N_10183,N_10237);
nand U11666 (N_11666,N_10373,N_9739);
nor U11667 (N_11667,N_9944,N_10262);
nand U11668 (N_11668,N_9888,N_10087);
or U11669 (N_11669,N_9980,N_10185);
nor U11670 (N_11670,N_10008,N_10428);
xnor U11671 (N_11671,N_10140,N_10064);
nand U11672 (N_11672,N_10081,N_9918);
or U11673 (N_11673,N_9086,N_9679);
xor U11674 (N_11674,N_9691,N_9873);
nor U11675 (N_11675,N_9830,N_9000);
and U11676 (N_11676,N_10171,N_10057);
nand U11677 (N_11677,N_9849,N_10093);
and U11678 (N_11678,N_9917,N_9563);
xor U11679 (N_11679,N_10131,N_9648);
nand U11680 (N_11680,N_10057,N_9754);
or U11681 (N_11681,N_10071,N_10192);
xor U11682 (N_11682,N_10092,N_9872);
nand U11683 (N_11683,N_10448,N_10423);
xnor U11684 (N_11684,N_9978,N_10083);
nand U11685 (N_11685,N_9744,N_9673);
or U11686 (N_11686,N_9086,N_9256);
xnor U11687 (N_11687,N_9217,N_9979);
and U11688 (N_11688,N_9701,N_9464);
nor U11689 (N_11689,N_9982,N_9471);
nand U11690 (N_11690,N_10231,N_10288);
nand U11691 (N_11691,N_10040,N_9337);
nand U11692 (N_11692,N_9962,N_9286);
and U11693 (N_11693,N_9593,N_9731);
and U11694 (N_11694,N_9896,N_9048);
nor U11695 (N_11695,N_10329,N_9778);
or U11696 (N_11696,N_10372,N_9386);
or U11697 (N_11697,N_9348,N_10490);
xnor U11698 (N_11698,N_10017,N_9528);
xor U11699 (N_11699,N_10411,N_9908);
and U11700 (N_11700,N_9245,N_9534);
and U11701 (N_11701,N_9527,N_9721);
or U11702 (N_11702,N_10412,N_9218);
or U11703 (N_11703,N_9370,N_10371);
or U11704 (N_11704,N_9929,N_9400);
or U11705 (N_11705,N_9127,N_9137);
and U11706 (N_11706,N_10469,N_9139);
and U11707 (N_11707,N_10111,N_9259);
or U11708 (N_11708,N_10436,N_10332);
xor U11709 (N_11709,N_10416,N_9775);
and U11710 (N_11710,N_9613,N_9601);
and U11711 (N_11711,N_10339,N_9405);
xor U11712 (N_11712,N_9723,N_10051);
xor U11713 (N_11713,N_9611,N_9403);
nor U11714 (N_11714,N_10278,N_10411);
and U11715 (N_11715,N_9891,N_10360);
nand U11716 (N_11716,N_9057,N_9236);
nand U11717 (N_11717,N_10026,N_10372);
nand U11718 (N_11718,N_9916,N_9458);
and U11719 (N_11719,N_9619,N_10149);
xnor U11720 (N_11720,N_9505,N_9017);
nand U11721 (N_11721,N_9463,N_10238);
and U11722 (N_11722,N_9179,N_10411);
or U11723 (N_11723,N_10314,N_10171);
and U11724 (N_11724,N_9579,N_10447);
nor U11725 (N_11725,N_9611,N_10159);
or U11726 (N_11726,N_9528,N_9750);
nand U11727 (N_11727,N_10213,N_9663);
nand U11728 (N_11728,N_9819,N_9623);
and U11729 (N_11729,N_10391,N_9700);
and U11730 (N_11730,N_9137,N_9403);
xnor U11731 (N_11731,N_9683,N_9348);
nand U11732 (N_11732,N_10309,N_9860);
nand U11733 (N_11733,N_9392,N_9583);
nand U11734 (N_11734,N_9342,N_10061);
or U11735 (N_11735,N_9311,N_9509);
xnor U11736 (N_11736,N_10464,N_9312);
or U11737 (N_11737,N_9034,N_9062);
nand U11738 (N_11738,N_10161,N_9748);
and U11739 (N_11739,N_9162,N_10097);
nor U11740 (N_11740,N_9441,N_9329);
or U11741 (N_11741,N_9598,N_10421);
xnor U11742 (N_11742,N_10425,N_9366);
or U11743 (N_11743,N_9634,N_9019);
or U11744 (N_11744,N_9794,N_9034);
nor U11745 (N_11745,N_10476,N_9663);
nor U11746 (N_11746,N_10197,N_9147);
and U11747 (N_11747,N_9472,N_9935);
nor U11748 (N_11748,N_9286,N_9103);
nor U11749 (N_11749,N_9910,N_9224);
and U11750 (N_11750,N_9045,N_10113);
and U11751 (N_11751,N_9403,N_9475);
nor U11752 (N_11752,N_9640,N_10419);
xor U11753 (N_11753,N_9653,N_9612);
nor U11754 (N_11754,N_10080,N_9839);
xor U11755 (N_11755,N_9050,N_10379);
nor U11756 (N_11756,N_9912,N_9876);
nand U11757 (N_11757,N_9633,N_9062);
and U11758 (N_11758,N_9289,N_9065);
or U11759 (N_11759,N_10276,N_9761);
xor U11760 (N_11760,N_9646,N_9013);
xnor U11761 (N_11761,N_10485,N_9558);
nand U11762 (N_11762,N_10247,N_10485);
and U11763 (N_11763,N_9719,N_9198);
and U11764 (N_11764,N_10359,N_9437);
and U11765 (N_11765,N_9029,N_10496);
and U11766 (N_11766,N_9475,N_10302);
nor U11767 (N_11767,N_9201,N_10218);
or U11768 (N_11768,N_10204,N_10060);
nor U11769 (N_11769,N_9654,N_10405);
nor U11770 (N_11770,N_10298,N_10085);
xnor U11771 (N_11771,N_9907,N_9012);
nand U11772 (N_11772,N_10375,N_9483);
and U11773 (N_11773,N_9791,N_9118);
nor U11774 (N_11774,N_9437,N_9264);
nor U11775 (N_11775,N_9085,N_10428);
nor U11776 (N_11776,N_9835,N_9313);
nand U11777 (N_11777,N_9689,N_9696);
and U11778 (N_11778,N_10375,N_9415);
and U11779 (N_11779,N_9122,N_9638);
nand U11780 (N_11780,N_9117,N_9008);
or U11781 (N_11781,N_9874,N_10280);
and U11782 (N_11782,N_9891,N_9901);
nor U11783 (N_11783,N_9959,N_9843);
and U11784 (N_11784,N_9387,N_10413);
nand U11785 (N_11785,N_9415,N_9900);
xor U11786 (N_11786,N_10335,N_9780);
nor U11787 (N_11787,N_9037,N_9346);
and U11788 (N_11788,N_9442,N_9379);
xor U11789 (N_11789,N_10146,N_9095);
or U11790 (N_11790,N_10294,N_10470);
or U11791 (N_11791,N_9773,N_9295);
xnor U11792 (N_11792,N_9851,N_10437);
and U11793 (N_11793,N_9402,N_9713);
nand U11794 (N_11794,N_10321,N_9326);
xor U11795 (N_11795,N_9063,N_10137);
xnor U11796 (N_11796,N_9627,N_9665);
nor U11797 (N_11797,N_10111,N_10325);
or U11798 (N_11798,N_9619,N_9521);
xor U11799 (N_11799,N_10179,N_9268);
nand U11800 (N_11800,N_10036,N_9107);
xor U11801 (N_11801,N_10079,N_9158);
nand U11802 (N_11802,N_10312,N_10189);
xnor U11803 (N_11803,N_10273,N_9406);
nor U11804 (N_11804,N_10428,N_9117);
xnor U11805 (N_11805,N_9449,N_9487);
nand U11806 (N_11806,N_9612,N_9641);
xnor U11807 (N_11807,N_9931,N_9090);
xor U11808 (N_11808,N_9174,N_10149);
xnor U11809 (N_11809,N_9657,N_10387);
nand U11810 (N_11810,N_10219,N_9766);
xor U11811 (N_11811,N_9535,N_9398);
or U11812 (N_11812,N_9447,N_10461);
nand U11813 (N_11813,N_9619,N_9495);
or U11814 (N_11814,N_9319,N_9907);
nand U11815 (N_11815,N_9780,N_9398);
or U11816 (N_11816,N_10470,N_9409);
nor U11817 (N_11817,N_9678,N_10109);
xor U11818 (N_11818,N_9676,N_9850);
nor U11819 (N_11819,N_9561,N_9814);
or U11820 (N_11820,N_9858,N_9280);
nor U11821 (N_11821,N_10123,N_10103);
xor U11822 (N_11822,N_9013,N_9057);
and U11823 (N_11823,N_9989,N_9480);
or U11824 (N_11824,N_9063,N_9309);
nand U11825 (N_11825,N_9215,N_9703);
or U11826 (N_11826,N_10257,N_9763);
or U11827 (N_11827,N_10174,N_9113);
nor U11828 (N_11828,N_9186,N_9195);
and U11829 (N_11829,N_9084,N_9273);
and U11830 (N_11830,N_10204,N_9190);
or U11831 (N_11831,N_9379,N_9104);
nor U11832 (N_11832,N_9369,N_9216);
nand U11833 (N_11833,N_10079,N_9550);
nor U11834 (N_11834,N_9031,N_9538);
xnor U11835 (N_11835,N_9156,N_9044);
nand U11836 (N_11836,N_9715,N_10263);
and U11837 (N_11837,N_9181,N_9903);
nand U11838 (N_11838,N_10027,N_9525);
nand U11839 (N_11839,N_10306,N_9462);
and U11840 (N_11840,N_9829,N_9720);
xnor U11841 (N_11841,N_10205,N_10148);
and U11842 (N_11842,N_10000,N_10098);
nor U11843 (N_11843,N_9455,N_9069);
or U11844 (N_11844,N_9573,N_9480);
or U11845 (N_11845,N_10314,N_9539);
nor U11846 (N_11846,N_9232,N_10469);
or U11847 (N_11847,N_9838,N_10311);
xor U11848 (N_11848,N_10494,N_10373);
and U11849 (N_11849,N_9944,N_9284);
nand U11850 (N_11850,N_9313,N_9995);
and U11851 (N_11851,N_9755,N_10181);
or U11852 (N_11852,N_9696,N_10429);
xor U11853 (N_11853,N_10263,N_9523);
or U11854 (N_11854,N_9571,N_10053);
or U11855 (N_11855,N_9160,N_10133);
nor U11856 (N_11856,N_9910,N_9562);
or U11857 (N_11857,N_9980,N_9427);
nor U11858 (N_11858,N_10197,N_9452);
and U11859 (N_11859,N_10105,N_10078);
or U11860 (N_11860,N_9622,N_9426);
and U11861 (N_11861,N_9204,N_9931);
nor U11862 (N_11862,N_10221,N_9782);
or U11863 (N_11863,N_9500,N_10143);
nand U11864 (N_11864,N_10307,N_10098);
xnor U11865 (N_11865,N_9154,N_9146);
nand U11866 (N_11866,N_9244,N_9215);
xor U11867 (N_11867,N_9102,N_9294);
and U11868 (N_11868,N_9514,N_9612);
and U11869 (N_11869,N_10474,N_10477);
nor U11870 (N_11870,N_9238,N_9507);
nor U11871 (N_11871,N_9264,N_9459);
xor U11872 (N_11872,N_10070,N_9333);
nor U11873 (N_11873,N_10120,N_9271);
or U11874 (N_11874,N_9999,N_9487);
nor U11875 (N_11875,N_10046,N_9990);
nor U11876 (N_11876,N_9852,N_9050);
and U11877 (N_11877,N_10474,N_10066);
xnor U11878 (N_11878,N_9818,N_10427);
or U11879 (N_11879,N_9315,N_9676);
or U11880 (N_11880,N_9053,N_9616);
nand U11881 (N_11881,N_9415,N_9573);
and U11882 (N_11882,N_9463,N_10117);
nand U11883 (N_11883,N_9670,N_10066);
xnor U11884 (N_11884,N_10139,N_9502);
nand U11885 (N_11885,N_10031,N_9362);
xor U11886 (N_11886,N_10306,N_9045);
or U11887 (N_11887,N_10030,N_9162);
nand U11888 (N_11888,N_10039,N_9974);
or U11889 (N_11889,N_9656,N_9517);
and U11890 (N_11890,N_9640,N_9302);
nand U11891 (N_11891,N_9988,N_9458);
xnor U11892 (N_11892,N_10429,N_10320);
nand U11893 (N_11893,N_9420,N_9506);
nor U11894 (N_11894,N_10001,N_9520);
xor U11895 (N_11895,N_10246,N_9658);
xor U11896 (N_11896,N_10357,N_9977);
nor U11897 (N_11897,N_10417,N_9761);
or U11898 (N_11898,N_9766,N_10388);
or U11899 (N_11899,N_10084,N_9203);
and U11900 (N_11900,N_9978,N_10132);
nor U11901 (N_11901,N_9536,N_9872);
or U11902 (N_11902,N_9854,N_9602);
xor U11903 (N_11903,N_9087,N_10299);
and U11904 (N_11904,N_10082,N_9246);
or U11905 (N_11905,N_10231,N_10199);
and U11906 (N_11906,N_10464,N_9244);
or U11907 (N_11907,N_9690,N_9478);
and U11908 (N_11908,N_9140,N_9889);
nor U11909 (N_11909,N_9449,N_10200);
xnor U11910 (N_11910,N_10310,N_10056);
nor U11911 (N_11911,N_9937,N_10021);
nor U11912 (N_11912,N_10385,N_9226);
nand U11913 (N_11913,N_10028,N_9323);
xnor U11914 (N_11914,N_9093,N_9076);
and U11915 (N_11915,N_9023,N_9184);
nor U11916 (N_11916,N_10204,N_9951);
xnor U11917 (N_11917,N_10483,N_9098);
xnor U11918 (N_11918,N_9006,N_9392);
and U11919 (N_11919,N_10178,N_9393);
xor U11920 (N_11920,N_10238,N_10047);
xor U11921 (N_11921,N_9235,N_9985);
xor U11922 (N_11922,N_9233,N_10053);
nor U11923 (N_11923,N_10159,N_10178);
nor U11924 (N_11924,N_9925,N_9830);
and U11925 (N_11925,N_9028,N_9356);
nor U11926 (N_11926,N_9482,N_9714);
and U11927 (N_11927,N_9825,N_10324);
and U11928 (N_11928,N_9848,N_9878);
or U11929 (N_11929,N_10405,N_9026);
or U11930 (N_11930,N_10428,N_10134);
nand U11931 (N_11931,N_10113,N_9864);
nor U11932 (N_11932,N_9090,N_9542);
nand U11933 (N_11933,N_10181,N_9527);
and U11934 (N_11934,N_9985,N_9848);
nand U11935 (N_11935,N_10012,N_9059);
and U11936 (N_11936,N_9101,N_10059);
nor U11937 (N_11937,N_9925,N_10028);
nand U11938 (N_11938,N_10315,N_10007);
xor U11939 (N_11939,N_10352,N_9004);
xor U11940 (N_11940,N_9907,N_9634);
nand U11941 (N_11941,N_9596,N_10008);
or U11942 (N_11942,N_10040,N_9373);
and U11943 (N_11943,N_9528,N_10083);
xor U11944 (N_11944,N_9648,N_10332);
or U11945 (N_11945,N_9192,N_9200);
xor U11946 (N_11946,N_10147,N_9045);
and U11947 (N_11947,N_10156,N_9509);
and U11948 (N_11948,N_9959,N_10316);
and U11949 (N_11949,N_10363,N_9410);
xnor U11950 (N_11950,N_9214,N_9872);
or U11951 (N_11951,N_10347,N_9641);
xor U11952 (N_11952,N_9776,N_9406);
nor U11953 (N_11953,N_9561,N_10475);
nor U11954 (N_11954,N_9164,N_10078);
and U11955 (N_11955,N_10405,N_9430);
nor U11956 (N_11956,N_9823,N_9901);
nor U11957 (N_11957,N_9159,N_10425);
and U11958 (N_11958,N_9663,N_9343);
or U11959 (N_11959,N_10256,N_9012);
nand U11960 (N_11960,N_9239,N_9318);
nor U11961 (N_11961,N_10212,N_10265);
or U11962 (N_11962,N_9924,N_10212);
xnor U11963 (N_11963,N_9209,N_9931);
nand U11964 (N_11964,N_10338,N_9840);
nand U11965 (N_11965,N_9694,N_10244);
nand U11966 (N_11966,N_9988,N_9686);
or U11967 (N_11967,N_9418,N_9433);
nand U11968 (N_11968,N_10188,N_9036);
nor U11969 (N_11969,N_10350,N_10189);
xor U11970 (N_11970,N_9694,N_9108);
xnor U11971 (N_11971,N_10190,N_9660);
nor U11972 (N_11972,N_10425,N_9878);
and U11973 (N_11973,N_10197,N_10342);
nand U11974 (N_11974,N_9230,N_10432);
xor U11975 (N_11975,N_9026,N_10399);
and U11976 (N_11976,N_9766,N_9246);
xor U11977 (N_11977,N_9300,N_9273);
xnor U11978 (N_11978,N_9346,N_9180);
nor U11979 (N_11979,N_9755,N_10083);
nor U11980 (N_11980,N_9578,N_10291);
and U11981 (N_11981,N_9044,N_9160);
nand U11982 (N_11982,N_9717,N_9404);
nor U11983 (N_11983,N_9129,N_9584);
or U11984 (N_11984,N_9780,N_10407);
nor U11985 (N_11985,N_9363,N_10185);
or U11986 (N_11986,N_9151,N_9066);
xor U11987 (N_11987,N_9500,N_9565);
nand U11988 (N_11988,N_10192,N_9834);
and U11989 (N_11989,N_10307,N_10266);
and U11990 (N_11990,N_9925,N_9094);
nor U11991 (N_11991,N_10397,N_10120);
nor U11992 (N_11992,N_10141,N_9113);
xor U11993 (N_11993,N_9788,N_10465);
nor U11994 (N_11994,N_9560,N_10107);
or U11995 (N_11995,N_10224,N_9448);
xor U11996 (N_11996,N_9638,N_9227);
and U11997 (N_11997,N_9448,N_10032);
xnor U11998 (N_11998,N_10465,N_9669);
xnor U11999 (N_11999,N_9548,N_9096);
nand U12000 (N_12000,N_10644,N_11522);
xor U12001 (N_12001,N_11206,N_10817);
and U12002 (N_12002,N_10830,N_11667);
nand U12003 (N_12003,N_11567,N_11038);
or U12004 (N_12004,N_11329,N_10931);
or U12005 (N_12005,N_11287,N_10752);
xnor U12006 (N_12006,N_10839,N_11128);
nand U12007 (N_12007,N_10678,N_11670);
nor U12008 (N_12008,N_10670,N_11968);
nor U12009 (N_12009,N_11118,N_10946);
xnor U12010 (N_12010,N_11074,N_10833);
nand U12011 (N_12011,N_10914,N_10733);
nand U12012 (N_12012,N_11191,N_11883);
nand U12013 (N_12013,N_11070,N_11894);
nor U12014 (N_12014,N_10951,N_11490);
nor U12015 (N_12015,N_11426,N_10840);
or U12016 (N_12016,N_10622,N_10763);
xor U12017 (N_12017,N_11729,N_10634);
or U12018 (N_12018,N_10732,N_10641);
nand U12019 (N_12019,N_10939,N_10881);
nand U12020 (N_12020,N_11900,N_10955);
nor U12021 (N_12021,N_10545,N_11173);
xor U12022 (N_12022,N_10675,N_11876);
nor U12023 (N_12023,N_11688,N_10919);
nor U12024 (N_12024,N_10554,N_10723);
xnor U12025 (N_12025,N_11882,N_10905);
nand U12026 (N_12026,N_11819,N_11907);
and U12027 (N_12027,N_11628,N_10618);
nand U12028 (N_12028,N_11460,N_10531);
and U12029 (N_12029,N_11004,N_11856);
nor U12030 (N_12030,N_11917,N_11775);
nand U12031 (N_12031,N_10954,N_11493);
and U12032 (N_12032,N_11923,N_11753);
xor U12033 (N_12033,N_11048,N_10528);
or U12034 (N_12034,N_11727,N_11802);
nor U12035 (N_12035,N_10661,N_11494);
and U12036 (N_12036,N_10606,N_10706);
nor U12037 (N_12037,N_11334,N_11615);
nand U12038 (N_12038,N_11060,N_11827);
nand U12039 (N_12039,N_11858,N_11218);
and U12040 (N_12040,N_11877,N_11152);
nand U12041 (N_12041,N_10530,N_11777);
or U12042 (N_12042,N_10875,N_11382);
or U12043 (N_12043,N_10988,N_11549);
xor U12044 (N_12044,N_11742,N_10681);
xor U12045 (N_12045,N_11353,N_10688);
nand U12046 (N_12046,N_11146,N_10886);
nor U12047 (N_12047,N_11464,N_10754);
or U12048 (N_12048,N_11491,N_11141);
xor U12049 (N_12049,N_10724,N_11295);
and U12050 (N_12050,N_10877,N_11706);
nor U12051 (N_12051,N_11869,N_10624);
nand U12052 (N_12052,N_11725,N_11662);
xor U12053 (N_12053,N_11367,N_10518);
nor U12054 (N_12054,N_11360,N_11849);
nand U12055 (N_12055,N_10802,N_10583);
nor U12056 (N_12056,N_10854,N_11838);
and U12057 (N_12057,N_11245,N_10811);
or U12058 (N_12058,N_11304,N_11941);
xor U12059 (N_12059,N_11342,N_11357);
xnor U12060 (N_12060,N_11904,N_11945);
xnor U12061 (N_12061,N_11145,N_10534);
nor U12062 (N_12062,N_11235,N_11219);
or U12063 (N_12063,N_11358,N_11373);
nor U12064 (N_12064,N_11880,N_11537);
xor U12065 (N_12065,N_11347,N_11162);
nand U12066 (N_12066,N_11398,N_11596);
nor U12067 (N_12067,N_11558,N_11392);
or U12068 (N_12068,N_11938,N_10985);
xnor U12069 (N_12069,N_10682,N_10717);
and U12070 (N_12070,N_11581,N_11899);
or U12071 (N_12071,N_11593,N_11181);
and U12072 (N_12072,N_11671,N_11437);
or U12073 (N_12073,N_10797,N_11773);
or U12074 (N_12074,N_11463,N_11477);
nand U12075 (N_12075,N_11469,N_11484);
and U12076 (N_12076,N_11974,N_10937);
or U12077 (N_12077,N_11552,N_11170);
nand U12078 (N_12078,N_11260,N_11489);
and U12079 (N_12079,N_10762,N_10798);
and U12080 (N_12080,N_11247,N_11632);
nor U12081 (N_12081,N_11485,N_10698);
xnor U12082 (N_12082,N_11750,N_11860);
and U12083 (N_12083,N_11175,N_11831);
nand U12084 (N_12084,N_10836,N_11378);
nor U12085 (N_12085,N_11798,N_10861);
or U12086 (N_12086,N_10805,N_10747);
xor U12087 (N_12087,N_11804,N_10761);
nor U12088 (N_12088,N_11545,N_11765);
nand U12089 (N_12089,N_11589,N_10753);
or U12090 (N_12090,N_10856,N_10775);
nor U12091 (N_12091,N_11099,N_11441);
nand U12092 (N_12092,N_11768,N_10578);
nor U12093 (N_12093,N_11957,N_11169);
and U12094 (N_12094,N_11063,N_10702);
xor U12095 (N_12095,N_11616,N_11417);
or U12096 (N_12096,N_11517,N_10832);
or U12097 (N_12097,N_11698,N_11403);
xnor U12098 (N_12098,N_11713,N_11034);
nor U12099 (N_12099,N_10859,N_11291);
nand U12100 (N_12100,N_10893,N_11212);
or U12101 (N_12101,N_11799,N_11525);
nand U12102 (N_12102,N_11959,N_11745);
nor U12103 (N_12103,N_10815,N_11423);
xnor U12104 (N_12104,N_11801,N_11220);
or U12105 (N_12105,N_10827,N_11842);
xnor U12106 (N_12106,N_11603,N_11609);
nand U12107 (N_12107,N_10695,N_11668);
and U12108 (N_12108,N_11861,N_11316);
nor U12109 (N_12109,N_11955,N_10599);
nor U12110 (N_12110,N_11190,N_11227);
nor U12111 (N_12111,N_10816,N_11009);
or U12112 (N_12112,N_11231,N_11649);
nand U12113 (N_12113,N_11530,N_11355);
or U12114 (N_12114,N_11859,N_10858);
nand U12115 (N_12115,N_11881,N_10851);
or U12116 (N_12116,N_10609,N_11285);
xnor U12117 (N_12117,N_11514,N_10971);
xor U12118 (N_12118,N_11018,N_11998);
nand U12119 (N_12119,N_11487,N_11035);
nor U12120 (N_12120,N_10607,N_11943);
nand U12121 (N_12121,N_10700,N_11021);
nand U12122 (N_12122,N_11951,N_10619);
nor U12123 (N_12123,N_10772,N_11721);
nor U12124 (N_12124,N_11416,N_10729);
nand U12125 (N_12125,N_10970,N_11215);
nand U12126 (N_12126,N_11259,N_10842);
nand U12127 (N_12127,N_11813,N_11226);
and U12128 (N_12128,N_10617,N_11174);
nor U12129 (N_12129,N_11273,N_11396);
xor U12130 (N_12130,N_10941,N_10591);
nand U12131 (N_12131,N_10625,N_11092);
nand U12132 (N_12132,N_11158,N_11014);
nor U12133 (N_12133,N_11663,N_11695);
nand U12134 (N_12134,N_11161,N_11409);
nor U12135 (N_12135,N_11027,N_10968);
nand U12136 (N_12136,N_11025,N_11254);
nand U12137 (N_12137,N_11049,N_10899);
nor U12138 (N_12138,N_10976,N_11851);
xnor U12139 (N_12139,N_10929,N_11139);
nor U12140 (N_12140,N_11167,N_11949);
nor U12141 (N_12141,N_11012,N_11751);
and U12142 (N_12142,N_11772,N_10902);
or U12143 (N_12143,N_10814,N_10913);
and U12144 (N_12144,N_10785,N_11731);
xnor U12145 (N_12145,N_10776,N_10669);
and U12146 (N_12146,N_11144,N_11846);
nor U12147 (N_12147,N_10662,N_11930);
or U12148 (N_12148,N_11269,N_10803);
nand U12149 (N_12149,N_11108,N_10793);
or U12150 (N_12150,N_11843,N_10848);
or U12151 (N_12151,N_10882,N_11529);
xnor U12152 (N_12152,N_11635,N_10909);
nor U12153 (N_12153,N_11915,N_11443);
xor U12154 (N_12154,N_10903,N_11116);
xor U12155 (N_12155,N_11771,N_10915);
xnor U12156 (N_12156,N_11780,N_11818);
nand U12157 (N_12157,N_11527,N_11913);
nand U12158 (N_12158,N_10787,N_11272);
xor U12159 (N_12159,N_10835,N_11870);
or U12160 (N_12160,N_10991,N_10818);
xor U12161 (N_12161,N_10580,N_11978);
and U12162 (N_12162,N_11189,N_10807);
xnor U12163 (N_12163,N_10849,N_11246);
nor U12164 (N_12164,N_11997,N_11733);
nor U12165 (N_12165,N_11248,N_10581);
nand U12166 (N_12166,N_10998,N_11944);
nor U12167 (N_12167,N_11637,N_11720);
nor U12168 (N_12168,N_11322,N_11408);
nor U12169 (N_12169,N_11950,N_10812);
nor U12170 (N_12170,N_11594,N_11202);
nand U12171 (N_12171,N_11420,N_11135);
or U12172 (N_12172,N_11061,N_11587);
nand U12173 (N_12173,N_10889,N_11574);
or U12174 (N_12174,N_10918,N_11440);
xnor U12175 (N_12175,N_10795,N_11987);
xnor U12176 (N_12176,N_10890,N_10749);
and U12177 (N_12177,N_10796,N_11762);
xor U12178 (N_12178,N_11747,N_11261);
or U12179 (N_12179,N_11712,N_11125);
and U12180 (N_12180,N_11318,N_11372);
nand U12181 (N_12181,N_10600,N_11433);
or U12182 (N_12182,N_10574,N_10713);
xnor U12183 (N_12183,N_11826,N_10718);
or U12184 (N_12184,N_11496,N_11257);
or U12185 (N_12185,N_11510,N_11891);
or U12186 (N_12186,N_11263,N_11107);
nand U12187 (N_12187,N_10895,N_11154);
or U12188 (N_12188,N_11787,N_11091);
xor U12189 (N_12189,N_11076,N_10509);
nand U12190 (N_12190,N_10642,N_11293);
or U12191 (N_12191,N_11149,N_11002);
and U12192 (N_12192,N_11728,N_11976);
nand U12193 (N_12193,N_11981,N_11391);
and U12194 (N_12194,N_10646,N_10694);
nor U12195 (N_12195,N_11965,N_11036);
and U12196 (N_12196,N_11647,N_11216);
nand U12197 (N_12197,N_10961,N_10917);
xor U12198 (N_12198,N_10879,N_11458);
nor U12199 (N_12199,N_10673,N_11228);
and U12200 (N_12200,N_11590,N_11873);
or U12201 (N_12201,N_11462,N_10935);
and U12202 (N_12202,N_10594,N_11112);
nor U12203 (N_12203,N_11362,N_10556);
or U12204 (N_12204,N_10623,N_11449);
xor U12205 (N_12205,N_11077,N_10683);
xor U12206 (N_12206,N_11363,N_11599);
and U12207 (N_12207,N_10628,N_11607);
nand U12208 (N_12208,N_11694,N_11124);
and U12209 (N_12209,N_11121,N_11068);
and U12210 (N_12210,N_10632,N_10711);
nand U12211 (N_12211,N_11303,N_11333);
or U12212 (N_12212,N_11833,N_10519);
nand U12213 (N_12213,N_11536,N_11364);
nor U12214 (N_12214,N_10779,N_11521);
and U12215 (N_12215,N_10928,N_10564);
nand U12216 (N_12216,N_11716,N_11889);
nand U12217 (N_12217,N_11914,N_11884);
xor U12218 (N_12218,N_10862,N_11715);
xnor U12219 (N_12219,N_11911,N_11905);
or U12220 (N_12220,N_11774,N_11701);
nor U12221 (N_12221,N_11645,N_11103);
nand U12222 (N_12222,N_11136,N_11090);
or U12223 (N_12223,N_10957,N_10789);
nor U12224 (N_12224,N_10728,N_11282);
or U12225 (N_12225,N_11138,N_10679);
xnor U12226 (N_12226,N_11678,N_11388);
or U12227 (N_12227,N_11868,N_11602);
or U12228 (N_12228,N_11932,N_11758);
or U12229 (N_12229,N_11126,N_11608);
and U12230 (N_12230,N_11646,N_11467);
and U12231 (N_12231,N_11019,N_11970);
or U12232 (N_12232,N_11283,N_11792);
and U12233 (N_12233,N_11642,N_11005);
xnor U12234 (N_12234,N_11520,N_11683);
or U12235 (N_12235,N_11199,N_10799);
nand U12236 (N_12236,N_11200,N_11194);
xor U12237 (N_12237,N_10967,N_10542);
and U12238 (N_12238,N_11150,N_11447);
or U12239 (N_12239,N_10739,N_11084);
and U12240 (N_12240,N_10503,N_11759);
or U12241 (N_12241,N_10500,N_11500);
nand U12242 (N_12242,N_10767,N_11814);
or U12243 (N_12243,N_11737,N_11007);
xnor U12244 (N_12244,N_11795,N_10965);
or U12245 (N_12245,N_10876,N_11515);
nand U12246 (N_12246,N_11708,N_10592);
nor U12247 (N_12247,N_10744,N_10565);
nand U12248 (N_12248,N_10691,N_11253);
nor U12249 (N_12249,N_11255,N_11381);
nor U12250 (N_12250,N_10950,N_11101);
and U12251 (N_12251,N_10819,N_10605);
or U12252 (N_12252,N_11058,N_10601);
and U12253 (N_12253,N_11390,N_11785);
and U12254 (N_12254,N_11625,N_10746);
nand U12255 (N_12255,N_11769,N_11898);
and U12256 (N_12256,N_11687,N_11102);
nand U12257 (N_12257,N_11298,N_11428);
xor U12258 (N_12258,N_11829,N_10692);
xor U12259 (N_12259,N_11523,N_10900);
and U12260 (N_12260,N_10778,N_11455);
or U12261 (N_12261,N_11832,N_10994);
or U12262 (N_12262,N_11677,N_10508);
nand U12263 (N_12263,N_10515,N_10852);
or U12264 (N_12264,N_10584,N_10921);
nand U12265 (N_12265,N_11928,N_11309);
xnor U12266 (N_12266,N_10635,N_10813);
nand U12267 (N_12267,N_10999,N_11993);
xor U12268 (N_12268,N_11643,N_11969);
or U12269 (N_12269,N_11601,N_10615);
nor U12270 (N_12270,N_11452,N_11177);
nand U12271 (N_12271,N_10510,N_10696);
or U12272 (N_12272,N_11296,N_11134);
or U12273 (N_12273,N_10888,N_10883);
and U12274 (N_12274,N_11985,N_11797);
nor U12275 (N_12275,N_11043,N_10532);
xor U12276 (N_12276,N_11271,N_11811);
nand U12277 (N_12277,N_11486,N_10620);
nor U12278 (N_12278,N_11623,N_10552);
xnor U12279 (N_12279,N_11760,N_10655);
nor U12280 (N_12280,N_11055,N_11057);
nand U12281 (N_12281,N_11680,N_11684);
nor U12282 (N_12282,N_11359,N_11280);
nand U12283 (N_12283,N_11539,N_10948);
and U12284 (N_12284,N_11654,N_10541);
or U12285 (N_12285,N_10756,N_10666);
nor U12286 (N_12286,N_11156,N_10667);
and U12287 (N_12287,N_11948,N_10631);
nor U12288 (N_12288,N_10514,N_11749);
or U12289 (N_12289,N_11561,N_11805);
or U12290 (N_12290,N_10588,N_10891);
or U12291 (N_12291,N_11661,N_11142);
and U12292 (N_12292,N_11165,N_10658);
nor U12293 (N_12293,N_11041,N_11187);
nor U12294 (N_12294,N_10603,N_10613);
or U12295 (N_12295,N_11502,N_11120);
xnor U12296 (N_12296,N_10575,N_11685);
xnor U12297 (N_12297,N_11188,N_10708);
or U12298 (N_12298,N_11383,N_11559);
nand U12299 (N_12299,N_11918,N_11746);
nand U12300 (N_12300,N_11171,N_11328);
nor U12301 (N_12301,N_11550,N_11032);
xor U12302 (N_12302,N_10627,N_10652);
nor U12303 (N_12303,N_10977,N_10922);
and U12304 (N_12304,N_11104,N_11979);
or U12305 (N_12305,N_11582,N_11300);
xnor U12306 (N_12306,N_10558,N_10853);
or U12307 (N_12307,N_11386,N_11453);
xnor U12308 (N_12308,N_10586,N_11553);
or U12309 (N_12309,N_11405,N_11779);
and U12310 (N_12310,N_11650,N_11130);
nand U12311 (N_12311,N_11479,N_10934);
or U12312 (N_12312,N_10726,N_11563);
and U12313 (N_12313,N_11585,N_10943);
xor U12314 (N_12314,N_11557,N_11538);
or U12315 (N_12315,N_11348,N_10551);
or U12316 (N_12316,N_11268,N_11906);
nor U12317 (N_12317,N_10958,N_10645);
nor U12318 (N_12318,N_11853,N_11903);
xnor U12319 (N_12319,N_10540,N_11376);
and U12320 (N_12320,N_11225,N_11474);
and U12321 (N_12321,N_11001,N_11690);
and U12322 (N_12322,N_10522,N_10822);
or U12323 (N_12323,N_11696,N_10649);
or U12324 (N_12324,N_11532,N_11224);
and U12325 (N_12325,N_11852,N_11666);
nor U12326 (N_12326,N_11665,N_10898);
xor U12327 (N_12327,N_11597,N_11109);
and U12328 (N_12328,N_10806,N_10533);
nand U12329 (N_12329,N_10986,N_11310);
and U12330 (N_12330,N_11823,N_10878);
nand U12331 (N_12331,N_11122,N_10869);
nor U12332 (N_12332,N_11178,N_11501);
and U12333 (N_12333,N_11572,N_11800);
or U12334 (N_12334,N_11864,N_11707);
nor U12335 (N_12335,N_11735,N_10731);
and U12336 (N_12336,N_11681,N_11085);
or U12337 (N_12337,N_11211,N_11312);
and U12338 (N_12338,N_11887,N_11972);
and U12339 (N_12339,N_11718,N_10982);
nand U12340 (N_12340,N_10926,N_11281);
nand U12341 (N_12341,N_10525,N_11850);
and U12342 (N_12342,N_11975,N_10945);
nor U12343 (N_12343,N_10870,N_10569);
nand U12344 (N_12344,N_10536,N_11472);
nand U12345 (N_12345,N_11789,N_10524);
or U12346 (N_12346,N_10927,N_11541);
xnor U12347 (N_12347,N_11468,N_11237);
xor U12348 (N_12348,N_11030,N_11208);
and U12349 (N_12349,N_10783,N_11096);
or U12350 (N_12350,N_11825,N_11262);
nor U12351 (N_12351,N_10582,N_10727);
and U12352 (N_12352,N_10944,N_10765);
nand U12353 (N_12353,N_10593,N_11986);
xnor U12354 (N_12354,N_11432,N_11548);
or U12355 (N_12355,N_11886,N_11193);
and U12356 (N_12356,N_10549,N_11321);
and U12357 (N_12357,N_10949,N_11505);
nor U12358 (N_12358,N_10940,N_11809);
nand U12359 (N_12359,N_11509,N_11323);
and U12360 (N_12360,N_10576,N_11822);
nand U12361 (N_12361,N_11697,N_11562);
nor U12362 (N_12362,N_11180,N_11153);
xnor U12363 (N_12363,N_11111,N_10804);
and U12364 (N_12364,N_11693,N_11929);
xnor U12365 (N_12365,N_11054,N_11198);
or U12366 (N_12366,N_10611,N_11042);
and U12367 (N_12367,N_10907,N_11613);
nand U12368 (N_12368,N_11098,N_10737);
xnor U12369 (N_12369,N_11223,N_11482);
or U12370 (N_12370,N_10942,N_11302);
nand U12371 (N_12371,N_10995,N_11573);
nor U12372 (N_12372,N_10637,N_11504);
and U12373 (N_12373,N_10665,N_11250);
and U12374 (N_12374,N_11791,N_10709);
or U12375 (N_12375,N_10897,N_10506);
nor U12376 (N_12376,N_11511,N_11412);
and U12377 (N_12377,N_11147,N_11406);
nand U12378 (N_12378,N_10626,N_11528);
xor U12379 (N_12379,N_11385,N_11963);
nor U12380 (N_12380,N_11794,N_10686);
nor U12381 (N_12381,N_11326,N_11577);
nand U12382 (N_12382,N_11470,N_11839);
nor U12383 (N_12383,N_11072,N_11411);
or U12384 (N_12384,N_11513,N_10938);
or U12385 (N_12385,N_11897,N_11937);
nand U12386 (N_12386,N_11531,N_11786);
nor U12387 (N_12387,N_11011,N_11000);
xnor U12388 (N_12388,N_10660,N_11422);
xor U12389 (N_12389,N_11790,N_11079);
xnor U12390 (N_12390,N_10884,N_10630);
and U12391 (N_12391,N_11784,N_11535);
or U12392 (N_12392,N_11570,N_11658);
nor U12393 (N_12393,N_10932,N_10638);
or U12394 (N_12394,N_11893,N_11875);
xnor U12395 (N_12395,N_10933,N_11892);
nor U12396 (N_12396,N_11370,N_11543);
nor U12397 (N_12397,N_11920,N_11029);
xor U12398 (N_12398,N_11380,N_10959);
or U12399 (N_12399,N_11705,N_11454);
and U12400 (N_12400,N_11604,N_10820);
nand U12401 (N_12401,N_11183,N_11127);
nor U12402 (N_12402,N_11922,N_11895);
xor U12403 (N_12403,N_11052,N_11620);
xor U12404 (N_12404,N_11350,N_11266);
or U12405 (N_12405,N_11744,N_11936);
nor U12406 (N_12406,N_10864,N_10894);
nand U12407 (N_12407,N_10790,N_10719);
or U12408 (N_12408,N_11429,N_11475);
nand U12409 (N_12409,N_10643,N_11995);
xnor U12410 (N_12410,N_10781,N_10755);
or U12411 (N_12411,N_11766,N_11095);
xnor U12412 (N_12412,N_11377,N_11080);
nand U12413 (N_12413,N_11075,N_11736);
nand U12414 (N_12414,N_10505,N_11176);
and U12415 (N_12415,N_10735,N_10771);
and U12416 (N_12416,N_11512,N_10561);
nand U12417 (N_12417,N_11393,N_11518);
nor U12418 (N_12418,N_11990,N_11954);
xnor U12419 (N_12419,N_11939,N_10750);
nand U12420 (N_12420,N_10676,N_11448);
and U12421 (N_12421,N_11952,N_11544);
nor U12422 (N_12422,N_10993,N_11820);
xor U12423 (N_12423,N_11461,N_10648);
nand U12424 (N_12424,N_11503,N_11065);
nor U12425 (N_12425,N_11916,N_10504);
xor U12426 (N_12426,N_11748,N_10748);
or U12427 (N_12427,N_10989,N_11947);
and U12428 (N_12428,N_11516,N_11934);
and U12429 (N_12429,N_11421,N_11793);
and U12430 (N_12430,N_11738,N_11401);
nand U12431 (N_12431,N_11431,N_10579);
and U12432 (N_12432,N_10722,N_11857);
or U12433 (N_12433,N_11931,N_11651);
nor U12434 (N_12434,N_10866,N_11240);
or U12435 (N_12435,N_10684,N_11093);
nor U12436 (N_12436,N_10828,N_11094);
and U12437 (N_12437,N_10837,N_11059);
or U12438 (N_12438,N_11368,N_11366);
xor U12439 (N_12439,N_11591,N_11466);
or U12440 (N_12440,N_11221,N_11151);
and U12441 (N_12441,N_10595,N_10912);
nand U12442 (N_12442,N_11569,N_11137);
nor U12443 (N_12443,N_11933,N_10992);
xnor U12444 (N_12444,N_10539,N_10910);
nand U12445 (N_12445,N_10960,N_11546);
and U12446 (N_12446,N_11534,N_11723);
and U12447 (N_12447,N_11692,N_11834);
or U12448 (N_12448,N_11547,N_11926);
or U12449 (N_12449,N_11424,N_11209);
nand U12450 (N_12450,N_11586,N_10701);
or U12451 (N_12451,N_11251,N_11560);
or U12452 (N_12452,N_11106,N_10996);
xnor U12453 (N_12453,N_11767,N_11069);
xor U12454 (N_12454,N_11324,N_11821);
or U12455 (N_12455,N_11415,N_11003);
nor U12456 (N_12456,N_11726,N_10687);
xor U12457 (N_12457,N_10952,N_11172);
nand U12458 (N_12458,N_10981,N_10857);
nand U12459 (N_12459,N_11022,N_11611);
or U12460 (N_12460,N_11294,N_11132);
xnor U12461 (N_12461,N_10768,N_11781);
and U12462 (N_12462,N_10734,N_10656);
nor U12463 (N_12463,N_10721,N_11710);
xnor U12464 (N_12464,N_11855,N_10930);
xnor U12465 (N_12465,N_10537,N_11100);
and U12466 (N_12466,N_11730,N_11439);
and U12467 (N_12467,N_11624,N_11430);
nand U12468 (N_12468,N_11155,N_11279);
nor U12469 (N_12469,N_11812,N_11444);
or U12470 (N_12470,N_11682,N_10571);
or U12471 (N_12471,N_11711,N_10757);
or U12472 (N_12472,N_11404,N_11921);
nor U12473 (N_12473,N_10526,N_11402);
nor U12474 (N_12474,N_11184,N_11305);
nand U12475 (N_12475,N_11568,N_11297);
nand U12476 (N_12476,N_11689,N_11579);
nor U12477 (N_12477,N_11277,N_11583);
xnor U12478 (N_12478,N_11770,N_11764);
xnor U12479 (N_12479,N_11714,N_11824);
or U12480 (N_12480,N_10826,N_11669);
xor U12481 (N_12481,N_10887,N_11992);
and U12482 (N_12482,N_11967,N_11047);
or U12483 (N_12483,N_11830,N_10544);
nand U12484 (N_12484,N_10801,N_11196);
and U12485 (N_12485,N_11473,N_11709);
nor U12486 (N_12486,N_11796,N_10604);
nor U12487 (N_12487,N_11033,N_11739);
and U12488 (N_12488,N_11044,N_11704);
or U12489 (N_12489,N_11761,N_11045);
nor U12490 (N_12490,N_11163,N_10527);
and U12491 (N_12491,N_11006,N_11964);
nor U12492 (N_12492,N_11195,N_11354);
or U12493 (N_12493,N_11081,N_11234);
or U12494 (N_12494,N_10653,N_11131);
or U12495 (N_12495,N_11427,N_11580);
or U12496 (N_12496,N_11129,N_10920);
and U12497 (N_12497,N_10543,N_10740);
nand U12498 (N_12498,N_10831,N_10969);
xnor U12499 (N_12499,N_10834,N_11284);
or U12500 (N_12500,N_10547,N_11204);
nand U12501 (N_12501,N_11352,N_11639);
nor U12502 (N_12502,N_11017,N_11308);
nand U12503 (N_12503,N_11407,N_11389);
and U12504 (N_12504,N_10784,N_10885);
or U12505 (N_12505,N_11595,N_11507);
or U12506 (N_12506,N_10825,N_10978);
nand U12507 (N_12507,N_11243,N_11630);
and U12508 (N_12508,N_10659,N_11841);
and U12509 (N_12509,N_10738,N_11909);
nor U12510 (N_12510,N_11148,N_11286);
xor U12511 (N_12511,N_11674,N_11087);
and U12512 (N_12512,N_10874,N_11425);
xnor U12513 (N_12513,N_11925,N_10697);
or U12514 (N_12514,N_11741,N_11275);
xnor U12515 (N_12515,N_11940,N_10689);
xnor U12516 (N_12516,N_11301,N_11332);
nor U12517 (N_12517,N_10529,N_11757);
xnor U12518 (N_12518,N_11657,N_11867);
nand U12519 (N_12519,N_10664,N_11871);
and U12520 (N_12520,N_11566,N_11258);
or U12521 (N_12521,N_11341,N_11369);
nor U12522 (N_12522,N_10873,N_10990);
and U12523 (N_12523,N_10788,N_10559);
xor U12524 (N_12524,N_10577,N_11166);
and U12525 (N_12525,N_10904,N_11242);
xnor U12526 (N_12526,N_11435,N_10855);
nand U12527 (N_12527,N_10838,N_11346);
or U12528 (N_12528,N_11644,N_10868);
or U12529 (N_12529,N_10521,N_11481);
or U12530 (N_12530,N_10629,N_10956);
nor U12531 (N_12531,N_11016,N_10865);
nand U12532 (N_12532,N_10716,N_10680);
nor U12533 (N_12533,N_10983,N_11276);
or U12534 (N_12534,N_10538,N_10850);
xor U12535 (N_12535,N_11946,N_11743);
nor U12536 (N_12536,N_10774,N_10513);
nand U12537 (N_12537,N_11588,N_11935);
and U12538 (N_12538,N_11629,N_10589);
or U12539 (N_12539,N_11319,N_10690);
nand U12540 (N_12540,N_10966,N_10548);
nand U12541 (N_12541,N_10636,N_11533);
and U12542 (N_12542,N_11140,N_10590);
xor U12543 (N_12543,N_10596,N_11434);
nor U12544 (N_12544,N_11256,N_11499);
xnor U12545 (N_12545,N_11008,N_10800);
nand U12546 (N_12546,N_11306,N_10560);
nand U12547 (N_12547,N_10770,N_11872);
or U12548 (N_12548,N_10936,N_11056);
xnor U12549 (N_12549,N_11717,N_10860);
nor U12550 (N_12550,N_11290,N_11083);
xor U12551 (N_12551,N_11110,N_10707);
nand U12552 (N_12552,N_11664,N_11213);
and U12553 (N_12553,N_11636,N_11648);
and U12554 (N_12554,N_11700,N_10911);
nor U12555 (N_12555,N_11384,N_11410);
xor U12556 (N_12556,N_10984,N_10657);
and U12557 (N_12557,N_10502,N_10616);
and U12558 (N_12558,N_11519,N_11752);
and U12559 (N_12559,N_11763,N_10880);
and U12560 (N_12560,N_10557,N_11483);
nand U12561 (N_12561,N_11854,N_11719);
nand U12562 (N_12562,N_11901,N_10963);
xor U12563 (N_12563,N_10871,N_10845);
and U12564 (N_12564,N_10760,N_11862);
nor U12565 (N_12565,N_11732,N_11605);
or U12566 (N_12566,N_11325,N_10745);
and U12567 (N_12567,N_11542,N_11331);
and U12568 (N_12568,N_11039,N_11564);
xor U12569 (N_12569,N_11612,N_11672);
nand U12570 (N_12570,N_11010,N_11064);
nor U12571 (N_12571,N_10997,N_11983);
nor U12572 (N_12572,N_11400,N_10567);
xnor U12573 (N_12573,N_11971,N_10896);
xor U12574 (N_12574,N_11927,N_10844);
xor U12575 (N_12575,N_11115,N_10563);
and U12576 (N_12576,N_11592,N_11641);
and U12577 (N_12577,N_11238,N_11186);
nand U12578 (N_12578,N_11088,N_11264);
nand U12579 (N_12579,N_11633,N_11980);
xnor U12580 (N_12580,N_11686,N_11201);
nand U12581 (N_12581,N_11179,N_11089);
and U12582 (N_12582,N_11879,N_11236);
or U12583 (N_12583,N_11336,N_11046);
nor U12584 (N_12584,N_10725,N_10925);
nand U12585 (N_12585,N_10973,N_10736);
or U12586 (N_12586,N_11724,N_11912);
nor U12587 (N_12587,N_11097,N_10979);
nand U12588 (N_12588,N_11270,N_11958);
xor U12589 (N_12589,N_11584,N_11627);
xor U12590 (N_12590,N_11863,N_11621);
and U12591 (N_12591,N_11526,N_10863);
xor U12592 (N_12592,N_11902,N_11292);
nand U12593 (N_12593,N_11977,N_11488);
and U12594 (N_12594,N_10550,N_10846);
or U12595 (N_12595,N_11026,N_11419);
nor U12596 (N_12596,N_11205,N_11631);
xnor U12597 (N_12597,N_10791,N_10710);
nor U12598 (N_12598,N_10650,N_11185);
and U12599 (N_12599,N_11960,N_11418);
or U12600 (N_12600,N_11249,N_11492);
nand U12601 (N_12601,N_10633,N_11614);
or U12602 (N_12602,N_10535,N_11314);
nand U12603 (N_12603,N_11442,N_10703);
and U12604 (N_12604,N_10810,N_11540);
xor U12605 (N_12605,N_10947,N_11086);
nor U12606 (N_12606,N_11015,N_11778);
and U12607 (N_12607,N_11640,N_11320);
or U12608 (N_12608,N_11807,N_11387);
nor U12609 (N_12609,N_11622,N_10867);
nor U12610 (N_12610,N_10570,N_10741);
nand U12611 (N_12611,N_10743,N_11289);
xor U12612 (N_12612,N_10555,N_11756);
nor U12613 (N_12613,N_10672,N_10674);
nor U12614 (N_12614,N_11066,N_11274);
and U12615 (N_12615,N_11217,N_11699);
or U12616 (N_12616,N_11233,N_11506);
or U12617 (N_12617,N_11267,N_11119);
nand U12618 (N_12618,N_11703,N_11626);
nor U12619 (N_12619,N_10668,N_11885);
xor U12620 (N_12620,N_11203,N_11299);
or U12621 (N_12621,N_11844,N_10553);
nand U12622 (N_12622,N_10712,N_11335);
nand U12623 (N_12623,N_11837,N_11555);
and U12624 (N_12624,N_11210,N_11078);
or U12625 (N_12625,N_11062,N_11013);
xor U12626 (N_12626,N_10516,N_11040);
nand U12627 (N_12627,N_11675,N_11252);
or U12628 (N_12628,N_11315,N_10780);
nand U12629 (N_12629,N_11456,N_11808);
nand U12630 (N_12630,N_11910,N_11828);
nor U12631 (N_12631,N_11192,N_11356);
nor U12632 (N_12632,N_11446,N_11618);
or U12633 (N_12633,N_11840,N_11123);
and U12634 (N_12634,N_11476,N_10808);
xnor U12635 (N_12635,N_11480,N_10794);
and U12636 (N_12636,N_11498,N_10705);
or U12637 (N_12637,N_11754,N_11339);
nand U12638 (N_12638,N_11037,N_11806);
or U12639 (N_12639,N_11679,N_11845);
and U12640 (N_12640,N_11067,N_11445);
or U12641 (N_12641,N_11722,N_10769);
or U12642 (N_12642,N_11330,N_11239);
xor U12643 (N_12643,N_11702,N_11288);
nor U12644 (N_12644,N_11020,N_11031);
or U12645 (N_12645,N_10568,N_11874);
and U12646 (N_12646,N_10663,N_11788);
xnor U12647 (N_12647,N_11374,N_10597);
nand U12648 (N_12648,N_11450,N_11113);
or U12649 (N_12649,N_11994,N_11214);
and U12650 (N_12650,N_11554,N_11890);
or U12651 (N_12651,N_10829,N_11556);
xnor U12652 (N_12652,N_11810,N_11164);
nor U12653 (N_12653,N_11338,N_11634);
nand U12654 (N_12654,N_11803,N_11024);
and U12655 (N_12655,N_10511,N_10699);
xor U12656 (N_12656,N_11071,N_11782);
nor U12657 (N_12657,N_11478,N_11465);
and U12658 (N_12658,N_10715,N_10610);
nand U12659 (N_12659,N_10786,N_11365);
xnor U12660 (N_12660,N_10654,N_10677);
xnor U12661 (N_12661,N_11157,N_11866);
nand U12662 (N_12662,N_10892,N_10720);
nor U12663 (N_12663,N_11229,N_11413);
and U12664 (N_12664,N_11691,N_11655);
or U12665 (N_12665,N_11956,N_11241);
and U12666 (N_12666,N_11606,N_11962);
nor U12667 (N_12667,N_10612,N_11344);
and U12668 (N_12668,N_11053,N_11740);
nand U12669 (N_12669,N_11232,N_10562);
and U12670 (N_12670,N_11652,N_10974);
xor U12671 (N_12671,N_11197,N_10501);
and U12672 (N_12672,N_11776,N_10507);
or U12673 (N_12673,N_10792,N_11961);
xor U12674 (N_12674,N_11617,N_10742);
xor U12675 (N_12675,N_10647,N_11371);
or U12676 (N_12676,N_10704,N_11953);
xor U12677 (N_12677,N_10758,N_11471);
xnor U12678 (N_12678,N_11143,N_11734);
and U12679 (N_12679,N_10841,N_10924);
xnor U12680 (N_12680,N_11619,N_11313);
xor U12681 (N_12681,N_11307,N_11497);
xor U12682 (N_12682,N_10517,N_11311);
and U12683 (N_12683,N_10809,N_10773);
and U12684 (N_12684,N_10766,N_10598);
or U12685 (N_12685,N_11375,N_11395);
nor U12686 (N_12686,N_10608,N_11551);
or U12687 (N_12687,N_11576,N_10821);
xnor U12688 (N_12688,N_11230,N_11327);
nor U12689 (N_12689,N_11815,N_10639);
or U12690 (N_12690,N_10759,N_11989);
or U12691 (N_12691,N_10962,N_11073);
nor U12692 (N_12692,N_11117,N_11848);
or U12693 (N_12693,N_11160,N_11343);
nor U12694 (N_12694,N_11459,N_11414);
xor U12695 (N_12695,N_11023,N_10730);
xor U12696 (N_12696,N_11379,N_11865);
xor U12697 (N_12697,N_11399,N_11351);
or U12698 (N_12698,N_10602,N_10546);
xnor U12699 (N_12699,N_11438,N_11361);
xor U12700 (N_12700,N_11991,N_10685);
nor U12701 (N_12701,N_11847,N_11999);
and U12702 (N_12702,N_10953,N_11524);
xnor U12703 (N_12703,N_10824,N_11638);
or U12704 (N_12704,N_10964,N_11114);
nand U12705 (N_12705,N_11836,N_11755);
or U12706 (N_12706,N_10566,N_11942);
or U12707 (N_12707,N_11265,N_11495);
nand U12708 (N_12708,N_10585,N_10573);
nor U12709 (N_12709,N_11919,N_10520);
nor U12710 (N_12710,N_11610,N_11966);
and U12711 (N_12711,N_10906,N_11924);
xor U12712 (N_12712,N_11451,N_11653);
and U12713 (N_12713,N_10847,N_11133);
and U12714 (N_12714,N_10843,N_11598);
nand U12715 (N_12715,N_11345,N_10621);
nor U12716 (N_12716,N_10587,N_10572);
or U12717 (N_12717,N_11896,N_10714);
or U12718 (N_12718,N_10640,N_11050);
nand U12719 (N_12719,N_11397,N_10523);
and U12720 (N_12720,N_11888,N_10980);
xnor U12721 (N_12721,N_11908,N_10782);
and U12722 (N_12722,N_11207,N_10777);
and U12723 (N_12723,N_10614,N_11982);
or U12724 (N_12724,N_11571,N_10923);
and U12725 (N_12725,N_11835,N_11222);
or U12726 (N_12726,N_11349,N_10872);
nand U12727 (N_12727,N_11105,N_11816);
nand U12728 (N_12728,N_11984,N_11051);
nand U12729 (N_12729,N_10671,N_11028);
xnor U12730 (N_12730,N_11656,N_11676);
nand U12731 (N_12731,N_11082,N_11673);
nand U12732 (N_12732,N_11337,N_11660);
xor U12733 (N_12733,N_10987,N_11168);
xor U12734 (N_12734,N_11996,N_10901);
or U12735 (N_12735,N_10512,N_11783);
and U12736 (N_12736,N_11278,N_11182);
and U12737 (N_12737,N_10916,N_11817);
nor U12738 (N_12738,N_11575,N_11159);
nand U12739 (N_12739,N_11973,N_11394);
nor U12740 (N_12740,N_10693,N_11340);
nor U12741 (N_12741,N_11988,N_11600);
and U12742 (N_12742,N_10764,N_11565);
or U12743 (N_12743,N_11659,N_10651);
and U12744 (N_12744,N_11508,N_11244);
or U12745 (N_12745,N_11317,N_10823);
and U12746 (N_12746,N_11436,N_11578);
xor U12747 (N_12747,N_11457,N_10751);
nor U12748 (N_12748,N_10975,N_11878);
and U12749 (N_12749,N_10972,N_10908);
xnor U12750 (N_12750,N_10836,N_11010);
or U12751 (N_12751,N_10890,N_11374);
or U12752 (N_12752,N_11700,N_11144);
xnor U12753 (N_12753,N_10602,N_10572);
or U12754 (N_12754,N_11425,N_11090);
and U12755 (N_12755,N_11094,N_11684);
nor U12756 (N_12756,N_11822,N_10738);
or U12757 (N_12757,N_10534,N_11908);
nand U12758 (N_12758,N_11753,N_11722);
and U12759 (N_12759,N_11047,N_11374);
or U12760 (N_12760,N_10727,N_11033);
xor U12761 (N_12761,N_11622,N_11666);
nand U12762 (N_12762,N_11673,N_10606);
nand U12763 (N_12763,N_11544,N_10897);
nor U12764 (N_12764,N_10531,N_10658);
or U12765 (N_12765,N_11628,N_11290);
xor U12766 (N_12766,N_11358,N_11066);
xnor U12767 (N_12767,N_10852,N_10619);
and U12768 (N_12768,N_11473,N_11646);
nand U12769 (N_12769,N_11583,N_10908);
or U12770 (N_12770,N_11150,N_11461);
or U12771 (N_12771,N_10660,N_11639);
xor U12772 (N_12772,N_11676,N_11669);
xnor U12773 (N_12773,N_11303,N_10748);
or U12774 (N_12774,N_10833,N_10624);
and U12775 (N_12775,N_11874,N_11571);
nand U12776 (N_12776,N_11344,N_11017);
or U12777 (N_12777,N_10980,N_10928);
xor U12778 (N_12778,N_11657,N_10554);
xor U12779 (N_12779,N_11745,N_11341);
and U12780 (N_12780,N_11314,N_11332);
nor U12781 (N_12781,N_10870,N_11724);
or U12782 (N_12782,N_10774,N_11229);
and U12783 (N_12783,N_10590,N_11142);
xnor U12784 (N_12784,N_11575,N_11672);
nor U12785 (N_12785,N_10868,N_11081);
and U12786 (N_12786,N_11522,N_10739);
nand U12787 (N_12787,N_11247,N_11445);
or U12788 (N_12788,N_10646,N_11469);
nor U12789 (N_12789,N_11524,N_10879);
xor U12790 (N_12790,N_10966,N_10962);
or U12791 (N_12791,N_11195,N_11867);
nand U12792 (N_12792,N_11244,N_10798);
and U12793 (N_12793,N_11179,N_11587);
or U12794 (N_12794,N_10605,N_11200);
nand U12795 (N_12795,N_11363,N_11535);
and U12796 (N_12796,N_11821,N_10747);
nor U12797 (N_12797,N_10629,N_11119);
nand U12798 (N_12798,N_10841,N_11477);
xor U12799 (N_12799,N_10698,N_10501);
nand U12800 (N_12800,N_10898,N_10833);
nand U12801 (N_12801,N_11787,N_11279);
xnor U12802 (N_12802,N_11916,N_10528);
xnor U12803 (N_12803,N_11051,N_10896);
nand U12804 (N_12804,N_11546,N_11909);
xnor U12805 (N_12805,N_10992,N_11167);
and U12806 (N_12806,N_11859,N_11904);
or U12807 (N_12807,N_10537,N_11862);
nor U12808 (N_12808,N_11922,N_11557);
and U12809 (N_12809,N_10858,N_11520);
nand U12810 (N_12810,N_10756,N_11587);
or U12811 (N_12811,N_11234,N_10710);
or U12812 (N_12812,N_11823,N_10858);
nor U12813 (N_12813,N_11556,N_11265);
nor U12814 (N_12814,N_10538,N_10825);
xor U12815 (N_12815,N_11170,N_11566);
nand U12816 (N_12816,N_11318,N_11434);
xnor U12817 (N_12817,N_11862,N_11876);
nor U12818 (N_12818,N_11317,N_11671);
xor U12819 (N_12819,N_11914,N_11599);
nand U12820 (N_12820,N_10837,N_11023);
or U12821 (N_12821,N_11066,N_11389);
nor U12822 (N_12822,N_10757,N_10879);
and U12823 (N_12823,N_11675,N_11360);
or U12824 (N_12824,N_11152,N_11908);
xor U12825 (N_12825,N_11746,N_11328);
and U12826 (N_12826,N_10728,N_11100);
and U12827 (N_12827,N_11879,N_11944);
or U12828 (N_12828,N_11646,N_10752);
xor U12829 (N_12829,N_11074,N_11006);
xnor U12830 (N_12830,N_10699,N_11537);
nor U12831 (N_12831,N_11535,N_11278);
nand U12832 (N_12832,N_11976,N_11329);
nand U12833 (N_12833,N_11009,N_10727);
xor U12834 (N_12834,N_11722,N_11250);
xnor U12835 (N_12835,N_10552,N_10546);
or U12836 (N_12836,N_10720,N_11221);
nand U12837 (N_12837,N_11195,N_10915);
and U12838 (N_12838,N_10797,N_10725);
nor U12839 (N_12839,N_11418,N_11387);
xor U12840 (N_12840,N_10711,N_11031);
xor U12841 (N_12841,N_11052,N_11532);
and U12842 (N_12842,N_11862,N_10768);
nand U12843 (N_12843,N_11820,N_11808);
and U12844 (N_12844,N_11670,N_10870);
nor U12845 (N_12845,N_10632,N_10674);
xor U12846 (N_12846,N_10505,N_11890);
nor U12847 (N_12847,N_11053,N_11842);
nor U12848 (N_12848,N_11859,N_10693);
xnor U12849 (N_12849,N_10848,N_11751);
nand U12850 (N_12850,N_11314,N_10526);
nand U12851 (N_12851,N_10818,N_11325);
nand U12852 (N_12852,N_11060,N_10528);
nand U12853 (N_12853,N_11730,N_10889);
or U12854 (N_12854,N_11076,N_10637);
nand U12855 (N_12855,N_11973,N_11794);
and U12856 (N_12856,N_11787,N_10989);
and U12857 (N_12857,N_11483,N_11285);
or U12858 (N_12858,N_10550,N_10505);
xnor U12859 (N_12859,N_10765,N_11006);
nor U12860 (N_12860,N_10757,N_11638);
or U12861 (N_12861,N_11963,N_11281);
xnor U12862 (N_12862,N_10905,N_11699);
nand U12863 (N_12863,N_11672,N_11611);
nor U12864 (N_12864,N_11618,N_11837);
or U12865 (N_12865,N_11438,N_10968);
and U12866 (N_12866,N_11694,N_11444);
and U12867 (N_12867,N_11535,N_10528);
and U12868 (N_12868,N_11495,N_11538);
or U12869 (N_12869,N_10562,N_11435);
and U12870 (N_12870,N_11098,N_11542);
nand U12871 (N_12871,N_11819,N_11064);
or U12872 (N_12872,N_11400,N_11768);
nand U12873 (N_12873,N_10995,N_11012);
or U12874 (N_12874,N_10749,N_11651);
nor U12875 (N_12875,N_11855,N_10810);
nor U12876 (N_12876,N_11236,N_11220);
and U12877 (N_12877,N_11190,N_10996);
or U12878 (N_12878,N_11479,N_11559);
or U12879 (N_12879,N_10867,N_11005);
and U12880 (N_12880,N_11845,N_11032);
nor U12881 (N_12881,N_11953,N_11484);
xnor U12882 (N_12882,N_11516,N_11461);
or U12883 (N_12883,N_10585,N_10765);
nor U12884 (N_12884,N_10821,N_11320);
xnor U12885 (N_12885,N_11349,N_10551);
or U12886 (N_12886,N_11732,N_10601);
nor U12887 (N_12887,N_10814,N_11066);
xnor U12888 (N_12888,N_11246,N_11545);
or U12889 (N_12889,N_11221,N_11466);
xnor U12890 (N_12890,N_11610,N_11797);
or U12891 (N_12891,N_11802,N_10754);
and U12892 (N_12892,N_10605,N_10928);
nand U12893 (N_12893,N_11302,N_11709);
and U12894 (N_12894,N_11904,N_10882);
xnor U12895 (N_12895,N_11509,N_10774);
nor U12896 (N_12896,N_10769,N_11872);
and U12897 (N_12897,N_11244,N_11887);
xor U12898 (N_12898,N_11559,N_11233);
nor U12899 (N_12899,N_11590,N_11203);
nor U12900 (N_12900,N_10556,N_10746);
xnor U12901 (N_12901,N_10564,N_11877);
and U12902 (N_12902,N_10503,N_11543);
nor U12903 (N_12903,N_11161,N_11088);
and U12904 (N_12904,N_11571,N_11710);
or U12905 (N_12905,N_10604,N_11114);
or U12906 (N_12906,N_11006,N_10545);
nand U12907 (N_12907,N_11264,N_10578);
or U12908 (N_12908,N_11729,N_10690);
or U12909 (N_12909,N_10511,N_10767);
or U12910 (N_12910,N_11950,N_11579);
nor U12911 (N_12911,N_11986,N_11450);
and U12912 (N_12912,N_11817,N_11810);
or U12913 (N_12913,N_10605,N_10515);
nor U12914 (N_12914,N_10585,N_10815);
and U12915 (N_12915,N_11939,N_10790);
and U12916 (N_12916,N_11012,N_11519);
nand U12917 (N_12917,N_11268,N_11669);
and U12918 (N_12918,N_10937,N_11074);
xnor U12919 (N_12919,N_10859,N_11416);
xor U12920 (N_12920,N_10806,N_11791);
xnor U12921 (N_12921,N_10976,N_10607);
nand U12922 (N_12922,N_11062,N_11708);
nand U12923 (N_12923,N_11752,N_10853);
xnor U12924 (N_12924,N_11801,N_11912);
and U12925 (N_12925,N_10753,N_11566);
xor U12926 (N_12926,N_10626,N_10637);
nand U12927 (N_12927,N_10511,N_11629);
and U12928 (N_12928,N_11697,N_11514);
nor U12929 (N_12929,N_11505,N_10785);
and U12930 (N_12930,N_11683,N_11557);
nand U12931 (N_12931,N_11764,N_11824);
and U12932 (N_12932,N_11459,N_11244);
nand U12933 (N_12933,N_10619,N_11372);
nand U12934 (N_12934,N_10689,N_11346);
or U12935 (N_12935,N_11192,N_11853);
or U12936 (N_12936,N_10966,N_11922);
and U12937 (N_12937,N_10904,N_11389);
xor U12938 (N_12938,N_11408,N_11546);
nor U12939 (N_12939,N_11230,N_10672);
or U12940 (N_12940,N_11825,N_10898);
nand U12941 (N_12941,N_11164,N_10871);
or U12942 (N_12942,N_10720,N_11280);
nor U12943 (N_12943,N_11043,N_11877);
nand U12944 (N_12944,N_10575,N_11021);
and U12945 (N_12945,N_11269,N_11527);
or U12946 (N_12946,N_10890,N_10799);
nand U12947 (N_12947,N_11654,N_11093);
and U12948 (N_12948,N_10753,N_11426);
nand U12949 (N_12949,N_11039,N_11952);
nand U12950 (N_12950,N_10541,N_10543);
and U12951 (N_12951,N_11774,N_11123);
and U12952 (N_12952,N_10872,N_10925);
and U12953 (N_12953,N_11492,N_11091);
and U12954 (N_12954,N_11512,N_11805);
nor U12955 (N_12955,N_10810,N_11984);
nand U12956 (N_12956,N_11006,N_11603);
nand U12957 (N_12957,N_10835,N_11777);
nor U12958 (N_12958,N_11580,N_10590);
nand U12959 (N_12959,N_10654,N_11689);
xnor U12960 (N_12960,N_11670,N_11215);
nor U12961 (N_12961,N_10884,N_11797);
nand U12962 (N_12962,N_10532,N_10775);
or U12963 (N_12963,N_10982,N_11676);
nor U12964 (N_12964,N_10822,N_11257);
and U12965 (N_12965,N_11833,N_11018);
or U12966 (N_12966,N_10902,N_11580);
nor U12967 (N_12967,N_11015,N_11463);
nand U12968 (N_12968,N_11243,N_11701);
or U12969 (N_12969,N_10536,N_11884);
nand U12970 (N_12970,N_11457,N_11907);
xor U12971 (N_12971,N_10961,N_11172);
nor U12972 (N_12972,N_11786,N_11687);
nor U12973 (N_12973,N_10950,N_10819);
and U12974 (N_12974,N_11505,N_10604);
or U12975 (N_12975,N_11234,N_11844);
nor U12976 (N_12976,N_11247,N_10525);
nand U12977 (N_12977,N_11271,N_10988);
and U12978 (N_12978,N_10770,N_11630);
nor U12979 (N_12979,N_11099,N_11577);
nor U12980 (N_12980,N_11824,N_10926);
or U12981 (N_12981,N_11259,N_11332);
xor U12982 (N_12982,N_11507,N_11363);
nor U12983 (N_12983,N_10848,N_11063);
and U12984 (N_12984,N_11511,N_11051);
xor U12985 (N_12985,N_11211,N_11926);
or U12986 (N_12986,N_10695,N_11839);
nor U12987 (N_12987,N_10674,N_11247);
nor U12988 (N_12988,N_11658,N_10663);
or U12989 (N_12989,N_11334,N_10966);
nand U12990 (N_12990,N_11773,N_11899);
or U12991 (N_12991,N_11481,N_11155);
xnor U12992 (N_12992,N_11856,N_11948);
and U12993 (N_12993,N_11838,N_11239);
nor U12994 (N_12994,N_11313,N_10773);
or U12995 (N_12995,N_11511,N_11174);
xor U12996 (N_12996,N_11548,N_11596);
or U12997 (N_12997,N_10994,N_10692);
nand U12998 (N_12998,N_10677,N_10873);
or U12999 (N_12999,N_11434,N_10647);
nor U13000 (N_13000,N_11596,N_11304);
xnor U13001 (N_13001,N_11168,N_11041);
nor U13002 (N_13002,N_11906,N_10986);
or U13003 (N_13003,N_11171,N_11509);
nor U13004 (N_13004,N_10909,N_10731);
and U13005 (N_13005,N_10879,N_11971);
nand U13006 (N_13006,N_10646,N_11882);
nand U13007 (N_13007,N_11379,N_10745);
xnor U13008 (N_13008,N_11262,N_10511);
and U13009 (N_13009,N_11101,N_11519);
nor U13010 (N_13010,N_11603,N_10868);
xor U13011 (N_13011,N_11435,N_11765);
and U13012 (N_13012,N_10536,N_10687);
nand U13013 (N_13013,N_10944,N_10889);
nor U13014 (N_13014,N_11511,N_11392);
nor U13015 (N_13015,N_10575,N_10555);
or U13016 (N_13016,N_10933,N_11989);
or U13017 (N_13017,N_11368,N_10658);
and U13018 (N_13018,N_11301,N_11068);
nand U13019 (N_13019,N_11133,N_11604);
or U13020 (N_13020,N_11571,N_10915);
or U13021 (N_13021,N_11934,N_11535);
or U13022 (N_13022,N_10688,N_11710);
xor U13023 (N_13023,N_11847,N_11936);
xor U13024 (N_13024,N_11416,N_11741);
nor U13025 (N_13025,N_11806,N_11288);
and U13026 (N_13026,N_11126,N_11149);
or U13027 (N_13027,N_11649,N_11820);
xor U13028 (N_13028,N_10506,N_10983);
xor U13029 (N_13029,N_11021,N_11325);
nand U13030 (N_13030,N_11163,N_11314);
nand U13031 (N_13031,N_10693,N_10975);
and U13032 (N_13032,N_10598,N_11409);
or U13033 (N_13033,N_10749,N_11948);
xnor U13034 (N_13034,N_11483,N_10586);
or U13035 (N_13035,N_10946,N_11080);
xnor U13036 (N_13036,N_11649,N_11582);
nor U13037 (N_13037,N_10935,N_10598);
nand U13038 (N_13038,N_10792,N_11038);
and U13039 (N_13039,N_11811,N_11731);
xor U13040 (N_13040,N_11412,N_11948);
nor U13041 (N_13041,N_10726,N_11649);
nand U13042 (N_13042,N_11001,N_11797);
or U13043 (N_13043,N_11503,N_11101);
and U13044 (N_13044,N_11858,N_11514);
or U13045 (N_13045,N_11130,N_10694);
nand U13046 (N_13046,N_11297,N_11940);
or U13047 (N_13047,N_11802,N_11100);
xor U13048 (N_13048,N_11021,N_11097);
or U13049 (N_13049,N_11378,N_10622);
or U13050 (N_13050,N_11845,N_10826);
or U13051 (N_13051,N_11401,N_10519);
and U13052 (N_13052,N_11038,N_11620);
nand U13053 (N_13053,N_11006,N_10741);
and U13054 (N_13054,N_11156,N_11209);
xnor U13055 (N_13055,N_11348,N_11799);
or U13056 (N_13056,N_11230,N_11682);
nand U13057 (N_13057,N_11659,N_11738);
or U13058 (N_13058,N_11494,N_10806);
or U13059 (N_13059,N_11299,N_11429);
and U13060 (N_13060,N_11856,N_11074);
nor U13061 (N_13061,N_11831,N_11653);
nor U13062 (N_13062,N_11814,N_10680);
or U13063 (N_13063,N_10772,N_10725);
or U13064 (N_13064,N_11728,N_10908);
nor U13065 (N_13065,N_10940,N_11930);
and U13066 (N_13066,N_11527,N_11375);
nor U13067 (N_13067,N_11845,N_11289);
xor U13068 (N_13068,N_10858,N_10714);
or U13069 (N_13069,N_11246,N_11752);
nor U13070 (N_13070,N_11292,N_11046);
and U13071 (N_13071,N_11807,N_11341);
and U13072 (N_13072,N_11823,N_10802);
and U13073 (N_13073,N_11716,N_11718);
and U13074 (N_13074,N_11492,N_11164);
and U13075 (N_13075,N_10501,N_11982);
nor U13076 (N_13076,N_11696,N_10956);
xor U13077 (N_13077,N_10907,N_10639);
nor U13078 (N_13078,N_11228,N_11781);
nor U13079 (N_13079,N_10999,N_10529);
and U13080 (N_13080,N_10538,N_11720);
xor U13081 (N_13081,N_10884,N_11237);
xnor U13082 (N_13082,N_11467,N_10771);
nand U13083 (N_13083,N_11162,N_10826);
or U13084 (N_13084,N_11384,N_11030);
and U13085 (N_13085,N_11679,N_10591);
or U13086 (N_13086,N_11288,N_10521);
or U13087 (N_13087,N_11386,N_10909);
nor U13088 (N_13088,N_10911,N_10733);
nand U13089 (N_13089,N_11736,N_11372);
or U13090 (N_13090,N_10501,N_10744);
nor U13091 (N_13091,N_11849,N_11282);
xnor U13092 (N_13092,N_11431,N_11919);
xnor U13093 (N_13093,N_11529,N_11144);
nand U13094 (N_13094,N_11718,N_11405);
xnor U13095 (N_13095,N_10789,N_11471);
nand U13096 (N_13096,N_10752,N_10726);
and U13097 (N_13097,N_11936,N_11099);
xor U13098 (N_13098,N_10750,N_10730);
xnor U13099 (N_13099,N_10573,N_10827);
nor U13100 (N_13100,N_11452,N_10736);
nand U13101 (N_13101,N_11629,N_11874);
and U13102 (N_13102,N_11540,N_10795);
nor U13103 (N_13103,N_11335,N_10558);
xor U13104 (N_13104,N_11457,N_11737);
and U13105 (N_13105,N_11741,N_11469);
nand U13106 (N_13106,N_11343,N_11088);
and U13107 (N_13107,N_10870,N_11349);
or U13108 (N_13108,N_10809,N_11861);
and U13109 (N_13109,N_11056,N_10897);
nor U13110 (N_13110,N_11933,N_11386);
nand U13111 (N_13111,N_11262,N_11322);
xnor U13112 (N_13112,N_11631,N_11908);
xnor U13113 (N_13113,N_11334,N_11180);
or U13114 (N_13114,N_11614,N_11432);
and U13115 (N_13115,N_10961,N_10676);
xnor U13116 (N_13116,N_11544,N_11877);
nand U13117 (N_13117,N_11595,N_11476);
and U13118 (N_13118,N_11792,N_11870);
and U13119 (N_13119,N_10599,N_11934);
or U13120 (N_13120,N_11938,N_11582);
and U13121 (N_13121,N_11705,N_11520);
nand U13122 (N_13122,N_11008,N_11363);
nor U13123 (N_13123,N_11990,N_11088);
or U13124 (N_13124,N_10858,N_11233);
nand U13125 (N_13125,N_11557,N_11074);
xor U13126 (N_13126,N_11764,N_11844);
nand U13127 (N_13127,N_11624,N_10628);
xnor U13128 (N_13128,N_11916,N_10782);
nor U13129 (N_13129,N_10623,N_11552);
nor U13130 (N_13130,N_10619,N_11482);
nand U13131 (N_13131,N_11498,N_10714);
and U13132 (N_13132,N_10619,N_11868);
xnor U13133 (N_13133,N_11018,N_10716);
or U13134 (N_13134,N_10831,N_11803);
nor U13135 (N_13135,N_10725,N_11703);
xnor U13136 (N_13136,N_10561,N_10760);
nand U13137 (N_13137,N_11702,N_11139);
and U13138 (N_13138,N_11276,N_11892);
nor U13139 (N_13139,N_11344,N_10534);
nand U13140 (N_13140,N_10962,N_11508);
or U13141 (N_13141,N_11468,N_11820);
nor U13142 (N_13142,N_10509,N_10593);
xnor U13143 (N_13143,N_10725,N_11118);
and U13144 (N_13144,N_10561,N_10774);
and U13145 (N_13145,N_11109,N_11537);
nand U13146 (N_13146,N_11844,N_11967);
and U13147 (N_13147,N_11323,N_11263);
or U13148 (N_13148,N_11424,N_10830);
xor U13149 (N_13149,N_11841,N_10517);
or U13150 (N_13150,N_10954,N_10952);
and U13151 (N_13151,N_11076,N_11997);
nor U13152 (N_13152,N_11742,N_11519);
and U13153 (N_13153,N_11389,N_11035);
nand U13154 (N_13154,N_11384,N_11287);
and U13155 (N_13155,N_11926,N_11617);
nor U13156 (N_13156,N_10835,N_11817);
or U13157 (N_13157,N_11460,N_11669);
nand U13158 (N_13158,N_11289,N_11250);
nand U13159 (N_13159,N_11600,N_11347);
nor U13160 (N_13160,N_10793,N_11324);
nand U13161 (N_13161,N_10833,N_10944);
and U13162 (N_13162,N_10681,N_11789);
and U13163 (N_13163,N_10891,N_10824);
nor U13164 (N_13164,N_11942,N_11723);
and U13165 (N_13165,N_10571,N_11318);
nor U13166 (N_13166,N_10850,N_11676);
nand U13167 (N_13167,N_10980,N_11595);
nand U13168 (N_13168,N_11853,N_10993);
or U13169 (N_13169,N_11335,N_10580);
or U13170 (N_13170,N_10708,N_11251);
or U13171 (N_13171,N_11920,N_10630);
nand U13172 (N_13172,N_11789,N_11018);
nor U13173 (N_13173,N_10868,N_11042);
or U13174 (N_13174,N_11222,N_11322);
or U13175 (N_13175,N_11571,N_10729);
nand U13176 (N_13176,N_11851,N_11687);
xnor U13177 (N_13177,N_11775,N_11039);
nor U13178 (N_13178,N_11116,N_11958);
nor U13179 (N_13179,N_10531,N_11659);
or U13180 (N_13180,N_10817,N_10576);
and U13181 (N_13181,N_10869,N_11053);
or U13182 (N_13182,N_11847,N_11567);
and U13183 (N_13183,N_11610,N_11479);
nor U13184 (N_13184,N_10868,N_11263);
and U13185 (N_13185,N_10811,N_10827);
nand U13186 (N_13186,N_10913,N_11884);
nand U13187 (N_13187,N_11719,N_11919);
nor U13188 (N_13188,N_11470,N_11731);
and U13189 (N_13189,N_11412,N_11428);
xor U13190 (N_13190,N_10650,N_11413);
nor U13191 (N_13191,N_11162,N_11135);
or U13192 (N_13192,N_11393,N_10520);
xor U13193 (N_13193,N_11662,N_10991);
nand U13194 (N_13194,N_11057,N_11813);
and U13195 (N_13195,N_11133,N_11271);
or U13196 (N_13196,N_11955,N_10724);
xor U13197 (N_13197,N_11712,N_11612);
and U13198 (N_13198,N_11830,N_11978);
nand U13199 (N_13199,N_10522,N_11781);
nor U13200 (N_13200,N_11167,N_11462);
nand U13201 (N_13201,N_11758,N_10508);
nand U13202 (N_13202,N_10979,N_10668);
nor U13203 (N_13203,N_10710,N_11914);
nor U13204 (N_13204,N_11871,N_11316);
and U13205 (N_13205,N_11877,N_10812);
and U13206 (N_13206,N_11333,N_11797);
or U13207 (N_13207,N_11666,N_11102);
nand U13208 (N_13208,N_11701,N_10637);
nor U13209 (N_13209,N_10986,N_11884);
nand U13210 (N_13210,N_10995,N_11133);
and U13211 (N_13211,N_11468,N_11076);
xnor U13212 (N_13212,N_11450,N_10956);
and U13213 (N_13213,N_10707,N_11723);
nand U13214 (N_13214,N_11009,N_11041);
and U13215 (N_13215,N_10640,N_10541);
nor U13216 (N_13216,N_10567,N_11443);
nand U13217 (N_13217,N_11702,N_11842);
and U13218 (N_13218,N_11732,N_11375);
xnor U13219 (N_13219,N_11277,N_11880);
and U13220 (N_13220,N_10634,N_11868);
nor U13221 (N_13221,N_11922,N_11027);
and U13222 (N_13222,N_11329,N_11347);
nor U13223 (N_13223,N_11729,N_11011);
or U13224 (N_13224,N_11742,N_11611);
xnor U13225 (N_13225,N_11973,N_11163);
nor U13226 (N_13226,N_11529,N_11874);
nand U13227 (N_13227,N_11866,N_11159);
xor U13228 (N_13228,N_11425,N_11245);
and U13229 (N_13229,N_11882,N_11521);
and U13230 (N_13230,N_11426,N_11605);
nand U13231 (N_13231,N_11212,N_10812);
nor U13232 (N_13232,N_11630,N_10660);
and U13233 (N_13233,N_10838,N_10922);
or U13234 (N_13234,N_10617,N_11451);
xnor U13235 (N_13235,N_11811,N_11740);
or U13236 (N_13236,N_11400,N_11617);
nand U13237 (N_13237,N_11688,N_10735);
nand U13238 (N_13238,N_11985,N_10834);
xor U13239 (N_13239,N_11896,N_10611);
xor U13240 (N_13240,N_11845,N_11585);
or U13241 (N_13241,N_11718,N_11626);
and U13242 (N_13242,N_11210,N_11427);
nand U13243 (N_13243,N_10998,N_10875);
xor U13244 (N_13244,N_10572,N_11297);
nand U13245 (N_13245,N_11661,N_11064);
and U13246 (N_13246,N_11007,N_10529);
and U13247 (N_13247,N_11810,N_11973);
nor U13248 (N_13248,N_10886,N_11735);
or U13249 (N_13249,N_11502,N_10590);
nand U13250 (N_13250,N_11110,N_11258);
nor U13251 (N_13251,N_11217,N_11881);
nand U13252 (N_13252,N_11029,N_11262);
and U13253 (N_13253,N_10596,N_11909);
nand U13254 (N_13254,N_11873,N_10569);
nor U13255 (N_13255,N_11821,N_10775);
xnor U13256 (N_13256,N_10556,N_10898);
and U13257 (N_13257,N_11986,N_10509);
and U13258 (N_13258,N_10985,N_11605);
or U13259 (N_13259,N_11410,N_11655);
nand U13260 (N_13260,N_11387,N_10561);
and U13261 (N_13261,N_11393,N_10913);
and U13262 (N_13262,N_11544,N_11892);
and U13263 (N_13263,N_10704,N_11982);
and U13264 (N_13264,N_11340,N_10510);
nor U13265 (N_13265,N_10809,N_11799);
nor U13266 (N_13266,N_10867,N_11737);
nor U13267 (N_13267,N_11513,N_11439);
or U13268 (N_13268,N_11820,N_11964);
nor U13269 (N_13269,N_11827,N_11059);
nor U13270 (N_13270,N_11248,N_11537);
or U13271 (N_13271,N_11113,N_10889);
nor U13272 (N_13272,N_10646,N_11611);
or U13273 (N_13273,N_11407,N_11990);
or U13274 (N_13274,N_11221,N_11230);
nor U13275 (N_13275,N_11524,N_11356);
xor U13276 (N_13276,N_11251,N_11142);
nor U13277 (N_13277,N_10532,N_11975);
and U13278 (N_13278,N_11417,N_11893);
or U13279 (N_13279,N_11306,N_11850);
nor U13280 (N_13280,N_11622,N_11024);
nand U13281 (N_13281,N_11472,N_11298);
nand U13282 (N_13282,N_11943,N_10767);
and U13283 (N_13283,N_11103,N_10520);
and U13284 (N_13284,N_10576,N_11483);
nor U13285 (N_13285,N_11607,N_11244);
xor U13286 (N_13286,N_11861,N_11480);
and U13287 (N_13287,N_11790,N_10600);
and U13288 (N_13288,N_11588,N_11967);
and U13289 (N_13289,N_11675,N_10738);
xor U13290 (N_13290,N_11020,N_10937);
or U13291 (N_13291,N_10915,N_11456);
xor U13292 (N_13292,N_10510,N_10574);
and U13293 (N_13293,N_11383,N_11218);
nor U13294 (N_13294,N_11563,N_11422);
or U13295 (N_13295,N_10694,N_11980);
xor U13296 (N_13296,N_11132,N_11660);
xor U13297 (N_13297,N_10719,N_10765);
nand U13298 (N_13298,N_11527,N_11266);
xor U13299 (N_13299,N_11513,N_10777);
or U13300 (N_13300,N_10771,N_10595);
and U13301 (N_13301,N_11847,N_11032);
xor U13302 (N_13302,N_10941,N_11235);
or U13303 (N_13303,N_10935,N_11564);
xnor U13304 (N_13304,N_10610,N_11419);
nor U13305 (N_13305,N_10732,N_10815);
or U13306 (N_13306,N_10860,N_10880);
xnor U13307 (N_13307,N_10598,N_11580);
and U13308 (N_13308,N_11907,N_11562);
xnor U13309 (N_13309,N_10703,N_11118);
nor U13310 (N_13310,N_11889,N_10809);
and U13311 (N_13311,N_10716,N_11139);
nor U13312 (N_13312,N_10567,N_11410);
nor U13313 (N_13313,N_11932,N_11452);
and U13314 (N_13314,N_11877,N_11721);
or U13315 (N_13315,N_10977,N_11051);
and U13316 (N_13316,N_10687,N_10647);
or U13317 (N_13317,N_11842,N_11952);
and U13318 (N_13318,N_10567,N_10940);
xor U13319 (N_13319,N_10507,N_11927);
xnor U13320 (N_13320,N_11248,N_10699);
or U13321 (N_13321,N_10928,N_10971);
xor U13322 (N_13322,N_11387,N_11365);
nand U13323 (N_13323,N_11990,N_11947);
or U13324 (N_13324,N_10702,N_11039);
and U13325 (N_13325,N_11624,N_11682);
nand U13326 (N_13326,N_11317,N_11700);
and U13327 (N_13327,N_11793,N_11840);
nand U13328 (N_13328,N_11393,N_11429);
nor U13329 (N_13329,N_11680,N_11308);
nor U13330 (N_13330,N_10828,N_10973);
and U13331 (N_13331,N_11670,N_11927);
xnor U13332 (N_13332,N_11768,N_11001);
and U13333 (N_13333,N_10758,N_10940);
nor U13334 (N_13334,N_11570,N_11701);
or U13335 (N_13335,N_11233,N_10690);
nor U13336 (N_13336,N_10772,N_11183);
nand U13337 (N_13337,N_11659,N_11436);
and U13338 (N_13338,N_11298,N_10905);
nor U13339 (N_13339,N_10608,N_11658);
or U13340 (N_13340,N_10654,N_10808);
nand U13341 (N_13341,N_11998,N_11893);
xnor U13342 (N_13342,N_10955,N_11324);
xnor U13343 (N_13343,N_11297,N_11283);
and U13344 (N_13344,N_10707,N_11174);
xnor U13345 (N_13345,N_11358,N_10774);
and U13346 (N_13346,N_11740,N_11058);
nand U13347 (N_13347,N_10917,N_11501);
and U13348 (N_13348,N_11769,N_11809);
nor U13349 (N_13349,N_11234,N_11120);
nand U13350 (N_13350,N_10950,N_11476);
nor U13351 (N_13351,N_11826,N_11399);
and U13352 (N_13352,N_11256,N_10916);
nand U13353 (N_13353,N_11785,N_11592);
nor U13354 (N_13354,N_11468,N_11409);
nand U13355 (N_13355,N_11804,N_11587);
or U13356 (N_13356,N_11916,N_11342);
nand U13357 (N_13357,N_10954,N_10633);
nor U13358 (N_13358,N_11563,N_11129);
xnor U13359 (N_13359,N_10807,N_10926);
or U13360 (N_13360,N_10881,N_10552);
and U13361 (N_13361,N_10662,N_10569);
xor U13362 (N_13362,N_11481,N_10557);
nor U13363 (N_13363,N_11527,N_11932);
xnor U13364 (N_13364,N_11049,N_11790);
and U13365 (N_13365,N_11776,N_10700);
xnor U13366 (N_13366,N_11689,N_10959);
and U13367 (N_13367,N_11568,N_11736);
nand U13368 (N_13368,N_10704,N_10539);
nand U13369 (N_13369,N_10649,N_10692);
nand U13370 (N_13370,N_10564,N_10974);
nand U13371 (N_13371,N_10615,N_11020);
and U13372 (N_13372,N_11882,N_10850);
xor U13373 (N_13373,N_10560,N_11689);
nand U13374 (N_13374,N_10763,N_11461);
and U13375 (N_13375,N_10821,N_10594);
and U13376 (N_13376,N_11760,N_10667);
and U13377 (N_13377,N_10786,N_11550);
nor U13378 (N_13378,N_11909,N_11610);
xnor U13379 (N_13379,N_11333,N_11942);
nand U13380 (N_13380,N_11296,N_10750);
nand U13381 (N_13381,N_11153,N_10564);
nor U13382 (N_13382,N_11909,N_11144);
nand U13383 (N_13383,N_11658,N_11480);
nand U13384 (N_13384,N_11603,N_10808);
nor U13385 (N_13385,N_11330,N_10908);
nor U13386 (N_13386,N_11805,N_11747);
xnor U13387 (N_13387,N_10585,N_11334);
xnor U13388 (N_13388,N_10831,N_10882);
nor U13389 (N_13389,N_11138,N_11934);
xor U13390 (N_13390,N_11891,N_11864);
nor U13391 (N_13391,N_10632,N_11764);
and U13392 (N_13392,N_11256,N_10893);
xor U13393 (N_13393,N_11684,N_11420);
xor U13394 (N_13394,N_11405,N_11062);
or U13395 (N_13395,N_10686,N_11547);
or U13396 (N_13396,N_11061,N_10753);
nand U13397 (N_13397,N_11930,N_11238);
and U13398 (N_13398,N_11761,N_11454);
xor U13399 (N_13399,N_10966,N_10910);
or U13400 (N_13400,N_11573,N_11549);
or U13401 (N_13401,N_11241,N_10618);
xnor U13402 (N_13402,N_10895,N_10885);
and U13403 (N_13403,N_10572,N_11717);
nand U13404 (N_13404,N_11494,N_11775);
nor U13405 (N_13405,N_11561,N_11335);
or U13406 (N_13406,N_11453,N_10777);
nor U13407 (N_13407,N_11154,N_11066);
nand U13408 (N_13408,N_11489,N_11218);
nand U13409 (N_13409,N_10912,N_10513);
nand U13410 (N_13410,N_11843,N_10687);
and U13411 (N_13411,N_11140,N_11557);
and U13412 (N_13412,N_11279,N_10987);
nor U13413 (N_13413,N_11256,N_11712);
nand U13414 (N_13414,N_11955,N_11542);
nand U13415 (N_13415,N_10675,N_11683);
nand U13416 (N_13416,N_11023,N_11353);
nor U13417 (N_13417,N_11286,N_11262);
nor U13418 (N_13418,N_11264,N_11314);
xnor U13419 (N_13419,N_10931,N_11338);
xnor U13420 (N_13420,N_11255,N_11531);
xnor U13421 (N_13421,N_11087,N_10627);
and U13422 (N_13422,N_11810,N_10555);
nand U13423 (N_13423,N_11892,N_11732);
nor U13424 (N_13424,N_11956,N_11624);
nand U13425 (N_13425,N_10946,N_11210);
or U13426 (N_13426,N_11535,N_11657);
nand U13427 (N_13427,N_11505,N_10688);
nand U13428 (N_13428,N_11719,N_10594);
or U13429 (N_13429,N_11386,N_11500);
nand U13430 (N_13430,N_11949,N_10673);
and U13431 (N_13431,N_10768,N_11577);
xor U13432 (N_13432,N_11868,N_11130);
nand U13433 (N_13433,N_11398,N_10898);
xor U13434 (N_13434,N_11777,N_10747);
xor U13435 (N_13435,N_10631,N_11190);
and U13436 (N_13436,N_11728,N_11155);
and U13437 (N_13437,N_11464,N_10616);
nor U13438 (N_13438,N_11500,N_11697);
nor U13439 (N_13439,N_10802,N_10803);
and U13440 (N_13440,N_10577,N_11613);
nand U13441 (N_13441,N_10825,N_10807);
nor U13442 (N_13442,N_11617,N_11572);
and U13443 (N_13443,N_10975,N_10504);
xor U13444 (N_13444,N_11386,N_10634);
nor U13445 (N_13445,N_11853,N_11773);
xor U13446 (N_13446,N_10559,N_11890);
and U13447 (N_13447,N_11276,N_11163);
or U13448 (N_13448,N_11884,N_11348);
and U13449 (N_13449,N_10745,N_10991);
or U13450 (N_13450,N_11526,N_11191);
or U13451 (N_13451,N_11703,N_11989);
xnor U13452 (N_13452,N_11324,N_11388);
nand U13453 (N_13453,N_11727,N_10585);
nor U13454 (N_13454,N_11286,N_11775);
nand U13455 (N_13455,N_10501,N_10954);
nand U13456 (N_13456,N_11621,N_11720);
xor U13457 (N_13457,N_11833,N_11117);
nand U13458 (N_13458,N_11475,N_11322);
nand U13459 (N_13459,N_11367,N_11058);
nand U13460 (N_13460,N_10638,N_10864);
xnor U13461 (N_13461,N_10607,N_10580);
nand U13462 (N_13462,N_11638,N_11713);
nand U13463 (N_13463,N_11206,N_11050);
or U13464 (N_13464,N_11222,N_10909);
nor U13465 (N_13465,N_10679,N_10510);
nor U13466 (N_13466,N_11619,N_11079);
nand U13467 (N_13467,N_10690,N_10695);
or U13468 (N_13468,N_11438,N_11672);
nor U13469 (N_13469,N_11896,N_11638);
and U13470 (N_13470,N_11416,N_11459);
nor U13471 (N_13471,N_11512,N_11946);
and U13472 (N_13472,N_11153,N_11662);
nand U13473 (N_13473,N_10644,N_11424);
nand U13474 (N_13474,N_10678,N_10518);
nand U13475 (N_13475,N_11467,N_10969);
and U13476 (N_13476,N_11864,N_10837);
nand U13477 (N_13477,N_11298,N_11116);
and U13478 (N_13478,N_10847,N_11181);
and U13479 (N_13479,N_10699,N_11487);
nand U13480 (N_13480,N_11061,N_11137);
nand U13481 (N_13481,N_11409,N_11734);
xor U13482 (N_13482,N_11647,N_10884);
nand U13483 (N_13483,N_11425,N_10668);
or U13484 (N_13484,N_11844,N_10501);
nor U13485 (N_13485,N_11752,N_11514);
or U13486 (N_13486,N_11778,N_10701);
nor U13487 (N_13487,N_11573,N_10888);
nand U13488 (N_13488,N_11153,N_11584);
and U13489 (N_13489,N_11370,N_11350);
nand U13490 (N_13490,N_11791,N_11918);
nor U13491 (N_13491,N_10811,N_11465);
nor U13492 (N_13492,N_10716,N_11124);
or U13493 (N_13493,N_11737,N_10939);
nor U13494 (N_13494,N_10643,N_11854);
xnor U13495 (N_13495,N_11869,N_11200);
nor U13496 (N_13496,N_10874,N_11976);
nor U13497 (N_13497,N_11365,N_11789);
nand U13498 (N_13498,N_11004,N_10682);
nand U13499 (N_13499,N_10868,N_11207);
xnor U13500 (N_13500,N_13250,N_12516);
or U13501 (N_13501,N_12287,N_13110);
xor U13502 (N_13502,N_12471,N_13465);
or U13503 (N_13503,N_13031,N_12401);
nor U13504 (N_13504,N_12804,N_12542);
or U13505 (N_13505,N_12129,N_12565);
nor U13506 (N_13506,N_12658,N_12829);
xor U13507 (N_13507,N_12189,N_12797);
nand U13508 (N_13508,N_12103,N_12692);
nand U13509 (N_13509,N_13446,N_12960);
nand U13510 (N_13510,N_12174,N_12119);
or U13511 (N_13511,N_12736,N_13231);
xor U13512 (N_13512,N_12980,N_13062);
and U13513 (N_13513,N_12904,N_13438);
and U13514 (N_13514,N_12262,N_13018);
or U13515 (N_13515,N_13156,N_13433);
and U13516 (N_13516,N_12579,N_12180);
or U13517 (N_13517,N_13176,N_12171);
or U13518 (N_13518,N_12237,N_13288);
and U13519 (N_13519,N_12780,N_12138);
xnor U13520 (N_13520,N_12790,N_12010);
nor U13521 (N_13521,N_12358,N_12774);
nand U13522 (N_13522,N_13450,N_12197);
or U13523 (N_13523,N_12686,N_13347);
and U13524 (N_13524,N_12803,N_12268);
nand U13525 (N_13525,N_13046,N_13320);
nor U13526 (N_13526,N_12207,N_13049);
nand U13527 (N_13527,N_12992,N_13361);
and U13528 (N_13528,N_12321,N_13030);
xnor U13529 (N_13529,N_12373,N_13101);
or U13530 (N_13530,N_13136,N_13096);
nand U13531 (N_13531,N_12532,N_12120);
or U13532 (N_13532,N_12559,N_12301);
nand U13533 (N_13533,N_12646,N_13319);
xor U13534 (N_13534,N_12061,N_13206);
or U13535 (N_13535,N_12648,N_12016);
nand U13536 (N_13536,N_12413,N_12640);
or U13537 (N_13537,N_12687,N_12914);
or U13538 (N_13538,N_12846,N_13190);
xor U13539 (N_13539,N_12680,N_12108);
xnor U13540 (N_13540,N_13473,N_13307);
and U13541 (N_13541,N_13374,N_13185);
and U13542 (N_13542,N_12372,N_12574);
or U13543 (N_13543,N_12758,N_12808);
and U13544 (N_13544,N_13195,N_13400);
or U13545 (N_13545,N_13172,N_12899);
xor U13546 (N_13546,N_13191,N_12799);
and U13547 (N_13547,N_13064,N_13067);
or U13548 (N_13548,N_13410,N_12578);
and U13549 (N_13549,N_13357,N_13302);
and U13550 (N_13550,N_12623,N_13178);
xor U13551 (N_13551,N_12481,N_13418);
and U13552 (N_13552,N_12206,N_12234);
xor U13553 (N_13553,N_12779,N_12344);
nand U13554 (N_13554,N_13069,N_12520);
xnor U13555 (N_13555,N_12946,N_12984);
xor U13556 (N_13556,N_13102,N_12932);
xnor U13557 (N_13557,N_13028,N_12998);
and U13558 (N_13558,N_13051,N_12053);
nor U13559 (N_13559,N_12540,N_12227);
nor U13560 (N_13560,N_12845,N_13128);
nor U13561 (N_13561,N_12606,N_13299);
nor U13562 (N_13562,N_12771,N_12494);
xor U13563 (N_13563,N_12558,N_13074);
xnor U13564 (N_13564,N_12722,N_12857);
xnor U13565 (N_13565,N_12734,N_12855);
nand U13566 (N_13566,N_12387,N_13164);
or U13567 (N_13567,N_12263,N_12751);
and U13568 (N_13568,N_12106,N_12560);
and U13569 (N_13569,N_13281,N_12918);
or U13570 (N_13570,N_13257,N_12209);
nor U13571 (N_13571,N_12659,N_13108);
and U13572 (N_13572,N_13114,N_12518);
nand U13573 (N_13573,N_12151,N_12312);
and U13574 (N_13574,N_13267,N_12726);
xor U13575 (N_13575,N_12337,N_13057);
nor U13576 (N_13576,N_12749,N_13032);
and U13577 (N_13577,N_12265,N_13271);
or U13578 (N_13578,N_13432,N_12419);
xor U13579 (N_13579,N_13039,N_12187);
and U13580 (N_13580,N_12205,N_12432);
and U13581 (N_13581,N_12110,N_12331);
and U13582 (N_13582,N_12698,N_12837);
and U13583 (N_13583,N_13423,N_12380);
xnor U13584 (N_13584,N_12477,N_12022);
xor U13585 (N_13585,N_13245,N_13447);
nor U13586 (N_13586,N_12224,N_13227);
and U13587 (N_13587,N_12140,N_12064);
nand U13588 (N_13588,N_12203,N_12328);
and U13589 (N_13589,N_13296,N_13263);
nand U13590 (N_13590,N_12299,N_12159);
xor U13591 (N_13591,N_12195,N_13265);
and U13592 (N_13592,N_12785,N_13020);
xor U13593 (N_13593,N_12585,N_12128);
nor U13594 (N_13594,N_12839,N_13088);
xor U13595 (N_13595,N_12525,N_12805);
or U13596 (N_13596,N_12100,N_13367);
xnor U13597 (N_13597,N_13170,N_12890);
xor U13598 (N_13598,N_13277,N_13181);
xor U13599 (N_13599,N_12356,N_13474);
xnor U13600 (N_13600,N_13397,N_12828);
xor U13601 (N_13601,N_12149,N_12215);
or U13602 (N_13602,N_12868,N_12063);
nor U13603 (N_13603,N_13480,N_13133);
nand U13604 (N_13604,N_13454,N_13405);
and U13605 (N_13605,N_13269,N_13255);
nand U13606 (N_13606,N_12915,N_13104);
or U13607 (N_13607,N_13484,N_12093);
nand U13608 (N_13608,N_13216,N_12427);
or U13609 (N_13609,N_12399,N_12541);
nand U13610 (N_13610,N_13158,N_13481);
and U13611 (N_13611,N_12647,N_12523);
or U13612 (N_13612,N_12367,N_12360);
nor U13613 (N_13613,N_12274,N_13217);
nor U13614 (N_13614,N_12934,N_12663);
nand U13615 (N_13615,N_13371,N_13065);
nand U13616 (N_13616,N_12694,N_12192);
and U13617 (N_13617,N_13463,N_12533);
nor U13618 (N_13618,N_12397,N_13370);
or U13619 (N_13619,N_12352,N_13259);
nor U13620 (N_13620,N_13122,N_13115);
and U13621 (N_13621,N_12261,N_12618);
nand U13622 (N_13622,N_13442,N_12143);
or U13623 (N_13623,N_12550,N_12690);
xor U13624 (N_13624,N_12544,N_12310);
and U13625 (N_13625,N_12019,N_12201);
and U13626 (N_13626,N_13396,N_12316);
xor U13627 (N_13627,N_13163,N_12089);
nor U13628 (N_13628,N_13013,N_12457);
and U13629 (N_13629,N_12404,N_12912);
nor U13630 (N_13630,N_12723,N_12188);
nand U13631 (N_13631,N_13244,N_13055);
and U13632 (N_13632,N_12843,N_12377);
or U13633 (N_13633,N_12666,N_13358);
and U13634 (N_13634,N_12077,N_12988);
nand U13635 (N_13635,N_12638,N_13381);
or U13636 (N_13636,N_12038,N_12292);
and U13637 (N_13637,N_13173,N_12220);
xor U13638 (N_13638,N_12500,N_12593);
nand U13639 (N_13639,N_12581,N_12873);
xor U13640 (N_13640,N_13016,N_12583);
nor U13641 (N_13641,N_13360,N_13386);
nor U13642 (N_13642,N_12236,N_13004);
or U13643 (N_13643,N_13017,N_12231);
or U13644 (N_13644,N_13006,N_12990);
nor U13645 (N_13645,N_12555,N_12929);
nand U13646 (N_13646,N_12625,N_12517);
nand U13647 (N_13647,N_12892,N_13313);
nor U13648 (N_13648,N_12153,N_12860);
nand U13649 (N_13649,N_12307,N_13027);
nand U13650 (N_13650,N_12003,N_13350);
and U13651 (N_13651,N_13434,N_12973);
xor U13652 (N_13652,N_12416,N_13234);
nor U13653 (N_13653,N_12080,N_12567);
nand U13654 (N_13654,N_12178,N_12341);
nand U13655 (N_13655,N_12781,N_12735);
nand U13656 (N_13656,N_12649,N_12591);
xnor U13657 (N_13657,N_12505,N_13311);
xor U13658 (N_13658,N_12452,N_13460);
or U13659 (N_13659,N_12357,N_12744);
or U13660 (N_13660,N_12166,N_13141);
xnor U13661 (N_13661,N_13127,N_12461);
nand U13662 (N_13662,N_12613,N_12114);
nor U13663 (N_13663,N_12628,N_13148);
nand U13664 (N_13664,N_12831,N_12139);
and U13665 (N_13665,N_12130,N_12013);
and U13666 (N_13666,N_12249,N_13002);
nor U13667 (N_13667,N_12497,N_13033);
and U13668 (N_13668,N_12813,N_12222);
nand U13669 (N_13669,N_12664,N_13470);
nand U13670 (N_13670,N_12524,N_12712);
nand U13671 (N_13671,N_13107,N_12051);
and U13672 (N_13672,N_12256,N_12414);
nand U13673 (N_13673,N_12821,N_12029);
xnor U13674 (N_13674,N_12798,N_12807);
or U13675 (N_13675,N_13284,N_12878);
or U13676 (N_13676,N_12296,N_13198);
nor U13677 (N_13677,N_12871,N_12162);
xnor U13678 (N_13678,N_12859,N_13214);
nand U13679 (N_13679,N_12463,N_13001);
nand U13680 (N_13680,N_12787,N_13278);
nor U13681 (N_13681,N_12247,N_13152);
nor U13682 (N_13682,N_12791,N_12651);
and U13683 (N_13683,N_12184,N_13196);
xnor U13684 (N_13684,N_12181,N_12782);
or U13685 (N_13685,N_13224,N_12097);
nor U13686 (N_13686,N_12396,N_12075);
xnor U13687 (N_13687,N_12848,N_12703);
nor U13688 (N_13688,N_12521,N_12656);
xnor U13689 (N_13689,N_12161,N_12048);
nand U13690 (N_13690,N_13455,N_12989);
or U13691 (N_13691,N_13329,N_12705);
or U13692 (N_13692,N_13022,N_12662);
nand U13693 (N_13693,N_12971,N_12271);
nand U13694 (N_13694,N_12800,N_13422);
and U13695 (N_13695,N_12102,N_12765);
or U13696 (N_13696,N_12823,N_13491);
or U13697 (N_13697,N_12354,N_13209);
nor U13698 (N_13698,N_12833,N_12176);
or U13699 (N_13699,N_13068,N_12275);
nor U13700 (N_13700,N_12928,N_12071);
nand U13701 (N_13701,N_12193,N_12109);
xor U13702 (N_13702,N_12952,N_12562);
and U13703 (N_13703,N_12154,N_13485);
nand U13704 (N_13704,N_12660,N_12789);
or U13705 (N_13705,N_13493,N_13382);
xor U13706 (N_13706,N_12281,N_12011);
nor U13707 (N_13707,N_12336,N_13315);
nand U13708 (N_13708,N_12076,N_12895);
or U13709 (N_13709,N_13186,N_12995);
xor U13710 (N_13710,N_12513,N_12055);
nor U13711 (N_13711,N_13406,N_12718);
and U13712 (N_13712,N_12598,N_12536);
nand U13713 (N_13713,N_12448,N_13026);
and U13714 (N_13714,N_12204,N_12910);
nor U13715 (N_13715,N_12374,N_12959);
nor U13716 (N_13716,N_13071,N_13183);
xnor U13717 (N_13717,N_13145,N_12592);
nand U13718 (N_13718,N_12887,N_13409);
xnor U13719 (N_13719,N_13317,N_12816);
and U13720 (N_13720,N_12641,N_12213);
nand U13721 (N_13721,N_12468,N_12293);
and U13722 (N_13722,N_13280,N_13407);
nor U13723 (N_13723,N_13160,N_12023);
xor U13724 (N_13724,N_12801,N_12759);
and U13725 (N_13725,N_13169,N_12398);
nand U13726 (N_13726,N_13476,N_12635);
and U13727 (N_13727,N_13308,N_12886);
nand U13728 (N_13728,N_12926,N_13075);
nor U13729 (N_13729,N_13008,N_12761);
nor U13730 (N_13730,N_12830,N_12072);
nand U13731 (N_13731,N_12720,N_12670);
and U13732 (N_13732,N_12724,N_13459);
or U13733 (N_13733,N_12573,N_12601);
nand U13734 (N_13734,N_12351,N_12556);
or U13735 (N_13735,N_12177,N_13356);
or U13736 (N_13736,N_12480,N_12936);
or U13737 (N_13737,N_12729,N_12627);
and U13738 (N_13738,N_12727,N_13045);
nand U13739 (N_13739,N_12920,N_12577);
nand U13740 (N_13740,N_13402,N_12543);
and U13741 (N_13741,N_13200,N_12449);
nand U13742 (N_13742,N_12502,N_12825);
nand U13743 (N_13743,N_13037,N_12393);
nor U13744 (N_13744,N_13330,N_12459);
nand U13745 (N_13745,N_12067,N_12589);
nor U13746 (N_13746,N_12665,N_13130);
nand U13747 (N_13747,N_13416,N_12552);
nand U13748 (N_13748,N_12507,N_13393);
xor U13749 (N_13749,N_12743,N_12697);
nor U13750 (N_13750,N_12933,N_12571);
nor U13751 (N_13751,N_12322,N_12991);
xnor U13752 (N_13752,N_12802,N_13249);
nor U13753 (N_13753,N_13398,N_12050);
nor U13754 (N_13754,N_12325,N_13229);
nand U13755 (N_13755,N_12242,N_12430);
nand U13756 (N_13756,N_12005,N_12603);
or U13757 (N_13757,N_12438,N_13380);
xnor U13758 (N_13758,N_13175,N_12794);
and U13759 (N_13759,N_12286,N_13235);
and U13760 (N_13760,N_12814,N_12849);
and U13761 (N_13761,N_13199,N_12669);
xor U13762 (N_13762,N_13328,N_13440);
or U13763 (N_13763,N_13488,N_12241);
nand U13764 (N_13764,N_12546,N_12388);
xnor U13765 (N_13765,N_13208,N_12060);
or U13766 (N_13766,N_12062,N_13044);
or U13767 (N_13767,N_13291,N_12002);
or U13768 (N_13768,N_13219,N_13349);
xor U13769 (N_13769,N_13243,N_12725);
and U13770 (N_13770,N_13090,N_13373);
nand U13771 (N_13771,N_12856,N_13477);
nand U13772 (N_13772,N_12007,N_12614);
nor U13773 (N_13773,N_13094,N_12018);
nor U13774 (N_13774,N_12302,N_13312);
nand U13775 (N_13775,N_12975,N_12600);
and U13776 (N_13776,N_13341,N_12496);
xor U13777 (N_13777,N_12526,N_13079);
nand U13778 (N_13778,N_12239,N_13368);
nor U13779 (N_13779,N_12355,N_13048);
xnor U13780 (N_13780,N_12183,N_13489);
xnor U13781 (N_13781,N_12342,N_13379);
and U13782 (N_13782,N_12210,N_13171);
nand U13783 (N_13783,N_13129,N_12644);
and U13784 (N_13784,N_13246,N_12366);
xnor U13785 (N_13785,N_13304,N_12754);
xor U13786 (N_13786,N_13273,N_12708);
nor U13787 (N_13787,N_13103,N_12295);
xor U13788 (N_13788,N_12145,N_13056);
nand U13789 (N_13789,N_12940,N_13408);
nand U13790 (N_13790,N_12806,N_12677);
xnor U13791 (N_13791,N_13012,N_13092);
or U13792 (N_13792,N_13035,N_13230);
xor U13793 (N_13793,N_12303,N_12172);
nand U13794 (N_13794,N_13137,N_13089);
or U13795 (N_13795,N_12259,N_13324);
and U13796 (N_13796,N_13097,N_13117);
nor U13797 (N_13797,N_13143,N_12068);
nand U13798 (N_13798,N_12530,N_13187);
nor U13799 (N_13799,N_13126,N_12458);
xnor U13800 (N_13800,N_13162,N_12551);
and U13801 (N_13801,N_13015,N_12065);
and U13802 (N_13802,N_12238,N_12314);
nor U13803 (N_13803,N_12599,N_12017);
or U13804 (N_13804,N_12999,N_12752);
or U13805 (N_13805,N_12012,N_13337);
xnor U13806 (N_13806,N_12225,N_12315);
and U13807 (N_13807,N_13326,N_12569);
nand U13808 (N_13808,N_12538,N_12326);
nand U13809 (N_13809,N_13276,N_13076);
or U13810 (N_13810,N_13305,N_12146);
or U13811 (N_13811,N_12136,N_12107);
and U13812 (N_13812,N_12441,N_12896);
nor U13813 (N_13813,N_12861,N_12112);
or U13814 (N_13814,N_12415,N_12453);
nand U13815 (N_13815,N_12616,N_12832);
or U13816 (N_13816,N_12961,N_13483);
nand U13817 (N_13817,N_12508,N_13268);
and U13818 (N_13818,N_13084,N_12852);
or U13819 (N_13819,N_12709,N_13105);
nand U13820 (N_13820,N_12707,N_12371);
nand U13821 (N_13821,N_13149,N_13077);
or U13822 (N_13822,N_12568,N_12594);
and U13823 (N_13823,N_12228,N_13142);
and U13824 (N_13824,N_12248,N_12696);
xnor U13825 (N_13825,N_12411,N_12588);
or U13826 (N_13826,N_13391,N_12810);
or U13827 (N_13827,N_13179,N_12820);
or U13828 (N_13828,N_13167,N_12913);
and U13829 (N_13829,N_12333,N_13232);
nor U13830 (N_13830,N_12309,N_12437);
nor U13831 (N_13831,N_13420,N_12731);
or U13832 (N_13832,N_13340,N_12086);
xnor U13833 (N_13833,N_13458,N_13369);
and U13834 (N_13834,N_13333,N_13325);
nor U13835 (N_13835,N_12710,N_12996);
nand U13836 (N_13836,N_12767,N_12620);
nand U13837 (N_13837,N_13377,N_13194);
nand U13838 (N_13838,N_12025,N_12092);
or U13839 (N_13839,N_13424,N_12898);
nand U13840 (N_13840,N_13496,N_12844);
xor U13841 (N_13841,N_12706,N_12020);
nand U13842 (N_13842,N_12445,N_13417);
and U13843 (N_13843,N_12446,N_13462);
nand U13844 (N_13844,N_12983,N_12611);
xor U13845 (N_13845,N_13060,N_13113);
nand U13846 (N_13846,N_12240,N_13439);
and U13847 (N_13847,N_12838,N_12211);
xor U13848 (N_13848,N_13073,N_12111);
nor U13849 (N_13849,N_13394,N_12436);
nand U13850 (N_13850,N_12379,N_12386);
and U13851 (N_13851,N_12041,N_12046);
xor U13852 (N_13852,N_12473,N_13025);
or U13853 (N_13853,N_13441,N_12035);
nand U13854 (N_13854,N_12911,N_12661);
nand U13855 (N_13855,N_12308,N_12243);
xor U13856 (N_13856,N_12987,N_12391);
xnor U13857 (N_13857,N_12784,N_13131);
xnor U13858 (N_13858,N_12363,N_12909);
nand U13859 (N_13859,N_12916,N_12777);
nand U13860 (N_13860,N_12897,N_13461);
or U13861 (N_13861,N_12853,N_13498);
nor U13862 (N_13862,N_12486,N_12157);
nand U13863 (N_13863,N_12006,N_12298);
nand U13864 (N_13864,N_12528,N_13335);
nor U13865 (N_13865,N_12941,N_12866);
nor U13866 (N_13866,N_13109,N_12908);
nor U13867 (N_13867,N_12748,N_12701);
xor U13868 (N_13868,N_13467,N_13411);
nor U13869 (N_13869,N_12052,N_12793);
and U13870 (N_13870,N_12300,N_13070);
xnor U13871 (N_13871,N_12462,N_12403);
nor U13872 (N_13872,N_13132,N_12327);
or U13873 (N_13873,N_12285,N_12037);
or U13874 (N_13874,N_13495,N_12294);
or U13875 (N_13875,N_12216,N_13262);
and U13876 (N_13876,N_13147,N_12182);
nor U13877 (N_13877,N_13286,N_13497);
xor U13878 (N_13878,N_12778,N_13429);
nand U13879 (N_13879,N_13189,N_12095);
nor U13880 (N_13880,N_13404,N_13323);
and U13881 (N_13881,N_12253,N_12950);
nand U13882 (N_13882,N_12847,N_12501);
and U13883 (N_13883,N_12255,N_12760);
nor U13884 (N_13884,N_12657,N_12740);
nand U13885 (N_13885,N_12117,N_12345);
and U13886 (N_13886,N_12590,N_12755);
or U13887 (N_13887,N_13295,N_12137);
or U13888 (N_13888,N_12503,N_12431);
xnor U13889 (N_13889,N_12084,N_12713);
nand U13890 (N_13890,N_13365,N_12190);
nand U13891 (N_13891,N_12083,N_12716);
xor U13892 (N_13892,N_13448,N_12000);
nor U13893 (N_13893,N_13203,N_13086);
or U13894 (N_13894,N_12633,N_12498);
xor U13895 (N_13895,N_12385,N_12066);
nor U13896 (N_13896,N_12185,N_13239);
xor U13897 (N_13897,N_12639,N_12214);
nor U13898 (N_13898,N_12059,N_13301);
or U13899 (N_13899,N_12854,N_13395);
nand U13900 (N_13900,N_13193,N_13233);
and U13901 (N_13901,N_12014,N_12375);
nor U13902 (N_13902,N_13161,N_12198);
xnor U13903 (N_13903,N_12434,N_13138);
nor U13904 (N_13904,N_12087,N_12484);
and U13905 (N_13905,N_13252,N_12226);
xor U13906 (N_13906,N_12824,N_12632);
nor U13907 (N_13907,N_12489,N_13024);
and U13908 (N_13908,N_12232,N_12483);
or U13909 (N_13909,N_12572,N_12700);
and U13910 (N_13910,N_12746,N_13344);
xor U13911 (N_13911,N_12124,N_13298);
and U13912 (N_13912,N_12098,N_12619);
and U13913 (N_13913,N_12131,N_12547);
and U13914 (N_13914,N_12745,N_13492);
xnor U13915 (N_13915,N_13184,N_13053);
nor U13916 (N_13916,N_12931,N_13345);
and U13917 (N_13917,N_12469,N_12631);
nand U13918 (N_13918,N_12796,N_12420);
and U13919 (N_13919,N_12200,N_13009);
or U13920 (N_13920,N_13425,N_12116);
xnor U13921 (N_13921,N_13014,N_12283);
xnor U13922 (N_13922,N_12605,N_12405);
and U13923 (N_13923,N_13052,N_12889);
nor U13924 (N_13924,N_12610,N_13083);
or U13925 (N_13925,N_12094,N_13352);
nand U13926 (N_13926,N_12815,N_13401);
nor U13927 (N_13927,N_13100,N_12905);
nand U13928 (N_13928,N_12564,N_12134);
nand U13929 (N_13929,N_13334,N_12575);
or U13930 (N_13930,N_12369,N_12142);
xnor U13931 (N_13931,N_12034,N_12683);
and U13932 (N_13932,N_12851,N_12495);
xor U13933 (N_13933,N_12049,N_13346);
nor U13934 (N_13934,N_12121,N_12245);
or U13935 (N_13935,N_12811,N_12877);
or U13936 (N_13936,N_12362,N_13359);
nor U13937 (N_13937,N_13019,N_13111);
or U13938 (N_13938,N_12548,N_12147);
nor U13939 (N_13939,N_12763,N_12948);
and U13940 (N_13940,N_12428,N_12338);
or U13941 (N_13941,N_12681,N_12862);
and U13942 (N_13942,N_12402,N_13174);
or U13943 (N_13943,N_13363,N_13378);
and U13944 (N_13944,N_12969,N_12876);
nand U13945 (N_13945,N_12615,N_12160);
nand U13946 (N_13946,N_12756,N_12630);
nor U13947 (N_13947,N_13210,N_12888);
nor U13948 (N_13948,N_12165,N_13310);
nor U13949 (N_13949,N_12334,N_13222);
nor U13950 (N_13950,N_12015,N_13011);
and U13951 (N_13951,N_13080,N_12747);
xor U13952 (N_13952,N_13287,N_13135);
and U13953 (N_13953,N_12024,N_13003);
xor U13954 (N_13954,N_13041,N_13157);
and U13955 (N_13955,N_12977,N_12343);
nand U13956 (N_13956,N_12135,N_12349);
xor U13957 (N_13957,N_12026,N_12244);
nand U13958 (N_13958,N_12361,N_12927);
nor U13959 (N_13959,N_12118,N_13412);
and U13960 (N_13960,N_12212,N_13202);
or U13961 (N_13961,N_13336,N_12655);
nand U13962 (N_13962,N_12865,N_13125);
xnor U13963 (N_13963,N_12587,N_12788);
nor U13964 (N_13964,N_12762,N_12368);
nand U13965 (N_13965,N_12297,N_13120);
xor U13966 (N_13966,N_12642,N_13499);
or U13967 (N_13967,N_13220,N_12464);
or U13968 (N_13968,N_12267,N_12152);
nor U13969 (N_13969,N_12218,N_13248);
nor U13970 (N_13970,N_13453,N_13058);
or U13971 (N_13971,N_13212,N_12967);
xnor U13972 (N_13972,N_12175,N_12650);
and U13973 (N_13973,N_12772,N_12289);
nor U13974 (N_13974,N_12406,N_13443);
or U13975 (N_13975,N_12284,N_13098);
or U13976 (N_13976,N_13043,N_12553);
and U13977 (N_13977,N_12893,N_12923);
nor U13978 (N_13978,N_12695,N_12879);
nand U13979 (N_13979,N_12675,N_13279);
nor U13980 (N_13980,N_12409,N_12291);
and U13981 (N_13981,N_12429,N_12539);
or U13982 (N_13982,N_12252,N_12250);
nor U13983 (N_13983,N_12260,N_13180);
and U13984 (N_13984,N_12976,N_12389);
or U13985 (N_13985,N_12410,N_12939);
or U13986 (N_13986,N_12730,N_12230);
or U13987 (N_13987,N_13112,N_12381);
and U13988 (N_13988,N_12515,N_12395);
nor U13989 (N_13989,N_12043,N_12088);
nand U13990 (N_13990,N_13155,N_13091);
or U13991 (N_13991,N_13085,N_12753);
or U13992 (N_13992,N_12602,N_12280);
nand U13993 (N_13993,N_13264,N_12425);
xor U13994 (N_13994,N_12702,N_12869);
nand U13995 (N_13995,N_13236,N_12907);
nor U13996 (N_13996,N_12882,N_12475);
and U13997 (N_13997,N_13293,N_13151);
xnor U13998 (N_13998,N_12317,N_13063);
nand U13999 (N_13999,N_13118,N_12186);
and U14000 (N_14000,N_13221,N_13413);
xor U14001 (N_14001,N_12346,N_12937);
nand U14002 (N_14002,N_12456,N_12306);
xor U14003 (N_14003,N_12074,N_12634);
nor U14004 (N_14004,N_12359,N_12981);
or U14005 (N_14005,N_12554,N_12001);
nor U14006 (N_14006,N_13426,N_12776);
and U14007 (N_14007,N_13300,N_12580);
nor U14008 (N_14008,N_12105,N_12217);
nand U14009 (N_14009,N_13192,N_12545);
nand U14010 (N_14010,N_12826,N_12506);
and U14011 (N_14011,N_12257,N_13294);
nor U14012 (N_14012,N_13099,N_13469);
xnor U14013 (N_14013,N_12509,N_12953);
or U14014 (N_14014,N_12764,N_13327);
xor U14015 (N_14015,N_12412,N_13188);
and U14016 (N_14016,N_13134,N_13456);
and U14017 (N_14017,N_13283,N_12123);
and U14018 (N_14018,N_12679,N_12418);
nand U14019 (N_14019,N_12609,N_13272);
nand U14020 (N_14020,N_12842,N_12277);
xnor U14021 (N_14021,N_13478,N_12104);
nand U14022 (N_14022,N_12085,N_12504);
nor U14023 (N_14023,N_12045,N_12672);
nand U14024 (N_14024,N_12563,N_12561);
or U14025 (N_14025,N_12965,N_13415);
and U14026 (N_14026,N_12421,N_12472);
or U14027 (N_14027,N_12944,N_12819);
nor U14028 (N_14028,N_12586,N_12290);
nor U14029 (N_14029,N_12676,N_13081);
or U14030 (N_14030,N_13095,N_13050);
xnor U14031 (N_14031,N_13471,N_13256);
and U14032 (N_14032,N_13399,N_12978);
or U14033 (N_14033,N_12979,N_12652);
xnor U14034 (N_14034,N_13007,N_13215);
nor U14035 (N_14035,N_12082,N_13182);
or U14036 (N_14036,N_13023,N_13106);
nand U14037 (N_14037,N_12070,N_12906);
or U14038 (N_14038,N_12493,N_12320);
nand U14039 (N_14039,N_12519,N_12125);
nor U14040 (N_14040,N_12208,N_12273);
or U14041 (N_14041,N_12440,N_12884);
xor U14042 (N_14042,N_13472,N_13331);
and U14043 (N_14043,N_12864,N_12451);
nor U14044 (N_14044,N_12678,N_13072);
nor U14045 (N_14045,N_12324,N_12466);
and U14046 (N_14046,N_13389,N_12750);
or U14047 (N_14047,N_13270,N_12935);
nand U14048 (N_14048,N_12770,N_12974);
xnor U14049 (N_14049,N_13342,N_12691);
or U14050 (N_14050,N_12318,N_13387);
nand U14051 (N_14051,N_13154,N_12841);
or U14052 (N_14052,N_13254,N_12942);
nor U14053 (N_14053,N_13314,N_12444);
nand U14054 (N_14054,N_12056,N_13464);
nand U14055 (N_14055,N_13242,N_12194);
or U14056 (N_14056,N_12537,N_12269);
or U14057 (N_14057,N_12685,N_13449);
nor U14058 (N_14058,N_12766,N_12492);
nand U14059 (N_14059,N_12557,N_12168);
and U14060 (N_14060,N_12096,N_12057);
nand U14061 (N_14061,N_13253,N_13468);
or U14062 (N_14062,N_12039,N_12997);
or U14063 (N_14063,N_12054,N_12031);
and U14064 (N_14064,N_13364,N_12246);
and U14065 (N_14065,N_13392,N_12266);
nand U14066 (N_14066,N_13201,N_12254);
and U14067 (N_14067,N_13414,N_12090);
nand U14068 (N_14068,N_12424,N_12741);
xor U14069 (N_14069,N_12009,N_12607);
or U14070 (N_14070,N_12400,N_12487);
nand U14071 (N_14071,N_12150,N_13436);
nor U14072 (N_14072,N_12783,N_12968);
and U14073 (N_14073,N_12966,N_13059);
nand U14074 (N_14074,N_12311,N_12527);
and U14075 (N_14075,N_13228,N_12229);
or U14076 (N_14076,N_12938,N_12867);
and U14077 (N_14077,N_13437,N_12924);
nand U14078 (N_14078,N_12221,N_12510);
xor U14079 (N_14079,N_12954,N_12417);
xnor U14080 (N_14080,N_12608,N_12951);
nor U14081 (N_14081,N_12881,N_12917);
nand U14082 (N_14082,N_12499,N_12167);
nand U14083 (N_14083,N_12902,N_13303);
or U14084 (N_14084,N_12383,N_13166);
xor U14085 (N_14085,N_12078,N_13384);
nor U14086 (N_14086,N_12689,N_12699);
nor U14087 (N_14087,N_12233,N_13061);
or U14088 (N_14088,N_13197,N_12040);
or U14089 (N_14089,N_12101,N_12957);
or U14090 (N_14090,N_12169,N_12454);
nor U14091 (N_14091,N_12382,N_12376);
or U14092 (N_14092,N_13479,N_12235);
and U14093 (N_14093,N_12570,N_13066);
nor U14094 (N_14094,N_12597,N_13123);
nand U14095 (N_14095,N_13475,N_12042);
and U14096 (N_14096,N_12994,N_12875);
nand U14097 (N_14097,N_13322,N_12113);
nor U14098 (N_14098,N_12993,N_12945);
nor U14099 (N_14099,N_12894,N_12335);
and U14100 (N_14100,N_12667,N_13078);
xnor U14101 (N_14101,N_12612,N_12353);
nand U14102 (N_14102,N_12901,N_12148);
nand U14103 (N_14103,N_13207,N_12956);
or U14104 (N_14104,N_12164,N_13318);
nor U14105 (N_14105,N_13038,N_13274);
or U14106 (N_14106,N_13218,N_12439);
nand U14107 (N_14107,N_13140,N_12282);
nor U14108 (N_14108,N_13421,N_12549);
nand U14109 (N_14109,N_13482,N_12476);
or U14110 (N_14110,N_12693,N_12115);
or U14111 (N_14111,N_12943,N_12714);
nand U14112 (N_14112,N_13403,N_13353);
nand U14113 (N_14113,N_12191,N_13223);
nand U14114 (N_14114,N_12482,N_12809);
and U14115 (N_14115,N_12365,N_12535);
and U14116 (N_14116,N_13388,N_12621);
or U14117 (N_14117,N_12624,N_12870);
xnor U14118 (N_14118,N_12595,N_12036);
nor U14119 (N_14119,N_13321,N_12455);
xor U14120 (N_14120,N_12529,N_13348);
and U14121 (N_14121,N_13494,N_12721);
xor U14122 (N_14122,N_13177,N_12460);
nand U14123 (N_14123,N_12478,N_12964);
or U14124 (N_14124,N_12390,N_12900);
nor U14125 (N_14125,N_12033,N_12047);
and U14126 (N_14126,N_13266,N_13226);
nand U14127 (N_14127,N_12426,N_13153);
and U14128 (N_14128,N_12442,N_12955);
and U14129 (N_14129,N_13431,N_13238);
nand U14130 (N_14130,N_12202,N_12949);
nor U14131 (N_14131,N_12407,N_12144);
nand U14132 (N_14132,N_12972,N_12044);
nand U14133 (N_14133,N_12850,N_13372);
nor U14134 (N_14134,N_12733,N_12279);
and U14135 (N_14135,N_12596,N_13251);
nor U14136 (N_14136,N_13289,N_13258);
or U14137 (N_14137,N_12323,N_12179);
nand U14138 (N_14138,N_12008,N_13351);
and U14139 (N_14139,N_12272,N_13355);
or U14140 (N_14140,N_12717,N_12433);
nand U14141 (N_14141,N_12156,N_12514);
or U14142 (N_14142,N_12921,N_13240);
or U14143 (N_14143,N_12488,N_13000);
nand U14144 (N_14144,N_12485,N_13285);
or U14145 (N_14145,N_12196,N_13144);
or U14146 (N_14146,N_12004,N_12576);
and U14147 (N_14147,N_12348,N_12835);
or U14148 (N_14148,N_12474,N_13435);
xor U14149 (N_14149,N_12947,N_12582);
or U14150 (N_14150,N_12126,N_12812);
xor U14151 (N_14151,N_12958,N_13047);
and U14152 (N_14152,N_12132,N_12674);
and U14153 (N_14153,N_12435,N_12688);
nor U14154 (N_14154,N_12738,N_12903);
nand U14155 (N_14155,N_13309,N_12339);
nand U14156 (N_14156,N_13204,N_12626);
and U14157 (N_14157,N_12021,N_12653);
nand U14158 (N_14158,N_12885,N_12027);
xnor U14159 (N_14159,N_12629,N_13121);
or U14160 (N_14160,N_12030,N_12872);
nor U14161 (N_14161,N_13124,N_12982);
xnor U14162 (N_14162,N_13419,N_12742);
or U14163 (N_14163,N_12258,N_13225);
or U14164 (N_14164,N_12673,N_12158);
nand U14165 (N_14165,N_13146,N_12715);
and U14166 (N_14166,N_12032,N_12643);
and U14167 (N_14167,N_12122,N_12636);
and U14168 (N_14168,N_12199,N_13486);
nor U14169 (N_14169,N_12925,N_12970);
nor U14170 (N_14170,N_12313,N_12450);
and U14171 (N_14171,N_12684,N_12883);
nor U14172 (N_14172,N_12732,N_12319);
and U14173 (N_14173,N_13021,N_12378);
nand U14174 (N_14174,N_12531,N_13029);
and U14175 (N_14175,N_13290,N_12340);
nand U14176 (N_14176,N_12818,N_13010);
and U14177 (N_14177,N_13385,N_12874);
and U14178 (N_14178,N_12511,N_12370);
nor U14179 (N_14179,N_12091,N_13275);
xnor U14180 (N_14180,N_13093,N_13451);
nand U14181 (N_14181,N_12737,N_13339);
or U14182 (N_14182,N_12073,N_12822);
nand U14183 (N_14183,N_13292,N_12584);
and U14184 (N_14184,N_13343,N_13205);
nor U14185 (N_14185,N_13036,N_12288);
nand U14186 (N_14186,N_12350,N_12566);
nor U14187 (N_14187,N_13390,N_13457);
nand U14188 (N_14188,N_12491,N_13165);
nor U14189 (N_14189,N_12604,N_13168);
nor U14190 (N_14190,N_12163,N_13427);
or U14191 (N_14191,N_12394,N_13490);
nor U14192 (N_14192,N_12270,N_12757);
and U14193 (N_14193,N_13362,N_12479);
and U14194 (N_14194,N_12817,N_13159);
or U14195 (N_14195,N_12773,N_12863);
nor U14196 (N_14196,N_12840,N_13430);
or U14197 (N_14197,N_13306,N_13444);
or U14198 (N_14198,N_12465,N_12170);
or U14199 (N_14199,N_12775,N_12223);
and U14200 (N_14200,N_13042,N_13034);
or U14201 (N_14201,N_12637,N_12447);
nand U14202 (N_14202,N_13211,N_12384);
xor U14203 (N_14203,N_12332,N_13116);
or U14204 (N_14204,N_12792,N_13087);
xor U14205 (N_14205,N_12617,N_13297);
or U14206 (N_14206,N_12304,N_12099);
or U14207 (N_14207,N_12081,N_13338);
xnor U14208 (N_14208,N_12141,N_13119);
xor U14209 (N_14209,N_12682,N_13260);
nand U14210 (N_14210,N_13428,N_12985);
and U14211 (N_14211,N_12962,N_12079);
or U14212 (N_14212,N_12827,N_13316);
or U14213 (N_14213,N_12408,N_12986);
nor U14214 (N_14214,N_12834,N_12858);
nor U14215 (N_14215,N_12654,N_12622);
nor U14216 (N_14216,N_12392,N_12305);
and U14217 (N_14217,N_13213,N_13082);
or U14218 (N_14218,N_12443,N_13332);
and U14219 (N_14219,N_12795,N_12534);
nor U14220 (N_14220,N_12329,N_12963);
and U14221 (N_14221,N_12768,N_13383);
nor U14222 (N_14222,N_12836,N_13366);
nor U14223 (N_14223,N_13150,N_12671);
and U14224 (N_14224,N_13376,N_13282);
nor U14225 (N_14225,N_13354,N_12423);
nor U14226 (N_14226,N_12251,N_12219);
and U14227 (N_14227,N_13241,N_12891);
and U14228 (N_14228,N_12512,N_12728);
and U14229 (N_14229,N_12704,N_12058);
nor U14230 (N_14230,N_12069,N_12711);
and U14231 (N_14231,N_13445,N_13247);
nor U14232 (N_14232,N_12930,N_12769);
and U14233 (N_14233,N_12422,N_12490);
nand U14234 (N_14234,N_12645,N_13261);
nand U14235 (N_14235,N_12173,N_13466);
nand U14236 (N_14236,N_12330,N_12880);
nand U14237 (N_14237,N_13054,N_12739);
nor U14238 (N_14238,N_12278,N_12127);
xor U14239 (N_14239,N_12522,N_12133);
nor U14240 (N_14240,N_12264,N_12719);
and U14241 (N_14241,N_13452,N_12155);
nor U14242 (N_14242,N_12028,N_12919);
or U14243 (N_14243,N_12786,N_13237);
xor U14244 (N_14244,N_12470,N_12276);
and U14245 (N_14245,N_13040,N_12467);
nand U14246 (N_14246,N_12364,N_13139);
xor U14247 (N_14247,N_13375,N_12922);
and U14248 (N_14248,N_12347,N_12668);
xor U14249 (N_14249,N_13005,N_13487);
or U14250 (N_14250,N_13428,N_12701);
nor U14251 (N_14251,N_12281,N_12480);
nand U14252 (N_14252,N_13020,N_12751);
nand U14253 (N_14253,N_12476,N_12182);
nor U14254 (N_14254,N_12541,N_12927);
nand U14255 (N_14255,N_12308,N_12303);
nor U14256 (N_14256,N_12874,N_12076);
nor U14257 (N_14257,N_13436,N_13451);
xnor U14258 (N_14258,N_12586,N_13160);
and U14259 (N_14259,N_13428,N_13221);
nand U14260 (N_14260,N_12240,N_13230);
nand U14261 (N_14261,N_13197,N_13269);
xor U14262 (N_14262,N_12107,N_12910);
nor U14263 (N_14263,N_12140,N_12796);
or U14264 (N_14264,N_12087,N_12047);
nand U14265 (N_14265,N_13373,N_12603);
nor U14266 (N_14266,N_12831,N_12415);
xnor U14267 (N_14267,N_13460,N_13343);
and U14268 (N_14268,N_12038,N_12256);
nand U14269 (N_14269,N_12590,N_12295);
nor U14270 (N_14270,N_13492,N_12764);
nand U14271 (N_14271,N_12522,N_12059);
xnor U14272 (N_14272,N_13455,N_13004);
xnor U14273 (N_14273,N_13143,N_12671);
and U14274 (N_14274,N_12633,N_12877);
nor U14275 (N_14275,N_12190,N_13341);
nor U14276 (N_14276,N_13184,N_12714);
and U14277 (N_14277,N_12187,N_13280);
nor U14278 (N_14278,N_12715,N_12893);
nand U14279 (N_14279,N_12958,N_12497);
xor U14280 (N_14280,N_12123,N_12636);
or U14281 (N_14281,N_13266,N_12737);
xnor U14282 (N_14282,N_13470,N_12219);
and U14283 (N_14283,N_12661,N_12984);
xor U14284 (N_14284,N_12338,N_12765);
xor U14285 (N_14285,N_12314,N_12340);
and U14286 (N_14286,N_12339,N_12373);
nor U14287 (N_14287,N_12790,N_12134);
and U14288 (N_14288,N_12527,N_12552);
and U14289 (N_14289,N_12982,N_12657);
nand U14290 (N_14290,N_12238,N_12337);
nand U14291 (N_14291,N_13410,N_13294);
or U14292 (N_14292,N_12526,N_12493);
and U14293 (N_14293,N_12224,N_12664);
and U14294 (N_14294,N_13463,N_12645);
xor U14295 (N_14295,N_12403,N_13456);
xnor U14296 (N_14296,N_12600,N_12658);
nand U14297 (N_14297,N_13373,N_13001);
nand U14298 (N_14298,N_13180,N_12768);
and U14299 (N_14299,N_12184,N_12759);
nand U14300 (N_14300,N_12259,N_12039);
nand U14301 (N_14301,N_12460,N_12513);
nor U14302 (N_14302,N_13123,N_12836);
nand U14303 (N_14303,N_12966,N_13188);
or U14304 (N_14304,N_13406,N_13385);
and U14305 (N_14305,N_13170,N_12432);
nor U14306 (N_14306,N_12683,N_12897);
nor U14307 (N_14307,N_12643,N_13307);
or U14308 (N_14308,N_12118,N_12956);
nor U14309 (N_14309,N_12878,N_12723);
xnor U14310 (N_14310,N_12647,N_12369);
nor U14311 (N_14311,N_13213,N_12423);
xnor U14312 (N_14312,N_13459,N_12312);
or U14313 (N_14313,N_12339,N_12723);
or U14314 (N_14314,N_12539,N_13217);
nor U14315 (N_14315,N_13235,N_13332);
xnor U14316 (N_14316,N_12772,N_12354);
nor U14317 (N_14317,N_13343,N_12073);
or U14318 (N_14318,N_13208,N_12730);
or U14319 (N_14319,N_13027,N_12509);
nand U14320 (N_14320,N_12516,N_13372);
nor U14321 (N_14321,N_13284,N_12078);
nor U14322 (N_14322,N_12721,N_12562);
or U14323 (N_14323,N_12489,N_12710);
xor U14324 (N_14324,N_12175,N_13137);
nor U14325 (N_14325,N_12711,N_12339);
or U14326 (N_14326,N_12533,N_13278);
nand U14327 (N_14327,N_12645,N_12364);
or U14328 (N_14328,N_13269,N_12592);
or U14329 (N_14329,N_13089,N_12206);
and U14330 (N_14330,N_12191,N_12670);
xnor U14331 (N_14331,N_12454,N_12448);
and U14332 (N_14332,N_12148,N_12189);
xor U14333 (N_14333,N_13275,N_13100);
and U14334 (N_14334,N_13017,N_13091);
or U14335 (N_14335,N_13315,N_12036);
and U14336 (N_14336,N_13318,N_12231);
nor U14337 (N_14337,N_13497,N_12824);
or U14338 (N_14338,N_12849,N_12367);
nand U14339 (N_14339,N_12646,N_12161);
and U14340 (N_14340,N_12043,N_12040);
and U14341 (N_14341,N_13074,N_13134);
and U14342 (N_14342,N_12492,N_13019);
nand U14343 (N_14343,N_13087,N_12724);
xnor U14344 (N_14344,N_13083,N_12274);
nor U14345 (N_14345,N_13484,N_13315);
and U14346 (N_14346,N_13052,N_13376);
nor U14347 (N_14347,N_13114,N_12179);
nand U14348 (N_14348,N_12091,N_12260);
nor U14349 (N_14349,N_13250,N_12717);
nor U14350 (N_14350,N_12208,N_13132);
nor U14351 (N_14351,N_13025,N_12406);
nand U14352 (N_14352,N_12366,N_12986);
nor U14353 (N_14353,N_12211,N_12150);
or U14354 (N_14354,N_13021,N_12289);
nor U14355 (N_14355,N_12391,N_12864);
nor U14356 (N_14356,N_13244,N_12094);
or U14357 (N_14357,N_13064,N_13314);
nand U14358 (N_14358,N_12463,N_13395);
and U14359 (N_14359,N_12034,N_12106);
nand U14360 (N_14360,N_12548,N_12119);
and U14361 (N_14361,N_12719,N_12926);
xor U14362 (N_14362,N_12470,N_12973);
or U14363 (N_14363,N_13470,N_13148);
or U14364 (N_14364,N_12260,N_12859);
xnor U14365 (N_14365,N_12475,N_13233);
nor U14366 (N_14366,N_13432,N_12735);
nand U14367 (N_14367,N_12290,N_13051);
or U14368 (N_14368,N_12895,N_12805);
nand U14369 (N_14369,N_12021,N_13467);
nand U14370 (N_14370,N_13115,N_12647);
nor U14371 (N_14371,N_12385,N_13224);
nand U14372 (N_14372,N_12978,N_13110);
nand U14373 (N_14373,N_12933,N_12920);
and U14374 (N_14374,N_12268,N_12871);
nand U14375 (N_14375,N_13000,N_12820);
nor U14376 (N_14376,N_12600,N_12548);
and U14377 (N_14377,N_13180,N_12397);
xnor U14378 (N_14378,N_13430,N_13228);
nor U14379 (N_14379,N_13002,N_12156);
nand U14380 (N_14380,N_12131,N_12738);
or U14381 (N_14381,N_12202,N_12787);
xnor U14382 (N_14382,N_13131,N_12447);
and U14383 (N_14383,N_13284,N_13025);
xnor U14384 (N_14384,N_13321,N_13105);
or U14385 (N_14385,N_13239,N_13081);
or U14386 (N_14386,N_12810,N_12183);
nor U14387 (N_14387,N_12169,N_12045);
or U14388 (N_14388,N_13171,N_12081);
nor U14389 (N_14389,N_13327,N_13031);
xnor U14390 (N_14390,N_13450,N_12969);
nor U14391 (N_14391,N_12484,N_12670);
xnor U14392 (N_14392,N_12730,N_12798);
and U14393 (N_14393,N_12106,N_12629);
xnor U14394 (N_14394,N_12632,N_13337);
xnor U14395 (N_14395,N_12973,N_12307);
xor U14396 (N_14396,N_12403,N_13239);
xnor U14397 (N_14397,N_12508,N_12107);
nand U14398 (N_14398,N_12386,N_12990);
nand U14399 (N_14399,N_12964,N_12446);
nand U14400 (N_14400,N_12113,N_13267);
nor U14401 (N_14401,N_12504,N_12237);
nand U14402 (N_14402,N_12687,N_13098);
nor U14403 (N_14403,N_12058,N_13253);
xnor U14404 (N_14404,N_12804,N_13184);
xor U14405 (N_14405,N_12862,N_12653);
or U14406 (N_14406,N_12396,N_12832);
nand U14407 (N_14407,N_13004,N_12208);
and U14408 (N_14408,N_12547,N_13467);
nand U14409 (N_14409,N_12440,N_12112);
or U14410 (N_14410,N_12735,N_13340);
nor U14411 (N_14411,N_12870,N_12693);
nand U14412 (N_14412,N_12165,N_12094);
or U14413 (N_14413,N_13358,N_13212);
nor U14414 (N_14414,N_12024,N_13326);
nand U14415 (N_14415,N_12403,N_12169);
and U14416 (N_14416,N_12150,N_12595);
or U14417 (N_14417,N_12738,N_13136);
nor U14418 (N_14418,N_12555,N_12599);
xnor U14419 (N_14419,N_13463,N_13429);
nor U14420 (N_14420,N_13425,N_12044);
nor U14421 (N_14421,N_13446,N_12322);
nand U14422 (N_14422,N_12698,N_12349);
nand U14423 (N_14423,N_12292,N_12869);
xnor U14424 (N_14424,N_13324,N_12088);
xor U14425 (N_14425,N_12429,N_12356);
xnor U14426 (N_14426,N_12891,N_12571);
nand U14427 (N_14427,N_12541,N_12058);
and U14428 (N_14428,N_13038,N_12871);
and U14429 (N_14429,N_12077,N_12742);
nor U14430 (N_14430,N_12785,N_13386);
and U14431 (N_14431,N_12858,N_12006);
nand U14432 (N_14432,N_12652,N_12908);
or U14433 (N_14433,N_13043,N_12936);
and U14434 (N_14434,N_13067,N_12866);
or U14435 (N_14435,N_12652,N_13429);
nor U14436 (N_14436,N_12218,N_12792);
nand U14437 (N_14437,N_12732,N_12328);
nor U14438 (N_14438,N_12990,N_13383);
nor U14439 (N_14439,N_12520,N_12886);
nor U14440 (N_14440,N_12410,N_12882);
xor U14441 (N_14441,N_12900,N_13122);
nand U14442 (N_14442,N_12003,N_13455);
nor U14443 (N_14443,N_12506,N_12168);
nand U14444 (N_14444,N_12434,N_13366);
or U14445 (N_14445,N_13303,N_12827);
nor U14446 (N_14446,N_12590,N_12152);
nor U14447 (N_14447,N_12019,N_12150);
xor U14448 (N_14448,N_12392,N_13312);
nor U14449 (N_14449,N_12700,N_12411);
or U14450 (N_14450,N_12484,N_12406);
or U14451 (N_14451,N_12138,N_13167);
and U14452 (N_14452,N_12118,N_12536);
nor U14453 (N_14453,N_12487,N_12836);
nand U14454 (N_14454,N_13421,N_12265);
or U14455 (N_14455,N_12314,N_12792);
xor U14456 (N_14456,N_13140,N_13303);
nor U14457 (N_14457,N_12316,N_12480);
nor U14458 (N_14458,N_13412,N_12895);
or U14459 (N_14459,N_12011,N_13044);
xor U14460 (N_14460,N_13001,N_12212);
and U14461 (N_14461,N_12825,N_12856);
and U14462 (N_14462,N_12029,N_12907);
and U14463 (N_14463,N_12462,N_13402);
nor U14464 (N_14464,N_12783,N_12463);
or U14465 (N_14465,N_12480,N_12140);
nor U14466 (N_14466,N_12644,N_12110);
nand U14467 (N_14467,N_12239,N_13233);
and U14468 (N_14468,N_12153,N_13273);
nor U14469 (N_14469,N_12063,N_13247);
nor U14470 (N_14470,N_12279,N_13193);
and U14471 (N_14471,N_12926,N_13495);
and U14472 (N_14472,N_13013,N_12779);
nor U14473 (N_14473,N_12553,N_12176);
nor U14474 (N_14474,N_13497,N_12262);
nand U14475 (N_14475,N_13001,N_13187);
xnor U14476 (N_14476,N_12948,N_12040);
xor U14477 (N_14477,N_12936,N_12017);
xor U14478 (N_14478,N_13176,N_13188);
nor U14479 (N_14479,N_12610,N_13009);
nand U14480 (N_14480,N_12500,N_12147);
nand U14481 (N_14481,N_12675,N_12133);
or U14482 (N_14482,N_12046,N_12844);
nor U14483 (N_14483,N_12851,N_12525);
xnor U14484 (N_14484,N_12063,N_12758);
nor U14485 (N_14485,N_12328,N_12672);
xnor U14486 (N_14486,N_12132,N_12417);
xnor U14487 (N_14487,N_12071,N_13154);
nand U14488 (N_14488,N_13065,N_13292);
and U14489 (N_14489,N_12922,N_12959);
nor U14490 (N_14490,N_12793,N_12599);
xnor U14491 (N_14491,N_12250,N_12331);
nor U14492 (N_14492,N_12335,N_12246);
nand U14493 (N_14493,N_12841,N_12736);
xor U14494 (N_14494,N_12341,N_12549);
and U14495 (N_14495,N_12616,N_13234);
nand U14496 (N_14496,N_12769,N_12367);
xnor U14497 (N_14497,N_12798,N_12162);
nor U14498 (N_14498,N_13060,N_13394);
nor U14499 (N_14499,N_12698,N_12120);
or U14500 (N_14500,N_13316,N_13002);
xnor U14501 (N_14501,N_13267,N_13358);
nor U14502 (N_14502,N_12594,N_12595);
and U14503 (N_14503,N_12870,N_12888);
or U14504 (N_14504,N_12117,N_13274);
nand U14505 (N_14505,N_12882,N_12337);
xnor U14506 (N_14506,N_12989,N_12215);
and U14507 (N_14507,N_13069,N_12401);
nor U14508 (N_14508,N_12572,N_12337);
nor U14509 (N_14509,N_12885,N_13193);
and U14510 (N_14510,N_12932,N_12456);
and U14511 (N_14511,N_12951,N_13475);
xnor U14512 (N_14512,N_12704,N_13373);
or U14513 (N_14513,N_13242,N_12373);
or U14514 (N_14514,N_12354,N_12515);
xor U14515 (N_14515,N_13381,N_12885);
xor U14516 (N_14516,N_12482,N_12031);
nor U14517 (N_14517,N_13181,N_12285);
nor U14518 (N_14518,N_13482,N_12246);
xor U14519 (N_14519,N_12915,N_12032);
and U14520 (N_14520,N_13172,N_13295);
nand U14521 (N_14521,N_13094,N_12249);
or U14522 (N_14522,N_12865,N_12186);
nor U14523 (N_14523,N_12481,N_12002);
nor U14524 (N_14524,N_13038,N_12578);
nand U14525 (N_14525,N_12121,N_13059);
and U14526 (N_14526,N_12174,N_12895);
or U14527 (N_14527,N_12927,N_12412);
nand U14528 (N_14528,N_12520,N_12148);
nand U14529 (N_14529,N_13327,N_13077);
nor U14530 (N_14530,N_13280,N_13421);
and U14531 (N_14531,N_12759,N_12120);
xor U14532 (N_14532,N_12837,N_13246);
nand U14533 (N_14533,N_13448,N_12002);
nor U14534 (N_14534,N_12368,N_13362);
or U14535 (N_14535,N_12089,N_12873);
xnor U14536 (N_14536,N_13075,N_13121);
and U14537 (N_14537,N_13320,N_12349);
nor U14538 (N_14538,N_13034,N_12624);
and U14539 (N_14539,N_12030,N_12656);
nand U14540 (N_14540,N_12171,N_13191);
nand U14541 (N_14541,N_12379,N_12460);
or U14542 (N_14542,N_12273,N_12055);
and U14543 (N_14543,N_12469,N_13304);
xnor U14544 (N_14544,N_13437,N_12156);
or U14545 (N_14545,N_12810,N_12828);
nand U14546 (N_14546,N_13486,N_12158);
or U14547 (N_14547,N_12430,N_13191);
xor U14548 (N_14548,N_13456,N_12929);
nand U14549 (N_14549,N_12745,N_12100);
and U14550 (N_14550,N_12404,N_13305);
nand U14551 (N_14551,N_12255,N_12951);
or U14552 (N_14552,N_12970,N_13488);
and U14553 (N_14553,N_13079,N_13464);
and U14554 (N_14554,N_12546,N_12246);
xor U14555 (N_14555,N_12687,N_12193);
or U14556 (N_14556,N_13038,N_12492);
or U14557 (N_14557,N_13106,N_12468);
and U14558 (N_14558,N_12722,N_13411);
xor U14559 (N_14559,N_12479,N_13320);
nand U14560 (N_14560,N_12476,N_12905);
and U14561 (N_14561,N_12719,N_12104);
nand U14562 (N_14562,N_12901,N_13340);
and U14563 (N_14563,N_12390,N_13354);
and U14564 (N_14564,N_12033,N_12314);
nor U14565 (N_14565,N_12259,N_12817);
nand U14566 (N_14566,N_12880,N_13345);
nor U14567 (N_14567,N_12147,N_12143);
nor U14568 (N_14568,N_12740,N_12895);
and U14569 (N_14569,N_12426,N_12260);
and U14570 (N_14570,N_12452,N_12519);
or U14571 (N_14571,N_12643,N_12846);
nand U14572 (N_14572,N_12024,N_12450);
or U14573 (N_14573,N_12114,N_12211);
nor U14574 (N_14574,N_13140,N_13016);
or U14575 (N_14575,N_13048,N_13040);
or U14576 (N_14576,N_13044,N_13267);
or U14577 (N_14577,N_12102,N_13262);
or U14578 (N_14578,N_12575,N_12085);
or U14579 (N_14579,N_13181,N_12923);
or U14580 (N_14580,N_13134,N_12561);
or U14581 (N_14581,N_12837,N_12343);
nand U14582 (N_14582,N_12596,N_12194);
or U14583 (N_14583,N_12883,N_13051);
nand U14584 (N_14584,N_12429,N_13347);
xor U14585 (N_14585,N_13493,N_13491);
nand U14586 (N_14586,N_12290,N_12722);
or U14587 (N_14587,N_13266,N_12547);
and U14588 (N_14588,N_13445,N_13248);
or U14589 (N_14589,N_12450,N_13145);
xnor U14590 (N_14590,N_12679,N_12647);
nor U14591 (N_14591,N_12742,N_12707);
or U14592 (N_14592,N_13303,N_12861);
xnor U14593 (N_14593,N_12992,N_13348);
or U14594 (N_14594,N_12210,N_12715);
xor U14595 (N_14595,N_12603,N_13361);
nor U14596 (N_14596,N_12507,N_12863);
nand U14597 (N_14597,N_12997,N_12604);
nor U14598 (N_14598,N_13008,N_12544);
or U14599 (N_14599,N_13127,N_12869);
nor U14600 (N_14600,N_13296,N_12440);
xor U14601 (N_14601,N_12677,N_13337);
or U14602 (N_14602,N_12214,N_12763);
xor U14603 (N_14603,N_13049,N_12873);
xor U14604 (N_14604,N_12401,N_13236);
nand U14605 (N_14605,N_12916,N_12786);
nand U14606 (N_14606,N_12830,N_13426);
or U14607 (N_14607,N_13321,N_12312);
nor U14608 (N_14608,N_12792,N_12982);
xor U14609 (N_14609,N_12476,N_13355);
nor U14610 (N_14610,N_13349,N_12270);
nand U14611 (N_14611,N_13370,N_12076);
or U14612 (N_14612,N_12779,N_12703);
nor U14613 (N_14613,N_12426,N_13197);
nand U14614 (N_14614,N_13239,N_13410);
or U14615 (N_14615,N_13326,N_12562);
nand U14616 (N_14616,N_12168,N_12298);
and U14617 (N_14617,N_12755,N_13489);
or U14618 (N_14618,N_13363,N_12137);
xor U14619 (N_14619,N_12671,N_13385);
xnor U14620 (N_14620,N_13113,N_12887);
xor U14621 (N_14621,N_12655,N_12040);
and U14622 (N_14622,N_12448,N_13286);
or U14623 (N_14623,N_12486,N_13072);
nand U14624 (N_14624,N_13239,N_12544);
and U14625 (N_14625,N_13407,N_12580);
nor U14626 (N_14626,N_12757,N_13123);
and U14627 (N_14627,N_12582,N_13273);
nor U14628 (N_14628,N_12707,N_12141);
nor U14629 (N_14629,N_13032,N_12466);
or U14630 (N_14630,N_12516,N_12762);
xnor U14631 (N_14631,N_12036,N_12420);
xor U14632 (N_14632,N_12039,N_12281);
and U14633 (N_14633,N_13003,N_12702);
or U14634 (N_14634,N_12867,N_13074);
and U14635 (N_14635,N_12379,N_12117);
xor U14636 (N_14636,N_13127,N_12119);
xnor U14637 (N_14637,N_12072,N_12716);
nor U14638 (N_14638,N_12019,N_12136);
or U14639 (N_14639,N_13342,N_13373);
nor U14640 (N_14640,N_13013,N_12735);
nand U14641 (N_14641,N_13390,N_12814);
xnor U14642 (N_14642,N_12573,N_12602);
nand U14643 (N_14643,N_12851,N_13116);
nand U14644 (N_14644,N_12597,N_12537);
or U14645 (N_14645,N_13310,N_12256);
and U14646 (N_14646,N_13338,N_13198);
and U14647 (N_14647,N_12733,N_13373);
nor U14648 (N_14648,N_13196,N_12056);
xnor U14649 (N_14649,N_12699,N_12627);
or U14650 (N_14650,N_13353,N_13304);
xor U14651 (N_14651,N_13209,N_13426);
xnor U14652 (N_14652,N_13391,N_12987);
xor U14653 (N_14653,N_13183,N_12621);
or U14654 (N_14654,N_13236,N_13379);
xnor U14655 (N_14655,N_12610,N_13484);
nand U14656 (N_14656,N_12770,N_13249);
nor U14657 (N_14657,N_12164,N_12794);
or U14658 (N_14658,N_13336,N_13179);
and U14659 (N_14659,N_12886,N_12223);
or U14660 (N_14660,N_12451,N_13339);
nor U14661 (N_14661,N_13373,N_12054);
or U14662 (N_14662,N_13104,N_12382);
and U14663 (N_14663,N_13161,N_13252);
nand U14664 (N_14664,N_13265,N_12918);
nand U14665 (N_14665,N_13397,N_12051);
or U14666 (N_14666,N_13190,N_13087);
or U14667 (N_14667,N_12896,N_13128);
and U14668 (N_14668,N_12022,N_12080);
or U14669 (N_14669,N_12958,N_13333);
and U14670 (N_14670,N_12638,N_13049);
or U14671 (N_14671,N_12754,N_12053);
xor U14672 (N_14672,N_13331,N_12193);
or U14673 (N_14673,N_12305,N_12855);
or U14674 (N_14674,N_12866,N_12293);
or U14675 (N_14675,N_12384,N_12615);
nor U14676 (N_14676,N_12270,N_12335);
nor U14677 (N_14677,N_13298,N_12553);
or U14678 (N_14678,N_12777,N_12910);
nor U14679 (N_14679,N_13490,N_12423);
and U14680 (N_14680,N_12080,N_13147);
nor U14681 (N_14681,N_12546,N_13197);
nand U14682 (N_14682,N_13063,N_12977);
and U14683 (N_14683,N_13020,N_12102);
xor U14684 (N_14684,N_13283,N_13360);
xnor U14685 (N_14685,N_13009,N_13357);
and U14686 (N_14686,N_12291,N_12403);
or U14687 (N_14687,N_13069,N_13480);
and U14688 (N_14688,N_13107,N_12973);
or U14689 (N_14689,N_12449,N_12701);
and U14690 (N_14690,N_13487,N_12823);
nand U14691 (N_14691,N_12603,N_12523);
nor U14692 (N_14692,N_12539,N_12245);
nor U14693 (N_14693,N_12632,N_12213);
or U14694 (N_14694,N_12729,N_12388);
nand U14695 (N_14695,N_12257,N_13093);
nand U14696 (N_14696,N_13117,N_12537);
xnor U14697 (N_14697,N_12686,N_12954);
or U14698 (N_14698,N_12153,N_12684);
xnor U14699 (N_14699,N_13069,N_12545);
and U14700 (N_14700,N_12799,N_13495);
nor U14701 (N_14701,N_13410,N_12368);
nand U14702 (N_14702,N_12126,N_12461);
or U14703 (N_14703,N_12550,N_12797);
and U14704 (N_14704,N_12271,N_12114);
nand U14705 (N_14705,N_12167,N_12826);
or U14706 (N_14706,N_12679,N_13130);
and U14707 (N_14707,N_13366,N_12583);
nand U14708 (N_14708,N_12163,N_12831);
xnor U14709 (N_14709,N_12763,N_12189);
xor U14710 (N_14710,N_12482,N_12565);
nand U14711 (N_14711,N_13183,N_12146);
xor U14712 (N_14712,N_12354,N_12881);
and U14713 (N_14713,N_12073,N_13413);
nand U14714 (N_14714,N_12162,N_12024);
xor U14715 (N_14715,N_12567,N_12501);
nand U14716 (N_14716,N_12125,N_13400);
nor U14717 (N_14717,N_12227,N_12393);
nor U14718 (N_14718,N_13243,N_13439);
xnor U14719 (N_14719,N_12442,N_12026);
xnor U14720 (N_14720,N_13377,N_12054);
nor U14721 (N_14721,N_13247,N_12369);
nand U14722 (N_14722,N_13187,N_12730);
nand U14723 (N_14723,N_13331,N_12557);
xor U14724 (N_14724,N_12223,N_13299);
or U14725 (N_14725,N_13370,N_12208);
xnor U14726 (N_14726,N_12470,N_13038);
and U14727 (N_14727,N_12695,N_13406);
nand U14728 (N_14728,N_12340,N_13412);
or U14729 (N_14729,N_12754,N_12700);
xor U14730 (N_14730,N_12667,N_12045);
or U14731 (N_14731,N_13249,N_13043);
nor U14732 (N_14732,N_12661,N_12652);
nand U14733 (N_14733,N_12614,N_13474);
nor U14734 (N_14734,N_12385,N_13099);
xor U14735 (N_14735,N_13056,N_12841);
nor U14736 (N_14736,N_13397,N_13220);
xor U14737 (N_14737,N_12094,N_13175);
or U14738 (N_14738,N_13256,N_12876);
nand U14739 (N_14739,N_12403,N_12370);
xor U14740 (N_14740,N_12340,N_12050);
or U14741 (N_14741,N_12214,N_12086);
nand U14742 (N_14742,N_12849,N_12389);
xor U14743 (N_14743,N_12468,N_13390);
nor U14744 (N_14744,N_12926,N_13066);
or U14745 (N_14745,N_12413,N_12718);
and U14746 (N_14746,N_12611,N_12168);
or U14747 (N_14747,N_12479,N_12428);
xnor U14748 (N_14748,N_12691,N_12491);
and U14749 (N_14749,N_13136,N_13015);
xor U14750 (N_14750,N_12772,N_13130);
nand U14751 (N_14751,N_13304,N_13166);
nand U14752 (N_14752,N_12884,N_12438);
xor U14753 (N_14753,N_12618,N_12555);
nor U14754 (N_14754,N_12151,N_12168);
nand U14755 (N_14755,N_13035,N_12083);
xnor U14756 (N_14756,N_13246,N_12265);
nor U14757 (N_14757,N_12439,N_12414);
or U14758 (N_14758,N_13191,N_12052);
nand U14759 (N_14759,N_13248,N_12992);
or U14760 (N_14760,N_12779,N_13088);
and U14761 (N_14761,N_12282,N_12023);
nand U14762 (N_14762,N_12422,N_12479);
xnor U14763 (N_14763,N_12497,N_13050);
and U14764 (N_14764,N_12321,N_13033);
and U14765 (N_14765,N_12963,N_12883);
or U14766 (N_14766,N_12653,N_13353);
and U14767 (N_14767,N_12151,N_13213);
nand U14768 (N_14768,N_13153,N_13380);
xnor U14769 (N_14769,N_13195,N_12224);
nand U14770 (N_14770,N_13173,N_12794);
nor U14771 (N_14771,N_12178,N_13166);
nand U14772 (N_14772,N_12552,N_12145);
or U14773 (N_14773,N_12272,N_12008);
and U14774 (N_14774,N_13366,N_12798);
nand U14775 (N_14775,N_12151,N_12244);
xor U14776 (N_14776,N_13027,N_12293);
nand U14777 (N_14777,N_12821,N_12823);
nand U14778 (N_14778,N_12555,N_12460);
nand U14779 (N_14779,N_12431,N_12248);
or U14780 (N_14780,N_13172,N_12203);
nand U14781 (N_14781,N_13282,N_12995);
xnor U14782 (N_14782,N_12438,N_12718);
and U14783 (N_14783,N_12733,N_12375);
xor U14784 (N_14784,N_13301,N_13212);
xor U14785 (N_14785,N_13139,N_13138);
xnor U14786 (N_14786,N_12592,N_13318);
nor U14787 (N_14787,N_12019,N_12738);
or U14788 (N_14788,N_12038,N_12815);
and U14789 (N_14789,N_12886,N_12586);
xnor U14790 (N_14790,N_13034,N_12497);
or U14791 (N_14791,N_12961,N_13017);
nor U14792 (N_14792,N_13290,N_12021);
and U14793 (N_14793,N_12837,N_12049);
and U14794 (N_14794,N_12330,N_12943);
nor U14795 (N_14795,N_12202,N_12518);
nor U14796 (N_14796,N_12223,N_12113);
nor U14797 (N_14797,N_12622,N_12639);
nor U14798 (N_14798,N_12318,N_13220);
or U14799 (N_14799,N_12247,N_12117);
or U14800 (N_14800,N_12485,N_13243);
nand U14801 (N_14801,N_13153,N_13174);
nand U14802 (N_14802,N_12652,N_12157);
and U14803 (N_14803,N_12079,N_12527);
and U14804 (N_14804,N_13474,N_13081);
nand U14805 (N_14805,N_12130,N_12880);
and U14806 (N_14806,N_13348,N_13294);
or U14807 (N_14807,N_12878,N_13261);
nand U14808 (N_14808,N_12325,N_12662);
nor U14809 (N_14809,N_13409,N_13192);
nor U14810 (N_14810,N_12473,N_13484);
xnor U14811 (N_14811,N_12096,N_13011);
and U14812 (N_14812,N_12247,N_12041);
or U14813 (N_14813,N_13489,N_13120);
nor U14814 (N_14814,N_13245,N_13243);
xor U14815 (N_14815,N_12197,N_13219);
xor U14816 (N_14816,N_13212,N_12433);
nor U14817 (N_14817,N_12163,N_12010);
nand U14818 (N_14818,N_13259,N_12669);
or U14819 (N_14819,N_13278,N_12401);
nor U14820 (N_14820,N_12713,N_12217);
or U14821 (N_14821,N_12757,N_12303);
and U14822 (N_14822,N_13188,N_12479);
and U14823 (N_14823,N_12960,N_13371);
and U14824 (N_14824,N_13304,N_12836);
or U14825 (N_14825,N_12268,N_12100);
xnor U14826 (N_14826,N_13034,N_13207);
and U14827 (N_14827,N_13371,N_13336);
xor U14828 (N_14828,N_13437,N_12084);
or U14829 (N_14829,N_13035,N_12133);
nand U14830 (N_14830,N_12690,N_13494);
nor U14831 (N_14831,N_13491,N_12316);
xor U14832 (N_14832,N_12048,N_13341);
or U14833 (N_14833,N_12516,N_13147);
xnor U14834 (N_14834,N_12569,N_13057);
nand U14835 (N_14835,N_13001,N_13109);
nand U14836 (N_14836,N_13317,N_12956);
nand U14837 (N_14837,N_12790,N_12144);
nand U14838 (N_14838,N_12881,N_12230);
or U14839 (N_14839,N_13441,N_12388);
and U14840 (N_14840,N_12705,N_12200);
nor U14841 (N_14841,N_12612,N_12582);
nor U14842 (N_14842,N_12746,N_12390);
nand U14843 (N_14843,N_12555,N_13149);
and U14844 (N_14844,N_12744,N_12071);
or U14845 (N_14845,N_12500,N_13030);
or U14846 (N_14846,N_13193,N_12126);
xor U14847 (N_14847,N_12139,N_12026);
and U14848 (N_14848,N_13083,N_12289);
nand U14849 (N_14849,N_13127,N_12985);
nor U14850 (N_14850,N_12811,N_12866);
xnor U14851 (N_14851,N_13156,N_13195);
xor U14852 (N_14852,N_13234,N_13370);
nor U14853 (N_14853,N_12097,N_12250);
xnor U14854 (N_14854,N_12143,N_12463);
nand U14855 (N_14855,N_12810,N_12940);
or U14856 (N_14856,N_12263,N_12881);
nand U14857 (N_14857,N_13332,N_12127);
xor U14858 (N_14858,N_12323,N_12549);
nand U14859 (N_14859,N_12223,N_13281);
or U14860 (N_14860,N_12907,N_12851);
and U14861 (N_14861,N_12305,N_13031);
nand U14862 (N_14862,N_13023,N_13377);
and U14863 (N_14863,N_13430,N_13487);
nor U14864 (N_14864,N_13152,N_13397);
xnor U14865 (N_14865,N_13083,N_12373);
and U14866 (N_14866,N_12670,N_13253);
and U14867 (N_14867,N_12430,N_12924);
or U14868 (N_14868,N_12823,N_13432);
or U14869 (N_14869,N_12016,N_13139);
and U14870 (N_14870,N_12944,N_12748);
and U14871 (N_14871,N_12632,N_12845);
nor U14872 (N_14872,N_12683,N_13307);
and U14873 (N_14873,N_12903,N_13374);
nor U14874 (N_14874,N_12935,N_13354);
xor U14875 (N_14875,N_12837,N_12392);
xor U14876 (N_14876,N_12057,N_13427);
or U14877 (N_14877,N_12277,N_12364);
or U14878 (N_14878,N_12258,N_12701);
nor U14879 (N_14879,N_12328,N_13444);
nor U14880 (N_14880,N_12976,N_12282);
nor U14881 (N_14881,N_12051,N_12060);
nand U14882 (N_14882,N_12746,N_13478);
nor U14883 (N_14883,N_13258,N_12725);
or U14884 (N_14884,N_12571,N_12616);
and U14885 (N_14885,N_13108,N_13380);
xnor U14886 (N_14886,N_12243,N_12412);
nor U14887 (N_14887,N_12077,N_12627);
xor U14888 (N_14888,N_12887,N_13207);
and U14889 (N_14889,N_13188,N_12440);
and U14890 (N_14890,N_12467,N_12179);
and U14891 (N_14891,N_13177,N_13184);
xnor U14892 (N_14892,N_13400,N_12980);
nand U14893 (N_14893,N_12899,N_12481);
and U14894 (N_14894,N_13120,N_12652);
and U14895 (N_14895,N_12964,N_13336);
nor U14896 (N_14896,N_13093,N_13284);
nor U14897 (N_14897,N_13492,N_13434);
xnor U14898 (N_14898,N_12820,N_12805);
and U14899 (N_14899,N_12635,N_12244);
nand U14900 (N_14900,N_12000,N_12959);
nor U14901 (N_14901,N_12682,N_12804);
nand U14902 (N_14902,N_13341,N_12026);
xor U14903 (N_14903,N_12951,N_13369);
and U14904 (N_14904,N_13441,N_12311);
or U14905 (N_14905,N_12432,N_12702);
or U14906 (N_14906,N_12851,N_12651);
nor U14907 (N_14907,N_12151,N_13137);
xnor U14908 (N_14908,N_13166,N_13066);
or U14909 (N_14909,N_13425,N_13289);
xor U14910 (N_14910,N_13060,N_12684);
and U14911 (N_14911,N_12932,N_12591);
nor U14912 (N_14912,N_13445,N_13411);
nor U14913 (N_14913,N_12426,N_12968);
nand U14914 (N_14914,N_13435,N_12249);
nor U14915 (N_14915,N_13452,N_13357);
nand U14916 (N_14916,N_12170,N_13493);
xnor U14917 (N_14917,N_12834,N_12034);
or U14918 (N_14918,N_12260,N_12858);
nor U14919 (N_14919,N_12625,N_12572);
xor U14920 (N_14920,N_12932,N_12253);
and U14921 (N_14921,N_13111,N_12985);
and U14922 (N_14922,N_12824,N_12221);
or U14923 (N_14923,N_12980,N_12669);
nand U14924 (N_14924,N_13275,N_12894);
or U14925 (N_14925,N_13285,N_12407);
xnor U14926 (N_14926,N_12238,N_12415);
and U14927 (N_14927,N_13439,N_13184);
nand U14928 (N_14928,N_13359,N_12200);
nor U14929 (N_14929,N_13129,N_13375);
and U14930 (N_14930,N_12275,N_12825);
or U14931 (N_14931,N_12763,N_12057);
nand U14932 (N_14932,N_12919,N_13122);
nand U14933 (N_14933,N_12380,N_12943);
xor U14934 (N_14934,N_13217,N_13171);
nand U14935 (N_14935,N_12524,N_12337);
or U14936 (N_14936,N_12220,N_13223);
nand U14937 (N_14937,N_13171,N_13373);
nor U14938 (N_14938,N_12743,N_13191);
or U14939 (N_14939,N_12550,N_12476);
and U14940 (N_14940,N_12643,N_13147);
and U14941 (N_14941,N_12085,N_12660);
and U14942 (N_14942,N_13180,N_13169);
nand U14943 (N_14943,N_13380,N_12111);
xor U14944 (N_14944,N_12096,N_13158);
nor U14945 (N_14945,N_12666,N_13447);
and U14946 (N_14946,N_12646,N_12028);
and U14947 (N_14947,N_13044,N_12114);
or U14948 (N_14948,N_12060,N_12497);
xor U14949 (N_14949,N_12618,N_12904);
and U14950 (N_14950,N_12773,N_13059);
or U14951 (N_14951,N_13470,N_12797);
nor U14952 (N_14952,N_12930,N_13110);
and U14953 (N_14953,N_12843,N_13041);
or U14954 (N_14954,N_13214,N_12171);
or U14955 (N_14955,N_12929,N_12080);
nor U14956 (N_14956,N_13186,N_12967);
and U14957 (N_14957,N_12024,N_13296);
nand U14958 (N_14958,N_13358,N_13447);
xor U14959 (N_14959,N_12131,N_12210);
and U14960 (N_14960,N_12774,N_12146);
and U14961 (N_14961,N_12196,N_13331);
xor U14962 (N_14962,N_12134,N_12737);
and U14963 (N_14963,N_13364,N_12342);
or U14964 (N_14964,N_13420,N_13173);
and U14965 (N_14965,N_12758,N_13291);
xnor U14966 (N_14966,N_13323,N_12714);
and U14967 (N_14967,N_13193,N_12037);
nor U14968 (N_14968,N_12443,N_12470);
and U14969 (N_14969,N_12921,N_12421);
or U14970 (N_14970,N_12637,N_12686);
or U14971 (N_14971,N_12335,N_12143);
nand U14972 (N_14972,N_12663,N_13327);
nor U14973 (N_14973,N_12926,N_13361);
nand U14974 (N_14974,N_12779,N_13225);
or U14975 (N_14975,N_13346,N_12500);
nand U14976 (N_14976,N_13039,N_12429);
xor U14977 (N_14977,N_12500,N_12076);
or U14978 (N_14978,N_12911,N_13444);
xor U14979 (N_14979,N_13406,N_12152);
nand U14980 (N_14980,N_12769,N_12911);
nand U14981 (N_14981,N_12532,N_12335);
xor U14982 (N_14982,N_12920,N_12948);
xor U14983 (N_14983,N_12837,N_12528);
nor U14984 (N_14984,N_12850,N_12047);
and U14985 (N_14985,N_12077,N_12483);
nor U14986 (N_14986,N_12196,N_12669);
xnor U14987 (N_14987,N_12092,N_12308);
or U14988 (N_14988,N_13371,N_13487);
xor U14989 (N_14989,N_13171,N_12705);
and U14990 (N_14990,N_12811,N_12119);
and U14991 (N_14991,N_12033,N_13060);
and U14992 (N_14992,N_12095,N_12957);
nor U14993 (N_14993,N_13107,N_13071);
or U14994 (N_14994,N_12515,N_12508);
or U14995 (N_14995,N_12764,N_12968);
or U14996 (N_14996,N_12586,N_12406);
and U14997 (N_14997,N_13398,N_13487);
nand U14998 (N_14998,N_13471,N_12483);
and U14999 (N_14999,N_13176,N_13187);
and UO_0 (O_0,N_13577,N_14496);
nand UO_1 (O_1,N_14346,N_14748);
nor UO_2 (O_2,N_14480,N_14033);
xnor UO_3 (O_3,N_14546,N_13591);
or UO_4 (O_4,N_14556,N_13961);
or UO_5 (O_5,N_14025,N_14693);
nor UO_6 (O_6,N_13754,N_14407);
nor UO_7 (O_7,N_13699,N_14666);
nand UO_8 (O_8,N_14517,N_14635);
and UO_9 (O_9,N_14044,N_14211);
and UO_10 (O_10,N_13599,N_13804);
or UO_11 (O_11,N_13942,N_13751);
xor UO_12 (O_12,N_14684,N_14854);
nor UO_13 (O_13,N_13904,N_13932);
xor UO_14 (O_14,N_13730,N_13877);
nand UO_15 (O_15,N_14241,N_14552);
and UO_16 (O_16,N_14973,N_14197);
nand UO_17 (O_17,N_13564,N_14622);
or UO_18 (O_18,N_14958,N_13663);
nor UO_19 (O_19,N_13802,N_14607);
xor UO_20 (O_20,N_13869,N_14390);
nor UO_21 (O_21,N_14833,N_14419);
or UO_22 (O_22,N_14555,N_14589);
or UO_23 (O_23,N_14142,N_13623);
and UO_24 (O_24,N_14041,N_14002);
nor UO_25 (O_25,N_14271,N_13974);
and UO_26 (O_26,N_14260,N_14006);
nand UO_27 (O_27,N_14929,N_14987);
and UO_28 (O_28,N_14813,N_14152);
and UO_29 (O_29,N_14986,N_14526);
xnor UO_30 (O_30,N_13905,N_14367);
and UO_31 (O_31,N_14151,N_14083);
xnor UO_32 (O_32,N_14847,N_14918);
and UO_33 (O_33,N_14363,N_14273);
nor UO_34 (O_34,N_13921,N_13502);
xnor UO_35 (O_35,N_13722,N_13925);
or UO_36 (O_36,N_14160,N_14902);
nor UO_37 (O_37,N_13727,N_14643);
nand UO_38 (O_38,N_14500,N_14722);
xnor UO_39 (O_39,N_14647,N_14482);
nand UO_40 (O_40,N_14043,N_14539);
nand UO_41 (O_41,N_14942,N_14625);
nor UO_42 (O_42,N_14699,N_13855);
or UO_43 (O_43,N_14711,N_14889);
nand UO_44 (O_44,N_14992,N_14375);
nand UO_45 (O_45,N_14327,N_13538);
nand UO_46 (O_46,N_14239,N_14365);
nor UO_47 (O_47,N_13648,N_14948);
xnor UO_48 (O_48,N_14282,N_13620);
or UO_49 (O_49,N_14131,N_13989);
nor UO_50 (O_50,N_14434,N_13830);
or UO_51 (O_51,N_14134,N_14921);
nand UO_52 (O_52,N_14513,N_14337);
or UO_53 (O_53,N_14310,N_13840);
or UO_54 (O_54,N_14528,N_14771);
xnor UO_55 (O_55,N_14252,N_14793);
xnor UO_56 (O_56,N_14183,N_14287);
and UO_57 (O_57,N_14386,N_14398);
nand UO_58 (O_58,N_13927,N_13769);
xnor UO_59 (O_59,N_13595,N_13934);
or UO_60 (O_60,N_13805,N_13558);
or UO_61 (O_61,N_14175,N_14069);
xnor UO_62 (O_62,N_14537,N_14877);
xnor UO_63 (O_63,N_13531,N_14037);
nand UO_64 (O_64,N_14976,N_14609);
or UO_65 (O_65,N_14218,N_14614);
and UO_66 (O_66,N_14162,N_14723);
xnor UO_67 (O_67,N_14068,N_13887);
nor UO_68 (O_68,N_13966,N_14270);
nor UO_69 (O_69,N_13860,N_14011);
xor UO_70 (O_70,N_14411,N_14096);
nand UO_71 (O_71,N_14313,N_14053);
nor UO_72 (O_72,N_14495,N_14220);
nand UO_73 (O_73,N_14424,N_14455);
xor UO_74 (O_74,N_13570,N_13912);
nor UO_75 (O_75,N_14339,N_14501);
nand UO_76 (O_76,N_14472,N_14089);
or UO_77 (O_77,N_13549,N_14538);
nor UO_78 (O_78,N_14626,N_14954);
and UO_79 (O_79,N_13718,N_14357);
xor UO_80 (O_80,N_13811,N_14791);
or UO_81 (O_81,N_14493,N_14226);
xor UO_82 (O_82,N_14276,N_13796);
nor UO_83 (O_83,N_14499,N_13775);
nor UO_84 (O_84,N_13627,N_13878);
nand UO_85 (O_85,N_14952,N_14412);
xor UO_86 (O_86,N_13828,N_14901);
nor UO_87 (O_87,N_14021,N_13682);
xnor UO_88 (O_88,N_14176,N_14370);
nand UO_89 (O_89,N_13884,N_14989);
or UO_90 (O_90,N_14497,N_14628);
or UO_91 (O_91,N_13504,N_14384);
nand UO_92 (O_92,N_14117,N_14303);
or UO_93 (O_93,N_13615,N_14332);
nor UO_94 (O_94,N_14017,N_14395);
nand UO_95 (O_95,N_13689,N_13665);
nand UO_96 (O_96,N_14124,N_14503);
xor UO_97 (O_97,N_14143,N_14478);
nor UO_98 (O_98,N_13528,N_14839);
nand UO_99 (O_99,N_14167,N_14560);
and UO_100 (O_100,N_14894,N_14979);
xor UO_101 (O_101,N_13894,N_13752);
xnor UO_102 (O_102,N_14893,N_13915);
and UO_103 (O_103,N_13953,N_13816);
nand UO_104 (O_104,N_13848,N_13794);
nand UO_105 (O_105,N_14774,N_14009);
xnor UO_106 (O_106,N_14476,N_14878);
and UO_107 (O_107,N_13960,N_14272);
or UO_108 (O_108,N_14563,N_14810);
and UO_109 (O_109,N_13566,N_14072);
xnor UO_110 (O_110,N_14757,N_14524);
or UO_111 (O_111,N_14465,N_14646);
nand UO_112 (O_112,N_13909,N_13980);
and UO_113 (O_113,N_13712,N_14030);
xnor UO_114 (O_114,N_13574,N_13922);
and UO_115 (O_115,N_13986,N_14582);
or UO_116 (O_116,N_14199,N_13500);
nor UO_117 (O_117,N_14330,N_13736);
or UO_118 (O_118,N_14277,N_13862);
nor UO_119 (O_119,N_13889,N_13814);
and UO_120 (O_120,N_13747,N_13834);
nand UO_121 (O_121,N_14026,N_14462);
or UO_122 (O_122,N_13990,N_13851);
nor UO_123 (O_123,N_14435,N_14071);
xor UO_124 (O_124,N_14566,N_14809);
nand UO_125 (O_125,N_13971,N_14007);
nand UO_126 (O_126,N_13749,N_14688);
nor UO_127 (O_127,N_14518,N_14221);
nand UO_128 (O_128,N_14141,N_13755);
or UO_129 (O_129,N_14704,N_13725);
nor UO_130 (O_130,N_13935,N_13688);
nor UO_131 (O_131,N_14819,N_13801);
and UO_132 (O_132,N_13588,N_14772);
or UO_133 (O_133,N_14597,N_13969);
or UO_134 (O_134,N_14746,N_14323);
and UO_135 (O_135,N_13673,N_13907);
nor UO_136 (O_136,N_14803,N_13544);
nor UO_137 (O_137,N_13982,N_14415);
nand UO_138 (O_138,N_13707,N_14629);
nand UO_139 (O_139,N_14144,N_14615);
nor UO_140 (O_140,N_13957,N_14898);
xor UO_141 (O_141,N_14210,N_14256);
or UO_142 (O_142,N_14737,N_14967);
and UO_143 (O_143,N_14110,N_13853);
xor UO_144 (O_144,N_13680,N_13551);
xor UO_145 (O_145,N_14799,N_14639);
or UO_146 (O_146,N_14675,N_14316);
nor UO_147 (O_147,N_13917,N_14579);
or UO_148 (O_148,N_13890,N_13738);
or UO_149 (O_149,N_13983,N_13653);
or UO_150 (O_150,N_14749,N_14300);
nor UO_151 (O_151,N_14381,N_13784);
and UO_152 (O_152,N_14269,N_14544);
xor UO_153 (O_153,N_14447,N_13555);
and UO_154 (O_154,N_14189,N_14119);
xnor UO_155 (O_155,N_13790,N_14155);
or UO_156 (O_156,N_13800,N_14397);
and UO_157 (O_157,N_14177,N_14742);
or UO_158 (O_158,N_13861,N_13618);
nor UO_159 (O_159,N_14296,N_14253);
nand UO_160 (O_160,N_13780,N_14448);
and UO_161 (O_161,N_13636,N_14264);
xor UO_162 (O_162,N_13501,N_14421);
nor UO_163 (O_163,N_13601,N_14568);
or UO_164 (O_164,N_14302,N_14374);
nand UO_165 (O_165,N_13526,N_14456);
nand UO_166 (O_166,N_14788,N_14662);
and UO_167 (O_167,N_14245,N_13582);
nand UO_168 (O_168,N_14993,N_14617);
or UO_169 (O_169,N_14288,N_14640);
or UO_170 (O_170,N_13692,N_14961);
nand UO_171 (O_171,N_14652,N_14618);
nor UO_172 (O_172,N_13603,N_13600);
and UO_173 (O_173,N_14777,N_14888);
and UO_174 (O_174,N_14161,N_14949);
nor UO_175 (O_175,N_13535,N_13676);
nand UO_176 (O_176,N_14984,N_14712);
xnor UO_177 (O_177,N_14977,N_14594);
nand UO_178 (O_178,N_13813,N_13946);
xnor UO_179 (O_179,N_14200,N_13624);
xor UO_180 (O_180,N_14743,N_14806);
or UO_181 (O_181,N_13687,N_13686);
xor UO_182 (O_182,N_14669,N_14511);
xor UO_183 (O_183,N_13879,N_14457);
nand UO_184 (O_184,N_14077,N_14733);
nor UO_185 (O_185,N_14172,N_14531);
xor UO_186 (O_186,N_13593,N_13553);
nand UO_187 (O_187,N_13576,N_14923);
nand UO_188 (O_188,N_14094,N_14202);
and UO_189 (O_189,N_13892,N_14912);
or UO_190 (O_190,N_13940,N_14157);
nand UO_191 (O_191,N_14631,N_14084);
and UO_192 (O_192,N_13773,N_13753);
or UO_193 (O_193,N_13675,N_14786);
and UO_194 (O_194,N_14734,N_13803);
or UO_195 (O_195,N_14763,N_14057);
nand UO_196 (O_196,N_14477,N_13881);
or UO_197 (O_197,N_14887,N_14858);
or UO_198 (O_198,N_14995,N_13785);
nand UO_199 (O_199,N_13737,N_14331);
nor UO_200 (O_200,N_13652,N_14473);
or UO_201 (O_201,N_14135,N_13674);
xnor UO_202 (O_202,N_14645,N_13695);
xor UO_203 (O_203,N_13525,N_14826);
or UO_204 (O_204,N_13509,N_14045);
nor UO_205 (O_205,N_13901,N_14054);
nor UO_206 (O_206,N_14228,N_14073);
nand UO_207 (O_207,N_14595,N_14613);
nor UO_208 (O_208,N_14933,N_14506);
and UO_209 (O_209,N_13864,N_14744);
xnor UO_210 (O_210,N_14321,N_14388);
xor UO_211 (O_211,N_14880,N_14778);
and UO_212 (O_212,N_14185,N_13584);
or UO_213 (O_213,N_14985,N_13654);
or UO_214 (O_214,N_13677,N_14554);
xnor UO_215 (O_215,N_14082,N_13931);
or UO_216 (O_216,N_14934,N_14076);
or UO_217 (O_217,N_14700,N_14947);
or UO_218 (O_218,N_13745,N_13507);
nor UO_219 (O_219,N_14845,N_14364);
and UO_220 (O_220,N_13741,N_13723);
or UO_221 (O_221,N_14204,N_14259);
and UO_222 (O_222,N_14716,N_13583);
and UO_223 (O_223,N_13939,N_13767);
nor UO_224 (O_224,N_14738,N_14962);
or UO_225 (O_225,N_13841,N_14516);
or UO_226 (O_226,N_14637,N_13575);
nand UO_227 (O_227,N_14638,N_14215);
and UO_228 (O_228,N_13602,N_14056);
or UO_229 (O_229,N_14023,N_13808);
or UO_230 (O_230,N_13956,N_13838);
and UO_231 (O_231,N_14400,N_14883);
nand UO_232 (O_232,N_13938,N_14405);
nand UO_233 (O_233,N_14341,N_13797);
or UO_234 (O_234,N_14348,N_13891);
or UO_235 (O_235,N_13944,N_14188);
and UO_236 (O_236,N_14896,N_14470);
nand UO_237 (O_237,N_14849,N_14207);
or UO_238 (O_238,N_14035,N_14095);
nor UO_239 (O_239,N_13798,N_14032);
nand UO_240 (O_240,N_14164,N_14728);
nor UO_241 (O_241,N_13916,N_14825);
or UO_242 (O_242,N_13857,N_14768);
xor UO_243 (O_243,N_13963,N_14389);
nor UO_244 (O_244,N_13572,N_13519);
and UO_245 (O_245,N_13569,N_14335);
xor UO_246 (O_246,N_14193,N_14593);
nand UO_247 (O_247,N_14471,N_13763);
nand UO_248 (O_248,N_14061,N_14147);
nor UO_249 (O_249,N_14740,N_14093);
and UO_250 (O_250,N_13899,N_13516);
and UO_251 (O_251,N_14286,N_13659);
nor UO_252 (O_252,N_14665,N_14240);
xor UO_253 (O_253,N_13985,N_13997);
or UO_254 (O_254,N_14369,N_14661);
nand UO_255 (O_255,N_14863,N_13945);
and UO_256 (O_256,N_14158,N_13691);
nor UO_257 (O_257,N_14146,N_14861);
or UO_258 (O_258,N_13896,N_13978);
or UO_259 (O_259,N_14201,N_14794);
and UO_260 (O_260,N_14275,N_14824);
nor UO_261 (O_261,N_13598,N_13678);
and UO_262 (O_262,N_14066,N_14100);
or UO_263 (O_263,N_14795,N_14567);
nor UO_264 (O_264,N_14013,N_14811);
or UO_265 (O_265,N_14319,N_14678);
and UO_266 (O_266,N_13868,N_14103);
nor UO_267 (O_267,N_13964,N_14289);
or UO_268 (O_268,N_13799,N_14092);
nor UO_269 (O_269,N_13776,N_14783);
xnor UO_270 (O_270,N_14611,N_14946);
or UO_271 (O_271,N_13850,N_14149);
xnor UO_272 (O_272,N_13642,N_14573);
nor UO_273 (O_273,N_14187,N_14692);
and UO_274 (O_274,N_14705,N_14163);
nor UO_275 (O_275,N_13537,N_13789);
or UO_276 (O_276,N_13721,N_14636);
nor UO_277 (O_277,N_14479,N_14928);
nand UO_278 (O_278,N_14311,N_13903);
nor UO_279 (O_279,N_14250,N_14868);
nor UO_280 (O_280,N_14802,N_14726);
or UO_281 (O_281,N_14616,N_14835);
nand UO_282 (O_282,N_13651,N_14760);
nor UO_283 (O_283,N_13510,N_14875);
xor UO_284 (O_284,N_14116,N_14966);
nor UO_285 (O_285,N_13703,N_14028);
nand UO_286 (O_286,N_14725,N_13882);
nor UO_287 (O_287,N_13836,N_14431);
or UO_288 (O_288,N_14841,N_13697);
nand UO_289 (O_289,N_14553,N_14590);
nor UO_290 (O_290,N_14104,N_14753);
nand UO_291 (O_291,N_14755,N_13949);
and UO_292 (O_292,N_14512,N_14800);
xor UO_293 (O_293,N_14106,N_14343);
and UO_294 (O_294,N_14342,N_13669);
nor UO_295 (O_295,N_14674,N_14340);
or UO_296 (O_296,N_14140,N_14680);
nand UO_297 (O_297,N_13585,N_14922);
nor UO_298 (O_298,N_13690,N_13829);
xnor UO_299 (O_299,N_14754,N_13512);
nand UO_300 (O_300,N_14360,N_14663);
or UO_301 (O_301,N_14925,N_14173);
nand UO_302 (O_302,N_14885,N_13567);
or UO_303 (O_303,N_14014,N_14322);
and UO_304 (O_304,N_14780,N_14294);
and UO_305 (O_305,N_14070,N_14548);
or UO_306 (O_306,N_13532,N_14458);
xnor UO_307 (O_307,N_14650,N_14366);
or UO_308 (O_308,N_14520,N_14871);
nor UO_309 (O_309,N_14058,N_14442);
xnor UO_310 (O_310,N_13505,N_14263);
or UO_311 (O_311,N_13756,N_14980);
nor UO_312 (O_312,N_13587,N_14078);
nor UO_313 (O_313,N_14644,N_13708);
nor UO_314 (O_314,N_14238,N_14790);
nor UO_315 (O_315,N_14295,N_14387);
and UO_316 (O_316,N_13958,N_13772);
or UO_317 (O_317,N_13818,N_14299);
nand UO_318 (O_318,N_13645,N_14706);
or UO_319 (O_319,N_14208,N_14102);
and UO_320 (O_320,N_14936,N_14990);
xnor UO_321 (O_321,N_13580,N_14019);
xor UO_322 (O_322,N_14246,N_14536);
nand UO_323 (O_323,N_14505,N_14336);
nor UO_324 (O_324,N_14569,N_13664);
nand UO_325 (O_325,N_14420,N_14660);
nand UO_326 (O_326,N_14565,N_13782);
xor UO_327 (O_327,N_14821,N_13760);
nor UO_328 (O_328,N_13911,N_14775);
nand UO_329 (O_329,N_14074,N_13993);
nor UO_330 (O_330,N_13906,N_13529);
xnor UO_331 (O_331,N_14174,N_13656);
nor UO_332 (O_332,N_13926,N_14181);
xnor UO_333 (O_333,N_14406,N_13614);
nand UO_334 (O_334,N_13571,N_13545);
xnor UO_335 (O_335,N_13795,N_14939);
nor UO_336 (O_336,N_14393,N_14996);
xor UO_337 (O_337,N_14133,N_13710);
or UO_338 (O_338,N_14975,N_14426);
nand UO_339 (O_339,N_14673,N_13846);
nand UO_340 (O_340,N_14399,N_13592);
xnor UO_341 (O_341,N_14600,N_14687);
nand UO_342 (O_342,N_14223,N_14087);
or UO_343 (O_343,N_14765,N_14641);
nor UO_344 (O_344,N_14128,N_14410);
nand UO_345 (O_345,N_14352,N_13701);
nor UO_346 (O_346,N_13876,N_14708);
xor UO_347 (O_347,N_14735,N_13641);
and UO_348 (O_348,N_14383,N_14099);
nor UO_349 (O_349,N_14664,N_14686);
nor UO_350 (O_350,N_14831,N_13959);
nor UO_351 (O_351,N_14186,N_14121);
xnor UO_352 (O_352,N_14535,N_14209);
or UO_353 (O_353,N_13568,N_13515);
nand UO_354 (O_354,N_14944,N_14670);
and UO_355 (O_355,N_14968,N_13565);
nor UO_356 (O_356,N_13597,N_14866);
nand UO_357 (O_357,N_13578,N_14750);
xor UO_358 (O_358,N_14971,N_14018);
and UO_359 (O_359,N_13820,N_14619);
and UO_360 (O_360,N_14697,N_14170);
nand UO_361 (O_361,N_13632,N_13518);
and UO_362 (O_362,N_13929,N_14585);
xnor UO_363 (O_363,N_14222,N_14759);
nand UO_364 (O_364,N_13542,N_14049);
nor UO_365 (O_365,N_14122,N_14864);
nand UO_366 (O_366,N_14558,N_14731);
nand UO_367 (O_367,N_13937,N_14764);
and UO_368 (O_368,N_14293,N_13606);
or UO_369 (O_369,N_14545,N_14191);
and UO_370 (O_370,N_13842,N_14145);
or UO_371 (O_371,N_14459,N_14432);
xor UO_372 (O_372,N_14509,N_14502);
or UO_373 (O_373,N_14599,N_14422);
or UO_374 (O_374,N_14235,N_13976);
and UO_375 (O_375,N_14257,N_14938);
and UO_376 (O_376,N_13886,N_14368);
xor UO_377 (O_377,N_14997,N_14039);
nand UO_378 (O_378,N_14691,N_14454);
nor UO_379 (O_379,N_14464,N_14540);
and UO_380 (O_380,N_13880,N_14521);
or UO_381 (O_381,N_14136,N_13661);
nand UO_382 (O_382,N_13660,N_14062);
nor UO_383 (O_383,N_14908,N_14409);
xnor UO_384 (O_384,N_13843,N_14358);
or UO_385 (O_385,N_13854,N_14654);
nor UO_386 (O_386,N_13508,N_14085);
and UO_387 (O_387,N_14168,N_14355);
nand UO_388 (O_388,N_13693,N_14634);
nand UO_389 (O_389,N_14040,N_14773);
nor UO_390 (O_390,N_14776,N_13920);
nor UO_391 (O_391,N_13536,N_14587);
nand UO_392 (O_392,N_13819,N_13607);
xor UO_393 (O_393,N_13524,N_14881);
and UO_394 (O_394,N_14874,N_13977);
nand UO_395 (O_395,N_14361,N_14460);
nand UO_396 (O_396,N_14891,N_13972);
and UO_397 (O_397,N_13766,N_13863);
and UO_398 (O_398,N_14904,N_14266);
xnor UO_399 (O_399,N_14015,N_14031);
xnor UO_400 (O_400,N_13655,N_14965);
or UO_401 (O_401,N_14862,N_14577);
xnor UO_402 (O_402,N_14159,N_13646);
xor UO_403 (O_403,N_13809,N_14262);
nor UO_404 (O_404,N_14817,N_14926);
nor UO_405 (O_405,N_14098,N_14394);
or UO_406 (O_406,N_14930,N_14667);
nand UO_407 (O_407,N_14672,N_14027);
nand UO_408 (O_408,N_13950,N_14886);
xnor UO_409 (O_409,N_14550,N_14510);
and UO_410 (O_410,N_14827,N_14808);
nand UO_411 (O_411,N_13506,N_14621);
or UO_412 (O_412,N_14236,N_13706);
or UO_413 (O_413,N_14329,N_13837);
or UO_414 (O_414,N_14055,N_14801);
or UO_415 (O_415,N_14605,N_14010);
nand UO_416 (O_416,N_13657,N_14446);
nor UO_417 (O_417,N_14689,N_13668);
and UO_418 (O_418,N_13771,N_14425);
and UO_419 (O_419,N_13812,N_14379);
nor UO_420 (O_420,N_13726,N_14829);
nand UO_421 (O_421,N_14060,N_14982);
nand UO_422 (O_422,N_14570,N_14385);
xnor UO_423 (O_423,N_14449,N_14433);
or UO_424 (O_424,N_14408,N_14450);
nor UO_425 (O_425,N_13557,N_14720);
or UO_426 (O_426,N_14752,N_14254);
nand UO_427 (O_427,N_13548,N_14000);
nor UO_428 (O_428,N_14581,N_14445);
xnor UO_429 (O_429,N_14972,N_13962);
nand UO_430 (O_430,N_14436,N_13617);
nand UO_431 (O_431,N_14414,N_14649);
xnor UO_432 (O_432,N_14789,N_14079);
nor UO_433 (O_433,N_13640,N_14856);
xor UO_434 (O_434,N_14113,N_14959);
nand UO_435 (O_435,N_14255,N_14701);
and UO_436 (O_436,N_14219,N_14047);
xor UO_437 (O_437,N_13541,N_13999);
nand UO_438 (O_438,N_13865,N_14378);
xor UO_439 (O_439,N_13832,N_14561);
nand UO_440 (O_440,N_13831,N_14999);
nand UO_441 (O_441,N_14953,N_14430);
nand UO_442 (O_442,N_13742,N_13630);
xnor UO_443 (O_443,N_13875,N_14022);
or UO_444 (O_444,N_14413,N_14530);
or UO_445 (O_445,N_14895,N_14782);
xor UO_446 (O_446,N_14490,N_14232);
and UO_447 (O_447,N_13589,N_13604);
nor UO_448 (O_448,N_14205,N_14848);
nor UO_449 (O_449,N_14278,N_13720);
or UO_450 (O_450,N_14130,N_14024);
or UO_451 (O_451,N_14249,N_13815);
xor UO_452 (O_452,N_14111,N_14108);
xnor UO_453 (O_453,N_13716,N_14052);
xnor UO_454 (O_454,N_14941,N_14867);
or UO_455 (O_455,N_14213,N_14080);
nor UO_456 (O_456,N_13822,N_14994);
nor UO_457 (O_457,N_14730,N_14940);
or UO_458 (O_458,N_14325,N_13947);
nand UO_459 (O_459,N_14350,N_14469);
nor UO_460 (O_460,N_14717,N_14907);
nor UO_461 (O_461,N_13765,N_14001);
or UO_462 (O_462,N_14372,N_14514);
xnor UO_463 (O_463,N_13625,N_14659);
or UO_464 (O_464,N_14551,N_14036);
nand UO_465 (O_465,N_13827,N_13670);
or UO_466 (O_466,N_14836,N_14951);
nor UO_467 (O_467,N_13513,N_13744);
xnor UO_468 (O_468,N_14620,N_13629);
nand UO_469 (O_469,N_13715,N_14345);
nor UO_470 (O_470,N_13779,N_13981);
and UO_471 (O_471,N_14244,N_14956);
or UO_472 (O_472,N_14486,N_14380);
nor UO_473 (O_473,N_14198,N_14091);
nand UO_474 (O_474,N_14129,N_14112);
nand UO_475 (O_475,N_14065,N_13761);
and UO_476 (O_476,N_13556,N_13893);
nor UO_477 (O_477,N_13919,N_14844);
and UO_478 (O_478,N_14237,N_13561);
and UO_479 (O_479,N_14171,N_14578);
nand UO_480 (O_480,N_13644,N_13866);
nor UO_481 (O_481,N_13874,N_14349);
nand UO_482 (O_482,N_13817,N_14927);
and UO_483 (O_483,N_13560,N_14008);
xor UO_484 (O_484,N_13543,N_14416);
xor UO_485 (O_485,N_14815,N_14932);
nand UO_486 (O_486,N_13954,N_13791);
or UO_487 (O_487,N_14429,N_14401);
nand UO_488 (O_488,N_13705,N_13996);
nor UO_489 (O_489,N_13979,N_14279);
and UO_490 (O_490,N_14224,N_14498);
or UO_491 (O_491,N_13534,N_13867);
and UO_492 (O_492,N_14899,N_14309);
xor UO_493 (O_493,N_14761,N_13895);
nand UO_494 (O_494,N_14707,N_14353);
xnor UO_495 (O_495,N_14557,N_13951);
and UO_496 (O_496,N_14306,N_14656);
or UO_497 (O_497,N_14156,N_14770);
nand UO_498 (O_498,N_14251,N_13762);
xor UO_499 (O_499,N_14830,N_14910);
nor UO_500 (O_500,N_14525,N_13672);
and UO_501 (O_501,N_13821,N_14214);
or UO_502 (O_502,N_14267,N_13998);
nand UO_503 (O_503,N_14182,N_13638);
nor UO_504 (O_504,N_14623,N_14767);
nand UO_505 (O_505,N_14217,N_14547);
nand UO_506 (O_506,N_14417,N_13666);
nand UO_507 (O_507,N_14724,N_13734);
and UO_508 (O_508,N_14179,N_14698);
and UO_509 (O_509,N_14114,N_14602);
nand UO_510 (O_510,N_14828,N_13770);
nor UO_511 (O_511,N_14846,N_13647);
xor UO_512 (O_512,N_13611,N_13872);
nand UO_513 (O_513,N_13847,N_14741);
nand UO_514 (O_514,N_14373,N_13984);
xnor UO_515 (O_515,N_13952,N_14120);
nand UO_516 (O_516,N_14481,N_14900);
nor UO_517 (O_517,N_14906,N_13936);
xnor UO_518 (O_518,N_14377,N_14890);
or UO_519 (O_519,N_14612,N_14822);
nand UO_520 (O_520,N_13724,N_13533);
or UO_521 (O_521,N_14586,N_13633);
nor UO_522 (O_522,N_13746,N_13540);
or UO_523 (O_523,N_14676,N_13667);
nand UO_524 (O_524,N_14729,N_14559);
xor UO_525 (O_525,N_13613,N_13750);
nor UO_526 (O_526,N_13844,N_13743);
xnor UO_527 (O_527,N_14153,N_14180);
nand UO_528 (O_528,N_14315,N_14491);
nor UO_529 (O_529,N_14920,N_14924);
nand UO_530 (O_530,N_13562,N_13987);
and UO_531 (O_531,N_13733,N_13658);
nand UO_532 (O_532,N_13530,N_14879);
xor UO_533 (O_533,N_14258,N_14284);
nor UO_534 (O_534,N_14067,N_13649);
xnor UO_535 (O_535,N_14583,N_13696);
nand UO_536 (O_536,N_14865,N_13973);
nor UO_537 (O_537,N_13704,N_14487);
and UO_538 (O_538,N_14630,N_13900);
and UO_539 (O_539,N_14709,N_14931);
nor UO_540 (O_540,N_13883,N_14837);
xnor UO_541 (O_541,N_13605,N_13590);
or UO_542 (O_542,N_14020,N_13910);
xnor UO_543 (O_543,N_14206,N_13941);
nand UO_544 (O_544,N_13596,N_14703);
nor UO_545 (O_545,N_14608,N_14362);
xnor UO_546 (O_546,N_14003,N_14184);
nand UO_547 (O_547,N_14969,N_14747);
xnor UO_548 (O_548,N_14571,N_14227);
xor UO_549 (O_549,N_14150,N_13825);
nor UO_550 (O_550,N_13873,N_14694);
nor UO_551 (O_551,N_14596,N_13559);
nor UO_552 (O_552,N_14842,N_14769);
and UO_553 (O_553,N_14632,N_13719);
nor UO_554 (O_554,N_14051,N_14653);
nand UO_555 (O_555,N_13870,N_14658);
and UO_556 (O_556,N_13807,N_14351);
and UO_557 (O_557,N_14816,N_14216);
xnor UO_558 (O_558,N_14005,N_13871);
nor UO_559 (O_559,N_14166,N_14766);
and UO_560 (O_560,N_14301,N_14466);
xor UO_561 (O_561,N_14376,N_13908);
nand UO_562 (O_562,N_14115,N_14542);
nand UO_563 (O_563,N_13554,N_14404);
or UO_564 (O_564,N_13731,N_14897);
xnor UO_565 (O_565,N_13550,N_14075);
xor UO_566 (O_566,N_14139,N_14718);
nand UO_567 (O_567,N_13924,N_13639);
xnor UO_568 (O_568,N_14840,N_14453);
nand UO_569 (O_569,N_14838,N_13918);
nand UO_570 (O_570,N_14034,N_13621);
xor UO_571 (O_571,N_14328,N_14798);
nor UO_572 (O_572,N_13823,N_13683);
nand UO_573 (O_573,N_13739,N_14012);
nor UO_574 (O_574,N_14657,N_14290);
nand UO_575 (O_575,N_14320,N_13759);
and UO_576 (O_576,N_14677,N_14248);
nand UO_577 (O_577,N_14721,N_13714);
nand UO_578 (O_578,N_13517,N_14307);
or UO_579 (O_579,N_14736,N_14437);
nand UO_580 (O_580,N_14523,N_13970);
or UO_581 (O_581,N_14988,N_14212);
and UO_582 (O_582,N_13631,N_14850);
nor UO_583 (O_583,N_14048,N_14195);
and UO_584 (O_584,N_14549,N_14088);
xnor UO_585 (O_585,N_14655,N_14648);
or UO_586 (O_586,N_14344,N_13758);
xor UO_587 (O_587,N_14126,N_14592);
or UO_588 (O_588,N_14683,N_13930);
xor UO_589 (O_589,N_14919,N_14601);
nand UO_590 (O_590,N_14713,N_13679);
nand UO_591 (O_591,N_14109,N_14468);
xor UO_592 (O_592,N_13662,N_14852);
nor UO_593 (O_593,N_13511,N_13622);
and UO_594 (O_594,N_14804,N_13539);
nor UO_595 (O_595,N_13523,N_14333);
xnor UO_596 (O_596,N_14974,N_14137);
nor UO_597 (O_597,N_13948,N_14960);
nor UO_598 (O_598,N_14857,N_13778);
and UO_599 (O_599,N_14543,N_14784);
xor UO_600 (O_600,N_14834,N_13933);
or UO_601 (O_601,N_13845,N_14064);
nor UO_602 (O_602,N_13635,N_14610);
xnor UO_603 (O_603,N_14681,N_14529);
and UO_604 (O_604,N_14326,N_14869);
and UO_605 (O_605,N_14955,N_14354);
xnor UO_606 (O_606,N_14461,N_14522);
nand UO_607 (O_607,N_13610,N_14945);
nand UO_608 (O_608,N_13579,N_14541);
nand UO_609 (O_609,N_14588,N_14983);
xnor UO_610 (O_610,N_14402,N_13728);
or UO_611 (O_611,N_14242,N_13681);
nand UO_612 (O_612,N_13988,N_14427);
or UO_613 (O_613,N_14562,N_14229);
xor UO_614 (O_614,N_14903,N_13700);
nand UO_615 (O_615,N_13849,N_14534);
and UO_616 (O_616,N_13806,N_13757);
xnor UO_617 (O_617,N_14046,N_14029);
or UO_618 (O_618,N_14265,N_14059);
or UO_619 (O_619,N_14312,N_14494);
and UO_620 (O_620,N_13740,N_14859);
nor UO_621 (O_621,N_14970,N_14624);
nor UO_622 (O_622,N_14853,N_14998);
or UO_623 (O_623,N_14564,N_14576);
xnor UO_624 (O_624,N_14533,N_14443);
xor UO_625 (O_625,N_14452,N_14905);
xor UO_626 (O_626,N_14696,N_14291);
xor UO_627 (O_627,N_13709,N_14132);
or UO_628 (O_628,N_14651,N_13902);
nor UO_629 (O_629,N_14710,N_14532);
or UO_630 (O_630,N_13943,N_14451);
and UO_631 (O_631,N_13968,N_14165);
and UO_632 (O_632,N_14261,N_14123);
nor UO_633 (O_633,N_14305,N_13888);
nand UO_634 (O_634,N_14127,N_14913);
or UO_635 (O_635,N_14484,N_14371);
or UO_636 (O_636,N_14475,N_14504);
or UO_637 (O_637,N_14463,N_14347);
or UO_638 (O_638,N_14148,N_13764);
xor UO_639 (O_639,N_13897,N_14507);
nand UO_640 (O_640,N_13732,N_14403);
and UO_641 (O_641,N_13694,N_14225);
or UO_642 (O_642,N_14914,N_14714);
xnor UO_643 (O_643,N_13852,N_14280);
or UO_644 (O_644,N_14101,N_14627);
nand UO_645 (O_645,N_13628,N_14283);
or UO_646 (O_646,N_14338,N_13546);
nor UO_647 (O_647,N_14230,N_13609);
nor UO_648 (O_648,N_14715,N_14758);
or UO_649 (O_649,N_14038,N_14178);
nor UO_650 (O_650,N_13833,N_14105);
nand UO_651 (O_651,N_14492,N_14820);
xnor UO_652 (O_652,N_13698,N_14382);
or UO_653 (O_653,N_13967,N_14807);
xor UO_654 (O_654,N_14702,N_13626);
xnor UO_655 (O_655,N_14584,N_14792);
xnor UO_656 (O_656,N_14274,N_14732);
nand UO_657 (O_657,N_13581,N_14935);
or UO_658 (O_658,N_13914,N_13684);
nand UO_659 (O_659,N_13735,N_14192);
nand UO_660 (O_660,N_13612,N_13898);
or UO_661 (O_661,N_13792,N_14527);
nand UO_662 (O_662,N_14392,N_13573);
xnor UO_663 (O_663,N_14474,N_14943);
or UO_664 (O_664,N_14297,N_14915);
or UO_665 (O_665,N_14359,N_14292);
nand UO_666 (O_666,N_13786,N_13991);
nand UO_667 (O_667,N_14063,N_14882);
nor UO_668 (O_668,N_14832,N_14428);
nand UO_669 (O_669,N_14851,N_14515);
nand UO_670 (O_670,N_14439,N_14884);
and UO_671 (O_671,N_14668,N_14818);
and UO_672 (O_672,N_14107,N_14308);
or UO_673 (O_673,N_13788,N_14756);
xnor UO_674 (O_674,N_14823,N_14916);
nor UO_675 (O_675,N_14785,N_14937);
or UO_676 (O_676,N_13594,N_13637);
and UO_677 (O_677,N_13616,N_14762);
nor UO_678 (O_678,N_13955,N_14719);
and UO_679 (O_679,N_14860,N_13503);
xnor UO_680 (O_680,N_14438,N_13859);
xnor UO_681 (O_681,N_14298,N_14281);
nand UO_682 (O_682,N_14418,N_14633);
or UO_683 (O_683,N_14781,N_14873);
and UO_684 (O_684,N_14805,N_14580);
or UO_685 (O_685,N_14314,N_14963);
nand UO_686 (O_686,N_14957,N_14485);
and UO_687 (O_687,N_13928,N_14190);
or UO_688 (O_688,N_14606,N_14981);
nor UO_689 (O_689,N_13522,N_14391);
nand UO_690 (O_690,N_14991,N_14050);
nor UO_691 (O_691,N_13514,N_14855);
nor UO_692 (O_692,N_14154,N_14488);
nor UO_693 (O_693,N_14796,N_14797);
nand UO_694 (O_694,N_13547,N_14489);
nand UO_695 (O_695,N_14285,N_13975);
xor UO_696 (O_696,N_14739,N_13650);
xnor UO_697 (O_697,N_14042,N_13994);
and UO_698 (O_698,N_14304,N_14234);
or UO_699 (O_699,N_14016,N_14444);
or UO_700 (O_700,N_14603,N_14572);
nand UO_701 (O_701,N_13885,N_14642);
xnor UO_702 (O_702,N_14870,N_14196);
and UO_703 (O_703,N_13729,N_14575);
and UO_704 (O_704,N_14591,N_13858);
and UO_705 (O_705,N_14125,N_14317);
and UO_706 (O_706,N_14909,N_14843);
and UO_707 (O_707,N_13995,N_13856);
or UO_708 (O_708,N_14876,N_13685);
nand UO_709 (O_709,N_14917,N_14243);
nand UO_710 (O_710,N_13527,N_13586);
nand UO_711 (O_711,N_14574,N_14081);
xor UO_712 (O_712,N_14231,N_14097);
xor UO_713 (O_713,N_13748,N_14138);
nor UO_714 (O_714,N_14194,N_13826);
xor UO_715 (O_715,N_13608,N_14814);
nand UO_716 (O_716,N_14118,N_14679);
nand UO_717 (O_717,N_14508,N_14318);
nor UO_718 (O_718,N_13787,N_13552);
or UO_719 (O_719,N_14086,N_13713);
or UO_720 (O_720,N_14751,N_14745);
and UO_721 (O_721,N_14324,N_13563);
and UO_722 (O_722,N_14682,N_14169);
nor UO_723 (O_723,N_13839,N_14695);
or UO_724 (O_724,N_14356,N_14441);
xnor UO_725 (O_725,N_14978,N_13521);
or UO_726 (O_726,N_13913,N_13992);
nand UO_727 (O_727,N_14483,N_14690);
or UO_728 (O_728,N_14519,N_13793);
nand UO_729 (O_729,N_13777,N_14727);
or UO_730 (O_730,N_13711,N_13824);
nor UO_731 (O_731,N_13768,N_13781);
xor UO_732 (O_732,N_14964,N_14787);
and UO_733 (O_733,N_13774,N_14203);
nand UO_734 (O_734,N_14440,N_14604);
and UO_735 (O_735,N_14911,N_14467);
or UO_736 (O_736,N_14812,N_14268);
xor UO_737 (O_737,N_13643,N_14334);
nand UO_738 (O_738,N_13520,N_13702);
and UO_739 (O_739,N_13671,N_14247);
nand UO_740 (O_740,N_14779,N_14892);
or UO_741 (O_741,N_13783,N_13965);
nand UO_742 (O_742,N_13619,N_14598);
and UO_743 (O_743,N_13923,N_13835);
and UO_744 (O_744,N_14872,N_13634);
nor UO_745 (O_745,N_14423,N_14671);
nand UO_746 (O_746,N_14396,N_14950);
nor UO_747 (O_747,N_14090,N_13810);
nand UO_748 (O_748,N_14004,N_14685);
xnor UO_749 (O_749,N_13717,N_14233);
or UO_750 (O_750,N_14130,N_14282);
nand UO_751 (O_751,N_14062,N_14704);
and UO_752 (O_752,N_14304,N_13589);
xnor UO_753 (O_753,N_13718,N_13890);
nand UO_754 (O_754,N_14207,N_13996);
nand UO_755 (O_755,N_14185,N_14998);
xnor UO_756 (O_756,N_14966,N_14300);
and UO_757 (O_757,N_14714,N_14039);
and UO_758 (O_758,N_13818,N_14777);
or UO_759 (O_759,N_13631,N_14187);
nor UO_760 (O_760,N_14011,N_13775);
xor UO_761 (O_761,N_14554,N_14431);
xor UO_762 (O_762,N_14486,N_13570);
nor UO_763 (O_763,N_14518,N_14879);
or UO_764 (O_764,N_13576,N_14546);
and UO_765 (O_765,N_13613,N_14092);
or UO_766 (O_766,N_14846,N_13837);
nand UO_767 (O_767,N_14063,N_14789);
nand UO_768 (O_768,N_14153,N_13818);
nand UO_769 (O_769,N_14667,N_14805);
or UO_770 (O_770,N_13949,N_14359);
nor UO_771 (O_771,N_13759,N_14924);
xor UO_772 (O_772,N_14622,N_14367);
nand UO_773 (O_773,N_14133,N_14480);
and UO_774 (O_774,N_14825,N_13737);
xor UO_775 (O_775,N_13825,N_13784);
and UO_776 (O_776,N_14495,N_14882);
nor UO_777 (O_777,N_14914,N_14092);
and UO_778 (O_778,N_14222,N_14048);
xnor UO_779 (O_779,N_14284,N_14432);
nand UO_780 (O_780,N_14186,N_13862);
or UO_781 (O_781,N_13649,N_13992);
xor UO_782 (O_782,N_13651,N_14161);
nor UO_783 (O_783,N_13640,N_14671);
or UO_784 (O_784,N_14336,N_14119);
nand UO_785 (O_785,N_14019,N_13501);
or UO_786 (O_786,N_14234,N_13639);
and UO_787 (O_787,N_14658,N_13656);
nand UO_788 (O_788,N_14598,N_13990);
and UO_789 (O_789,N_14210,N_14569);
or UO_790 (O_790,N_13679,N_14780);
nand UO_791 (O_791,N_14271,N_13890);
nand UO_792 (O_792,N_14823,N_13566);
nand UO_793 (O_793,N_14180,N_14833);
or UO_794 (O_794,N_14045,N_14713);
or UO_795 (O_795,N_14053,N_14172);
and UO_796 (O_796,N_13932,N_13598);
or UO_797 (O_797,N_14193,N_14081);
or UO_798 (O_798,N_14217,N_14233);
nor UO_799 (O_799,N_14198,N_14047);
nand UO_800 (O_800,N_13893,N_14517);
nor UO_801 (O_801,N_14545,N_13884);
nor UO_802 (O_802,N_14984,N_14397);
nor UO_803 (O_803,N_13622,N_14665);
xor UO_804 (O_804,N_14738,N_14849);
nor UO_805 (O_805,N_14642,N_14525);
nand UO_806 (O_806,N_13718,N_13529);
nand UO_807 (O_807,N_14634,N_14427);
nor UO_808 (O_808,N_14988,N_13734);
or UO_809 (O_809,N_13557,N_13671);
nor UO_810 (O_810,N_13654,N_13594);
xor UO_811 (O_811,N_14084,N_14028);
or UO_812 (O_812,N_13640,N_14411);
or UO_813 (O_813,N_13902,N_14390);
nor UO_814 (O_814,N_14476,N_14070);
nand UO_815 (O_815,N_14226,N_13846);
nand UO_816 (O_816,N_13635,N_14712);
nor UO_817 (O_817,N_13696,N_14264);
nand UO_818 (O_818,N_14814,N_14671);
or UO_819 (O_819,N_13794,N_14322);
xor UO_820 (O_820,N_13928,N_13610);
and UO_821 (O_821,N_14312,N_14231);
or UO_822 (O_822,N_14700,N_13695);
xor UO_823 (O_823,N_14084,N_14365);
and UO_824 (O_824,N_14272,N_14951);
xor UO_825 (O_825,N_14140,N_14148);
and UO_826 (O_826,N_14688,N_13701);
nor UO_827 (O_827,N_14762,N_14374);
xor UO_828 (O_828,N_14194,N_14692);
xor UO_829 (O_829,N_13846,N_14432);
nor UO_830 (O_830,N_13860,N_14959);
nand UO_831 (O_831,N_13900,N_14212);
nand UO_832 (O_832,N_14514,N_13644);
xor UO_833 (O_833,N_14415,N_13664);
or UO_834 (O_834,N_14334,N_14611);
or UO_835 (O_835,N_14021,N_13955);
or UO_836 (O_836,N_13905,N_14127);
nor UO_837 (O_837,N_13673,N_13717);
or UO_838 (O_838,N_13886,N_14388);
xnor UO_839 (O_839,N_14713,N_14546);
nand UO_840 (O_840,N_14406,N_14697);
nand UO_841 (O_841,N_14768,N_14681);
and UO_842 (O_842,N_14439,N_14805);
nand UO_843 (O_843,N_14140,N_13743);
or UO_844 (O_844,N_14609,N_14657);
nand UO_845 (O_845,N_13556,N_14473);
and UO_846 (O_846,N_14752,N_13500);
nor UO_847 (O_847,N_14484,N_14119);
nand UO_848 (O_848,N_13711,N_14143);
or UO_849 (O_849,N_13680,N_14277);
nor UO_850 (O_850,N_14678,N_14789);
nand UO_851 (O_851,N_14684,N_14269);
xnor UO_852 (O_852,N_14214,N_14983);
or UO_853 (O_853,N_14404,N_14281);
or UO_854 (O_854,N_14699,N_14693);
nand UO_855 (O_855,N_13519,N_13541);
xnor UO_856 (O_856,N_14641,N_14818);
or UO_857 (O_857,N_13613,N_14238);
or UO_858 (O_858,N_14745,N_14324);
and UO_859 (O_859,N_14725,N_14272);
nor UO_860 (O_860,N_14130,N_13998);
and UO_861 (O_861,N_14454,N_14358);
xnor UO_862 (O_862,N_13924,N_14828);
nand UO_863 (O_863,N_14419,N_13656);
or UO_864 (O_864,N_14908,N_14737);
nand UO_865 (O_865,N_14199,N_14256);
and UO_866 (O_866,N_13555,N_14960);
and UO_867 (O_867,N_14633,N_13875);
nor UO_868 (O_868,N_14647,N_14381);
and UO_869 (O_869,N_14971,N_14622);
nor UO_870 (O_870,N_14316,N_14666);
nor UO_871 (O_871,N_14358,N_13562);
xnor UO_872 (O_872,N_14867,N_14323);
xor UO_873 (O_873,N_13713,N_14269);
or UO_874 (O_874,N_14000,N_13967);
and UO_875 (O_875,N_13569,N_14337);
and UO_876 (O_876,N_13762,N_13866);
nand UO_877 (O_877,N_13637,N_14501);
and UO_878 (O_878,N_14675,N_13670);
nand UO_879 (O_879,N_14632,N_13760);
nor UO_880 (O_880,N_13500,N_14324);
xor UO_881 (O_881,N_14157,N_13626);
or UO_882 (O_882,N_14940,N_13959);
and UO_883 (O_883,N_13628,N_14624);
xor UO_884 (O_884,N_14023,N_14505);
and UO_885 (O_885,N_13599,N_14909);
nor UO_886 (O_886,N_13503,N_13978);
nor UO_887 (O_887,N_14123,N_14567);
xor UO_888 (O_888,N_14003,N_14543);
and UO_889 (O_889,N_14699,N_14896);
and UO_890 (O_890,N_14738,N_14522);
and UO_891 (O_891,N_13683,N_14796);
or UO_892 (O_892,N_13698,N_14619);
nand UO_893 (O_893,N_13973,N_14098);
xnor UO_894 (O_894,N_13877,N_14439);
nand UO_895 (O_895,N_14490,N_13740);
xnor UO_896 (O_896,N_14177,N_13807);
and UO_897 (O_897,N_14834,N_13962);
and UO_898 (O_898,N_14513,N_14052);
and UO_899 (O_899,N_14602,N_14393);
xnor UO_900 (O_900,N_13787,N_14043);
nor UO_901 (O_901,N_14986,N_13901);
or UO_902 (O_902,N_14331,N_13980);
and UO_903 (O_903,N_13596,N_13787);
or UO_904 (O_904,N_14288,N_14997);
and UO_905 (O_905,N_13611,N_14508);
or UO_906 (O_906,N_13773,N_13928);
xnor UO_907 (O_907,N_14868,N_14295);
xnor UO_908 (O_908,N_13824,N_14512);
nor UO_909 (O_909,N_14940,N_13585);
xnor UO_910 (O_910,N_13644,N_13634);
or UO_911 (O_911,N_14071,N_14449);
nor UO_912 (O_912,N_14724,N_13526);
nand UO_913 (O_913,N_13510,N_13759);
nand UO_914 (O_914,N_14086,N_14052);
nand UO_915 (O_915,N_14332,N_14919);
or UO_916 (O_916,N_13563,N_13971);
nor UO_917 (O_917,N_14070,N_14006);
and UO_918 (O_918,N_14756,N_14841);
xor UO_919 (O_919,N_14620,N_14510);
nor UO_920 (O_920,N_14607,N_14447);
xor UO_921 (O_921,N_13741,N_14592);
xor UO_922 (O_922,N_14693,N_14225);
or UO_923 (O_923,N_13836,N_13544);
xor UO_924 (O_924,N_14115,N_14923);
and UO_925 (O_925,N_14346,N_14059);
xnor UO_926 (O_926,N_14159,N_14190);
and UO_927 (O_927,N_14107,N_13703);
and UO_928 (O_928,N_14513,N_14258);
xnor UO_929 (O_929,N_14056,N_14196);
nor UO_930 (O_930,N_14769,N_14283);
nand UO_931 (O_931,N_14492,N_13980);
and UO_932 (O_932,N_14640,N_14213);
xnor UO_933 (O_933,N_14394,N_14859);
nand UO_934 (O_934,N_14457,N_14886);
and UO_935 (O_935,N_13811,N_13943);
nor UO_936 (O_936,N_14911,N_13738);
xnor UO_937 (O_937,N_14039,N_14237);
or UO_938 (O_938,N_13967,N_14323);
and UO_939 (O_939,N_14785,N_14670);
nand UO_940 (O_940,N_14644,N_14130);
nor UO_941 (O_941,N_14777,N_13869);
nor UO_942 (O_942,N_13794,N_14004);
nand UO_943 (O_943,N_13659,N_13540);
xor UO_944 (O_944,N_13868,N_14900);
nor UO_945 (O_945,N_14773,N_14087);
and UO_946 (O_946,N_13976,N_14044);
nand UO_947 (O_947,N_14173,N_14582);
nor UO_948 (O_948,N_13861,N_14550);
nand UO_949 (O_949,N_13656,N_13636);
xor UO_950 (O_950,N_14832,N_14840);
nand UO_951 (O_951,N_14402,N_14825);
nor UO_952 (O_952,N_14617,N_13914);
nor UO_953 (O_953,N_14063,N_13915);
or UO_954 (O_954,N_14701,N_13717);
and UO_955 (O_955,N_14848,N_14190);
and UO_956 (O_956,N_13950,N_14490);
nand UO_957 (O_957,N_14852,N_14646);
and UO_958 (O_958,N_14615,N_14862);
or UO_959 (O_959,N_13910,N_13624);
nand UO_960 (O_960,N_13703,N_14211);
nor UO_961 (O_961,N_14838,N_14634);
xnor UO_962 (O_962,N_13608,N_14278);
nand UO_963 (O_963,N_14861,N_14547);
nor UO_964 (O_964,N_13648,N_13768);
nand UO_965 (O_965,N_14018,N_14314);
xor UO_966 (O_966,N_13940,N_14112);
or UO_967 (O_967,N_14997,N_13641);
or UO_968 (O_968,N_14054,N_13603);
or UO_969 (O_969,N_14531,N_14486);
nand UO_970 (O_970,N_13823,N_14375);
or UO_971 (O_971,N_14660,N_14415);
nand UO_972 (O_972,N_13669,N_14076);
nor UO_973 (O_973,N_13763,N_13767);
or UO_974 (O_974,N_14019,N_13546);
and UO_975 (O_975,N_14355,N_14555);
or UO_976 (O_976,N_14840,N_14992);
nor UO_977 (O_977,N_14526,N_14350);
xnor UO_978 (O_978,N_14187,N_14634);
nand UO_979 (O_979,N_14810,N_14717);
or UO_980 (O_980,N_13677,N_14550);
or UO_981 (O_981,N_13764,N_14159);
or UO_982 (O_982,N_14966,N_14660);
nand UO_983 (O_983,N_14216,N_13877);
or UO_984 (O_984,N_14818,N_13724);
nand UO_985 (O_985,N_13688,N_13619);
nor UO_986 (O_986,N_13635,N_14179);
nor UO_987 (O_987,N_14065,N_14672);
xor UO_988 (O_988,N_14081,N_14340);
and UO_989 (O_989,N_13844,N_14439);
xor UO_990 (O_990,N_14901,N_14801);
or UO_991 (O_991,N_14136,N_14503);
and UO_992 (O_992,N_14810,N_14536);
or UO_993 (O_993,N_14216,N_14160);
nand UO_994 (O_994,N_14230,N_14413);
nand UO_995 (O_995,N_13894,N_14027);
nand UO_996 (O_996,N_14416,N_14068);
nor UO_997 (O_997,N_13833,N_13894);
nand UO_998 (O_998,N_13632,N_14400);
xnor UO_999 (O_999,N_14216,N_14961);
and UO_1000 (O_1000,N_14730,N_14472);
nand UO_1001 (O_1001,N_13648,N_13674);
nor UO_1002 (O_1002,N_13858,N_14992);
xor UO_1003 (O_1003,N_14678,N_13542);
nand UO_1004 (O_1004,N_13764,N_14000);
and UO_1005 (O_1005,N_14368,N_14010);
nand UO_1006 (O_1006,N_14900,N_13978);
nor UO_1007 (O_1007,N_13644,N_13558);
and UO_1008 (O_1008,N_14147,N_14004);
or UO_1009 (O_1009,N_14974,N_13580);
or UO_1010 (O_1010,N_14762,N_14199);
xnor UO_1011 (O_1011,N_14527,N_14395);
nand UO_1012 (O_1012,N_13889,N_14224);
and UO_1013 (O_1013,N_13923,N_14830);
and UO_1014 (O_1014,N_14663,N_14242);
xor UO_1015 (O_1015,N_14170,N_14519);
and UO_1016 (O_1016,N_14067,N_13686);
nand UO_1017 (O_1017,N_14512,N_13738);
nand UO_1018 (O_1018,N_14741,N_13656);
nand UO_1019 (O_1019,N_14465,N_14812);
xor UO_1020 (O_1020,N_13962,N_14341);
and UO_1021 (O_1021,N_14898,N_14448);
xnor UO_1022 (O_1022,N_13653,N_13878);
and UO_1023 (O_1023,N_14989,N_13657);
nor UO_1024 (O_1024,N_14391,N_14826);
or UO_1025 (O_1025,N_13641,N_14658);
and UO_1026 (O_1026,N_13988,N_13778);
or UO_1027 (O_1027,N_13842,N_14401);
nor UO_1028 (O_1028,N_13765,N_13507);
or UO_1029 (O_1029,N_14068,N_14794);
and UO_1030 (O_1030,N_14716,N_14460);
xnor UO_1031 (O_1031,N_13954,N_14510);
xor UO_1032 (O_1032,N_14702,N_14400);
and UO_1033 (O_1033,N_13512,N_14474);
or UO_1034 (O_1034,N_14253,N_14423);
or UO_1035 (O_1035,N_14621,N_14313);
or UO_1036 (O_1036,N_14350,N_13881);
or UO_1037 (O_1037,N_14928,N_13716);
and UO_1038 (O_1038,N_14978,N_14562);
nor UO_1039 (O_1039,N_13782,N_14539);
or UO_1040 (O_1040,N_14007,N_14268);
and UO_1041 (O_1041,N_13528,N_14864);
xor UO_1042 (O_1042,N_14104,N_14124);
nand UO_1043 (O_1043,N_14496,N_13506);
xor UO_1044 (O_1044,N_14550,N_14849);
and UO_1045 (O_1045,N_14159,N_13552);
xnor UO_1046 (O_1046,N_14805,N_14008);
nor UO_1047 (O_1047,N_14864,N_14790);
and UO_1048 (O_1048,N_14914,N_14809);
nand UO_1049 (O_1049,N_14978,N_14551);
nand UO_1050 (O_1050,N_13602,N_14913);
nor UO_1051 (O_1051,N_13860,N_13704);
nor UO_1052 (O_1052,N_13907,N_14952);
or UO_1053 (O_1053,N_13917,N_14870);
nor UO_1054 (O_1054,N_13754,N_14852);
xnor UO_1055 (O_1055,N_14204,N_14965);
and UO_1056 (O_1056,N_14049,N_14127);
nand UO_1057 (O_1057,N_14584,N_13726);
or UO_1058 (O_1058,N_14741,N_14910);
xor UO_1059 (O_1059,N_14754,N_14348);
nand UO_1060 (O_1060,N_14600,N_14044);
xnor UO_1061 (O_1061,N_14000,N_13559);
nand UO_1062 (O_1062,N_14934,N_14981);
or UO_1063 (O_1063,N_14099,N_13804);
nor UO_1064 (O_1064,N_13723,N_13990);
nand UO_1065 (O_1065,N_14469,N_14620);
or UO_1066 (O_1066,N_14288,N_14409);
nand UO_1067 (O_1067,N_14868,N_14396);
and UO_1068 (O_1068,N_13983,N_13771);
nand UO_1069 (O_1069,N_14090,N_14097);
and UO_1070 (O_1070,N_14634,N_14320);
xor UO_1071 (O_1071,N_13553,N_14548);
or UO_1072 (O_1072,N_14862,N_14453);
nand UO_1073 (O_1073,N_14854,N_13894);
or UO_1074 (O_1074,N_14000,N_14620);
and UO_1075 (O_1075,N_14667,N_14082);
and UO_1076 (O_1076,N_14827,N_13616);
or UO_1077 (O_1077,N_14889,N_14122);
or UO_1078 (O_1078,N_14696,N_13684);
nand UO_1079 (O_1079,N_14677,N_13879);
or UO_1080 (O_1080,N_14014,N_14667);
xor UO_1081 (O_1081,N_14062,N_14060);
xor UO_1082 (O_1082,N_14857,N_14992);
nor UO_1083 (O_1083,N_14514,N_14583);
nor UO_1084 (O_1084,N_13722,N_14595);
xor UO_1085 (O_1085,N_14825,N_14093);
xor UO_1086 (O_1086,N_14856,N_13748);
or UO_1087 (O_1087,N_14380,N_13522);
or UO_1088 (O_1088,N_13701,N_14323);
and UO_1089 (O_1089,N_14681,N_14789);
and UO_1090 (O_1090,N_14242,N_14009);
or UO_1091 (O_1091,N_14411,N_14656);
nand UO_1092 (O_1092,N_13609,N_14922);
nand UO_1093 (O_1093,N_14048,N_14995);
and UO_1094 (O_1094,N_14378,N_14596);
nand UO_1095 (O_1095,N_14885,N_14738);
nor UO_1096 (O_1096,N_14423,N_13959);
or UO_1097 (O_1097,N_14306,N_13535);
xnor UO_1098 (O_1098,N_14921,N_14689);
nor UO_1099 (O_1099,N_14347,N_14741);
nor UO_1100 (O_1100,N_14945,N_14033);
nor UO_1101 (O_1101,N_13685,N_13571);
and UO_1102 (O_1102,N_14044,N_14380);
nand UO_1103 (O_1103,N_14032,N_14687);
xnor UO_1104 (O_1104,N_14674,N_14298);
and UO_1105 (O_1105,N_14746,N_14571);
nor UO_1106 (O_1106,N_13595,N_14600);
nor UO_1107 (O_1107,N_14335,N_13993);
and UO_1108 (O_1108,N_14837,N_13995);
or UO_1109 (O_1109,N_13509,N_14959);
or UO_1110 (O_1110,N_13696,N_14754);
and UO_1111 (O_1111,N_13764,N_14272);
and UO_1112 (O_1112,N_13749,N_14124);
and UO_1113 (O_1113,N_14074,N_14923);
xor UO_1114 (O_1114,N_14852,N_14671);
nor UO_1115 (O_1115,N_13822,N_13502);
nor UO_1116 (O_1116,N_13752,N_14047);
xnor UO_1117 (O_1117,N_14820,N_14181);
nand UO_1118 (O_1118,N_14125,N_14590);
nor UO_1119 (O_1119,N_13537,N_14530);
and UO_1120 (O_1120,N_13679,N_14046);
and UO_1121 (O_1121,N_14571,N_13619);
nand UO_1122 (O_1122,N_13809,N_13838);
nor UO_1123 (O_1123,N_14386,N_13674);
or UO_1124 (O_1124,N_14613,N_14713);
or UO_1125 (O_1125,N_13696,N_13646);
and UO_1126 (O_1126,N_14982,N_14283);
nor UO_1127 (O_1127,N_13624,N_14994);
nand UO_1128 (O_1128,N_14038,N_14717);
nand UO_1129 (O_1129,N_13874,N_14140);
xor UO_1130 (O_1130,N_14301,N_14507);
and UO_1131 (O_1131,N_14797,N_14000);
and UO_1132 (O_1132,N_13792,N_13556);
and UO_1133 (O_1133,N_14625,N_14548);
nor UO_1134 (O_1134,N_13927,N_14493);
or UO_1135 (O_1135,N_14414,N_13889);
or UO_1136 (O_1136,N_13657,N_13918);
xnor UO_1137 (O_1137,N_14340,N_14024);
and UO_1138 (O_1138,N_14634,N_13574);
nand UO_1139 (O_1139,N_14895,N_14678);
nand UO_1140 (O_1140,N_14404,N_13723);
or UO_1141 (O_1141,N_14132,N_14984);
and UO_1142 (O_1142,N_14810,N_14829);
nor UO_1143 (O_1143,N_14950,N_14168);
nand UO_1144 (O_1144,N_14022,N_14097);
nand UO_1145 (O_1145,N_14894,N_14985);
nand UO_1146 (O_1146,N_14459,N_13807);
xor UO_1147 (O_1147,N_14471,N_13586);
nand UO_1148 (O_1148,N_14082,N_14270);
or UO_1149 (O_1149,N_14602,N_14055);
nand UO_1150 (O_1150,N_13900,N_14730);
and UO_1151 (O_1151,N_14288,N_14028);
nor UO_1152 (O_1152,N_13917,N_14060);
xor UO_1153 (O_1153,N_14981,N_13928);
or UO_1154 (O_1154,N_14300,N_13625);
nor UO_1155 (O_1155,N_14617,N_13522);
xor UO_1156 (O_1156,N_14059,N_14494);
and UO_1157 (O_1157,N_13516,N_14261);
nand UO_1158 (O_1158,N_14871,N_13623);
or UO_1159 (O_1159,N_13742,N_14996);
xnor UO_1160 (O_1160,N_14478,N_14096);
nor UO_1161 (O_1161,N_14662,N_14573);
and UO_1162 (O_1162,N_14682,N_13707);
xnor UO_1163 (O_1163,N_14383,N_14186);
or UO_1164 (O_1164,N_14443,N_14007);
xor UO_1165 (O_1165,N_14470,N_14409);
xnor UO_1166 (O_1166,N_14794,N_13970);
and UO_1167 (O_1167,N_14210,N_13927);
and UO_1168 (O_1168,N_13943,N_14323);
xor UO_1169 (O_1169,N_14820,N_13828);
or UO_1170 (O_1170,N_14010,N_13841);
or UO_1171 (O_1171,N_14210,N_13569);
nor UO_1172 (O_1172,N_13526,N_14094);
or UO_1173 (O_1173,N_13734,N_13751);
nand UO_1174 (O_1174,N_14450,N_14652);
xor UO_1175 (O_1175,N_13750,N_14856);
nand UO_1176 (O_1176,N_14725,N_13561);
nor UO_1177 (O_1177,N_14823,N_14635);
nand UO_1178 (O_1178,N_13831,N_14906);
nor UO_1179 (O_1179,N_13636,N_14882);
xor UO_1180 (O_1180,N_13733,N_14871);
or UO_1181 (O_1181,N_13984,N_13936);
nand UO_1182 (O_1182,N_14842,N_14037);
nor UO_1183 (O_1183,N_14684,N_14172);
nand UO_1184 (O_1184,N_14614,N_14792);
or UO_1185 (O_1185,N_14874,N_13809);
and UO_1186 (O_1186,N_14878,N_14048);
and UO_1187 (O_1187,N_14806,N_13909);
nand UO_1188 (O_1188,N_14050,N_14262);
nand UO_1189 (O_1189,N_14781,N_14221);
xor UO_1190 (O_1190,N_14405,N_14216);
nor UO_1191 (O_1191,N_13994,N_14340);
and UO_1192 (O_1192,N_14500,N_13538);
nand UO_1193 (O_1193,N_14228,N_13519);
and UO_1194 (O_1194,N_14233,N_14969);
and UO_1195 (O_1195,N_14360,N_14815);
nand UO_1196 (O_1196,N_14588,N_14171);
xor UO_1197 (O_1197,N_14128,N_14147);
xor UO_1198 (O_1198,N_13993,N_14231);
or UO_1199 (O_1199,N_14476,N_14602);
and UO_1200 (O_1200,N_14348,N_14271);
nor UO_1201 (O_1201,N_13945,N_14346);
nor UO_1202 (O_1202,N_14474,N_13830);
nand UO_1203 (O_1203,N_13633,N_14211);
and UO_1204 (O_1204,N_14666,N_14442);
nor UO_1205 (O_1205,N_14951,N_14261);
nand UO_1206 (O_1206,N_14605,N_14437);
and UO_1207 (O_1207,N_14698,N_14399);
and UO_1208 (O_1208,N_14707,N_13528);
xnor UO_1209 (O_1209,N_14000,N_13756);
nand UO_1210 (O_1210,N_13954,N_13717);
or UO_1211 (O_1211,N_13679,N_13847);
nand UO_1212 (O_1212,N_14374,N_14476);
or UO_1213 (O_1213,N_14611,N_14293);
nor UO_1214 (O_1214,N_13555,N_14079);
nand UO_1215 (O_1215,N_14421,N_14791);
xnor UO_1216 (O_1216,N_14992,N_14547);
nand UO_1217 (O_1217,N_14478,N_14351);
and UO_1218 (O_1218,N_13933,N_13652);
and UO_1219 (O_1219,N_14308,N_14265);
and UO_1220 (O_1220,N_14890,N_14187);
and UO_1221 (O_1221,N_14851,N_14262);
nand UO_1222 (O_1222,N_13968,N_13697);
xnor UO_1223 (O_1223,N_13658,N_14040);
nand UO_1224 (O_1224,N_14515,N_14301);
or UO_1225 (O_1225,N_14976,N_14875);
nor UO_1226 (O_1226,N_13652,N_14461);
nor UO_1227 (O_1227,N_13580,N_14857);
nor UO_1228 (O_1228,N_14501,N_13844);
or UO_1229 (O_1229,N_14396,N_13523);
and UO_1230 (O_1230,N_13617,N_14426);
or UO_1231 (O_1231,N_13662,N_14979);
xor UO_1232 (O_1232,N_13740,N_14470);
and UO_1233 (O_1233,N_14414,N_13776);
and UO_1234 (O_1234,N_14790,N_14522);
or UO_1235 (O_1235,N_13755,N_13588);
and UO_1236 (O_1236,N_14340,N_14756);
nand UO_1237 (O_1237,N_14570,N_14771);
xor UO_1238 (O_1238,N_14525,N_13689);
or UO_1239 (O_1239,N_14418,N_14849);
xor UO_1240 (O_1240,N_14232,N_14264);
or UO_1241 (O_1241,N_13946,N_14684);
or UO_1242 (O_1242,N_14088,N_13848);
or UO_1243 (O_1243,N_14021,N_14503);
or UO_1244 (O_1244,N_14251,N_13551);
nor UO_1245 (O_1245,N_14644,N_13527);
xnor UO_1246 (O_1246,N_13699,N_14169);
and UO_1247 (O_1247,N_13704,N_14402);
nand UO_1248 (O_1248,N_14359,N_14087);
xnor UO_1249 (O_1249,N_14416,N_14214);
nand UO_1250 (O_1250,N_14065,N_14957);
nand UO_1251 (O_1251,N_13688,N_14153);
and UO_1252 (O_1252,N_14239,N_14234);
xor UO_1253 (O_1253,N_14245,N_13944);
nand UO_1254 (O_1254,N_14356,N_14202);
xor UO_1255 (O_1255,N_13730,N_13785);
nor UO_1256 (O_1256,N_14738,N_14534);
nand UO_1257 (O_1257,N_14943,N_14330);
nor UO_1258 (O_1258,N_13882,N_14718);
nand UO_1259 (O_1259,N_13826,N_13774);
nand UO_1260 (O_1260,N_14293,N_14944);
nand UO_1261 (O_1261,N_14374,N_13527);
nand UO_1262 (O_1262,N_14446,N_13575);
and UO_1263 (O_1263,N_14543,N_14498);
and UO_1264 (O_1264,N_13803,N_14655);
nor UO_1265 (O_1265,N_13896,N_14092);
nor UO_1266 (O_1266,N_14008,N_14385);
nor UO_1267 (O_1267,N_13708,N_14459);
nand UO_1268 (O_1268,N_14609,N_13539);
xnor UO_1269 (O_1269,N_13877,N_13565);
xor UO_1270 (O_1270,N_13597,N_13853);
nor UO_1271 (O_1271,N_13553,N_13989);
nand UO_1272 (O_1272,N_14216,N_13915);
nor UO_1273 (O_1273,N_14445,N_14997);
nand UO_1274 (O_1274,N_14433,N_14350);
nand UO_1275 (O_1275,N_13506,N_14604);
xor UO_1276 (O_1276,N_13649,N_13552);
or UO_1277 (O_1277,N_13942,N_14811);
and UO_1278 (O_1278,N_13712,N_14938);
nor UO_1279 (O_1279,N_14882,N_14499);
and UO_1280 (O_1280,N_13960,N_14981);
nand UO_1281 (O_1281,N_13632,N_13679);
and UO_1282 (O_1282,N_14053,N_14096);
and UO_1283 (O_1283,N_14198,N_13587);
nor UO_1284 (O_1284,N_14897,N_14316);
nand UO_1285 (O_1285,N_14996,N_13971);
and UO_1286 (O_1286,N_14922,N_14764);
and UO_1287 (O_1287,N_14278,N_13706);
nand UO_1288 (O_1288,N_14947,N_14238);
xor UO_1289 (O_1289,N_13937,N_14838);
or UO_1290 (O_1290,N_14713,N_13511);
nand UO_1291 (O_1291,N_14272,N_13709);
or UO_1292 (O_1292,N_14066,N_13561);
nand UO_1293 (O_1293,N_14387,N_14592);
and UO_1294 (O_1294,N_13537,N_14339);
xor UO_1295 (O_1295,N_14541,N_14011);
xnor UO_1296 (O_1296,N_14920,N_14970);
and UO_1297 (O_1297,N_13550,N_13924);
and UO_1298 (O_1298,N_14295,N_13930);
nor UO_1299 (O_1299,N_14831,N_14120);
and UO_1300 (O_1300,N_13705,N_13510);
nor UO_1301 (O_1301,N_13532,N_13687);
nand UO_1302 (O_1302,N_14455,N_14548);
nand UO_1303 (O_1303,N_14446,N_14199);
nand UO_1304 (O_1304,N_14235,N_13800);
nor UO_1305 (O_1305,N_14537,N_14224);
nor UO_1306 (O_1306,N_13578,N_14917);
nand UO_1307 (O_1307,N_14935,N_14771);
or UO_1308 (O_1308,N_14287,N_14213);
nor UO_1309 (O_1309,N_14093,N_14920);
nor UO_1310 (O_1310,N_14615,N_14601);
xnor UO_1311 (O_1311,N_14043,N_14502);
and UO_1312 (O_1312,N_14193,N_13849);
xor UO_1313 (O_1313,N_14152,N_14989);
xor UO_1314 (O_1314,N_14815,N_14973);
nand UO_1315 (O_1315,N_13984,N_13574);
nand UO_1316 (O_1316,N_14891,N_14769);
nand UO_1317 (O_1317,N_13964,N_13615);
nor UO_1318 (O_1318,N_13890,N_14072);
or UO_1319 (O_1319,N_14824,N_14749);
or UO_1320 (O_1320,N_13850,N_13599);
xor UO_1321 (O_1321,N_14918,N_14453);
nor UO_1322 (O_1322,N_13580,N_14107);
xnor UO_1323 (O_1323,N_14404,N_14528);
nand UO_1324 (O_1324,N_14956,N_13752);
or UO_1325 (O_1325,N_14193,N_13514);
xor UO_1326 (O_1326,N_14556,N_14783);
and UO_1327 (O_1327,N_14952,N_14381);
and UO_1328 (O_1328,N_14176,N_14405);
or UO_1329 (O_1329,N_14138,N_13846);
or UO_1330 (O_1330,N_13673,N_14273);
xor UO_1331 (O_1331,N_14054,N_14159);
nand UO_1332 (O_1332,N_13747,N_13509);
nand UO_1333 (O_1333,N_13553,N_13703);
nand UO_1334 (O_1334,N_14887,N_14384);
nor UO_1335 (O_1335,N_14395,N_13869);
xor UO_1336 (O_1336,N_14842,N_14282);
nand UO_1337 (O_1337,N_13820,N_13528);
and UO_1338 (O_1338,N_14688,N_14984);
nor UO_1339 (O_1339,N_14793,N_14127);
and UO_1340 (O_1340,N_13822,N_13911);
nand UO_1341 (O_1341,N_14991,N_14386);
xnor UO_1342 (O_1342,N_14389,N_14748);
nor UO_1343 (O_1343,N_14027,N_14050);
nor UO_1344 (O_1344,N_14982,N_13632);
and UO_1345 (O_1345,N_13582,N_14589);
or UO_1346 (O_1346,N_13839,N_13886);
nand UO_1347 (O_1347,N_13701,N_13559);
xor UO_1348 (O_1348,N_14609,N_14415);
nand UO_1349 (O_1349,N_13930,N_14699);
xnor UO_1350 (O_1350,N_13581,N_14391);
or UO_1351 (O_1351,N_14709,N_14673);
or UO_1352 (O_1352,N_14300,N_14256);
or UO_1353 (O_1353,N_14538,N_14830);
or UO_1354 (O_1354,N_13687,N_13770);
and UO_1355 (O_1355,N_13849,N_14517);
or UO_1356 (O_1356,N_13527,N_14838);
nand UO_1357 (O_1357,N_13635,N_13970);
and UO_1358 (O_1358,N_14916,N_14322);
nand UO_1359 (O_1359,N_13711,N_13607);
nand UO_1360 (O_1360,N_14482,N_13509);
nor UO_1361 (O_1361,N_14965,N_13666);
nand UO_1362 (O_1362,N_14241,N_13633);
and UO_1363 (O_1363,N_14993,N_13971);
xnor UO_1364 (O_1364,N_13958,N_14725);
and UO_1365 (O_1365,N_14541,N_14390);
nand UO_1366 (O_1366,N_13571,N_14189);
nand UO_1367 (O_1367,N_13741,N_13792);
nor UO_1368 (O_1368,N_14721,N_14409);
nand UO_1369 (O_1369,N_14089,N_14441);
xnor UO_1370 (O_1370,N_14488,N_13522);
nor UO_1371 (O_1371,N_14453,N_14788);
xnor UO_1372 (O_1372,N_14191,N_14118);
nor UO_1373 (O_1373,N_14857,N_14828);
or UO_1374 (O_1374,N_14265,N_13656);
nor UO_1375 (O_1375,N_13982,N_14690);
nand UO_1376 (O_1376,N_13711,N_13631);
xor UO_1377 (O_1377,N_14233,N_13869);
nor UO_1378 (O_1378,N_13709,N_13759);
nor UO_1379 (O_1379,N_14656,N_14365);
nor UO_1380 (O_1380,N_14932,N_13701);
or UO_1381 (O_1381,N_13817,N_14503);
xor UO_1382 (O_1382,N_13892,N_13887);
nor UO_1383 (O_1383,N_14297,N_13740);
nor UO_1384 (O_1384,N_14564,N_14131);
and UO_1385 (O_1385,N_13756,N_13855);
nand UO_1386 (O_1386,N_14132,N_14091);
nor UO_1387 (O_1387,N_14636,N_13512);
or UO_1388 (O_1388,N_14277,N_14889);
or UO_1389 (O_1389,N_14301,N_13652);
or UO_1390 (O_1390,N_13885,N_13924);
nor UO_1391 (O_1391,N_13906,N_14614);
nand UO_1392 (O_1392,N_14586,N_13626);
nand UO_1393 (O_1393,N_13916,N_14637);
nand UO_1394 (O_1394,N_13885,N_14899);
and UO_1395 (O_1395,N_14375,N_13617);
or UO_1396 (O_1396,N_14110,N_13679);
or UO_1397 (O_1397,N_13793,N_14081);
and UO_1398 (O_1398,N_14572,N_13708);
nand UO_1399 (O_1399,N_13965,N_14100);
or UO_1400 (O_1400,N_13918,N_14886);
nand UO_1401 (O_1401,N_14267,N_14669);
nand UO_1402 (O_1402,N_13908,N_13912);
nor UO_1403 (O_1403,N_14162,N_13524);
xor UO_1404 (O_1404,N_13792,N_14098);
nor UO_1405 (O_1405,N_14259,N_14115);
or UO_1406 (O_1406,N_13813,N_13693);
xor UO_1407 (O_1407,N_13508,N_14316);
and UO_1408 (O_1408,N_13810,N_14287);
xnor UO_1409 (O_1409,N_13633,N_13736);
nor UO_1410 (O_1410,N_13774,N_14637);
nor UO_1411 (O_1411,N_14118,N_14398);
xor UO_1412 (O_1412,N_14321,N_14833);
xor UO_1413 (O_1413,N_14319,N_14301);
or UO_1414 (O_1414,N_14209,N_13693);
nand UO_1415 (O_1415,N_14755,N_14434);
or UO_1416 (O_1416,N_13711,N_14596);
nor UO_1417 (O_1417,N_14460,N_14900);
nand UO_1418 (O_1418,N_14120,N_13923);
or UO_1419 (O_1419,N_14168,N_14740);
xnor UO_1420 (O_1420,N_14475,N_14836);
nand UO_1421 (O_1421,N_14329,N_13881);
nand UO_1422 (O_1422,N_13813,N_14563);
and UO_1423 (O_1423,N_14917,N_13889);
or UO_1424 (O_1424,N_14287,N_14334);
and UO_1425 (O_1425,N_13708,N_13882);
and UO_1426 (O_1426,N_14294,N_13537);
or UO_1427 (O_1427,N_13910,N_13592);
nand UO_1428 (O_1428,N_14371,N_14434);
xnor UO_1429 (O_1429,N_14792,N_14567);
nor UO_1430 (O_1430,N_14478,N_14197);
nor UO_1431 (O_1431,N_14673,N_14293);
and UO_1432 (O_1432,N_14907,N_14007);
nor UO_1433 (O_1433,N_14916,N_14887);
xor UO_1434 (O_1434,N_13972,N_14245);
nand UO_1435 (O_1435,N_13906,N_14250);
nor UO_1436 (O_1436,N_13859,N_14505);
or UO_1437 (O_1437,N_13916,N_13678);
or UO_1438 (O_1438,N_14688,N_14612);
or UO_1439 (O_1439,N_13933,N_13582);
or UO_1440 (O_1440,N_14734,N_13766);
nand UO_1441 (O_1441,N_14491,N_14517);
nor UO_1442 (O_1442,N_14010,N_14707);
xnor UO_1443 (O_1443,N_14127,N_14161);
and UO_1444 (O_1444,N_13541,N_14119);
or UO_1445 (O_1445,N_14686,N_14114);
nand UO_1446 (O_1446,N_14248,N_14584);
or UO_1447 (O_1447,N_13521,N_14272);
xor UO_1448 (O_1448,N_14603,N_13962);
xor UO_1449 (O_1449,N_14927,N_14547);
or UO_1450 (O_1450,N_13512,N_13670);
or UO_1451 (O_1451,N_14416,N_13623);
nand UO_1452 (O_1452,N_14323,N_14948);
nand UO_1453 (O_1453,N_14441,N_13634);
and UO_1454 (O_1454,N_13666,N_14356);
or UO_1455 (O_1455,N_14608,N_14525);
nor UO_1456 (O_1456,N_14134,N_14678);
nand UO_1457 (O_1457,N_14445,N_13648);
or UO_1458 (O_1458,N_13599,N_14068);
and UO_1459 (O_1459,N_14458,N_14352);
and UO_1460 (O_1460,N_13590,N_14365);
xor UO_1461 (O_1461,N_14379,N_14293);
nand UO_1462 (O_1462,N_14515,N_14575);
and UO_1463 (O_1463,N_13896,N_14936);
and UO_1464 (O_1464,N_14984,N_13522);
or UO_1465 (O_1465,N_14716,N_14063);
or UO_1466 (O_1466,N_14135,N_13788);
nand UO_1467 (O_1467,N_13718,N_13762);
nor UO_1468 (O_1468,N_13686,N_14793);
nor UO_1469 (O_1469,N_14099,N_14849);
and UO_1470 (O_1470,N_13781,N_14738);
nand UO_1471 (O_1471,N_13729,N_14760);
nand UO_1472 (O_1472,N_14215,N_14356);
or UO_1473 (O_1473,N_14816,N_14891);
xnor UO_1474 (O_1474,N_14118,N_13835);
and UO_1475 (O_1475,N_14308,N_14895);
nor UO_1476 (O_1476,N_13572,N_14698);
xnor UO_1477 (O_1477,N_14916,N_13665);
nand UO_1478 (O_1478,N_13650,N_14727);
or UO_1479 (O_1479,N_14367,N_14569);
nand UO_1480 (O_1480,N_14206,N_13940);
xor UO_1481 (O_1481,N_14650,N_14883);
nand UO_1482 (O_1482,N_14376,N_14705);
nand UO_1483 (O_1483,N_14538,N_13777);
or UO_1484 (O_1484,N_14187,N_14215);
xnor UO_1485 (O_1485,N_13592,N_13633);
nor UO_1486 (O_1486,N_14702,N_13567);
nand UO_1487 (O_1487,N_14380,N_13889);
nand UO_1488 (O_1488,N_13828,N_14856);
nand UO_1489 (O_1489,N_14990,N_13837);
and UO_1490 (O_1490,N_13751,N_14346);
or UO_1491 (O_1491,N_14320,N_13726);
nand UO_1492 (O_1492,N_13900,N_14209);
or UO_1493 (O_1493,N_14677,N_14603);
xor UO_1494 (O_1494,N_14839,N_14998);
nand UO_1495 (O_1495,N_14361,N_13708);
nand UO_1496 (O_1496,N_13769,N_13587);
and UO_1497 (O_1497,N_13532,N_14374);
nor UO_1498 (O_1498,N_13536,N_14981);
xnor UO_1499 (O_1499,N_14442,N_13761);
or UO_1500 (O_1500,N_14039,N_13974);
xor UO_1501 (O_1501,N_14045,N_14143);
nand UO_1502 (O_1502,N_14777,N_14221);
nor UO_1503 (O_1503,N_14842,N_14066);
nor UO_1504 (O_1504,N_14292,N_14325);
or UO_1505 (O_1505,N_14228,N_14306);
xnor UO_1506 (O_1506,N_13968,N_14396);
or UO_1507 (O_1507,N_14114,N_14048);
xnor UO_1508 (O_1508,N_14667,N_13821);
nor UO_1509 (O_1509,N_14445,N_13977);
and UO_1510 (O_1510,N_13653,N_14776);
and UO_1511 (O_1511,N_14715,N_13958);
nand UO_1512 (O_1512,N_13517,N_14138);
or UO_1513 (O_1513,N_14918,N_13856);
nor UO_1514 (O_1514,N_13555,N_14228);
nor UO_1515 (O_1515,N_13964,N_14840);
xor UO_1516 (O_1516,N_14813,N_14223);
and UO_1517 (O_1517,N_14860,N_14269);
nor UO_1518 (O_1518,N_14465,N_13803);
nor UO_1519 (O_1519,N_13825,N_14723);
nor UO_1520 (O_1520,N_14790,N_13790);
nor UO_1521 (O_1521,N_14834,N_13978);
and UO_1522 (O_1522,N_14716,N_14891);
and UO_1523 (O_1523,N_13902,N_13635);
nand UO_1524 (O_1524,N_13637,N_13906);
nand UO_1525 (O_1525,N_14842,N_13853);
nand UO_1526 (O_1526,N_13800,N_13860);
and UO_1527 (O_1527,N_14647,N_13635);
and UO_1528 (O_1528,N_14222,N_14145);
and UO_1529 (O_1529,N_14706,N_14952);
and UO_1530 (O_1530,N_13698,N_14208);
nor UO_1531 (O_1531,N_13751,N_14522);
nand UO_1532 (O_1532,N_14749,N_14996);
xnor UO_1533 (O_1533,N_13760,N_14131);
and UO_1534 (O_1534,N_14881,N_13865);
nor UO_1535 (O_1535,N_13852,N_13909);
and UO_1536 (O_1536,N_13618,N_13799);
xnor UO_1537 (O_1537,N_14684,N_14532);
or UO_1538 (O_1538,N_14794,N_14034);
nand UO_1539 (O_1539,N_13902,N_14288);
nor UO_1540 (O_1540,N_13641,N_13884);
and UO_1541 (O_1541,N_14627,N_13942);
nor UO_1542 (O_1542,N_13603,N_14419);
nand UO_1543 (O_1543,N_14668,N_14297);
xor UO_1544 (O_1544,N_14600,N_14628);
xor UO_1545 (O_1545,N_14229,N_13605);
and UO_1546 (O_1546,N_14199,N_13586);
nor UO_1547 (O_1547,N_13852,N_14527);
xnor UO_1548 (O_1548,N_14932,N_14698);
and UO_1549 (O_1549,N_13754,N_14261);
xnor UO_1550 (O_1550,N_14412,N_13961);
xor UO_1551 (O_1551,N_14107,N_14137);
nor UO_1552 (O_1552,N_13612,N_14598);
or UO_1553 (O_1553,N_14342,N_14816);
and UO_1554 (O_1554,N_13815,N_13700);
nand UO_1555 (O_1555,N_14021,N_14758);
nand UO_1556 (O_1556,N_13770,N_14466);
nand UO_1557 (O_1557,N_14731,N_14658);
xor UO_1558 (O_1558,N_14571,N_14802);
and UO_1559 (O_1559,N_14829,N_14678);
nand UO_1560 (O_1560,N_13702,N_13790);
xnor UO_1561 (O_1561,N_14792,N_13990);
nand UO_1562 (O_1562,N_13968,N_13796);
nor UO_1563 (O_1563,N_14247,N_13652);
xnor UO_1564 (O_1564,N_14122,N_14610);
xnor UO_1565 (O_1565,N_14760,N_14465);
xor UO_1566 (O_1566,N_13556,N_13542);
or UO_1567 (O_1567,N_14167,N_14644);
nor UO_1568 (O_1568,N_13939,N_14140);
and UO_1569 (O_1569,N_13708,N_13919);
and UO_1570 (O_1570,N_13738,N_14104);
nand UO_1571 (O_1571,N_14457,N_14654);
or UO_1572 (O_1572,N_14153,N_14557);
nand UO_1573 (O_1573,N_14791,N_14911);
nand UO_1574 (O_1574,N_14949,N_13898);
xor UO_1575 (O_1575,N_14935,N_13631);
and UO_1576 (O_1576,N_13639,N_13741);
or UO_1577 (O_1577,N_13539,N_14008);
or UO_1578 (O_1578,N_14716,N_13559);
nand UO_1579 (O_1579,N_14016,N_14189);
nand UO_1580 (O_1580,N_14195,N_13644);
or UO_1581 (O_1581,N_14996,N_14404);
or UO_1582 (O_1582,N_13592,N_14066);
nor UO_1583 (O_1583,N_14210,N_14640);
and UO_1584 (O_1584,N_14711,N_13624);
or UO_1585 (O_1585,N_14236,N_14822);
nor UO_1586 (O_1586,N_14895,N_13510);
nand UO_1587 (O_1587,N_14268,N_14378);
nand UO_1588 (O_1588,N_14322,N_14188);
nor UO_1589 (O_1589,N_13897,N_14522);
or UO_1590 (O_1590,N_14128,N_14308);
or UO_1591 (O_1591,N_13768,N_14376);
nand UO_1592 (O_1592,N_14421,N_13613);
nand UO_1593 (O_1593,N_14146,N_14246);
nand UO_1594 (O_1594,N_14254,N_14259);
nor UO_1595 (O_1595,N_14648,N_13970);
and UO_1596 (O_1596,N_13609,N_13844);
or UO_1597 (O_1597,N_13991,N_13773);
or UO_1598 (O_1598,N_14900,N_14212);
nor UO_1599 (O_1599,N_13883,N_14535);
and UO_1600 (O_1600,N_13556,N_13967);
nor UO_1601 (O_1601,N_14365,N_14363);
nor UO_1602 (O_1602,N_14436,N_14816);
xor UO_1603 (O_1603,N_13861,N_13920);
nor UO_1604 (O_1604,N_13652,N_14290);
xnor UO_1605 (O_1605,N_14959,N_14870);
nor UO_1606 (O_1606,N_14042,N_13932);
and UO_1607 (O_1607,N_13927,N_14190);
and UO_1608 (O_1608,N_13949,N_14846);
and UO_1609 (O_1609,N_14048,N_13610);
nor UO_1610 (O_1610,N_14570,N_14628);
nand UO_1611 (O_1611,N_14830,N_13939);
or UO_1612 (O_1612,N_14224,N_13870);
xor UO_1613 (O_1613,N_14433,N_14832);
and UO_1614 (O_1614,N_13578,N_14649);
xor UO_1615 (O_1615,N_14323,N_14437);
or UO_1616 (O_1616,N_13708,N_14060);
or UO_1617 (O_1617,N_14556,N_13759);
nor UO_1618 (O_1618,N_14591,N_13612);
or UO_1619 (O_1619,N_13607,N_14411);
and UO_1620 (O_1620,N_14161,N_14827);
nand UO_1621 (O_1621,N_14578,N_13699);
or UO_1622 (O_1622,N_13820,N_14201);
xnor UO_1623 (O_1623,N_14646,N_13649);
nand UO_1624 (O_1624,N_13753,N_14919);
nand UO_1625 (O_1625,N_14301,N_14736);
and UO_1626 (O_1626,N_14412,N_14409);
nand UO_1627 (O_1627,N_14254,N_14008);
or UO_1628 (O_1628,N_14577,N_14194);
nor UO_1629 (O_1629,N_14540,N_14777);
or UO_1630 (O_1630,N_13914,N_14797);
nor UO_1631 (O_1631,N_14920,N_13907);
and UO_1632 (O_1632,N_14060,N_14923);
nor UO_1633 (O_1633,N_14418,N_14581);
or UO_1634 (O_1634,N_13606,N_14955);
and UO_1635 (O_1635,N_14930,N_13514);
or UO_1636 (O_1636,N_14005,N_14826);
and UO_1637 (O_1637,N_13754,N_14796);
nand UO_1638 (O_1638,N_14722,N_13588);
nand UO_1639 (O_1639,N_14882,N_14715);
nand UO_1640 (O_1640,N_13575,N_13755);
nand UO_1641 (O_1641,N_14940,N_14201);
or UO_1642 (O_1642,N_13709,N_13919);
xnor UO_1643 (O_1643,N_13544,N_14118);
nand UO_1644 (O_1644,N_14447,N_13557);
nor UO_1645 (O_1645,N_14310,N_14809);
nand UO_1646 (O_1646,N_13741,N_13609);
nor UO_1647 (O_1647,N_13741,N_14596);
nand UO_1648 (O_1648,N_13861,N_14865);
xnor UO_1649 (O_1649,N_14495,N_13655);
nand UO_1650 (O_1650,N_14754,N_14545);
nand UO_1651 (O_1651,N_13821,N_13536);
nand UO_1652 (O_1652,N_14759,N_14323);
and UO_1653 (O_1653,N_13696,N_14076);
nand UO_1654 (O_1654,N_13637,N_14999);
nor UO_1655 (O_1655,N_13904,N_14915);
nor UO_1656 (O_1656,N_14963,N_13867);
nor UO_1657 (O_1657,N_14692,N_14948);
or UO_1658 (O_1658,N_14947,N_14106);
nand UO_1659 (O_1659,N_14078,N_13555);
nand UO_1660 (O_1660,N_14246,N_13923);
and UO_1661 (O_1661,N_14198,N_13785);
and UO_1662 (O_1662,N_14392,N_13997);
nand UO_1663 (O_1663,N_14277,N_14832);
or UO_1664 (O_1664,N_13856,N_13918);
nor UO_1665 (O_1665,N_13937,N_13950);
or UO_1666 (O_1666,N_14765,N_14646);
nand UO_1667 (O_1667,N_14987,N_14297);
nand UO_1668 (O_1668,N_13920,N_14865);
xnor UO_1669 (O_1669,N_14414,N_14593);
and UO_1670 (O_1670,N_13626,N_14075);
or UO_1671 (O_1671,N_14639,N_14329);
or UO_1672 (O_1672,N_14658,N_14873);
or UO_1673 (O_1673,N_14141,N_14475);
nand UO_1674 (O_1674,N_13776,N_13630);
and UO_1675 (O_1675,N_14318,N_13690);
or UO_1676 (O_1676,N_13597,N_14139);
xor UO_1677 (O_1677,N_13760,N_13792);
nand UO_1678 (O_1678,N_13549,N_14219);
or UO_1679 (O_1679,N_13551,N_14976);
or UO_1680 (O_1680,N_14582,N_14112);
xor UO_1681 (O_1681,N_14009,N_14900);
and UO_1682 (O_1682,N_13719,N_14799);
or UO_1683 (O_1683,N_13829,N_13932);
or UO_1684 (O_1684,N_14336,N_13654);
xor UO_1685 (O_1685,N_14957,N_13807);
and UO_1686 (O_1686,N_14594,N_13584);
nand UO_1687 (O_1687,N_13952,N_14753);
nand UO_1688 (O_1688,N_14272,N_14982);
and UO_1689 (O_1689,N_14361,N_14544);
nand UO_1690 (O_1690,N_14534,N_13884);
or UO_1691 (O_1691,N_13708,N_14504);
or UO_1692 (O_1692,N_14743,N_14372);
nand UO_1693 (O_1693,N_14257,N_14856);
nand UO_1694 (O_1694,N_14777,N_14793);
nand UO_1695 (O_1695,N_14772,N_14648);
or UO_1696 (O_1696,N_13619,N_13872);
nand UO_1697 (O_1697,N_14954,N_14614);
nand UO_1698 (O_1698,N_14957,N_13767);
nor UO_1699 (O_1699,N_14410,N_14636);
or UO_1700 (O_1700,N_13521,N_14124);
and UO_1701 (O_1701,N_14338,N_14255);
nor UO_1702 (O_1702,N_13706,N_13517);
xor UO_1703 (O_1703,N_14521,N_14356);
or UO_1704 (O_1704,N_14046,N_13776);
and UO_1705 (O_1705,N_14548,N_13818);
and UO_1706 (O_1706,N_14790,N_14074);
xnor UO_1707 (O_1707,N_13956,N_14902);
xnor UO_1708 (O_1708,N_14681,N_14870);
nand UO_1709 (O_1709,N_14481,N_14639);
xor UO_1710 (O_1710,N_13975,N_13544);
and UO_1711 (O_1711,N_14225,N_14102);
nor UO_1712 (O_1712,N_14802,N_14751);
and UO_1713 (O_1713,N_14298,N_14292);
nor UO_1714 (O_1714,N_14795,N_14740);
nand UO_1715 (O_1715,N_14689,N_14368);
nand UO_1716 (O_1716,N_14952,N_14758);
nor UO_1717 (O_1717,N_14844,N_14565);
nand UO_1718 (O_1718,N_14210,N_14610);
nor UO_1719 (O_1719,N_14519,N_14147);
and UO_1720 (O_1720,N_14415,N_14716);
xnor UO_1721 (O_1721,N_14478,N_14898);
nor UO_1722 (O_1722,N_14910,N_14556);
or UO_1723 (O_1723,N_14693,N_14511);
and UO_1724 (O_1724,N_14658,N_13752);
nand UO_1725 (O_1725,N_13823,N_14812);
xnor UO_1726 (O_1726,N_13522,N_13767);
nor UO_1727 (O_1727,N_13681,N_14671);
or UO_1728 (O_1728,N_14074,N_14016);
xnor UO_1729 (O_1729,N_14046,N_14044);
nor UO_1730 (O_1730,N_13744,N_14739);
and UO_1731 (O_1731,N_14942,N_14070);
and UO_1732 (O_1732,N_14968,N_14320);
and UO_1733 (O_1733,N_13724,N_14637);
and UO_1734 (O_1734,N_13516,N_13628);
or UO_1735 (O_1735,N_14817,N_14930);
nand UO_1736 (O_1736,N_13927,N_14308);
nand UO_1737 (O_1737,N_14833,N_14162);
nand UO_1738 (O_1738,N_14048,N_14898);
or UO_1739 (O_1739,N_14883,N_14153);
and UO_1740 (O_1740,N_14232,N_14384);
nor UO_1741 (O_1741,N_14270,N_14517);
or UO_1742 (O_1742,N_14008,N_14930);
xnor UO_1743 (O_1743,N_14671,N_14938);
nand UO_1744 (O_1744,N_13995,N_13817);
or UO_1745 (O_1745,N_14567,N_14391);
nand UO_1746 (O_1746,N_14689,N_13679);
and UO_1747 (O_1747,N_13568,N_13749);
nor UO_1748 (O_1748,N_14395,N_13523);
xnor UO_1749 (O_1749,N_14623,N_14274);
nor UO_1750 (O_1750,N_14527,N_14528);
or UO_1751 (O_1751,N_13876,N_14094);
and UO_1752 (O_1752,N_14127,N_13854);
nand UO_1753 (O_1753,N_13624,N_14308);
or UO_1754 (O_1754,N_13602,N_14112);
nand UO_1755 (O_1755,N_13596,N_14553);
xnor UO_1756 (O_1756,N_13959,N_14849);
or UO_1757 (O_1757,N_14169,N_14466);
nand UO_1758 (O_1758,N_14653,N_14098);
nor UO_1759 (O_1759,N_14069,N_13528);
nand UO_1760 (O_1760,N_14527,N_14499);
nor UO_1761 (O_1761,N_14903,N_14356);
nand UO_1762 (O_1762,N_13703,N_13606);
nand UO_1763 (O_1763,N_13671,N_14891);
nand UO_1764 (O_1764,N_13585,N_14564);
nand UO_1765 (O_1765,N_13530,N_14059);
and UO_1766 (O_1766,N_14365,N_14459);
nand UO_1767 (O_1767,N_13767,N_14987);
and UO_1768 (O_1768,N_14787,N_13859);
or UO_1769 (O_1769,N_14984,N_14508);
or UO_1770 (O_1770,N_14430,N_14706);
xnor UO_1771 (O_1771,N_13631,N_13957);
and UO_1772 (O_1772,N_14577,N_13745);
and UO_1773 (O_1773,N_13540,N_14874);
or UO_1774 (O_1774,N_13806,N_14277);
and UO_1775 (O_1775,N_14581,N_14262);
nor UO_1776 (O_1776,N_14247,N_14406);
or UO_1777 (O_1777,N_14855,N_14748);
or UO_1778 (O_1778,N_14702,N_14229);
or UO_1779 (O_1779,N_14606,N_14396);
and UO_1780 (O_1780,N_14272,N_13971);
xor UO_1781 (O_1781,N_14734,N_14315);
or UO_1782 (O_1782,N_14443,N_13990);
xor UO_1783 (O_1783,N_14498,N_14838);
nand UO_1784 (O_1784,N_14711,N_14213);
nor UO_1785 (O_1785,N_13640,N_14509);
nand UO_1786 (O_1786,N_14000,N_13976);
or UO_1787 (O_1787,N_14619,N_13780);
and UO_1788 (O_1788,N_13581,N_13641);
or UO_1789 (O_1789,N_14060,N_14160);
nor UO_1790 (O_1790,N_14761,N_14015);
nor UO_1791 (O_1791,N_14202,N_14737);
or UO_1792 (O_1792,N_14159,N_14914);
and UO_1793 (O_1793,N_14072,N_13809);
nor UO_1794 (O_1794,N_14757,N_14136);
xnor UO_1795 (O_1795,N_14613,N_13867);
and UO_1796 (O_1796,N_13851,N_14907);
nor UO_1797 (O_1797,N_14544,N_13750);
or UO_1798 (O_1798,N_13529,N_14076);
or UO_1799 (O_1799,N_14682,N_14990);
and UO_1800 (O_1800,N_14589,N_14323);
xor UO_1801 (O_1801,N_13636,N_14323);
nor UO_1802 (O_1802,N_14528,N_13664);
and UO_1803 (O_1803,N_14999,N_14625);
or UO_1804 (O_1804,N_14494,N_13585);
nor UO_1805 (O_1805,N_13518,N_14633);
or UO_1806 (O_1806,N_14516,N_14784);
nand UO_1807 (O_1807,N_14119,N_13805);
nand UO_1808 (O_1808,N_14952,N_14825);
and UO_1809 (O_1809,N_13689,N_14970);
xnor UO_1810 (O_1810,N_14365,N_14152);
and UO_1811 (O_1811,N_14901,N_14713);
nand UO_1812 (O_1812,N_13609,N_14705);
and UO_1813 (O_1813,N_14219,N_13795);
nor UO_1814 (O_1814,N_14180,N_14062);
or UO_1815 (O_1815,N_14367,N_14241);
nor UO_1816 (O_1816,N_14854,N_13596);
xnor UO_1817 (O_1817,N_14663,N_14889);
and UO_1818 (O_1818,N_13874,N_14943);
nor UO_1819 (O_1819,N_14280,N_14555);
or UO_1820 (O_1820,N_13793,N_13873);
or UO_1821 (O_1821,N_13762,N_14666);
nor UO_1822 (O_1822,N_14440,N_14601);
xor UO_1823 (O_1823,N_14380,N_14018);
nor UO_1824 (O_1824,N_14423,N_13911);
nand UO_1825 (O_1825,N_14247,N_14076);
xor UO_1826 (O_1826,N_13659,N_14969);
and UO_1827 (O_1827,N_14443,N_14447);
and UO_1828 (O_1828,N_14489,N_14367);
nor UO_1829 (O_1829,N_14859,N_14261);
or UO_1830 (O_1830,N_13615,N_14578);
nor UO_1831 (O_1831,N_14645,N_13772);
xor UO_1832 (O_1832,N_13921,N_13621);
or UO_1833 (O_1833,N_13754,N_14959);
nor UO_1834 (O_1834,N_13868,N_14011);
and UO_1835 (O_1835,N_13917,N_14366);
and UO_1836 (O_1836,N_14599,N_14132);
nor UO_1837 (O_1837,N_14484,N_14866);
and UO_1838 (O_1838,N_14344,N_14352);
or UO_1839 (O_1839,N_13575,N_14998);
xnor UO_1840 (O_1840,N_13851,N_14383);
nor UO_1841 (O_1841,N_13821,N_13607);
nand UO_1842 (O_1842,N_13560,N_13847);
xor UO_1843 (O_1843,N_14205,N_14441);
nor UO_1844 (O_1844,N_14657,N_14438);
nor UO_1845 (O_1845,N_13639,N_14482);
xnor UO_1846 (O_1846,N_14933,N_13607);
xnor UO_1847 (O_1847,N_14883,N_13686);
nor UO_1848 (O_1848,N_13573,N_14295);
xor UO_1849 (O_1849,N_14031,N_13732);
or UO_1850 (O_1850,N_14536,N_14894);
nand UO_1851 (O_1851,N_14928,N_14158);
xnor UO_1852 (O_1852,N_13910,N_14274);
xnor UO_1853 (O_1853,N_13773,N_14509);
nor UO_1854 (O_1854,N_14263,N_14948);
nand UO_1855 (O_1855,N_14919,N_13920);
xnor UO_1856 (O_1856,N_14965,N_14342);
nand UO_1857 (O_1857,N_14485,N_14546);
nand UO_1858 (O_1858,N_14221,N_14802);
nor UO_1859 (O_1859,N_14640,N_14930);
xor UO_1860 (O_1860,N_13645,N_14001);
xnor UO_1861 (O_1861,N_14646,N_13943);
nand UO_1862 (O_1862,N_14429,N_14104);
nand UO_1863 (O_1863,N_14246,N_13679);
and UO_1864 (O_1864,N_13837,N_13750);
nor UO_1865 (O_1865,N_14532,N_13818);
xor UO_1866 (O_1866,N_14017,N_14937);
and UO_1867 (O_1867,N_13993,N_13715);
nand UO_1868 (O_1868,N_13957,N_14487);
nand UO_1869 (O_1869,N_14646,N_14126);
and UO_1870 (O_1870,N_14837,N_14180);
nand UO_1871 (O_1871,N_14551,N_14991);
nand UO_1872 (O_1872,N_13648,N_13982);
and UO_1873 (O_1873,N_14434,N_14068);
xor UO_1874 (O_1874,N_13530,N_14715);
and UO_1875 (O_1875,N_13734,N_14449);
nand UO_1876 (O_1876,N_13823,N_13565);
nor UO_1877 (O_1877,N_14599,N_14035);
nor UO_1878 (O_1878,N_13549,N_13648);
xnor UO_1879 (O_1879,N_13902,N_14528);
xor UO_1880 (O_1880,N_14930,N_14306);
and UO_1881 (O_1881,N_14935,N_14223);
nor UO_1882 (O_1882,N_14818,N_13732);
and UO_1883 (O_1883,N_13507,N_13713);
xnor UO_1884 (O_1884,N_13703,N_14692);
and UO_1885 (O_1885,N_13739,N_14472);
and UO_1886 (O_1886,N_14118,N_13520);
nand UO_1887 (O_1887,N_14854,N_14556);
nand UO_1888 (O_1888,N_14652,N_13624);
and UO_1889 (O_1889,N_13733,N_14411);
nor UO_1890 (O_1890,N_14593,N_14929);
or UO_1891 (O_1891,N_14498,N_13641);
nand UO_1892 (O_1892,N_14146,N_13795);
xnor UO_1893 (O_1893,N_13988,N_14120);
or UO_1894 (O_1894,N_14752,N_14404);
xnor UO_1895 (O_1895,N_13536,N_14296);
xor UO_1896 (O_1896,N_14700,N_14501);
or UO_1897 (O_1897,N_13548,N_13873);
nand UO_1898 (O_1898,N_14201,N_14246);
xnor UO_1899 (O_1899,N_14058,N_14946);
and UO_1900 (O_1900,N_14034,N_14778);
xnor UO_1901 (O_1901,N_14505,N_14654);
or UO_1902 (O_1902,N_14466,N_14729);
xnor UO_1903 (O_1903,N_14919,N_13966);
or UO_1904 (O_1904,N_14184,N_14480);
and UO_1905 (O_1905,N_14275,N_14167);
and UO_1906 (O_1906,N_14166,N_14801);
or UO_1907 (O_1907,N_14322,N_14424);
nand UO_1908 (O_1908,N_14856,N_14434);
nor UO_1909 (O_1909,N_13579,N_13855);
or UO_1910 (O_1910,N_13619,N_14796);
nand UO_1911 (O_1911,N_13903,N_13767);
xor UO_1912 (O_1912,N_14566,N_14950);
nor UO_1913 (O_1913,N_13513,N_14921);
nand UO_1914 (O_1914,N_14686,N_13517);
or UO_1915 (O_1915,N_14773,N_14251);
nor UO_1916 (O_1916,N_13603,N_14850);
nor UO_1917 (O_1917,N_14092,N_13758);
nand UO_1918 (O_1918,N_14756,N_14755);
and UO_1919 (O_1919,N_14231,N_14810);
nor UO_1920 (O_1920,N_14308,N_13810);
nor UO_1921 (O_1921,N_14637,N_13666);
nand UO_1922 (O_1922,N_14985,N_14276);
nand UO_1923 (O_1923,N_14310,N_14336);
or UO_1924 (O_1924,N_13934,N_14021);
nor UO_1925 (O_1925,N_14204,N_13642);
nor UO_1926 (O_1926,N_14372,N_13733);
and UO_1927 (O_1927,N_13983,N_14142);
xnor UO_1928 (O_1928,N_14810,N_14203);
nand UO_1929 (O_1929,N_13581,N_14728);
xor UO_1930 (O_1930,N_14925,N_14994);
nand UO_1931 (O_1931,N_14487,N_14091);
or UO_1932 (O_1932,N_14629,N_14119);
and UO_1933 (O_1933,N_14094,N_14079);
or UO_1934 (O_1934,N_14978,N_13668);
nand UO_1935 (O_1935,N_13687,N_14150);
or UO_1936 (O_1936,N_13963,N_14795);
xor UO_1937 (O_1937,N_13879,N_14866);
or UO_1938 (O_1938,N_14778,N_13897);
or UO_1939 (O_1939,N_13955,N_14616);
or UO_1940 (O_1940,N_13524,N_14293);
or UO_1941 (O_1941,N_14118,N_14965);
or UO_1942 (O_1942,N_14955,N_14986);
and UO_1943 (O_1943,N_14385,N_13675);
nor UO_1944 (O_1944,N_14234,N_14151);
xor UO_1945 (O_1945,N_13659,N_14278);
or UO_1946 (O_1946,N_13665,N_14147);
nand UO_1947 (O_1947,N_14645,N_14365);
or UO_1948 (O_1948,N_14102,N_14313);
and UO_1949 (O_1949,N_13668,N_13923);
nand UO_1950 (O_1950,N_14592,N_14182);
nand UO_1951 (O_1951,N_14842,N_14529);
xor UO_1952 (O_1952,N_14781,N_14320);
nand UO_1953 (O_1953,N_13908,N_14083);
and UO_1954 (O_1954,N_14894,N_14551);
or UO_1955 (O_1955,N_14665,N_14610);
and UO_1956 (O_1956,N_14781,N_14182);
and UO_1957 (O_1957,N_14683,N_13611);
nand UO_1958 (O_1958,N_14567,N_13837);
nand UO_1959 (O_1959,N_13977,N_13513);
and UO_1960 (O_1960,N_14614,N_13649);
or UO_1961 (O_1961,N_14522,N_14291);
xnor UO_1962 (O_1962,N_14609,N_14047);
or UO_1963 (O_1963,N_14724,N_13990);
and UO_1964 (O_1964,N_13829,N_14776);
nor UO_1965 (O_1965,N_13625,N_13947);
nand UO_1966 (O_1966,N_14495,N_13854);
and UO_1967 (O_1967,N_14401,N_14901);
xor UO_1968 (O_1968,N_14189,N_14883);
nand UO_1969 (O_1969,N_14150,N_13974);
nor UO_1970 (O_1970,N_14405,N_14558);
nand UO_1971 (O_1971,N_14848,N_14239);
and UO_1972 (O_1972,N_13962,N_14741);
nor UO_1973 (O_1973,N_14411,N_14173);
or UO_1974 (O_1974,N_14852,N_14833);
or UO_1975 (O_1975,N_14015,N_13915);
nand UO_1976 (O_1976,N_14062,N_13778);
or UO_1977 (O_1977,N_14798,N_13527);
and UO_1978 (O_1978,N_14034,N_14365);
xnor UO_1979 (O_1979,N_13929,N_14628);
nand UO_1980 (O_1980,N_13902,N_14361);
nor UO_1981 (O_1981,N_13880,N_14502);
xnor UO_1982 (O_1982,N_14224,N_13790);
or UO_1983 (O_1983,N_14646,N_13907);
and UO_1984 (O_1984,N_14283,N_13730);
and UO_1985 (O_1985,N_13599,N_14431);
or UO_1986 (O_1986,N_13640,N_13936);
xnor UO_1987 (O_1987,N_14726,N_14833);
xor UO_1988 (O_1988,N_14101,N_13625);
nand UO_1989 (O_1989,N_14187,N_14141);
nand UO_1990 (O_1990,N_14233,N_14935);
and UO_1991 (O_1991,N_14707,N_14232);
and UO_1992 (O_1992,N_14195,N_13721);
xnor UO_1993 (O_1993,N_14780,N_14688);
nand UO_1994 (O_1994,N_14884,N_13825);
nor UO_1995 (O_1995,N_14308,N_14549);
xnor UO_1996 (O_1996,N_14769,N_14880);
or UO_1997 (O_1997,N_14414,N_14030);
xnor UO_1998 (O_1998,N_14296,N_13921);
nor UO_1999 (O_1999,N_14515,N_14887);
endmodule